* SPICE3 file created from MUX2X1.ext - technology: sky130A

.subckt MUX2X1 Y A0 A1 S VDD GND
M1000 Y.t3 a_1327_1050.t5 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VDD.t13 A0.t0 a_661_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t2 a_185_209.t3 a_1327_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_185_209.t2 S.t2 VDD.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_661_1050.t0 A0.t1 VDD.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VDD.t12 A1.t1 a_1327_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_661_1050.t4 S.t3 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_1327_1050.t0 a_185_209.t4 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VDD.t4 a_1327_1050.t6 Y.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 GND a_661_1050.t6 a_1888_101.t0 nshort w=-1.605u l=1.765u
+  ad=1.6781p pd=12.81u as=0p ps=0u
M1010 GND a_185_209.t5 a_1222_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1011 VDD.t9 S.t4 a_661_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VDD.t3 a_661_1050.t5 Y.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1327_1050.t3 A1.t2 VDD.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y a_1327_1050.t7 a_1888_101.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1015 VDD.t6 S.t5 a_185_209.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y.t0 a_661_1050.t7 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 GND S.t1 a_556_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
C0 VDD S 0.20fF
C1 VDD A0 0.07fF
C2 VDD A1 0.07fF
C3 VDD Y 1.36fF
C4 A0 S 0.27fF
R0 S.n2 S.t5 512.525
R1 S.n0 S.t4 480.392
R2 S.n0 S.t3 403.272
R3 S.n2 S.t2 371.139
R4 S.n1 S.t1 230.374
R5 S.n3 S.n2 199.753
R6 S.n3 S.t0 183.881
R7 S.n1 S.n0 151.553
R8 S.n4 S.n1 77.859
R9 S.n4 S.n3 76
R10 S.n4 S 0.046
R11 GND.n26 GND.n24 219.745
R12 GND.n85 GND.n84 219.745
R13 GND.n118 GND.n117 219.745
R14 GND.n26 GND.n25 85.529
R15 GND.n85 GND.n83 85.529
R16 GND.n118 GND.n116 85.529
R17 GND.n14 GND.n13 84.842
R18 GND.n44 GND.n43 84.842
R19 GND.n53 GND.n52 76
R20 GND.n12 GND.n11 76
R21 GND.n17 GND.n16 76
R22 GND.n20 GND.n19 76
R23 GND.n23 GND.n22 76
R24 GND.n30 GND.n29 76
R25 GND.n33 GND.n32 76
R26 GND.n36 GND.n35 76
R27 GND.n39 GND.n38 76
R28 GND.n42 GND.n41 76
R29 GND.n47 GND.n46 76
R30 GND.n50 GND.n49 76
R31 GND.n121 GND.n120 76
R32 GND.n114 GND.n113 76
R33 GND.n111 GND.n110 76
R34 GND.n108 GND.n107 76
R35 GND.n105 GND.n104 76
R36 GND.n102 GND.n101 76
R37 GND.n99 GND.n98 76
R38 GND.n91 GND.n90 76
R39 GND.n88 GND.n87 76
R40 GND.n81 GND.n80 76
R41 GND.n78 GND.n77 76
R42 GND.n70 GND.n69 76
R43 GND.n62 GND.n61 76
R44 GND.n96 GND.n95 63.835
R45 GND.n58 GND.t2 39.412
R46 GND.n74 GND.n73 35.01
R47 GND.n8 GND.n7 34.942
R48 GND.n95 GND.n94 28.421
R49 GND.n95 GND.n93 25.263
R50 GND.n93 GND.n92 24.383
R51 GND.n75 GND.n74 19.735
R52 GND.n67 GND.n66 19.735
R53 GND.n60 GND.n59 19.735
R54 GND.n74 GND.n72 19.017
R55 GND.n58 GND.n57 17.185
R56 GND.n6 GND.n5 14.167
R57 GND.n5 GND.n4 14.167
R58 GND.n29 GND.n27 14.167
R59 GND.n120 GND.n119 14.167
R60 GND.n87 GND.n86 14.167
R61 GND.n61 GND.n54 13.653
R62 GND.n69 GND.n68 13.653
R63 GND.n77 GND.n76 13.653
R64 GND.n80 GND.n79 13.653
R65 GND.n87 GND.n82 13.653
R66 GND.n90 GND.n89 13.653
R67 GND.n98 GND.n97 13.653
R68 GND.n101 GND.n100 13.653
R69 GND.n104 GND.n103 13.653
R70 GND.n107 GND.n106 13.653
R71 GND.n110 GND.n109 13.653
R72 GND.n113 GND.n112 13.653
R73 GND.n120 GND.n115 13.653
R74 GND.n49 GND.n48 13.653
R75 GND.n46 GND.n45 13.653
R76 GND.n41 GND.n40 13.653
R77 GND.n38 GND.n37 13.653
R78 GND.n35 GND.n34 13.653
R79 GND.n32 GND.n31 13.653
R80 GND.n29 GND.n28 13.653
R81 GND.n22 GND.n21 13.653
R82 GND.n19 GND.n18 13.653
R83 GND.n16 GND.n15 13.653
R84 GND.n11 GND.n10 13.653
R85 GND.n4 GND.n3 13.653
R86 GND.n5 GND.n2 13.653
R87 GND.n6 GND.n1 13.653
R88 GND.n72 GND.n71 7.5
R89 GND.n65 GND.n64 7.5
R90 GND.n27 GND.n26 7.312
R91 GND.n86 GND.n85 7.312
R92 GND.n119 GND.n118 7.312
R93 GND.n7 GND.n0 7.083
R94 GND.n7 GND.n6 6.474
R95 GND.n59 GND.n58 6.139
R96 GND.n56 GND.n55 4.551
R97 GND.n16 GND.n14 3.935
R98 GND.n46 GND.n44 3.935
R99 GND.n98 GND.n96 3.935
R100 GND.n77 GND.n75 3.935
R101 GND.n61 GND.n60 3.541
R102 GND.t2 GND.n56 2.238
R103 GND.n64 GND.n63 1.935
R104 GND.n52 GND.n51 0.596
R105 GND.n66 GND.n65 0.358
R106 GND.n30 GND.n23 0.29
R107 GND.n121 GND.n114 0.29
R108 GND.n88 GND.n81 0.29
R109 GND.n53 GND 0.207
R110 GND.n69 GND.n67 0.196
R111 GND.n12 GND.n9 0.181
R112 GND.n42 GND.n39 0.181
R113 GND.n105 GND.n102 0.181
R114 GND.n78 GND.n70 0.157
R115 GND.n70 GND.n62 0.157
R116 GND.n9 GND.n8 0.145
R117 GND.n17 GND.n12 0.145
R118 GND.n20 GND.n17 0.145
R119 GND.n23 GND.n20 0.145
R120 GND.n33 GND.n30 0.145
R121 GND.n36 GND.n33 0.145
R122 GND.n39 GND.n36 0.145
R123 GND.n47 GND.n42 0.145
R124 GND.n50 GND.n47 0.145
R125 GND.n114 GND.n111 0.145
R126 GND.n111 GND.n108 0.145
R127 GND.n108 GND.n105 0.145
R128 GND.n102 GND.n99 0.145
R129 GND.n99 GND.n91 0.145
R130 GND.n91 GND.n88 0.145
R131 GND.n81 GND.n78 0.145
R132 GND.n62 GND.n53 0.145
R133 GND GND.n121 0.078
R134 GND GND.n50 0.066
R135 a_185_209.n1 a_185_209.t3 480.392
R136 a_185_209.n1 a_185_209.t4 403.272
R137 a_185_209.n2 a_185_209.t5 256.927
R138 a_185_209.n5 a_185_209.n3 185.537
R139 a_185_209.n3 a_185_209.n0 184.007
R140 a_185_209.n3 a_185_209.n2 155.763
R141 a_185_209.n2 a_185_209.n1 125
R142 a_185_209.n5 a_185_209.n4 15.218
R143 a_185_209.n0 a_185_209.t1 14.282
R144 a_185_209.n0 a_185_209.t2 14.282
R145 a_185_209.n6 a_185_209.n5 12.014
R146 a_556_101.n12 a_556_101.n11 26.811
R147 a_556_101.n6 a_556_101.n5 24.977
R148 a_556_101.n2 a_556_101.n1 24.877
R149 a_556_101.t0 a_556_101.n2 12.677
R150 a_556_101.t0 a_556_101.n3 11.595
R151 a_556_101.t1 a_556_101.n8 8.137
R152 a_556_101.t0 a_556_101.n4 7.273
R153 a_556_101.t0 a_556_101.n0 6.109
R154 a_556_101.t1 a_556_101.n7 4.864
R155 a_556_101.t0 a_556_101.n12 2.074
R156 a_556_101.n7 a_556_101.n6 1.13
R157 a_556_101.n12 a_556_101.t1 0.937
R158 a_556_101.t1 a_556_101.n10 0.804
R159 a_556_101.n10 a_556_101.n9 0.136
R160 a_1327_1050.n3 a_1327_1050.t6 472.359
R161 a_1327_1050.n3 a_1327_1050.t5 384.527
R162 a_1327_1050.n4 a_1327_1050.t7 214.619
R163 a_1327_1050.n7 a_1327_1050.n5 190.561
R164 a_1327_1050.n5 a_1327_1050.n2 179.052
R165 a_1327_1050.n5 a_1327_1050.n4 153.859
R166 a_1327_1050.n4 a_1327_1050.n3 136.613
R167 a_1327_1050.n2 a_1327_1050.n1 76.002
R168 a_1327_1050.n7 a_1327_1050.n6 15.218
R169 a_1327_1050.n0 a_1327_1050.t4 14.282
R170 a_1327_1050.n0 a_1327_1050.t3 14.282
R171 a_1327_1050.n1 a_1327_1050.t1 14.282
R172 a_1327_1050.n1 a_1327_1050.t0 14.282
R173 a_1327_1050.n2 a_1327_1050.n0 12.85
R174 a_1327_1050.n8 a_1327_1050.n7 12.014
R175 VDD.n162 VDD.n160 144.705
R176 VDD.n83 VDD.n81 144.705
R177 VDD.n224 VDD.n222 144.705
R178 VDD.n152 VDD.n151 77.792
R179 VDD.n141 VDD.n140 77.792
R180 VDD.n44 VDD.n43 76
R181 VDD.n49 VDD.n48 76
R182 VDD.n54 VDD.n53 76
R183 VDD.n58 VDD.n57 76
R184 VDD.n85 VDD.n84 76
R185 VDD.n90 VDD.n89 76
R186 VDD.n95 VDD.n94 76
R187 VDD.n101 VDD.n100 76
R188 VDD.n106 VDD.n105 76
R189 VDD.n111 VDD.n110 76
R190 VDD.n116 VDD.n115 76
R191 VDD.n247 VDD.n246 76
R192 VDD.n221 VDD.n220 76
R193 VDD.n217 VDD.n216 76
R194 VDD.n212 VDD.n211 76
R195 VDD.n207 VDD.n206 76
R196 VDD.n201 VDD.n200 76
R197 VDD.n196 VDD.n195 76
R198 VDD.n191 VDD.n190 76
R199 VDD.n186 VDD.n185 76
R200 VDD.n159 VDD.n158 76
R201 VDD.n155 VDD.n154 76
R202 VDD.n149 VDD.n148 76
R203 VDD.n145 VDD.n144 76
R204 VDD.n139 VDD.n138 76
R205 VDD.n143 VDD.t7 55.106
R206 VDD.n150 VDD.t6 55.106
R207 VDD.n187 VDD.t8 55.106
R208 VDD.n112 VDD.t1 55.106
R209 VDD.n50 VDD.t0 55.106
R210 VDD.n215 VDD.t13 55.106
R211 VDD.n88 VDD.t12 55.106
R212 VDD.n35 VDD.t4 55.106
R213 VDD.n205 VDD.n204 40.824
R214 VDD.n99 VDD.n98 40.824
R215 VDD.n29 VDD.n28 40.824
R216 VDD.n229 VDD.n228 36.774
R217 VDD.n63 VDD.n62 36.774
R218 VDD.n178 VDD.n177 36.774
R219 VDD.n32 VDD.n31 36.608
R220 VDD.n92 VDD.n91 36.608
R221 VDD.n209 VDD.n208 36.608
R222 VDD.n38 VDD.n37 34.942
R223 VDD.n46 VDD.n45 32.032
R224 VDD.n108 VDD.n107 32.032
R225 VDD.n193 VDD.n192 32.032
R226 VDD.n138 VDD.n135 21.841
R227 VDD.n23 VDD.n20 21.841
R228 VDD.n204 VDD.t10 14.282
R229 VDD.n204 VDD.t9 14.282
R230 VDD.n98 VDD.t11 14.282
R231 VDD.n98 VDD.t2 14.282
R232 VDD.n28 VDD.t5 14.282
R233 VDD.n28 VDD.t3 14.282
R234 VDD.n135 VDD.n118 14.167
R235 VDD.n118 VDD.n117 14.167
R236 VDD.n244 VDD.n226 14.167
R237 VDD.n226 VDD.n225 14.167
R238 VDD.n79 VDD.n60 14.167
R239 VDD.n60 VDD.n59 14.167
R240 VDD.n183 VDD.n164 14.167
R241 VDD.n164 VDD.n163 14.167
R242 VDD.n20 VDD.n19 14.167
R243 VDD.n19 VDD.n17 14.167
R244 VDD.n34 VDD.n30 14.167
R245 VDD.n84 VDD.n80 14.167
R246 VDD.n246 VDD.n245 14.167
R247 VDD.n185 VDD.n184 14.167
R248 VDD.n23 VDD.n22 13.653
R249 VDD.n22 VDD.n21 13.653
R250 VDD.n36 VDD.n25 13.653
R251 VDD.n25 VDD.n24 13.653
R252 VDD.n34 VDD.n33 13.653
R253 VDD.n33 VDD.n32 13.653
R254 VDD.n30 VDD.n27 13.653
R255 VDD.n27 VDD.n26 13.653
R256 VDD.n43 VDD.n42 13.653
R257 VDD.n42 VDD.n41 13.653
R258 VDD.n48 VDD.n47 13.653
R259 VDD.n47 VDD.n46 13.653
R260 VDD.n53 VDD.n52 13.653
R261 VDD.n52 VDD.n51 13.653
R262 VDD.n57 VDD.n56 13.653
R263 VDD.n56 VDD.n55 13.653
R264 VDD.n84 VDD.n83 13.653
R265 VDD.n83 VDD.n82 13.653
R266 VDD.n89 VDD.n87 13.653
R267 VDD.n87 VDD.n86 13.653
R268 VDD.n94 VDD.n93 13.653
R269 VDD.n93 VDD.n92 13.653
R270 VDD.n100 VDD.n97 13.653
R271 VDD.n97 VDD.n96 13.653
R272 VDD.n105 VDD.n104 13.653
R273 VDD.n104 VDD.n103 13.653
R274 VDD.n110 VDD.n109 13.653
R275 VDD.n109 VDD.n108 13.653
R276 VDD.n115 VDD.n114 13.653
R277 VDD.n114 VDD.n113 13.653
R278 VDD.n246 VDD.n224 13.653
R279 VDD.n224 VDD.n223 13.653
R280 VDD.n220 VDD.n219 13.653
R281 VDD.n219 VDD.n218 13.653
R282 VDD.n216 VDD.n214 13.653
R283 VDD.n214 VDD.n213 13.653
R284 VDD.n211 VDD.n210 13.653
R285 VDD.n210 VDD.n209 13.653
R286 VDD.n206 VDD.n203 13.653
R287 VDD.n203 VDD.n202 13.653
R288 VDD.n200 VDD.n199 13.653
R289 VDD.n199 VDD.n198 13.653
R290 VDD.n195 VDD.n194 13.653
R291 VDD.n194 VDD.n193 13.653
R292 VDD.n190 VDD.n189 13.653
R293 VDD.n189 VDD.n188 13.653
R294 VDD.n185 VDD.n162 13.653
R295 VDD.n162 VDD.n161 13.653
R296 VDD.n158 VDD.n157 13.653
R297 VDD.n157 VDD.n156 13.653
R298 VDD.n154 VDD.n153 13.653
R299 VDD.n153 VDD.n152 13.653
R300 VDD.n148 VDD.n147 13.653
R301 VDD.n147 VDD.n146 13.653
R302 VDD.n144 VDD.n142 13.653
R303 VDD.n142 VDD.n141 13.653
R304 VDD.n138 VDD.n137 13.653
R305 VDD.n137 VDD.n136 13.653
R306 VDD.n4 VDD.n2 12.915
R307 VDD.n4 VDD.n3 12.66
R308 VDD.n12 VDD.n11 12.343
R309 VDD.n8 VDD.n7 12.343
R310 VDD.n12 VDD.n9 12.343
R311 VDD.n35 VDD.n34 11.806
R312 VDD.n30 VDD.n29 8.658
R313 VDD.n100 VDD.n99 8.658
R314 VDD.n206 VDD.n205 8.658
R315 VDD.n245 VDD.n244 7.674
R316 VDD.n80 VDD.n79 7.674
R317 VDD.n184 VDD.n183 7.674
R318 VDD.n74 VDD.n73 7.5
R319 VDD.n68 VDD.n67 7.5
R320 VDD.n70 VDD.n69 7.5
R321 VDD.n65 VDD.n64 7.5
R322 VDD.n79 VDD.n78 7.5
R323 VDD.n239 VDD.n238 7.5
R324 VDD.n233 VDD.n232 7.5
R325 VDD.n235 VDD.n234 7.5
R326 VDD.n241 VDD.n231 7.5
R327 VDD.n241 VDD.n229 7.5
R328 VDD.n244 VDD.n243 7.5
R329 VDD.n168 VDD.n167 7.5
R330 VDD.n171 VDD.n170 7.5
R331 VDD.n173 VDD.n172 7.5
R332 VDD.n176 VDD.n175 7.5
R333 VDD.n183 VDD.n182 7.5
R334 VDD.n130 VDD.n129 7.5
R335 VDD.n124 VDD.n123 7.5
R336 VDD.n126 VDD.n125 7.5
R337 VDD.n132 VDD.n122 7.5
R338 VDD.n132 VDD.n120 7.5
R339 VDD.n135 VDD.n134 7.5
R340 VDD.n20 VDD.n16 7.5
R341 VDD.n2 VDD.n1 7.5
R342 VDD.n7 VDD.n6 7.5
R343 VDD.n11 VDD.n10 7.5
R344 VDD.n19 VDD.n18 7.5
R345 VDD.n14 VDD.n0 7.5
R346 VDD.n66 VDD.n63 6.772
R347 VDD.n77 VDD.n61 6.772
R348 VDD.n75 VDD.n72 6.772
R349 VDD.n71 VDD.n68 6.772
R350 VDD.n242 VDD.n227 6.772
R351 VDD.n240 VDD.n237 6.772
R352 VDD.n236 VDD.n233 6.772
R353 VDD.n133 VDD.n119 6.772
R354 VDD.n131 VDD.n128 6.772
R355 VDD.n127 VDD.n124 6.772
R356 VDD.n66 VDD.n65 6.772
R357 VDD.n71 VDD.n70 6.772
R358 VDD.n75 VDD.n74 6.772
R359 VDD.n78 VDD.n77 6.772
R360 VDD.n236 VDD.n235 6.772
R361 VDD.n240 VDD.n239 6.772
R362 VDD.n243 VDD.n242 6.772
R363 VDD.n127 VDD.n126 6.772
R364 VDD.n131 VDD.n130 6.772
R365 VDD.n134 VDD.n133 6.772
R366 VDD.n182 VDD.n181 6.772
R367 VDD.n169 VDD.n166 6.772
R368 VDD.n174 VDD.n171 6.772
R369 VDD.n179 VDD.n176 6.772
R370 VDD.n179 VDD.n178 6.772
R371 VDD.n174 VDD.n173 6.772
R372 VDD.n169 VDD.n168 6.772
R373 VDD.n181 VDD.n165 6.772
R374 VDD.n37 VDD.n23 6.487
R375 VDD.n37 VDD.n36 6.475
R376 VDD.n16 VDD.n15 6.458
R377 VDD.n231 VDD.n230 6.202
R378 VDD.n122 VDD.n121 6.202
R379 VDD.n41 VDD.n40 4.576
R380 VDD.n103 VDD.n102 4.576
R381 VDD.n198 VDD.n197 4.576
R382 VDD.n53 VDD.n50 2.754
R383 VDD.n115 VDD.n112 2.754
R384 VDD.n190 VDD.n187 2.754
R385 VDD.n36 VDD.n35 2.361
R386 VDD.n89 VDD.n88 2.361
R387 VDD.n216 VDD.n215 2.361
R388 VDD.n154 VDD.n150 1.967
R389 VDD.n144 VDD.n143 1.967
R390 VDD.n14 VDD.n5 1.329
R391 VDD.n14 VDD.n8 1.329
R392 VDD.n14 VDD.n12 1.329
R393 VDD.n14 VDD.n13 1.329
R394 VDD.n15 VDD.n14 0.696
R395 VDD.n14 VDD.n4 0.696
R396 VDD.n76 VDD.n75 0.365
R397 VDD.n76 VDD.n71 0.365
R398 VDD.n76 VDD.n66 0.365
R399 VDD.n77 VDD.n76 0.365
R400 VDD.n241 VDD.n240 0.365
R401 VDD.n241 VDD.n236 0.365
R402 VDD.n242 VDD.n241 0.365
R403 VDD.n132 VDD.n131 0.365
R404 VDD.n132 VDD.n127 0.365
R405 VDD.n133 VDD.n132 0.365
R406 VDD.n180 VDD.n179 0.365
R407 VDD.n180 VDD.n174 0.365
R408 VDD.n180 VDD.n169 0.365
R409 VDD.n181 VDD.n180 0.365
R410 VDD.n85 VDD.n58 0.29
R411 VDD.n247 VDD.n221 0.29
R412 VDD.n186 VDD.n159 0.29
R413 VDD.n139 VDD 0.207
R414 VDD.n44 VDD.n39 0.181
R415 VDD.n106 VDD.n101 0.181
R416 VDD.n207 VDD.n201 0.181
R417 VDD.n155 VDD.n149 0.157
R418 VDD.n149 VDD.n145 0.157
R419 VDD.n39 VDD.n38 0.145
R420 VDD.n49 VDD.n44 0.145
R421 VDD.n54 VDD.n49 0.145
R422 VDD.n58 VDD.n54 0.145
R423 VDD.n90 VDD.n85 0.145
R424 VDD.n95 VDD.n90 0.145
R425 VDD.n101 VDD.n95 0.145
R426 VDD.n111 VDD.n106 0.145
R427 VDD.n116 VDD.n111 0.145
R428 VDD.n221 VDD.n217 0.145
R429 VDD.n217 VDD.n212 0.145
R430 VDD.n212 VDD.n207 0.145
R431 VDD.n201 VDD.n196 0.145
R432 VDD.n196 VDD.n191 0.145
R433 VDD.n191 VDD.n186 0.145
R434 VDD.n159 VDD.n155 0.145
R435 VDD.n145 VDD.n139 0.145
R436 VDD VDD.n247 0.078
R437 VDD VDD.n116 0.066
R438 Y.n7 Y.n6 184.039
R439 Y.n7 Y.n2 179.052
R440 Y.n2 Y.n1 76.002
R441 Y.n8 Y.n7 76
R442 Y.n6 Y.n5 30
R443 Y.n4 Y.n3 24.383
R444 Y.n6 Y.n4 23.684
R445 Y.n0 Y.t2 14.282
R446 Y.n0 Y.t3 14.282
R447 Y.n1 Y.t1 14.282
R448 Y.n1 Y.t0 14.282
R449 Y.n2 Y.n0 12.85
R450 Y.n8 Y 0.046
R451 A0.n0 A0.t0 472.359
R452 A0.n0 A0.t1 384.527
R453 A0.n1 A0.t2 241.172
R454 A0.n1 A0.n0 110.06
R455 A0.n2 A0.n1 76
R456 A0.n2 A0 0.046
R457 a_661_1050.n0 a_661_1050.t5 480.392
R458 a_661_1050.n0 a_661_1050.t7 403.272
R459 a_661_1050.n1 a_661_1050.t6 230.374
R460 a_661_1050.n5 a_661_1050.n3 205.605
R461 a_661_1050.n3 a_661_1050.n2 179.225
R462 a_661_1050.n3 a_661_1050.n1 155.763
R463 a_661_1050.n1 a_661_1050.n0 151.553
R464 a_661_1050.n5 a_661_1050.n4 76.002
R465 a_661_1050.n4 a_661_1050.t3 14.282
R466 a_661_1050.n4 a_661_1050.t4 14.282
R467 a_661_1050.t1 a_661_1050.n6 14.282
R468 a_661_1050.n6 a_661_1050.t0 14.282
R469 a_661_1050.n6 a_661_1050.n5 12.848
R470 A1.n0 A1.t1 472.359
R471 A1.n0 A1.t2 384.527
R472 A1.n1 A1.t0 267.725
R473 A1.n1 A1.n0 83.507
R474 A1.n2 A1.n1 76
R475 A1.n2 A1 0.046
R476 a_1222_101.n12 a_1222_101.n11 26.811
R477 a_1222_101.n6 a_1222_101.n5 24.977
R478 a_1222_101.n2 a_1222_101.n1 24.877
R479 a_1222_101.t0 a_1222_101.n2 12.677
R480 a_1222_101.t0 a_1222_101.n3 11.595
R481 a_1222_101.t1 a_1222_101.n8 8.137
R482 a_1222_101.t0 a_1222_101.n4 7.273
R483 a_1222_101.t0 a_1222_101.n0 6.109
R484 a_1222_101.t1 a_1222_101.n7 4.864
R485 a_1222_101.t0 a_1222_101.n12 2.074
R486 a_1222_101.n7 a_1222_101.n6 1.13
R487 a_1222_101.n12 a_1222_101.t1 0.937
R488 a_1222_101.t1 a_1222_101.n10 0.804
R489 a_1222_101.n10 a_1222_101.n9 0.136
R490 a_1888_101.n12 a_1888_101.n11 26.811
R491 a_1888_101.n6 a_1888_101.n5 24.977
R492 a_1888_101.n2 a_1888_101.n1 24.877
R493 a_1888_101.t0 a_1888_101.n2 12.677
R494 a_1888_101.t0 a_1888_101.n3 11.595
R495 a_1888_101.t1 a_1888_101.n8 8.137
R496 a_1888_101.t0 a_1888_101.n4 7.273
R497 a_1888_101.t0 a_1888_101.n0 6.109
R498 a_1888_101.t1 a_1888_101.n7 4.864
R499 a_1888_101.t0 a_1888_101.n12 2.074
R500 a_1888_101.n7 a_1888_101.n6 1.13
R501 a_1888_101.n12 a_1888_101.t1 0.937
R502 a_1888_101.t1 a_1888_101.n10 0.804
R503 a_1888_101.n10 a_1888_101.n9 0.136
C5 S GND 1.50fF
C6 VDD GND 9.87fF
C7 a_1888_101.n0 GND 0.02fF
C8 a_1888_101.n1 GND 0.10fF
C9 a_1888_101.n2 GND 0.06fF
C10 a_1888_101.n3 GND 0.06fF
C11 a_1888_101.n4 GND 0.00fF
C12 a_1888_101.n5 GND 0.04fF
C13 a_1888_101.n6 GND 0.05fF
C14 a_1888_101.n7 GND 0.02fF
C15 a_1888_101.n8 GND 0.05fF
C16 a_1888_101.n9 GND 0.07fF
C17 a_1888_101.n10 GND 0.17fF
C18 a_1888_101.n11 GND 0.09fF
C19 a_1888_101.n12 GND 0.00fF
C20 a_1222_101.n0 GND 0.02fF
C21 a_1222_101.n1 GND 0.10fF
C22 a_1222_101.n2 GND 0.06fF
C23 a_1222_101.n3 GND 0.06fF
C24 a_1222_101.n4 GND 0.00fF
C25 a_1222_101.n5 GND 0.04fF
C26 a_1222_101.n6 GND 0.05fF
C27 a_1222_101.n7 GND 0.02fF
C28 a_1222_101.n8 GND 0.05fF
C29 a_1222_101.n9 GND 0.08fF
C30 a_1222_101.n10 GND 0.17fF
C31 a_1222_101.t1 GND 0.23fF
C32 a_1222_101.n11 GND 0.09fF
C33 a_1222_101.n12 GND 0.00fF
C34 a_661_1050.n0 GND 0.43fF
C35 a_661_1050.n1 GND 0.82fF
C36 a_661_1050.n2 GND 0.33fF
C37 a_661_1050.n3 GND 0.90fF
C38 a_661_1050.n4 GND 0.62fF
C39 a_661_1050.n5 GND 0.36fF
C40 a_661_1050.n6 GND 0.53fF
C41 Y.n0 GND 0.48fF
C42 Y.n1 GND 0.57fF
C43 Y.n2 GND 0.31fF
C44 Y.n3 GND 0.04fF
C45 Y.n4 GND 0.05fF
C46 Y.n5 GND 0.03fF
C47 Y.n6 GND 0.24fF
C48 Y.n7 GND 0.39fF
C49 Y.n8 GND 0.01fF
C50 VDD.n0 GND 0.14fF
C51 VDD.n1 GND 0.02fF
C52 VDD.n2 GND 0.02fF
C53 VDD.n3 GND 0.04fF
C54 VDD.n4 GND 0.01fF
C55 VDD.n6 GND 0.02fF
C56 VDD.n7 GND 0.02fF
C57 VDD.n9 GND 0.02fF
C58 VDD.n10 GND 0.02fF
C59 VDD.n11 GND 0.02fF
C60 VDD.n14 GND 0.42fF
C61 VDD.n16 GND 0.03fF
C62 VDD.n17 GND 0.02fF
C63 VDD.n18 GND 0.02fF
C64 VDD.n19 GND 0.02fF
C65 VDD.n20 GND 0.03fF
C66 VDD.n21 GND 0.25fF
C67 VDD.n22 GND 0.02fF
C68 VDD.n23 GND 0.03fF
C69 VDD.n24 GND 0.22fF
C70 VDD.n25 GND 0.01fF
C71 VDD.n26 GND 0.28fF
C72 VDD.n27 GND 0.01fF
C73 VDD.n28 GND 0.10fF
C74 VDD.n29 GND 0.02fF
C75 VDD.n30 GND 0.02fF
C76 VDD.n31 GND 0.13fF
C77 VDD.n32 GND 0.15fF
C78 VDD.n33 GND 0.01fF
C79 VDD.n34 GND 0.02fF
C80 VDD.n35 GND 0.05fF
C81 VDD.n36 GND 0.01fF
C82 VDD.n37 GND 0.00fF
C83 VDD.n38 GND 0.08fF
C84 VDD.n39 GND 0.02fF
C85 VDD.n40 GND 0.16fF
C86 VDD.n41 GND 0.13fF
C87 VDD.n42 GND 0.01fF
C88 VDD.n43 GND 0.02fF
C89 VDD.n44 GND 0.02fF
C90 VDD.n45 GND 0.13fF
C91 VDD.n46 GND 0.15fF
C92 VDD.n47 GND 0.01fF
C93 VDD.n48 GND 0.02fF
C94 VDD.n49 GND 0.02fF
C95 VDD.n50 GND 0.06fF
C96 VDD.n51 GND 0.23fF
C97 VDD.n52 GND 0.01fF
C98 VDD.n53 GND 0.01fF
C99 VDD.n54 GND 0.02fF
C100 VDD.n55 GND 0.25fF
C101 VDD.n56 GND 0.01fF
C102 VDD.n57 GND 0.02fF
C103 VDD.n58 GND 0.03fF
C104 VDD.n59 GND 0.02fF
C105 VDD.n60 GND 0.02fF
C106 VDD.n61 GND 0.02fF
C107 VDD.n62 GND 0.20fF
C108 VDD.n63 GND 0.04fF
C109 VDD.n64 GND 0.03fF
C110 VDD.n65 GND 0.02fF
C111 VDD.n67 GND 0.02fF
C112 VDD.n68 GND 0.02fF
C113 VDD.n69 GND 0.02fF
C114 VDD.n70 GND 0.02fF
C115 VDD.n72 GND 0.02fF
C116 VDD.n73 GND 0.02fF
C117 VDD.n74 GND 0.02fF
C118 VDD.n76 GND 0.25fF
C119 VDD.n78 GND 0.02fF
C120 VDD.n79 GND 0.02fF
C121 VDD.n80 GND 0.03fF
C122 VDD.n81 GND 0.02fF
C123 VDD.n82 GND 0.25fF
C124 VDD.n83 GND 0.01fF
C125 VDD.n84 GND 0.02fF
C126 VDD.n85 GND 0.03fF
C127 VDD.n86 GND 0.22fF
C128 VDD.n87 GND 0.01fF
C129 VDD.n88 GND 0.05fF
C130 VDD.n89 GND 0.01fF
C131 VDD.n90 GND 0.02fF
C132 VDD.n91 GND 0.13fF
C133 VDD.n92 GND 0.15fF
C134 VDD.n93 GND 0.01fF
C135 VDD.n94 GND 0.02fF
C136 VDD.n95 GND 0.02fF
C137 VDD.n96 GND 0.28fF
C138 VDD.n97 GND 0.01fF
C139 VDD.n98 GND 0.10fF
C140 VDD.n99 GND 0.02fF
C141 VDD.n100 GND 0.02fF
C142 VDD.n101 GND 0.02fF
C143 VDD.n102 GND 0.16fF
C144 VDD.n103 GND 0.13fF
C145 VDD.n104 GND 0.01fF
C146 VDD.n105 GND 0.02fF
C147 VDD.n106 GND 0.02fF
C148 VDD.n107 GND 0.13fF
C149 VDD.n108 GND 0.15fF
C150 VDD.n109 GND 0.01fF
C151 VDD.n110 GND 0.02fF
C152 VDD.n111 GND 0.02fF
C153 VDD.n112 GND 0.06fF
C154 VDD.n113 GND 0.23fF
C155 VDD.n114 GND 0.01fF
C156 VDD.n115 GND 0.01fF
C157 VDD.n116 GND 0.02fF
C158 VDD.n117 GND 0.02fF
C159 VDD.n118 GND 0.02fF
C160 VDD.n119 GND 0.02fF
C161 VDD.n120 GND 0.11fF
C162 VDD.n121 GND 0.03fF
C163 VDD.n122 GND 0.02fF
C164 VDD.n123 GND 0.02fF
C165 VDD.n124 GND 0.02fF
C166 VDD.n125 GND 0.02fF
C167 VDD.n126 GND 0.02fF
C168 VDD.n128 GND 0.02fF
C169 VDD.n129 GND 0.02fF
C170 VDD.n130 GND 0.02fF
C171 VDD.n132 GND 0.42fF
C172 VDD.n134 GND 0.03fF
C173 VDD.n135 GND 0.03fF
C174 VDD.n136 GND 0.25fF
C175 VDD.n137 GND 0.02fF
C176 VDD.n138 GND 0.03fF
C177 VDD.n139 GND 0.03fF
C178 VDD.n140 GND 0.14fF
C179 VDD.n141 GND 0.19fF
C180 VDD.n142 GND 0.01fF
C181 VDD.n143 GND 0.06fF
C182 VDD.n144 GND 0.01fF
C183 VDD.n145 GND 0.02fF
C184 VDD.n146 GND 0.15fF
C185 VDD.n147 GND 0.01fF
C186 VDD.n148 GND 0.02fF
C187 VDD.n149 GND 0.02fF
C188 VDD.n150 GND 0.05fF
C189 VDD.n151 GND 0.14fF
C190 VDD.n152 GND 0.19fF
C191 VDD.n153 GND 0.01fF
C192 VDD.n154 GND 0.01fF
C193 VDD.n155 GND 0.02fF
C194 VDD.n156 GND 0.25fF
C195 VDD.n157 GND 0.01fF
C196 VDD.n158 GND 0.02fF
C197 VDD.n159 GND 0.03fF
C198 VDD.n160 GND 0.02fF
C199 VDD.n161 GND 0.25fF
C200 VDD.n162 GND 0.01fF
C201 VDD.n163 GND 0.02fF
C202 VDD.n164 GND 0.02fF
C203 VDD.n165 GND 0.02fF
C204 VDD.n166 GND 0.02fF
C205 VDD.n167 GND 0.02fF
C206 VDD.n168 GND 0.02fF
C207 VDD.n170 GND 0.02fF
C208 VDD.n171 GND 0.02fF
C209 VDD.n172 GND 0.02fF
C210 VDD.n173 GND 0.02fF
C211 VDD.n175 GND 0.03fF
C212 VDD.n176 GND 0.02fF
C213 VDD.n177 GND 0.17fF
C214 VDD.n178 GND 0.04fF
C215 VDD.n180 GND 0.25fF
C216 VDD.n182 GND 0.02fF
C217 VDD.n183 GND 0.02fF
C218 VDD.n184 GND 0.03fF
C219 VDD.n185 GND 0.02fF
C220 VDD.n186 GND 0.03fF
C221 VDD.n187 GND 0.06fF
C222 VDD.n188 GND 0.23fF
C223 VDD.n189 GND 0.01fF
C224 VDD.n190 GND 0.01fF
C225 VDD.n191 GND 0.02fF
C226 VDD.n192 GND 0.13fF
C227 VDD.n193 GND 0.15fF
C228 VDD.n194 GND 0.01fF
C229 VDD.n195 GND 0.02fF
C230 VDD.n196 GND 0.02fF
C231 VDD.n197 GND 0.16fF
C232 VDD.n198 GND 0.13fF
C233 VDD.n199 GND 0.01fF
C234 VDD.n200 GND 0.02fF
C235 VDD.n201 GND 0.02fF
C236 VDD.n202 GND 0.28fF
C237 VDD.n203 GND 0.01fF
C238 VDD.n204 GND 0.10fF
C239 VDD.n205 GND 0.02fF
C240 VDD.n206 GND 0.02fF
C241 VDD.n207 GND 0.02fF
C242 VDD.n208 GND 0.13fF
C243 VDD.n209 GND 0.15fF
C244 VDD.n210 GND 0.01fF
C245 VDD.n211 GND 0.02fF
C246 VDD.n212 GND 0.02fF
C247 VDD.n213 GND 0.22fF
C248 VDD.n214 GND 0.01fF
C249 VDD.n215 GND 0.05fF
C250 VDD.n216 GND 0.01fF
C251 VDD.n217 GND 0.02fF
C252 VDD.n218 GND 0.25fF
C253 VDD.n219 GND 0.01fF
C254 VDD.n220 GND 0.02fF
C255 VDD.n221 GND 0.03fF
C256 VDD.n222 GND 0.02fF
C257 VDD.n223 GND 0.25fF
C258 VDD.n224 GND 0.01fF
C259 VDD.n225 GND 0.02fF
C260 VDD.n226 GND 0.02fF
C261 VDD.n227 GND 0.02fF
C262 VDD.n228 GND 0.20fF
C263 VDD.n229 GND 0.04fF
C264 VDD.n230 GND 0.03fF
C265 VDD.n231 GND 0.02fF
C266 VDD.n232 GND 0.02fF
C267 VDD.n233 GND 0.02fF
C268 VDD.n234 GND 0.02fF
C269 VDD.n235 GND 0.02fF
C270 VDD.n237 GND 0.02fF
C271 VDD.n238 GND 0.02fF
C272 VDD.n239 GND 0.02fF
C273 VDD.n241 GND 0.25fF
C274 VDD.n243 GND 0.02fF
C275 VDD.n244 GND 0.02fF
C276 VDD.n245 GND 0.03fF
C277 VDD.n246 GND 0.02fF
C278 VDD.n247 GND 0.03fF
C279 a_1327_1050.n0 GND 0.49fF
C280 a_1327_1050.n1 GND 0.58fF
C281 a_1327_1050.n2 GND 0.31fF
C282 a_1327_1050.n3 GND 0.34fF
C283 a_1327_1050.n4 GND 0.57fF
C284 a_1327_1050.n5 GND 0.62fF
C285 a_1327_1050.n6 GND 0.08fF
C286 a_1327_1050.n7 GND 0.24fF
C287 a_1327_1050.n8 GND 0.04fF
C288 a_556_101.n0 GND 0.02fF
C289 a_556_101.n1 GND 0.10fF
C290 a_556_101.n2 GND 0.06fF
C291 a_556_101.n3 GND 0.06fF
C292 a_556_101.n4 GND 0.00fF
C293 a_556_101.n5 GND 0.04fF
C294 a_556_101.n6 GND 0.05fF
C295 a_556_101.n7 GND 0.02fF
C296 a_556_101.n8 GND 0.05fF
C297 a_556_101.n9 GND 0.08fF
C298 a_556_101.n10 GND 0.18fF
C299 a_556_101.t1 GND 0.24fF
C300 a_556_101.n11 GND 0.09fF
C301 a_556_101.n12 GND 0.00fF
C302 a_185_209.n0 GND 0.82fF
C303 a_185_209.n1 GND 0.44fF
C304 a_185_209.n2 GND 0.91fF
C305 a_185_209.n3 GND 0.97fF
C306 a_185_209.n4 GND 0.09fF
C307 a_185_209.n5 GND 0.27fF
C308 a_185_209.n6 GND 0.05fF
C309 S.n0 GND 0.33fF
C310 S.n1 GND 0.30fF
C311 S.n2 GND 0.31fF
C312 S.t0 GND 0.37fF
C313 S.n3 GND 0.33fF
C314 S.n4 GND 0.35fF
.ends
