// File: DLATCHN.spi.pex
// Created: Tue Oct 15 15:48:39 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_DLATCHN\%GND ( 1 38 50 54 62 68 76 80 83 88 92 100 108 111 116 120 \
 123 128 134 140 146 151 156 160 180 184 192 196 204 210 218 222 230 234 245 \
 248 259 271 273 285 288 300 320 340 341 342 343 344 345 346 347 )
c307 ( 347 0 ) capacitor c=0.0706776f //x=19.43 //y=0.365
c308 ( 346 0 ) capacitor c=0.0706539f //x=16.1 //y=0.365
c309 ( 345 0 ) capacitor c=0.0578714f //x=13.815 //y=0.37
c310 ( 344 0 ) capacitor c=0.0207878f //x=10.98 //y=0.865
c311 ( 343 0 ) capacitor c=0.0572693f //x=8.265 //y=0.37
c312 ( 342 0 ) capacitor c=0.0207873f //x=5.43 //y=0.865
c313 ( 341 0 ) capacitor c=0.0572693f //x=2.715 //y=0.37
c314 ( 340 0 ) capacitor c=0.0589324f //x=0.495 //y=0.37
c315 ( 320 0 ) capacitor c=0.10534f //x=18.87 //y=0
c316 ( 300 0 ) capacitor c=0.103812f //x=15.54 //y=0
c317 ( 288 0 ) capacitor c=0.10149f //x=13.32 //y=0
c318 ( 287 0 ) capacitor c=0.00440095f //x=11.1 //y=0
c319 ( 285 0 ) capacitor c=0.102231f //x=9.99 //y=0
c320 ( 273 0 ) capacitor c=0.10097f //x=7.77 //y=0
c321 ( 272 0 ) capacitor c=0.00440095f //x=5.62 //y=0
c322 ( 271 0 ) capacitor c=0.102231f //x=4.44 //y=0
c323 ( 259 0 ) capacitor c=0.0966579f //x=2.22 //y=0
c324 ( 248 0 ) capacitor c=0.192978f //x=0.63 //y=0
c325 ( 245 0 ) capacitor c=0.204536f //x=21.83 //y=0
c326 ( 243 0 ) capacitor c=0.0659517f //x=21.59 //y=0
c327 ( 237 0 ) capacitor c=0.00609805f //x=21.505 //y=0.445
c328 ( 234 0 ) capacitor c=0.00505637f //x=21.42 //y=0.53
c329 ( 233 0 ) capacitor c=0.00468234f //x=21.02 //y=0.445
c330 ( 230 0 ) capacitor c=0.00537084f //x=20.935 //y=0.53
c331 ( 225 0 ) capacitor c=0.00468234f //x=20.535 //y=0.445
c332 ( 222 0 ) capacitor c=0.00537084f //x=20.45 //y=0.53
c333 ( 221 0 ) capacitor c=0.00468234f //x=20.05 //y=0.445
c334 ( 218 0 ) capacitor c=0.00634502f //x=19.965 //y=0.53
c335 ( 213 0 ) capacitor c=0.00609805f //x=19.565 //y=0.445
c336 ( 210 0 ) capacitor c=0.0195795f //x=19.48 //y=0
c337 ( 205 0 ) capacitor c=0.0659516f //x=18.26 //y=0
c338 ( 204 0 ) capacitor c=0.0195795f //x=18.7 //y=0
c339 ( 199 0 ) capacitor c=0.00609805f //x=18.175 //y=0.445
c340 ( 196 0 ) capacitor c=0.00505127f //x=18.09 //y=0.53
c341 ( 195 0 ) capacitor c=0.00468234f //x=17.69 //y=0.445
c342 ( 192 0 ) capacitor c=0.00537002f //x=17.605 //y=0.53
c343 ( 187 0 ) capacitor c=0.00468234f //x=17.205 //y=0.445
c344 ( 184 0 ) capacitor c=0.00556167f //x=17.12 //y=0.53
c345 ( 183 0 ) capacitor c=0.00468234f //x=16.72 //y=0.445
c346 ( 180 0 ) capacitor c=0.00642891f //x=16.635 //y=0.53
c347 ( 175 0 ) capacitor c=0.00609805f //x=16.235 //y=0.445
c348 ( 172 0 ) capacitor c=0.0227441f //x=16.15 //y=0
c349 ( 169 0 ) capacitor c=0.0360689f //x=15.005 //y=0
c350 ( 168 0 ) capacitor c=0.0184787f //x=15.37 //y=0
c351 ( 163 0 ) capacitor c=0.00583665f //x=14.92 //y=0.45
c352 ( 160 0 ) capacitor c=0.00536917f //x=14.835 //y=0.535
c353 ( 159 0 ) capacitor c=0.00479856f //x=14.435 //y=0.45
c354 ( 156 0 ) capacitor c=0.00640467f //x=14.35 //y=0.535
c355 ( 151 0 ) capacitor c=0.00588377f //x=13.95 //y=0.45
c356 ( 146 0 ) capacitor c=0.0164879f //x=13.865 //y=0
c357 ( 140 0 ) capacitor c=0.0720403f //x=13.15 //y=0
c358 ( 134 0 ) capacitor c=0.0389171f //x=11.085 //y=0
c359 ( 129 0 ) capacitor c=0.0360881f //x=9.455 //y=0
c360 ( 128 0 ) capacitor c=0.0160123f //x=9.82 //y=0
c361 ( 123 0 ) capacitor c=0.00583665f //x=9.37 //y=0.45
c362 ( 120 0 ) capacitor c=0.00531808f //x=9.285 //y=0.535
c363 ( 119 0 ) capacitor c=0.00479856f //x=8.885 //y=0.45
c364 ( 116 0 ) capacitor c=0.006266f //x=8.8 //y=0.535
c365 ( 111 0 ) capacitor c=0.00588377f //x=8.4 //y=0.45
c366 ( 108 0 ) capacitor c=0.0164879f //x=8.315 //y=0
c367 ( 100 0 ) capacitor c=0.0720721f //x=7.6 //y=0
c368 ( 92 0 ) capacitor c=0.0389171f //x=5.535 //y=0
c369 ( 89 0 ) capacitor c=0.0360881f //x=3.905 //y=0
c370 ( 88 0 ) capacitor c=0.0160123f //x=4.27 //y=0
c371 ( 83 0 ) capacitor c=0.00583665f //x=3.82 //y=0.45
c372 ( 80 0 ) capacitor c=0.00531808f //x=3.735 //y=0.535
c373 ( 79 0 ) capacitor c=0.00479856f //x=3.335 //y=0.45
c374 ( 76 0 ) capacitor c=0.006266f //x=3.25 //y=0.535
c375 ( 71 0 ) capacitor c=0.00592191f //x=2.85 //y=0.45
c376 ( 68 0 ) capacitor c=0.0164879f //x=2.765 //y=0
c377 ( 63 0 ) capacitor c=0.0360681f //x=1.685 //y=0
c378 ( 62 0 ) capacitor c=0.0160123f //x=2.05 //y=0
c379 ( 57 0 ) capacitor c=0.00587411f //x=1.6 //y=0.45
c380 ( 54 0 ) capacitor c=0.00536604f //x=1.515 //y=0.535
c381 ( 53 0 ) capacitor c=0.00479856f //x=1.115 //y=0.45
c382 ( 50 0 ) capacitor c=0.00707849f //x=1.03 //y=0.535
c383 ( 45 0 ) capacitor c=0.00592191f //x=0.63 //y=0.45
c384 ( 38 0 ) capacitor c=0.748287f //x=21.83 //y=0
r385 (  328 329 ) resistor r=14.8796 //w=0.357 //l=0.415 //layer=li \
 //thickness=0.1 //x=21.09 //y=0 //x2=21.505 //y2=0
r386 (  326 328 ) resistor r=2.5098 //w=0.357 //l=0.07 //layer=li \
 //thickness=0.1 //x=21.02 //y=0 //x2=21.09 //y2=0
r387 (  325 326 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.535 //y=0 //x2=21.02 //y2=0
r388 (  324 325 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.05 //y=0 //x2=20.535 //y2=0
r389 (  323 324 ) resistor r=2.5098 //w=0.357 //l=0.07 //layer=li \
 //thickness=0.1 //x=19.98 //y=0 //x2=20.05 //y2=0
r390 (  321 323 ) resistor r=14.8796 //w=0.357 //l=0.415 //layer=li \
 //thickness=0.1 //x=19.565 //y=0 //x2=19.98 //y2=0
r391 (  308 309 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.69 //y=0 //x2=18.175 //y2=0
r392 (  307 308 ) resistor r=10.7563 //w=0.357 //l=0.3 //layer=li \
 //thickness=0.1 //x=17.39 //y=0 //x2=17.69 //y2=0
r393 (  305 307 ) resistor r=6.63305 //w=0.357 //l=0.185 //layer=li \
 //thickness=0.1 //x=17.205 //y=0 //x2=17.39 //y2=0
r394 (  304 305 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.72 //y=0 //x2=17.205 //y2=0
r395 (  303 304 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=16.28 //y=0 //x2=16.72 //y2=0
r396 (  301 303 ) resistor r=1.61345 //w=0.357 //l=0.045 //layer=li \
 //thickness=0.1 //x=16.235 //y=0 //x2=16.28 //y2=0
r397 (  292 293 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=14.8 //y=0 //x2=14.92 //y2=0
r398 (  290 292 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=14.435 //y=0 //x2=14.8 //y2=0
r399 (  289 290 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=13.95 //y=0 //x2=14.435 //y2=0
r400 (  277 278 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.885 //y=0 //x2=9.37 //y2=0
r401 (  276 277 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=8.51 //y=0 //x2=8.885 //y2=0
r402 (  274 276 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=8.4 //y=0 //x2=8.51 //y2=0
r403 (  263 264 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.335 //y=0 //x2=3.82 //y2=0
r404 (  262 263 ) resistor r=0.179272 //w=0.357 //l=0.005 //layer=li \
 //thickness=0.1 //x=3.33 //y=0 //x2=3.335 //y2=0
r405 (  260 262 ) resistor r=17.2101 //w=0.357 //l=0.48 //layer=li \
 //thickness=0.1 //x=2.85 //y=0 //x2=3.33 //y2=0
r406 (  251 252 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.115 //y=0 //x2=1.6 //y2=0
r407 (  250 251 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.115 //y2=0
r408 (  248 250 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=0.63 //y=0 //x2=0.74 //y2=0
r409 (  243 329 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.59 //y=0 //x2=21.505 //y2=0
r410 (  243 245 ) resistor r=8.60504 //w=0.357 //l=0.24 //layer=li \
 //thickness=0.1 //x=21.59 //y=0 //x2=21.83 //y2=0
r411 (  238 347 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.505 //y=0.615 //x2=21.505 //y2=0.53
r412 (  238 347 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=21.505 //y=0.615 //x2=21.505 //y2=0.88
r413 (  237 347 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.505 //y=0.445 //x2=21.505 //y2=0.53
r414 (  236 329 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.505 //y=0.17 //x2=21.505 //y2=0
r415 (  236 237 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=21.505 //y=0.17 //x2=21.505 //y2=0.445
r416 (  235 347 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.105 //y=0.53 //x2=21.02 //y2=0.53
r417 (  234 347 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.42 //y=0.53 //x2=21.505 //y2=0.53
r418 (  234 235 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=21.42 //y=0.53 //x2=21.105 //y2=0.53
r419 (  233 347 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.02 //y=0.445 //x2=21.02 //y2=0.53
r420 (  232 326 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.02 //y=0.17 //x2=21.02 //y2=0
r421 (  232 233 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=21.02 //y=0.17 //x2=21.02 //y2=0.445
r422 (  231 347 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.62 //y=0.53 //x2=20.535 //y2=0.53
r423 (  230 347 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.935 //y=0.53 //x2=21.02 //y2=0.53
r424 (  230 231 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=20.935 //y=0.53 //x2=20.62 //y2=0.53
r425 (  226 347 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.535 //y=0.615 //x2=20.535 //y2=0.53
r426 (  226 347 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=20.535 //y=0.615 //x2=20.535 //y2=0.88
r427 (  225 347 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.535 //y=0.445 //x2=20.535 //y2=0.53
r428 (  224 325 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.535 //y=0.17 //x2=20.535 //y2=0
r429 (  224 225 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=20.535 //y=0.17 //x2=20.535 //y2=0.445
r430 (  223 347 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.135 //y=0.53 //x2=20.05 //y2=0.53
r431 (  222 347 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.45 //y=0.53 //x2=20.535 //y2=0.53
r432 (  222 223 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=20.45 //y=0.53 //x2=20.135 //y2=0.53
r433 (  221 347 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.05 //y=0.445 //x2=20.05 //y2=0.53
r434 (  220 324 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.05 //y=0.17 //x2=20.05 //y2=0
r435 (  220 221 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=20.05 //y=0.17 //x2=20.05 //y2=0.445
r436 (  219 347 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.65 //y=0.53 //x2=19.565 //y2=0.53
r437 (  218 347 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.965 //y=0.53 //x2=20.05 //y2=0.53
r438 (  218 219 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=19.965 //y=0.53 //x2=19.65 //y2=0.53
r439 (  214 347 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.565 //y=0.615 //x2=19.565 //y2=0.53
r440 (  214 347 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=19.565 //y=0.615 //x2=19.565 //y2=1.22
r441 (  213 347 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.565 //y=0.445 //x2=19.565 //y2=0.53
r442 (  212 321 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.565 //y=0.17 //x2=19.565 //y2=0
r443 (  212 213 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=19.565 //y=0.17 //x2=19.565 //y2=0.445
r444 (  211 320 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.04 //y=0 //x2=18.87 //y2=0
r445 (  210 321 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.48 //y=0 //x2=19.565 //y2=0
r446 (  210 211 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=19.48 //y=0 //x2=19.04 //y2=0
r447 (  205 309 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.26 //y=0 //x2=18.175 //y2=0
r448 (  205 207 ) resistor r=8.60504 //w=0.357 //l=0.24 //layer=li \
 //thickness=0.1 //x=18.26 //y=0 //x2=18.5 //y2=0
r449 (  204 320 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.7 //y=0 //x2=18.87 //y2=0
r450 (  204 207 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=18.7 //y=0 //x2=18.5 //y2=0
r451 (  200 346 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.175 //y=0.615 //x2=18.175 //y2=0.53
r452 (  200 346 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=18.175 //y=0.615 //x2=18.175 //y2=0.88
r453 (  199 346 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.175 //y=0.445 //x2=18.175 //y2=0.53
r454 (  198 309 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.175 //y=0.17 //x2=18.175 //y2=0
r455 (  198 199 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=18.175 //y=0.17 //x2=18.175 //y2=0.445
r456 (  197 346 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.775 //y=0.53 //x2=17.69 //y2=0.53
r457 (  196 346 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.09 //y=0.53 //x2=18.175 //y2=0.53
r458 (  196 197 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=18.09 //y=0.53 //x2=17.775 //y2=0.53
r459 (  195 346 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.69 //y=0.445 //x2=17.69 //y2=0.53
r460 (  194 308 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.69 //y=0.17 //x2=17.69 //y2=0
r461 (  194 195 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=17.69 //y=0.17 //x2=17.69 //y2=0.445
r462 (  193 346 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.29 //y=0.53 //x2=17.205 //y2=0.53
r463 (  192 346 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.605 //y=0.53 //x2=17.69 //y2=0.53
r464 (  192 193 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=17.605 //y=0.53 //x2=17.29 //y2=0.53
r465 (  188 346 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.205 //y=0.615 //x2=17.205 //y2=0.53
r466 (  188 346 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=17.205 //y=0.615 //x2=17.205 //y2=0.88
r467 (  187 346 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.205 //y=0.445 //x2=17.205 //y2=0.53
r468 (  186 305 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.205 //y=0.17 //x2=17.205 //y2=0
r469 (  186 187 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=17.205 //y=0.17 //x2=17.205 //y2=0.445
r470 (  185 346 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.805 //y=0.53 //x2=16.72 //y2=0.53
r471 (  184 346 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.12 //y=0.53 //x2=17.205 //y2=0.53
r472 (  184 185 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=17.12 //y=0.53 //x2=16.805 //y2=0.53
r473 (  183 346 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.72 //y=0.445 //x2=16.72 //y2=0.53
r474 (  182 304 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.72 //y=0.17 //x2=16.72 //y2=0
r475 (  182 183 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=16.72 //y=0.17 //x2=16.72 //y2=0.445
r476 (  181 346 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.32 //y=0.53 //x2=16.235 //y2=0.53
r477 (  180 346 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.635 //y=0.53 //x2=16.72 //y2=0.53
r478 (  180 181 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=16.635 //y=0.53 //x2=16.32 //y2=0.53
r479 (  176 346 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.235 //y=0.615 //x2=16.235 //y2=0.53
r480 (  176 346 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=16.235 //y=0.615 //x2=16.235 //y2=1.22
r481 (  175 346 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.235 //y=0.445 //x2=16.235 //y2=0.53
r482 (  174 301 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.235 //y=0.17 //x2=16.235 //y2=0
r483 (  174 175 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=16.235 //y=0.17 //x2=16.235 //y2=0.445
r484 (  173 300 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.71 //y=0 //x2=15.54 //y2=0
r485 (  172 301 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.15 //y=0 //x2=16.235 //y2=0
r486 (  172 173 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=16.15 //y=0 //x2=15.71 //y2=0
r487 (  169 293 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.005 //y=0 //x2=14.92 //y2=0
r488 (  168 300 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.37 //y=0 //x2=15.54 //y2=0
r489 (  168 169 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=15.37 //y=0 //x2=15.005 //y2=0
r490 (  164 345 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.92 //y=0.62 //x2=14.92 //y2=0.535
r491 (  164 345 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=14.92 //y=0.62 //x2=14.92 //y2=1.225
r492 (  163 345 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.92 //y=0.45 //x2=14.92 //y2=0.535
r493 (  162 293 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.92 //y=0.17 //x2=14.92 //y2=0
r494 (  162 163 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=14.92 //y=0.17 //x2=14.92 //y2=0.45
r495 (  161 345 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.52 //y=0.535 //x2=14.435 //y2=0.535
r496 (  160 345 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.835 //y=0.535 //x2=14.92 //y2=0.535
r497 (  160 161 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=14.835 //y=0.535 //x2=14.52 //y2=0.535
r498 (  159 345 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.435 //y=0.45 //x2=14.435 //y2=0.535
r499 (  158 290 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.435 //y=0.17 //x2=14.435 //y2=0
r500 (  158 159 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=14.435 //y=0.17 //x2=14.435 //y2=0.45
r501 (  157 345 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.035 //y=0.535 //x2=13.95 //y2=0.535
r502 (  156 345 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.35 //y=0.535 //x2=14.435 //y2=0.535
r503 (  156 157 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=14.35 //y=0.535 //x2=14.035 //y2=0.535
r504 (  152 345 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.95 //y=0.62 //x2=13.95 //y2=0.535
r505 (  152 345 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=13.95 //y=0.62 //x2=13.95 //y2=1.225
r506 (  151 345 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.95 //y=0.45 //x2=13.95 //y2=0.535
r507 (  150 289 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.95 //y=0.17 //x2=13.95 //y2=0
r508 (  150 151 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=13.95 //y=0.17 //x2=13.95 //y2=0.45
r509 (  147 288 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.49 //y=0 //x2=13.32 //y2=0
r510 (  147 149 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=13.49 //y=0 //x2=13.69 //y2=0
r511 (  146 289 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.865 //y=0 //x2=13.95 //y2=0
r512 (  146 149 ) resistor r=6.27451 //w=0.357 //l=0.175 //layer=li \
 //thickness=0.1 //x=13.865 //y=0 //x2=13.69 //y2=0
r513 (  141 287 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.255 //y=0 //x2=11.17 //y2=0
r514 (  141 143 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=11.255 //y=0 //x2=12.21 //y2=0
r515 (  140 288 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.15 //y=0 //x2=13.32 //y2=0
r516 (  140 143 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=13.15 //y=0 //x2=12.21 //y2=0
r517 (  136 287 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.17 //y=0.17 //x2=11.17 //y2=0
r518 (  136 344 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=11.17 //y=0.17 //x2=11.17 //y2=0.955
r519 (  135 285 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.16 //y=0 //x2=9.99 //y2=0
r520 (  134 287 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.085 //y=0 //x2=11.17 //y2=0
r521 (  134 135 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=11.085 //y=0 //x2=10.16 //y2=0
r522 (  129 278 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.455 //y=0 //x2=9.37 //y2=0
r523 (  129 131 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=9.455 //y=0 //x2=9.62 //y2=0
r524 (  128 285 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.82 //y=0 //x2=9.99 //y2=0
r525 (  128 131 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=9.82 //y=0 //x2=9.62 //y2=0
r526 (  124 343 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.37 //y=0.62 //x2=9.37 //y2=0.535
r527 (  124 343 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=9.37 //y=0.62 //x2=9.37 //y2=1.225
r528 (  123 343 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.37 //y=0.45 //x2=9.37 //y2=0.535
r529 (  122 278 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.37 //y=0.17 //x2=9.37 //y2=0
r530 (  122 123 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=9.37 //y=0.17 //x2=9.37 //y2=0.45
r531 (  121 343 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.97 //y=0.535 //x2=8.885 //y2=0.535
r532 (  120 343 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.285 //y=0.535 //x2=9.37 //y2=0.535
r533 (  120 121 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=9.285 //y=0.535 //x2=8.97 //y2=0.535
r534 (  119 343 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.885 //y=0.45 //x2=8.885 //y2=0.535
r535 (  118 277 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.885 //y=0.17 //x2=8.885 //y2=0
r536 (  118 119 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=8.885 //y=0.17 //x2=8.885 //y2=0.45
r537 (  117 343 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.485 //y=0.535 //x2=8.4 //y2=0.535
r538 (  116 343 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.8 //y=0.535 //x2=8.885 //y2=0.535
r539 (  116 117 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=8.8 //y=0.535 //x2=8.485 //y2=0.535
r540 (  112 343 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.4 //y=0.62 //x2=8.4 //y2=0.535
r541 (  112 343 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=8.4 //y=0.62 //x2=8.4 //y2=1.225
r542 (  111 343 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.4 //y=0.45 //x2=8.4 //y2=0.535
r543 (  110 274 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.4 //y=0.17 //x2=8.4 //y2=0
r544 (  110 111 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=8.4 //y=0.17 //x2=8.4 //y2=0.45
r545 (  109 273 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.94 //y=0 //x2=7.77 //y2=0
r546 (  108 274 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.315 //y=0 //x2=8.4 //y2=0
r547 (  108 109 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=8.315 //y=0 //x2=7.94 //y2=0
r548 (  103 105 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=5.92 //y=0 //x2=7.03 //y2=0
r549 (  101 272 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.705 //y=0 //x2=5.62 //y2=0
r550 (  101 103 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=5.705 //y=0 //x2=5.92 //y2=0
r551 (  100 273 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.6 //y=0 //x2=7.77 //y2=0
r552 (  100 105 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=7.6 //y=0 //x2=7.03 //y2=0
r553 (  96 272 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.62 //y=0.17 //x2=5.62 //y2=0
r554 (  96 342 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=5.62 //y=0.17 //x2=5.62 //y2=0.955
r555 (  93 271 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.61 //y=0 //x2=4.44 //y2=0
r556 (  93 95 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=4.61 //y=0 //x2=4.81 //y2=0
r557 (  92 272 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.535 //y=0 //x2=5.62 //y2=0
r558 (  92 95 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=5.535 //y=0 //x2=4.81 //y2=0
r559 (  89 264 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.905 //y=0 //x2=3.82 //y2=0
r560 (  88 271 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.27 //y=0 //x2=4.44 //y2=0
r561 (  88 89 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=4.27 //y=0 //x2=3.905 //y2=0
r562 (  84 341 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.82 //y=0.62 //x2=3.82 //y2=0.535
r563 (  84 341 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=3.82 //y=0.62 //x2=3.82 //y2=1.225
r564 (  83 341 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.82 //y=0.45 //x2=3.82 //y2=0.535
r565 (  82 264 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.82 //y=0.17 //x2=3.82 //y2=0
r566 (  82 83 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=3.82 //y=0.17 //x2=3.82 //y2=0.45
r567 (  81 341 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.42 //y=0.535 //x2=3.335 //y2=0.535
r568 (  80 341 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.735 //y=0.535 //x2=3.82 //y2=0.535
r569 (  80 81 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.735 //y=0.535 //x2=3.42 //y2=0.535
r570 (  79 341 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.335 //y=0.45 //x2=3.335 //y2=0.535
r571 (  78 263 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.335 //y=0.17 //x2=3.335 //y2=0
r572 (  78 79 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=3.335 //y=0.17 //x2=3.335 //y2=0.45
r573 (  77 341 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=0.535 //x2=2.85 //y2=0.535
r574 (  76 341 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.25 //y=0.535 //x2=3.335 //y2=0.535
r575 (  76 77 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.25 //y=0.535 //x2=2.935 //y2=0.535
r576 (  72 341 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.85 //y=0.62 //x2=2.85 //y2=0.535
r577 (  72 341 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=2.85 //y=0.62 //x2=2.85 //y2=1.225
r578 (  71 341 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.85 //y=0.45 //x2=2.85 //y2=0.535
r579 (  70 260 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.85 //y=0.17 //x2=2.85 //y2=0
r580 (  70 71 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=2.85 //y=0.17 //x2=2.85 //y2=0.45
r581 (  69 259 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.39 //y=0 //x2=2.22 //y2=0
r582 (  68 260 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=0 //x2=2.85 //y2=0
r583 (  68 69 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=2.765 //y=0 //x2=2.39 //y2=0
r584 (  63 252 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.685 //y=0 //x2=1.6 //y2=0
r585 (  63 65 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=1.685 //y=0 //x2=1.85 //y2=0
r586 (  62 259 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.05 //y=0 //x2=2.22 //y2=0
r587 (  62 65 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=2.05 //y=0 //x2=1.85 //y2=0
r588 (  58 340 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=0.535
r589 (  58 340 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=1.225
r590 (  57 340 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.45 //x2=1.6 //y2=0.535
r591 (  56 252 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0
r592 (  56 57 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0.45
r593 (  55 340 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.2 //y=0.535 //x2=1.115 //y2=0.535
r594 (  54 340 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.6 //y2=0.535
r595 (  54 55 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.2 //y2=0.535
r596 (  53 340 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.45 //x2=1.115 //y2=0.535
r597 (  52 251 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0
r598 (  52 53 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0.45
r599 (  51 340 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.715 //y=0.535 //x2=0.63 //y2=0.535
r600 (  50 340 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=1.115 //y2=0.535
r601 (  50 51 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=0.715 //y2=0.535
r602 (  46 340 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=0.535
r603 (  46 340 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=1.225
r604 (  45 340 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.45 //x2=0.63 //y2=0.535
r605 (  44 248 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0
r606 (  44 45 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0.45
r607 (  38 245 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.83 //y=0 //x2=21.83 //y2=0
r608 (  36 328 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=0 //x2=21.09 //y2=0
r609 (  36 38 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=0 //x2=21.83 //y2=0
r610 (  34 323 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=0 //x2=19.98 //y2=0
r611 (  34 36 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=0 //x2=21.09 //y2=0
r612 (  32 207 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=0 //x2=18.5 //y2=0
r613 (  32 34 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=0 //x2=19.98 //y2=0
r614 (  30 307 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=0 //x2=17.39 //y2=0
r615 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=0 //x2=18.5 //y2=0
r616 (  28 303 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=0 //x2=16.28 //y2=0
r617 (  28 30 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=0 //x2=17.39 //y2=0
r618 (  26 292 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.8 //y=0 //x2=14.8 //y2=0
r619 (  26 28 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=14.8 //y=0 //x2=16.28 //y2=0
r620 (  24 149 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=0 //x2=13.69 //y2=0
r621 (  24 26 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=13.69 //y=0 //x2=14.8 //y2=0
r622 (  22 143 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.21 //y=0 //x2=12.21 //y2=0
r623 (  22 24 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.21 //y=0 //x2=13.69 //y2=0
r624 (  18 131 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.62 //y=0 //x2=9.62 //y2=0
r625 (  16 276 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.51 //y=0 //x2=8.51 //y2=0
r626 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=8.51 //y=0 //x2=9.62 //y2=0
r627 (  14 105 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=0 //x2=7.03 //y2=0
r628 (  14 16 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=0 //x2=8.51 //y2=0
r629 (  12 103 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.92 //y=0 //x2=5.92 //y2=0
r630 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.92 //y=0 //x2=7.03 //y2=0
r631 (  10 95 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.81 //y=0 //x2=4.81 //y2=0
r632 (  10 12 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.81 //y=0 //x2=5.92 //y2=0
r633 (  8 262 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=3.33 //y=0 //x2=3.33 //y2=0
r634 (  8 10 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=0 //x2=4.81 //y2=0
r635 (  6 65 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r636 (  6 8 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=3.33 //y2=0
r637 (  3 250 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r638 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r639 (  1 287 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.1 //y=0 //x2=11.1 //y2=0
r640 (  1 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.1 //y=0 //x2=12.21 //y2=0
r641 (  1 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=11.1 //y=0 //x2=9.62 //y2=0
ends PM_DLATCHN\%GND

subckt PM_DLATCHN\%VDD ( 1 38 50 72 82 86 96 106 114 118 126 134 140 148 158 \
 182 190 194 204 212 227 231 233 236 241 245 249 253 255 257 258 259 260 261 \
 262 263 264 265 266 267 268 269 270 271 272 )
c295 ( 272 0 ) capacitor c=0.0255388f //x=19.955 //y=5.025
c296 ( 271 0 ) capacitor c=0.0255739f //x=16.625 //y=5.025
c297 ( 270 0 ) capacitor c=0.0433929f //x=14.73 //y=5.02
c298 ( 269 0 ) capacitor c=0.0422979f //x=13.86 //y=5.02
c299 ( 268 0 ) capacitor c=0.0382117f //x=12.395 //y=5.02
c300 ( 267 0 ) capacitor c=0.0240874f //x=11.515 //y=5.02
c301 ( 266 0 ) capacitor c=0.0494569f //x=10.645 //y=5.02
c302 ( 265 0 ) capacitor c=0.0432963f //x=9.18 //y=5.02
c303 ( 264 0 ) capacitor c=0.0422219f //x=8.31 //y=5.02
c304 ( 263 0 ) capacitor c=0.0381505f //x=6.845 //y=5.02
c305 ( 262 0 ) capacitor c=0.0240879f //x=5.965 //y=5.02
c306 ( 261 0 ) capacitor c=0.0494569f //x=5.095 //y=5.02
c307 ( 260 0 ) capacitor c=0.0432963f //x=3.63 //y=5.02
c308 ( 259 0 ) capacitor c=0.0421596f //x=2.76 //y=5.02
c309 ( 258 0 ) capacitor c=0.0438108f //x=1.41 //y=5.02
c310 ( 257 0 ) capacitor c=0.0427416f //x=0.54 //y=5.02
c311 ( 256 0 ) capacitor c=0.00591168f //x=20.1 //y=7.4
c312 ( 255 0 ) capacitor c=0.111374f //x=18.87 //y=7.4
c313 ( 254 0 ) capacitor c=0.00591168f //x=16.77 //y=7.4
c314 ( 253 0 ) capacitor c=0.109883f //x=15.54 //y=7.4
c315 ( 252 0 ) capacitor c=0.00591168f //x=14.8 //y=7.4
c316 ( 250 0 ) capacitor c=0.00591168f //x=13.995 //y=7.4
c317 ( 249 0 ) capacitor c=0.109921f //x=13.32 //y=7.4
c318 ( 248 0 ) capacitor c=0.00591168f //x=12.54 //y=7.4
c319 ( 247 0 ) capacitor c=0.00591168f //x=11.66 //y=7.4
c320 ( 246 0 ) capacitor c=0.00591168f //x=10.78 //y=7.4
c321 ( 245 0 ) capacitor c=0.114228f //x=9.99 //y=7.4
c322 ( 244 0 ) capacitor c=0.00591168f //x=9.325 //y=7.4
c323 ( 243 0 ) capacitor c=0.00591168f //x=8.51 //y=7.4
c324 ( 241 0 ) capacitor c=0.108342f //x=7.77 //y=7.4
c325 ( 240 0 ) capacitor c=0.00591168f //x=7.03 //y=7.4
c326 ( 238 0 ) capacitor c=0.00591168f //x=6.11 //y=7.4
c327 ( 237 0 ) capacitor c=0.00591168f //x=5.23 //y=7.4
c328 ( 236 0 ) capacitor c=0.114226f //x=4.44 //y=7.4
c329 ( 235 0 ) capacitor c=0.00591168f //x=3.775 //y=7.4
c330 ( 234 0 ) capacitor c=0.00591168f //x=2.895 //y=7.4
c331 ( 233 0 ) capacitor c=0.108542f //x=2.22 //y=7.4
c332 ( 232 0 ) capacitor c=0.00591168f //x=1.555 //y=7.4
c333 ( 231 0 ) capacitor c=0.23322f //x=0.74 //y=7.4
c334 ( 227 0 ) capacitor c=0.287249f //x=21.83 //y=7.4
c335 ( 212 0 ) capacitor c=0.0427882f //x=20.015 //y=7.4
c336 ( 204 0 ) capacitor c=0.074729f //x=18.7 //y=7.4
c337 ( 194 0 ) capacitor c=0.0427882f //x=16.685 //y=7.4
c338 ( 190 0 ) capacitor c=0.0181526f //x=15.37 //y=7.4
c339 ( 182 0 ) capacitor c=0.0288426f //x=14.79 //y=7.4
c340 ( 172 0 ) capacitor c=0.0216067f //x=13.91 //y=7.4
c341 ( 168 0 ) capacitor c=0.0275781f //x=13.15 //y=7.4
c342 ( 158 0 ) capacitor c=0.0284327f //x=12.455 //y=7.4
c343 ( 148 0 ) capacitor c=0.0288633f //x=11.575 //y=7.4
c344 ( 140 0 ) capacitor c=0.0240981f //x=10.695 //y=7.4
c345 ( 134 0 ) capacitor c=0.0181526f //x=9.82 //y=7.4
c346 ( 126 0 ) capacitor c=0.0289624f //x=9.24 //y=7.4
c347 ( 118 0 ) capacitor c=0.0186283f //x=8.36 //y=7.4
c348 ( 114 0 ) capacitor c=0.0236224f //x=7.6 //y=7.4
c349 ( 106 0 ) capacitor c=0.0288639f //x=6.905 //y=7.4
c350 ( 96 0 ) capacitor c=0.0288633f //x=6.025 //y=7.4
c351 ( 86 0 ) capacitor c=0.0240981f //x=5.145 //y=7.4
c352 ( 82 0 ) capacitor c=0.0181526f //x=4.27 //y=7.4
c353 ( 72 0 ) capacitor c=0.0291066f //x=3.69 //y=7.4
c354 ( 64 0 ) capacitor c=0.0216067f //x=2.81 //y=7.4
c355 ( 58 0 ) capacitor c=0.0210379f //x=2.05 //y=7.4
c356 ( 50 0 ) capacitor c=0.0287207f //x=1.47 //y=7.4
c357 ( 38 0 ) capacitor c=0.768357f //x=21.83 //y=7.4
r358 (  225 227 ) resistor r=26.5322 //w=0.357 //l=0.74 //layer=li \
 //thickness=0.1 //x=21.09 //y=7.4 //x2=21.83 //y2=7.4
r359 (  223 256 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.185 //y=7.4 //x2=20.1 //y2=7.4
r360 (  223 225 ) resistor r=32.4482 //w=0.357 //l=0.905 //layer=li \
 //thickness=0.1 //x=20.185 //y=7.4 //x2=21.09 //y2=7.4
r361 (  216 256 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.1 //y=7.23 //x2=20.1 //y2=7.4
r362 (  216 272 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=20.1 //y=7.23 //x2=20.1 //y2=6.74
r363 (  213 255 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.04 //y=7.4 //x2=18.87 //y2=7.4
r364 (  213 215 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=19.04 //y=7.4 //x2=19.98 //y2=7.4
r365 (  212 256 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.015 //y=7.4 //x2=20.1 //y2=7.4
r366 (  212 215 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=20.015 //y=7.4 //x2=19.98 //y2=7.4
r367 (  207 209 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=17.39 //y=7.4 //x2=18.5 //y2=7.4
r368 (  205 254 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.855 //y=7.4 //x2=16.77 //y2=7.4
r369 (  205 207 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=16.855 //y=7.4 //x2=17.39 //y2=7.4
r370 (  204 255 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.7 //y=7.4 //x2=18.87 //y2=7.4
r371 (  204 209 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=18.7 //y=7.4 //x2=18.5 //y2=7.4
r372 (  198 254 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.77 //y=7.23 //x2=16.77 //y2=7.4
r373 (  198 271 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=16.77 //y=7.23 //x2=16.77 //y2=6.74
r374 (  195 253 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.71 //y=7.4 //x2=15.54 //y2=7.4
r375 (  195 197 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=15.71 //y=7.4 //x2=16.28 //y2=7.4
r376 (  194 254 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.685 //y=7.4 //x2=16.77 //y2=7.4
r377 (  194 197 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=16.685 //y=7.4 //x2=16.28 //y2=7.4
r378 (  191 252 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.96 //y=7.4 //x2=14.875 //y2=7.4
r379 (  190 253 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.37 //y=7.4 //x2=15.54 //y2=7.4
r380 (  190 191 ) resistor r=14.7003 //w=0.357 //l=0.41 //layer=li \
 //thickness=0.1 //x=15.37 //y=7.4 //x2=14.96 //y2=7.4
r381 (  184 252 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.875 //y=7.23 //x2=14.875 //y2=7.4
r382 (  184 270 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=14.875 //y=7.23 //x2=14.875 //y2=6.405
r383 (  183 250 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.08 //y=7.4 //x2=13.995 //y2=7.4
r384 (  182 252 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.79 //y=7.4 //x2=14.875 //y2=7.4
r385 (  182 183 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=14.79 //y=7.4 //x2=14.08 //y2=7.4
r386 (  176 250 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.995 //y=7.23 //x2=13.995 //y2=7.4
r387 (  176 269 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=13.995 //y=7.23 //x2=13.995 //y2=6.405
r388 (  173 249 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.49 //y=7.4 //x2=13.32 //y2=7.4
r389 (  173 175 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=13.49 //y=7.4 //x2=13.69 //y2=7.4
r390 (  172 250 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.91 //y=7.4 //x2=13.995 //y2=7.4
r391 (  172 175 ) resistor r=7.88796 //w=0.357 //l=0.22 //layer=li \
 //thickness=0.1 //x=13.91 //y=7.4 //x2=13.69 //y2=7.4
r392 (  169 248 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.625 //y=7.4 //x2=12.54 //y2=7.4
r393 (  168 249 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.15 //y=7.4 //x2=13.32 //y2=7.4
r394 (  168 169 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=13.15 //y=7.4 //x2=12.625 //y2=7.4
r395 (  162 248 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.54 //y=7.23 //x2=12.54 //y2=7.4
r396 (  162 268 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.54 //y=7.23 //x2=12.54 //y2=6.745
r397 (  159 247 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.745 //y=7.4 //x2=11.66 //y2=7.4
r398 (  159 161 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=11.745 //y=7.4 //x2=12.21 //y2=7.4
r399 (  158 248 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.455 //y=7.4 //x2=12.54 //y2=7.4
r400 (  158 161 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=12.455 //y=7.4 //x2=12.21 //y2=7.4
r401 (  152 247 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.66 //y=7.23 //x2=11.66 //y2=7.4
r402 (  152 267 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.66 //y=7.23 //x2=11.66 //y2=6.745
r403 (  149 246 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.865 //y=7.4 //x2=10.78 //y2=7.4
r404 (  149 151 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=10.865 //y=7.4 //x2=11.1 //y2=7.4
r405 (  148 247 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.575 //y=7.4 //x2=11.66 //y2=7.4
r406 (  148 151 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=11.575 //y=7.4 //x2=11.1 //y2=7.4
r407 (  142 246 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.78 //y=7.23 //x2=10.78 //y2=7.4
r408 (  142 266 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=10.78 //y=7.23 //x2=10.78 //y2=6.405
r409 (  141 245 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.16 //y=7.4 //x2=9.99 //y2=7.4
r410 (  140 246 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.695 //y=7.4 //x2=10.78 //y2=7.4
r411 (  140 141 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=10.695 //y=7.4 //x2=10.16 //y2=7.4
r412 (  135 244 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.41 //y=7.4 //x2=9.325 //y2=7.4
r413 (  135 137 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=9.41 //y=7.4 //x2=9.62 //y2=7.4
r414 (  134 245 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.82 //y=7.4 //x2=9.99 //y2=7.4
r415 (  134 137 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=9.82 //y=7.4 //x2=9.62 //y2=7.4
r416 (  128 244 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.325 //y=7.23 //x2=9.325 //y2=7.4
r417 (  128 265 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=9.325 //y=7.23 //x2=9.325 //y2=6.405
r418 (  127 243 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.53 //y=7.4 //x2=8.445 //y2=7.4
r419 (  126 244 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.24 //y=7.4 //x2=9.325 //y2=7.4
r420 (  126 127 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=9.24 //y=7.4 //x2=8.53 //y2=7.4
r421 (  120 243 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.445 //y=7.23 //x2=8.445 //y2=7.4
r422 (  120 264 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=8.445 //y=7.23 //x2=8.445 //y2=6.405
r423 (  119 241 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.94 //y=7.4 //x2=7.77 //y2=7.4
r424 (  118 243 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.36 //y=7.4 //x2=8.445 //y2=7.4
r425 (  118 119 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=8.36 //y=7.4 //x2=7.94 //y2=7.4
r426 (  115 240 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.075 //y=7.4 //x2=6.99 //y2=7.4
r427 (  114 241 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.6 //y=7.4 //x2=7.77 //y2=7.4
r428 (  114 115 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=7.6 //y=7.4 //x2=7.075 //y2=7.4
r429 (  108 240 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.99 //y=7.23 //x2=6.99 //y2=7.4
r430 (  108 263 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.99 //y=7.23 //x2=6.99 //y2=6.745
r431 (  107 238 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.195 //y=7.4 //x2=6.11 //y2=7.4
r432 (  106 240 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.905 //y=7.4 //x2=6.99 //y2=7.4
r433 (  106 107 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=6.905 //y=7.4 //x2=6.195 //y2=7.4
r434 (  100 238 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.11 //y=7.23 //x2=6.11 //y2=7.4
r435 (  100 262 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.11 //y=7.23 //x2=6.11 //y2=6.745
r436 (  97 237 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.315 //y=7.4 //x2=5.23 //y2=7.4
r437 (  97 99 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=5.315 //y=7.4 //x2=5.92 //y2=7.4
r438 (  96 238 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.025 //y=7.4 //x2=6.11 //y2=7.4
r439 (  96 99 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=6.025 //y=7.4 //x2=5.92 //y2=7.4
r440 (  90 237 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.23 //y=7.23 //x2=5.23 //y2=7.4
r441 (  90 261 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=5.23 //y=7.23 //x2=5.23 //y2=6.405
r442 (  87 236 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.61 //y=7.4 //x2=4.44 //y2=7.4
r443 (  87 89 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=4.61 //y=7.4 //x2=4.81 //y2=7.4
r444 (  86 237 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.145 //y=7.4 //x2=5.23 //y2=7.4
r445 (  86 89 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=5.145 //y=7.4 //x2=4.81 //y2=7.4
r446 (  83 235 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.86 //y=7.4 //x2=3.775 //y2=7.4
r447 (  82 236 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.27 //y=7.4 //x2=4.44 //y2=7.4
r448 (  82 83 ) resistor r=14.7003 //w=0.357 //l=0.41 //layer=li \
 //thickness=0.1 //x=4.27 //y=7.4 //x2=3.86 //y2=7.4
r449 (  76 235 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.775 //y=7.23 //x2=3.775 //y2=7.4
r450 (  76 260 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=3.775 //y=7.23 //x2=3.775 //y2=6.405
r451 (  73 234 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.98 //y=7.4 //x2=2.895 //y2=7.4
r452 (  73 75 ) resistor r=12.549 //w=0.357 //l=0.35 //layer=li \
 //thickness=0.1 //x=2.98 //y=7.4 //x2=3.33 //y2=7.4
r453 (  72 235 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.69 //y=7.4 //x2=3.775 //y2=7.4
r454 (  72 75 ) resistor r=12.9076 //w=0.357 //l=0.36 //layer=li \
 //thickness=0.1 //x=3.69 //y=7.4 //x2=3.33 //y2=7.4
r455 (  66 234 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.895 //y=7.23 //x2=2.895 //y2=7.4
r456 (  66 259 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=2.895 //y=7.23 //x2=2.895 //y2=6.405
r457 (  65 233 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.39 //y=7.4 //x2=2.22 //y2=7.4
r458 (  64 234 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.81 //y=7.4 //x2=2.895 //y2=7.4
r459 (  64 65 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=2.81 //y=7.4 //x2=2.39 //y2=7.4
r460 (  59 232 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.64 //y=7.4 //x2=1.555 //y2=7.4
r461 (  59 61 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=1.64 //y=7.4 //x2=1.85 //y2=7.4
r462 (  58 233 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.05 //y=7.4 //x2=2.22 //y2=7.4
r463 (  58 61 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=2.05 //y=7.4 //x2=1.85 //y2=7.4
r464 (  52 232 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=7.4
r465 (  52 258 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=6.405
r466 (  51 231 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.76 //y=7.4 //x2=0.675 //y2=7.4
r467 (  50 232 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=1.555 //y2=7.4
r468 (  50 51 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=0.76 //y2=7.4
r469 (  44 231 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=7.4
r470 (  44 257 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=6.405
r471 (  38 227 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.83 //y=7.4 //x2=21.83 //y2=7.4
r472 (  36 225 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=7.4 //x2=21.09 //y2=7.4
r473 (  36 38 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=7.4 //x2=21.83 //y2=7.4
r474 (  34 215 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=7.4 //x2=19.98 //y2=7.4
r475 (  34 36 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=7.4 //x2=21.09 //y2=7.4
r476 (  32 209 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=7.4 //x2=18.5 //y2=7.4
r477 (  32 34 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=7.4 //x2=19.98 //y2=7.4
r478 (  30 207 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=7.4 //x2=17.39 //y2=7.4
r479 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=7.4 //x2=18.5 //y2=7.4
r480 (  28 197 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=7.4 //x2=16.28 //y2=7.4
r481 (  28 30 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=7.4 //x2=17.39 //y2=7.4
r482 (  26 252 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.8 //y=7.4 //x2=14.8 //y2=7.4
r483 (  26 28 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=14.8 //y=7.4 //x2=16.28 //y2=7.4
r484 (  24 175 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=7.4 //x2=13.69 //y2=7.4
r485 (  24 26 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=13.69 //y=7.4 //x2=14.8 //y2=7.4
r486 (  22 161 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.21 //y=7.4 //x2=12.21 //y2=7.4
r487 (  22 24 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.21 //y=7.4 //x2=13.69 //y2=7.4
r488 (  18 137 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.62 //y=7.4 //x2=9.62 //y2=7.4
r489 (  16 243 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.51 //y=7.4 //x2=8.51 //y2=7.4
r490 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=8.51 //y=7.4 //x2=9.62 //y2=7.4
r491 (  14 240 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=7.4 //x2=7.03 //y2=7.4
r492 (  14 16 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=7.4 //x2=8.51 //y2=7.4
r493 (  12 99 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.92 //y=7.4 //x2=5.92 //y2=7.4
r494 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.92 //y=7.4 //x2=7.03 //y2=7.4
r495 (  10 89 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.81 //y=7.4 //x2=4.81 //y2=7.4
r496 (  10 12 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.81 //y=7.4 //x2=5.92 //y2=7.4
r497 (  8 75 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=3.33 //y=7.4 //x2=3.33 //y2=7.4
r498 (  8 10 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=7.4 //x2=4.81 //y2=7.4
r499 (  6 61 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r500 (  6 8 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=3.33 //y2=7.4
r501 (  3 231 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r502 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r503 (  1 151 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.1 //y=7.4 //x2=11.1 //y2=7.4
r504 (  1 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.1 //y=7.4 //x2=12.21 //y2=7.4
r505 (  1 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=11.1 //y=7.4 //x2=9.62 //y2=7.4
ends PM_DLATCHN\%VDD

subckt PM_DLATCHN\%noxref_3 ( 1 2 17 18 19 20 24 26 33 34 35 36 37 38 39 43 45 \
 48 49 59 62 64 )
c117 ( 64 0 ) capacitor c=0.0288745f //x=3.19 //y=5.02
c118 ( 62 0 ) capacitor c=0.0173218f //x=3.145 //y=0.91
c119 ( 59 0 ) capacitor c=0.0593152f //x=5.55 //y=4.7
c120 ( 49 0 ) capacitor c=0.0318948f //x=5.885 //y=1.21
c121 ( 48 0 ) capacitor c=0.0187384f //x=5.885 //y=0.865
c122 ( 45 0 ) capacitor c=0.0141798f //x=5.73 //y=1.365
c123 ( 43 0 ) capacitor c=0.0149844f //x=5.73 //y=0.71
c124 ( 39 0 ) capacitor c=0.0819799f //x=5.355 //y=1.915
c125 ( 38 0 ) capacitor c=0.0229722f //x=5.355 //y=1.52
c126 ( 37 0 ) capacitor c=0.0234352f //x=5.355 //y=1.21
c127 ( 36 0 ) capacitor c=0.0199343f //x=5.355 //y=0.865
c128 ( 35 0 ) capacitor c=0.110275f //x=5.89 //y=6.02
c129 ( 34 0 ) capacitor c=0.154305f //x=5.45 //y=6.02
c130 ( 26 0 ) capacitor c=0.0930091f //x=5.55 //y=2.08
c131 ( 24 0 ) capacitor c=0.083023f //x=3.7 //y=3.7
c132 ( 20 0 ) capacitor c=0.00417404f //x=3.42 //y=4.58
c133 ( 19 0 ) capacitor c=0.0118896f //x=3.615 //y=4.58
c134 ( 18 0 ) capacitor c=0.00549299f //x=3.415 //y=2.08
c135 ( 17 0 ) capacitor c=0.013178f //x=3.615 //y=2.08
c136 ( 2 0 ) capacitor c=0.0123469f //x=3.815 //y=3.7
c137 ( 1 0 ) capacitor c=0.0440072f //x=5.435 //y=3.7
r138 (  57 59 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=5.45 //y=4.7 //x2=5.55 //y2=4.7
r139 (  50 59 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=5.89 //y=4.865 //x2=5.55 //y2=4.7
r140 (  49 61 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.21 //x2=5.845 //y2=1.365
r141 (  48 60 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.885 //y=0.865 //x2=5.845 //y2=0.71
r142 (  48 49 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.885 //y=0.865 //x2=5.885 //y2=1.21
r143 (  46 56 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.51 //y=1.365 //x2=5.395 //y2=1.365
r144 (  45 61 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.73 //y=1.365 //x2=5.845 //y2=1.365
r145 (  44 55 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.51 //y=0.71 //x2=5.395 //y2=0.71
r146 (  43 60 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.73 //y=0.71 //x2=5.845 //y2=0.71
r147 (  43 44 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=5.73 //y=0.71 //x2=5.51 //y2=0.71
r148 (  40 57 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=5.45 //y=4.865 //x2=5.45 //y2=4.7
r149 (  39 54 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=5.355 //y=1.915 //x2=5.55 //y2=2.08
r150 (  38 56 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.355 //y=1.52 //x2=5.395 //y2=1.365
r151 (  38 39 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=5.355 //y=1.52 //x2=5.355 //y2=1.915
r152 (  37 56 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.355 //y=1.21 //x2=5.395 //y2=1.365
r153 (  36 55 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.355 //y=0.865 //x2=5.395 //y2=0.71
r154 (  36 37 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.355 //y=0.865 //x2=5.355 //y2=1.21
r155 (  35 50 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.89 //y=6.02 //x2=5.89 //y2=4.865
r156 (  34 40 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.45 //y=6.02 //x2=5.45 //y2=4.865
r157 (  33 45 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.365 //x2=5.73 //y2=1.365
r158 (  33 46 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.365 //x2=5.51 //y2=1.365
r159 (  31 59 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.55 //y=4.7 //x2=5.55 //y2=4.7
r160 (  29 31 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=5.55 //y=3.7 //x2=5.55 //y2=4.7
r161 (  26 54 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.55 //y=2.08 //x2=5.55 //y2=2.08
r162 (  26 29 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=5.55 //y=2.08 //x2=5.55 //y2=3.7
r163 (  22 24 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=3.7 //y=4.495 //x2=3.7 //y2=3.7
r164 (  21 24 ) resistor r=105.07 //w=0.187 //l=1.535 //layer=li \
 //thickness=0.1 //x=3.7 //y=2.165 //x2=3.7 //y2=3.7
r165 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.615 //y=4.58 //x2=3.7 //y2=4.495
r166 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=3.615 //y=4.58 //x2=3.42 //y2=4.58
r167 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.615 //y=2.08 //x2=3.7 //y2=2.165
r168 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.615 //y=2.08 //x2=3.415 //y2=2.08
r169 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.335 //y=4.665 //x2=3.42 //y2=4.58
r170 (  11 64 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=3.335 //y=4.665 //x2=3.335 //y2=5.725
r171 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.33 //y=1.995 //x2=3.415 //y2=2.08
r172 (  7 62 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=3.33 //y=1.995 //x2=3.33 //y2=1.005
r173 (  6 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.55 //y=3.7 //x2=5.55 //y2=3.7
r174 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=3.7 \
 //y=3.7 //x2=3.7 //y2=3.7
r175 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.815 //y=3.7 //x2=3.7 //y2=3.7
r176 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.435 //y=3.7 //x2=5.55 //y2=3.7
r177 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=5.435 //y=3.7 //x2=3.815 //y2=3.7
ends PM_DLATCHN\%noxref_3

subckt PM_DLATCHN\%noxref_4 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 48 \
 52 53 54 56 62 63 65 73 75 76 )
c134 ( 76 0 ) capacitor c=0.0220291f //x=6.405 //y=5.02
c135 ( 75 0 ) capacitor c=0.0217503f //x=5.525 //y=5.02
c136 ( 73 0 ) capacitor c=0.0084702f //x=6.4 //y=0.905
c137 ( 65 0 ) capacitor c=0.0511458f //x=8.51 //y=2.085
c138 ( 63 0 ) capacitor c=0.0435629f //x=9.15 //y=1.255
c139 ( 62 0 ) capacitor c=0.0200386f //x=9.15 //y=0.91
c140 ( 56 0 ) capacitor c=0.0152946f //x=8.995 //y=1.41
c141 ( 54 0 ) capacitor c=0.0157804f //x=8.995 //y=0.755
c142 ( 53 0 ) capacitor c=0.0490829f //x=8.74 //y=4.79
c143 ( 52 0 ) capacitor c=0.0303096f //x=9.03 //y=4.79
c144 ( 48 0 ) capacitor c=0.0290017f //x=8.62 //y=1.92
c145 ( 47 0 ) capacitor c=0.0250027f //x=8.62 //y=1.565
c146 ( 46 0 ) capacitor c=0.0234316f //x=8.62 //y=1.255
c147 ( 45 0 ) capacitor c=0.0200596f //x=8.62 //y=0.91
c148 ( 44 0 ) capacitor c=0.154218f //x=9.105 //y=6.02
c149 ( 43 0 ) capacitor c=0.154243f //x=8.665 //y=6.02
c150 ( 41 0 ) capacitor c=0.0023043f //x=6.55 //y=5.2
c151 ( 34 0 ) capacitor c=0.0884603f //x=8.51 //y=2.085
c152 ( 32 0 ) capacitor c=0.10682f //x=7.03 //y=3.33
c153 ( 28 0 ) capacitor c=0.00468667f //x=6.675 //y=1.655
c154 ( 27 0 ) capacitor c=0.0131863f //x=6.945 //y=1.655
c155 ( 25 0 ) capacitor c=0.0141863f //x=6.945 //y=5.2
c156 ( 14 0 ) capacitor c=0.00265825f //x=5.755 //y=5.2
c157 ( 13 0 ) capacitor c=0.0149089f //x=6.465 //y=5.2
c158 ( 2 0 ) capacitor c=0.0120846f //x=7.145 //y=3.33
c159 ( 1 0 ) capacitor c=0.0361557f //x=8.395 //y=3.33
r160 (  65 66 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.51 //y=2.085 //x2=8.62 //y2=2.085
r161 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.15 //y=1.255 //x2=9.11 //y2=1.41
r162 (  62 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.15 //y=0.91 //x2=9.11 //y2=0.755
r163 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.15 //y=0.91 //x2=9.15 //y2=1.255
r164 (  57 70 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.775 //y=1.41 //x2=8.66 //y2=1.41
r165 (  56 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.995 //y=1.41 //x2=9.11 //y2=1.41
r166 (  55 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.775 //y=0.755 //x2=8.66 //y2=0.755
r167 (  54 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.995 //y=0.755 //x2=9.11 //y2=0.755
r168 (  54 55 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=8.995 //y=0.755 //x2=8.775 //y2=0.755
r169 (  52 59 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=9.03 //y=4.79 //x2=9.105 //y2=4.865
r170 (  52 53 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=9.03 //y=4.79 //x2=8.74 //y2=4.79
r171 (  49 53 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=8.665 //y=4.865 //x2=8.74 //y2=4.79
r172 (  49 68 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=8.665 //y=4.865 //x2=8.51 //y2=4.7
r173 (  48 66 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=8.62 //y=1.92 //x2=8.62 //y2=2.085
r174 (  47 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.62 //y=1.565 //x2=8.66 //y2=1.41
r175 (  47 48 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=8.62 //y=1.565 //x2=8.62 //y2=1.92
r176 (  46 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.62 //y=1.255 //x2=8.66 //y2=1.41
r177 (  45 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.62 //y=0.91 //x2=8.66 //y2=0.755
r178 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.62 //y=0.91 //x2=8.62 //y2=1.255
r179 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.105 //y=6.02 //x2=9.105 //y2=4.865
r180 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.665 //y=6.02 //x2=8.665 //y2=4.865
r181 (  42 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.885 //y=1.41 //x2=8.995 //y2=1.41
r182 (  42 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.885 //y=1.41 //x2=8.775 //y2=1.41
r183 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.51 //y=4.7 //x2=8.51 //y2=4.7
r184 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=8.51 //y=3.33 //x2=8.51 //y2=4.7
r185 (  34 65 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.51 //y=2.085 //x2=8.51 //y2=2.085
r186 (  34 37 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=8.51 //y=2.085 //x2=8.51 //y2=3.33
r187 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=7.03 //y=5.115 //x2=7.03 //y2=3.33
r188 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=7.03 //y=1.74 //x2=7.03 //y2=3.33
r189 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.945 //y=1.655 //x2=7.03 //y2=1.74
r190 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=6.945 //y=1.655 //x2=6.675 //y2=1.655
r191 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.635 //y=5.2 //x2=6.55 //y2=5.2
r192 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.945 //y=5.2 //x2=7.03 //y2=5.115
r193 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=6.945 //y=5.2 //x2=6.635 //y2=5.2
r194 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.59 //y=1.57 //x2=6.675 //y2=1.655
r195 (  21 73 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=6.59 //y=1.57 //x2=6.59 //y2=1
r196 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.55 //y=5.285 //x2=6.55 //y2=5.2
r197 (  15 76 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=6.55 //y=5.285 //x2=6.55 //y2=5.725
r198 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.465 //y=5.2 //x2=6.55 //y2=5.2
r199 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=6.465 //y=5.2 //x2=5.755 //y2=5.2
r200 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5.67 //y=5.285 //x2=5.755 //y2=5.2
r201 (  7 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=5.67 //y=5.285 //x2=5.67 //y2=5.725
r202 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.51 //y=3.33 //x2=8.51 //y2=3.33
r203 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.03 //y=3.33 //x2=7.03 //y2=3.33
r204 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.145 //y=3.33 //x2=7.03 //y2=3.33
r205 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.395 //y=3.33 //x2=8.51 //y2=3.33
r206 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=8.395 //y=3.33 //x2=7.145 //y2=3.33
ends PM_DLATCHN\%noxref_4

subckt PM_DLATCHN\%noxref_5 ( 1 2 3 4 21 22 23 24 28 29 31 36 45 46 47 48 49 \
 50 51 52 53 58 60 62 68 69 70 71 72 73 77 79 82 83 88 89 92 106 109 111 )
c238 ( 111 0 ) capacitor c=0.028734f //x=0.97 //y=5.02
c239 ( 109 0 ) capacitor c=0.0173218f //x=0.925 //y=0.91
c240 ( 106 0 ) capacitor c=0.0593152f //x=11.1 //y=4.7
c241 ( 92 0 ) capacitor c=0.0331552f //x=6.32 //y=4.7
c242 ( 89 0 ) capacitor c=0.0279499f //x=6.29 //y=1.915
c243 ( 88 0 ) capacitor c=0.0422509f //x=6.29 //y=2.08
c244 ( 83 0 ) capacitor c=0.0318948f //x=11.435 //y=1.21
c245 ( 82 0 ) capacitor c=0.0187384f //x=11.435 //y=0.865
c246 ( 79 0 ) capacitor c=0.0141798f //x=11.28 //y=1.365
c247 ( 77 0 ) capacitor c=0.0149844f //x=11.28 //y=0.71
c248 ( 73 0 ) capacitor c=0.0819722f //x=10.905 //y=1.915
c249 ( 72 0 ) capacitor c=0.0229722f //x=10.905 //y=1.52
c250 ( 71 0 ) capacitor c=0.0234352f //x=10.905 //y=1.21
c251 ( 70 0 ) capacitor c=0.0199343f //x=10.905 //y=0.865
c252 ( 69 0 ) capacitor c=0.0429696f //x=6.855 //y=1.25
c253 ( 68 0 ) capacitor c=0.0192208f //x=6.855 //y=0.905
c254 ( 62 0 ) capacitor c=0.0158629f //x=6.7 //y=1.405
c255 ( 60 0 ) capacitor c=0.0157803f //x=6.7 //y=0.75
c256 ( 58 0 ) capacitor c=0.0300505f //x=6.695 //y=4.79
c257 ( 53 0 ) capacitor c=0.0205163f //x=6.325 //y=1.56
c258 ( 52 0 ) capacitor c=0.0168481f //x=6.325 //y=1.25
c259 ( 51 0 ) capacitor c=0.0174783f //x=6.325 //y=0.905
c260 ( 50 0 ) capacitor c=0.110275f //x=11.44 //y=6.02
c261 ( 49 0 ) capacitor c=0.154305f //x=11 //y=6.02
c262 ( 48 0 ) capacitor c=0.15358f //x=6.77 //y=6.02
c263 ( 47 0 ) capacitor c=0.110281f //x=6.33 //y=6.02
c264 ( 36 0 ) capacitor c=0.0925986f //x=11.1 //y=2.08
c265 ( 31 0 ) capacitor c=0.0756836f //x=6.29 //y=2.08
c266 ( 29 0 ) capacitor c=0.00453889f //x=6.29 //y=4.535
c267 ( 28 0 ) capacitor c=0.0850308f //x=1.48 //y=2.96
c268 ( 24 0 ) capacitor c=0.00575887f //x=1.2 //y=4.58
c269 ( 23 0 ) capacitor c=0.0136332f //x=1.395 //y=4.58
c270 ( 22 0 ) capacitor c=0.00636159f //x=1.195 //y=2.08
c271 ( 21 0 ) capacitor c=0.0137907f //x=1.395 //y=2.08
c272 ( 4 0 ) capacitor c=0.00779117f //x=6.405 //y=2.96
c273 ( 3 0 ) capacitor c=0.14924f //x=10.985 //y=2.96
c274 ( 2 0 ) capacitor c=0.0176065f //x=1.595 //y=2.96
c275 ( 1 0 ) capacitor c=0.158168f //x=6.175 //y=2.96
r276 (  104 106 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=11 //y=4.7 //x2=11.1 //y2=4.7
r277 (  94 95 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=6.32 //y=4.79 //x2=6.32 //y2=4.865
r278 (  92 94 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=6.32 //y=4.7 //x2=6.32 //y2=4.79
r279 (  88 89 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.29 //y=2.08 //x2=6.29 //y2=1.915
r280 (  84 106 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=11.44 //y=4.865 //x2=11.1 //y2=4.7
r281 (  83 108 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.435 //y=1.21 //x2=11.395 //y2=1.365
r282 (  82 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.435 //y=0.865 //x2=11.395 //y2=0.71
r283 (  82 83 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.435 //y=0.865 //x2=11.435 //y2=1.21
r284 (  80 103 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.06 //y=1.365 //x2=10.945 //y2=1.365
r285 (  79 108 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.28 //y=1.365 //x2=11.395 //y2=1.365
r286 (  78 102 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.06 //y=0.71 //x2=10.945 //y2=0.71
r287 (  77 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.28 //y=0.71 //x2=11.395 //y2=0.71
r288 (  77 78 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=11.28 //y=0.71 //x2=11.06 //y2=0.71
r289 (  74 104 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=11 //y=4.865 //x2=11 //y2=4.7
r290 (  73 101 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=10.905 //y=1.915 //x2=11.1 //y2=2.08
r291 (  72 103 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.905 //y=1.52 //x2=10.945 //y2=1.365
r292 (  72 73 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=10.905 //y=1.52 //x2=10.905 //y2=1.915
r293 (  71 103 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.905 //y=1.21 //x2=10.945 //y2=1.365
r294 (  70 102 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.905 //y=0.865 //x2=10.945 //y2=0.71
r295 (  70 71 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.905 //y=0.865 //x2=10.905 //y2=1.21
r296 (  69 99 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.855 //y=1.25 //x2=6.815 //y2=1.405
r297 (  68 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.855 //y=0.905 //x2=6.815 //y2=0.75
r298 (  68 69 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.855 //y=0.905 //x2=6.855 //y2=1.25
r299 (  63 97 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.48 //y=1.405 //x2=6.365 //y2=1.405
r300 (  62 99 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.7 //y=1.405 //x2=6.815 //y2=1.405
r301 (  61 96 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.48 //y=0.75 //x2=6.365 //y2=0.75
r302 (  60 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.7 //y=0.75 //x2=6.815 //y2=0.75
r303 (  60 61 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=6.7 //y=0.75 //x2=6.48 //y2=0.75
r304 (  59 94 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=6.455 //y=4.79 //x2=6.32 //y2=4.79
r305 (  58 65 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.695 //y=4.79 //x2=6.77 //y2=4.865
r306 (  58 59 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=6.695 //y=4.79 //x2=6.455 //y2=4.79
r307 (  53 97 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.325 //y=1.56 //x2=6.365 //y2=1.405
r308 (  53 89 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=6.325 //y=1.56 //x2=6.325 //y2=1.915
r309 (  52 97 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.325 //y=1.25 //x2=6.365 //y2=1.405
r310 (  51 96 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.325 //y=0.905 //x2=6.365 //y2=0.75
r311 (  51 52 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.325 //y=0.905 //x2=6.325 //y2=1.25
r312 (  50 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.44 //y=6.02 //x2=11.44 //y2=4.865
r313 (  49 74 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11 //y=6.02 //x2=11 //y2=4.865
r314 (  48 65 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.77 //y=6.02 //x2=6.77 //y2=4.865
r315 (  47 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.33 //y=6.02 //x2=6.33 //y2=4.865
r316 (  46 79 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.17 //y=1.365 //x2=11.28 //y2=1.365
r317 (  46 80 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.17 //y=1.365 //x2=11.06 //y2=1.365
r318 (  45 62 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.59 //y=1.405 //x2=6.7 //y2=1.405
r319 (  45 63 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.59 //y=1.405 //x2=6.48 //y2=1.405
r320 (  44 92 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.32 //y=4.7 //x2=6.32 //y2=4.7
r321 (  41 106 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.1 //y=4.7 //x2=11.1 //y2=4.7
r322 (  39 41 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=11.1 //y=2.96 //x2=11.1 //y2=4.7
r323 (  36 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.1 //y=2.08 //x2=11.1 //y2=2.08
r324 (  36 39 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=11.1 //y=2.08 //x2=11.1 //y2=2.96
r325 (  31 88 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.29 //y=2.08 //x2=6.29 //y2=2.08
r326 (  31 34 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=6.29 //y=2.08 //x2=6.29 //y2=2.96
r327 (  29 44 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=6.29 //y=4.535 //x2=6.305 //y2=4.7
r328 (  29 34 ) resistor r=107.807 //w=0.187 //l=1.575 //layer=li \
 //thickness=0.1 //x=6.29 //y=4.535 //x2=6.29 //y2=2.96
r329 (  26 28 ) resistor r=105.07 //w=0.187 //l=1.535 //layer=li \
 //thickness=0.1 //x=1.48 //y=4.495 //x2=1.48 //y2=2.96
r330 (  25 28 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=1.48 //y=2.165 //x2=1.48 //y2=2.96
r331 (  23 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.48 //y2=4.495
r332 (  23 24 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.2 //y2=4.58
r333 (  21 25 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.48 //y2=2.165
r334 (  21 22 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.195 //y2=2.08
r335 (  15 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.2 //y2=4.58
r336 (  15 111 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.115 //y2=5.725
r337 (  11 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.195 //y2=2.08
r338 (  11 109 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.11 //y2=1.005
r339 (  10 39 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.1 //y=2.96 //x2=11.1 //y2=2.96
r340 (  8 34 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.29 //y=2.96 //x2=6.29 //y2=2.96
r341 (  6 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.48 //y=2.96 //x2=1.48 //y2=2.96
r342 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.405 //y=2.96 //x2=6.29 //y2=2.96
r343 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.985 //y=2.96 //x2=11.1 //y2=2.96
r344 (  3 4 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=10.985 //y=2.96 //x2=6.405 //y2=2.96
r345 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.595 //y=2.96 //x2=1.48 //y2=2.96
r346 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.175 //y=2.96 //x2=6.29 //y2=2.96
r347 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=6.175 //y=2.96 //x2=1.595 //y2=2.96
ends PM_DLATCHN\%noxref_5

subckt PM_DLATCHN\%D ( 1 2 7 8 9 10 11 12 13 14 15 16 18 29 31 41 42 43 44 45 \
 46 47 48 49 50 54 55 56 58 64 65 66 67 68 73 75 77 83 84 86 95 96 99 )
c179 ( 99 0 ) capacitor c=0.0331844f //x=11.87 //y=4.7
c180 ( 96 0 ) capacitor c=0.0279499f //x=11.84 //y=1.915
c181 ( 95 0 ) capacitor c=0.0437302f //x=11.84 //y=2.08
c182 ( 86 0 ) capacitor c=0.0511458f //x=2.96 //y=2.085
c183 ( 84 0 ) capacitor c=0.0429696f //x=12.405 //y=1.25
c184 ( 83 0 ) capacitor c=0.0192208f //x=12.405 //y=0.905
c185 ( 77 0 ) capacitor c=0.0158629f //x=12.25 //y=1.405
c186 ( 75 0 ) capacitor c=0.0157803f //x=12.25 //y=0.75
c187 ( 73 0 ) capacitor c=0.0307199f //x=12.245 //y=4.79
c188 ( 68 0 ) capacitor c=0.0205163f //x=11.875 //y=1.56
c189 ( 67 0 ) capacitor c=0.0168481f //x=11.875 //y=1.25
c190 ( 66 0 ) capacitor c=0.0174783f //x=11.875 //y=0.905
c191 ( 65 0 ) capacitor c=0.0435629f //x=3.6 //y=1.255
c192 ( 64 0 ) capacitor c=0.0200386f //x=3.6 //y=0.91
c193 ( 58 0 ) capacitor c=0.0152946f //x=3.445 //y=1.41
c194 ( 56 0 ) capacitor c=0.0157804f //x=3.445 //y=0.755
c195 ( 55 0 ) capacitor c=0.0490957f //x=3.19 //y=4.79
c196 ( 54 0 ) capacitor c=0.0303096f //x=3.48 //y=4.79
c197 ( 50 0 ) capacitor c=0.0290017f //x=3.07 //y=1.92
c198 ( 49 0 ) capacitor c=0.0250027f //x=3.07 //y=1.565
c199 ( 48 0 ) capacitor c=0.0234316f //x=3.07 //y=1.255
c200 ( 47 0 ) capacitor c=0.0200596f //x=3.07 //y=0.91
c201 ( 46 0 ) capacitor c=0.15358f //x=12.32 //y=6.02
c202 ( 45 0 ) capacitor c=0.110281f //x=11.88 //y=6.02
c203 ( 44 0 ) capacitor c=0.154218f //x=3.555 //y=6.02
c204 ( 43 0 ) capacitor c=0.154243f //x=3.115 //y=6.02
c205 ( 31 0 ) capacitor c=0.0762219f //x=11.84 //y=2.08
c206 ( 29 0 ) capacitor c=0.00453889f //x=11.84 //y=4.535
c207 ( 18 0 ) capacitor c=0.0910566f //x=2.96 //y=2.085
c208 ( 2 0 ) capacitor c=0.0168127f //x=3.075 //y=4.07
c209 ( 1 0 ) capacitor c=0.246212f //x=11.725 //y=4.07
r210 (  101 102 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=11.87 //y=4.79 //x2=11.87 //y2=4.865
r211 (  99 101 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=11.87 //y=4.7 //x2=11.87 //y2=4.79
r212 (  95 96 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=11.84 //y=2.08 //x2=11.84 //y2=1.915
r213 (  86 87 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.96 //y=2.085 //x2=3.07 //y2=2.085
r214 (  84 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.405 //y=1.25 //x2=12.365 //y2=1.405
r215 (  83 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.405 //y=0.905 //x2=12.365 //y2=0.75
r216 (  83 84 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.405 //y=0.905 //x2=12.405 //y2=1.25
r217 (  78 104 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.03 //y=1.405 //x2=11.915 //y2=1.405
r218 (  77 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.25 //y=1.405 //x2=12.365 //y2=1.405
r219 (  76 103 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.03 //y=0.75 //x2=11.915 //y2=0.75
r220 (  75 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.25 //y=0.75 //x2=12.365 //y2=0.75
r221 (  75 76 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=12.25 //y=0.75 //x2=12.03 //y2=0.75
r222 (  74 101 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=12.005 //y=4.79 //x2=11.87 //y2=4.79
r223 (  73 80 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=12.245 //y=4.79 //x2=12.32 //y2=4.865
r224 (  73 74 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=12.245 //y=4.79 //x2=12.005 //y2=4.79
r225 (  68 104 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.875 //y=1.56 //x2=11.915 //y2=1.405
r226 (  68 96 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=11.875 //y=1.56 //x2=11.875 //y2=1.915
r227 (  67 104 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.875 //y=1.25 //x2=11.915 //y2=1.405
r228 (  66 103 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.875 //y=0.905 //x2=11.915 //y2=0.75
r229 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.875 //y=0.905 //x2=11.875 //y2=1.25
r230 (  65 93 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.6 //y=1.255 //x2=3.56 //y2=1.41
r231 (  64 92 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.6 //y=0.91 //x2=3.56 //y2=0.755
r232 (  64 65 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.6 //y=0.91 //x2=3.6 //y2=1.255
r233 (  59 91 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.225 //y=1.41 //x2=3.11 //y2=1.41
r234 (  58 93 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.445 //y=1.41 //x2=3.56 //y2=1.41
r235 (  57 90 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.225 //y=0.755 //x2=3.11 //y2=0.755
r236 (  56 92 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.445 //y=0.755 //x2=3.56 //y2=0.755
r237 (  56 57 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.445 //y=0.755 //x2=3.225 //y2=0.755
r238 (  54 61 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=3.48 //y=4.79 //x2=3.555 //y2=4.865
r239 (  54 55 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=3.48 //y=4.79 //x2=3.19 //y2=4.79
r240 (  51 55 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=3.115 //y=4.865 //x2=3.19 //y2=4.79
r241 (  51 89 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=3.115 //y=4.865 //x2=2.96 //y2=4.7
r242 (  50 87 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.07 //y=1.92 //x2=3.07 //y2=2.085
r243 (  49 91 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.07 //y=1.565 //x2=3.11 //y2=1.41
r244 (  49 50 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=3.07 //y=1.565 //x2=3.07 //y2=1.92
r245 (  48 91 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.07 //y=1.255 //x2=3.11 //y2=1.41
r246 (  47 90 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.07 //y=0.91 //x2=3.11 //y2=0.755
r247 (  47 48 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.07 //y=0.91 //x2=3.07 //y2=1.255
r248 (  46 80 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.32 //y=6.02 //x2=12.32 //y2=4.865
r249 (  45 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.88 //y=6.02 //x2=11.88 //y2=4.865
r250 (  44 61 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.555 //y=6.02 //x2=3.555 //y2=4.865
r251 (  43 51 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.115 //y=6.02 //x2=3.115 //y2=4.865
r252 (  42 77 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.14 //y=1.405 //x2=12.25 //y2=1.405
r253 (  42 78 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.14 //y=1.405 //x2=12.03 //y2=1.405
r254 (  41 58 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.335 //y=1.41 //x2=3.445 //y2=1.41
r255 (  41 59 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.335 //y=1.41 //x2=3.225 //y2=1.41
r256 (  40 99 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.87 //y=4.7 //x2=11.87 //y2=4.7
r257 (  31 95 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=2.08 //x2=11.84 //y2=2.08
r258 (  29 40 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=11.84 //y=4.535 //x2=11.855 //y2=4.7
r259 (  27 89 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.96 //y=4.7 //x2=2.96 //y2=4.7
r260 (  18 86 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.96 //y=2.085 //x2=2.96 //y2=2.085
r261 (  16 29 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=11.84 //y=4.44 //x2=11.84 //y2=4.535
r262 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=11.84 //y=4.07 //x2=11.84 //y2=4.44
r263 (  14 15 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=11.84 //y=3.33 //x2=11.84 //y2=4.07
r264 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.96 //x2=11.84 //y2=3.33
r265 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.59 //x2=11.84 //y2=2.96
r266 (  12 31 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.59 //x2=11.84 //y2=2.08
r267 (  11 27 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=2.96 //y=4.44 //x2=2.96 //y2=4.7
r268 (  10 11 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.96 //y=4.07 //x2=2.96 //y2=4.44
r269 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.96 //y=3.7 //x2=2.96 //y2=4.07
r270 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=2.96 //y=3.33 //x2=2.96 //y2=3.7
r271 (  7 8 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li //thickness=0.1 \
 //x=2.96 //y=2.59 //x2=2.96 //y2=3.33
r272 (  7 18 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=2.96 //y=2.59 //x2=2.96 //y2=2.085
r273 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.84 //y=4.07 //x2=11.84 //y2=4.07
r274 (  4 10 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.96 //y=4.07 //x2=2.96 //y2=4.07
r275 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.075 //y=4.07 //x2=2.96 //y2=4.07
r276 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.725 //y=4.07 //x2=11.84 //y2=4.07
r277 (  1 2 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=11.725 //y=4.07 //x2=3.075 //y2=4.07
ends PM_DLATCHN\%D

subckt PM_DLATCHN\%noxref_7 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 48 \
 52 53 54 56 62 63 65 73 75 76 )
c139 ( 76 0 ) capacitor c=0.0220291f //x=11.955 //y=5.02
c140 ( 75 0 ) capacitor c=0.0217503f //x=11.075 //y=5.02
c141 ( 73 0 ) capacitor c=0.0084702f //x=11.95 //y=0.905
c142 ( 65 0 ) capacitor c=0.0528806f //x=14.06 //y=2.085
c143 ( 63 0 ) capacitor c=0.0435629f //x=14.7 //y=1.255
c144 ( 62 0 ) capacitor c=0.0200386f //x=14.7 //y=0.91
c145 ( 56 0 ) capacitor c=0.0152946f //x=14.545 //y=1.41
c146 ( 54 0 ) capacitor c=0.0157804f //x=14.545 //y=0.755
c147 ( 53 0 ) capacitor c=0.0493989f //x=14.29 //y=4.79
c148 ( 52 0 ) capacitor c=0.0304843f //x=14.58 //y=4.79
c149 ( 48 0 ) capacitor c=0.0290017f //x=14.17 //y=1.92
c150 ( 47 0 ) capacitor c=0.0250027f //x=14.17 //y=1.565
c151 ( 46 0 ) capacitor c=0.0234316f //x=14.17 //y=1.255
c152 ( 45 0 ) capacitor c=0.0200596f //x=14.17 //y=0.91
c153 ( 44 0 ) capacitor c=0.154218f //x=14.655 //y=6.02
c154 ( 43 0 ) capacitor c=0.154243f //x=14.215 //y=6.02
c155 ( 41 0 ) capacitor c=0.0024826f //x=12.1 //y=5.2
c156 ( 34 0 ) capacitor c=0.0908493f //x=14.06 //y=2.085
c157 ( 32 0 ) capacitor c=0.108527f //x=12.58 //y=3.33
c158 ( 28 0 ) capacitor c=0.00525782f //x=12.225 //y=1.655
c159 ( 27 0 ) capacitor c=0.0139525f //x=12.495 //y=1.655
c160 ( 25 0 ) capacitor c=0.0144648f //x=12.495 //y=5.2
c161 ( 14 0 ) capacitor c=0.00265825f //x=11.305 //y=5.2
c162 ( 13 0 ) capacitor c=0.0150834f //x=12.015 //y=5.2
c163 ( 2 0 ) capacitor c=0.0111324f //x=12.695 //y=3.33
c164 ( 1 0 ) capacitor c=0.0522233f //x=13.945 //y=3.33
r165 (  65 66 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.06 //y=2.085 //x2=14.17 //y2=2.085
r166 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.7 //y=1.255 //x2=14.66 //y2=1.41
r167 (  62 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.7 //y=0.91 //x2=14.66 //y2=0.755
r168 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.7 //y=0.91 //x2=14.7 //y2=1.255
r169 (  57 70 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.325 //y=1.41 //x2=14.21 //y2=1.41
r170 (  56 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.545 //y=1.41 //x2=14.66 //y2=1.41
r171 (  55 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.325 //y=0.755 //x2=14.21 //y2=0.755
r172 (  54 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.545 //y=0.755 //x2=14.66 //y2=0.755
r173 (  54 55 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=14.545 //y=0.755 //x2=14.325 //y2=0.755
r174 (  52 59 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=14.58 //y=4.79 //x2=14.655 //y2=4.865
r175 (  52 53 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=14.58 //y=4.79 //x2=14.29 //y2=4.79
r176 (  49 53 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=14.215 //y=4.865 //x2=14.29 //y2=4.79
r177 (  49 68 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=14.215 //y=4.865 //x2=14.06 //y2=4.7
r178 (  48 66 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=14.17 //y=1.92 //x2=14.17 //y2=2.085
r179 (  47 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.17 //y=1.565 //x2=14.21 //y2=1.41
r180 (  47 48 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=14.17 //y=1.565 //x2=14.17 //y2=1.92
r181 (  46 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.17 //y=1.255 //x2=14.21 //y2=1.41
r182 (  45 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.17 //y=0.91 //x2=14.21 //y2=0.755
r183 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.17 //y=0.91 //x2=14.17 //y2=1.255
r184 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.655 //y=6.02 //x2=14.655 //y2=4.865
r185 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.215 //y=6.02 //x2=14.215 //y2=4.865
r186 (  42 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.435 //y=1.41 //x2=14.545 //y2=1.41
r187 (  42 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.435 //y=1.41 //x2=14.325 //y2=1.41
r188 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=4.7 //x2=14.06 //y2=4.7
r189 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=14.06 //y=3.33 //x2=14.06 //y2=4.7
r190 (  34 65 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=2.085 //x2=14.06 //y2=2.085
r191 (  34 37 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=14.06 //y=2.085 //x2=14.06 //y2=3.33
r192 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=12.58 //y=5.115 //x2=12.58 //y2=3.33
r193 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=12.58 //y=1.74 //x2=12.58 //y2=3.33
r194 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.495 //y=1.655 //x2=12.58 //y2=1.74
r195 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=12.495 //y=1.655 //x2=12.225 //y2=1.655
r196 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.185 //y=5.2 //x2=12.1 //y2=5.2
r197 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.495 //y=5.2 //x2=12.58 //y2=5.115
r198 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=12.495 //y=5.2 //x2=12.185 //y2=5.2
r199 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.14 //y=1.57 //x2=12.225 //y2=1.655
r200 (  21 73 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=12.14 //y=1.57 //x2=12.14 //y2=1
r201 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.1 //y=5.285 //x2=12.1 //y2=5.2
r202 (  15 76 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=12.1 //y=5.285 //x2=12.1 //y2=5.725
r203 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.015 //y=5.2 //x2=12.1 //y2=5.2
r204 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=12.015 //y=5.2 //x2=11.305 //y2=5.2
r205 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.22 //y=5.285 //x2=11.305 //y2=5.2
r206 (  7 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=11.22 //y=5.285 //x2=11.22 //y2=5.725
r207 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.06 //y=3.33 //x2=14.06 //y2=3.33
r208 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.58 //y=3.33 //x2=12.58 //y2=3.33
r209 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.695 //y=3.33 //x2=12.58 //y2=3.33
r210 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=3.33 //x2=14.06 //y2=3.33
r211 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=3.33 //x2=12.695 //y2=3.33
ends PM_DLATCHN\%noxref_7

subckt PM_DLATCHN\%noxref_8 ( 1 2 17 18 19 20 24 27 32 34 35 36 37 38 39 40 44 \
 46 49 51 52 57 67 69 )
c164 ( 69 0 ) capacitor c=0.0288745f //x=8.74 //y=5.02
c165 ( 67 0 ) capacitor c=0.0173218f //x=8.695 //y=0.91
c166 ( 57 0 ) capacitor c=0.0403405f //x=16.495 //y=4.705
c167 ( 52 0 ) capacitor c=0.0321911f //x=16.985 //y=1.25
c168 ( 51 0 ) capacitor c=0.0185201f //x=16.985 //y=0.905
c169 ( 49 0 ) capacitor c=0.0288104f //x=16.915 //y=4.795
c170 ( 46 0 ) capacitor c=0.0133656f //x=16.83 //y=1.405
c171 ( 44 0 ) capacitor c=0.0157804f //x=16.83 //y=0.75
c172 ( 40 0 ) capacitor c=0.0828832f //x=16.455 //y=1.915
c173 ( 39 0 ) capacitor c=0.022867f //x=16.455 //y=1.56
c174 ( 38 0 ) capacitor c=0.0234318f //x=16.455 //y=1.25
c175 ( 37 0 ) capacitor c=0.0192004f //x=16.455 //y=0.905
c176 ( 36 0 ) capacitor c=0.110795f //x=16.99 //y=6.025
c177 ( 35 0 ) capacitor c=0.153847f //x=16.55 //y=6.025
c178 ( 32 0 ) capacitor c=0.00993392f //x=16.495 //y=4.705
c179 ( 27 0 ) capacitor c=0.0921227f //x=16.65 //y=2.08
c180 ( 24 0 ) capacitor c=0.0820607f //x=9.25 //y=3.7
c181 ( 20 0 ) capacitor c=0.00417404f //x=8.97 //y=4.58
c182 ( 19 0 ) capacitor c=0.0118896f //x=9.165 //y=4.58
c183 ( 18 0 ) capacitor c=0.00549299f //x=8.965 //y=2.08
c184 ( 17 0 ) capacitor c=0.013178f //x=9.165 //y=2.08
c185 ( 2 0 ) capacitor c=0.0108199f //x=9.365 //y=3.7
c186 ( 1 0 ) capacitor c=0.214055f //x=16.535 //y=3.7
r187 (  59 60 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=16.495 //y=4.795 //x2=16.495 //y2=4.87
r188 (  57 59 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=16.495 //y=4.705 //x2=16.495 //y2=4.795
r189 (  52 66 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.985 //y=1.25 //x2=16.945 //y2=1.405
r190 (  51 65 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.985 //y=0.905 //x2=16.945 //y2=0.75
r191 (  51 52 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.985 //y=0.905 //x2=16.985 //y2=1.25
r192 (  50 59 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=16.63 //y=4.795 //x2=16.495 //y2=4.795
r193 (  49 53 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=16.915 //y=4.795 //x2=16.99 //y2=4.87
r194 (  49 50 ) resistor r=146.138 //w=0.094 //l=0.285 //layer=ply \
 //thickness=0.18 //x=16.915 //y=4.795 //x2=16.63 //y2=4.795
r195 (  47 64 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.61 //y=1.405 //x2=16.495 //y2=1.405
r196 (  46 66 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.83 //y=1.405 //x2=16.945 //y2=1.405
r197 (  45 63 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.61 //y=0.75 //x2=16.495 //y2=0.75
r198 (  44 65 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.83 //y=0.75 //x2=16.945 //y2=0.75
r199 (  44 45 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=16.83 //y=0.75 //x2=16.61 //y2=0.75
r200 (  40 62 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=16.455 //y=1.915 //x2=16.65 //y2=2.08
r201 (  39 64 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.455 //y=1.56 //x2=16.495 //y2=1.405
r202 (  39 40 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=16.455 //y=1.56 //x2=16.455 //y2=1.915
r203 (  38 64 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.455 //y=1.25 //x2=16.495 //y2=1.405
r204 (  37 63 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.455 //y=0.905 //x2=16.495 //y2=0.75
r205 (  37 38 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.455 //y=0.905 //x2=16.455 //y2=1.25
r206 (  36 53 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.99 //y=6.025 //x2=16.99 //y2=4.87
r207 (  35 60 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.55 //y=6.025 //x2=16.55 //y2=4.87
r208 (  34 46 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=16.72 //y=1.405 //x2=16.83 //y2=1.405
r209 (  34 47 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=16.72 //y=1.405 //x2=16.61 //y2=1.405
r210 (  32 57 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.495 //y=4.705 //x2=16.495 //y2=4.705
r211 (  32 33 ) resistor r=7.81102 //w=0.254 //l=0.155 //layer=li \
 //thickness=0.1 //x=16.495 //y=4.705 //x2=16.65 //y2=4.705
r212 (  27 62 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.65 //y=2.08 //x2=16.65 //y2=2.08
r213 (  27 30 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=16.65 //y=2.08 //x2=16.65 //y2=3.7
r214 (  25 33 ) resistor r=3.23951 //w=0.254 //l=0.165 //layer=li \
 //thickness=0.1 //x=16.65 //y=4.54 //x2=16.65 //y2=4.705
r215 (  25 30 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=16.65 //y=4.54 //x2=16.65 //y2=3.7
r216 (  22 24 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=9.25 //y=4.495 //x2=9.25 //y2=3.7
r217 (  21 24 ) resistor r=105.07 //w=0.187 //l=1.535 //layer=li \
 //thickness=0.1 //x=9.25 //y=2.165 //x2=9.25 //y2=3.7
r218 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.165 //y=4.58 //x2=9.25 //y2=4.495
r219 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=9.165 //y=4.58 //x2=8.97 //y2=4.58
r220 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.165 //y=2.08 //x2=9.25 //y2=2.165
r221 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=9.165 //y=2.08 //x2=8.965 //y2=2.08
r222 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.885 //y=4.665 //x2=8.97 //y2=4.58
r223 (  11 69 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=8.885 //y=4.665 //x2=8.885 //y2=5.725
r224 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.88 //y=1.995 //x2=8.965 //y2=2.08
r225 (  7 67 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=8.88 //y=1.995 //x2=8.88 //y2=1.005
r226 (  6 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=16.65 //y=3.7 //x2=16.65 //y2=3.7
r227 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.25 //y=3.7 //x2=9.25 //y2=3.7
r228 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.365 //y=3.7 //x2=9.25 //y2=3.7
r229 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.535 //y=3.7 //x2=16.65 //y2=3.7
r230 (  1 2 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=16.535 //y=3.7 //x2=9.365 //y2=3.7
ends PM_DLATCHN\%noxref_8

subckt PM_DLATCHN\%Q ( 1 2 7 8 9 10 11 12 13 14 15 16 21 22 33 34 35 47 57 59 \
 60 61 62 63 64 65 69 71 74 76 77 82 92 93 96 )
c167 ( 96 0 ) capacitor c=0.0159573f //x=17.505 //y=5.025
c168 ( 93 0 ) capacitor c=0.00923651f //x=17.5 //y=0.905
c169 ( 92 0 ) capacitor c=0.007684f //x=16.53 //y=0.905
c170 ( 82 0 ) capacitor c=0.0402699f //x=19.825 //y=4.705
c171 ( 77 0 ) capacitor c=0.0321911f //x=20.315 //y=1.25
c172 ( 76 0 ) capacitor c=0.0185201f //x=20.315 //y=0.905
c173 ( 74 0 ) capacitor c=0.0288104f //x=20.245 //y=4.795
c174 ( 71 0 ) capacitor c=0.0133656f //x=20.16 //y=1.405
c175 ( 69 0 ) capacitor c=0.0157804f //x=20.16 //y=0.75
c176 ( 65 0 ) capacitor c=0.0822075f //x=19.785 //y=1.915
c177 ( 64 0 ) capacitor c=0.022867f //x=19.785 //y=1.56
c178 ( 63 0 ) capacitor c=0.0234318f //x=19.785 //y=1.25
c179 ( 62 0 ) capacitor c=0.0192004f //x=19.785 //y=0.905
c180 ( 61 0 ) capacitor c=0.110795f //x=20.32 //y=6.025
c181 ( 60 0 ) capacitor c=0.153847f //x=19.88 //y=6.025
c182 ( 57 0 ) capacitor c=0.00993392f //x=19.825 //y=4.705
c183 ( 55 0 ) capacitor c=0.00454201f //x=17.69 //y=1.655
c184 ( 47 0 ) capacitor c=0.0893171f //x=19.98 //y=2.08
c185 ( 35 0 ) capacitor c=0.0140918f //x=18.045 //y=1.655
c186 ( 34 0 ) capacitor c=0.00308317f //x=17.735 //y=5.21
c187 ( 33 0 ) capacitor c=0.0137261f //x=18.045 //y=5.21
c188 ( 22 0 ) capacitor c=0.00224268f //x=16.805 //y=1.655
c189 ( 21 0 ) capacitor c=0.0218623f //x=17.605 //y=1.655
c190 ( 7 0 ) capacitor c=0.110461f //x=18.13 //y=2.22
c191 ( 2 0 ) capacitor c=0.0112178f //x=18.245 //y=3.33
c192 ( 1 0 ) capacitor c=0.0678125f //x=19.865 //y=3.33
r193 (  84 85 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=19.825 //y=4.795 //x2=19.825 //y2=4.87
r194 (  82 84 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=19.825 //y=4.705 //x2=19.825 //y2=4.795
r195 (  77 91 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.315 //y=1.25 //x2=20.275 //y2=1.405
r196 (  76 90 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.315 //y=0.905 //x2=20.275 //y2=0.75
r197 (  76 77 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.315 //y=0.905 //x2=20.315 //y2=1.25
r198 (  75 84 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=19.96 //y=4.795 //x2=19.825 //y2=4.795
r199 (  74 78 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.245 //y=4.795 //x2=20.32 //y2=4.87
r200 (  74 75 ) resistor r=146.138 //w=0.094 //l=0.285 //layer=ply \
 //thickness=0.18 //x=20.245 //y=4.795 //x2=19.96 //y2=4.795
r201 (  72 89 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.94 //y=1.405 //x2=19.825 //y2=1.405
r202 (  71 91 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.16 //y=1.405 //x2=20.275 //y2=1.405
r203 (  70 88 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.94 //y=0.75 //x2=19.825 //y2=0.75
r204 (  69 90 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.16 //y=0.75 //x2=20.275 //y2=0.75
r205 (  69 70 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=20.16 //y=0.75 //x2=19.94 //y2=0.75
r206 (  65 87 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=19.785 //y=1.915 //x2=19.98 //y2=2.08
r207 (  64 89 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.785 //y=1.56 //x2=19.825 //y2=1.405
r208 (  64 65 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=19.785 //y=1.56 //x2=19.785 //y2=1.915
r209 (  63 89 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.785 //y=1.25 //x2=19.825 //y2=1.405
r210 (  62 88 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.785 //y=0.905 //x2=19.825 //y2=0.75
r211 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=19.785 //y=0.905 //x2=19.785 //y2=1.25
r212 (  61 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.32 //y=6.025 //x2=20.32 //y2=4.87
r213 (  60 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.88 //y=6.025 //x2=19.88 //y2=4.87
r214 (  59 71 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.405 //x2=20.16 //y2=1.405
r215 (  59 72 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.405 //x2=19.94 //y2=1.405
r216 (  57 82 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.825 //y=4.705 //x2=19.825 //y2=4.705
r217 (  57 58 ) resistor r=7.81102 //w=0.254 //l=0.155 //layer=li \
 //thickness=0.1 //x=19.825 //y=4.705 //x2=19.98 //y2=4.705
r218 (  47 87 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.98 //y=2.08 //x2=19.98 //y2=2.08
r219 (  45 58 ) resistor r=3.23951 //w=0.254 //l=0.165 //layer=li \
 //thickness=0.1 //x=19.98 //y=4.54 //x2=19.98 //y2=4.705
r220 (  36 55 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.775 //y=1.655 //x2=17.69 //y2=1.655
r221 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.045 //y=1.655 //x2=18.13 //y2=1.74
r222 (  35 36 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=18.045 //y=1.655 //x2=17.775 //y2=1.655
r223 (  33 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.045 //y=5.21 //x2=18.13 //y2=5.125
r224 (  33 34 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=18.045 //y=5.21 //x2=17.735 //y2=5.21
r225 (  29 55 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.69 //y=1.57 //x2=17.69 //y2=1.655
r226 (  29 93 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=17.69 //y=1.57 //x2=17.69 //y2=1
r227 (  23 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.65 //y=5.295 //x2=17.735 //y2=5.21
r228 (  23 96 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=17.65 //y=5.295 //x2=17.65 //y2=5.72
r229 (  21 55 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.605 //y=1.655 //x2=17.69 //y2=1.655
r230 (  21 22 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li \
 //thickness=0.1 //x=17.605 //y=1.655 //x2=16.805 //y2=1.655
r231 (  17 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.72 //y=1.57 //x2=16.805 //y2=1.655
r232 (  17 92 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=16.72 //y=1.57 //x2=16.72 //y2=1
r233 (  16 45 ) resistor r=6.84492 //w=0.187 //l=0.1 //layer=li \
 //thickness=0.1 //x=19.98 //y=4.44 //x2=19.98 //y2=4.54
r234 (  15 16 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=19.98 //y=3.33 //x2=19.98 //y2=4.44
r235 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.96 //x2=19.98 //y2=3.33
r236 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.59 //x2=19.98 //y2=2.96
r237 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.22 //x2=19.98 //y2=2.59
r238 (  12 47 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.22 //x2=19.98 //y2=2.08
r239 (  11 38 ) resistor r=46.8877 //w=0.187 //l=0.685 //layer=li \
 //thickness=0.1 //x=18.13 //y=4.44 //x2=18.13 //y2=5.125
r240 (  10 11 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=18.13 //y=3.33 //x2=18.13 //y2=4.44
r241 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=18.13 //y=2.96 //x2=18.13 //y2=3.33
r242 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=18.13 //y=2.59 //x2=18.13 //y2=2.96
r243 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=18.13 //y=2.22 //x2=18.13 //y2=2.59
r244 (  7 37 ) resistor r=32.8556 //w=0.187 //l=0.48 //layer=li \
 //thickness=0.1 //x=18.13 //y=2.22 //x2=18.13 //y2=1.74
r245 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=19.98 //y=3.33 //x2=19.98 //y2=3.33
r246 (  4 10 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.13 //y=3.33 //x2=18.13 //y2=3.33
r247 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.245 //y=3.33 //x2=18.13 //y2=3.33
r248 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=19.865 //y=3.33 //x2=19.98 //y2=3.33
r249 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=19.865 //y=3.33 //x2=18.245 //y2=3.33
ends PM_DLATCHN\%Q

subckt PM_DLATCHN\%noxref_10 ( 1 2 17 18 19 20 24 25 27 33 34 35 36 37 38 43 \
 45 47 53 54 56 57 60 68 70 )
c162 ( 70 0 ) capacitor c=0.028853f //x=14.29 //y=5.02
c163 ( 68 0 ) capacitor c=0.0173218f //x=14.245 //y=0.91
c164 ( 60 0 ) capacitor c=0.0354945f //x=20.755 //y=4.705
c165 ( 57 0 ) capacitor c=0.0279572f //x=20.72 //y=1.915
c166 ( 56 0 ) capacitor c=0.0422144f //x=20.72 //y=2.08
c167 ( 54 0 ) capacitor c=0.0237734f //x=21.285 //y=1.255
c168 ( 53 0 ) capacitor c=0.0191782f //x=21.285 //y=0.905
c169 ( 47 0 ) capacitor c=0.0346941f //x=21.13 //y=1.405
c170 ( 45 0 ) capacitor c=0.0157803f //x=21.13 //y=0.75
c171 ( 43 0 ) capacitor c=0.030194f //x=21.125 //y=4.795
c172 ( 38 0 ) capacitor c=0.0199921f //x=20.755 //y=1.56
c173 ( 37 0 ) capacitor c=0.0169608f //x=20.755 //y=1.255
c174 ( 36 0 ) capacitor c=0.0185462f //x=20.755 //y=0.905
c175 ( 35 0 ) capacitor c=0.15325f //x=21.2 //y=6.025
c176 ( 34 0 ) capacitor c=0.110232f //x=20.76 //y=6.025
c177 ( 27 0 ) capacitor c=0.0760752f //x=20.72 //y=2.08
c178 ( 25 0 ) capacitor c=0.00514985f //x=20.72 //y=4.54
c179 ( 24 0 ) capacitor c=0.0855616f //x=14.8 //y=4.07
c180 ( 20 0 ) capacitor c=0.00497659f //x=14.52 //y=4.58
c181 ( 19 0 ) capacitor c=0.012509f //x=14.715 //y=4.58
c182 ( 18 0 ) capacitor c=0.00612032f //x=14.515 //y=2.08
c183 ( 17 0 ) capacitor c=0.0138937f //x=14.715 //y=2.08
c184 ( 2 0 ) capacitor c=0.0119148f //x=14.915 //y=4.07
c185 ( 1 0 ) capacitor c=0.169542f //x=20.605 //y=4.07
r186 (  62 63 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=20.755 //y=4.795 //x2=20.755 //y2=4.87
r187 (  60 62 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=20.755 //y=4.705 //x2=20.755 //y2=4.795
r188 (  56 57 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=20.72 //y=2.08 //x2=20.72 //y2=1.915
r189 (  54 67 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=21.285 //y=1.255 //x2=21.285 //y2=1.367
r190 (  53 66 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.285 //y=0.905 //x2=21.245 //y2=0.75
r191 (  53 54 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=21.285 //y=0.905 //x2=21.285 //y2=1.255
r192 (  48 65 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.91 //y=1.405 //x2=20.795 //y2=1.405
r193 (  47 67 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=21.13 //y=1.405 //x2=21.285 //y2=1.367
r194 (  46 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.91 //y=0.75 //x2=20.795 //y2=0.75
r195 (  45 66 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.13 //y=0.75 //x2=21.245 //y2=0.75
r196 (  45 46 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=21.13 //y=0.75 //x2=20.91 //y2=0.75
r197 (  44 62 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=20.89 //y=4.795 //x2=20.755 //y2=4.795
r198 (  43 50 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=21.125 //y=4.795 //x2=21.2 //y2=4.87
r199 (  43 44 ) resistor r=120.5 //w=0.094 //l=0.235 //layer=ply \
 //thickness=0.18 //x=21.125 //y=4.795 //x2=20.89 //y2=4.795
r200 (  38 65 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.755 //y=1.56 //x2=20.795 //y2=1.405
r201 (  38 57 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=20.755 //y=1.56 //x2=20.755 //y2=1.915
r202 (  37 65 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=20.755 //y=1.255 //x2=20.795 //y2=1.405
r203 (  36 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.755 //y=0.905 //x2=20.795 //y2=0.75
r204 (  36 37 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=20.755 //y=0.905 //x2=20.755 //y2=1.255
r205 (  35 50 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.2 //y=6.025 //x2=21.2 //y2=4.87
r206 (  34 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.76 //y=6.025 //x2=20.76 //y2=4.87
r207 (  33 47 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=21.02 //y=1.405 //x2=21.13 //y2=1.405
r208 (  33 48 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=21.02 //y=1.405 //x2=20.91 //y2=1.405
r209 (  32 60 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.755 //y=4.705 //x2=20.755 //y2=4.705
r210 (  27 56 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.72 //y=2.08 //x2=20.72 //y2=2.08
r211 (  27 30 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=20.72 //y=2.08 //x2=20.72 //y2=4.07
r212 (  25 32 ) resistor r=11.332 //w=0.189 //l=0.173292 //layer=li \
 //thickness=0.1 //x=20.72 //y=4.54 //x2=20.737 //y2=4.705
r213 (  25 30 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=20.72 //y=4.54 //x2=20.72 //y2=4.07
r214 (  22 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=14.8 //y=4.495 //x2=14.8 //y2=4.07
r215 (  21 24 ) resistor r=130.396 //w=0.187 //l=1.905 //layer=li \
 //thickness=0.1 //x=14.8 //y=2.165 //x2=14.8 //y2=4.07
r216 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.715 //y=4.58 //x2=14.8 //y2=4.495
r217 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=14.715 //y=4.58 //x2=14.52 //y2=4.58
r218 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.715 //y=2.08 //x2=14.8 //y2=2.165
r219 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=14.715 //y=2.08 //x2=14.515 //y2=2.08
r220 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.435 //y=4.665 //x2=14.52 //y2=4.58
r221 (  11 70 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=14.435 //y=4.665 //x2=14.435 //y2=5.725
r222 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.43 //y=1.995 //x2=14.515 //y2=2.08
r223 (  7 68 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=14.43 //y=1.995 //x2=14.43 //y2=1.005
r224 (  6 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=20.72 //y=4.07 //x2=20.72 //y2=4.07
r225 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.8 //y=4.07 //x2=14.8 //y2=4.07
r226 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=14.915 //y=4.07 //x2=14.8 //y2=4.07
r227 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=4.07 //x2=20.72 //y2=4.07
r228 (  1 2 ) resistor r=5.42939 //w=0.131 //l=5.69 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=4.07 //x2=14.915 //y2=4.07
ends PM_DLATCHN\%noxref_10

subckt PM_DLATCHN\%noxref_11 ( 1 2 7 9 17 18 29 30 31 36 40 41 42 43 44 45 50 \
 52 54 60 61 63 64 67 75 76 79 )
c162 ( 79 0 ) capacitor c=0.0159573f //x=20.835 //y=5.025
c163 ( 76 0 ) capacitor c=0.00905936f //x=20.83 //y=0.905
c164 ( 75 0 ) capacitor c=0.007684f //x=19.86 //y=0.905
c165 ( 67 0 ) capacitor c=0.0354569f //x=17.425 //y=4.705
c166 ( 64 0 ) capacitor c=0.0279572f //x=17.39 //y=1.915
c167 ( 63 0 ) capacitor c=0.0422144f //x=17.39 //y=2.08
c168 ( 61 0 ) capacitor c=0.0237734f //x=17.955 //y=1.255
c169 ( 60 0 ) capacitor c=0.0191782f //x=17.955 //y=0.905
c170 ( 54 0 ) capacitor c=0.0346941f //x=17.8 //y=1.405
c171 ( 52 0 ) capacitor c=0.0157803f //x=17.8 //y=0.75
c172 ( 50 0 ) capacitor c=0.0295389f //x=17.795 //y=4.795
c173 ( 45 0 ) capacitor c=0.0199921f //x=17.425 //y=1.56
c174 ( 44 0 ) capacitor c=0.0169608f //x=17.425 //y=1.255
c175 ( 43 0 ) capacitor c=0.0185462f //x=17.425 //y=0.905
c176 ( 42 0 ) capacitor c=0.15325f //x=17.87 //y=6.025
c177 ( 41 0 ) capacitor c=0.110232f //x=17.43 //y=6.025
c178 ( 39 0 ) capacitor c=0.00454201f //x=21.02 //y=1.655
c179 ( 36 0 ) capacitor c=0.128643f //x=21.46 //y=3.7
c180 ( 31 0 ) capacitor c=0.0141769f //x=21.375 //y=1.655
c181 ( 30 0 ) capacitor c=0.00326058f //x=21.065 //y=5.21
c182 ( 29 0 ) capacitor c=0.014f //x=21.375 //y=5.21
c183 ( 18 0 ) capacitor c=0.00217843f //x=20.135 //y=1.655
c184 ( 17 0 ) capacitor c=0.0212471f //x=20.935 //y=1.655
c185 ( 9 0 ) capacitor c=0.0762833f //x=17.39 //y=2.08
c186 ( 7 0 ) capacitor c=0.00514991f //x=17.39 //y=4.54
c187 ( 2 0 ) capacitor c=0.00669602f //x=17.505 //y=3.7
c188 ( 1 0 ) capacitor c=0.100901f //x=21.345 //y=3.7
r189 (  69 70 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=17.425 //y=4.795 //x2=17.425 //y2=4.87
r190 (  67 69 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=17.425 //y=4.705 //x2=17.425 //y2=4.795
r191 (  63 64 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=17.39 //y=2.08 //x2=17.39 //y2=1.915
r192 (  61 74 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=17.955 //y=1.255 //x2=17.955 //y2=1.367
r193 (  60 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.955 //y=0.905 //x2=17.915 //y2=0.75
r194 (  60 61 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=17.955 //y=0.905 //x2=17.955 //y2=1.255
r195 (  55 72 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.58 //y=1.405 //x2=17.465 //y2=1.405
r196 (  54 74 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=17.8 //y=1.405 //x2=17.955 //y2=1.367
r197 (  53 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.58 //y=0.75 //x2=17.465 //y2=0.75
r198 (  52 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.8 //y=0.75 //x2=17.915 //y2=0.75
r199 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=17.8 //y=0.75 //x2=17.58 //y2=0.75
r200 (  51 69 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=17.56 //y=4.795 //x2=17.425 //y2=4.795
r201 (  50 57 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=17.795 //y=4.795 //x2=17.87 //y2=4.87
r202 (  50 51 ) resistor r=120.5 //w=0.094 //l=0.235 //layer=ply \
 //thickness=0.18 //x=17.795 //y=4.795 //x2=17.56 //y2=4.795
r203 (  45 72 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.425 //y=1.56 //x2=17.465 //y2=1.405
r204 (  45 64 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=17.425 //y=1.56 //x2=17.425 //y2=1.915
r205 (  44 72 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=17.425 //y=1.255 //x2=17.465 //y2=1.405
r206 (  43 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.425 //y=0.905 //x2=17.465 //y2=0.75
r207 (  43 44 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=17.425 //y=0.905 //x2=17.425 //y2=1.255
r208 (  42 57 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.87 //y=6.025 //x2=17.87 //y2=4.87
r209 (  41 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.43 //y=6.025 //x2=17.43 //y2=4.87
r210 (  40 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.69 //y=1.405 //x2=17.8 //y2=1.405
r211 (  40 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.69 //y=1.405 //x2=17.58 //y2=1.405
r212 (  38 67 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.425 //y=4.705 //x2=17.425 //y2=4.705
r213 (  34 36 ) resistor r=97.5401 //w=0.187 //l=1.425 //layer=li \
 //thickness=0.1 //x=21.46 //y=5.125 //x2=21.46 //y2=3.7
r214 (  33 36 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=21.46 //y=1.74 //x2=21.46 //y2=3.7
r215 (  32 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.105 //y=1.655 //x2=21.02 //y2=1.655
r216 (  31 33 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.375 //y=1.655 //x2=21.46 //y2=1.74
r217 (  31 32 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=21.375 //y=1.655 //x2=21.105 //y2=1.655
r218 (  29 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.375 //y=5.21 //x2=21.46 //y2=5.125
r219 (  29 30 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=21.375 //y=5.21 //x2=21.065 //y2=5.21
r220 (  25 39 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.02 //y=1.57 //x2=21.02 //y2=1.655
r221 (  25 76 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=21.02 //y=1.57 //x2=21.02 //y2=1
r222 (  19 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.98 //y=5.295 //x2=21.065 //y2=5.21
r223 (  19 79 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=20.98 //y=5.295 //x2=20.98 //y2=5.72
r224 (  17 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.935 //y=1.655 //x2=21.02 //y2=1.655
r225 (  17 18 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li \
 //thickness=0.1 //x=20.935 //y=1.655 //x2=20.135 //y2=1.655
r226 (  13 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.05 //y=1.57 //x2=20.135 //y2=1.655
r227 (  13 75 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=20.05 //y=1.57 //x2=20.05 //y2=1
r228 (  9 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.39 //y=2.08 //x2=17.39 //y2=2.08
r229 (  9 12 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=17.39 //y=2.08 //x2=17.39 //y2=3.7
r230 (  7 38 ) resistor r=11.332 //w=0.189 //l=0.173292 //layer=li \
 //thickness=0.1 //x=17.39 //y=4.54 //x2=17.407 //y2=4.705
r231 (  7 12 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=17.39 //y=4.54 //x2=17.39 //y2=3.7
r232 (  6 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.46 //y=3.7 //x2=21.46 //y2=3.7
r233 (  4 12 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.39 //y=3.7 //x2=17.39 //y2=3.7
r234 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.505 //y=3.7 //x2=17.39 //y2=3.7
r235 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=3.7 //x2=21.46 //y2=3.7
r236 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=3.7 //x2=17.505 //y2=3.7
ends PM_DLATCHN\%noxref_11

subckt PM_DLATCHN\%GATE_N ( 1 2 3 4 5 6 8 19 20 21 22 23 24 25 29 30 31 33 39 \
 40 42 )
c49 ( 42 0 ) capacitor c=0.0537799f //x=0.74 //y=2.085
c50 ( 40 0 ) capacitor c=0.0435629f //x=1.38 //y=1.255
c51 ( 39 0 ) capacitor c=0.0200386f //x=1.38 //y=0.91
c52 ( 33 0 ) capacitor c=0.0152946f //x=1.225 //y=1.41
c53 ( 31 0 ) capacitor c=0.0157804f //x=1.225 //y=0.755
c54 ( 30 0 ) capacitor c=0.0524167f //x=0.97 //y=4.79
c55 ( 29 0 ) capacitor c=0.0323991f //x=1.26 //y=4.79
c56 ( 25 0 ) capacitor c=0.0290017f //x=0.85 //y=1.92
c57 ( 24 0 ) capacitor c=0.0250027f //x=0.85 //y=1.565
c58 ( 23 0 ) capacitor c=0.0234316f //x=0.85 //y=1.255
c59 ( 22 0 ) capacitor c=0.0200596f //x=0.85 //y=0.91
c60 ( 21 0 ) capacitor c=0.154218f //x=1.335 //y=6.02
c61 ( 20 0 ) capacitor c=0.154243f //x=0.895 //y=6.02
c62 ( 8 0 ) capacitor c=0.114231f //x=0.74 //y=2.085
r63 (  42 43 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=0.74 //y=2.085 //x2=0.85 //y2=2.085
r64 (  40 49 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=1.255 //x2=1.34 //y2=1.41
r65 (  39 48 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.34 //y2=0.755
r66 (  39 40 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.38 //y2=1.255
r67 (  34 47 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=1.41 //x2=0.89 //y2=1.41
r68 (  33 49 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=1.41 //x2=1.34 //y2=1.41
r69 (  32 46 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=0.755 //x2=0.89 //y2=0.755
r70 (  31 48 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.34 //y2=0.755
r71 (  31 32 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.005 //y2=0.755
r72 (  29 36 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=1.335 //y2=4.865
r73 (  29 30 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=0.97 //y2=4.79
r74 (  26 30 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.97 //y2=4.79
r75 (  26 45 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.74 //y2=4.7
r76 (  25 43 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.92 //x2=0.85 //y2=2.085
r77 (  24 47 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.89 //y2=1.41
r78 (  24 25 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.85 //y2=1.92
r79 (  23 47 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.255 //x2=0.89 //y2=1.41
r80 (  22 46 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.89 //y2=0.755
r81 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.85 //y2=1.255
r82 (  21 36 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.335 //y=6.02 //x2=1.335 //y2=4.865
r83 (  20 26 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=0.895 //y=6.02 //x2=0.895 //y2=4.865
r84 (  19 33 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.225 //y2=1.41
r85 (  19 34 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.005 //y2=1.41
r86 (  17 45 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=4.7 //x2=0.74 //y2=4.7
r87 (  8 42 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=2.085 //x2=0.74 //y2=2.085
r88 (  6 17 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li //thickness=0.1 \
 //x=0.74 //y=4.44 //x2=0.74 //y2=4.7
r89 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=4.07 //x2=0.74 //y2=4.44
r90 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=3.7 //x2=0.74 //y2=4.07
r91 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=3.33 //x2=0.74 //y2=3.7
r92 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.96 //x2=0.74 //y2=3.33
r93 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.59 //x2=0.74 //y2=2.96
r94 (  1 8 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.59 //x2=0.74 //y2=2.085
ends PM_DLATCHN\%GATE_N

subckt PM_DLATCHN\%noxref_13 ( 1 5 9 10 13 17 29 )
c54 ( 29 0 ) capacitor c=0.0631306f //x=5 //y=0.365
c55 ( 17 0 ) capacitor c=0.00722223f //x=7.075 //y=0.615
c56 ( 13 0 ) capacitor c=0.0149611f //x=6.99 //y=0.53
c57 ( 10 0 ) capacitor c=0.00638024f //x=6.105 //y=1.495
c58 ( 9 0 ) capacitor c=0.006761f //x=6.105 //y=0.615
c59 ( 5 0 ) capacitor c=0.0189075f //x=6.02 //y=1.58
c60 ( 1 0 ) capacitor c=0.00798521f //x=5.135 //y=1.495
r61 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=7.075 //y=0.615 //x2=7.075 //y2=0.49
r62 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=7.075 //y=0.615 //x2=7.075 //y2=0.88
r63 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.19 //y=0.53 //x2=6.105 //y2=0.49
r64 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.19 //y=0.53 //x2=6.59 //y2=0.53
r65 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.99 //y=0.53 //x2=7.075 //y2=0.49
r66 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.99 //y=0.53 //x2=6.59 //y2=0.53
r67 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=6.105 //y=1.495 //x2=6.105 //y2=1.62
r68 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.105 //y=1.495 //x2=6.105 //y2=0.88
r69 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.105 //y=0.615 //x2=6.105 //y2=0.49
r70 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.105 //y=0.615 //x2=6.105 //y2=0.88
r71 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.22 //y=1.58 //x2=5.135 //y2=1.62
r72 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.22 //y=1.58 //x2=5.62 //y2=1.58
r73 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.02 //y=1.58 //x2=6.105 //y2=1.62
r74 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.02 //y=1.58 //x2=5.62 //y2=1.58
r75 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=5.135 //y=1.495 //x2=5.135 //y2=1.62
r76 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=5.135 //y=1.495 //x2=5.135 //y2=0.88
ends PM_DLATCHN\%noxref_13

subckt PM_DLATCHN\%noxref_14 ( 1 5 9 10 13 17 29 )
c54 ( 29 0 ) capacitor c=0.0633899f //x=10.55 //y=0.365
c55 ( 17 0 ) capacitor c=0.00722223f //x=12.625 //y=0.615
c56 ( 13 0 ) capacitor c=0.0149613f //x=12.54 //y=0.53
c57 ( 10 0 ) capacitor c=0.00687696f //x=11.655 //y=1.495
c58 ( 9 0 ) capacitor c=0.006761f //x=11.655 //y=0.615
c59 ( 5 0 ) capacitor c=0.0199444f //x=11.57 //y=1.58
c60 ( 1 0 ) capacitor c=0.00798521f //x=10.685 //y=1.495
r61 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=12.625 //y=0.615 //x2=12.625 //y2=0.49
r62 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=12.625 //y=0.615 //x2=12.625 //y2=0.88
r63 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.74 //y=0.53 //x2=11.655 //y2=0.49
r64 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.74 //y=0.53 //x2=12.14 //y2=0.53
r65 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.54 //y=0.53 //x2=12.625 //y2=0.49
r66 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.54 //y=0.53 //x2=12.14 //y2=0.53
r67 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=11.655 //y=1.495 //x2=11.655 //y2=1.62
r68 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=11.655 //y=1.495 //x2=11.655 //y2=0.88
r69 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=11.655 //y=0.615 //x2=11.655 //y2=0.49
r70 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=11.655 //y=0.615 //x2=11.655 //y2=0.88
r71 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.77 //y=1.58 //x2=10.685 //y2=1.62
r72 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.77 //y=1.58 //x2=11.17 //y2=1.58
r73 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.57 //y=1.58 //x2=11.655 //y2=1.62
r74 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.57 //y=1.58 //x2=11.17 //y2=1.58
r75 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=10.685 //y=1.495 //x2=10.685 //y2=1.62
r76 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=10.685 //y=1.495 //x2=10.685 //y2=0.88
ends PM_DLATCHN\%noxref_14

subckt PM_DLATCHN\%noxref_15 ( 7 8 15 16 23 24 25 )
c43 ( 25 0 ) capacitor c=0.0306628f //x=17.945 //y=5.025
c44 ( 24 0 ) capacitor c=0.0185379f //x=17.065 //y=5.025
c45 ( 23 0 ) capacitor c=0.0409962f //x=16.195 //y=5.025
c46 ( 16 0 ) capacitor c=0.00193672f //x=17.295 //y=6.91
c47 ( 15 0 ) capacitor c=0.0129692f //x=18.005 //y=6.91
c48 ( 8 0 ) capacitor c=0.00576007f //x=16.415 //y=5.21
c49 ( 7 0 ) capacitor c=0.0170172f //x=17.125 //y=5.21
r50 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.09 //y=6.825 //x2=18.09 //y2=6.74
r51 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.005 //y=6.91 //x2=18.09 //y2=6.825
r52 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=18.005 //y=6.91 //x2=17.295 //y2=6.91
r53 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.21 //y=6.825 //x2=17.295 //y2=6.91
r54 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=17.21 //y=6.825 //x2=17.21 //y2=6.4
r55 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=17.21 //y=5.295 //x2=17.21 //y2=5.72
r56 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.125 //y=5.21 //x2=17.21 //y2=5.295
r57 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=17.125 //y=5.21 //x2=16.415 //y2=5.21
r58 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.33 //y=5.295 //x2=16.415 //y2=5.21
r59 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=16.33 //y=5.295 //x2=16.33 //y2=5.72
ends PM_DLATCHN\%noxref_15

subckt PM_DLATCHN\%noxref_16 ( 7 8 15 16 23 24 25 )
c42 ( 25 0 ) capacitor c=0.0307189f //x=21.275 //y=5.025
c43 ( 24 0 ) capacitor c=0.0185379f //x=20.395 //y=5.025
c44 ( 23 0 ) capacitor c=0.0410313f //x=19.525 //y=5.025
c45 ( 16 0 ) capacitor c=0.00193672f //x=20.625 //y=6.91
c46 ( 15 0 ) capacitor c=0.0132919f //x=21.335 //y=6.91
c47 ( 8 0 ) capacitor c=0.0056411f //x=19.745 //y=5.21
c48 ( 7 0 ) capacitor c=0.0169676f //x=20.455 //y=5.21
r49 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.42 //y=6.825 //x2=21.42 //y2=6.74
r50 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.335 //y=6.91 //x2=21.42 //y2=6.825
r51 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=21.335 //y=6.91 //x2=20.625 //y2=6.91
r52 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.54 //y=6.825 //x2=20.625 //y2=6.91
r53 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=20.54 //y=6.825 //x2=20.54 //y2=6.4
r54 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=20.54 //y=5.295 //x2=20.54 //y2=5.72
r55 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.455 //y=5.21 //x2=20.54 //y2=5.295
r56 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=20.455 //y=5.21 //x2=19.745 //y2=5.21
r57 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=19.66 //y=5.295 //x2=19.745 //y2=5.21
r58 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=19.66 //y=5.295 //x2=19.66 //y2=5.72
ends PM_DLATCHN\%noxref_16

