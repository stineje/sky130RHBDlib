magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 2522 582
<< pwell >>
rect 99 201 2483 203
rect 1 23 2483 201
rect 1 21 344 23
rect 610 21 1116 23
rect 2011 21 2483 23
rect 29 -17 63 21
<< locali >>
rect 190 215 268 255
rect 1340 335 1374 357
rect 1320 185 1374 335
rect 1320 151 1385 185
rect 1351 119 1385 151
rect 2400 357 2467 493
rect 2104 215 2193 255
rect 2425 165 2467 357
rect 2399 51 2467 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 17 402 86 493
rect 120 436 154 527
rect 343 477 703 493
rect 188 459 703 477
rect 188 443 394 459
rect 188 402 222 443
rect 649 422 692 459
rect 17 368 222 402
rect 256 391 290 409
rect 17 300 88 368
rect 256 357 410 391
rect 513 357 579 409
rect 256 334 290 357
rect 122 300 290 334
rect 17 161 51 300
rect 122 265 156 300
rect 444 270 478 357
rect 85 199 156 265
rect 122 181 156 199
rect 302 187 348 265
rect 17 147 86 161
rect 122 147 265 181
rect 20 51 86 147
rect 126 17 160 109
rect 199 93 265 147
rect 302 153 305 187
rect 339 153 348 187
rect 302 133 348 153
rect 397 135 478 270
rect 590 253 624 323
rect 560 249 624 253
rect 528 219 624 249
rect 528 215 594 219
rect 658 185 692 422
rect 742 458 1013 492
rect 742 264 776 458
rect 816 339 889 424
rect 963 413 1013 458
rect 1052 447 1118 527
rect 1165 459 1590 493
rect 1165 413 1199 459
rect 963 379 1199 413
rect 1240 391 1442 425
rect 1240 379 1306 391
rect 1240 345 1274 379
rect 938 277 1034 345
rect 1127 311 1274 345
rect 966 265 1034 277
rect 742 230 814 264
rect 611 181 746 185
rect 444 119 478 135
rect 524 151 746 181
rect 524 147 627 151
rect 524 131 605 147
rect 643 93 678 117
rect 199 85 420 93
rect 503 85 678 93
rect 199 51 678 85
rect 712 85 746 151
rect 780 119 814 230
rect 848 187 898 265
rect 848 153 857 187
rect 891 153 898 187
rect 848 129 898 153
rect 966 199 1126 265
rect 966 102 1000 199
rect 1160 163 1194 311
rect 848 85 914 95
rect 712 51 914 85
rect 1036 17 1102 161
rect 1136 76 1194 163
rect 1228 148 1285 265
rect 1408 246 1442 391
rect 1476 306 1510 425
rect 1556 344 1590 459
rect 1644 459 1882 493
rect 1644 391 1678 459
rect 1712 357 1778 425
rect 1556 310 1607 344
rect 1476 272 1522 306
rect 1488 258 1522 272
rect 1408 212 1454 246
rect 1488 221 1539 258
rect 1420 185 1454 212
rect 1420 119 1470 185
rect 1251 85 1317 114
rect 1504 85 1539 221
rect 1573 199 1607 310
rect 1675 306 1778 357
rect 1848 409 1882 459
rect 2038 439 2072 527
rect 1848 408 2021 409
rect 1848 407 2024 408
rect 1848 406 2026 407
rect 1848 405 2029 406
rect 2107 405 2177 493
rect 1848 375 2177 405
rect 1675 289 1734 306
rect 1675 185 1711 289
rect 1767 199 1814 265
rect 1251 51 1539 85
rect 1573 85 1607 148
rect 1661 119 1711 185
rect 1848 153 1882 375
rect 2011 374 2177 375
rect 2014 373 2177 374
rect 2017 372 2177 373
rect 2020 371 2177 372
rect 1745 119 1882 153
rect 1928 307 2002 341
rect 1928 165 1962 307
rect 2036 289 2177 371
rect 2215 291 2281 493
rect 2315 357 2366 527
rect 2036 265 2070 289
rect 1996 199 2070 265
rect 2036 181 2070 199
rect 1928 85 1996 165
rect 2036 147 2182 181
rect 1573 51 1996 85
rect 2036 17 2070 113
rect 2106 57 2182 147
rect 2231 136 2281 291
rect 2329 199 2391 323
rect 2231 54 2265 136
rect 2299 17 2365 102
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 305 153 339 187
rect 857 153 891 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
<< metal1 >>
rect 0 561 2484 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2484 561
rect 0 496 2484 527
rect 293 187 351 193
rect 293 153 305 187
rect 339 184 351 187
rect 845 187 903 193
rect 845 184 857 187
rect 339 156 857 184
rect 339 153 351 156
rect 293 147 351 153
rect 845 153 857 156
rect 891 153 903 187
rect 845 147 903 153
rect 0 17 2484 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2484 17
rect 0 -48 2484 -17
<< obsm1 >>
rect 364 388 422 397
rect 502 388 560 397
rect 816 388 874 397
rect 364 360 874 388
rect 364 351 422 360
rect 502 351 560 360
rect 816 351 874 360
rect 578 320 636 329
rect 940 320 998 329
rect 578 292 998 320
rect 578 283 636 292
rect 940 283 998 292
rect 1676 320 1734 329
rect 2324 320 2382 329
rect 1676 292 2382 320
rect 1676 283 1734 292
rect 2324 283 2382 292
rect 385 252 443 261
rect 1216 252 1274 261
rect 1768 252 1826 261
rect 385 224 1826 252
rect 385 215 443 224
rect 1216 215 1274 224
rect 1768 215 1826 224
rect 1492 184 1550 193
rect 2232 184 2290 193
rect 1492 156 2290 184
rect 1492 147 1550 156
rect 2232 147 2290 156
<< labels >>
rlabel locali s 190 215 268 255 6 A
port 1 nsew signal input
rlabel metal1 s 845 147 903 156 6 B
port 2 nsew signal input
rlabel metal1 s 293 147 351 156 6 B
port 2 nsew signal input
rlabel metal1 s 293 156 903 184 6 B
port 2 nsew signal input
rlabel metal1 s 845 184 903 193 6 B
port 2 nsew signal input
rlabel metal1 s 293 184 351 193 6 B
port 2 nsew signal input
rlabel locali s 2104 215 2193 255 6 CIN
port 3 nsew signal input
rlabel metal1 s 0 -48 2484 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 2011 21 2483 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 610 21 1116 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 344 23 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 23 2483 201 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 99 201 2483 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 2522 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2484 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1351 119 1385 151 6 COUT
port 8 nsew signal output
rlabel locali s 1320 151 1385 185 6 COUT
port 8 nsew signal output
rlabel locali s 1320 185 1374 335 6 COUT
port 8 nsew signal output
rlabel locali s 1340 335 1374 357 6 COUT
port 8 nsew signal output
rlabel locali s 2399 51 2467 165 6 SUM
port 9 nsew signal output
rlabel locali s 2425 165 2467 357 6 SUM
port 9 nsew signal output
rlabel locali s 2400 357 2467 493 6 SUM
port 9 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2484 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 2132810
string GDS_START 2113526
<< end >>
