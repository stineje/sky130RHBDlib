magic
tech sky130A
magscale 1 2
timestamp 1652332156
<< nwell >>
rect 531 1532 1689 1550
rect 528 1514 1026 1532
rect 1194 1514 1692 1532
rect 478 1446 1076 1514
rect 1144 1446 1742 1514
rect 528 1439 1026 1446
rect 528 968 539 1439
rect 585 1330 619 1364
rect 1015 968 1026 1439
rect 528 825 1026 968
rect 1194 1440 1692 1446
rect 1194 968 1205 1440
rect 1681 968 1692 1440
rect 1194 825 1692 968
rect 531 786 1689 825
<< pwell >>
rect -34 -34 2254 544
<< pdiffc >>
rect 585 1330 619 1364
rect 761 1330 795 1364
rect 937 1330 971 1364
rect 1251 1330 1285 1364
rect 1427 1330 1461 1364
rect 1603 1330 1637 1364
rect 585 1058 619 1092
rect 761 1058 795 1092
rect 849 1058 883 1092
rect 1251 1058 1285 1092
rect 1427 1058 1461 1092
rect 1515 1058 1549 1092
<< psubdiff >>
rect 478 482 1079 544
rect 1141 482 1742 544
rect 478 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1076 17
rect 478 -34 1076 -17
rect 1144 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1742 17
rect 1144 -34 1742 -17
<< nsubdiff >>
rect 478 1497 1076 1514
rect 478 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1076 1497
rect 1144 1497 1742 1514
rect 1144 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1742 1497
rect 478 822 1079 884
rect 1141 822 1742 884
<< psubdiffcont >>
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
<< nsubdiffcont >>
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
<< poly >>
rect 612 383 639 413
rect 806 383 861 413
rect 1278 383 1305 413
rect 1472 383 1527 413
rect 612 375 642 383
rect 806 382 836 383
rect 1278 375 1308 383
rect 1472 382 1502 383
<< locali >>
rect 478 1497 1076 1514
rect 478 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1076 1497
rect 478 1446 1076 1463
rect 1144 1497 1742 1514
rect 1144 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1742 1497
rect 1144 1446 1742 1463
rect 585 1364 619 1380
rect 585 1312 619 1330
rect 673 1312 707 1446
rect 761 1364 971 1398
rect 761 1312 795 1330
rect 937 1312 971 1330
rect 1251 1364 1285 1380
rect 1251 1312 1285 1330
rect 1339 1312 1373 1446
rect 1427 1364 1637 1398
rect 1427 1312 1461 1330
rect 1603 1312 1637 1330
rect 585 1092 619 1110
rect 761 1092 795 1110
rect 585 1024 795 1058
rect 849 1092 883 1110
rect 1251 1092 1285 1110
rect 1427 1092 1461 1110
rect 849 1024 979 1058
rect 1251 1024 1461 1058
rect 1515 1092 1549 1110
rect 1515 1024 1645 1058
rect 649 447 683 907
rect 871 825 905 907
rect 871 449 905 617
rect 945 347 979 1024
rect 1315 862 1349 907
rect 1315 444 1349 634
rect 1537 448 1571 907
rect 1611 347 1645 1024
rect 857 313 979 347
rect 1523 313 1645 347
rect 857 216 891 313
rect 1523 216 1557 313
rect 663 34 697 174
rect 1329 34 1363 174
rect 478 17 1076 34
rect 478 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1076 17
rect 478 -34 1076 -17
rect 1144 17 1742 34
rect 1144 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1742 17
rect 1144 -34 1742 -17
<< viali >>
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
<< metal1 >>
rect 478 1497 1076 1514
rect 478 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1076 1497
rect 478 1446 1076 1463
rect 1144 1497 1742 1514
rect 1144 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1742 1497
rect 1144 1446 1742 1463
rect 1378 871 1905 905
rect 187 797 623 831
rect 939 797 2022 831
rect 981 723 1586 757
rect 1372 649 2053 683
rect 905 575 1882 609
rect 315 501 1512 535
rect 478 17 1076 34
rect 478 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1076 17
rect 478 -34 1076 -17
rect 1144 17 1742 34
rect 1144 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1742 17
rect 1144 -34 1742 -17
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 148 0 -1 814
box -53 -33 29 33
use invx1_pcell  invx1_pcell_0
timestamp 1652329846
transform 1 0 0 0 1 0
box -87 -34 531 1550
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform -1 0 296 0 -1 518
box -53 -33 29 33
use diff_ring_side  diff_ring_side_1
timestamp 1652319726
transform 1 0 444 0 1 0
box -87 -34 87 1550
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 666 0 1 814
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_0
timestamp 1648060378
transform 0 1 667 -1 0 941
box -32 -28 34 26
use pmos2_1  pmos2_1_0
timestamp 1647326732
transform 1 0 487 0 1 1403
box 52 -460 352 37
use pmos2_1  pmos2_1_1
timestamp 1647326732
transform 1 0 663 0 1 1403
box 52 -460 352 37
use poly_li1_contact  poly_li1_contact_1
timestamp 1648060378
transform 0 1 667 -1 0 417
box -32 -28 34 26
use nmos_top_trim1  nmos_top_trim1_0
timestamp 1651256895
transform -1 0 998 0 1 73
box 0 0 248 309
use nmos_bottom  nmos_bottom_0
timestamp 1651256857
transform -1 0 804 0 1 73
box 0 0 248 302
use diff_ring_side  diff_ring_side_0
timestamp 1652319726
transform 1 0 1110 0 1 0
box -87 -34 87 1550
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 888 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform -1 0 962 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform -1 0 888 0 -1 592
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_3
timestamp 1648060378
transform 0 1 889 -1 0 941
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_2
timestamp 1648060378
transform 0 1 889 -1 0 417
box -32 -28 34 26
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform -1 0 1332 0 -1 666
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_5
timestamp 1648060378
transform 0 1 1333 -1 0 941
box -32 -28 34 26
use pmos2_1  pmos2_1_3
timestamp 1647326732
transform 1 0 1329 0 1 1403
box 52 -460 352 37
use pmos2_1  pmos2_1_2
timestamp 1647326732
transform 1 0 1153 0 1 1403
box 52 -460 352 37
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform -1 0 1332 0 -1 888
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_4
timestamp 1648060378
transform 0 1 1333 -1 0 417
box -32 -28 34 26
use nmos_top_trim1  nmos_top_trim1_1
timestamp 1651256895
transform -1 0 1664 0 1 73
box 0 0 248 309
use nmos_bottom  nmos_bottom_1
timestamp 1651256857
transform -1 0 1470 0 1 73
box 0 0 248 302
use diff_ring_side  diff_ring_side_3
timestamp 1652319726
transform 1 0 1776 0 1 0
box -87 -34 87 1550
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 1628 0 1 740
box -53 -33 29 33
use poly_li1_contact  poly_li1_contact_7
timestamp 1648060378
transform 0 1 1555 -1 0 941
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_6
timestamp 1648060378
transform 0 1 1555 -1 0 417
box -32 -28 34 26
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform 1 0 1554 0 1 518
box -53 -33 29 33
use invx1_pcell  invx1_pcell_1
timestamp 1652329846
transform -1 0 2220 0 1 0
box -87 -34 531 1550
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform 1 0 1924 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform 1 0 2072 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform 1 0 2072 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 1924 0 1 592
box -53 -33 29 33
<< end >>
