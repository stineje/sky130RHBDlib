magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1931 203
rect 29 -17 63 21
<< scnmos >>
rect 86 47 116 177
rect 170 47 200 177
rect 271 47 301 177
rect 507 47 537 177
rect 591 47 621 177
rect 675 47 705 177
rect 759 47 789 177
rect 843 47 873 177
rect 927 47 957 177
rect 1011 47 1041 177
rect 1095 47 1125 177
rect 1231 47 1261 177
rect 1315 47 1345 177
rect 1399 47 1429 177
rect 1483 47 1513 177
rect 1567 47 1597 177
rect 1651 47 1681 177
rect 1735 47 1765 177
rect 1819 47 1849 177
<< scpmoshvt >>
rect 86 297 116 497
rect 170 297 200 497
rect 271 297 301 497
rect 459 309 489 497
rect 543 309 573 497
rect 627 309 657 497
rect 711 309 741 497
rect 795 309 825 497
rect 879 309 909 497
rect 963 309 993 497
rect 1047 309 1077 497
rect 1231 297 1261 497
rect 1315 297 1345 497
rect 1399 297 1429 497
rect 1483 297 1513 497
rect 1567 297 1597 497
rect 1651 297 1681 497
rect 1735 297 1765 497
rect 1819 297 1849 497
<< ndiff >>
rect 27 157 86 177
rect 27 123 39 157
rect 73 123 86 157
rect 27 89 86 123
rect 27 55 39 89
rect 73 55 86 89
rect 27 47 86 55
rect 116 106 170 177
rect 116 72 126 106
rect 160 72 170 106
rect 116 47 170 72
rect 200 89 271 177
rect 200 55 210 89
rect 244 55 271 89
rect 200 47 271 55
rect 301 129 353 177
rect 301 95 311 129
rect 345 95 353 129
rect 301 47 353 95
rect 455 129 507 177
rect 455 95 463 129
rect 497 95 507 129
rect 455 47 507 95
rect 537 89 591 177
rect 537 55 547 89
rect 581 55 591 89
rect 537 47 591 55
rect 621 129 675 177
rect 621 95 631 129
rect 665 95 675 129
rect 621 47 675 95
rect 705 89 759 177
rect 705 55 715 89
rect 749 55 759 89
rect 705 47 759 55
rect 789 129 843 177
rect 789 95 799 129
rect 833 95 843 129
rect 789 47 843 95
rect 873 89 927 177
rect 873 55 883 89
rect 917 55 927 89
rect 873 47 927 55
rect 957 129 1011 177
rect 957 95 967 129
rect 1001 95 1011 129
rect 957 47 1011 95
rect 1041 89 1095 177
rect 1041 55 1051 89
rect 1085 55 1095 89
rect 1041 47 1095 55
rect 1125 129 1231 177
rect 1125 95 1162 129
rect 1196 95 1231 129
rect 1125 47 1231 95
rect 1261 169 1315 177
rect 1261 135 1271 169
rect 1305 135 1315 169
rect 1261 47 1315 135
rect 1345 89 1399 177
rect 1345 55 1355 89
rect 1389 55 1399 89
rect 1345 47 1399 55
rect 1429 169 1483 177
rect 1429 135 1439 169
rect 1473 135 1483 169
rect 1429 47 1483 135
rect 1513 89 1567 177
rect 1513 55 1523 89
rect 1557 55 1567 89
rect 1513 47 1567 55
rect 1597 169 1651 177
rect 1597 135 1607 169
rect 1641 135 1651 169
rect 1597 47 1651 135
rect 1681 89 1735 177
rect 1681 55 1691 89
rect 1725 55 1735 89
rect 1681 47 1735 55
rect 1765 169 1819 177
rect 1765 135 1775 169
rect 1809 135 1819 169
rect 1765 47 1819 135
rect 1849 89 1905 177
rect 1849 55 1859 89
rect 1893 55 1905 89
rect 1849 47 1905 55
<< pdiff >>
rect 27 489 86 497
rect 27 455 39 489
rect 73 455 86 489
rect 27 421 86 455
rect 27 387 39 421
rect 73 387 86 421
rect 27 297 86 387
rect 116 461 170 497
rect 116 427 126 461
rect 160 427 170 461
rect 116 297 170 427
rect 200 489 271 497
rect 200 455 210 489
rect 244 455 271 489
rect 200 421 271 455
rect 200 387 210 421
rect 244 387 271 421
rect 200 297 271 387
rect 301 479 353 497
rect 301 445 311 479
rect 345 445 353 479
rect 301 411 353 445
rect 301 377 311 411
rect 345 377 353 411
rect 301 343 353 377
rect 301 309 311 343
rect 345 309 353 343
rect 407 477 459 497
rect 407 443 415 477
rect 449 443 459 477
rect 407 309 459 443
rect 489 489 543 497
rect 489 455 499 489
rect 533 455 543 489
rect 489 309 543 455
rect 573 477 627 497
rect 573 443 583 477
rect 617 443 627 477
rect 573 309 627 443
rect 657 489 711 497
rect 657 455 667 489
rect 701 455 711 489
rect 657 309 711 455
rect 741 477 795 497
rect 741 443 751 477
rect 785 443 795 477
rect 741 309 795 443
rect 825 489 879 497
rect 825 455 835 489
rect 869 455 879 489
rect 825 309 879 455
rect 909 477 963 497
rect 909 443 919 477
rect 953 443 963 477
rect 909 309 963 443
rect 993 489 1047 497
rect 993 455 1003 489
rect 1037 455 1047 489
rect 993 309 1047 455
rect 1077 477 1231 497
rect 1077 443 1104 477
rect 1138 443 1172 477
rect 1206 443 1231 477
rect 1077 309 1231 443
rect 301 297 353 309
rect 1092 297 1231 309
rect 1261 345 1315 497
rect 1261 311 1271 345
rect 1305 311 1315 345
rect 1261 297 1315 311
rect 1345 489 1399 497
rect 1345 455 1355 489
rect 1389 455 1399 489
rect 1345 421 1399 455
rect 1345 387 1355 421
rect 1389 387 1399 421
rect 1345 297 1399 387
rect 1429 345 1483 497
rect 1429 311 1439 345
rect 1473 311 1483 345
rect 1429 297 1483 311
rect 1513 489 1567 497
rect 1513 455 1523 489
rect 1557 455 1567 489
rect 1513 421 1567 455
rect 1513 387 1523 421
rect 1557 387 1567 421
rect 1513 297 1567 387
rect 1597 345 1651 497
rect 1597 311 1607 345
rect 1641 311 1651 345
rect 1597 297 1651 311
rect 1681 489 1735 497
rect 1681 455 1691 489
rect 1725 455 1735 489
rect 1681 421 1735 455
rect 1681 387 1691 421
rect 1725 387 1735 421
rect 1681 297 1735 387
rect 1765 345 1819 497
rect 1765 311 1775 345
rect 1809 311 1819 345
rect 1765 297 1819 311
rect 1849 489 1905 497
rect 1849 455 1859 489
rect 1893 455 1905 489
rect 1849 421 1905 455
rect 1849 387 1859 421
rect 1893 387 1905 421
rect 1849 297 1905 387
<< ndiffc >>
rect 39 123 73 157
rect 39 55 73 89
rect 126 72 160 106
rect 210 55 244 89
rect 311 95 345 129
rect 463 95 497 129
rect 547 55 581 89
rect 631 95 665 129
rect 715 55 749 89
rect 799 95 833 129
rect 883 55 917 89
rect 967 95 1001 129
rect 1051 55 1085 89
rect 1162 95 1196 129
rect 1271 135 1305 169
rect 1355 55 1389 89
rect 1439 135 1473 169
rect 1523 55 1557 89
rect 1607 135 1641 169
rect 1691 55 1725 89
rect 1775 135 1809 169
rect 1859 55 1893 89
<< pdiffc >>
rect 39 455 73 489
rect 39 387 73 421
rect 126 427 160 461
rect 210 455 244 489
rect 210 387 244 421
rect 311 445 345 479
rect 311 377 345 411
rect 311 309 345 343
rect 415 443 449 477
rect 499 455 533 489
rect 583 443 617 477
rect 667 455 701 489
rect 751 443 785 477
rect 835 455 869 489
rect 919 443 953 477
rect 1003 455 1037 489
rect 1104 443 1138 477
rect 1172 443 1206 477
rect 1271 311 1305 345
rect 1355 455 1389 489
rect 1355 387 1389 421
rect 1439 311 1473 345
rect 1523 455 1557 489
rect 1523 387 1557 421
rect 1607 311 1641 345
rect 1691 455 1725 489
rect 1691 387 1725 421
rect 1775 311 1809 345
rect 1859 455 1893 489
rect 1859 387 1893 421
<< poly >>
rect 86 497 116 523
rect 170 497 200 523
rect 271 497 301 523
rect 459 497 489 523
rect 543 497 573 523
rect 627 497 657 523
rect 711 497 741 523
rect 795 497 825 523
rect 879 497 909 523
rect 963 497 993 523
rect 1047 497 1077 523
rect 1231 497 1261 523
rect 1315 497 1345 523
rect 1399 497 1429 523
rect 1483 497 1513 523
rect 1567 497 1597 523
rect 1651 497 1681 523
rect 1735 497 1765 523
rect 1819 497 1849 523
rect 86 265 116 297
rect 32 259 116 265
rect 170 259 200 297
rect 271 265 301 297
rect 459 294 489 309
rect 543 294 573 309
rect 627 294 657 309
rect 711 294 741 309
rect 795 294 825 309
rect 879 294 909 309
rect 963 294 993 309
rect 1047 294 1077 309
rect 384 265 1077 294
rect 32 249 200 259
rect 32 215 42 249
rect 76 215 200 249
rect 32 205 200 215
rect 32 199 116 205
rect 86 177 116 199
rect 170 177 200 205
rect 242 264 1077 265
rect 242 249 414 264
rect 1231 259 1261 297
rect 1315 259 1345 297
rect 1399 259 1429 297
rect 1483 259 1513 297
rect 1567 259 1597 297
rect 1651 259 1681 297
rect 1735 259 1765 297
rect 1819 259 1849 297
rect 242 215 252 249
rect 286 215 414 249
rect 1119 249 1185 259
rect 1119 222 1135 249
rect 242 199 414 215
rect 507 215 1135 222
rect 1169 215 1185 249
rect 271 177 301 199
rect 507 192 1185 215
rect 1231 249 1849 259
rect 1231 215 1255 249
rect 1289 215 1323 249
rect 1357 215 1391 249
rect 1425 215 1459 249
rect 1493 215 1527 249
rect 1561 215 1595 249
rect 1629 215 1663 249
rect 1697 215 1731 249
rect 1765 215 1849 249
rect 1231 205 1849 215
rect 507 177 537 192
rect 591 177 621 192
rect 675 177 705 192
rect 759 177 789 192
rect 843 177 873 192
rect 927 177 957 192
rect 1011 177 1041 192
rect 1095 177 1125 192
rect 1231 177 1261 205
rect 1315 177 1345 205
rect 1399 177 1429 205
rect 1483 177 1513 205
rect 1567 177 1597 205
rect 1651 177 1681 205
rect 1735 177 1765 205
rect 1819 177 1849 205
rect 86 21 116 47
rect 170 21 200 47
rect 271 21 301 47
rect 507 21 537 47
rect 591 21 621 47
rect 675 21 705 47
rect 759 21 789 47
rect 843 21 873 47
rect 927 21 957 47
rect 1011 21 1041 47
rect 1095 21 1125 47
rect 1231 21 1261 47
rect 1315 21 1345 47
rect 1399 21 1429 47
rect 1483 21 1513 47
rect 1567 21 1597 47
rect 1651 21 1681 47
rect 1735 21 1765 47
rect 1819 21 1849 47
<< polycont >>
rect 42 215 76 249
rect 252 215 286 249
rect 1135 215 1169 249
rect 1255 215 1289 249
rect 1323 215 1357 249
rect 1391 215 1425 249
rect 1459 215 1493 249
rect 1527 215 1561 249
rect 1595 215 1629 249
rect 1663 215 1697 249
rect 1731 215 1765 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 17 489 89 527
rect 17 455 39 489
rect 73 455 89 489
rect 17 421 89 455
rect 17 387 39 421
rect 73 387 89 421
rect 17 357 89 387
rect 123 461 160 493
rect 123 427 126 461
rect 123 323 160 427
rect 194 489 261 527
rect 194 455 210 489
rect 244 455 261 489
rect 194 421 261 455
rect 194 387 210 421
rect 244 387 261 421
rect 194 373 261 387
rect 295 479 365 493
rect 295 445 311 479
rect 345 445 365 479
rect 295 411 365 445
rect 295 377 311 411
rect 345 377 365 411
rect 399 477 449 493
rect 399 443 415 477
rect 483 489 549 527
rect 483 455 499 489
rect 533 455 549 489
rect 483 447 549 455
rect 583 477 617 493
rect 399 413 449 443
rect 651 489 717 527
rect 651 455 667 489
rect 701 455 717 489
rect 651 447 717 455
rect 751 477 785 493
rect 583 413 617 443
rect 819 489 885 527
rect 819 455 835 489
rect 869 455 885 489
rect 819 447 885 455
rect 919 477 953 493
rect 751 413 785 443
rect 987 489 1053 527
rect 987 455 1003 489
rect 1037 455 1053 489
rect 987 447 1053 455
rect 1087 489 1915 493
rect 1087 477 1355 489
rect 919 413 953 443
rect 1087 443 1104 477
rect 1138 443 1172 477
rect 1206 455 1355 477
rect 1389 455 1523 489
rect 1557 455 1691 489
rect 1725 455 1859 489
rect 1893 455 1915 489
rect 1206 443 1915 455
rect 1087 421 1915 443
rect 1087 413 1355 421
rect 399 387 1355 413
rect 1389 387 1523 421
rect 1557 387 1691 421
rect 1725 387 1859 421
rect 1893 387 1915 421
rect 399 379 1915 387
rect 295 343 365 377
rect 17 249 86 323
rect 17 215 42 249
rect 76 215 86 249
rect 17 199 86 215
rect 120 255 160 323
rect 120 221 121 255
rect 155 221 160 255
rect 120 199 160 221
rect 17 157 89 165
rect 17 123 39 157
rect 73 123 89 157
rect 17 89 89 123
rect 17 55 39 89
rect 73 55 89 89
rect 123 106 160 199
rect 194 265 261 339
rect 295 309 311 343
rect 345 309 365 343
rect 295 299 365 309
rect 194 249 286 265
rect 194 215 252 249
rect 194 199 286 215
rect 320 255 365 299
rect 399 311 1271 345
rect 1305 311 1439 345
rect 1473 311 1607 345
rect 1641 311 1775 345
rect 1809 311 1915 345
rect 399 289 1915 311
rect 320 249 1185 255
rect 320 215 1135 249
rect 1169 215 1185 249
rect 320 205 1185 215
rect 1235 249 1316 255
rect 1350 249 1831 255
rect 1235 215 1255 249
rect 1289 221 1316 249
rect 1289 215 1323 221
rect 1357 215 1391 249
rect 1425 215 1459 249
rect 1493 215 1527 249
rect 1561 215 1595 249
rect 1629 215 1663 249
rect 1697 215 1731 249
rect 1765 215 1831 249
rect 1235 205 1831 215
rect 194 124 261 199
rect 320 165 397 205
rect 1865 171 1915 289
rect 295 129 397 165
rect 123 72 126 106
rect 295 95 311 129
rect 345 95 397 129
rect 123 56 160 72
rect 17 17 89 55
rect 194 55 210 89
rect 244 55 261 89
rect 194 17 261 55
rect 295 51 397 95
rect 431 131 1221 171
rect 431 129 497 131
rect 431 95 463 129
rect 631 129 665 131
rect 431 51 497 95
rect 531 89 597 97
rect 531 55 547 89
rect 581 55 597 89
rect 799 129 833 131
rect 631 55 665 95
rect 699 89 765 97
rect 699 55 715 89
rect 749 55 765 89
rect 531 17 597 55
rect 699 17 765 55
rect 967 129 1001 131
rect 799 51 833 95
rect 867 89 933 97
rect 867 55 883 89
rect 917 55 933 89
rect 1135 129 1221 131
rect 967 55 1001 95
rect 1035 89 1101 97
rect 1035 55 1051 89
rect 1085 55 1101 89
rect 867 17 933 55
rect 1035 17 1101 55
rect 1135 95 1162 129
rect 1196 95 1221 129
rect 1255 169 1915 171
rect 1255 135 1271 169
rect 1305 135 1439 169
rect 1473 135 1607 169
rect 1641 135 1775 169
rect 1809 135 1915 169
rect 1255 123 1915 135
rect 1135 89 1221 95
rect 1135 55 1355 89
rect 1389 55 1523 89
rect 1557 55 1691 89
rect 1725 55 1859 89
rect 1893 55 1915 89
rect 1135 51 1915 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 121 221 155 255
rect 1316 249 1350 255
rect 1316 221 1323 249
rect 1323 221 1350 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 109 255 167 261
rect 109 221 121 255
rect 155 252 167 255
rect 1304 255 1362 261
rect 1304 252 1316 255
rect 155 224 1316 252
rect 155 221 167 224
rect 109 215 167 221
rect 1304 221 1316 224
rect 1350 221 1362 255
rect 1304 215 1362 221
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 1868 153 1902 187 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1868 221 1902 255 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 857 289 891 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 949 289 983 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1041 289 1075 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1133 289 1167 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 489 289 523 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 581 289 615 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 673 289 707 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 765 289 799 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 213 153 247 187 0 FreeSans 200 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 1224 289 1258 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1408 289 1442 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 213 289 247 323 0 FreeSans 200 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 1868 289 1902 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1776 289 1810 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1500 289 1534 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1592 289 1626 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 1684 289 1718 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 ebufn_8
rlabel metal1 s 0 -48 1932 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1932 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 2970756
string GDS_START 2956844
<< end >>
