* SPICE3 file created from TMRDFFQNX1.ext - technology: sky130A

.subckt TMRDFFQNX1 QN D CLK VDD GND
M1000 GND a_7469_1050.t5 a_8030_101.t0 nshort w=-1.605u l=1.765u
+  ad=3.7611p pd=32.97u as=0p ps=0u
M1001 a_599_989.t4 D.t0 VDD.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t81 a_10429_1050.t5 a_8731_187.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 QN.t4 a_7595_411.t5 a_13757_1051.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_10429_1050.t4 a_8731_187.t5 VDD.t70 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_7469_1050.t3 a_7595_411.t7 VDD.t74 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VDD.t26 a_9183_989.t5 a_8861_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 GND a_1845_1050.t5 a_2406_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_4569_1050.t1 CLK.t0 VDD.t80 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VDD.t64 a_4439_187.t5 a_6137_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1845_1050.t1 a_599_989.t5 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VDD.t73 a_8861_1050.t7 a_9183_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_8861_1050.t2 CLK.t1 VDD.t39 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 GND a_8861_1050.t8 a_9658_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_13093_1051.t3 a_11887_411.t5 VDD.t40 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VDD.t14 a_147_187.t6 a_1845_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_6137_1050.t0 a_4891_989.t5 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VDD.t62 a_4569_1050.t7 a_4891_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_13093_1051.t1 a_11887_411.t6 a_13757_1051.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VDD.t32 a_4439_187.t6 a_7595_411.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 VDD.t42 a_147_187.t7 a_277_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VDD.t27 a_6137_1050.t5 a_4439_187.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VDD.t69 a_8731_187.t8 a_8861_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 GND a_147_187.t8 a_91_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_3177_1050.t4 a_277_1050.t7 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 VDD.t2 a_1845_1050.t6 a_147_187.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_11887_411.t4 a_11761_1050.t5 VDD.t35 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VDD.t7 D.t2 a_9183_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 QN a_7595_411.t9 a_14320_101.t0 nshort w=-1.83u l=2.06u
+  ad=0.5373p pd=4.72u as=0p ps=0u
M1029 GND a_8861_1050.t9 a_11656_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1030 VDD.t12 D.t3 a_4891_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 GND a_10429_1050.t6 a_10990_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1032 GND a_4439_187.t8 a_4383_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1033 VDD.t43 a_7469_1050.t6 a_7595_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 VDD.t61 CLK.t2 a_277_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_13757_1051.t5 a_7595_411.t8 QN.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_3177_1050.t1 a_3303_411.t7 VDD.t44 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VDD.t21 CLK.t5 a_147_187.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_11887_411.t2 a_8731_187.t10 VDD.t68 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 GND a_599_989.t8 a_1740_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1040 VDD.t16 a_11887_411.t7 a_11761_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 GND a_4569_1050.t9 a_5366_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1042 VDD.t38 CLK.t6 a_4439_187.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1043 GND a_11887_411.t8 a_13654_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_9183_989.t1 D.t4 VDD.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_3303_411.t2 a_3177_1050.t5 VDD.t37 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 GND a_11887_411.t10 a_12988_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1047 VDD.t33 a_599_989.t7 a_277_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 VDD.t1 a_277_1050.t8 a_599_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_8731_187.t2 a_10429_1050.t7 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_4569_1050.t2 a_4891_989.t7 VDD.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_13757_1051.t3 a_3303_411.t8 QN.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 VDD.t23 a_9183_989.t6 a_10429_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 VDD.t41 a_147_187.t9 a_3303_411.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_7595_411.t3 a_7469_1050.t7 VDD.t56 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 VDD.t28 a_4569_1050.t8 a_7469_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 QN a_3303_411.t13 a_13654_101.t0 nshort w=-1.235u l=1.535u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_4439_187.t1 CLK.t7 VDD.t60 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_1845_1050.t2 a_147_187.t10 VDD.t75 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1059 a_8861_1050.t3 a_9183_989.t7 VDD.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1060 VDD.t31 a_4439_187.t10 a_4569_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 a_6137_1050.t2 a_4439_187.t11 VDD.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 GND a_3177_1050.t6 a_3738_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1063 GND a_4569_1050.t10 a_7364_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1064 a_9183_989.t3 a_8861_1050.t10 VDD.t57 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 GND a_9183_989.t8 a_10324_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1066 a_13093_1051.t5 a_3303_411.t9 a_13757_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_11761_1050.t1 a_11887_411.t9 VDD.t51 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_3303_411.t0 a_147_187.t11 VDD.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 VDD.t47 a_7595_411.t10 a_13093_1051.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 VDD.t11 D.t5 a_599_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 a_8731_187.t1 CLK.t9 VDD.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1072 a_13757_1051.t4 a_11887_411.t11 a_13093_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1073 VDD.t67 a_8731_187.t11 a_10429_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1074 a_277_1050.t5 a_147_187.t12 VDD.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 VDD.t55 a_7595_411.t11 a_7469_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1076 a_4439_187.t4 a_6137_1050.t6 VDD.t36 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 GND a_277_1050.t9 a_1074_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1078 VDD.t59 CLK.t12 a_4569_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 VDD.t45 a_599_989.t9 a_1845_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 a_11761_1050.t4 a_8861_1050.t11 VDD.t72 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 VDD.t54 a_11887_411.t12 a_13093_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1082 a_4891_989.t0 D.t7 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 GND a_11761_1050.t7 a_12322_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1084 a_13757_1051.t0 a_3303_411.t10 a_13093_1051.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 a_277_1050.t0 CLK.t13 VDD.t79 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 VDD.t52 a_4891_989.t8 a_4569_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 VDD.t77 a_277_1050.t10 a_3177_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 a_147_187.t2 CLK.t15 VDD.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 VDD.t29 a_11761_1050.t6 a_11887_411.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 GND a_6137_1050.t7 a_6698_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1091 QN a_7595_411.t12 a_12988_101.t1 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1092 GND a_277_1050.t12 a_3072_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1093 a_4891_989.t3 a_4569_1050.t11 VDD.t53 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 a_7595_411.t2 a_4439_187.t12 VDD.t50 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1095 GND a_4891_989.t10 a_6032_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1096 a_277_1050.t3 a_599_989.t10 VDD.t71 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 a_599_989.t1 a_277_1050.t11 VDD.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 GND a_3303_411.t5 a_14320_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1099 QN.t1 a_3303_411.t11 a_13757_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 a_8861_1050.t0 a_8731_187.t12 VDD.t66 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1101 VDD.t48 CLK.t16 a_8731_187.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 a_10429_1050.t1 a_9183_989.t10 VDD.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_7469_1050.t4 a_4569_1050.t12 VDD.t49 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 a_147_187.t1 a_1845_1050.t7 VDD.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 VDD.t46 a_3303_411.t12 a_3177_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 VDD.t65 a_8731_187.t13 a_11887_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 VDD.t58 CLK.t17 a_8861_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 a_4569_1050.t5 a_4439_187.t13 VDD.t63 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 VDD.t76 a_4891_989.t9 a_6137_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 VDD.t15 a_8861_1050.t12 a_11761_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 GND a_8731_187.t7 a_8675_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1112 VDD.t78 a_3177_1050.t7 a_3303_411.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1113 a_13093_1051.t6 a_7595_411.t13 VDD.t34 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VDD CLK 1.74fF
C1 VDD D 0.22fF
C2 VDD QN 0.29fF
C3 CLK D 0.45fF
R0 D.n5 D.t5 472.359
R1 D.n2 D.t3 472.359
R2 D.n0 D.t2 472.359
R3 D.n5 D.t0 384.527
R4 D.n2 D.t7 384.527
R5 D.n0 D.t4 384.527
R6 D.n6 D.n5 216.272
R7 D.n3 D.n2 216.272
R8 D.n1 D.n0 216.272
R9 D.n6 D.t1 141.114
R10 D.n3 D.t8 141.114
R11 D.n1 D.t6 141.114
R12 D.n4 D.n1 91.734
R13 D.n4 D.n3 76
R14 D.n7 D.n6 76
R15 D.n7 D.n4 15.734
R16 D.n7 D 0.046
R17 VDD.n769 VDD.n767 144.705
R18 VDD.n830 VDD.n828 144.705
R19 VDD.n891 VDD.n889 144.705
R20 VDD.n952 VDD.n950 144.705
R21 VDD.n1013 VDD.n1011 144.705
R22 VDD.n1074 VDD.n1072 144.705
R23 VDD.n1155 VDD.n1153 144.705
R24 VDD.n1216 VDD.n1214 144.705
R25 VDD.n1277 VDD.n1275 144.705
R26 VDD.n638 VDD.n636 144.705
R27 VDD.n1338 VDD.n1336 144.705
R28 VDD.n577 VDD.n575 144.705
R29 VDD.n496 VDD.n494 144.705
R30 VDD.n435 VDD.n433 144.705
R31 VDD.n374 VDD.n372 144.705
R32 VDD.n313 VDD.n311 144.705
R33 VDD.n252 VDD.n250 144.705
R34 VDD.n191 VDD.n189 144.705
R35 VDD.n130 VDD.n128 144.705
R36 VDD.n76 VDD.n74 144.705
R37 VDD.n39 VDD.n38 76
R38 VDD.n43 VDD.n42 76
R39 VDD.n47 VDD.n46 76
R40 VDD.n51 VDD.n50 76
R41 VDD.n78 VDD.n77 76
R42 VDD.n82 VDD.n81 76
R43 VDD.n86 VDD.n85 76
R44 VDD.n90 VDD.n89 76
R45 VDD.n94 VDD.n93 76
R46 VDD.n98 VDD.n97 76
R47 VDD.n102 VDD.n101 76
R48 VDD.n106 VDD.n105 76
R49 VDD.n132 VDD.n131 76
R50 VDD.n137 VDD.n136 76
R51 VDD.n142 VDD.n141 76
R52 VDD.n148 VDD.n147 76
R53 VDD.n153 VDD.n152 76
R54 VDD.n158 VDD.n157 76
R55 VDD.n163 VDD.n162 76
R56 VDD.n167 VDD.n166 76
R57 VDD.n193 VDD.n192 76
R58 VDD.n198 VDD.n197 76
R59 VDD.n203 VDD.n202 76
R60 VDD.n209 VDD.n208 76
R61 VDD.n214 VDD.n213 76
R62 VDD.n219 VDD.n218 76
R63 VDD.n224 VDD.n223 76
R64 VDD.n228 VDD.n227 76
R65 VDD.n254 VDD.n253 76
R66 VDD.n259 VDD.n258 76
R67 VDD.n264 VDD.n263 76
R68 VDD.n270 VDD.n269 76
R69 VDD.n275 VDD.n274 76
R70 VDD.n280 VDD.n279 76
R71 VDD.n285 VDD.n284 76
R72 VDD.n289 VDD.n288 76
R73 VDD.n315 VDD.n314 76
R74 VDD.n320 VDD.n319 76
R75 VDD.n325 VDD.n324 76
R76 VDD.n331 VDD.n330 76
R77 VDD.n336 VDD.n335 76
R78 VDD.n341 VDD.n340 76
R79 VDD.n346 VDD.n345 76
R80 VDD.n350 VDD.n349 76
R81 VDD.n376 VDD.n375 76
R82 VDD.n381 VDD.n380 76
R83 VDD.n386 VDD.n385 76
R84 VDD.n392 VDD.n391 76
R85 VDD.n397 VDD.n396 76
R86 VDD.n402 VDD.n401 76
R87 VDD.n407 VDD.n406 76
R88 VDD.n411 VDD.n410 76
R89 VDD.n437 VDD.n436 76
R90 VDD.n442 VDD.n441 76
R91 VDD.n447 VDD.n446 76
R92 VDD.n453 VDD.n452 76
R93 VDD.n458 VDD.n457 76
R94 VDD.n463 VDD.n462 76
R95 VDD.n468 VDD.n467 76
R96 VDD.n472 VDD.n471 76
R97 VDD.n498 VDD.n497 76
R98 VDD.n502 VDD.n501 76
R99 VDD.n506 VDD.n505 76
R100 VDD.n511 VDD.n510 76
R101 VDD.n518 VDD.n517 76
R102 VDD.n523 VDD.n522 76
R103 VDD.n528 VDD.n527 76
R104 VDD.n535 VDD.n534 76
R105 VDD.n540 VDD.n539 76
R106 VDD.n545 VDD.n544 76
R107 VDD.n549 VDD.n548 76
R108 VDD.n553 VDD.n552 76
R109 VDD.n579 VDD.n578 76
R110 VDD.n584 VDD.n583 76
R111 VDD.n589 VDD.n588 76
R112 VDD.n595 VDD.n594 76
R113 VDD.n600 VDD.n599 76
R114 VDD.n605 VDD.n604 76
R115 VDD.n610 VDD.n609 76
R116 VDD.n614 VDD.n613 76
R117 VDD.n640 VDD.n639 76
R118 VDD.n645 VDD.n644 76
R119 VDD.n650 VDD.n649 76
R120 VDD.n656 VDD.n655 76
R121 VDD.n661 VDD.n660 76
R122 VDD.n666 VDD.n665 76
R123 VDD.n1345 VDD.n1344 76
R124 VDD.n1340 VDD.n1339 76
R125 VDD.n1314 VDD.n1313 76
R126 VDD.n1310 VDD.n1309 76
R127 VDD.n1305 VDD.n1304 76
R128 VDD.n1300 VDD.n1299 76
R129 VDD.n1294 VDD.n1293 76
R130 VDD.n1289 VDD.n1288 76
R131 VDD.n1284 VDD.n1283 76
R132 VDD.n1279 VDD.n1278 76
R133 VDD.n1253 VDD.n1252 76
R134 VDD.n1249 VDD.n1248 76
R135 VDD.n1244 VDD.n1243 76
R136 VDD.n1239 VDD.n1238 76
R137 VDD.n1233 VDD.n1232 76
R138 VDD.n1228 VDD.n1227 76
R139 VDD.n1223 VDD.n1222 76
R140 VDD.n1218 VDD.n1217 76
R141 VDD.n1192 VDD.n1191 76
R142 VDD.n1188 VDD.n1187 76
R143 VDD.n1183 VDD.n1182 76
R144 VDD.n1178 VDD.n1177 76
R145 VDD.n1172 VDD.n1171 76
R146 VDD.n1167 VDD.n1166 76
R147 VDD.n1162 VDD.n1161 76
R148 VDD.n1157 VDD.n1156 76
R149 VDD.n1131 VDD.n1130 76
R150 VDD.n1127 VDD.n1126 76
R151 VDD.n1123 VDD.n1122 76
R152 VDD.n1119 VDD.n1118 76
R153 VDD.n1114 VDD.n1113 76
R154 VDD.n1107 VDD.n1106 76
R155 VDD.n1102 VDD.n1101 76
R156 VDD.n1097 VDD.n1096 76
R157 VDD.n1090 VDD.n1089 76
R158 VDD.n1085 VDD.n1084 76
R159 VDD.n1080 VDD.n1079 76
R160 VDD.n1076 VDD.n1075 76
R161 VDD.n1050 VDD.n1049 76
R162 VDD.n1046 VDD.n1045 76
R163 VDD.n1041 VDD.n1040 76
R164 VDD.n1036 VDD.n1035 76
R165 VDD.n1030 VDD.n1029 76
R166 VDD.n1025 VDD.n1024 76
R167 VDD.n1020 VDD.n1019 76
R168 VDD.n1015 VDD.n1014 76
R169 VDD.n989 VDD.n988 76
R170 VDD.n985 VDD.n984 76
R171 VDD.n980 VDD.n979 76
R172 VDD.n975 VDD.n974 76
R173 VDD.n969 VDD.n968 76
R174 VDD.n964 VDD.n963 76
R175 VDD.n959 VDD.n958 76
R176 VDD.n954 VDD.n953 76
R177 VDD.n928 VDD.n927 76
R178 VDD.n924 VDD.n923 76
R179 VDD.n919 VDD.n918 76
R180 VDD.n914 VDD.n913 76
R181 VDD.n908 VDD.n907 76
R182 VDD.n903 VDD.n902 76
R183 VDD.n898 VDD.n897 76
R184 VDD.n893 VDD.n892 76
R185 VDD.n867 VDD.n866 76
R186 VDD.n863 VDD.n862 76
R187 VDD.n858 VDD.n857 76
R188 VDD.n853 VDD.n852 76
R189 VDD.n847 VDD.n846 76
R190 VDD.n842 VDD.n841 76
R191 VDD.n837 VDD.n836 76
R192 VDD.n832 VDD.n831 76
R193 VDD.n806 VDD.n805 76
R194 VDD.n802 VDD.n801 76
R195 VDD.n797 VDD.n796 76
R196 VDD.n792 VDD.n791 76
R197 VDD.n786 VDD.n785 76
R198 VDD.n781 VDD.n780 76
R199 VDD.n776 VDD.n775 76
R200 VDD.n771 VDD.n770 76
R201 VDD.n744 VDD.n743 76
R202 VDD.n740 VDD.n739 76
R203 VDD.n736 VDD.n735 76
R204 VDD.n732 VDD.n731 76
R205 VDD.n727 VDD.n726 76
R206 VDD.n720 VDD.n719 76
R207 VDD.n715 VDD.n714 76
R208 VDD.n710 VDD.n709 76
R209 VDD.n703 VDD.n702 76
R210 VDD.n698 VDD.n697 76
R211 VDD.n693 VDD.n692 76
R212 VDD.n689 VDD.n688 76
R213 VDD.n508 VDD.n507 64.064
R214 VDD.n1116 VDD.n1115 64.064
R215 VDD.n729 VDD.n728 64.064
R216 VDD.n537 VDD.n536 59.488
R217 VDD.n1087 VDD.n1086 59.488
R218 VDD.n700 VDD.n699 59.488
R219 VDD.n159 VDD.t40 55.465
R220 VDD.n133 VDD.t47 55.465
R221 VDD.n694 VDD.t13 55.106
R222 VDD.n772 VDD.t6 55.106
R223 VDD.n833 VDD.t3 55.106
R224 VDD.n894 VDD.t19 55.106
R225 VDD.n955 VDD.t18 55.106
R226 VDD.n1016 VDD.t37 55.106
R227 VDD.n1081 VDD.t63 55.106
R228 VDD.n1158 VDD.t53 55.106
R229 VDD.n1219 VDD.t0 55.106
R230 VDD.n1280 VDD.t36 55.106
R231 VDD.n1341 VDD.t49 55.106
R232 VDD.n606 VDD.t56 55.106
R233 VDD.n541 VDD.t66 55.106
R234 VDD.n464 VDD.t57 55.106
R235 VDD.n403 VDD.t24 55.106
R236 VDD.n342 VDD.t5 55.106
R237 VDD.n281 VDD.t72 55.106
R238 VDD.n220 VDD.t35 55.106
R239 VDD.n735 VDD.t33 55.106
R240 VDD.n1122 VDD.t52 55.106
R241 VDD.n505 VDD.t26 55.106
R242 VDD.n798 VDD.t11 55.106
R243 VDD.n859 VDD.t14 55.106
R244 VDD.n920 VDD.t21 55.106
R245 VDD.n981 VDD.t46 55.106
R246 VDD.n1042 VDD.t41 55.106
R247 VDD.n1184 VDD.t12 55.106
R248 VDD.n1245 VDD.t64 55.106
R249 VDD.n1306 VDD.t38 55.106
R250 VDD.n641 VDD.t55 55.106
R251 VDD.n580 VDD.t32 55.106
R252 VDD.n438 VDD.t7 55.106
R253 VDD.n377 VDD.t67 55.106
R254 VDD.n316 VDD.t48 55.106
R255 VDD.n255 VDD.t16 55.106
R256 VDD.n194 VDD.t65 55.106
R257 VDD.n144 VDD.n143 41.183
R258 VDD.n705 VDD.n704 40.824
R259 VDD.n725 VDD.n724 40.824
R260 VDD.n788 VDD.n787 40.824
R261 VDD.n849 VDD.n848 40.824
R262 VDD.n910 VDD.n909 40.824
R263 VDD.n971 VDD.n970 40.824
R264 VDD.n1032 VDD.n1031 40.824
R265 VDD.n1092 VDD.n1091 40.824
R266 VDD.n1112 VDD.n1111 40.824
R267 VDD.n1174 VDD.n1173 40.824
R268 VDD.n1235 VDD.n1234 40.824
R269 VDD.n1296 VDD.n1295 40.824
R270 VDD.n652 VDD.n651 40.824
R271 VDD.n591 VDD.n590 40.824
R272 VDD.n530 VDD.n529 40.824
R273 VDD.n516 VDD.n515 40.824
R274 VDD.n449 VDD.n448 40.824
R275 VDD.n388 VDD.n387 40.824
R276 VDD.n327 VDD.n326 40.824
R277 VDD.n266 VDD.n265 40.824
R278 VDD.n205 VDD.n204 40.824
R279 VDD.n811 VDD.n810 36.774
R280 VDD.n872 VDD.n871 36.774
R281 VDD.n933 VDD.n932 36.774
R282 VDD.n994 VDD.n993 36.774
R283 VDD.n1055 VDD.n1054 36.774
R284 VDD.n1136 VDD.n1135 36.774
R285 VDD.n1197 VDD.n1196 36.774
R286 VDD.n1258 VDD.n1257 36.774
R287 VDD.n1319 VDD.n1318 36.774
R288 VDD.n619 VDD.n618 36.774
R289 VDD.n558 VDD.n557 36.774
R290 VDD.n477 VDD.n476 36.774
R291 VDD.n416 VDD.n415 36.774
R292 VDD.n355 VDD.n354 36.774
R293 VDD.n294 VDD.n293 36.774
R294 VDD.n233 VDD.n232 36.774
R295 VDD.n172 VDD.n171 36.774
R296 VDD.n111 VDD.n110 36.774
R297 VDD.n56 VDD.n55 36.774
R298 VDD.n760 VDD.n759 36.774
R299 VDD.n139 VDD.n138 36.608
R300 VDD.n200 VDD.n199 36.608
R301 VDD.n261 VDD.n260 36.608
R302 VDD.n322 VDD.n321 36.608
R303 VDD.n383 VDD.n382 36.608
R304 VDD.n444 VDD.n443 36.608
R305 VDD.n586 VDD.n585 36.608
R306 VDD.n647 VDD.n646 36.608
R307 VDD.n1302 VDD.n1301 36.608
R308 VDD.n1241 VDD.n1240 36.608
R309 VDD.n1180 VDD.n1179 36.608
R310 VDD.n1038 VDD.n1037 36.608
R311 VDD.n977 VDD.n976 36.608
R312 VDD.n916 VDD.n915 36.608
R313 VDD.n855 VDD.n854 36.608
R314 VDD.n794 VDD.n793 36.608
R315 VDD.n34 VDD.n33 34.942
R316 VDD.n155 VDD.n154 32.032
R317 VDD.n216 VDD.n215 32.032
R318 VDD.n277 VDD.n276 32.032
R319 VDD.n338 VDD.n337 32.032
R320 VDD.n399 VDD.n398 32.032
R321 VDD.n460 VDD.n459 32.032
R322 VDD.n602 VDD.n601 32.032
R323 VDD.n663 VDD.n662 32.032
R324 VDD.n1286 VDD.n1285 32.032
R325 VDD.n1225 VDD.n1224 32.032
R326 VDD.n1164 VDD.n1163 32.032
R327 VDD.n1022 VDD.n1021 32.032
R328 VDD.n961 VDD.n960 32.032
R329 VDD.n900 VDD.n899 32.032
R330 VDD.n839 VDD.n838 32.032
R331 VDD.n778 VDD.n777 32.032
R332 VDD.n513 VDD.n512 27.456
R333 VDD.n1109 VDD.n1108 27.456
R334 VDD.n722 VDD.n721 27.456
R335 VDD.n532 VDD.n531 22.88
R336 VDD.n1094 VDD.n1093 22.88
R337 VDD.n707 VDD.n706 22.88
R338 VDD.n688 VDD.n685 21.841
R339 VDD.n23 VDD.n20 21.841
R340 VDD.n704 VDD.t79 14.282
R341 VDD.n704 VDD.t42 14.282
R342 VDD.n724 VDD.t71 14.282
R343 VDD.n724 VDD.t61 14.282
R344 VDD.n787 VDD.t10 14.282
R345 VDD.n787 VDD.t1 14.282
R346 VDD.n848 VDD.t75 14.282
R347 VDD.n848 VDD.t45 14.282
R348 VDD.n909 VDD.t20 14.282
R349 VDD.n909 VDD.t2 14.282
R350 VDD.n970 VDD.t44 14.282
R351 VDD.n970 VDD.t77 14.282
R352 VDD.n1031 VDD.t4 14.282
R353 VDD.n1031 VDD.t78 14.282
R354 VDD.n1091 VDD.t80 14.282
R355 VDD.n1091 VDD.t31 14.282
R356 VDD.n1111 VDD.t17 14.282
R357 VDD.n1111 VDD.t59 14.282
R358 VDD.n1173 VDD.t8 14.282
R359 VDD.n1173 VDD.t62 14.282
R360 VDD.n1234 VDD.t22 14.282
R361 VDD.n1234 VDD.t76 14.282
R362 VDD.n1295 VDD.t60 14.282
R363 VDD.n1295 VDD.t27 14.282
R364 VDD.n651 VDD.t74 14.282
R365 VDD.n651 VDD.t28 14.282
R366 VDD.n590 VDD.t50 14.282
R367 VDD.n590 VDD.t43 14.282
R368 VDD.n529 VDD.t39 14.282
R369 VDD.n529 VDD.t69 14.282
R370 VDD.n515 VDD.t25 14.282
R371 VDD.n515 VDD.t58 14.282
R372 VDD.n448 VDD.t9 14.282
R373 VDD.n448 VDD.t73 14.282
R374 VDD.n387 VDD.t70 14.282
R375 VDD.n387 VDD.t23 14.282
R376 VDD.n326 VDD.t30 14.282
R377 VDD.n326 VDD.t81 14.282
R378 VDD.n265 VDD.t51 14.282
R379 VDD.n265 VDD.t15 14.282
R380 VDD.n204 VDD.t68 14.282
R381 VDD.n204 VDD.t29 14.282
R382 VDD.n143 VDD.t34 14.282
R383 VDD.n143 VDD.t54 14.282
R384 VDD.n685 VDD.n668 14.167
R385 VDD.n668 VDD.n667 14.167
R386 VDD.n826 VDD.n808 14.167
R387 VDD.n808 VDD.n807 14.167
R388 VDD.n887 VDD.n869 14.167
R389 VDD.n869 VDD.n868 14.167
R390 VDD.n948 VDD.n930 14.167
R391 VDD.n930 VDD.n929 14.167
R392 VDD.n1009 VDD.n991 14.167
R393 VDD.n991 VDD.n990 14.167
R394 VDD.n1070 VDD.n1052 14.167
R395 VDD.n1052 VDD.n1051 14.167
R396 VDD.n1151 VDD.n1133 14.167
R397 VDD.n1133 VDD.n1132 14.167
R398 VDD.n1212 VDD.n1194 14.167
R399 VDD.n1194 VDD.n1193 14.167
R400 VDD.n1273 VDD.n1255 14.167
R401 VDD.n1255 VDD.n1254 14.167
R402 VDD.n1334 VDD.n1316 14.167
R403 VDD.n1316 VDD.n1315 14.167
R404 VDD.n634 VDD.n616 14.167
R405 VDD.n616 VDD.n615 14.167
R406 VDD.n573 VDD.n555 14.167
R407 VDD.n555 VDD.n554 14.167
R408 VDD.n492 VDD.n474 14.167
R409 VDD.n474 VDD.n473 14.167
R410 VDD.n431 VDD.n413 14.167
R411 VDD.n413 VDD.n412 14.167
R412 VDD.n370 VDD.n352 14.167
R413 VDD.n352 VDD.n351 14.167
R414 VDD.n309 VDD.n291 14.167
R415 VDD.n291 VDD.n290 14.167
R416 VDD.n248 VDD.n230 14.167
R417 VDD.n230 VDD.n229 14.167
R418 VDD.n187 VDD.n169 14.167
R419 VDD.n169 VDD.n168 14.167
R420 VDD.n126 VDD.n108 14.167
R421 VDD.n108 VDD.n107 14.167
R422 VDD.n72 VDD.n53 14.167
R423 VDD.n53 VDD.n52 14.167
R424 VDD.n765 VDD.n746 14.167
R425 VDD.n746 VDD.n745 14.167
R426 VDD.n20 VDD.n19 14.167
R427 VDD.n19 VDD.n17 14.167
R428 VDD.n32 VDD.n29 14.167
R429 VDD.n29 VDD.n28 14.167
R430 VDD.n77 VDD.n73 14.167
R431 VDD.n131 VDD.n127 14.167
R432 VDD.n192 VDD.n188 14.167
R433 VDD.n253 VDD.n249 14.167
R434 VDD.n314 VDD.n310 14.167
R435 VDD.n375 VDD.n371 14.167
R436 VDD.n436 VDD.n432 14.167
R437 VDD.n497 VDD.n493 14.167
R438 VDD.n578 VDD.n574 14.167
R439 VDD.n639 VDD.n635 14.167
R440 VDD.n1339 VDD.n1335 14.167
R441 VDD.n1278 VDD.n1274 14.167
R442 VDD.n1217 VDD.n1213 14.167
R443 VDD.n1156 VDD.n1152 14.167
R444 VDD.n1075 VDD.n1071 14.167
R445 VDD.n1014 VDD.n1010 14.167
R446 VDD.n953 VDD.n949 14.167
R447 VDD.n892 VDD.n888 14.167
R448 VDD.n831 VDD.n827 14.167
R449 VDD.n770 VDD.n766 14.167
R450 VDD.n525 VDD.n524 13.728
R451 VDD.n1099 VDD.n1098 13.728
R452 VDD.n712 VDD.n711 13.728
R453 VDD.n23 VDD.n22 13.653
R454 VDD.n22 VDD.n21 13.653
R455 VDD.n32 VDD.n31 13.653
R456 VDD.n31 VDD.n30 13.653
R457 VDD.n29 VDD.n25 13.653
R458 VDD.n25 VDD.n24 13.653
R459 VDD.n28 VDD.n27 13.653
R460 VDD.n27 VDD.n26 13.653
R461 VDD.n38 VDD.n37 13.653
R462 VDD.n37 VDD.n36 13.653
R463 VDD.n42 VDD.n41 13.653
R464 VDD.n41 VDD.n40 13.653
R465 VDD.n46 VDD.n45 13.653
R466 VDD.n45 VDD.n44 13.653
R467 VDD.n50 VDD.n49 13.653
R468 VDD.n49 VDD.n48 13.653
R469 VDD.n77 VDD.n76 13.653
R470 VDD.n76 VDD.n75 13.653
R471 VDD.n81 VDD.n80 13.653
R472 VDD.n80 VDD.n79 13.653
R473 VDD.n85 VDD.n84 13.653
R474 VDD.n84 VDD.n83 13.653
R475 VDD.n89 VDD.n88 13.653
R476 VDD.n88 VDD.n87 13.653
R477 VDD.n93 VDD.n92 13.653
R478 VDD.n92 VDD.n91 13.653
R479 VDD.n97 VDD.n96 13.653
R480 VDD.n96 VDD.n95 13.653
R481 VDD.n101 VDD.n100 13.653
R482 VDD.n100 VDD.n99 13.653
R483 VDD.n105 VDD.n104 13.653
R484 VDD.n104 VDD.n103 13.653
R485 VDD.n131 VDD.n130 13.653
R486 VDD.n130 VDD.n129 13.653
R487 VDD.n136 VDD.n135 13.653
R488 VDD.n135 VDD.n134 13.653
R489 VDD.n141 VDD.n140 13.653
R490 VDD.n140 VDD.n139 13.653
R491 VDD.n147 VDD.n146 13.653
R492 VDD.n146 VDD.n145 13.653
R493 VDD.n152 VDD.n151 13.653
R494 VDD.n151 VDD.n150 13.653
R495 VDD.n157 VDD.n156 13.653
R496 VDD.n156 VDD.n155 13.653
R497 VDD.n162 VDD.n161 13.653
R498 VDD.n161 VDD.n160 13.653
R499 VDD.n166 VDD.n165 13.653
R500 VDD.n165 VDD.n164 13.653
R501 VDD.n192 VDD.n191 13.653
R502 VDD.n191 VDD.n190 13.653
R503 VDD.n197 VDD.n196 13.653
R504 VDD.n196 VDD.n195 13.653
R505 VDD.n202 VDD.n201 13.653
R506 VDD.n201 VDD.n200 13.653
R507 VDD.n208 VDD.n207 13.653
R508 VDD.n207 VDD.n206 13.653
R509 VDD.n213 VDD.n212 13.653
R510 VDD.n212 VDD.n211 13.653
R511 VDD.n218 VDD.n217 13.653
R512 VDD.n217 VDD.n216 13.653
R513 VDD.n223 VDD.n222 13.653
R514 VDD.n222 VDD.n221 13.653
R515 VDD.n227 VDD.n226 13.653
R516 VDD.n226 VDD.n225 13.653
R517 VDD.n253 VDD.n252 13.653
R518 VDD.n252 VDD.n251 13.653
R519 VDD.n258 VDD.n257 13.653
R520 VDD.n257 VDD.n256 13.653
R521 VDD.n263 VDD.n262 13.653
R522 VDD.n262 VDD.n261 13.653
R523 VDD.n269 VDD.n268 13.653
R524 VDD.n268 VDD.n267 13.653
R525 VDD.n274 VDD.n273 13.653
R526 VDD.n273 VDD.n272 13.653
R527 VDD.n279 VDD.n278 13.653
R528 VDD.n278 VDD.n277 13.653
R529 VDD.n284 VDD.n283 13.653
R530 VDD.n283 VDD.n282 13.653
R531 VDD.n288 VDD.n287 13.653
R532 VDD.n287 VDD.n286 13.653
R533 VDD.n314 VDD.n313 13.653
R534 VDD.n313 VDD.n312 13.653
R535 VDD.n319 VDD.n318 13.653
R536 VDD.n318 VDD.n317 13.653
R537 VDD.n324 VDD.n323 13.653
R538 VDD.n323 VDD.n322 13.653
R539 VDD.n330 VDD.n329 13.653
R540 VDD.n329 VDD.n328 13.653
R541 VDD.n335 VDD.n334 13.653
R542 VDD.n334 VDD.n333 13.653
R543 VDD.n340 VDD.n339 13.653
R544 VDD.n339 VDD.n338 13.653
R545 VDD.n345 VDD.n344 13.653
R546 VDD.n344 VDD.n343 13.653
R547 VDD.n349 VDD.n348 13.653
R548 VDD.n348 VDD.n347 13.653
R549 VDD.n375 VDD.n374 13.653
R550 VDD.n374 VDD.n373 13.653
R551 VDD.n380 VDD.n379 13.653
R552 VDD.n379 VDD.n378 13.653
R553 VDD.n385 VDD.n384 13.653
R554 VDD.n384 VDD.n383 13.653
R555 VDD.n391 VDD.n390 13.653
R556 VDD.n390 VDD.n389 13.653
R557 VDD.n396 VDD.n395 13.653
R558 VDD.n395 VDD.n394 13.653
R559 VDD.n401 VDD.n400 13.653
R560 VDD.n400 VDD.n399 13.653
R561 VDD.n406 VDD.n405 13.653
R562 VDD.n405 VDD.n404 13.653
R563 VDD.n410 VDD.n409 13.653
R564 VDD.n409 VDD.n408 13.653
R565 VDD.n436 VDD.n435 13.653
R566 VDD.n435 VDD.n434 13.653
R567 VDD.n441 VDD.n440 13.653
R568 VDD.n440 VDD.n439 13.653
R569 VDD.n446 VDD.n445 13.653
R570 VDD.n445 VDD.n444 13.653
R571 VDD.n452 VDD.n451 13.653
R572 VDD.n451 VDD.n450 13.653
R573 VDD.n457 VDD.n456 13.653
R574 VDD.n456 VDD.n455 13.653
R575 VDD.n462 VDD.n461 13.653
R576 VDD.n461 VDD.n460 13.653
R577 VDD.n467 VDD.n466 13.653
R578 VDD.n466 VDD.n465 13.653
R579 VDD.n471 VDD.n470 13.653
R580 VDD.n470 VDD.n469 13.653
R581 VDD.n497 VDD.n496 13.653
R582 VDD.n496 VDD.n495 13.653
R583 VDD.n501 VDD.n500 13.653
R584 VDD.n500 VDD.n499 13.653
R585 VDD.n505 VDD.n504 13.653
R586 VDD.n504 VDD.n503 13.653
R587 VDD.n510 VDD.n509 13.653
R588 VDD.n509 VDD.n508 13.653
R589 VDD.n517 VDD.n514 13.653
R590 VDD.n514 VDD.n513 13.653
R591 VDD.n522 VDD.n521 13.653
R592 VDD.n521 VDD.n520 13.653
R593 VDD.n527 VDD.n526 13.653
R594 VDD.n526 VDD.n525 13.653
R595 VDD.n534 VDD.n533 13.653
R596 VDD.n533 VDD.n532 13.653
R597 VDD.n539 VDD.n538 13.653
R598 VDD.n538 VDD.n537 13.653
R599 VDD.n544 VDD.n543 13.653
R600 VDD.n543 VDD.n542 13.653
R601 VDD.n548 VDD.n547 13.653
R602 VDD.n547 VDD.n546 13.653
R603 VDD.n552 VDD.n551 13.653
R604 VDD.n551 VDD.n550 13.653
R605 VDD.n578 VDD.n577 13.653
R606 VDD.n577 VDD.n576 13.653
R607 VDD.n583 VDD.n582 13.653
R608 VDD.n582 VDD.n581 13.653
R609 VDD.n588 VDD.n587 13.653
R610 VDD.n587 VDD.n586 13.653
R611 VDD.n594 VDD.n593 13.653
R612 VDD.n593 VDD.n592 13.653
R613 VDD.n599 VDD.n598 13.653
R614 VDD.n598 VDD.n597 13.653
R615 VDD.n604 VDD.n603 13.653
R616 VDD.n603 VDD.n602 13.653
R617 VDD.n609 VDD.n608 13.653
R618 VDD.n608 VDD.n607 13.653
R619 VDD.n613 VDD.n612 13.653
R620 VDD.n612 VDD.n611 13.653
R621 VDD.n639 VDD.n638 13.653
R622 VDD.n638 VDD.n637 13.653
R623 VDD.n644 VDD.n643 13.653
R624 VDD.n643 VDD.n642 13.653
R625 VDD.n649 VDD.n648 13.653
R626 VDD.n648 VDD.n647 13.653
R627 VDD.n655 VDD.n654 13.653
R628 VDD.n654 VDD.n653 13.653
R629 VDD.n660 VDD.n659 13.653
R630 VDD.n659 VDD.n658 13.653
R631 VDD.n665 VDD.n664 13.653
R632 VDD.n664 VDD.n663 13.653
R633 VDD.n1344 VDD.n1343 13.653
R634 VDD.n1343 VDD.n1342 13.653
R635 VDD.n1339 VDD.n1338 13.653
R636 VDD.n1338 VDD.n1337 13.653
R637 VDD.n1313 VDD.n1312 13.653
R638 VDD.n1312 VDD.n1311 13.653
R639 VDD.n1309 VDD.n1308 13.653
R640 VDD.n1308 VDD.n1307 13.653
R641 VDD.n1304 VDD.n1303 13.653
R642 VDD.n1303 VDD.n1302 13.653
R643 VDD.n1299 VDD.n1298 13.653
R644 VDD.n1298 VDD.n1297 13.653
R645 VDD.n1293 VDD.n1292 13.653
R646 VDD.n1292 VDD.n1291 13.653
R647 VDD.n1288 VDD.n1287 13.653
R648 VDD.n1287 VDD.n1286 13.653
R649 VDD.n1283 VDD.n1282 13.653
R650 VDD.n1282 VDD.n1281 13.653
R651 VDD.n1278 VDD.n1277 13.653
R652 VDD.n1277 VDD.n1276 13.653
R653 VDD.n1252 VDD.n1251 13.653
R654 VDD.n1251 VDD.n1250 13.653
R655 VDD.n1248 VDD.n1247 13.653
R656 VDD.n1247 VDD.n1246 13.653
R657 VDD.n1243 VDD.n1242 13.653
R658 VDD.n1242 VDD.n1241 13.653
R659 VDD.n1238 VDD.n1237 13.653
R660 VDD.n1237 VDD.n1236 13.653
R661 VDD.n1232 VDD.n1231 13.653
R662 VDD.n1231 VDD.n1230 13.653
R663 VDD.n1227 VDD.n1226 13.653
R664 VDD.n1226 VDD.n1225 13.653
R665 VDD.n1222 VDD.n1221 13.653
R666 VDD.n1221 VDD.n1220 13.653
R667 VDD.n1217 VDD.n1216 13.653
R668 VDD.n1216 VDD.n1215 13.653
R669 VDD.n1191 VDD.n1190 13.653
R670 VDD.n1190 VDD.n1189 13.653
R671 VDD.n1187 VDD.n1186 13.653
R672 VDD.n1186 VDD.n1185 13.653
R673 VDD.n1182 VDD.n1181 13.653
R674 VDD.n1181 VDD.n1180 13.653
R675 VDD.n1177 VDD.n1176 13.653
R676 VDD.n1176 VDD.n1175 13.653
R677 VDD.n1171 VDD.n1170 13.653
R678 VDD.n1170 VDD.n1169 13.653
R679 VDD.n1166 VDD.n1165 13.653
R680 VDD.n1165 VDD.n1164 13.653
R681 VDD.n1161 VDD.n1160 13.653
R682 VDD.n1160 VDD.n1159 13.653
R683 VDD.n1156 VDD.n1155 13.653
R684 VDD.n1155 VDD.n1154 13.653
R685 VDD.n1130 VDD.n1129 13.653
R686 VDD.n1129 VDD.n1128 13.653
R687 VDD.n1126 VDD.n1125 13.653
R688 VDD.n1125 VDD.n1124 13.653
R689 VDD.n1122 VDD.n1121 13.653
R690 VDD.n1121 VDD.n1120 13.653
R691 VDD.n1118 VDD.n1117 13.653
R692 VDD.n1117 VDD.n1116 13.653
R693 VDD.n1113 VDD.n1110 13.653
R694 VDD.n1110 VDD.n1109 13.653
R695 VDD.n1106 VDD.n1105 13.653
R696 VDD.n1105 VDD.n1104 13.653
R697 VDD.n1101 VDD.n1100 13.653
R698 VDD.n1100 VDD.n1099 13.653
R699 VDD.n1096 VDD.n1095 13.653
R700 VDD.n1095 VDD.n1094 13.653
R701 VDD.n1089 VDD.n1088 13.653
R702 VDD.n1088 VDD.n1087 13.653
R703 VDD.n1084 VDD.n1083 13.653
R704 VDD.n1083 VDD.n1082 13.653
R705 VDD.n1079 VDD.n1078 13.653
R706 VDD.n1078 VDD.n1077 13.653
R707 VDD.n1075 VDD.n1074 13.653
R708 VDD.n1074 VDD.n1073 13.653
R709 VDD.n1049 VDD.n1048 13.653
R710 VDD.n1048 VDD.n1047 13.653
R711 VDD.n1045 VDD.n1044 13.653
R712 VDD.n1044 VDD.n1043 13.653
R713 VDD.n1040 VDD.n1039 13.653
R714 VDD.n1039 VDD.n1038 13.653
R715 VDD.n1035 VDD.n1034 13.653
R716 VDD.n1034 VDD.n1033 13.653
R717 VDD.n1029 VDD.n1028 13.653
R718 VDD.n1028 VDD.n1027 13.653
R719 VDD.n1024 VDD.n1023 13.653
R720 VDD.n1023 VDD.n1022 13.653
R721 VDD.n1019 VDD.n1018 13.653
R722 VDD.n1018 VDD.n1017 13.653
R723 VDD.n1014 VDD.n1013 13.653
R724 VDD.n1013 VDD.n1012 13.653
R725 VDD.n988 VDD.n987 13.653
R726 VDD.n987 VDD.n986 13.653
R727 VDD.n984 VDD.n983 13.653
R728 VDD.n983 VDD.n982 13.653
R729 VDD.n979 VDD.n978 13.653
R730 VDD.n978 VDD.n977 13.653
R731 VDD.n974 VDD.n973 13.653
R732 VDD.n973 VDD.n972 13.653
R733 VDD.n968 VDD.n967 13.653
R734 VDD.n967 VDD.n966 13.653
R735 VDD.n963 VDD.n962 13.653
R736 VDD.n962 VDD.n961 13.653
R737 VDD.n958 VDD.n957 13.653
R738 VDD.n957 VDD.n956 13.653
R739 VDD.n953 VDD.n952 13.653
R740 VDD.n952 VDD.n951 13.653
R741 VDD.n927 VDD.n926 13.653
R742 VDD.n926 VDD.n925 13.653
R743 VDD.n923 VDD.n922 13.653
R744 VDD.n922 VDD.n921 13.653
R745 VDD.n918 VDD.n917 13.653
R746 VDD.n917 VDD.n916 13.653
R747 VDD.n913 VDD.n912 13.653
R748 VDD.n912 VDD.n911 13.653
R749 VDD.n907 VDD.n906 13.653
R750 VDD.n906 VDD.n905 13.653
R751 VDD.n902 VDD.n901 13.653
R752 VDD.n901 VDD.n900 13.653
R753 VDD.n897 VDD.n896 13.653
R754 VDD.n896 VDD.n895 13.653
R755 VDD.n892 VDD.n891 13.653
R756 VDD.n891 VDD.n890 13.653
R757 VDD.n866 VDD.n865 13.653
R758 VDD.n865 VDD.n864 13.653
R759 VDD.n862 VDD.n861 13.653
R760 VDD.n861 VDD.n860 13.653
R761 VDD.n857 VDD.n856 13.653
R762 VDD.n856 VDD.n855 13.653
R763 VDD.n852 VDD.n851 13.653
R764 VDD.n851 VDD.n850 13.653
R765 VDD.n846 VDD.n845 13.653
R766 VDD.n845 VDD.n844 13.653
R767 VDD.n841 VDD.n840 13.653
R768 VDD.n840 VDD.n839 13.653
R769 VDD.n836 VDD.n835 13.653
R770 VDD.n835 VDD.n834 13.653
R771 VDD.n831 VDD.n830 13.653
R772 VDD.n830 VDD.n829 13.653
R773 VDD.n805 VDD.n804 13.653
R774 VDD.n804 VDD.n803 13.653
R775 VDD.n801 VDD.n800 13.653
R776 VDD.n800 VDD.n799 13.653
R777 VDD.n796 VDD.n795 13.653
R778 VDD.n795 VDD.n794 13.653
R779 VDD.n791 VDD.n790 13.653
R780 VDD.n790 VDD.n789 13.653
R781 VDD.n785 VDD.n784 13.653
R782 VDD.n784 VDD.n783 13.653
R783 VDD.n780 VDD.n779 13.653
R784 VDD.n779 VDD.n778 13.653
R785 VDD.n775 VDD.n774 13.653
R786 VDD.n774 VDD.n773 13.653
R787 VDD.n770 VDD.n769 13.653
R788 VDD.n769 VDD.n768 13.653
R789 VDD.n743 VDD.n742 13.653
R790 VDD.n742 VDD.n741 13.653
R791 VDD.n739 VDD.n738 13.653
R792 VDD.n738 VDD.n737 13.653
R793 VDD.n735 VDD.n734 13.653
R794 VDD.n734 VDD.n733 13.653
R795 VDD.n731 VDD.n730 13.653
R796 VDD.n730 VDD.n729 13.653
R797 VDD.n726 VDD.n723 13.653
R798 VDD.n723 VDD.n722 13.653
R799 VDD.n719 VDD.n718 13.653
R800 VDD.n718 VDD.n717 13.653
R801 VDD.n714 VDD.n713 13.653
R802 VDD.n713 VDD.n712 13.653
R803 VDD.n709 VDD.n708 13.653
R804 VDD.n708 VDD.n707 13.653
R805 VDD.n702 VDD.n701 13.653
R806 VDD.n701 VDD.n700 13.653
R807 VDD.n697 VDD.n696 13.653
R808 VDD.n696 VDD.n695 13.653
R809 VDD.n692 VDD.n691 13.653
R810 VDD.n691 VDD.n690 13.653
R811 VDD.n688 VDD.n687 13.653
R812 VDD.n687 VDD.n686 13.653
R813 VDD.n4 VDD.n2 12.915
R814 VDD.n4 VDD.n3 12.66
R815 VDD.n13 VDD.n12 12.343
R816 VDD.n10 VDD.n9 12.343
R817 VDD.n7 VDD.n6 12.343
R818 VDD.n520 VDD.n519 9.152
R819 VDD.n1104 VDD.n1103 9.152
R820 VDD.n717 VDD.n716 9.152
R821 VDD.n147 VDD.n144 8.658
R822 VDD.n208 VDD.n205 8.658
R823 VDD.n269 VDD.n266 8.658
R824 VDD.n330 VDD.n327 8.658
R825 VDD.n391 VDD.n388 8.658
R826 VDD.n452 VDD.n449 8.658
R827 VDD.n594 VDD.n591 8.658
R828 VDD.n655 VDD.n652 8.658
R829 VDD.n1299 VDD.n1296 8.658
R830 VDD.n1238 VDD.n1235 8.658
R831 VDD.n1177 VDD.n1174 8.658
R832 VDD.n1035 VDD.n1032 8.658
R833 VDD.n974 VDD.n971 8.658
R834 VDD.n913 VDD.n910 8.658
R835 VDD.n852 VDD.n849 8.658
R836 VDD.n791 VDD.n788 8.658
R837 VDD.n827 VDD.n826 7.674
R838 VDD.n888 VDD.n887 7.674
R839 VDD.n949 VDD.n948 7.674
R840 VDD.n1010 VDD.n1009 7.674
R841 VDD.n1071 VDD.n1070 7.674
R842 VDD.n1152 VDD.n1151 7.674
R843 VDD.n1213 VDD.n1212 7.674
R844 VDD.n1274 VDD.n1273 7.674
R845 VDD.n1335 VDD.n1334 7.674
R846 VDD.n635 VDD.n634 7.674
R847 VDD.n574 VDD.n573 7.674
R848 VDD.n493 VDD.n492 7.674
R849 VDD.n432 VDD.n431 7.674
R850 VDD.n371 VDD.n370 7.674
R851 VDD.n310 VDD.n309 7.674
R852 VDD.n249 VDD.n248 7.674
R853 VDD.n188 VDD.n187 7.674
R854 VDD.n127 VDD.n126 7.674
R855 VDD.n73 VDD.n72 7.674
R856 VDD.n766 VDD.n765 7.674
R857 VDD.n67 VDD.n66 7.5
R858 VDD.n61 VDD.n60 7.5
R859 VDD.n63 VDD.n62 7.5
R860 VDD.n58 VDD.n57 7.5
R861 VDD.n72 VDD.n71 7.5
R862 VDD.n121 VDD.n120 7.5
R863 VDD.n115 VDD.n114 7.5
R864 VDD.n117 VDD.n116 7.5
R865 VDD.n123 VDD.n113 7.5
R866 VDD.n123 VDD.n111 7.5
R867 VDD.n126 VDD.n125 7.5
R868 VDD.n182 VDD.n181 7.5
R869 VDD.n176 VDD.n175 7.5
R870 VDD.n178 VDD.n177 7.5
R871 VDD.n184 VDD.n174 7.5
R872 VDD.n184 VDD.n172 7.5
R873 VDD.n187 VDD.n186 7.5
R874 VDD.n243 VDD.n242 7.5
R875 VDD.n237 VDD.n236 7.5
R876 VDD.n239 VDD.n238 7.5
R877 VDD.n245 VDD.n235 7.5
R878 VDD.n245 VDD.n233 7.5
R879 VDD.n248 VDD.n247 7.5
R880 VDD.n304 VDD.n303 7.5
R881 VDD.n298 VDD.n297 7.5
R882 VDD.n300 VDD.n299 7.5
R883 VDD.n306 VDD.n296 7.5
R884 VDD.n306 VDD.n294 7.5
R885 VDD.n309 VDD.n308 7.5
R886 VDD.n365 VDD.n364 7.5
R887 VDD.n359 VDD.n358 7.5
R888 VDD.n361 VDD.n360 7.5
R889 VDD.n367 VDD.n357 7.5
R890 VDD.n367 VDD.n355 7.5
R891 VDD.n370 VDD.n369 7.5
R892 VDD.n426 VDD.n425 7.5
R893 VDD.n420 VDD.n419 7.5
R894 VDD.n422 VDD.n421 7.5
R895 VDD.n428 VDD.n418 7.5
R896 VDD.n428 VDD.n416 7.5
R897 VDD.n431 VDD.n430 7.5
R898 VDD.n487 VDD.n486 7.5
R899 VDD.n481 VDD.n480 7.5
R900 VDD.n483 VDD.n482 7.5
R901 VDD.n489 VDD.n479 7.5
R902 VDD.n489 VDD.n477 7.5
R903 VDD.n492 VDD.n491 7.5
R904 VDD.n568 VDD.n567 7.5
R905 VDD.n562 VDD.n561 7.5
R906 VDD.n564 VDD.n563 7.5
R907 VDD.n570 VDD.n560 7.5
R908 VDD.n570 VDD.n558 7.5
R909 VDD.n573 VDD.n572 7.5
R910 VDD.n629 VDD.n628 7.5
R911 VDD.n623 VDD.n622 7.5
R912 VDD.n625 VDD.n624 7.5
R913 VDD.n631 VDD.n621 7.5
R914 VDD.n631 VDD.n619 7.5
R915 VDD.n634 VDD.n633 7.5
R916 VDD.n1329 VDD.n1328 7.5
R917 VDD.n1323 VDD.n1322 7.5
R918 VDD.n1325 VDD.n1324 7.5
R919 VDD.n1331 VDD.n1321 7.5
R920 VDD.n1331 VDD.n1319 7.5
R921 VDD.n1334 VDD.n1333 7.5
R922 VDD.n1268 VDD.n1267 7.5
R923 VDD.n1262 VDD.n1261 7.5
R924 VDD.n1264 VDD.n1263 7.5
R925 VDD.n1270 VDD.n1260 7.5
R926 VDD.n1270 VDD.n1258 7.5
R927 VDD.n1273 VDD.n1272 7.5
R928 VDD.n1207 VDD.n1206 7.5
R929 VDD.n1201 VDD.n1200 7.5
R930 VDD.n1203 VDD.n1202 7.5
R931 VDD.n1209 VDD.n1199 7.5
R932 VDD.n1209 VDD.n1197 7.5
R933 VDD.n1212 VDD.n1211 7.5
R934 VDD.n1146 VDD.n1145 7.5
R935 VDD.n1140 VDD.n1139 7.5
R936 VDD.n1142 VDD.n1141 7.5
R937 VDD.n1148 VDD.n1138 7.5
R938 VDD.n1148 VDD.n1136 7.5
R939 VDD.n1151 VDD.n1150 7.5
R940 VDD.n1065 VDD.n1064 7.5
R941 VDD.n1059 VDD.n1058 7.5
R942 VDD.n1061 VDD.n1060 7.5
R943 VDD.n1067 VDD.n1057 7.5
R944 VDD.n1067 VDD.n1055 7.5
R945 VDD.n1070 VDD.n1069 7.5
R946 VDD.n1004 VDD.n1003 7.5
R947 VDD.n998 VDD.n997 7.5
R948 VDD.n1000 VDD.n999 7.5
R949 VDD.n1006 VDD.n996 7.5
R950 VDD.n1006 VDD.n994 7.5
R951 VDD.n1009 VDD.n1008 7.5
R952 VDD.n943 VDD.n942 7.5
R953 VDD.n937 VDD.n936 7.5
R954 VDD.n939 VDD.n938 7.5
R955 VDD.n945 VDD.n935 7.5
R956 VDD.n945 VDD.n933 7.5
R957 VDD.n948 VDD.n947 7.5
R958 VDD.n882 VDD.n881 7.5
R959 VDD.n876 VDD.n875 7.5
R960 VDD.n878 VDD.n877 7.5
R961 VDD.n884 VDD.n874 7.5
R962 VDD.n884 VDD.n872 7.5
R963 VDD.n887 VDD.n886 7.5
R964 VDD.n821 VDD.n820 7.5
R965 VDD.n815 VDD.n814 7.5
R966 VDD.n817 VDD.n816 7.5
R967 VDD.n823 VDD.n813 7.5
R968 VDD.n823 VDD.n811 7.5
R969 VDD.n826 VDD.n825 7.5
R970 VDD.n750 VDD.n749 7.5
R971 VDD.n753 VDD.n752 7.5
R972 VDD.n755 VDD.n754 7.5
R973 VDD.n758 VDD.n757 7.5
R974 VDD.n765 VDD.n764 7.5
R975 VDD.n680 VDD.n679 7.5
R976 VDD.n674 VDD.n673 7.5
R977 VDD.n676 VDD.n675 7.5
R978 VDD.n682 VDD.n672 7.5
R979 VDD.n682 VDD.n670 7.5
R980 VDD.n685 VDD.n684 7.5
R981 VDD.n20 VDD.n16 7.5
R982 VDD.n2 VDD.n1 7.5
R983 VDD.n6 VDD.n5 7.5
R984 VDD.n9 VDD.n8 7.5
R985 VDD.n19 VDD.n18 7.5
R986 VDD.n14 VDD.n0 7.5
R987 VDD.n59 VDD.n56 6.772
R988 VDD.n70 VDD.n54 6.772
R989 VDD.n68 VDD.n65 6.772
R990 VDD.n64 VDD.n61 6.772
R991 VDD.n124 VDD.n109 6.772
R992 VDD.n122 VDD.n119 6.772
R993 VDD.n118 VDD.n115 6.772
R994 VDD.n185 VDD.n170 6.772
R995 VDD.n183 VDD.n180 6.772
R996 VDD.n179 VDD.n176 6.772
R997 VDD.n246 VDD.n231 6.772
R998 VDD.n244 VDD.n241 6.772
R999 VDD.n240 VDD.n237 6.772
R1000 VDD.n307 VDD.n292 6.772
R1001 VDD.n305 VDD.n302 6.772
R1002 VDD.n301 VDD.n298 6.772
R1003 VDD.n368 VDD.n353 6.772
R1004 VDD.n366 VDD.n363 6.772
R1005 VDD.n362 VDD.n359 6.772
R1006 VDD.n429 VDD.n414 6.772
R1007 VDD.n427 VDD.n424 6.772
R1008 VDD.n423 VDD.n420 6.772
R1009 VDD.n490 VDD.n475 6.772
R1010 VDD.n488 VDD.n485 6.772
R1011 VDD.n484 VDD.n481 6.772
R1012 VDD.n571 VDD.n556 6.772
R1013 VDD.n569 VDD.n566 6.772
R1014 VDD.n565 VDD.n562 6.772
R1015 VDD.n632 VDD.n617 6.772
R1016 VDD.n630 VDD.n627 6.772
R1017 VDD.n626 VDD.n623 6.772
R1018 VDD.n1332 VDD.n1317 6.772
R1019 VDD.n1330 VDD.n1327 6.772
R1020 VDD.n1326 VDD.n1323 6.772
R1021 VDD.n1271 VDD.n1256 6.772
R1022 VDD.n1269 VDD.n1266 6.772
R1023 VDD.n1265 VDD.n1262 6.772
R1024 VDD.n1210 VDD.n1195 6.772
R1025 VDD.n1208 VDD.n1205 6.772
R1026 VDD.n1204 VDD.n1201 6.772
R1027 VDD.n1149 VDD.n1134 6.772
R1028 VDD.n1147 VDD.n1144 6.772
R1029 VDD.n1143 VDD.n1140 6.772
R1030 VDD.n1068 VDD.n1053 6.772
R1031 VDD.n1066 VDD.n1063 6.772
R1032 VDD.n1062 VDD.n1059 6.772
R1033 VDD.n1007 VDD.n992 6.772
R1034 VDD.n1005 VDD.n1002 6.772
R1035 VDD.n1001 VDD.n998 6.772
R1036 VDD.n946 VDD.n931 6.772
R1037 VDD.n944 VDD.n941 6.772
R1038 VDD.n940 VDD.n937 6.772
R1039 VDD.n885 VDD.n870 6.772
R1040 VDD.n883 VDD.n880 6.772
R1041 VDD.n879 VDD.n876 6.772
R1042 VDD.n824 VDD.n809 6.772
R1043 VDD.n822 VDD.n819 6.772
R1044 VDD.n818 VDD.n815 6.772
R1045 VDD.n683 VDD.n669 6.772
R1046 VDD.n681 VDD.n678 6.772
R1047 VDD.n677 VDD.n674 6.772
R1048 VDD.n59 VDD.n58 6.772
R1049 VDD.n64 VDD.n63 6.772
R1050 VDD.n68 VDD.n67 6.772
R1051 VDD.n71 VDD.n70 6.772
R1052 VDD.n118 VDD.n117 6.772
R1053 VDD.n122 VDD.n121 6.772
R1054 VDD.n125 VDD.n124 6.772
R1055 VDD.n179 VDD.n178 6.772
R1056 VDD.n183 VDD.n182 6.772
R1057 VDD.n186 VDD.n185 6.772
R1058 VDD.n240 VDD.n239 6.772
R1059 VDD.n244 VDD.n243 6.772
R1060 VDD.n247 VDD.n246 6.772
R1061 VDD.n301 VDD.n300 6.772
R1062 VDD.n305 VDD.n304 6.772
R1063 VDD.n308 VDD.n307 6.772
R1064 VDD.n362 VDD.n361 6.772
R1065 VDD.n366 VDD.n365 6.772
R1066 VDD.n369 VDD.n368 6.772
R1067 VDD.n423 VDD.n422 6.772
R1068 VDD.n427 VDD.n426 6.772
R1069 VDD.n430 VDD.n429 6.772
R1070 VDD.n484 VDD.n483 6.772
R1071 VDD.n488 VDD.n487 6.772
R1072 VDD.n491 VDD.n490 6.772
R1073 VDD.n565 VDD.n564 6.772
R1074 VDD.n569 VDD.n568 6.772
R1075 VDD.n572 VDD.n571 6.772
R1076 VDD.n626 VDD.n625 6.772
R1077 VDD.n630 VDD.n629 6.772
R1078 VDD.n633 VDD.n632 6.772
R1079 VDD.n1326 VDD.n1325 6.772
R1080 VDD.n1330 VDD.n1329 6.772
R1081 VDD.n1333 VDD.n1332 6.772
R1082 VDD.n1265 VDD.n1264 6.772
R1083 VDD.n1269 VDD.n1268 6.772
R1084 VDD.n1272 VDD.n1271 6.772
R1085 VDD.n1204 VDD.n1203 6.772
R1086 VDD.n1208 VDD.n1207 6.772
R1087 VDD.n1211 VDD.n1210 6.772
R1088 VDD.n1143 VDD.n1142 6.772
R1089 VDD.n1147 VDD.n1146 6.772
R1090 VDD.n1150 VDD.n1149 6.772
R1091 VDD.n1062 VDD.n1061 6.772
R1092 VDD.n1066 VDD.n1065 6.772
R1093 VDD.n1069 VDD.n1068 6.772
R1094 VDD.n1001 VDD.n1000 6.772
R1095 VDD.n1005 VDD.n1004 6.772
R1096 VDD.n1008 VDD.n1007 6.772
R1097 VDD.n940 VDD.n939 6.772
R1098 VDD.n944 VDD.n943 6.772
R1099 VDD.n947 VDD.n946 6.772
R1100 VDD.n879 VDD.n878 6.772
R1101 VDD.n883 VDD.n882 6.772
R1102 VDD.n886 VDD.n885 6.772
R1103 VDD.n818 VDD.n817 6.772
R1104 VDD.n822 VDD.n821 6.772
R1105 VDD.n825 VDD.n824 6.772
R1106 VDD.n677 VDD.n676 6.772
R1107 VDD.n681 VDD.n680 6.772
R1108 VDD.n684 VDD.n683 6.772
R1109 VDD.n764 VDD.n763 6.772
R1110 VDD.n751 VDD.n748 6.772
R1111 VDD.n756 VDD.n753 6.772
R1112 VDD.n761 VDD.n758 6.772
R1113 VDD.n761 VDD.n760 6.772
R1114 VDD.n756 VDD.n755 6.772
R1115 VDD.n751 VDD.n750 6.772
R1116 VDD.n763 VDD.n747 6.772
R1117 VDD.n534 VDD.n530 6.69
R1118 VDD.n1096 VDD.n1092 6.69
R1119 VDD.n709 VDD.n705 6.69
R1120 VDD.n33 VDD.n23 6.487
R1121 VDD.n33 VDD.n32 6.475
R1122 VDD.n16 VDD.n15 6.458
R1123 VDD.n517 VDD.n516 6.296
R1124 VDD.n1113 VDD.n1112 6.296
R1125 VDD.n726 VDD.n725 6.296
R1126 VDD.n113 VDD.n112 6.202
R1127 VDD.n174 VDD.n173 6.202
R1128 VDD.n235 VDD.n234 6.202
R1129 VDD.n296 VDD.n295 6.202
R1130 VDD.n357 VDD.n356 6.202
R1131 VDD.n418 VDD.n417 6.202
R1132 VDD.n479 VDD.n478 6.202
R1133 VDD.n560 VDD.n559 6.202
R1134 VDD.n621 VDD.n620 6.202
R1135 VDD.n1321 VDD.n1320 6.202
R1136 VDD.n1260 VDD.n1259 6.202
R1137 VDD.n1199 VDD.n1198 6.202
R1138 VDD.n1138 VDD.n1137 6.202
R1139 VDD.n1057 VDD.n1056 6.202
R1140 VDD.n996 VDD.n995 6.202
R1141 VDD.n935 VDD.n934 6.202
R1142 VDD.n874 VDD.n873 6.202
R1143 VDD.n813 VDD.n812 6.202
R1144 VDD.n672 VDD.n671 6.202
R1145 VDD.n150 VDD.n149 4.576
R1146 VDD.n211 VDD.n210 4.576
R1147 VDD.n272 VDD.n271 4.576
R1148 VDD.n333 VDD.n332 4.576
R1149 VDD.n394 VDD.n393 4.576
R1150 VDD.n455 VDD.n454 4.576
R1151 VDD.n597 VDD.n596 4.576
R1152 VDD.n658 VDD.n657 4.576
R1153 VDD.n1291 VDD.n1290 4.576
R1154 VDD.n1230 VDD.n1229 4.576
R1155 VDD.n1169 VDD.n1168 4.576
R1156 VDD.n1027 VDD.n1026 4.576
R1157 VDD.n966 VDD.n965 4.576
R1158 VDD.n905 VDD.n904 4.576
R1159 VDD.n844 VDD.n843 4.576
R1160 VDD.n783 VDD.n782 4.576
R1161 VDD.n162 VDD.n159 2.754
R1162 VDD.n223 VDD.n220 2.754
R1163 VDD.n284 VDD.n281 2.754
R1164 VDD.n345 VDD.n342 2.754
R1165 VDD.n406 VDD.n403 2.754
R1166 VDD.n467 VDD.n464 2.754
R1167 VDD.n609 VDD.n606 2.754
R1168 VDD.n1344 VDD.n1341 2.754
R1169 VDD.n1283 VDD.n1280 2.754
R1170 VDD.n1222 VDD.n1219 2.754
R1171 VDD.n1161 VDD.n1158 2.754
R1172 VDD.n1019 VDD.n1016 2.754
R1173 VDD.n958 VDD.n955 2.754
R1174 VDD.n897 VDD.n894 2.754
R1175 VDD.n836 VDD.n833 2.754
R1176 VDD.n775 VDD.n772 2.754
R1177 VDD.n136 VDD.n133 2.361
R1178 VDD.n197 VDD.n194 2.361
R1179 VDD.n258 VDD.n255 2.361
R1180 VDD.n319 VDD.n316 2.361
R1181 VDD.n380 VDD.n377 2.361
R1182 VDD.n441 VDD.n438 2.361
R1183 VDD.n583 VDD.n580 2.361
R1184 VDD.n644 VDD.n641 2.361
R1185 VDD.n1309 VDD.n1306 2.361
R1186 VDD.n1248 VDD.n1245 2.361
R1187 VDD.n1187 VDD.n1184 2.361
R1188 VDD.n1045 VDD.n1042 2.361
R1189 VDD.n984 VDD.n981 2.361
R1190 VDD.n923 VDD.n920 2.361
R1191 VDD.n862 VDD.n859 2.361
R1192 VDD.n801 VDD.n798 2.361
R1193 VDD.n14 VDD.n7 1.329
R1194 VDD.n14 VDD.n10 1.329
R1195 VDD.n14 VDD.n11 1.329
R1196 VDD.n14 VDD.n13 1.329
R1197 VDD.n15 VDD.n14 0.696
R1198 VDD.n14 VDD.n4 0.696
R1199 VDD.n544 VDD.n541 0.393
R1200 VDD.n1084 VDD.n1081 0.393
R1201 VDD.n697 VDD.n694 0.393
R1202 VDD.n69 VDD.n68 0.365
R1203 VDD.n69 VDD.n64 0.365
R1204 VDD.n69 VDD.n59 0.365
R1205 VDD.n70 VDD.n69 0.365
R1206 VDD.n123 VDD.n122 0.365
R1207 VDD.n123 VDD.n118 0.365
R1208 VDD.n124 VDD.n123 0.365
R1209 VDD.n184 VDD.n183 0.365
R1210 VDD.n184 VDD.n179 0.365
R1211 VDD.n185 VDD.n184 0.365
R1212 VDD.n245 VDD.n244 0.365
R1213 VDD.n245 VDD.n240 0.365
R1214 VDD.n246 VDD.n245 0.365
R1215 VDD.n306 VDD.n305 0.365
R1216 VDD.n306 VDD.n301 0.365
R1217 VDD.n307 VDD.n306 0.365
R1218 VDD.n367 VDD.n366 0.365
R1219 VDD.n367 VDD.n362 0.365
R1220 VDD.n368 VDD.n367 0.365
R1221 VDD.n428 VDD.n427 0.365
R1222 VDD.n428 VDD.n423 0.365
R1223 VDD.n429 VDD.n428 0.365
R1224 VDD.n489 VDD.n488 0.365
R1225 VDD.n489 VDD.n484 0.365
R1226 VDD.n490 VDD.n489 0.365
R1227 VDD.n570 VDD.n569 0.365
R1228 VDD.n570 VDD.n565 0.365
R1229 VDD.n571 VDD.n570 0.365
R1230 VDD.n631 VDD.n630 0.365
R1231 VDD.n631 VDD.n626 0.365
R1232 VDD.n632 VDD.n631 0.365
R1233 VDD.n1331 VDD.n1330 0.365
R1234 VDD.n1331 VDD.n1326 0.365
R1235 VDD.n1332 VDD.n1331 0.365
R1236 VDD.n1270 VDD.n1269 0.365
R1237 VDD.n1270 VDD.n1265 0.365
R1238 VDD.n1271 VDD.n1270 0.365
R1239 VDD.n1209 VDD.n1208 0.365
R1240 VDD.n1209 VDD.n1204 0.365
R1241 VDD.n1210 VDD.n1209 0.365
R1242 VDD.n1148 VDD.n1147 0.365
R1243 VDD.n1148 VDD.n1143 0.365
R1244 VDD.n1149 VDD.n1148 0.365
R1245 VDD.n1067 VDD.n1066 0.365
R1246 VDD.n1067 VDD.n1062 0.365
R1247 VDD.n1068 VDD.n1067 0.365
R1248 VDD.n1006 VDD.n1005 0.365
R1249 VDD.n1006 VDD.n1001 0.365
R1250 VDD.n1007 VDD.n1006 0.365
R1251 VDD.n945 VDD.n944 0.365
R1252 VDD.n945 VDD.n940 0.365
R1253 VDD.n946 VDD.n945 0.365
R1254 VDD.n884 VDD.n883 0.365
R1255 VDD.n884 VDD.n879 0.365
R1256 VDD.n885 VDD.n884 0.365
R1257 VDD.n823 VDD.n822 0.365
R1258 VDD.n823 VDD.n818 0.365
R1259 VDD.n824 VDD.n823 0.365
R1260 VDD.n682 VDD.n681 0.365
R1261 VDD.n682 VDD.n677 0.365
R1262 VDD.n683 VDD.n682 0.365
R1263 VDD.n762 VDD.n761 0.365
R1264 VDD.n762 VDD.n756 0.365
R1265 VDD.n762 VDD.n751 0.365
R1266 VDD.n763 VDD.n762 0.365
R1267 VDD.n78 VDD.n51 0.29
R1268 VDD.n132 VDD.n106 0.29
R1269 VDD.n193 VDD.n167 0.29
R1270 VDD.n254 VDD.n228 0.29
R1271 VDD.n315 VDD.n289 0.29
R1272 VDD.n376 VDD.n350 0.29
R1273 VDD.n437 VDD.n411 0.29
R1274 VDD.n498 VDD.n472 0.29
R1275 VDD.n579 VDD.n553 0.29
R1276 VDD.n640 VDD.n614 0.29
R1277 VDD.n1340 VDD.n1314 0.29
R1278 VDD.n1279 VDD.n1253 0.29
R1279 VDD.n1218 VDD.n1192 0.29
R1280 VDD.n1157 VDD.n1131 0.29
R1281 VDD.n1076 VDD.n1050 0.29
R1282 VDD.n1015 VDD.n989 0.29
R1283 VDD.n954 VDD.n928 0.29
R1284 VDD.n893 VDD.n867 0.29
R1285 VDD.n832 VDD.n806 0.29
R1286 VDD.n771 VDD.n744 0.29
R1287 VDD.n689 VDD 0.207
R1288 VDD.n528 VDD.n523 0.197
R1289 VDD.n1107 VDD.n1102 0.197
R1290 VDD.n720 VDD.n715 0.197
R1291 VDD.n39 VDD.n35 0.181
R1292 VDD.n94 VDD.n90 0.181
R1293 VDD.n153 VDD.n148 0.181
R1294 VDD.n214 VDD.n209 0.181
R1295 VDD.n275 VDD.n270 0.181
R1296 VDD.n336 VDD.n331 0.181
R1297 VDD.n397 VDD.n392 0.181
R1298 VDD.n458 VDD.n453 0.181
R1299 VDD.n600 VDD.n595 0.181
R1300 VDD.n661 VDD.n656 0.181
R1301 VDD.n1300 VDD.n1294 0.181
R1302 VDD.n1239 VDD.n1233 0.181
R1303 VDD.n1178 VDD.n1172 0.181
R1304 VDD.n1036 VDD.n1030 0.181
R1305 VDD.n975 VDD.n969 0.181
R1306 VDD.n914 VDD.n908 0.181
R1307 VDD.n853 VDD.n847 0.181
R1308 VDD.n792 VDD.n786 0.181
R1309 VDD.n35 VDD.n34 0.145
R1310 VDD.n43 VDD.n39 0.145
R1311 VDD.n47 VDD.n43 0.145
R1312 VDD.n51 VDD.n47 0.145
R1313 VDD.n82 VDD.n78 0.145
R1314 VDD.n86 VDD.n82 0.145
R1315 VDD.n90 VDD.n86 0.145
R1316 VDD.n98 VDD.n94 0.145
R1317 VDD.n102 VDD.n98 0.145
R1318 VDD.n106 VDD.n102 0.145
R1319 VDD.n137 VDD.n132 0.145
R1320 VDD.n142 VDD.n137 0.145
R1321 VDD.n148 VDD.n142 0.145
R1322 VDD.n158 VDD.n153 0.145
R1323 VDD.n163 VDD.n158 0.145
R1324 VDD.n167 VDD.n163 0.145
R1325 VDD.n198 VDD.n193 0.145
R1326 VDD.n203 VDD.n198 0.145
R1327 VDD.n209 VDD.n203 0.145
R1328 VDD.n219 VDD.n214 0.145
R1329 VDD.n224 VDD.n219 0.145
R1330 VDD.n228 VDD.n224 0.145
R1331 VDD.n259 VDD.n254 0.145
R1332 VDD.n264 VDD.n259 0.145
R1333 VDD.n270 VDD.n264 0.145
R1334 VDD.n280 VDD.n275 0.145
R1335 VDD.n285 VDD.n280 0.145
R1336 VDD.n289 VDD.n285 0.145
R1337 VDD.n320 VDD.n315 0.145
R1338 VDD.n325 VDD.n320 0.145
R1339 VDD.n331 VDD.n325 0.145
R1340 VDD.n341 VDD.n336 0.145
R1341 VDD.n346 VDD.n341 0.145
R1342 VDD.n350 VDD.n346 0.145
R1343 VDD.n381 VDD.n376 0.145
R1344 VDD.n386 VDD.n381 0.145
R1345 VDD.n392 VDD.n386 0.145
R1346 VDD.n402 VDD.n397 0.145
R1347 VDD.n407 VDD.n402 0.145
R1348 VDD.n411 VDD.n407 0.145
R1349 VDD.n442 VDD.n437 0.145
R1350 VDD.n447 VDD.n442 0.145
R1351 VDD.n453 VDD.n447 0.145
R1352 VDD.n463 VDD.n458 0.145
R1353 VDD.n468 VDD.n463 0.145
R1354 VDD.n472 VDD.n468 0.145
R1355 VDD.n502 VDD.n498 0.145
R1356 VDD.n506 VDD.n502 0.145
R1357 VDD.n511 VDD.n506 0.145
R1358 VDD.n518 VDD.n511 0.145
R1359 VDD.n523 VDD.n518 0.145
R1360 VDD.n535 VDD.n528 0.145
R1361 VDD.n540 VDD.n535 0.145
R1362 VDD.n545 VDD.n540 0.145
R1363 VDD.n549 VDD.n545 0.145
R1364 VDD.n553 VDD.n549 0.145
R1365 VDD.n584 VDD.n579 0.145
R1366 VDD.n589 VDD.n584 0.145
R1367 VDD.n595 VDD.n589 0.145
R1368 VDD.n605 VDD.n600 0.145
R1369 VDD.n610 VDD.n605 0.145
R1370 VDD.n614 VDD.n610 0.145
R1371 VDD.n645 VDD.n640 0.145
R1372 VDD.n650 VDD.n645 0.145
R1373 VDD.n656 VDD.n650 0.145
R1374 VDD.n666 VDD.n661 0.145
R1375 VDD.n1345 VDD.n1340 0.145
R1376 VDD.n1314 VDD.n1310 0.145
R1377 VDD.n1310 VDD.n1305 0.145
R1378 VDD.n1305 VDD.n1300 0.145
R1379 VDD.n1294 VDD.n1289 0.145
R1380 VDD.n1289 VDD.n1284 0.145
R1381 VDD.n1284 VDD.n1279 0.145
R1382 VDD.n1253 VDD.n1249 0.145
R1383 VDD.n1249 VDD.n1244 0.145
R1384 VDD.n1244 VDD.n1239 0.145
R1385 VDD.n1233 VDD.n1228 0.145
R1386 VDD.n1228 VDD.n1223 0.145
R1387 VDD.n1223 VDD.n1218 0.145
R1388 VDD.n1192 VDD.n1188 0.145
R1389 VDD.n1188 VDD.n1183 0.145
R1390 VDD.n1183 VDD.n1178 0.145
R1391 VDD.n1172 VDD.n1167 0.145
R1392 VDD.n1167 VDD.n1162 0.145
R1393 VDD.n1162 VDD.n1157 0.145
R1394 VDD.n1131 VDD.n1127 0.145
R1395 VDD.n1127 VDD.n1123 0.145
R1396 VDD.n1123 VDD.n1119 0.145
R1397 VDD.n1119 VDD.n1114 0.145
R1398 VDD.n1114 VDD.n1107 0.145
R1399 VDD.n1102 VDD.n1097 0.145
R1400 VDD.n1097 VDD.n1090 0.145
R1401 VDD.n1090 VDD.n1085 0.145
R1402 VDD.n1085 VDD.n1080 0.145
R1403 VDD.n1080 VDD.n1076 0.145
R1404 VDD.n1050 VDD.n1046 0.145
R1405 VDD.n1046 VDD.n1041 0.145
R1406 VDD.n1041 VDD.n1036 0.145
R1407 VDD.n1030 VDD.n1025 0.145
R1408 VDD.n1025 VDD.n1020 0.145
R1409 VDD.n1020 VDD.n1015 0.145
R1410 VDD.n989 VDD.n985 0.145
R1411 VDD.n985 VDD.n980 0.145
R1412 VDD.n980 VDD.n975 0.145
R1413 VDD.n969 VDD.n964 0.145
R1414 VDD.n964 VDD.n959 0.145
R1415 VDD.n959 VDD.n954 0.145
R1416 VDD.n928 VDD.n924 0.145
R1417 VDD.n924 VDD.n919 0.145
R1418 VDD.n919 VDD.n914 0.145
R1419 VDD.n908 VDD.n903 0.145
R1420 VDD.n903 VDD.n898 0.145
R1421 VDD.n898 VDD.n893 0.145
R1422 VDD.n867 VDD.n863 0.145
R1423 VDD.n863 VDD.n858 0.145
R1424 VDD.n858 VDD.n853 0.145
R1425 VDD.n847 VDD.n842 0.145
R1426 VDD.n842 VDD.n837 0.145
R1427 VDD.n837 VDD.n832 0.145
R1428 VDD.n806 VDD.n802 0.145
R1429 VDD.n802 VDD.n797 0.145
R1430 VDD.n797 VDD.n792 0.145
R1431 VDD.n786 VDD.n781 0.145
R1432 VDD.n781 VDD.n776 0.145
R1433 VDD.n776 VDD.n771 0.145
R1434 VDD.n744 VDD.n740 0.145
R1435 VDD.n740 VDD.n736 0.145
R1436 VDD.n736 VDD.n732 0.145
R1437 VDD.n732 VDD.n727 0.145
R1438 VDD.n727 VDD.n720 0.145
R1439 VDD.n715 VDD.n710 0.145
R1440 VDD.n710 VDD.n703 0.145
R1441 VDD.n703 VDD.n698 0.145
R1442 VDD.n698 VDD.n693 0.145
R1443 VDD.n693 VDD.n689 0.145
R1444 VDD VDD.n1345 0.082
R1445 VDD VDD.n666 0.062
R1446 a_599_989.n0 a_599_989.t9 480.392
R1447 a_599_989.n2 a_599_989.t10 454.685
R1448 a_599_989.n2 a_599_989.t7 428.979
R1449 a_599_989.n0 a_599_989.t5 403.272
R1450 a_599_989.n1 a_599_989.t8 283.48
R1451 a_599_989.n3 a_599_989.t6 237.959
R1452 a_599_989.n9 a_599_989.n8 210.592
R1453 a_599_989.n11 a_599_989.n9 152.499
R1454 a_599_989.n3 a_599_989.n2 98.447
R1455 a_599_989.n1 a_599_989.n0 98.447
R1456 a_599_989.n4 a_599_989.n3 78.947
R1457 a_599_989.n4 a_599_989.n1 77.315
R1458 a_599_989.n11 a_599_989.n10 76.002
R1459 a_599_989.n9 a_599_989.n4 76
R1460 a_599_989.n8 a_599_989.n7 30
R1461 a_599_989.n6 a_599_989.n5 24.383
R1462 a_599_989.n8 a_599_989.n6 23.684
R1463 a_599_989.n10 a_599_989.t0 14.282
R1464 a_599_989.n10 a_599_989.t1 14.282
R1465 a_599_989.n12 a_599_989.t3 14.282
R1466 a_599_989.t4 a_599_989.n12 14.282
R1467 a_599_989.n12 a_599_989.n11 12.848
R1468 a_3303_411.n4 a_3303_411.t8 512.525
R1469 a_3303_411.n3 a_3303_411.t10 512.525
R1470 a_3303_411.n8 a_3303_411.t12 472.359
R1471 a_3303_411.n8 a_3303_411.t7 384.527
R1472 a_3303_411.n4 a_3303_411.t11 371.139
R1473 a_3303_411.n3 a_3303_411.t9 371.139
R1474 a_3303_411.n5 a_3303_411.n4 265.439
R1475 a_3303_411.n9 a_3303_411.t6 214.619
R1476 a_3303_411.n13 a_3303_411.n11 190.561
R1477 a_3303_411.n7 a_3303_411.n3 185.78
R1478 a_3303_411.n11 a_3303_411.n2 179.052
R1479 a_3303_411.n5 a_3303_411.t5 176.995
R1480 a_3303_411.n6 a_3303_411.t13 170.569
R1481 a_3303_411.n6 a_3303_411.n5 153.043
R1482 a_3303_411.n9 a_3303_411.n8 136.613
R1483 a_3303_411.n10 a_3303_411.n7 112.41
R1484 a_3303_411.n7 a_3303_411.n6 79.658
R1485 a_3303_411.n10 a_3303_411.n9 78.947
R1486 a_3303_411.n2 a_3303_411.n1 76.002
R1487 a_3303_411.n11 a_3303_411.n10 76
R1488 a_3303_411.n13 a_3303_411.n12 15.218
R1489 a_3303_411.n0 a_3303_411.t3 14.282
R1490 a_3303_411.n0 a_3303_411.t0 14.282
R1491 a_3303_411.n1 a_3303_411.t4 14.282
R1492 a_3303_411.n1 a_3303_411.t2 14.282
R1493 a_3303_411.n2 a_3303_411.n0 12.85
R1494 a_3303_411.n14 a_3303_411.n13 12.014
R1495 a_14320_101.t0 a_14320_101.n1 93.333
R1496 a_14320_101.n4 a_14320_101.n2 55.07
R1497 a_14320_101.t0 a_14320_101.n0 8.137
R1498 a_14320_101.n4 a_14320_101.n3 4.619
R1499 a_14320_101.t0 a_14320_101.n4 0.071
R1500 GND.n26 GND.n24 219.745
R1501 GND.n56 GND.n54 219.745
R1502 GND.n380 GND.n379 219.745
R1503 GND.n413 GND.n411 219.745
R1504 GND.n446 GND.n444 219.745
R1505 GND.n476 GND.n474 219.745
R1506 GND.n506 GND.n504 219.745
R1507 GND.n539 GND.n537 219.745
R1508 GND.n581 GND.n579 219.745
R1509 GND.n611 GND.n609 219.745
R1510 GND.n641 GND.n639 219.745
R1511 GND.n671 GND.n669 219.745
R1512 GND.n314 GND.n312 219.745
R1513 GND.n284 GND.n282 219.745
R1514 GND.n242 GND.n240 219.745
R1515 GND.n212 GND.n210 219.745
R1516 GND.n179 GND.n177 219.745
R1517 GND.n149 GND.n147 219.745
R1518 GND.n119 GND.n117 219.745
R1519 GND.n86 GND.n85 219.745
R1520 GND.n273 GND.n272 85.559
R1521 GND.n548 GND.n547 85.559
R1522 GND.n347 GND.n346 85.559
R1523 GND.n26 GND.n25 85.529
R1524 GND.n56 GND.n55 85.529
R1525 GND.n380 GND.n378 85.529
R1526 GND.n413 GND.n412 85.529
R1527 GND.n446 GND.n445 85.529
R1528 GND.n476 GND.n475 85.529
R1529 GND.n506 GND.n505 85.529
R1530 GND.n539 GND.n538 85.529
R1531 GND.n581 GND.n580 85.529
R1532 GND.n611 GND.n610 85.529
R1533 GND.n641 GND.n640 85.529
R1534 GND.n671 GND.n670 85.529
R1535 GND.n314 GND.n313 85.529
R1536 GND.n284 GND.n283 85.529
R1537 GND.n242 GND.n241 85.529
R1538 GND.n212 GND.n211 85.529
R1539 GND.n179 GND.n178 85.529
R1540 GND.n149 GND.n148 85.529
R1541 GND.n119 GND.n118 85.529
R1542 GND.n86 GND.n84 85.529
R1543 GND.n44 GND.n43 84.842
R1544 GND.n74 GND.n73 84.842
R1545 GND.n137 GND.n136 84.842
R1546 GND.n167 GND.n166 84.842
R1547 GND.n230 GND.n229 84.842
R1548 GND.n302 GND.n301 84.842
R1549 GND.n649 GND.n648 84.842
R1550 GND.n619 GND.n618 84.842
R1551 GND.n589 GND.n588 84.842
R1552 GND.n484 GND.n483 84.842
R1553 GND.n454 GND.n453 84.842
R1554 GND.n14 GND.n13 84.842
R1555 GND.n341 GND.n340 76
R1556 GND.n39 GND.n38 76
R1557 GND.n42 GND.n41 76
R1558 GND.n47 GND.n46 76
R1559 GND.n50 GND.n49 76
R1560 GND.n53 GND.n52 76
R1561 GND.n60 GND.n59 76
R1562 GND.n63 GND.n62 76
R1563 GND.n66 GND.n65 76
R1564 GND.n69 GND.n68 76
R1565 GND.n72 GND.n71 76
R1566 GND.n77 GND.n76 76
R1567 GND.n80 GND.n79 76
R1568 GND.n83 GND.n82 76
R1569 GND.n90 GND.n89 76
R1570 GND.n93 GND.n92 76
R1571 GND.n96 GND.n95 76
R1572 GND.n99 GND.n98 76
R1573 GND.n102 GND.n101 76
R1574 GND.n110 GND.n109 76
R1575 GND.n113 GND.n112 76
R1576 GND.n116 GND.n115 76
R1577 GND.n123 GND.n122 76
R1578 GND.n126 GND.n125 76
R1579 GND.n129 GND.n128 76
R1580 GND.n132 GND.n131 76
R1581 GND.n135 GND.n134 76
R1582 GND.n140 GND.n139 76
R1583 GND.n143 GND.n142 76
R1584 GND.n146 GND.n145 76
R1585 GND.n153 GND.n152 76
R1586 GND.n156 GND.n155 76
R1587 GND.n159 GND.n158 76
R1588 GND.n162 GND.n161 76
R1589 GND.n165 GND.n164 76
R1590 GND.n170 GND.n169 76
R1591 GND.n173 GND.n172 76
R1592 GND.n176 GND.n175 76
R1593 GND.n183 GND.n182 76
R1594 GND.n186 GND.n185 76
R1595 GND.n189 GND.n188 76
R1596 GND.n192 GND.n191 76
R1597 GND.n195 GND.n194 76
R1598 GND.n203 GND.n202 76
R1599 GND.n206 GND.n205 76
R1600 GND.n209 GND.n208 76
R1601 GND.n216 GND.n215 76
R1602 GND.n219 GND.n218 76
R1603 GND.n222 GND.n221 76
R1604 GND.n225 GND.n224 76
R1605 GND.n228 GND.n227 76
R1606 GND.n233 GND.n232 76
R1607 GND.n236 GND.n235 76
R1608 GND.n239 GND.n238 76
R1609 GND.n246 GND.n245 76
R1610 GND.n249 GND.n248 76
R1611 GND.n252 GND.n251 76
R1612 GND.n255 GND.n254 76
R1613 GND.n258 GND.n257 76
R1614 GND.n261 GND.n260 76
R1615 GND.n264 GND.n263 76
R1616 GND.n267 GND.n266 76
R1617 GND.n270 GND.n269 76
R1618 GND.n275 GND.n274 76
R1619 GND.n278 GND.n277 76
R1620 GND.n281 GND.n280 76
R1621 GND.n288 GND.n287 76
R1622 GND.n291 GND.n290 76
R1623 GND.n294 GND.n293 76
R1624 GND.n297 GND.n296 76
R1625 GND.n300 GND.n299 76
R1626 GND.n305 GND.n304 76
R1627 GND.n308 GND.n307 76
R1628 GND.n311 GND.n310 76
R1629 GND.n318 GND.n317 76
R1630 GND.n321 GND.n320 76
R1631 GND.n324 GND.n323 76
R1632 GND.n327 GND.n326 76
R1633 GND.n330 GND.n329 76
R1634 GND.n338 GND.n337 76
R1635 GND.n677 GND.n676 76
R1636 GND.n674 GND.n673 76
R1637 GND.n667 GND.n666 76
R1638 GND.n664 GND.n663 76
R1639 GND.n661 GND.n660 76
R1640 GND.n658 GND.n657 76
R1641 GND.n655 GND.n654 76
R1642 GND.n652 GND.n651 76
R1643 GND.n647 GND.n646 76
R1644 GND.n644 GND.n643 76
R1645 GND.n637 GND.n636 76
R1646 GND.n634 GND.n633 76
R1647 GND.n631 GND.n630 76
R1648 GND.n628 GND.n627 76
R1649 GND.n625 GND.n624 76
R1650 GND.n622 GND.n621 76
R1651 GND.n617 GND.n616 76
R1652 GND.n614 GND.n613 76
R1653 GND.n607 GND.n606 76
R1654 GND.n604 GND.n603 76
R1655 GND.n601 GND.n600 76
R1656 GND.n598 GND.n597 76
R1657 GND.n595 GND.n594 76
R1658 GND.n592 GND.n591 76
R1659 GND.n587 GND.n586 76
R1660 GND.n584 GND.n583 76
R1661 GND.n577 GND.n576 76
R1662 GND.n574 GND.n573 76
R1663 GND.n571 GND.n570 76
R1664 GND.n568 GND.n567 76
R1665 GND.n565 GND.n564 76
R1666 GND.n562 GND.n561 76
R1667 GND.n559 GND.n558 76
R1668 GND.n556 GND.n555 76
R1669 GND.n553 GND.n552 76
R1670 GND.n550 GND.n549 76
R1671 GND.n545 GND.n544 76
R1672 GND.n542 GND.n541 76
R1673 GND.n535 GND.n534 76
R1674 GND.n532 GND.n531 76
R1675 GND.n529 GND.n528 76
R1676 GND.n526 GND.n525 76
R1677 GND.n523 GND.n522 76
R1678 GND.n520 GND.n519 76
R1679 GND.n512 GND.n511 76
R1680 GND.n509 GND.n508 76
R1681 GND.n502 GND.n501 76
R1682 GND.n499 GND.n498 76
R1683 GND.n496 GND.n495 76
R1684 GND.n493 GND.n492 76
R1685 GND.n490 GND.n489 76
R1686 GND.n487 GND.n486 76
R1687 GND.n482 GND.n481 76
R1688 GND.n479 GND.n478 76
R1689 GND.n472 GND.n471 76
R1690 GND.n469 GND.n468 76
R1691 GND.n466 GND.n465 76
R1692 GND.n463 GND.n462 76
R1693 GND.n460 GND.n459 76
R1694 GND.n457 GND.n456 76
R1695 GND.n452 GND.n451 76
R1696 GND.n449 GND.n448 76
R1697 GND.n442 GND.n441 76
R1698 GND.n439 GND.n438 76
R1699 GND.n436 GND.n435 76
R1700 GND.n433 GND.n432 76
R1701 GND.n430 GND.n429 76
R1702 GND.n427 GND.n426 76
R1703 GND.n419 GND.n418 76
R1704 GND.n416 GND.n415 76
R1705 GND.n409 GND.n408 76
R1706 GND.n406 GND.n405 76
R1707 GND.n403 GND.n402 76
R1708 GND.n400 GND.n399 76
R1709 GND.n397 GND.n396 76
R1710 GND.n394 GND.n393 76
R1711 GND.n386 GND.n385 76
R1712 GND.n383 GND.n382 76
R1713 GND.n376 GND.n375 76
R1714 GND.n373 GND.n372 76
R1715 GND.n370 GND.n369 76
R1716 GND.n367 GND.n366 76
R1717 GND.n364 GND.n363 76
R1718 GND.n361 GND.n360 76
R1719 GND.n358 GND.n357 76
R1720 GND.n355 GND.n354 76
R1721 GND.n352 GND.n351 76
R1722 GND.n349 GND.n348 76
R1723 GND.n344 GND.n343 76
R1724 GND.n12 GND.n11 76
R1725 GND.n17 GND.n16 76
R1726 GND.n20 GND.n19 76
R1727 GND.n23 GND.n22 76
R1728 GND.n30 GND.n29 76
R1729 GND.n33 GND.n32 76
R1730 GND.n36 GND.n35 76
R1731 GND.n107 GND.n106 63.835
R1732 GND.n200 GND.n199 63.835
R1733 GND.n335 GND.n334 63.835
R1734 GND.n517 GND.n516 63.835
R1735 GND.n424 GND.n423 63.835
R1736 GND.n391 GND.n390 63.835
R1737 GND.n8 GND.n7 34.942
R1738 GND.n106 GND.n105 28.421
R1739 GND.n199 GND.n198 28.421
R1740 GND.n334 GND.n333 28.421
R1741 GND.n516 GND.n515 28.421
R1742 GND.n423 GND.n422 28.421
R1743 GND.n390 GND.n389 28.421
R1744 GND.n106 GND.n104 25.263
R1745 GND.n199 GND.n197 25.263
R1746 GND.n334 GND.n332 25.263
R1747 GND.n516 GND.n514 25.263
R1748 GND.n423 GND.n421 25.263
R1749 GND.n390 GND.n388 25.263
R1750 GND.n104 GND.n103 24.383
R1751 GND.n197 GND.n196 24.383
R1752 GND.n332 GND.n331 24.383
R1753 GND.n514 GND.n513 24.383
R1754 GND.n421 GND.n420 24.383
R1755 GND.n388 GND.n387 24.383
R1756 GND.n5 GND.n4 14.167
R1757 GND.n4 GND.n2 14.167
R1758 GND.n29 GND.n27 14.167
R1759 GND.n59 GND.n57 14.167
R1760 GND.n89 GND.n87 14.167
R1761 GND.n122 GND.n120 14.167
R1762 GND.n152 GND.n150 14.167
R1763 GND.n182 GND.n180 14.167
R1764 GND.n215 GND.n213 14.167
R1765 GND.n245 GND.n243 14.167
R1766 GND.n287 GND.n285 14.167
R1767 GND.n317 GND.n315 14.167
R1768 GND.n673 GND.n672 14.167
R1769 GND.n643 GND.n642 14.167
R1770 GND.n613 GND.n612 14.167
R1771 GND.n583 GND.n582 14.167
R1772 GND.n541 GND.n540 14.167
R1773 GND.n508 GND.n507 14.167
R1774 GND.n478 GND.n477 14.167
R1775 GND.n448 GND.n447 14.167
R1776 GND.n415 GND.n414 14.167
R1777 GND.n382 GND.n381 14.167
R1778 GND.n343 GND.n342 13.653
R1779 GND.n348 GND.n345 13.653
R1780 GND.n351 GND.n350 13.653
R1781 GND.n354 GND.n353 13.653
R1782 GND.n357 GND.n356 13.653
R1783 GND.n360 GND.n359 13.653
R1784 GND.n363 GND.n362 13.653
R1785 GND.n366 GND.n365 13.653
R1786 GND.n369 GND.n368 13.653
R1787 GND.n372 GND.n371 13.653
R1788 GND.n375 GND.n374 13.653
R1789 GND.n382 GND.n377 13.653
R1790 GND.n385 GND.n384 13.653
R1791 GND.n393 GND.n392 13.653
R1792 GND.n396 GND.n395 13.653
R1793 GND.n399 GND.n398 13.653
R1794 GND.n402 GND.n401 13.653
R1795 GND.n405 GND.n404 13.653
R1796 GND.n408 GND.n407 13.653
R1797 GND.n415 GND.n410 13.653
R1798 GND.n418 GND.n417 13.653
R1799 GND.n426 GND.n425 13.653
R1800 GND.n429 GND.n428 13.653
R1801 GND.n432 GND.n431 13.653
R1802 GND.n435 GND.n434 13.653
R1803 GND.n438 GND.n437 13.653
R1804 GND.n441 GND.n440 13.653
R1805 GND.n448 GND.n443 13.653
R1806 GND.n451 GND.n450 13.653
R1807 GND.n456 GND.n455 13.653
R1808 GND.n459 GND.n458 13.653
R1809 GND.n462 GND.n461 13.653
R1810 GND.n465 GND.n464 13.653
R1811 GND.n468 GND.n467 13.653
R1812 GND.n471 GND.n470 13.653
R1813 GND.n478 GND.n473 13.653
R1814 GND.n481 GND.n480 13.653
R1815 GND.n486 GND.n485 13.653
R1816 GND.n489 GND.n488 13.653
R1817 GND.n492 GND.n491 13.653
R1818 GND.n495 GND.n494 13.653
R1819 GND.n498 GND.n497 13.653
R1820 GND.n501 GND.n500 13.653
R1821 GND.n508 GND.n503 13.653
R1822 GND.n511 GND.n510 13.653
R1823 GND.n519 GND.n518 13.653
R1824 GND.n522 GND.n521 13.653
R1825 GND.n525 GND.n524 13.653
R1826 GND.n528 GND.n527 13.653
R1827 GND.n531 GND.n530 13.653
R1828 GND.n534 GND.n533 13.653
R1829 GND.n541 GND.n536 13.653
R1830 GND.n544 GND.n543 13.653
R1831 GND.n549 GND.n546 13.653
R1832 GND.n552 GND.n551 13.653
R1833 GND.n555 GND.n554 13.653
R1834 GND.n558 GND.n557 13.653
R1835 GND.n561 GND.n560 13.653
R1836 GND.n564 GND.n563 13.653
R1837 GND.n567 GND.n566 13.653
R1838 GND.n570 GND.n569 13.653
R1839 GND.n573 GND.n572 13.653
R1840 GND.n576 GND.n575 13.653
R1841 GND.n583 GND.n578 13.653
R1842 GND.n586 GND.n585 13.653
R1843 GND.n591 GND.n590 13.653
R1844 GND.n594 GND.n593 13.653
R1845 GND.n597 GND.n596 13.653
R1846 GND.n600 GND.n599 13.653
R1847 GND.n603 GND.n602 13.653
R1848 GND.n606 GND.n605 13.653
R1849 GND.n613 GND.n608 13.653
R1850 GND.n616 GND.n615 13.653
R1851 GND.n621 GND.n620 13.653
R1852 GND.n624 GND.n623 13.653
R1853 GND.n627 GND.n626 13.653
R1854 GND.n630 GND.n629 13.653
R1855 GND.n633 GND.n632 13.653
R1856 GND.n636 GND.n635 13.653
R1857 GND.n643 GND.n638 13.653
R1858 GND.n646 GND.n645 13.653
R1859 GND.n651 GND.n650 13.653
R1860 GND.n654 GND.n653 13.653
R1861 GND.n657 GND.n656 13.653
R1862 GND.n660 GND.n659 13.653
R1863 GND.n663 GND.n662 13.653
R1864 GND.n666 GND.n665 13.653
R1865 GND.n673 GND.n668 13.653
R1866 GND.n676 GND.n675 13.653
R1867 GND.n337 GND.n336 13.653
R1868 GND.n329 GND.n328 13.653
R1869 GND.n326 GND.n325 13.653
R1870 GND.n323 GND.n322 13.653
R1871 GND.n320 GND.n319 13.653
R1872 GND.n317 GND.n316 13.653
R1873 GND.n310 GND.n309 13.653
R1874 GND.n307 GND.n306 13.653
R1875 GND.n304 GND.n303 13.653
R1876 GND.n299 GND.n298 13.653
R1877 GND.n296 GND.n295 13.653
R1878 GND.n293 GND.n292 13.653
R1879 GND.n290 GND.n289 13.653
R1880 GND.n287 GND.n286 13.653
R1881 GND.n280 GND.n279 13.653
R1882 GND.n277 GND.n276 13.653
R1883 GND.n274 GND.n271 13.653
R1884 GND.n269 GND.n268 13.653
R1885 GND.n266 GND.n265 13.653
R1886 GND.n263 GND.n262 13.653
R1887 GND.n260 GND.n259 13.653
R1888 GND.n257 GND.n256 13.653
R1889 GND.n254 GND.n253 13.653
R1890 GND.n251 GND.n250 13.653
R1891 GND.n248 GND.n247 13.653
R1892 GND.n245 GND.n244 13.653
R1893 GND.n238 GND.n237 13.653
R1894 GND.n235 GND.n234 13.653
R1895 GND.n232 GND.n231 13.653
R1896 GND.n227 GND.n226 13.653
R1897 GND.n224 GND.n223 13.653
R1898 GND.n221 GND.n220 13.653
R1899 GND.n218 GND.n217 13.653
R1900 GND.n215 GND.n214 13.653
R1901 GND.n208 GND.n207 13.653
R1902 GND.n205 GND.n204 13.653
R1903 GND.n202 GND.n201 13.653
R1904 GND.n194 GND.n193 13.653
R1905 GND.n191 GND.n190 13.653
R1906 GND.n188 GND.n187 13.653
R1907 GND.n185 GND.n184 13.653
R1908 GND.n182 GND.n181 13.653
R1909 GND.n175 GND.n174 13.653
R1910 GND.n172 GND.n171 13.653
R1911 GND.n169 GND.n168 13.653
R1912 GND.n164 GND.n163 13.653
R1913 GND.n161 GND.n160 13.653
R1914 GND.n158 GND.n157 13.653
R1915 GND.n155 GND.n154 13.653
R1916 GND.n152 GND.n151 13.653
R1917 GND.n145 GND.n144 13.653
R1918 GND.n142 GND.n141 13.653
R1919 GND.n139 GND.n138 13.653
R1920 GND.n134 GND.n133 13.653
R1921 GND.n131 GND.n130 13.653
R1922 GND.n128 GND.n127 13.653
R1923 GND.n125 GND.n124 13.653
R1924 GND.n122 GND.n121 13.653
R1925 GND.n115 GND.n114 13.653
R1926 GND.n112 GND.n111 13.653
R1927 GND.n109 GND.n108 13.653
R1928 GND.n101 GND.n100 13.653
R1929 GND.n98 GND.n97 13.653
R1930 GND.n95 GND.n94 13.653
R1931 GND.n92 GND.n91 13.653
R1932 GND.n89 GND.n88 13.653
R1933 GND.n82 GND.n81 13.653
R1934 GND.n79 GND.n78 13.653
R1935 GND.n76 GND.n75 13.653
R1936 GND.n71 GND.n70 13.653
R1937 GND.n68 GND.n67 13.653
R1938 GND.n65 GND.n64 13.653
R1939 GND.n62 GND.n61 13.653
R1940 GND.n59 GND.n58 13.653
R1941 GND.n52 GND.n51 13.653
R1942 GND.n49 GND.n48 13.653
R1943 GND.n46 GND.n45 13.653
R1944 GND.n41 GND.n40 13.653
R1945 GND.n38 GND.n37 13.653
R1946 GND.n5 GND.n0 13.653
R1947 GND.n4 GND.n3 13.653
R1948 GND.n2 GND.n1 13.653
R1949 GND.n11 GND.n10 13.653
R1950 GND.n16 GND.n15 13.653
R1951 GND.n19 GND.n18 13.653
R1952 GND.n22 GND.n21 13.653
R1953 GND.n29 GND.n28 13.653
R1954 GND.n32 GND.n31 13.653
R1955 GND.n35 GND.n34 13.653
R1956 GND.n27 GND.n26 7.312
R1957 GND.n57 GND.n56 7.312
R1958 GND.n381 GND.n380 7.312
R1959 GND.n414 GND.n413 7.312
R1960 GND.n447 GND.n446 7.312
R1961 GND.n477 GND.n476 7.312
R1962 GND.n507 GND.n506 7.312
R1963 GND.n540 GND.n539 7.312
R1964 GND.n582 GND.n581 7.312
R1965 GND.n612 GND.n611 7.312
R1966 GND.n642 GND.n641 7.312
R1967 GND.n672 GND.n671 7.312
R1968 GND.n315 GND.n314 7.312
R1969 GND.n285 GND.n284 7.312
R1970 GND.n243 GND.n242 7.312
R1971 GND.n213 GND.n212 7.312
R1972 GND.n180 GND.n179 7.312
R1973 GND.n150 GND.n149 7.312
R1974 GND.n120 GND.n119 7.312
R1975 GND.n87 GND.n86 7.312
R1976 GND.n7 GND.n6 7.084
R1977 GND.n7 GND.n5 6.475
R1978 GND.n16 GND.n14 3.935
R1979 GND.n46 GND.n44 3.935
R1980 GND.n76 GND.n74 3.935
R1981 GND.n109 GND.n107 3.935
R1982 GND.n139 GND.n137 3.935
R1983 GND.n169 GND.n167 3.935
R1984 GND.n202 GND.n200 3.935
R1985 GND.n232 GND.n230 3.935
R1986 GND.n304 GND.n302 3.935
R1987 GND.n337 GND.n335 3.935
R1988 GND.n651 GND.n649 3.935
R1989 GND.n621 GND.n619 3.935
R1990 GND.n591 GND.n589 3.935
R1991 GND.n519 GND.n517 3.935
R1992 GND.n486 GND.n484 3.935
R1993 GND.n456 GND.n454 3.935
R1994 GND.n426 GND.n424 3.935
R1995 GND.n393 GND.n391 3.935
R1996 GND.n340 GND.n339 0.596
R1997 GND.n30 GND.n23 0.29
R1998 GND.n60 GND.n53 0.29
R1999 GND.n90 GND.n83 0.29
R2000 GND.n123 GND.n116 0.29
R2001 GND.n153 GND.n146 0.29
R2002 GND.n183 GND.n176 0.29
R2003 GND.n216 GND.n209 0.29
R2004 GND.n246 GND.n239 0.29
R2005 GND.n288 GND.n281 0.29
R2006 GND.n318 GND.n311 0.29
R2007 GND.n674 GND.n667 0.29
R2008 GND.n644 GND.n637 0.29
R2009 GND.n614 GND.n607 0.29
R2010 GND.n584 GND.n577 0.29
R2011 GND.n542 GND.n535 0.29
R2012 GND.n509 GND.n502 0.29
R2013 GND.n479 GND.n472 0.29
R2014 GND.n449 GND.n442 0.29
R2015 GND.n416 GND.n409 0.29
R2016 GND.n383 GND.n376 0.29
R2017 GND.n341 GND 0.207
R2018 GND.n264 GND.n261 0.197
R2019 GND.n562 GND.n559 0.197
R2020 GND.n361 GND.n358 0.197
R2021 GND.n274 GND.n273 0.196
R2022 GND.n549 GND.n548 0.196
R2023 GND.n348 GND.n347 0.196
R2024 GND.n12 GND.n9 0.181
R2025 GND.n42 GND.n39 0.181
R2026 GND.n72 GND.n69 0.181
R2027 GND.n102 GND.n99 0.181
R2028 GND.n135 GND.n132 0.181
R2029 GND.n165 GND.n162 0.181
R2030 GND.n195 GND.n192 0.181
R2031 GND.n228 GND.n225 0.181
R2032 GND.n300 GND.n297 0.181
R2033 GND.n330 GND.n327 0.181
R2034 GND.n658 GND.n655 0.181
R2035 GND.n628 GND.n625 0.181
R2036 GND.n598 GND.n595 0.181
R2037 GND.n526 GND.n523 0.181
R2038 GND.n493 GND.n490 0.181
R2039 GND.n463 GND.n460 0.181
R2040 GND.n433 GND.n430 0.181
R2041 GND.n400 GND.n397 0.181
R2042 GND.n9 GND.n8 0.145
R2043 GND.n17 GND.n12 0.145
R2044 GND.n20 GND.n17 0.145
R2045 GND.n23 GND.n20 0.145
R2046 GND.n33 GND.n30 0.145
R2047 GND.n36 GND.n33 0.145
R2048 GND.n39 GND.n36 0.145
R2049 GND.n47 GND.n42 0.145
R2050 GND.n50 GND.n47 0.145
R2051 GND.n53 GND.n50 0.145
R2052 GND.n63 GND.n60 0.145
R2053 GND.n66 GND.n63 0.145
R2054 GND.n69 GND.n66 0.145
R2055 GND.n77 GND.n72 0.145
R2056 GND.n80 GND.n77 0.145
R2057 GND.n83 GND.n80 0.145
R2058 GND.n93 GND.n90 0.145
R2059 GND.n96 GND.n93 0.145
R2060 GND.n99 GND.n96 0.145
R2061 GND.n110 GND.n102 0.145
R2062 GND.n113 GND.n110 0.145
R2063 GND.n116 GND.n113 0.145
R2064 GND.n126 GND.n123 0.145
R2065 GND.n129 GND.n126 0.145
R2066 GND.n132 GND.n129 0.145
R2067 GND.n140 GND.n135 0.145
R2068 GND.n143 GND.n140 0.145
R2069 GND.n146 GND.n143 0.145
R2070 GND.n156 GND.n153 0.145
R2071 GND.n159 GND.n156 0.145
R2072 GND.n162 GND.n159 0.145
R2073 GND.n170 GND.n165 0.145
R2074 GND.n173 GND.n170 0.145
R2075 GND.n176 GND.n173 0.145
R2076 GND.n186 GND.n183 0.145
R2077 GND.n189 GND.n186 0.145
R2078 GND.n192 GND.n189 0.145
R2079 GND.n203 GND.n195 0.145
R2080 GND.n206 GND.n203 0.145
R2081 GND.n209 GND.n206 0.145
R2082 GND.n219 GND.n216 0.145
R2083 GND.n222 GND.n219 0.145
R2084 GND.n225 GND.n222 0.145
R2085 GND.n233 GND.n228 0.145
R2086 GND.n236 GND.n233 0.145
R2087 GND.n239 GND.n236 0.145
R2088 GND.n249 GND.n246 0.145
R2089 GND.n252 GND.n249 0.145
R2090 GND.n255 GND.n252 0.145
R2091 GND.n258 GND.n255 0.145
R2092 GND.n261 GND.n258 0.145
R2093 GND.n267 GND.n264 0.145
R2094 GND.n270 GND.n267 0.145
R2095 GND.n275 GND.n270 0.145
R2096 GND.n278 GND.n275 0.145
R2097 GND.n281 GND.n278 0.145
R2098 GND.n291 GND.n288 0.145
R2099 GND.n294 GND.n291 0.145
R2100 GND.n297 GND.n294 0.145
R2101 GND.n305 GND.n300 0.145
R2102 GND.n308 GND.n305 0.145
R2103 GND.n311 GND.n308 0.145
R2104 GND.n321 GND.n318 0.145
R2105 GND.n324 GND.n321 0.145
R2106 GND.n327 GND.n324 0.145
R2107 GND.n338 GND.n330 0.145
R2108 GND.n677 GND.n674 0.145
R2109 GND.n667 GND.n664 0.145
R2110 GND.n664 GND.n661 0.145
R2111 GND.n661 GND.n658 0.145
R2112 GND.n655 GND.n652 0.145
R2113 GND.n652 GND.n647 0.145
R2114 GND.n647 GND.n644 0.145
R2115 GND.n637 GND.n634 0.145
R2116 GND.n634 GND.n631 0.145
R2117 GND.n631 GND.n628 0.145
R2118 GND.n625 GND.n622 0.145
R2119 GND.n622 GND.n617 0.145
R2120 GND.n617 GND.n614 0.145
R2121 GND.n607 GND.n604 0.145
R2122 GND.n604 GND.n601 0.145
R2123 GND.n601 GND.n598 0.145
R2124 GND.n595 GND.n592 0.145
R2125 GND.n592 GND.n587 0.145
R2126 GND.n587 GND.n584 0.145
R2127 GND.n577 GND.n574 0.145
R2128 GND.n574 GND.n571 0.145
R2129 GND.n571 GND.n568 0.145
R2130 GND.n568 GND.n565 0.145
R2131 GND.n565 GND.n562 0.145
R2132 GND.n559 GND.n556 0.145
R2133 GND.n556 GND.n553 0.145
R2134 GND.n553 GND.n550 0.145
R2135 GND.n550 GND.n545 0.145
R2136 GND.n545 GND.n542 0.145
R2137 GND.n535 GND.n532 0.145
R2138 GND.n532 GND.n529 0.145
R2139 GND.n529 GND.n526 0.145
R2140 GND.n523 GND.n520 0.145
R2141 GND.n520 GND.n512 0.145
R2142 GND.n512 GND.n509 0.145
R2143 GND.n502 GND.n499 0.145
R2144 GND.n499 GND.n496 0.145
R2145 GND.n496 GND.n493 0.145
R2146 GND.n490 GND.n487 0.145
R2147 GND.n487 GND.n482 0.145
R2148 GND.n482 GND.n479 0.145
R2149 GND.n472 GND.n469 0.145
R2150 GND.n469 GND.n466 0.145
R2151 GND.n466 GND.n463 0.145
R2152 GND.n460 GND.n457 0.145
R2153 GND.n457 GND.n452 0.145
R2154 GND.n452 GND.n449 0.145
R2155 GND.n442 GND.n439 0.145
R2156 GND.n439 GND.n436 0.145
R2157 GND.n436 GND.n433 0.145
R2158 GND.n430 GND.n427 0.145
R2159 GND.n427 GND.n419 0.145
R2160 GND.n419 GND.n416 0.145
R2161 GND.n409 GND.n406 0.145
R2162 GND.n406 GND.n403 0.145
R2163 GND.n403 GND.n400 0.145
R2164 GND.n397 GND.n394 0.145
R2165 GND.n394 GND.n386 0.145
R2166 GND.n386 GND.n383 0.145
R2167 GND.n376 GND.n373 0.145
R2168 GND.n373 GND.n370 0.145
R2169 GND.n370 GND.n367 0.145
R2170 GND.n367 GND.n364 0.145
R2171 GND.n364 GND.n361 0.145
R2172 GND.n358 GND.n355 0.145
R2173 GND.n355 GND.n352 0.145
R2174 GND.n352 GND.n349 0.145
R2175 GND.n349 GND.n344 0.145
R2176 GND.n344 GND.n341 0.145
R2177 GND GND.n677 0.082
R2178 GND GND.n338 0.062
R2179 a_10429_1050.n3 a_10429_1050.t5 480.392
R2180 a_10429_1050.n3 a_10429_1050.t7 403.272
R2181 a_10429_1050.n4 a_10429_1050.t6 283.48
R2182 a_10429_1050.n7 a_10429_1050.n5 217.114
R2183 a_10429_1050.n5 a_10429_1050.n4 153.315
R2184 a_10429_1050.n5 a_10429_1050.n2 152.499
R2185 a_10429_1050.n4 a_10429_1050.n3 98.447
R2186 a_10429_1050.n2 a_10429_1050.n1 76.002
R2187 a_10429_1050.n7 a_10429_1050.n6 15.218
R2188 a_10429_1050.n0 a_10429_1050.t2 14.282
R2189 a_10429_1050.n0 a_10429_1050.t4 14.282
R2190 a_10429_1050.n1 a_10429_1050.t0 14.282
R2191 a_10429_1050.n1 a_10429_1050.t1 14.282
R2192 a_10429_1050.n2 a_10429_1050.n0 12.85
R2193 a_10429_1050.n8 a_10429_1050.n7 12.014
R2194 a_8731_187.n5 a_8731_187.t8 512.525
R2195 a_8731_187.n3 a_8731_187.t11 472.359
R2196 a_8731_187.n1 a_8731_187.t13 472.359
R2197 a_8731_187.n3 a_8731_187.t5 384.527
R2198 a_8731_187.n1 a_8731_187.t10 384.527
R2199 a_8731_187.n5 a_8731_187.t12 371.139
R2200 a_8731_187.n6 a_8731_187.t7 340.774
R2201 a_8731_187.n4 a_8731_187.t6 294.278
R2202 a_8731_187.n2 a_8731_187.t9 294.278
R2203 a_8731_187.n10 a_8731_187.n9 285.437
R2204 a_8731_187.n6 a_8731_187.n5 109.607
R2205 a_8731_187.n11 a_8731_187.n10 99.394
R2206 a_8731_187.n7 a_8731_187.n6 82.484
R2207 a_8731_187.n8 a_8731_187.n2 80.307
R2208 a_8731_187.n12 a_8731_187.n11 76.001
R2209 a_8731_187.n7 a_8731_187.n4 76
R2210 a_8731_187.n10 a_8731_187.n8 76
R2211 a_8731_187.n4 a_8731_187.n3 56.954
R2212 a_8731_187.n2 a_8731_187.n1 56.954
R2213 a_8731_187.n0 a_8731_187.t4 14.282
R2214 a_8731_187.n0 a_8731_187.t1 14.282
R2215 a_8731_187.t3 a_8731_187.n12 14.282
R2216 a_8731_187.n12 a_8731_187.t2 14.282
R2217 a_8731_187.n11 a_8731_187.n0 12.85
R2218 a_8731_187.n8 a_8731_187.n7 2.947
R2219 a_7595_411.n4 a_7595_411.t8 475.572
R2220 a_7595_411.n8 a_7595_411.t11 472.359
R2221 a_7595_411.n3 a_7595_411.t10 469.145
R2222 a_7595_411.n8 a_7595_411.t7 384.527
R2223 a_7595_411.n4 a_7595_411.t5 384.527
R2224 a_7595_411.n3 a_7595_411.t13 384.527
R2225 a_7595_411.n5 a_7595_411.t9 294.278
R2226 a_7595_411.n11 a_7595_411.n2 232.158
R2227 a_7595_411.n9 a_7595_411.n8 189.719
R2228 a_7595_411.n9 a_7595_411.t6 161.513
R2229 a_7595_411.n7 a_7595_411.t12 161.513
R2230 a_7595_411.n6 a_7595_411.n5 156.851
R2231 a_7595_411.n13 a_7595_411.n11 137.455
R2232 a_7595_411.n7 a_7595_411.n6 132.764
R2233 a_7595_411.n10 a_7595_411.n7 93.638
R2234 a_7595_411.n10 a_7595_411.n9 78.947
R2235 a_7595_411.n2 a_7595_411.n1 76.002
R2236 a_7595_411.n11 a_7595_411.n10 76
R2237 a_7595_411.n5 a_7595_411.n4 57.842
R2238 a_7595_411.n6 a_7595_411.n3 56.833
R2239 a_7595_411.n13 a_7595_411.n12 15.218
R2240 a_7595_411.n0 a_7595_411.t0 14.282
R2241 a_7595_411.n0 a_7595_411.t2 14.282
R2242 a_7595_411.n1 a_7595_411.t1 14.282
R2243 a_7595_411.n1 a_7595_411.t3 14.282
R2244 a_7595_411.n2 a_7595_411.n0 12.85
R2245 a_7595_411.n14 a_7595_411.n13 12.014
R2246 a_13757_1051.n4 a_13757_1051.n3 196.002
R2247 a_13757_1051.n2 a_13757_1051.t5 89.553
R2248 a_13757_1051.n4 a_13757_1051.n0 75.271
R2249 a_13757_1051.n3 a_13757_1051.n2 75.214
R2250 a_13757_1051.n5 a_13757_1051.n4 36.519
R2251 a_13757_1051.n3 a_13757_1051.t1 14.338
R2252 a_13757_1051.n1 a_13757_1051.t6 14.282
R2253 a_13757_1051.n1 a_13757_1051.t3 14.282
R2254 a_13757_1051.n0 a_13757_1051.t7 14.282
R2255 a_13757_1051.n0 a_13757_1051.t4 14.282
R2256 a_13757_1051.n5 a_13757_1051.t2 14.282
R2257 a_13757_1051.t0 a_13757_1051.n5 14.282
R2258 a_13757_1051.n2 a_13757_1051.n1 12.119
R2259 QN.n14 QN.n13 216.728
R2260 QN.n14 QN.n2 126.664
R2261 QN.n11 QN.n10 98.501
R2262 QN.n11 QN.n6 96.417
R2263 QN.n13 QN.n11 78.403
R2264 QN.n15 QN.n14 76
R2265 QN.n2 QN.n1 75.271
R2266 QN.n13 QN.n12 42.274
R2267 QN.n6 QN.n5 30
R2268 QN.n10 QN.n9 30
R2269 QN.n4 QN.n3 24.383
R2270 QN.n8 QN.n7 24.383
R2271 QN.n6 QN.n4 23.684
R2272 QN.n10 QN.n8 23.684
R2273 QN.n0 QN.t3 14.282
R2274 QN.n0 QN.t4 14.282
R2275 QN.n1 QN.t2 14.282
R2276 QN.n1 QN.t1 14.282
R2277 QN.n2 QN.n0 12.119
R2278 QN.n15 QN 0.046
R2279 a_147_187.n7 a_147_187.t7 512.525
R2280 a_147_187.n5 a_147_187.t6 472.359
R2281 a_147_187.n3 a_147_187.t9 472.359
R2282 a_147_187.n5 a_147_187.t10 384.527
R2283 a_147_187.n3 a_147_187.t11 384.527
R2284 a_147_187.n7 a_147_187.t12 371.139
R2285 a_147_187.n8 a_147_187.t8 340.774
R2286 a_147_187.n6 a_147_187.t13 294.278
R2287 a_147_187.n4 a_147_187.t5 294.278
R2288 a_147_187.n13 a_147_187.n11 270.22
R2289 a_147_187.n8 a_147_187.n7 109.607
R2290 a_147_187.n11 a_147_187.n2 99.394
R2291 a_147_187.n9 a_147_187.n8 82.484
R2292 a_147_187.n10 a_147_187.n4 80.307
R2293 a_147_187.n2 a_147_187.n1 76.002
R2294 a_147_187.n9 a_147_187.n6 76
R2295 a_147_187.n11 a_147_187.n10 76
R2296 a_147_187.n6 a_147_187.n5 56.954
R2297 a_147_187.n4 a_147_187.n3 56.954
R2298 a_147_187.n13 a_147_187.n12 15.218
R2299 a_147_187.n0 a_147_187.t4 14.282
R2300 a_147_187.n0 a_147_187.t2 14.282
R2301 a_147_187.n1 a_147_187.t0 14.282
R2302 a_147_187.n1 a_147_187.t1 14.282
R2303 a_147_187.n2 a_147_187.n0 12.85
R2304 a_147_187.n14 a_147_187.n13 12.014
R2305 a_147_187.n10 a_147_187.n9 2.947
R2306 a_3738_101.n12 a_3738_101.n11 26.811
R2307 a_3738_101.n6 a_3738_101.n5 24.977
R2308 a_3738_101.n2 a_3738_101.n1 24.877
R2309 a_3738_101.t0 a_3738_101.n2 12.677
R2310 a_3738_101.t0 a_3738_101.n3 11.595
R2311 a_3738_101.t1 a_3738_101.n8 8.137
R2312 a_3738_101.t0 a_3738_101.n4 7.273
R2313 a_3738_101.t0 a_3738_101.n0 6.109
R2314 a_3738_101.t1 a_3738_101.n7 4.864
R2315 a_3738_101.t0 a_3738_101.n12 2.074
R2316 a_3738_101.n7 a_3738_101.n6 1.13
R2317 a_3738_101.n12 a_3738_101.t1 0.937
R2318 a_3738_101.t1 a_3738_101.n10 0.804
R2319 a_3738_101.n10 a_3738_101.n9 0.136
R2320 a_7364_101.n5 a_7364_101.n4 24.877
R2321 a_7364_101.t0 a_7364_101.n5 12.677
R2322 a_7364_101.t0 a_7364_101.n3 11.595
R2323 a_7364_101.t0 a_7364_101.n6 8.137
R2324 a_7364_101.n2 a_7364_101.n0 4.031
R2325 a_7364_101.n2 a_7364_101.n1 3.644
R2326 a_7364_101.t0 a_7364_101.n2 1.093
R2327 a_7469_1050.n0 a_7469_1050.t6 480.392
R2328 a_7469_1050.n0 a_7469_1050.t7 403.272
R2329 a_7469_1050.n1 a_7469_1050.t5 310.033
R2330 a_7469_1050.n3 a_7469_1050.n2 258.884
R2331 a_7469_1050.n3 a_7469_1050.n1 153.315
R2332 a_7469_1050.n5 a_7469_1050.n3 125.947
R2333 a_7469_1050.n5 a_7469_1050.n4 76.002
R2334 a_7469_1050.n1 a_7469_1050.n0 71.894
R2335 a_7469_1050.n4 a_7469_1050.t0 14.282
R2336 a_7469_1050.n4 a_7469_1050.t4 14.282
R2337 a_7469_1050.n6 a_7469_1050.t2 14.282
R2338 a_7469_1050.t3 a_7469_1050.n6 14.282
R2339 a_7469_1050.n6 a_7469_1050.n5 12.848
R2340 a_10324_101.n12 a_10324_101.n11 26.811
R2341 a_10324_101.n6 a_10324_101.n5 24.977
R2342 a_10324_101.n2 a_10324_101.n1 24.877
R2343 a_10324_101.t0 a_10324_101.n2 12.677
R2344 a_10324_101.t0 a_10324_101.n3 11.595
R2345 a_10324_101.t1 a_10324_101.n8 8.137
R2346 a_10324_101.t0 a_10324_101.n4 7.273
R2347 a_10324_101.t0 a_10324_101.n0 6.109
R2348 a_10324_101.t1 a_10324_101.n7 4.864
R2349 a_10324_101.t0 a_10324_101.n12 2.074
R2350 a_10324_101.n7 a_10324_101.n6 1.13
R2351 a_10324_101.n12 a_10324_101.t1 0.937
R2352 a_10324_101.t1 a_10324_101.n10 0.804
R2353 a_10324_101.n10 a_10324_101.n9 0.136
R2354 a_9183_989.n0 a_9183_989.t6 480.392
R2355 a_9183_989.n2 a_9183_989.t7 454.685
R2356 a_9183_989.n2 a_9183_989.t5 428.979
R2357 a_9183_989.n0 a_9183_989.t10 403.272
R2358 a_9183_989.n1 a_9183_989.t8 283.48
R2359 a_9183_989.n3 a_9183_989.t9 237.959
R2360 a_9183_989.n9 a_9183_989.n8 210.592
R2361 a_9183_989.n11 a_9183_989.n9 152.499
R2362 a_9183_989.n3 a_9183_989.n2 98.447
R2363 a_9183_989.n1 a_9183_989.n0 98.447
R2364 a_9183_989.n4 a_9183_989.n3 78.947
R2365 a_9183_989.n4 a_9183_989.n1 77.315
R2366 a_9183_989.n11 a_9183_989.n10 76.002
R2367 a_9183_989.n9 a_9183_989.n4 76
R2368 a_9183_989.n8 a_9183_989.n7 30
R2369 a_9183_989.n6 a_9183_989.n5 24.383
R2370 a_9183_989.n8 a_9183_989.n6 23.684
R2371 a_9183_989.n10 a_9183_989.t4 14.282
R2372 a_9183_989.n10 a_9183_989.t3 14.282
R2373 a_9183_989.t2 a_9183_989.n12 14.282
R2374 a_9183_989.n12 a_9183_989.t1 14.282
R2375 a_9183_989.n12 a_9183_989.n11 12.848
R2376 a_8861_1050.n4 a_8861_1050.t7 480.392
R2377 a_8861_1050.n2 a_8861_1050.t12 480.392
R2378 a_8861_1050.n4 a_8861_1050.t10 403.272
R2379 a_8861_1050.n2 a_8861_1050.t11 403.272
R2380 a_8861_1050.n5 a_8861_1050.t8 310.033
R2381 a_8861_1050.n3 a_8861_1050.t9 310.033
R2382 a_8861_1050.n11 a_8861_1050.n10 239.657
R2383 a_8861_1050.n12 a_8861_1050.n11 144.246
R2384 a_8861_1050.n6 a_8861_1050.n3 83.3
R2385 a_8861_1050.n14 a_8861_1050.n13 79.231
R2386 a_8861_1050.n11 a_8861_1050.n6 77.315
R2387 a_8861_1050.n6 a_8861_1050.n5 76
R2388 a_8861_1050.n5 a_8861_1050.n4 71.894
R2389 a_8861_1050.n3 a_8861_1050.n2 71.894
R2390 a_8861_1050.n13 a_8861_1050.n12 63.152
R2391 a_8861_1050.n10 a_8861_1050.n9 30
R2392 a_8861_1050.n8 a_8861_1050.n7 24.383
R2393 a_8861_1050.n10 a_8861_1050.n8 23.684
R2394 a_8861_1050.n12 a_8861_1050.n1 16.08
R2395 a_8861_1050.n13 a_8861_1050.n0 16.08
R2396 a_8861_1050.n1 a_8861_1050.t4 14.282
R2397 a_8861_1050.n1 a_8861_1050.t3 14.282
R2398 a_8861_1050.n0 a_8861_1050.t6 14.282
R2399 a_8861_1050.n0 a_8861_1050.t2 14.282
R2400 a_8861_1050.t1 a_8861_1050.n14 14.282
R2401 a_8861_1050.n14 a_8861_1050.t0 14.282
R2402 CLK.n15 CLK.t5 472.359
R2403 CLK.n6 CLK.t6 472.359
R2404 CLK.n0 CLK.t16 472.359
R2405 CLK.n20 CLK.t2 459.505
R2406 CLK.n11 CLK.t12 459.505
R2407 CLK.n2 CLK.t17 459.505
R2408 CLK.n20 CLK.t13 384.527
R2409 CLK.n15 CLK.t15 384.527
R2410 CLK.n11 CLK.t0 384.527
R2411 CLK.n6 CLK.t7 384.527
R2412 CLK.n2 CLK.t1 384.527
R2413 CLK.n0 CLK.t9 384.527
R2414 CLK.n21 CLK.t8 322.152
R2415 CLK.n12 CLK.t11 322.151
R2416 CLK.n3 CLK.t4 322.151
R2417 CLK.n1 CLK.t14 321.724
R2418 CLK.n17 CLK.t10 319.581
R2419 CLK.n8 CLK.t3 319.581
R2420 CLK.n9 CLK.n8 75.621
R2421 CLK.n18 CLK.n17 75.621
R2422 CLK.n22 CLK.n21 49.342
R2423 CLK.n4 CLK.n3 49.342
R2424 CLK.n13 CLK.n12 49.342
R2425 CLK.n4 CLK.n1 44.933
R2426 CLK.n21 CLK.n20 27.599
R2427 CLK.n3 CLK.n2 27.599
R2428 CLK.n12 CLK.n11 27.599
R2429 CLK.n1 CLK.n0 23.329
R2430 CLK.n16 CLK.n15 21.176
R2431 CLK.n7 CLK.n6 21.176
R2432 CLK.n13 CLK.n10 8.078
R2433 CLK.n22 CLK.n19 8.078
R2434 CLK.n14 CLK.n13 7.797
R2435 CLK.n5 CLK.n4 7.564
R2436 CLK.n17 CLK.n16 4.419
R2437 CLK.n8 CLK.n7 4.419
R2438 CLK.n22 CLK 0.046
R2439 CLK.n10 CLK.n9 0.038
R2440 CLK.n19 CLK.n18 0.038
R2441 CLK.n9 CLK.n5 0.008
R2442 CLK.n18 CLK.n14 0.008
R2443 a_4569_1050.n3 a_4569_1050.t7 480.392
R2444 a_4569_1050.n1 a_4569_1050.t8 480.392
R2445 a_4569_1050.n3 a_4569_1050.t11 403.272
R2446 a_4569_1050.n1 a_4569_1050.t12 403.272
R2447 a_4569_1050.n4 a_4569_1050.t9 310.033
R2448 a_4569_1050.n2 a_4569_1050.t10 310.033
R2449 a_4569_1050.n7 a_4569_1050.n6 261.396
R2450 a_4569_1050.n8 a_4569_1050.n7 144.246
R2451 a_4569_1050.n5 a_4569_1050.n2 83.3
R2452 a_4569_1050.n10 a_4569_1050.n9 79.232
R2453 a_4569_1050.n7 a_4569_1050.n5 77.315
R2454 a_4569_1050.n5 a_4569_1050.n4 76
R2455 a_4569_1050.n4 a_4569_1050.n3 71.894
R2456 a_4569_1050.n2 a_4569_1050.n1 71.894
R2457 a_4569_1050.n10 a_4569_1050.n8 63.152
R2458 a_4569_1050.n8 a_4569_1050.n0 16.08
R2459 a_4569_1050.n11 a_4569_1050.n10 16.078
R2460 a_4569_1050.n0 a_4569_1050.t4 14.282
R2461 a_4569_1050.n0 a_4569_1050.t2 14.282
R2462 a_4569_1050.n9 a_4569_1050.t3 14.282
R2463 a_4569_1050.n9 a_4569_1050.t5 14.282
R2464 a_4569_1050.n11 a_4569_1050.t0 14.282
R2465 a_4569_1050.t1 a_4569_1050.n11 14.282
R2466 a_4439_187.n4 a_4439_187.t10 512.525
R2467 a_4439_187.n2 a_4439_187.t5 472.359
R2468 a_4439_187.n0 a_4439_187.t6 472.359
R2469 a_4439_187.n2 a_4439_187.t11 384.527
R2470 a_4439_187.n0 a_4439_187.t12 384.527
R2471 a_4439_187.n4 a_4439_187.t13 371.139
R2472 a_4439_187.n5 a_4439_187.t8 340.774
R2473 a_4439_187.n3 a_4439_187.t7 294.278
R2474 a_4439_187.n1 a_4439_187.t9 294.278
R2475 a_4439_187.n12 a_4439_187.n11 263.698
R2476 a_4439_187.n5 a_4439_187.n4 109.607
R2477 a_4439_187.n14 a_4439_187.n12 99.394
R2478 a_4439_187.n6 a_4439_187.n5 82.484
R2479 a_4439_187.n7 a_4439_187.n1 80.307
R2480 a_4439_187.n14 a_4439_187.n13 76.002
R2481 a_4439_187.n6 a_4439_187.n3 76
R2482 a_4439_187.n12 a_4439_187.n7 76
R2483 a_4439_187.n3 a_4439_187.n2 56.954
R2484 a_4439_187.n1 a_4439_187.n0 56.954
R2485 a_4439_187.n11 a_4439_187.n10 30
R2486 a_4439_187.n9 a_4439_187.n8 24.383
R2487 a_4439_187.n11 a_4439_187.n9 23.684
R2488 a_4439_187.n13 a_4439_187.t3 14.282
R2489 a_4439_187.n13 a_4439_187.t4 14.282
R2490 a_4439_187.t2 a_4439_187.n15 14.282
R2491 a_4439_187.n15 a_4439_187.t1 14.282
R2492 a_4439_187.n15 a_4439_187.n14 12.848
R2493 a_4439_187.n7 a_4439_187.n6 2.947
R2494 a_6137_1050.n0 a_6137_1050.t5 480.392
R2495 a_6137_1050.n0 a_6137_1050.t6 403.272
R2496 a_6137_1050.n1 a_6137_1050.t7 283.48
R2497 a_6137_1050.n6 a_6137_1050.n5 210.592
R2498 a_6137_1050.n6 a_6137_1050.n1 153.315
R2499 a_6137_1050.n8 a_6137_1050.n6 152.499
R2500 a_6137_1050.n1 a_6137_1050.n0 98.447
R2501 a_6137_1050.n8 a_6137_1050.n7 76.002
R2502 a_6137_1050.n5 a_6137_1050.n4 30
R2503 a_6137_1050.n3 a_6137_1050.n2 24.383
R2504 a_6137_1050.n5 a_6137_1050.n3 23.684
R2505 a_6137_1050.n7 a_6137_1050.t4 14.282
R2506 a_6137_1050.n7 a_6137_1050.t0 14.282
R2507 a_6137_1050.t3 a_6137_1050.n9 14.282
R2508 a_6137_1050.n9 a_6137_1050.t2 14.282
R2509 a_6137_1050.n9 a_6137_1050.n8 12.848
R2510 a_1845_1050.n1 a_1845_1050.t6 480.392
R2511 a_1845_1050.n1 a_1845_1050.t7 403.272
R2512 a_1845_1050.n2 a_1845_1050.t5 283.48
R2513 a_1845_1050.n7 a_1845_1050.n6 210.592
R2514 a_1845_1050.n7 a_1845_1050.n2 153.315
R2515 a_1845_1050.n8 a_1845_1050.n7 152.499
R2516 a_1845_1050.n2 a_1845_1050.n1 98.447
R2517 a_1845_1050.n9 a_1845_1050.n8 76.001
R2518 a_1845_1050.n6 a_1845_1050.n5 30
R2519 a_1845_1050.n4 a_1845_1050.n3 24.383
R2520 a_1845_1050.n6 a_1845_1050.n4 23.684
R2521 a_1845_1050.n0 a_1845_1050.t3 14.282
R2522 a_1845_1050.n0 a_1845_1050.t2 14.282
R2523 a_1845_1050.n9 a_1845_1050.t0 14.282
R2524 a_1845_1050.t1 a_1845_1050.n9 14.282
R2525 a_1845_1050.n8 a_1845_1050.n0 12.85
R2526 a_8675_103.n1 a_8675_103.n0 25.576
R2527 a_8675_103.n3 a_8675_103.n2 9.111
R2528 a_8675_103.n7 a_8675_103.n5 7.859
R2529 a_8675_103.t0 a_8675_103.n7 3.034
R2530 a_8675_103.n5 a_8675_103.n3 1.964
R2531 a_8675_103.n5 a_8675_103.n4 1.964
R2532 a_8675_103.t0 a_8675_103.n1 1.871
R2533 a_8675_103.n7 a_8675_103.n6 0.443
R2534 a_11887_411.n2 a_11887_411.t12 512.525
R2535 a_11887_411.n0 a_11887_411.t6 477.179
R2536 a_11887_411.n5 a_11887_411.t7 472.359
R2537 a_11887_411.n0 a_11887_411.t11 406.485
R2538 a_11887_411.n5 a_11887_411.t9 384.527
R2539 a_11887_411.n2 a_11887_411.t5 371.139
R2540 a_11887_411.n1 a_11887_411.t8 363.924
R2541 a_11887_411.n4 a_11887_411.t10 303.606
R2542 a_11887_411.n6 a_11887_411.t13 267.725
R2543 a_11887_411.n12 a_11887_411.n11 237.145
R2544 a_11887_411.n14 a_11887_411.n12 125.947
R2545 a_11887_411.n3 a_11887_411.n1 101.359
R2546 a_11887_411.n6 a_11887_411.n5 83.507
R2547 a_11887_411.n7 a_11887_411.n6 78.947
R2548 a_11887_411.n7 a_11887_411.n4 77.043
R2549 a_11887_411.n14 a_11887_411.n13 76.002
R2550 a_11887_411.n12 a_11887_411.n7 76
R2551 a_11887_411.n3 a_11887_411.n2 71.88
R2552 a_11887_411.n4 a_11887_411.n3 53.891
R2553 a_11887_411.n11 a_11887_411.n10 30
R2554 a_11887_411.n9 a_11887_411.n8 24.383
R2555 a_11887_411.n11 a_11887_411.n9 23.684
R2556 a_11887_411.n1 a_11887_411.n0 15.776
R2557 a_11887_411.n13 a_11887_411.t0 14.282
R2558 a_11887_411.n13 a_11887_411.t4 14.282
R2559 a_11887_411.n15 a_11887_411.t1 14.282
R2560 a_11887_411.t2 a_11887_411.n15 14.282
R2561 a_11887_411.n15 a_11887_411.n14 12.848
R2562 a_13093_1051.n3 a_13093_1051.n2 195.987
R2563 a_13093_1051.n4 a_13093_1051.t5 89.553
R2564 a_13093_1051.n2 a_13093_1051.n1 75.271
R2565 a_13093_1051.n4 a_13093_1051.n3 75.214
R2566 a_13093_1051.n2 a_13093_1051.n0 36.519
R2567 a_13093_1051.n3 a_13093_1051.t0 14.338
R2568 a_13093_1051.n0 a_13093_1051.t7 14.282
R2569 a_13093_1051.n0 a_13093_1051.t6 14.282
R2570 a_13093_1051.n1 a_13093_1051.t2 14.282
R2571 a_13093_1051.n1 a_13093_1051.t3 14.282
R2572 a_13093_1051.n5 a_13093_1051.t4 14.282
R2573 a_13093_1051.t1 a_13093_1051.n5 14.282
R2574 a_13093_1051.n5 a_13093_1051.n4 12.122
R2575 a_4891_989.n0 a_4891_989.t9 480.392
R2576 a_4891_989.n2 a_4891_989.t7 454.685
R2577 a_4891_989.n2 a_4891_989.t8 428.979
R2578 a_4891_989.n0 a_4891_989.t5 403.272
R2579 a_4891_989.n1 a_4891_989.t10 283.48
R2580 a_4891_989.n3 a_4891_989.t6 237.959
R2581 a_4891_989.n9 a_4891_989.n8 210.592
R2582 a_4891_989.n11 a_4891_989.n9 152.499
R2583 a_4891_989.n3 a_4891_989.n2 98.447
R2584 a_4891_989.n1 a_4891_989.n0 98.447
R2585 a_4891_989.n4 a_4891_989.n3 78.947
R2586 a_4891_989.n4 a_4891_989.n1 77.315
R2587 a_4891_989.n11 a_4891_989.n10 76.002
R2588 a_4891_989.n9 a_4891_989.n4 76
R2589 a_4891_989.n8 a_4891_989.n7 30
R2590 a_4891_989.n6 a_4891_989.n5 24.383
R2591 a_4891_989.n8 a_4891_989.n6 23.684
R2592 a_4891_989.n10 a_4891_989.t4 14.282
R2593 a_4891_989.n10 a_4891_989.t3 14.282
R2594 a_4891_989.t1 a_4891_989.n12 14.282
R2595 a_4891_989.n12 a_4891_989.t0 14.282
R2596 a_4891_989.n12 a_4891_989.n11 12.848
R2597 a_8030_101.t0 a_8030_101.n1 34.62
R2598 a_8030_101.t0 a_8030_101.n0 8.137
R2599 a_8030_101.t0 a_8030_101.n2 4.69
R2600 a_1074_101.t0 a_1074_101.n1 34.62
R2601 a_1074_101.t0 a_1074_101.n0 8.137
R2602 a_1074_101.t0 a_1074_101.n2 4.69
R2603 a_277_1050.n3 a_277_1050.t8 480.392
R2604 a_277_1050.n1 a_277_1050.t10 480.392
R2605 a_277_1050.n3 a_277_1050.t11 403.272
R2606 a_277_1050.n1 a_277_1050.t7 403.272
R2607 a_277_1050.n4 a_277_1050.t9 310.033
R2608 a_277_1050.n2 a_277_1050.t12 310.033
R2609 a_277_1050.n10 a_277_1050.n9 239.657
R2610 a_277_1050.n11 a_277_1050.n10 144.246
R2611 a_277_1050.n5 a_277_1050.n2 83.3
R2612 a_277_1050.n13 a_277_1050.n12 79.232
R2613 a_277_1050.n10 a_277_1050.n5 77.315
R2614 a_277_1050.n5 a_277_1050.n4 76
R2615 a_277_1050.n4 a_277_1050.n3 71.894
R2616 a_277_1050.n2 a_277_1050.n1 71.894
R2617 a_277_1050.n13 a_277_1050.n11 63.152
R2618 a_277_1050.n9 a_277_1050.n8 30
R2619 a_277_1050.n7 a_277_1050.n6 24.383
R2620 a_277_1050.n9 a_277_1050.n7 23.684
R2621 a_277_1050.n11 a_277_1050.n0 16.08
R2622 a_277_1050.n14 a_277_1050.n13 16.078
R2623 a_277_1050.n0 a_277_1050.t4 14.282
R2624 a_277_1050.n0 a_277_1050.t3 14.282
R2625 a_277_1050.n12 a_277_1050.t6 14.282
R2626 a_277_1050.n12 a_277_1050.t5 14.282
R2627 a_277_1050.t1 a_277_1050.n14 14.282
R2628 a_277_1050.n14 a_277_1050.t0 14.282
R2629 a_3177_1050.n0 a_3177_1050.t7 480.392
R2630 a_3177_1050.n0 a_3177_1050.t5 403.272
R2631 a_3177_1050.n1 a_3177_1050.t6 310.033
R2632 a_3177_1050.n6 a_3177_1050.n5 237.145
R2633 a_3177_1050.n6 a_3177_1050.n1 153.315
R2634 a_3177_1050.n8 a_3177_1050.n6 125.947
R2635 a_3177_1050.n8 a_3177_1050.n7 76.002
R2636 a_3177_1050.n1 a_3177_1050.n0 71.894
R2637 a_3177_1050.n5 a_3177_1050.n4 30
R2638 a_3177_1050.n3 a_3177_1050.n2 24.383
R2639 a_3177_1050.n5 a_3177_1050.n3 23.684
R2640 a_3177_1050.n7 a_3177_1050.t3 14.282
R2641 a_3177_1050.n7 a_3177_1050.t4 14.282
R2642 a_3177_1050.n9 a_3177_1050.t0 14.282
R2643 a_3177_1050.t1 a_3177_1050.n9 14.282
R2644 a_3177_1050.n9 a_3177_1050.n8 12.848
R2645 a_12322_101.t0 a_12322_101.n1 34.62
R2646 a_12322_101.t0 a_12322_101.n0 8.137
R2647 a_12322_101.t0 a_12322_101.n2 4.69
R2648 a_2406_101.n12 a_2406_101.n11 26.811
R2649 a_2406_101.n6 a_2406_101.n5 24.977
R2650 a_2406_101.n2 a_2406_101.n1 24.877
R2651 a_2406_101.t0 a_2406_101.n2 12.677
R2652 a_2406_101.t0 a_2406_101.n3 11.595
R2653 a_2406_101.t1 a_2406_101.n8 8.137
R2654 a_2406_101.t0 a_2406_101.n4 7.273
R2655 a_2406_101.t0 a_2406_101.n0 6.109
R2656 a_2406_101.t1 a_2406_101.n7 4.864
R2657 a_2406_101.t0 a_2406_101.n12 2.074
R2658 a_2406_101.n7 a_2406_101.n6 1.13
R2659 a_2406_101.n12 a_2406_101.t1 0.937
R2660 a_2406_101.t1 a_2406_101.n10 0.804
R2661 a_2406_101.n10 a_2406_101.n9 0.136
R2662 a_372_210.n10 a_372_210.n8 82.852
R2663 a_372_210.n7 a_372_210.n6 32.833
R2664 a_372_210.n8 a_372_210.t1 32.416
R2665 a_372_210.n10 a_372_210.n9 27.2
R2666 a_372_210.n11 a_372_210.n0 23.498
R2667 a_372_210.n3 a_372_210.n2 23.284
R2668 a_372_210.n11 a_372_210.n10 22.4
R2669 a_372_210.n7 a_372_210.n4 19.017
R2670 a_372_210.n6 a_372_210.n5 13.494
R2671 a_372_210.t1 a_372_210.n1 7.04
R2672 a_372_210.t1 a_372_210.n3 5.727
R2673 a_372_210.n8 a_372_210.n7 1.435
R2674 a_11761_1050.n0 a_11761_1050.t6 480.392
R2675 a_11761_1050.n0 a_11761_1050.t5 403.272
R2676 a_11761_1050.n1 a_11761_1050.t7 363.924
R2677 a_11761_1050.n6 a_11761_1050.n5 290.251
R2678 a_11761_1050.n6 a_11761_1050.n1 126.657
R2679 a_11761_1050.n8 a_11761_1050.n7 76.002
R2680 a_11761_1050.n8 a_11761_1050.n6 72.841
R2681 a_11761_1050.n5 a_11761_1050.n4 30
R2682 a_11761_1050.n3 a_11761_1050.n2 24.383
R2683 a_11761_1050.n5 a_11761_1050.n3 23.684
R2684 a_11761_1050.n1 a_11761_1050.n0 15.545
R2685 a_11761_1050.n7 a_11761_1050.t3 14.282
R2686 a_11761_1050.n7 a_11761_1050.t4 14.282
R2687 a_11761_1050.t2 a_11761_1050.n9 14.282
R2688 a_11761_1050.n9 a_11761_1050.t1 14.282
R2689 a_11761_1050.n9 a_11761_1050.n8 12.848
R2690 a_9658_101.t0 a_9658_101.n1 34.62
R2691 a_9658_101.t0 a_9658_101.n0 8.137
R2692 a_9658_101.t0 a_9658_101.n2 4.69
R2693 a_4664_210.n9 a_4664_210.n7 82.852
R2694 a_4664_210.n3 a_4664_210.n1 44.628
R2695 a_4664_210.t0 a_4664_210.n9 32.417
R2696 a_4664_210.n7 a_4664_210.n6 27.2
R2697 a_4664_210.n5 a_4664_210.n4 23.498
R2698 a_4664_210.n3 a_4664_210.n2 23.284
R2699 a_4664_210.n7 a_4664_210.n5 22.4
R2700 a_4664_210.t0 a_4664_210.n11 20.241
R2701 a_4664_210.n11 a_4664_210.n10 13.494
R2702 a_4664_210.t0 a_4664_210.n0 8.137
R2703 a_4664_210.t0 a_4664_210.n3 5.727
R2704 a_4664_210.n9 a_4664_210.n8 1.435
R2705 a_3072_101.t0 a_3072_101.n1 34.62
R2706 a_3072_101.t0 a_3072_101.n0 8.137
R2707 a_3072_101.t0 a_3072_101.n2 4.69
R2708 a_6698_101.n12 a_6698_101.n11 26.811
R2709 a_6698_101.n6 a_6698_101.n5 24.977
R2710 a_6698_101.n2 a_6698_101.n1 24.877
R2711 a_6698_101.t0 a_6698_101.n2 12.677
R2712 a_6698_101.t0 a_6698_101.n3 11.595
R2713 a_6698_101.t1 a_6698_101.n8 8.137
R2714 a_6698_101.t0 a_6698_101.n4 7.273
R2715 a_6698_101.t0 a_6698_101.n0 6.109
R2716 a_6698_101.t1 a_6698_101.n7 4.864
R2717 a_6698_101.t0 a_6698_101.n12 2.074
R2718 a_6698_101.n7 a_6698_101.n6 1.13
R2719 a_6698_101.n12 a_6698_101.t1 0.937
R2720 a_6698_101.t1 a_6698_101.n10 0.804
R2721 a_6698_101.n10 a_6698_101.n9 0.136
R2722 a_6032_101.t0 a_6032_101.n1 34.62
R2723 a_6032_101.t0 a_6032_101.n0 8.137
R2724 a_6032_101.t0 a_6032_101.n2 4.69
R2725 a_91_103.n1 a_91_103.n0 25.576
R2726 a_91_103.n3 a_91_103.n2 9.111
R2727 a_91_103.n7 a_91_103.n6 2.455
R2728 a_91_103.n5 a_91_103.n3 1.964
R2729 a_91_103.n5 a_91_103.n4 1.964
R2730 a_91_103.t0 a_91_103.n1 1.871
R2731 a_91_103.n7 a_91_103.n5 0.636
R2732 a_91_103.t0 a_91_103.n7 0.246
R2733 a_8956_210.n10 a_8956_210.n8 82.852
R2734 a_8956_210.n11 a_8956_210.n0 49.6
R2735 a_8956_210.n7 a_8956_210.n6 32.833
R2736 a_8956_210.n8 a_8956_210.t1 32.416
R2737 a_8956_210.n10 a_8956_210.n9 27.2
R2738 a_8956_210.n3 a_8956_210.n2 23.284
R2739 a_8956_210.n11 a_8956_210.n10 22.4
R2740 a_8956_210.n7 a_8956_210.n4 19.017
R2741 a_8956_210.n6 a_8956_210.n5 13.494
R2742 a_8956_210.t1 a_8956_210.n1 7.04
R2743 a_8956_210.t1 a_8956_210.n3 5.727
R2744 a_8956_210.n8 a_8956_210.n7 1.435
R2745 a_11656_101.t0 a_11656_101.n1 34.62
R2746 a_11656_101.t0 a_11656_101.n0 8.137
R2747 a_11656_101.t0 a_11656_101.n2 4.69
R2748 a_10990_101.t0 a_10990_101.n1 34.62
R2749 a_10990_101.t0 a_10990_101.n0 8.137
R2750 a_10990_101.t0 a_10990_101.n2 4.69
R2751 a_4383_103.n5 a_4383_103.n4 19.724
R2752 a_4383_103.t0 a_4383_103.n3 11.595
R2753 a_4383_103.t0 a_4383_103.n5 9.207
R2754 a_4383_103.n2 a_4383_103.n1 2.455
R2755 a_4383_103.n2 a_4383_103.n0 1.32
R2756 a_4383_103.t0 a_4383_103.n2 0.246
R2757 a_5366_101.t0 a_5366_101.n1 34.62
R2758 a_5366_101.t0 a_5366_101.n0 8.137
R2759 a_5366_101.t0 a_5366_101.n2 4.69
R2760 a_1740_101.n12 a_1740_101.n11 26.811
R2761 a_1740_101.n6 a_1740_101.n5 24.977
R2762 a_1740_101.n2 a_1740_101.n1 24.877
R2763 a_1740_101.t0 a_1740_101.n2 12.677
R2764 a_1740_101.t0 a_1740_101.n3 11.595
R2765 a_1740_101.t1 a_1740_101.n8 8.137
R2766 a_1740_101.t0 a_1740_101.n4 7.273
R2767 a_1740_101.t0 a_1740_101.n0 6.109
R2768 a_1740_101.t1 a_1740_101.n7 4.864
R2769 a_1740_101.t0 a_1740_101.n12 2.074
R2770 a_1740_101.n7 a_1740_101.n6 1.13
R2771 a_1740_101.n12 a_1740_101.t1 0.937
R2772 a_1740_101.t1 a_1740_101.n10 0.804
R2773 a_1740_101.n10 a_1740_101.n9 0.136
R2774 a_13654_101.t0 a_13654_101.n0 34.602
R2775 a_13654_101.t0 a_13654_101.n1 2.138
R2776 a_12988_101.n13 a_12988_101.n12 26.811
R2777 a_12988_101.n6 a_12988_101.n5 24.977
R2778 a_12988_101.n2 a_12988_101.n1 24.877
R2779 a_12988_101.t0 a_12988_101.n2 12.677
R2780 a_12988_101.t0 a_12988_101.n3 11.595
R2781 a_12988_101.n11 a_12988_101.n10 8.561
R2782 a_12988_101.t0 a_12988_101.n4 7.273
R2783 a_12988_101.n9 a_12988_101.n8 7.066
R2784 a_12988_101.t0 a_12988_101.n0 6.109
R2785 a_12988_101.t1 a_12988_101.n7 4.864
R2786 a_12988_101.t0 a_12988_101.n13 2.074
R2787 a_12988_101.n7 a_12988_101.n6 1.13
R2788 a_12988_101.t1 a_12988_101.n11 0.958
R2789 a_12988_101.n13 a_12988_101.t1 0.937
R2790 a_12988_101.t1 a_12988_101.n9 0.86
C4 VDD GND 54.79fF
C5 a_12988_101.n0 GND 0.02fF
C6 a_12988_101.n1 GND 0.09fF
C7 a_12988_101.n2 GND 0.05fF
C8 a_12988_101.n3 GND 0.06fF
C9 a_12988_101.n4 GND 0.00fF
C10 a_12988_101.n5 GND 0.04fF
C11 a_12988_101.n6 GND 0.05fF
C12 a_12988_101.n7 GND 0.02fF
C13 a_12988_101.n8 GND 0.05fF
C14 a_12988_101.n9 GND 0.09fF
C15 a_12988_101.n10 GND 0.21fF
C16 a_12988_101.n11 GND 0.07fF
C17 a_12988_101.n12 GND 0.04fF
C18 a_12988_101.n13 GND 0.00fF
C19 a_13654_101.n0 GND 0.13fF
C20 a_13654_101.n1 GND 0.13fF
C21 a_1740_101.n0 GND 0.02fF
C22 a_1740_101.n1 GND 0.10fF
C23 a_1740_101.n2 GND 0.06fF
C24 a_1740_101.n3 GND 0.06fF
C25 a_1740_101.n4 GND 0.00fF
C26 a_1740_101.n5 GND 0.04fF
C27 a_1740_101.n6 GND 0.05fF
C28 a_1740_101.n7 GND 0.02fF
C29 a_1740_101.n8 GND 0.05fF
C30 a_1740_101.n9 GND 0.08fF
C31 a_1740_101.n10 GND 0.17fF
C32 a_1740_101.t1 GND 0.23fF
C33 a_1740_101.n11 GND 0.09fF
C34 a_1740_101.n12 GND 0.00fF
C35 a_5366_101.n0 GND 0.05fF
C36 a_5366_101.n1 GND 0.12fF
C37 a_5366_101.n2 GND 0.04fF
C38 a_4383_103.n0 GND 0.10fF
C39 a_4383_103.n1 GND 0.04fF
C40 a_4383_103.n2 GND 0.03fF
C41 a_4383_103.n3 GND 0.07fF
C42 a_4383_103.n4 GND 0.08fF
C43 a_4383_103.n5 GND 0.06fF
C44 a_10990_101.n0 GND 0.05fF
C45 a_10990_101.n1 GND 0.12fF
C46 a_10990_101.n2 GND 0.04fF
C47 a_11656_101.n0 GND 0.05fF
C48 a_11656_101.n1 GND 0.12fF
C49 a_11656_101.n2 GND 0.04fF
C50 a_8956_210.n0 GND 0.02fF
C51 a_8956_210.n1 GND 0.09fF
C52 a_8956_210.n2 GND 0.13fF
C53 a_8956_210.n3 GND 0.11fF
C54 a_8956_210.t1 GND 0.30fF
C55 a_8956_210.n4 GND 0.09fF
C56 a_8956_210.n5 GND 0.06fF
C57 a_8956_210.n6 GND 0.01fF
C58 a_8956_210.n7 GND 0.03fF
C59 a_8956_210.n8 GND 0.11fF
C60 a_8956_210.n9 GND 0.02fF
C61 a_8956_210.n10 GND 0.05fF
C62 a_8956_210.n11 GND 0.02fF
C63 a_91_103.n0 GND 0.09fF
C64 a_91_103.n1 GND 0.09fF
C65 a_91_103.n2 GND 0.04fF
C66 a_91_103.n3 GND 0.03fF
C67 a_91_103.n4 GND 0.04fF
C68 a_91_103.n5 GND 0.03fF
C69 a_91_103.n6 GND 0.04fF
C70 a_6032_101.n0 GND 0.05fF
C71 a_6032_101.n1 GND 0.12fF
C72 a_6032_101.n2 GND 0.04fF
C73 a_6698_101.n0 GND 0.02fF
C74 a_6698_101.n1 GND 0.10fF
C75 a_6698_101.n2 GND 0.06fF
C76 a_6698_101.n3 GND 0.06fF
C77 a_6698_101.n4 GND 0.00fF
C78 a_6698_101.n5 GND 0.04fF
C79 a_6698_101.n6 GND 0.05fF
C80 a_6698_101.n7 GND 0.02fF
C81 a_6698_101.n8 GND 0.05fF
C82 a_6698_101.n9 GND 0.08fF
C83 a_6698_101.n10 GND 0.17fF
C84 a_6698_101.t1 GND 0.23fF
C85 a_6698_101.n11 GND 0.09fF
C86 a_6698_101.n12 GND 0.00fF
C87 a_3072_101.n0 GND 0.05fF
C88 a_3072_101.n1 GND 0.12fF
C89 a_3072_101.n2 GND 0.04fF
C90 a_4664_210.n0 GND 0.07fF
C91 a_4664_210.n1 GND 0.09fF
C92 a_4664_210.n2 GND 0.13fF
C93 a_4664_210.n3 GND 0.11fF
C94 a_4664_210.n4 GND 0.02fF
C95 a_4664_210.n5 GND 0.03fF
C96 a_4664_210.n6 GND 0.02fF
C97 a_4664_210.n7 GND 0.05fF
C98 a_4664_210.n8 GND 0.03fF
C99 a_4664_210.n9 GND 0.11fF
C100 a_4664_210.n10 GND 0.06fF
C101 a_4664_210.n11 GND 0.01fF
C102 a_4664_210.t0 GND 0.33fF
C103 a_9658_101.n0 GND 0.05fF
C104 a_9658_101.n1 GND 0.12fF
C105 a_9658_101.n2 GND 0.04fF
C106 a_11761_1050.n0 GND 0.27fF
C107 a_11761_1050.n1 GND 0.62fF
C108 a_11761_1050.n2 GND 0.04fF
C109 a_11761_1050.n3 GND 0.05fF
C110 a_11761_1050.n4 GND 0.03fF
C111 a_11761_1050.n5 GND 0.39fF
C112 a_11761_1050.n6 GND 0.56fF
C113 a_11761_1050.n7 GND 0.62fF
C114 a_11761_1050.n8 GND 0.21fF
C115 a_11761_1050.n9 GND 0.53fF
C116 a_372_210.n0 GND 0.02fF
C117 a_372_210.n1 GND 0.09fF
C118 a_372_210.n2 GND 0.13fF
C119 a_372_210.n3 GND 0.11fF
C120 a_372_210.t1 GND 0.30fF
C121 a_372_210.n4 GND 0.09fF
C122 a_372_210.n5 GND 0.06fF
C123 a_372_210.n6 GND 0.01fF
C124 a_372_210.n7 GND 0.03fF
C125 a_372_210.n8 GND 0.11fF
C126 a_372_210.n9 GND 0.02fF
C127 a_372_210.n10 GND 0.05fF
C128 a_372_210.n11 GND 0.03fF
C129 a_2406_101.n0 GND 0.02fF
C130 a_2406_101.n1 GND 0.10fF
C131 a_2406_101.n2 GND 0.06fF
C132 a_2406_101.n3 GND 0.06fF
C133 a_2406_101.n4 GND 0.00fF
C134 a_2406_101.n5 GND 0.04fF
C135 a_2406_101.n6 GND 0.05fF
C136 a_2406_101.n7 GND 0.02fF
C137 a_2406_101.n8 GND 0.05fF
C138 a_2406_101.n9 GND 0.08fF
C139 a_2406_101.n10 GND 0.17fF
C140 a_2406_101.t1 GND 0.23fF
C141 a_2406_101.n11 GND 0.09fF
C142 a_2406_101.n12 GND 0.00fF
C143 a_12322_101.n0 GND 0.05fF
C144 a_12322_101.n1 GND 0.12fF
C145 a_12322_101.n2 GND 0.04fF
C146 a_3177_1050.n0 GND 0.36fF
C147 a_3177_1050.n1 GND 0.60fF
C148 a_3177_1050.n2 GND 0.04fF
C149 a_3177_1050.n3 GND 0.06fF
C150 a_3177_1050.n4 GND 0.04fF
C151 a_3177_1050.n5 GND 0.34fF
C152 a_3177_1050.n6 GND 0.62fF
C153 a_3177_1050.n7 GND 0.65fF
C154 a_3177_1050.n8 GND 0.29fF
C155 a_3177_1050.n9 GND 0.55fF
C156 a_277_1050.n0 GND 0.72fF
C157 a_277_1050.n1 GND 0.46fF
C158 a_277_1050.n2 GND 0.64fF
C159 a_277_1050.n3 GND 0.46fF
C160 a_277_1050.n4 GND 0.54fF
C161 a_277_1050.n5 GND 2.59fF
C162 a_277_1050.n6 GND 0.05fF
C163 a_277_1050.n7 GND 0.07fF
C164 a_277_1050.n8 GND 0.05fF
C165 a_277_1050.n9 GND 0.45fF
C166 a_277_1050.n10 GND 0.61fF
C167 a_277_1050.n11 GND 0.37fF
C168 a_277_1050.n12 GND 0.85fF
C169 a_277_1050.n13 GND 0.27fF
C170 a_277_1050.n14 GND 0.72fF
C171 a_1074_101.n0 GND 0.05fF
C172 a_1074_101.n1 GND 0.12fF
C173 a_1074_101.n2 GND 0.04fF
C174 a_8030_101.n0 GND 0.05fF
C175 a_8030_101.n1 GND 0.12fF
C176 a_8030_101.n2 GND 0.04fF
C177 a_4891_989.n0 GND 0.49fF
C178 a_4891_989.n1 GND 0.52fF
C179 a_4891_989.n2 GND 0.49fF
C180 a_4891_989.t6 GND 0.69fF
C181 a_4891_989.n3 GND 0.50fF
C182 a_4891_989.n4 GND 1.33fF
C183 a_4891_989.n5 GND 0.05fF
C184 a_4891_989.n6 GND 0.07fF
C185 a_4891_989.n7 GND 0.04fF
C186 a_4891_989.n8 GND 0.39fF
C187 a_4891_989.n9 GND 0.56fF
C188 a_4891_989.n10 GND 0.82fF
C189 a_4891_989.n11 GND 0.40fF
C190 a_4891_989.n12 GND 0.69fF
C191 a_13093_1051.n0 GND 0.37fF
C192 a_13093_1051.n1 GND 0.41fF
C193 a_13093_1051.n2 GND 0.28fF
C194 a_13093_1051.n3 GND 0.63fF
C195 a_13093_1051.n4 GND 0.24fF
C196 a_13093_1051.n5 GND 0.33fF
C197 a_11887_411.n0 GND 0.28fF
C198 a_11887_411.n1 GND 0.74fF
C199 a_11887_411.n2 GND 0.25fF
C200 a_11887_411.n3 GND 0.50fF
C201 a_11887_411.n4 GND 0.37fF
C202 a_11887_411.n5 GND 0.31fF
C203 a_11887_411.t13 GND 0.56fF
C204 a_11887_411.n6 GND 0.40fF
C205 a_11887_411.n7 GND 0.96fF
C206 a_11887_411.n8 GND 0.04fF
C207 a_11887_411.n9 GND 0.05fF
C208 a_11887_411.n10 GND 0.03fF
C209 a_11887_411.n11 GND 0.33fF
C210 a_11887_411.n12 GND 0.43fF
C211 a_11887_411.n13 GND 0.63fF
C212 a_11887_411.n14 GND 0.28fF
C213 a_11887_411.n15 GND 0.53fF
C214 a_8675_103.n0 GND 0.09fF
C215 a_8675_103.n1 GND 0.10fF
C216 a_8675_103.n2 GND 0.05fF
C217 a_8675_103.n3 GND 0.03fF
C218 a_8675_103.n4 GND 0.04fF
C219 a_8675_103.n5 GND 0.11fF
C220 a_8675_103.n6 GND 0.04fF
C221 a_1845_1050.n0 GND 0.54fF
C222 a_1845_1050.n1 GND 0.39fF
C223 a_1845_1050.n2 GND 0.59fF
C224 a_1845_1050.n3 GND 0.04fF
C225 a_1845_1050.n4 GND 0.06fF
C226 a_1845_1050.n5 GND 0.04fF
C227 a_1845_1050.n6 GND 0.31fF
C228 a_1845_1050.n7 GND 0.62fF
C229 a_1845_1050.n8 GND 0.31fF
C230 a_1845_1050.n9 GND 0.64fF
C231 a_6137_1050.n0 GND 0.43fF
C232 a_6137_1050.n1 GND 0.65fF
C233 a_6137_1050.n2 GND 0.05fF
C234 a_6137_1050.n3 GND 0.06fF
C235 a_6137_1050.n4 GND 0.04fF
C236 a_6137_1050.n5 GND 0.34fF
C237 a_6137_1050.n6 GND 0.69fF
C238 a_6137_1050.n7 GND 0.71fF
C239 a_6137_1050.n8 GND 0.35fF
C240 a_6137_1050.n9 GND 0.60fF
C241 a_4439_187.n0 GND 0.45fF
C242 a_4439_187.t9 GND 0.96fF
C243 a_4439_187.n1 GND 0.66fF
C244 a_4439_187.n2 GND 0.45fF
C245 a_4439_187.t7 GND 0.96fF
C246 a_4439_187.n3 GND 0.62fF
C247 a_4439_187.n4 GND 0.44fF
C248 a_4439_187.n5 GND 0.88fF
C249 a_4439_187.n6 GND 2.85fF
C250 a_4439_187.n7 GND 2.12fF
C251 a_4439_187.n8 GND 0.07fF
C252 a_4439_187.n9 GND 0.09fF
C253 a_4439_187.n10 GND 0.06fF
C254 a_4439_187.n11 GND 0.58fF
C255 a_4439_187.n12 GND 0.69fF
C256 a_4439_187.n13 GND 1.01fF
C257 a_4439_187.n14 GND 0.40fF
C258 a_4439_187.n15 GND 0.86fF
C259 a_4569_1050.n0 GND 0.79fF
C260 a_4569_1050.n1 GND 0.51fF
C261 a_4569_1050.n2 GND 0.70fF
C262 a_4569_1050.n3 GND 0.51fF
C263 a_4569_1050.n4 GND 0.59fF
C264 a_4569_1050.n5 GND 2.84fF
C265 a_4569_1050.n6 GND 0.64fF
C266 a_4569_1050.n7 GND 0.71fF
C267 a_4569_1050.n8 GND 0.41fF
C268 a_4569_1050.n9 GND 0.93fF
C269 a_4569_1050.n10 GND 0.29fF
C270 a_4569_1050.n11 GND 0.79fF
C271 a_8861_1050.n0 GND 0.79fF
C272 a_8861_1050.n1 GND 0.79fF
C273 a_8861_1050.n2 GND 0.51fF
C274 a_8861_1050.n3 GND 0.69fF
C275 a_8861_1050.n4 GND 0.51fF
C276 a_8861_1050.n5 GND 0.59fF
C277 a_8861_1050.n6 GND 2.83fF
C278 a_8861_1050.n7 GND 0.06fF
C279 a_8861_1050.n8 GND 0.08fF
C280 a_8861_1050.n9 GND 0.05fF
C281 a_8861_1050.n10 GND 0.49fF
C282 a_8861_1050.n11 GND 0.67fF
C283 a_8861_1050.n12 GND 0.41fF
C284 a_8861_1050.n13 GND 0.29fF
C285 a_8861_1050.n14 GND 0.93fF
C286 a_9183_989.n0 GND 0.50fF
C287 a_9183_989.n1 GND 0.53fF
C288 a_9183_989.n2 GND 0.50fF
C289 a_9183_989.t9 GND 0.71fF
C290 a_9183_989.n3 GND 0.51fF
C291 a_9183_989.n4 GND 1.36fF
C292 a_9183_989.n5 GND 0.05fF
C293 a_9183_989.n6 GND 0.07fF
C294 a_9183_989.n7 GND 0.05fF
C295 a_9183_989.n8 GND 0.40fF
C296 a_9183_989.n9 GND 0.57fF
C297 a_9183_989.n10 GND 0.84fF
C298 a_9183_989.n11 GND 0.41fF
C299 a_9183_989.n12 GND 0.71fF
C300 a_10324_101.n0 GND 0.02fF
C301 a_10324_101.n1 GND 0.10fF
C302 a_10324_101.n2 GND 0.06fF
C303 a_10324_101.n3 GND 0.06fF
C304 a_10324_101.n4 GND 0.00fF
C305 a_10324_101.n5 GND 0.04fF
C306 a_10324_101.n6 GND 0.05fF
C307 a_10324_101.n7 GND 0.02fF
C308 a_10324_101.n8 GND 0.05fF
C309 a_10324_101.n9 GND 0.08fF
C310 a_10324_101.n10 GND 0.17fF
C311 a_10324_101.t1 GND 0.23fF
C312 a_10324_101.n11 GND 0.09fF
C313 a_10324_101.n12 GND 0.00fF
C314 a_7469_1050.n0 GND 0.37fF
C315 a_7469_1050.n1 GND 0.61fF
C316 a_7469_1050.n2 GND 0.46fF
C317 a_7469_1050.n3 GND 0.67fF
C318 a_7469_1050.n4 GND 0.67fF
C319 a_7469_1050.n5 GND 0.29fF
C320 a_7469_1050.n6 GND 0.56fF
C321 a_7364_101.n0 GND 0.08fF
C322 a_7364_101.n1 GND 0.02fF
C323 a_7364_101.n2 GND 0.01fF
C324 a_7364_101.n3 GND 0.06fF
C325 a_7364_101.n4 GND 0.10fF
C326 a_7364_101.n5 GND 0.06fF
C327 a_7364_101.n6 GND 0.05fF
C328 a_3738_101.n0 GND 0.02fF
C329 a_3738_101.n1 GND 0.10fF
C330 a_3738_101.n2 GND 0.06fF
C331 a_3738_101.n3 GND 0.06fF
C332 a_3738_101.n4 GND 0.00fF
C333 a_3738_101.n5 GND 0.04fF
C334 a_3738_101.n6 GND 0.05fF
C335 a_3738_101.n7 GND 0.02fF
C336 a_3738_101.n8 GND 0.05fF
C337 a_3738_101.n9 GND 0.08fF
C338 a_3738_101.n10 GND 0.17fF
C339 a_3738_101.t1 GND 0.23fF
C340 a_3738_101.n11 GND 0.09fF
C341 a_3738_101.n12 GND 0.00fF
C342 a_147_187.n0 GND 0.79fF
C343 a_147_187.n1 GND 0.93fF
C344 a_147_187.n2 GND 0.36fF
C345 a_147_187.n3 GND 0.41fF
C346 a_147_187.t5 GND 0.88fF
C347 a_147_187.n4 GND 0.61fF
C348 a_147_187.n5 GND 0.41fF
C349 a_147_187.t13 GND 0.88fF
C350 a_147_187.n6 GND 0.57fF
C351 a_147_187.n7 GND 0.41fF
C352 a_147_187.n8 GND 0.81fF
C353 a_147_187.n9 GND 2.62fF
C354 a_147_187.n10 GND 1.95fF
C355 a_147_187.n11 GND 0.64fF
C356 a_147_187.n12 GND 0.12fF
C357 a_147_187.n13 GND 0.52fF
C358 a_147_187.n14 GND 0.07fF
C359 QN.n0 GND 0.42fF
C360 QN.n1 GND 0.51fF
C361 QN.n2 GND 0.25fF
C362 QN.n3 GND 0.04fF
C363 QN.n4 GND 0.05fF
C364 QN.n5 GND 0.03fF
C365 QN.n6 GND 0.09fF
C366 QN.n7 GND 0.04fF
C367 QN.n8 GND 0.05fF
C368 QN.n9 GND 0.03fF
C369 QN.n10 GND 0.10fF
C370 QN.n11 GND 1.06fF
C371 QN.n12 GND 0.13fF
C372 QN.n13 GND 0.32fF
C373 QN.n14 GND 0.37fF
C374 QN.n15 GND 0.01fF
C375 a_13757_1051.n0 GND 0.35fF
C376 a_13757_1051.n1 GND 0.29fF
C377 a_13757_1051.n2 GND 0.20fF
C378 a_13757_1051.n3 GND 0.56fF
C379 a_13757_1051.n4 GND 0.25fF
C380 a_13757_1051.n5 GND 0.28fF
C381 a_7595_411.n0 GND 0.69fF
C382 a_7595_411.n1 GND 0.81fF
C383 a_7595_411.n2 GND 0.52fF
C384 a_7595_411.n3 GND 0.36fF
C385 a_7595_411.n4 GND 0.40fF
C386 a_7595_411.n5 GND 1.26fF
C387 a_7595_411.n6 GND 1.02fF
C388 a_7595_411.n7 GND 0.88fF
C389 a_7595_411.n8 GND 0.55fF
C390 a_7595_411.t6 GND 0.59fF
C391 a_7595_411.n9 GND 0.50fF
C392 a_7595_411.n10 GND 5.53fF
C393 a_7595_411.n11 GND 0.57fF
C394 a_7595_411.n12 GND 0.11fF
C395 a_7595_411.n13 GND 0.25fF
C396 a_7595_411.n14 GND 0.06fF
C397 a_8731_187.n0 GND 0.84fF
C398 a_8731_187.n1 GND 0.44fF
C399 a_8731_187.t9 GND 0.94fF
C400 a_8731_187.n2 GND 0.65fF
C401 a_8731_187.n3 GND 0.44fF
C402 a_8731_187.t6 GND 0.94fF
C403 a_8731_187.n4 GND 0.61fF
C404 a_8731_187.n5 GND 0.43fF
C405 a_8731_187.n6 GND 0.86fF
C406 a_8731_187.n7 GND 2.79fF
C407 a_8731_187.n8 GND 2.08fF
C408 a_8731_187.n9 GND 0.73fF
C409 a_8731_187.n10 GND 0.72fF
C410 a_8731_187.n11 GND 0.39fF
C411 a_8731_187.n12 GND 0.99fF
C412 a_10429_1050.n0 GND 0.60fF
C413 a_10429_1050.n1 GND 0.71fF
C414 a_10429_1050.n2 GND 0.35fF
C415 a_10429_1050.n3 GND 0.43fF
C416 a_10429_1050.n4 GND 0.65fF
C417 a_10429_1050.n5 GND 0.69fF
C418 a_10429_1050.n6 GND 0.09fF
C419 a_10429_1050.n7 GND 0.33fF
C420 a_10429_1050.n8 GND 0.05fF
C421 a_14320_101.n0 GND 0.06fF
C422 a_14320_101.n1 GND 0.03fF
C423 a_14320_101.n2 GND 0.13fF
C424 a_14320_101.n3 GND 0.04fF
C425 a_14320_101.n4 GND 0.18fF
C426 a_3303_411.n0 GND 0.81fF
C427 a_3303_411.n1 GND 0.96fF
C428 a_3303_411.n2 GND 0.52fF
C429 a_3303_411.n3 GND 0.58fF
C430 a_3303_411.n4 GND 0.73fF
C431 a_3303_411.n5 GND 0.89fF
C432 a_3303_411.n6 GND 0.56fF
C433 a_3303_411.n7 GND 2.50fF
C434 a_3303_411.n8 GND 0.56fF
C435 a_3303_411.t6 GND 0.78fF
C436 a_3303_411.n9 GND 0.60fF
C437 a_3303_411.n10 GND 11.50fF
C438 a_3303_411.n11 GND 0.67fF
C439 a_3303_411.n12 GND 0.13fF
C440 a_3303_411.n13 GND 0.40fF
C441 a_3303_411.n14 GND 0.07fF
C442 a_599_989.n0 GND 0.40fF
C443 a_599_989.n1 GND 0.43fF
C444 a_599_989.n2 GND 0.40fF
C445 a_599_989.t6 GND 0.57fF
C446 a_599_989.n3 GND 0.41fF
C447 a_599_989.n4 GND 1.09fF
C448 a_599_989.n5 GND 0.04fF
C449 a_599_989.n6 GND 0.06fF
C450 a_599_989.n7 GND 0.04fF
C451 a_599_989.n8 GND 0.32fF
C452 a_599_989.n9 GND 0.46fF
C453 a_599_989.n10 GND 0.67fF
C454 a_599_989.n11 GND 0.33fF
C455 a_599_989.n12 GND 0.57fF
C456 VDD.n0 GND 0.16fF
C457 VDD.n1 GND 0.03fF
C458 VDD.n2 GND 0.02fF
C459 VDD.n3 GND 0.05fF
C460 VDD.n4 GND 0.01fF
C461 VDD.n5 GND 0.02fF
C462 VDD.n6 GND 0.02fF
C463 VDD.n8 GND 0.02fF
C464 VDD.n9 GND 0.02fF
C465 VDD.n12 GND 0.02fF
C466 VDD.n14 GND 0.47fF
C467 VDD.n16 GND 0.03fF
C468 VDD.n17 GND 0.02fF
C469 VDD.n18 GND 0.02fF
C470 VDD.n19 GND 0.02fF
C471 VDD.n20 GND 0.04fF
C472 VDD.n21 GND 0.28fF
C473 VDD.n22 GND 0.02fF
C474 VDD.n23 GND 0.03fF
C475 VDD.n24 GND 0.28fF
C476 VDD.n25 GND 0.01fF
C477 VDD.n26 GND 0.32fF
C478 VDD.n27 GND 0.01fF
C479 VDD.n28 GND 0.03fF
C480 VDD.n29 GND 0.02fF
C481 VDD.n30 GND 0.28fF
C482 VDD.n31 GND 0.01fF
C483 VDD.n32 GND 0.02fF
C484 VDD.n33 GND 0.00fF
C485 VDD.n34 GND 0.09fF
C486 VDD.n35 GND 0.03fF
C487 VDD.n36 GND 0.32fF
C488 VDD.n37 GND 0.01fF
C489 VDD.n38 GND 0.03fF
C490 VDD.n39 GND 0.03fF
C491 VDD.n40 GND 0.28fF
C492 VDD.n41 GND 0.01fF
C493 VDD.n42 GND 0.02fF
C494 VDD.n43 GND 0.02fF
C495 VDD.n44 GND 0.28fF
C496 VDD.n45 GND 0.01fF
C497 VDD.n46 GND 0.02fF
C498 VDD.n47 GND 0.02fF
C499 VDD.n48 GND 0.28fF
C500 VDD.n49 GND 0.01fF
C501 VDD.n50 GND 0.02fF
C502 VDD.n51 GND 0.04fF
C503 VDD.n52 GND 0.02fF
C504 VDD.n53 GND 0.02fF
C505 VDD.n54 GND 0.02fF
C506 VDD.n55 GND 0.22fF
C507 VDD.n56 GND 0.04fF
C508 VDD.n57 GND 0.04fF
C509 VDD.n58 GND 0.02fF
C510 VDD.n60 GND 0.02fF
C511 VDD.n61 GND 0.02fF
C512 VDD.n62 GND 0.02fF
C513 VDD.n63 GND 0.02fF
C514 VDD.n65 GND 0.02fF
C515 VDD.n66 GND 0.02fF
C516 VDD.n67 GND 0.02fF
C517 VDD.n69 GND 0.28fF
C518 VDD.n71 GND 0.02fF
C519 VDD.n72 GND 0.02fF
C520 VDD.n73 GND 0.03fF
C521 VDD.n74 GND 0.02fF
C522 VDD.n75 GND 0.28fF
C523 VDD.n76 GND 0.01fF
C524 VDD.n77 GND 0.02fF
C525 VDD.n78 GND 0.04fF
C526 VDD.n79 GND 0.28fF
C527 VDD.n80 GND 0.01fF
C528 VDD.n81 GND 0.02fF
C529 VDD.n82 GND 0.02fF
C530 VDD.n83 GND 0.28fF
C531 VDD.n84 GND 0.01fF
C532 VDD.n85 GND 0.02fF
C533 VDD.n86 GND 0.02fF
C534 VDD.n87 GND 0.32fF
C535 VDD.n88 GND 0.01fF
C536 VDD.n89 GND 0.03fF
C537 VDD.n90 GND 0.03fF
C538 VDD.n91 GND 0.32fF
C539 VDD.n92 GND 0.01fF
C540 VDD.n93 GND 0.03fF
C541 VDD.n94 GND 0.03fF
C542 VDD.n95 GND 0.28fF
C543 VDD.n96 GND 0.01fF
C544 VDD.n97 GND 0.02fF
C545 VDD.n98 GND 0.02fF
C546 VDD.n99 GND 0.28fF
C547 VDD.n100 GND 0.01fF
C548 VDD.n101 GND 0.02fF
C549 VDD.n102 GND 0.02fF
C550 VDD.n103 GND 0.28fF
C551 VDD.n104 GND 0.01fF
C552 VDD.n105 GND 0.02fF
C553 VDD.n106 GND 0.04fF
C554 VDD.n107 GND 0.02fF
C555 VDD.n108 GND 0.02fF
C556 VDD.n109 GND 0.02fF
C557 VDD.n110 GND 0.22fF
C558 VDD.n111 GND 0.04fF
C559 VDD.n112 GND 0.03fF
C560 VDD.n113 GND 0.02fF
C561 VDD.n114 GND 0.02fF
C562 VDD.n115 GND 0.02fF
C563 VDD.n116 GND 0.03fF
C564 VDD.n117 GND 0.02fF
C565 VDD.n119 GND 0.02fF
C566 VDD.n120 GND 0.02fF
C567 VDD.n121 GND 0.02fF
C568 VDD.n123 GND 0.28fF
C569 VDD.n125 GND 0.02fF
C570 VDD.n126 GND 0.02fF
C571 VDD.n127 GND 0.03fF
C572 VDD.n128 GND 0.02fF
C573 VDD.n129 GND 0.28fF
C574 VDD.n130 GND 0.01fF
C575 VDD.n131 GND 0.02fF
C576 VDD.n132 GND 0.04fF
C577 VDD.n133 GND 0.06fF
C578 VDD.n134 GND 0.25fF
C579 VDD.n135 GND 0.01fF
C580 VDD.n136 GND 0.01fF
C581 VDD.n137 GND 0.02fF
C582 VDD.n138 GND 0.14fF
C583 VDD.n139 GND 0.17fF
C584 VDD.n140 GND 0.01fF
C585 VDD.n141 GND 0.02fF
C586 VDD.n142 GND 0.02fF
C587 VDD.n143 GND 0.11fF
C588 VDD.n144 GND 0.03fF
C589 VDD.n145 GND 0.31fF
C590 VDD.n146 GND 0.01fF
C591 VDD.n147 GND 0.02fF
C592 VDD.n148 GND 0.03fF
C593 VDD.n149 GND 0.18fF
C594 VDD.n150 GND 0.14fF
C595 VDD.n151 GND 0.01fF
C596 VDD.n152 GND 0.02fF
C597 VDD.n153 GND 0.03fF
C598 VDD.n154 GND 0.14fF
C599 VDD.n155 GND 0.17fF
C600 VDD.n156 GND 0.01fF
C601 VDD.n157 GND 0.02fF
C602 VDD.n158 GND 0.02fF
C603 VDD.n159 GND 0.06fF
C604 VDD.n160 GND 0.25fF
C605 VDD.n161 GND 0.01fF
C606 VDD.n162 GND 0.01fF
C607 VDD.n163 GND 0.02fF
C608 VDD.n164 GND 0.28fF
C609 VDD.n165 GND 0.01fF
C610 VDD.n166 GND 0.02fF
C611 VDD.n167 GND 0.04fF
C612 VDD.n168 GND 0.02fF
C613 VDD.n169 GND 0.02fF
C614 VDD.n170 GND 0.02fF
C615 VDD.n171 GND 0.22fF
C616 VDD.n172 GND 0.04fF
C617 VDD.n173 GND 0.03fF
C618 VDD.n174 GND 0.02fF
C619 VDD.n175 GND 0.02fF
C620 VDD.n176 GND 0.02fF
C621 VDD.n177 GND 0.03fF
C622 VDD.n178 GND 0.02fF
C623 VDD.n180 GND 0.02fF
C624 VDD.n181 GND 0.02fF
C625 VDD.n182 GND 0.02fF
C626 VDD.n184 GND 0.28fF
C627 VDD.n186 GND 0.02fF
C628 VDD.n187 GND 0.02fF
C629 VDD.n188 GND 0.03fF
C630 VDD.n189 GND 0.02fF
C631 VDD.n190 GND 0.28fF
C632 VDD.n191 GND 0.01fF
C633 VDD.n192 GND 0.02fF
C634 VDD.n193 GND 0.04fF
C635 VDD.n194 GND 0.06fF
C636 VDD.n195 GND 0.25fF
C637 VDD.n196 GND 0.01fF
C638 VDD.n197 GND 0.01fF
C639 VDD.n198 GND 0.02fF
C640 VDD.n199 GND 0.14fF
C641 VDD.n200 GND 0.17fF
C642 VDD.n201 GND 0.01fF
C643 VDD.n202 GND 0.02fF
C644 VDD.n203 GND 0.02fF
C645 VDD.n204 GND 0.11fF
C646 VDD.n205 GND 0.03fF
C647 VDD.n206 GND 0.31fF
C648 VDD.n207 GND 0.01fF
C649 VDD.n208 GND 0.02fF
C650 VDD.n209 GND 0.03fF
C651 VDD.n210 GND 0.18fF
C652 VDD.n211 GND 0.14fF
C653 VDD.n212 GND 0.01fF
C654 VDD.n213 GND 0.02fF
C655 VDD.n214 GND 0.03fF
C656 VDD.n215 GND 0.14fF
C657 VDD.n216 GND 0.17fF
C658 VDD.n217 GND 0.01fF
C659 VDD.n218 GND 0.02fF
C660 VDD.n219 GND 0.02fF
C661 VDD.n220 GND 0.06fF
C662 VDD.n221 GND 0.25fF
C663 VDD.n222 GND 0.01fF
C664 VDD.n223 GND 0.01fF
C665 VDD.n224 GND 0.02fF
C666 VDD.n225 GND 0.28fF
C667 VDD.n226 GND 0.01fF
C668 VDD.n227 GND 0.02fF
C669 VDD.n228 GND 0.04fF
C670 VDD.n229 GND 0.02fF
C671 VDD.n230 GND 0.02fF
C672 VDD.n231 GND 0.02fF
C673 VDD.n232 GND 0.22fF
C674 VDD.n233 GND 0.04fF
C675 VDD.n234 GND 0.03fF
C676 VDD.n235 GND 0.02fF
C677 VDD.n236 GND 0.02fF
C678 VDD.n237 GND 0.02fF
C679 VDD.n238 GND 0.03fF
C680 VDD.n239 GND 0.02fF
C681 VDD.n241 GND 0.02fF
C682 VDD.n242 GND 0.02fF
C683 VDD.n243 GND 0.02fF
C684 VDD.n245 GND 0.28fF
C685 VDD.n247 GND 0.02fF
C686 VDD.n248 GND 0.02fF
C687 VDD.n249 GND 0.03fF
C688 VDD.n250 GND 0.02fF
C689 VDD.n251 GND 0.28fF
C690 VDD.n252 GND 0.01fF
C691 VDD.n253 GND 0.02fF
C692 VDD.n254 GND 0.04fF
C693 VDD.n255 GND 0.06fF
C694 VDD.n256 GND 0.25fF
C695 VDD.n257 GND 0.01fF
C696 VDD.n258 GND 0.01fF
C697 VDD.n259 GND 0.02fF
C698 VDD.n260 GND 0.14fF
C699 VDD.n261 GND 0.17fF
C700 VDD.n262 GND 0.01fF
C701 VDD.n263 GND 0.02fF
C702 VDD.n264 GND 0.02fF
C703 VDD.n265 GND 0.11fF
C704 VDD.n266 GND 0.03fF
C705 VDD.n267 GND 0.31fF
C706 VDD.n268 GND 0.01fF
C707 VDD.n269 GND 0.02fF
C708 VDD.n270 GND 0.03fF
C709 VDD.n271 GND 0.18fF
C710 VDD.n272 GND 0.14fF
C711 VDD.n273 GND 0.01fF
C712 VDD.n274 GND 0.02fF
C713 VDD.n275 GND 0.03fF
C714 VDD.n276 GND 0.14fF
C715 VDD.n277 GND 0.17fF
C716 VDD.n278 GND 0.01fF
C717 VDD.n279 GND 0.02fF
C718 VDD.n280 GND 0.02fF
C719 VDD.n281 GND 0.06fF
C720 VDD.n282 GND 0.25fF
C721 VDD.n283 GND 0.01fF
C722 VDD.n284 GND 0.01fF
C723 VDD.n285 GND 0.02fF
C724 VDD.n286 GND 0.28fF
C725 VDD.n287 GND 0.01fF
C726 VDD.n288 GND 0.02fF
C727 VDD.n289 GND 0.04fF
C728 VDD.n290 GND 0.02fF
C729 VDD.n291 GND 0.02fF
C730 VDD.n292 GND 0.02fF
C731 VDD.n293 GND 0.22fF
C732 VDD.n294 GND 0.04fF
C733 VDD.n295 GND 0.03fF
C734 VDD.n296 GND 0.02fF
C735 VDD.n297 GND 0.02fF
C736 VDD.n298 GND 0.02fF
C737 VDD.n299 GND 0.03fF
C738 VDD.n300 GND 0.02fF
C739 VDD.n302 GND 0.02fF
C740 VDD.n303 GND 0.02fF
C741 VDD.n304 GND 0.02fF
C742 VDD.n306 GND 0.28fF
C743 VDD.n308 GND 0.02fF
C744 VDD.n309 GND 0.02fF
C745 VDD.n310 GND 0.03fF
C746 VDD.n311 GND 0.02fF
C747 VDD.n312 GND 0.28fF
C748 VDD.n313 GND 0.01fF
C749 VDD.n314 GND 0.02fF
C750 VDD.n315 GND 0.04fF
C751 VDD.n316 GND 0.06fF
C752 VDD.n317 GND 0.25fF
C753 VDD.n318 GND 0.01fF
C754 VDD.n319 GND 0.01fF
C755 VDD.n320 GND 0.02fF
C756 VDD.n321 GND 0.14fF
C757 VDD.n322 GND 0.17fF
C758 VDD.n323 GND 0.01fF
C759 VDD.n324 GND 0.02fF
C760 VDD.n325 GND 0.02fF
C761 VDD.n326 GND 0.11fF
C762 VDD.n327 GND 0.03fF
C763 VDD.n328 GND 0.31fF
C764 VDD.n329 GND 0.01fF
C765 VDD.n330 GND 0.02fF
C766 VDD.n331 GND 0.03fF
C767 VDD.n332 GND 0.18fF
C768 VDD.n333 GND 0.14fF
C769 VDD.n334 GND 0.01fF
C770 VDD.n335 GND 0.02fF
C771 VDD.n336 GND 0.03fF
C772 VDD.n337 GND 0.14fF
C773 VDD.n338 GND 0.17fF
C774 VDD.n339 GND 0.01fF
C775 VDD.n340 GND 0.02fF
C776 VDD.n341 GND 0.02fF
C777 VDD.n342 GND 0.06fF
C778 VDD.n343 GND 0.25fF
C779 VDD.n344 GND 0.01fF
C780 VDD.n345 GND 0.01fF
C781 VDD.n346 GND 0.02fF
C782 VDD.n347 GND 0.28fF
C783 VDD.n348 GND 0.01fF
C784 VDD.n349 GND 0.02fF
C785 VDD.n350 GND 0.04fF
C786 VDD.n351 GND 0.02fF
C787 VDD.n352 GND 0.02fF
C788 VDD.n353 GND 0.02fF
C789 VDD.n354 GND 0.22fF
C790 VDD.n355 GND 0.04fF
C791 VDD.n356 GND 0.03fF
C792 VDD.n357 GND 0.02fF
C793 VDD.n358 GND 0.02fF
C794 VDD.n359 GND 0.02fF
C795 VDD.n360 GND 0.03fF
C796 VDD.n361 GND 0.02fF
C797 VDD.n363 GND 0.02fF
C798 VDD.n364 GND 0.02fF
C799 VDD.n365 GND 0.02fF
C800 VDD.n367 GND 0.28fF
C801 VDD.n369 GND 0.02fF
C802 VDD.n370 GND 0.02fF
C803 VDD.n371 GND 0.03fF
C804 VDD.n372 GND 0.02fF
C805 VDD.n373 GND 0.28fF
C806 VDD.n374 GND 0.01fF
C807 VDD.n375 GND 0.02fF
C808 VDD.n376 GND 0.04fF
C809 VDD.n377 GND 0.06fF
C810 VDD.n378 GND 0.25fF
C811 VDD.n379 GND 0.01fF
C812 VDD.n380 GND 0.01fF
C813 VDD.n381 GND 0.02fF
C814 VDD.n382 GND 0.14fF
C815 VDD.n383 GND 0.17fF
C816 VDD.n384 GND 0.01fF
C817 VDD.n385 GND 0.02fF
C818 VDD.n386 GND 0.02fF
C819 VDD.n387 GND 0.11fF
C820 VDD.n388 GND 0.03fF
C821 VDD.n389 GND 0.31fF
C822 VDD.n390 GND 0.01fF
C823 VDD.n391 GND 0.02fF
C824 VDD.n392 GND 0.03fF
C825 VDD.n393 GND 0.18fF
C826 VDD.n394 GND 0.14fF
C827 VDD.n395 GND 0.01fF
C828 VDD.n396 GND 0.02fF
C829 VDD.n397 GND 0.03fF
C830 VDD.n398 GND 0.14fF
C831 VDD.n399 GND 0.17fF
C832 VDD.n400 GND 0.01fF
C833 VDD.n401 GND 0.02fF
C834 VDD.n402 GND 0.02fF
C835 VDD.n403 GND 0.06fF
C836 VDD.n404 GND 0.25fF
C837 VDD.n405 GND 0.01fF
C838 VDD.n406 GND 0.01fF
C839 VDD.n407 GND 0.02fF
C840 VDD.n408 GND 0.28fF
C841 VDD.n409 GND 0.01fF
C842 VDD.n410 GND 0.02fF
C843 VDD.n411 GND 0.04fF
C844 VDD.n412 GND 0.02fF
C845 VDD.n413 GND 0.02fF
C846 VDD.n414 GND 0.02fF
C847 VDD.n415 GND 0.22fF
C848 VDD.n416 GND 0.04fF
C849 VDD.n417 GND 0.03fF
C850 VDD.n418 GND 0.02fF
C851 VDD.n419 GND 0.02fF
C852 VDD.n420 GND 0.02fF
C853 VDD.n421 GND 0.03fF
C854 VDD.n422 GND 0.02fF
C855 VDD.n424 GND 0.02fF
C856 VDD.n425 GND 0.02fF
C857 VDD.n426 GND 0.02fF
C858 VDD.n428 GND 0.28fF
C859 VDD.n430 GND 0.02fF
C860 VDD.n431 GND 0.02fF
C861 VDD.n432 GND 0.03fF
C862 VDD.n433 GND 0.02fF
C863 VDD.n434 GND 0.28fF
C864 VDD.n435 GND 0.01fF
C865 VDD.n436 GND 0.02fF
C866 VDD.n437 GND 0.04fF
C867 VDD.n438 GND 0.06fF
C868 VDD.n439 GND 0.25fF
C869 VDD.n440 GND 0.01fF
C870 VDD.n441 GND 0.01fF
C871 VDD.n442 GND 0.02fF
C872 VDD.n443 GND 0.14fF
C873 VDD.n444 GND 0.17fF
C874 VDD.n445 GND 0.01fF
C875 VDD.n446 GND 0.02fF
C876 VDD.n447 GND 0.02fF
C877 VDD.n448 GND 0.11fF
C878 VDD.n449 GND 0.03fF
C879 VDD.n450 GND 0.31fF
C880 VDD.n451 GND 0.01fF
C881 VDD.n452 GND 0.02fF
C882 VDD.n453 GND 0.03fF
C883 VDD.n454 GND 0.18fF
C884 VDD.n455 GND 0.14fF
C885 VDD.n456 GND 0.01fF
C886 VDD.n457 GND 0.02fF
C887 VDD.n458 GND 0.03fF
C888 VDD.n459 GND 0.14fF
C889 VDD.n460 GND 0.17fF
C890 VDD.n461 GND 0.01fF
C891 VDD.n462 GND 0.02fF
C892 VDD.n463 GND 0.02fF
C893 VDD.n464 GND 0.06fF
C894 VDD.n465 GND 0.25fF
C895 VDD.n466 GND 0.01fF
C896 VDD.n467 GND 0.01fF
C897 VDD.n468 GND 0.02fF
C898 VDD.n469 GND 0.28fF
C899 VDD.n470 GND 0.01fF
C900 VDD.n471 GND 0.02fF
C901 VDD.n472 GND 0.04fF
C902 VDD.n473 GND 0.02fF
C903 VDD.n474 GND 0.02fF
C904 VDD.n475 GND 0.02fF
C905 VDD.n476 GND 0.27fF
C906 VDD.n477 GND 0.04fF
C907 VDD.n478 GND 0.03fF
C908 VDD.n479 GND 0.02fF
C909 VDD.n480 GND 0.02fF
C910 VDD.n481 GND 0.02fF
C911 VDD.n482 GND 0.03fF
C912 VDD.n483 GND 0.02fF
C913 VDD.n485 GND 0.02fF
C914 VDD.n486 GND 0.02fF
C915 VDD.n487 GND 0.02fF
C916 VDD.n489 GND 0.28fF
C917 VDD.n491 GND 0.02fF
C918 VDD.n492 GND 0.02fF
C919 VDD.n493 GND 0.03fF
C920 VDD.n494 GND 0.02fF
C921 VDD.n495 GND 0.28fF
C922 VDD.n496 GND 0.01fF
C923 VDD.n497 GND 0.02fF
C924 VDD.n498 GND 0.04fF
C925 VDD.n499 GND 0.28fF
C926 VDD.n500 GND 0.01fF
C927 VDD.n501 GND 0.02fF
C928 VDD.n502 GND 0.02fF
C929 VDD.n503 GND 0.23fF
C930 VDD.n504 GND 0.01fF
C931 VDD.n505 GND 0.07fF
C932 VDD.n506 GND 0.02fF
C933 VDD.n507 GND 0.14fF
C934 VDD.n508 GND 0.17fF
C935 VDD.n509 GND 0.01fF
C936 VDD.n510 GND 0.02fF
C937 VDD.n511 GND 0.02fF
C938 VDD.n512 GND 0.14fF
C939 VDD.n513 GND 0.16fF
C940 VDD.n514 GND 0.01fF
C941 VDD.n515 GND 0.11fF
C942 VDD.n516 GND 0.02fF
C943 VDD.n517 GND 0.02fF
C944 VDD.n518 GND 0.02fF
C945 VDD.n519 GND 0.18fF
C946 VDD.n520 GND 0.15fF
C947 VDD.n521 GND 0.02fF
C948 VDD.n522 GND 0.02fF
C949 VDD.n523 GND 0.03fF
C950 VDD.n524 GND 0.18fF
C951 VDD.n525 GND 0.15fF
C952 VDD.n526 GND 0.02fF
C953 VDD.n527 GND 0.02fF
C954 VDD.n528 GND 0.03fF
C955 VDD.n529 GND 0.11fF
C956 VDD.n530 GND 0.02fF
C957 VDD.n531 GND 0.14fF
C958 VDD.n532 GND 0.16fF
C959 VDD.n533 GND 0.01fF
C960 VDD.n534 GND 0.02fF
C961 VDD.n535 GND 0.02fF
C962 VDD.n536 GND 0.14fF
C963 VDD.n537 GND 0.17fF
C964 VDD.n538 GND 0.01fF
C965 VDD.n539 GND 0.02fF
C966 VDD.n540 GND 0.02fF
C967 VDD.n541 GND 0.06fF
C968 VDD.n542 GND 0.23fF
C969 VDD.n543 GND 0.01fF
C970 VDD.n544 GND 0.01fF
C971 VDD.n545 GND 0.02fF
C972 VDD.n546 GND 0.28fF
C973 VDD.n547 GND 0.01fF
C974 VDD.n548 GND 0.02fF
C975 VDD.n549 GND 0.02fF
C976 VDD.n550 GND 0.28fF
C977 VDD.n551 GND 0.01fF
C978 VDD.n552 GND 0.02fF
C979 VDD.n553 GND 0.04fF
C980 VDD.n554 GND 0.02fF
C981 VDD.n555 GND 0.02fF
C982 VDD.n556 GND 0.02fF
C983 VDD.n557 GND 0.27fF
C984 VDD.n558 GND 0.04fF
C985 VDD.n559 GND 0.03fF
C986 VDD.n560 GND 0.02fF
C987 VDD.n561 GND 0.02fF
C988 VDD.n562 GND 0.02fF
C989 VDD.n563 GND 0.03fF
C990 VDD.n564 GND 0.02fF
C991 VDD.n566 GND 0.02fF
C992 VDD.n567 GND 0.02fF
C993 VDD.n568 GND 0.02fF
C994 VDD.n570 GND 0.28fF
C995 VDD.n572 GND 0.02fF
C996 VDD.n573 GND 0.02fF
C997 VDD.n574 GND 0.03fF
C998 VDD.n575 GND 0.02fF
C999 VDD.n576 GND 0.28fF
C1000 VDD.n577 GND 0.01fF
C1001 VDD.n578 GND 0.02fF
C1002 VDD.n579 GND 0.04fF
C1003 VDD.n580 GND 0.06fF
C1004 VDD.n581 GND 0.25fF
C1005 VDD.n582 GND 0.01fF
C1006 VDD.n583 GND 0.01fF
C1007 VDD.n584 GND 0.02fF
C1008 VDD.n585 GND 0.14fF
C1009 VDD.n586 GND 0.17fF
C1010 VDD.n587 GND 0.01fF
C1011 VDD.n588 GND 0.02fF
C1012 VDD.n589 GND 0.02fF
C1013 VDD.n590 GND 0.11fF
C1014 VDD.n591 GND 0.03fF
C1015 VDD.n592 GND 0.31fF
C1016 VDD.n593 GND 0.01fF
C1017 VDD.n594 GND 0.02fF
C1018 VDD.n595 GND 0.03fF
C1019 VDD.n596 GND 0.18fF
C1020 VDD.n597 GND 0.14fF
C1021 VDD.n598 GND 0.01fF
C1022 VDD.n599 GND 0.02fF
C1023 VDD.n600 GND 0.03fF
C1024 VDD.n601 GND 0.14fF
C1025 VDD.n602 GND 0.17fF
C1026 VDD.n603 GND 0.01fF
C1027 VDD.n604 GND 0.02fF
C1028 VDD.n605 GND 0.02fF
C1029 VDD.n606 GND 0.06fF
C1030 VDD.n607 GND 0.25fF
C1031 VDD.n608 GND 0.01fF
C1032 VDD.n609 GND 0.01fF
C1033 VDD.n610 GND 0.02fF
C1034 VDD.n611 GND 0.28fF
C1035 VDD.n612 GND 0.01fF
C1036 VDD.n613 GND 0.02fF
C1037 VDD.n614 GND 0.04fF
C1038 VDD.n615 GND 0.02fF
C1039 VDD.n616 GND 0.02fF
C1040 VDD.n617 GND 0.02fF
C1041 VDD.n618 GND 0.22fF
C1042 VDD.n619 GND 0.04fF
C1043 VDD.n620 GND 0.03fF
C1044 VDD.n621 GND 0.02fF
C1045 VDD.n622 GND 0.02fF
C1046 VDD.n623 GND 0.02fF
C1047 VDD.n624 GND 0.03fF
C1048 VDD.n625 GND 0.02fF
C1049 VDD.n627 GND 0.02fF
C1050 VDD.n628 GND 0.02fF
C1051 VDD.n629 GND 0.02fF
C1052 VDD.n631 GND 0.28fF
C1053 VDD.n633 GND 0.02fF
C1054 VDD.n634 GND 0.02fF
C1055 VDD.n635 GND 0.03fF
C1056 VDD.n636 GND 0.02fF
C1057 VDD.n637 GND 0.28fF
C1058 VDD.n638 GND 0.01fF
C1059 VDD.n639 GND 0.02fF
C1060 VDD.n640 GND 0.04fF
C1061 VDD.n641 GND 0.06fF
C1062 VDD.n642 GND 0.25fF
C1063 VDD.n643 GND 0.01fF
C1064 VDD.n644 GND 0.01fF
C1065 VDD.n645 GND 0.02fF
C1066 VDD.n646 GND 0.14fF
C1067 VDD.n647 GND 0.17fF
C1068 VDD.n648 GND 0.01fF
C1069 VDD.n649 GND 0.02fF
C1070 VDD.n650 GND 0.02fF
C1071 VDD.n651 GND 0.11fF
C1072 VDD.n652 GND 0.03fF
C1073 VDD.n653 GND 0.31fF
C1074 VDD.n654 GND 0.01fF
C1075 VDD.n655 GND 0.02fF
C1076 VDD.n656 GND 0.03fF
C1077 VDD.n657 GND 0.18fF
C1078 VDD.n658 GND 0.14fF
C1079 VDD.n659 GND 0.01fF
C1080 VDD.n660 GND 0.02fF
C1081 VDD.n661 GND 0.03fF
C1082 VDD.n662 GND 0.14fF
C1083 VDD.n663 GND 0.17fF
C1084 VDD.n664 GND 0.01fF
C1085 VDD.n665 GND 0.02fF
C1086 VDD.n666 GND 0.02fF
C1087 VDD.n667 GND 0.02fF
C1088 VDD.n668 GND 0.02fF
C1089 VDD.n669 GND 0.02fF
C1090 VDD.n670 GND 0.21fF
C1091 VDD.n671 GND 0.03fF
C1092 VDD.n672 GND 0.02fF
C1093 VDD.n673 GND 0.02fF
C1094 VDD.n674 GND 0.02fF
C1095 VDD.n675 GND 0.03fF
C1096 VDD.n676 GND 0.02fF
C1097 VDD.n678 GND 0.02fF
C1098 VDD.n679 GND 0.02fF
C1099 VDD.n680 GND 0.02fF
C1100 VDD.n682 GND 0.47fF
C1101 VDD.n684 GND 0.03fF
C1102 VDD.n685 GND 0.04fF
C1103 VDD.n686 GND 0.28fF
C1104 VDD.n687 GND 0.02fF
C1105 VDD.n688 GND 0.03fF
C1106 VDD.n689 GND 0.03fF
C1107 VDD.n690 GND 0.28fF
C1108 VDD.n691 GND 0.01fF
C1109 VDD.n692 GND 0.02fF
C1110 VDD.n693 GND 0.02fF
C1111 VDD.n694 GND 0.06fF
C1112 VDD.n695 GND 0.23fF
C1113 VDD.n696 GND 0.01fF
C1114 VDD.n697 GND 0.01fF
C1115 VDD.n698 GND 0.02fF
C1116 VDD.n699 GND 0.14fF
C1117 VDD.n700 GND 0.17fF
C1118 VDD.n701 GND 0.01fF
C1119 VDD.n702 GND 0.02fF
C1120 VDD.n703 GND 0.02fF
C1121 VDD.n704 GND 0.11fF
C1122 VDD.n705 GND 0.02fF
C1123 VDD.n706 GND 0.14fF
C1124 VDD.n707 GND 0.16fF
C1125 VDD.n708 GND 0.01fF
C1126 VDD.n709 GND 0.02fF
C1127 VDD.n710 GND 0.02fF
C1128 VDD.n711 GND 0.18fF
C1129 VDD.n712 GND 0.15fF
C1130 VDD.n713 GND 0.02fF
C1131 VDD.n714 GND 0.02fF
C1132 VDD.n715 GND 0.03fF
C1133 VDD.n716 GND 0.18fF
C1134 VDD.n717 GND 0.15fF
C1135 VDD.n718 GND 0.02fF
C1136 VDD.n719 GND 0.02fF
C1137 VDD.n720 GND 0.03fF
C1138 VDD.n721 GND 0.14fF
C1139 VDD.n722 GND 0.16fF
C1140 VDD.n723 GND 0.01fF
C1141 VDD.n724 GND 0.11fF
C1142 VDD.n725 GND 0.02fF
C1143 VDD.n726 GND 0.02fF
C1144 VDD.n727 GND 0.02fF
C1145 VDD.n728 GND 0.14fF
C1146 VDD.n729 GND 0.17fF
C1147 VDD.n730 GND 0.01fF
C1148 VDD.n731 GND 0.02fF
C1149 VDD.n732 GND 0.02fF
C1150 VDD.n733 GND 0.23fF
C1151 VDD.n734 GND 0.01fF
C1152 VDD.n735 GND 0.07fF
C1153 VDD.n736 GND 0.02fF
C1154 VDD.n737 GND 0.28fF
C1155 VDD.n738 GND 0.01fF
C1156 VDD.n739 GND 0.02fF
C1157 VDD.n740 GND 0.02fF
C1158 VDD.n741 GND 0.28fF
C1159 VDD.n742 GND 0.01fF
C1160 VDD.n743 GND 0.02fF
C1161 VDD.n744 GND 0.04fF
C1162 VDD.n745 GND 0.02fF
C1163 VDD.n746 GND 0.02fF
C1164 VDD.n747 GND 0.02fF
C1165 VDD.n748 GND 0.02fF
C1166 VDD.n749 GND 0.02fF
C1167 VDD.n750 GND 0.02fF
C1168 VDD.n752 GND 0.02fF
C1169 VDD.n753 GND 0.02fF
C1170 VDD.n754 GND 0.02fF
C1171 VDD.n755 GND 0.02fF
C1172 VDD.n757 GND 0.04fF
C1173 VDD.n758 GND 0.02fF
C1174 VDD.n759 GND 0.27fF
C1175 VDD.n760 GND 0.04fF
C1176 VDD.n762 GND 0.28fF
C1177 VDD.n764 GND 0.02fF
C1178 VDD.n765 GND 0.02fF
C1179 VDD.n766 GND 0.03fF
C1180 VDD.n767 GND 0.02fF
C1181 VDD.n768 GND 0.28fF
C1182 VDD.n769 GND 0.01fF
C1183 VDD.n770 GND 0.02fF
C1184 VDD.n771 GND 0.04fF
C1185 VDD.n772 GND 0.06fF
C1186 VDD.n773 GND 0.25fF
C1187 VDD.n774 GND 0.01fF
C1188 VDD.n775 GND 0.01fF
C1189 VDD.n776 GND 0.02fF
C1190 VDD.n777 GND 0.14fF
C1191 VDD.n778 GND 0.17fF
C1192 VDD.n779 GND 0.01fF
C1193 VDD.n780 GND 0.02fF
C1194 VDD.n781 GND 0.02fF
C1195 VDD.n782 GND 0.18fF
C1196 VDD.n783 GND 0.14fF
C1197 VDD.n784 GND 0.01fF
C1198 VDD.n785 GND 0.02fF
C1199 VDD.n786 GND 0.03fF
C1200 VDD.n787 GND 0.11fF
C1201 VDD.n788 GND 0.03fF
C1202 VDD.n789 GND 0.31fF
C1203 VDD.n790 GND 0.01fF
C1204 VDD.n791 GND 0.02fF
C1205 VDD.n792 GND 0.03fF
C1206 VDD.n793 GND 0.14fF
C1207 VDD.n794 GND 0.17fF
C1208 VDD.n795 GND 0.01fF
C1209 VDD.n796 GND 0.02fF
C1210 VDD.n797 GND 0.02fF
C1211 VDD.n798 GND 0.06fF
C1212 VDD.n799 GND 0.25fF
C1213 VDD.n800 GND 0.01fF
C1214 VDD.n801 GND 0.01fF
C1215 VDD.n802 GND 0.02fF
C1216 VDD.n803 GND 0.28fF
C1217 VDD.n804 GND 0.01fF
C1218 VDD.n805 GND 0.02fF
C1219 VDD.n806 GND 0.04fF
C1220 VDD.n807 GND 0.02fF
C1221 VDD.n808 GND 0.02fF
C1222 VDD.n809 GND 0.02fF
C1223 VDD.n810 GND 0.22fF
C1224 VDD.n811 GND 0.04fF
C1225 VDD.n812 GND 0.03fF
C1226 VDD.n813 GND 0.02fF
C1227 VDD.n814 GND 0.02fF
C1228 VDD.n815 GND 0.02fF
C1229 VDD.n816 GND 0.03fF
C1230 VDD.n817 GND 0.02fF
C1231 VDD.n819 GND 0.02fF
C1232 VDD.n820 GND 0.02fF
C1233 VDD.n821 GND 0.02fF
C1234 VDD.n823 GND 0.28fF
C1235 VDD.n825 GND 0.02fF
C1236 VDD.n826 GND 0.02fF
C1237 VDD.n827 GND 0.03fF
C1238 VDD.n828 GND 0.02fF
C1239 VDD.n829 GND 0.28fF
C1240 VDD.n830 GND 0.01fF
C1241 VDD.n831 GND 0.02fF
C1242 VDD.n832 GND 0.04fF
C1243 VDD.n833 GND 0.06fF
C1244 VDD.n834 GND 0.25fF
C1245 VDD.n835 GND 0.01fF
C1246 VDD.n836 GND 0.01fF
C1247 VDD.n837 GND 0.02fF
C1248 VDD.n838 GND 0.14fF
C1249 VDD.n839 GND 0.17fF
C1250 VDD.n840 GND 0.01fF
C1251 VDD.n841 GND 0.02fF
C1252 VDD.n842 GND 0.02fF
C1253 VDD.n843 GND 0.18fF
C1254 VDD.n844 GND 0.14fF
C1255 VDD.n845 GND 0.01fF
C1256 VDD.n846 GND 0.02fF
C1257 VDD.n847 GND 0.03fF
C1258 VDD.n848 GND 0.11fF
C1259 VDD.n849 GND 0.03fF
C1260 VDD.n850 GND 0.31fF
C1261 VDD.n851 GND 0.01fF
C1262 VDD.n852 GND 0.02fF
C1263 VDD.n853 GND 0.03fF
C1264 VDD.n854 GND 0.14fF
C1265 VDD.n855 GND 0.17fF
C1266 VDD.n856 GND 0.01fF
C1267 VDD.n857 GND 0.02fF
C1268 VDD.n858 GND 0.02fF
C1269 VDD.n859 GND 0.06fF
C1270 VDD.n860 GND 0.25fF
C1271 VDD.n861 GND 0.01fF
C1272 VDD.n862 GND 0.01fF
C1273 VDD.n863 GND 0.02fF
C1274 VDD.n864 GND 0.28fF
C1275 VDD.n865 GND 0.01fF
C1276 VDD.n866 GND 0.02fF
C1277 VDD.n867 GND 0.04fF
C1278 VDD.n868 GND 0.02fF
C1279 VDD.n869 GND 0.02fF
C1280 VDD.n870 GND 0.02fF
C1281 VDD.n871 GND 0.22fF
C1282 VDD.n872 GND 0.04fF
C1283 VDD.n873 GND 0.03fF
C1284 VDD.n874 GND 0.02fF
C1285 VDD.n875 GND 0.02fF
C1286 VDD.n876 GND 0.02fF
C1287 VDD.n877 GND 0.03fF
C1288 VDD.n878 GND 0.02fF
C1289 VDD.n880 GND 0.02fF
C1290 VDD.n881 GND 0.02fF
C1291 VDD.n882 GND 0.02fF
C1292 VDD.n884 GND 0.28fF
C1293 VDD.n886 GND 0.02fF
C1294 VDD.n887 GND 0.02fF
C1295 VDD.n888 GND 0.03fF
C1296 VDD.n889 GND 0.02fF
C1297 VDD.n890 GND 0.28fF
C1298 VDD.n891 GND 0.01fF
C1299 VDD.n892 GND 0.02fF
C1300 VDD.n893 GND 0.04fF
C1301 VDD.n894 GND 0.06fF
C1302 VDD.n895 GND 0.25fF
C1303 VDD.n896 GND 0.01fF
C1304 VDD.n897 GND 0.01fF
C1305 VDD.n898 GND 0.02fF
C1306 VDD.n899 GND 0.14fF
C1307 VDD.n900 GND 0.17fF
C1308 VDD.n901 GND 0.01fF
C1309 VDD.n902 GND 0.02fF
C1310 VDD.n903 GND 0.02fF
C1311 VDD.n904 GND 0.18fF
C1312 VDD.n905 GND 0.14fF
C1313 VDD.n906 GND 0.01fF
C1314 VDD.n907 GND 0.02fF
C1315 VDD.n908 GND 0.03fF
C1316 VDD.n909 GND 0.11fF
C1317 VDD.n910 GND 0.03fF
C1318 VDD.n911 GND 0.31fF
C1319 VDD.n912 GND 0.01fF
C1320 VDD.n913 GND 0.02fF
C1321 VDD.n914 GND 0.03fF
C1322 VDD.n915 GND 0.14fF
C1323 VDD.n916 GND 0.17fF
C1324 VDD.n917 GND 0.01fF
C1325 VDD.n918 GND 0.02fF
C1326 VDD.n919 GND 0.02fF
C1327 VDD.n920 GND 0.06fF
C1328 VDD.n921 GND 0.25fF
C1329 VDD.n922 GND 0.01fF
C1330 VDD.n923 GND 0.01fF
C1331 VDD.n924 GND 0.02fF
C1332 VDD.n925 GND 0.28fF
C1333 VDD.n926 GND 0.01fF
C1334 VDD.n927 GND 0.02fF
C1335 VDD.n928 GND 0.04fF
C1336 VDD.n929 GND 0.02fF
C1337 VDD.n930 GND 0.02fF
C1338 VDD.n931 GND 0.02fF
C1339 VDD.n932 GND 0.22fF
C1340 VDD.n933 GND 0.04fF
C1341 VDD.n934 GND 0.03fF
C1342 VDD.n935 GND 0.02fF
C1343 VDD.n936 GND 0.02fF
C1344 VDD.n937 GND 0.02fF
C1345 VDD.n938 GND 0.03fF
C1346 VDD.n939 GND 0.02fF
C1347 VDD.n941 GND 0.02fF
C1348 VDD.n942 GND 0.02fF
C1349 VDD.n943 GND 0.02fF
C1350 VDD.n945 GND 0.28fF
C1351 VDD.n947 GND 0.02fF
C1352 VDD.n948 GND 0.02fF
C1353 VDD.n949 GND 0.03fF
C1354 VDD.n950 GND 0.02fF
C1355 VDD.n951 GND 0.28fF
C1356 VDD.n952 GND 0.01fF
C1357 VDD.n953 GND 0.02fF
C1358 VDD.n954 GND 0.04fF
C1359 VDD.n955 GND 0.06fF
C1360 VDD.n956 GND 0.25fF
C1361 VDD.n957 GND 0.01fF
C1362 VDD.n958 GND 0.01fF
C1363 VDD.n959 GND 0.02fF
C1364 VDD.n960 GND 0.14fF
C1365 VDD.n961 GND 0.17fF
C1366 VDD.n962 GND 0.01fF
C1367 VDD.n963 GND 0.02fF
C1368 VDD.n964 GND 0.02fF
C1369 VDD.n965 GND 0.18fF
C1370 VDD.n966 GND 0.14fF
C1371 VDD.n967 GND 0.01fF
C1372 VDD.n968 GND 0.02fF
C1373 VDD.n969 GND 0.03fF
C1374 VDD.n970 GND 0.11fF
C1375 VDD.n971 GND 0.03fF
C1376 VDD.n972 GND 0.31fF
C1377 VDD.n973 GND 0.01fF
C1378 VDD.n974 GND 0.02fF
C1379 VDD.n975 GND 0.03fF
C1380 VDD.n976 GND 0.14fF
C1381 VDD.n977 GND 0.17fF
C1382 VDD.n978 GND 0.01fF
C1383 VDD.n979 GND 0.02fF
C1384 VDD.n980 GND 0.02fF
C1385 VDD.n981 GND 0.06fF
C1386 VDD.n982 GND 0.25fF
C1387 VDD.n983 GND 0.01fF
C1388 VDD.n984 GND 0.01fF
C1389 VDD.n985 GND 0.02fF
C1390 VDD.n986 GND 0.28fF
C1391 VDD.n987 GND 0.01fF
C1392 VDD.n988 GND 0.02fF
C1393 VDD.n989 GND 0.04fF
C1394 VDD.n990 GND 0.02fF
C1395 VDD.n991 GND 0.02fF
C1396 VDD.n992 GND 0.02fF
C1397 VDD.n993 GND 0.22fF
C1398 VDD.n994 GND 0.04fF
C1399 VDD.n995 GND 0.03fF
C1400 VDD.n996 GND 0.02fF
C1401 VDD.n997 GND 0.02fF
C1402 VDD.n998 GND 0.02fF
C1403 VDD.n999 GND 0.03fF
C1404 VDD.n1000 GND 0.02fF
C1405 VDD.n1002 GND 0.02fF
C1406 VDD.n1003 GND 0.02fF
C1407 VDD.n1004 GND 0.02fF
C1408 VDD.n1006 GND 0.28fF
C1409 VDD.n1008 GND 0.02fF
C1410 VDD.n1009 GND 0.02fF
C1411 VDD.n1010 GND 0.03fF
C1412 VDD.n1011 GND 0.02fF
C1413 VDD.n1012 GND 0.28fF
C1414 VDD.n1013 GND 0.01fF
C1415 VDD.n1014 GND 0.02fF
C1416 VDD.n1015 GND 0.04fF
C1417 VDD.n1016 GND 0.06fF
C1418 VDD.n1017 GND 0.25fF
C1419 VDD.n1018 GND 0.01fF
C1420 VDD.n1019 GND 0.01fF
C1421 VDD.n1020 GND 0.02fF
C1422 VDD.n1021 GND 0.14fF
C1423 VDD.n1022 GND 0.17fF
C1424 VDD.n1023 GND 0.01fF
C1425 VDD.n1024 GND 0.02fF
C1426 VDD.n1025 GND 0.02fF
C1427 VDD.n1026 GND 0.18fF
C1428 VDD.n1027 GND 0.14fF
C1429 VDD.n1028 GND 0.01fF
C1430 VDD.n1029 GND 0.02fF
C1431 VDD.n1030 GND 0.03fF
C1432 VDD.n1031 GND 0.11fF
C1433 VDD.n1032 GND 0.03fF
C1434 VDD.n1033 GND 0.31fF
C1435 VDD.n1034 GND 0.01fF
C1436 VDD.n1035 GND 0.02fF
C1437 VDD.n1036 GND 0.03fF
C1438 VDD.n1037 GND 0.14fF
C1439 VDD.n1038 GND 0.17fF
C1440 VDD.n1039 GND 0.01fF
C1441 VDD.n1040 GND 0.02fF
C1442 VDD.n1041 GND 0.02fF
C1443 VDD.n1042 GND 0.06fF
C1444 VDD.n1043 GND 0.25fF
C1445 VDD.n1044 GND 0.01fF
C1446 VDD.n1045 GND 0.01fF
C1447 VDD.n1046 GND 0.02fF
C1448 VDD.n1047 GND 0.28fF
C1449 VDD.n1048 GND 0.01fF
C1450 VDD.n1049 GND 0.02fF
C1451 VDD.n1050 GND 0.04fF
C1452 VDD.n1051 GND 0.02fF
C1453 VDD.n1052 GND 0.02fF
C1454 VDD.n1053 GND 0.02fF
C1455 VDD.n1054 GND 0.27fF
C1456 VDD.n1055 GND 0.04fF
C1457 VDD.n1056 GND 0.03fF
C1458 VDD.n1057 GND 0.02fF
C1459 VDD.n1058 GND 0.02fF
C1460 VDD.n1059 GND 0.02fF
C1461 VDD.n1060 GND 0.03fF
C1462 VDD.n1061 GND 0.02fF
C1463 VDD.n1063 GND 0.02fF
C1464 VDD.n1064 GND 0.02fF
C1465 VDD.n1065 GND 0.02fF
C1466 VDD.n1067 GND 0.28fF
C1467 VDD.n1069 GND 0.02fF
C1468 VDD.n1070 GND 0.02fF
C1469 VDD.n1071 GND 0.03fF
C1470 VDD.n1072 GND 0.02fF
C1471 VDD.n1073 GND 0.28fF
C1472 VDD.n1074 GND 0.01fF
C1473 VDD.n1075 GND 0.02fF
C1474 VDD.n1076 GND 0.04fF
C1475 VDD.n1077 GND 0.28fF
C1476 VDD.n1078 GND 0.01fF
C1477 VDD.n1079 GND 0.02fF
C1478 VDD.n1080 GND 0.02fF
C1479 VDD.n1081 GND 0.06fF
C1480 VDD.n1082 GND 0.23fF
C1481 VDD.n1083 GND 0.01fF
C1482 VDD.n1084 GND 0.01fF
C1483 VDD.n1085 GND 0.02fF
C1484 VDD.n1086 GND 0.14fF
C1485 VDD.n1087 GND 0.17fF
C1486 VDD.n1088 GND 0.01fF
C1487 VDD.n1089 GND 0.02fF
C1488 VDD.n1090 GND 0.02fF
C1489 VDD.n1091 GND 0.11fF
C1490 VDD.n1092 GND 0.02fF
C1491 VDD.n1093 GND 0.14fF
C1492 VDD.n1094 GND 0.16fF
C1493 VDD.n1095 GND 0.01fF
C1494 VDD.n1096 GND 0.02fF
C1495 VDD.n1097 GND 0.02fF
C1496 VDD.n1098 GND 0.18fF
C1497 VDD.n1099 GND 0.15fF
C1498 VDD.n1100 GND 0.02fF
C1499 VDD.n1101 GND 0.02fF
C1500 VDD.n1102 GND 0.03fF
C1501 VDD.n1103 GND 0.18fF
C1502 VDD.n1104 GND 0.15fF
C1503 VDD.n1105 GND 0.02fF
C1504 VDD.n1106 GND 0.02fF
C1505 VDD.n1107 GND 0.03fF
C1506 VDD.n1108 GND 0.14fF
C1507 VDD.n1109 GND 0.16fF
C1508 VDD.n1110 GND 0.01fF
C1509 VDD.n1111 GND 0.11fF
C1510 VDD.n1112 GND 0.02fF
C1511 VDD.n1113 GND 0.02fF
C1512 VDD.n1114 GND 0.02fF
C1513 VDD.n1115 GND 0.14fF
C1514 VDD.n1116 GND 0.17fF
C1515 VDD.n1117 GND 0.01fF
C1516 VDD.n1118 GND 0.02fF
C1517 VDD.n1119 GND 0.02fF
C1518 VDD.n1120 GND 0.23fF
C1519 VDD.n1121 GND 0.01fF
C1520 VDD.n1122 GND 0.07fF
C1521 VDD.n1123 GND 0.02fF
C1522 VDD.n1124 GND 0.28fF
C1523 VDD.n1125 GND 0.01fF
C1524 VDD.n1126 GND 0.02fF
C1525 VDD.n1127 GND 0.02fF
C1526 VDD.n1128 GND 0.28fF
C1527 VDD.n1129 GND 0.01fF
C1528 VDD.n1130 GND 0.02fF
C1529 VDD.n1131 GND 0.04fF
C1530 VDD.n1132 GND 0.02fF
C1531 VDD.n1133 GND 0.02fF
C1532 VDD.n1134 GND 0.02fF
C1533 VDD.n1135 GND 0.27fF
C1534 VDD.n1136 GND 0.04fF
C1535 VDD.n1137 GND 0.03fF
C1536 VDD.n1138 GND 0.02fF
C1537 VDD.n1139 GND 0.02fF
C1538 VDD.n1140 GND 0.02fF
C1539 VDD.n1141 GND 0.03fF
C1540 VDD.n1142 GND 0.02fF
C1541 VDD.n1144 GND 0.02fF
C1542 VDD.n1145 GND 0.02fF
C1543 VDD.n1146 GND 0.02fF
C1544 VDD.n1148 GND 0.28fF
C1545 VDD.n1150 GND 0.02fF
C1546 VDD.n1151 GND 0.02fF
C1547 VDD.n1152 GND 0.03fF
C1548 VDD.n1153 GND 0.02fF
C1549 VDD.n1154 GND 0.28fF
C1550 VDD.n1155 GND 0.01fF
C1551 VDD.n1156 GND 0.02fF
C1552 VDD.n1157 GND 0.04fF
C1553 VDD.n1158 GND 0.06fF
C1554 VDD.n1159 GND 0.25fF
C1555 VDD.n1160 GND 0.01fF
C1556 VDD.n1161 GND 0.01fF
C1557 VDD.n1162 GND 0.02fF
C1558 VDD.n1163 GND 0.14fF
C1559 VDD.n1164 GND 0.17fF
C1560 VDD.n1165 GND 0.01fF
C1561 VDD.n1166 GND 0.02fF
C1562 VDD.n1167 GND 0.02fF
C1563 VDD.n1168 GND 0.18fF
C1564 VDD.n1169 GND 0.14fF
C1565 VDD.n1170 GND 0.01fF
C1566 VDD.n1171 GND 0.02fF
C1567 VDD.n1172 GND 0.03fF
C1568 VDD.n1173 GND 0.11fF
C1569 VDD.n1174 GND 0.03fF
C1570 VDD.n1175 GND 0.31fF
C1571 VDD.n1176 GND 0.01fF
C1572 VDD.n1177 GND 0.02fF
C1573 VDD.n1178 GND 0.03fF
C1574 VDD.n1179 GND 0.14fF
C1575 VDD.n1180 GND 0.17fF
C1576 VDD.n1181 GND 0.01fF
C1577 VDD.n1182 GND 0.02fF
C1578 VDD.n1183 GND 0.02fF
C1579 VDD.n1184 GND 0.06fF
C1580 VDD.n1185 GND 0.25fF
C1581 VDD.n1186 GND 0.01fF
C1582 VDD.n1187 GND 0.01fF
C1583 VDD.n1188 GND 0.02fF
C1584 VDD.n1189 GND 0.28fF
C1585 VDD.n1190 GND 0.01fF
C1586 VDD.n1191 GND 0.02fF
C1587 VDD.n1192 GND 0.04fF
C1588 VDD.n1193 GND 0.02fF
C1589 VDD.n1194 GND 0.02fF
C1590 VDD.n1195 GND 0.02fF
C1591 VDD.n1196 GND 0.22fF
C1592 VDD.n1197 GND 0.04fF
C1593 VDD.n1198 GND 0.03fF
C1594 VDD.n1199 GND 0.02fF
C1595 VDD.n1200 GND 0.02fF
C1596 VDD.n1201 GND 0.02fF
C1597 VDD.n1202 GND 0.03fF
C1598 VDD.n1203 GND 0.02fF
C1599 VDD.n1205 GND 0.02fF
C1600 VDD.n1206 GND 0.02fF
C1601 VDD.n1207 GND 0.02fF
C1602 VDD.n1209 GND 0.28fF
C1603 VDD.n1211 GND 0.02fF
C1604 VDD.n1212 GND 0.02fF
C1605 VDD.n1213 GND 0.03fF
C1606 VDD.n1214 GND 0.02fF
C1607 VDD.n1215 GND 0.28fF
C1608 VDD.n1216 GND 0.01fF
C1609 VDD.n1217 GND 0.02fF
C1610 VDD.n1218 GND 0.04fF
C1611 VDD.n1219 GND 0.06fF
C1612 VDD.n1220 GND 0.25fF
C1613 VDD.n1221 GND 0.01fF
C1614 VDD.n1222 GND 0.01fF
C1615 VDD.n1223 GND 0.02fF
C1616 VDD.n1224 GND 0.14fF
C1617 VDD.n1225 GND 0.17fF
C1618 VDD.n1226 GND 0.01fF
C1619 VDD.n1227 GND 0.02fF
C1620 VDD.n1228 GND 0.02fF
C1621 VDD.n1229 GND 0.18fF
C1622 VDD.n1230 GND 0.14fF
C1623 VDD.n1231 GND 0.01fF
C1624 VDD.n1232 GND 0.02fF
C1625 VDD.n1233 GND 0.03fF
C1626 VDD.n1234 GND 0.11fF
C1627 VDD.n1235 GND 0.03fF
C1628 VDD.n1236 GND 0.31fF
C1629 VDD.n1237 GND 0.01fF
C1630 VDD.n1238 GND 0.02fF
C1631 VDD.n1239 GND 0.03fF
C1632 VDD.n1240 GND 0.14fF
C1633 VDD.n1241 GND 0.17fF
C1634 VDD.n1242 GND 0.01fF
C1635 VDD.n1243 GND 0.02fF
C1636 VDD.n1244 GND 0.02fF
C1637 VDD.n1245 GND 0.06fF
C1638 VDD.n1246 GND 0.25fF
C1639 VDD.n1247 GND 0.01fF
C1640 VDD.n1248 GND 0.01fF
C1641 VDD.n1249 GND 0.02fF
C1642 VDD.n1250 GND 0.28fF
C1643 VDD.n1251 GND 0.01fF
C1644 VDD.n1252 GND 0.02fF
C1645 VDD.n1253 GND 0.04fF
C1646 VDD.n1254 GND 0.02fF
C1647 VDD.n1255 GND 0.02fF
C1648 VDD.n1256 GND 0.02fF
C1649 VDD.n1257 GND 0.22fF
C1650 VDD.n1258 GND 0.04fF
C1651 VDD.n1259 GND 0.03fF
C1652 VDD.n1260 GND 0.02fF
C1653 VDD.n1261 GND 0.02fF
C1654 VDD.n1262 GND 0.02fF
C1655 VDD.n1263 GND 0.03fF
C1656 VDD.n1264 GND 0.02fF
C1657 VDD.n1266 GND 0.02fF
C1658 VDD.n1267 GND 0.02fF
C1659 VDD.n1268 GND 0.02fF
C1660 VDD.n1270 GND 0.28fF
C1661 VDD.n1272 GND 0.02fF
C1662 VDD.n1273 GND 0.02fF
C1663 VDD.n1274 GND 0.03fF
C1664 VDD.n1275 GND 0.02fF
C1665 VDD.n1276 GND 0.28fF
C1666 VDD.n1277 GND 0.01fF
C1667 VDD.n1278 GND 0.02fF
C1668 VDD.n1279 GND 0.04fF
C1669 VDD.n1280 GND 0.06fF
C1670 VDD.n1281 GND 0.25fF
C1671 VDD.n1282 GND 0.01fF
C1672 VDD.n1283 GND 0.01fF
C1673 VDD.n1284 GND 0.02fF
C1674 VDD.n1285 GND 0.14fF
C1675 VDD.n1286 GND 0.17fF
C1676 VDD.n1287 GND 0.01fF
C1677 VDD.n1288 GND 0.02fF
C1678 VDD.n1289 GND 0.02fF
C1679 VDD.n1290 GND 0.18fF
C1680 VDD.n1291 GND 0.14fF
C1681 VDD.n1292 GND 0.01fF
C1682 VDD.n1293 GND 0.02fF
C1683 VDD.n1294 GND 0.03fF
C1684 VDD.n1295 GND 0.11fF
C1685 VDD.n1296 GND 0.03fF
C1686 VDD.n1297 GND 0.31fF
C1687 VDD.n1298 GND 0.01fF
C1688 VDD.n1299 GND 0.02fF
C1689 VDD.n1300 GND 0.03fF
C1690 VDD.n1301 GND 0.14fF
C1691 VDD.n1302 GND 0.17fF
C1692 VDD.n1303 GND 0.01fF
C1693 VDD.n1304 GND 0.02fF
C1694 VDD.n1305 GND 0.02fF
C1695 VDD.n1306 GND 0.06fF
C1696 VDD.n1307 GND 0.25fF
C1697 VDD.n1308 GND 0.01fF
C1698 VDD.n1309 GND 0.01fF
C1699 VDD.n1310 GND 0.02fF
C1700 VDD.n1311 GND 0.28fF
C1701 VDD.n1312 GND 0.01fF
C1702 VDD.n1313 GND 0.02fF
C1703 VDD.n1314 GND 0.04fF
C1704 VDD.n1315 GND 0.02fF
C1705 VDD.n1316 GND 0.02fF
C1706 VDD.n1317 GND 0.02fF
C1707 VDD.n1318 GND 0.22fF
C1708 VDD.n1319 GND 0.04fF
C1709 VDD.n1320 GND 0.03fF
C1710 VDD.n1321 GND 0.02fF
C1711 VDD.n1322 GND 0.02fF
C1712 VDD.n1323 GND 0.02fF
C1713 VDD.n1324 GND 0.03fF
C1714 VDD.n1325 GND 0.02fF
C1715 VDD.n1327 GND 0.02fF
C1716 VDD.n1328 GND 0.02fF
C1717 VDD.n1329 GND 0.02fF
C1718 VDD.n1331 GND 0.28fF
C1719 VDD.n1333 GND 0.02fF
C1720 VDD.n1334 GND 0.02fF
C1721 VDD.n1335 GND 0.03fF
C1722 VDD.n1336 GND 0.02fF
C1723 VDD.n1337 GND 0.28fF
C1724 VDD.n1338 GND 0.01fF
C1725 VDD.n1339 GND 0.02fF
C1726 VDD.n1340 GND 0.04fF
C1727 VDD.n1341 GND 0.06fF
C1728 VDD.n1342 GND 0.25fF
C1729 VDD.n1343 GND 0.01fF
C1730 VDD.n1344 GND 0.01fF
C1731 VDD.n1345 GND 0.02fF
.ends
