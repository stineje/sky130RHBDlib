magic
tech sky130A
magscale 1 2
timestamp 1670281673
<< nwell >>
rect -87 786 14961 1550
<< pwell >>
rect -34 -34 14908 544
<< nmos >>
rect 147 290 177 351
tri 177 290 193 306 sw
rect 447 290 477 351
rect 147 260 253 290
tri 253 260 283 290 sw
rect 147 159 177 260
tri 177 244 193 260 nw
tri 237 244 253 260 ne
tri 177 159 193 175 sw
tri 237 159 253 175 se
rect 253 159 283 260
tri 342 260 372 290 se
rect 372 260 477 290
rect 342 166 372 260
tri 372 244 388 260 nw
tri 431 244 447 260 ne
tri 372 166 388 182 sw
tri 431 166 447 182 se
rect 447 166 477 260
tri 147 129 177 159 ne
rect 177 129 253 159
tri 253 129 283 159 nw
tri 342 136 372 166 ne
rect 372 136 447 166
tri 447 136 477 166 nw
rect 649 298 679 351
tri 679 298 695 314 sw
rect 649 268 755 298
tri 755 268 785 298 sw
rect 649 167 679 268
tri 679 252 695 268 nw
tri 739 252 755 268 ne
tri 679 167 695 183 sw
tri 739 167 755 183 se
rect 755 167 785 268
tri 649 137 679 167 ne
rect 679 137 755 167
tri 755 137 785 167 nw
rect 1130 288 1160 349
tri 1160 288 1176 304 sw
rect 1324 296 1354 349
tri 1354 296 1370 312 sw
rect 1130 258 1236 288
tri 1236 258 1266 288 sw
rect 1324 266 1430 296
tri 1430 266 1460 296 sw
rect 1130 157 1160 258
tri 1160 242 1176 258 nw
tri 1220 242 1236 258 ne
tri 1160 157 1176 173 sw
tri 1220 157 1236 173 se
rect 1236 157 1266 258
rect 1324 165 1354 266
tri 1354 250 1370 266 nw
tri 1414 250 1430 266 ne
tri 1354 165 1370 181 sw
tri 1414 165 1430 181 se
rect 1430 165 1460 266
tri 1130 127 1160 157 ne
rect 1160 127 1236 157
tri 1236 127 1266 157 nw
tri 1324 135 1354 165 ne
rect 1354 135 1430 165
tri 1430 135 1460 165 nw
rect 1796 288 1826 349
tri 1826 288 1842 304 sw
rect 1990 296 2020 349
tri 2020 296 2036 312 sw
rect 1796 258 1902 288
tri 1902 258 1932 288 sw
rect 1990 266 2096 296
tri 2096 266 2126 296 sw
rect 1796 157 1826 258
tri 1826 242 1842 258 nw
tri 1886 242 1902 258 ne
tri 1826 157 1842 173 sw
tri 1886 157 1902 173 se
rect 1902 157 1932 258
rect 1990 165 2020 266
tri 2020 250 2036 266 nw
tri 2080 250 2096 266 ne
tri 2020 165 2036 181 sw
tri 2080 165 2096 181 se
rect 2096 165 2126 266
tri 1796 127 1826 157 ne
rect 1826 127 1902 157
tri 1902 127 1932 157 nw
tri 1990 135 2020 165 ne
rect 2020 135 2096 165
tri 2096 135 2126 165 nw
rect 2462 288 2492 349
tri 2492 288 2508 304 sw
rect 2656 296 2686 349
tri 2686 296 2702 312 sw
rect 2462 258 2568 288
tri 2568 258 2598 288 sw
rect 2656 266 2762 296
tri 2762 266 2792 296 sw
rect 2462 157 2492 258
tri 2492 242 2508 258 nw
tri 2552 242 2568 258 ne
tri 2492 157 2508 173 sw
tri 2552 157 2568 173 se
rect 2568 157 2598 258
rect 2656 165 2686 266
tri 2686 250 2702 266 nw
tri 2746 250 2762 266 ne
tri 2686 165 2702 181 sw
tri 2746 165 2762 181 se
rect 2762 165 2792 266
tri 2462 127 2492 157 ne
rect 2492 127 2568 157
tri 2568 127 2598 157 nw
tri 2656 135 2686 165 ne
rect 2686 135 2762 165
tri 2762 135 2792 165 nw
rect 3128 288 3158 349
tri 3158 288 3174 304 sw
rect 3322 296 3352 349
tri 3352 296 3368 312 sw
rect 3128 258 3234 288
tri 3234 258 3264 288 sw
rect 3322 266 3428 296
tri 3428 266 3458 296 sw
rect 3128 157 3158 258
tri 3158 242 3174 258 nw
tri 3218 242 3234 258 ne
tri 3158 157 3174 173 sw
tri 3218 157 3234 173 se
rect 3234 157 3264 258
rect 3322 165 3352 266
tri 3352 250 3368 266 nw
tri 3412 250 3428 266 ne
tri 3352 165 3368 181 sw
tri 3412 165 3428 181 se
rect 3428 165 3458 266
tri 3128 127 3158 157 ne
rect 3158 127 3234 157
tri 3234 127 3264 157 nw
tri 3322 135 3352 165 ne
rect 3352 135 3428 165
tri 3428 135 3458 165 nw
rect 3794 288 3824 349
tri 3824 288 3840 304 sw
rect 3988 296 4018 349
tri 4018 296 4034 312 sw
rect 3794 258 3900 288
tri 3900 258 3930 288 sw
rect 3988 266 4094 296
tri 4094 266 4124 296 sw
rect 3794 157 3824 258
tri 3824 242 3840 258 nw
tri 3884 242 3900 258 ne
tri 3824 157 3840 173 sw
tri 3884 157 3900 173 se
rect 3900 157 3930 258
rect 3988 165 4018 266
tri 4018 250 4034 266 nw
tri 4078 250 4094 266 ne
tri 4018 165 4034 181 sw
tri 4078 165 4094 181 se
rect 4094 165 4124 266
tri 3794 127 3824 157 ne
rect 3824 127 3900 157
tri 3900 127 3930 157 nw
tri 3988 135 4018 165 ne
rect 4018 135 4094 165
tri 4094 135 4124 165 nw
rect 4439 290 4469 351
tri 4469 290 4485 306 sw
rect 4739 290 4769 351
rect 4439 260 4545 290
tri 4545 260 4575 290 sw
rect 4439 159 4469 260
tri 4469 244 4485 260 nw
tri 4529 244 4545 260 ne
tri 4469 159 4485 175 sw
tri 4529 159 4545 175 se
rect 4545 159 4575 260
tri 4634 260 4664 290 se
rect 4664 260 4769 290
rect 4634 166 4664 260
tri 4664 244 4680 260 nw
tri 4723 244 4739 260 ne
tri 4664 166 4680 182 sw
tri 4723 166 4739 182 se
rect 4739 166 4769 260
tri 4439 129 4469 159 ne
rect 4469 129 4545 159
tri 4545 129 4575 159 nw
tri 4634 136 4664 166 ne
rect 4664 136 4739 166
tri 4739 136 4769 166 nw
rect 4941 298 4971 351
tri 4971 298 4987 314 sw
rect 4941 268 5047 298
tri 5047 268 5077 298 sw
rect 4941 167 4971 268
tri 4971 252 4987 268 nw
tri 5031 252 5047 268 ne
tri 4971 167 4987 183 sw
tri 5031 167 5047 183 se
rect 5047 167 5077 268
tri 4941 137 4971 167 ne
rect 4971 137 5047 167
tri 5047 137 5077 167 nw
rect 5422 288 5452 349
tri 5452 288 5468 304 sw
rect 5616 296 5646 349
tri 5646 296 5662 312 sw
rect 5422 258 5528 288
tri 5528 258 5558 288 sw
rect 5616 266 5722 296
tri 5722 266 5752 296 sw
rect 5422 157 5452 258
tri 5452 242 5468 258 nw
tri 5512 242 5528 258 ne
tri 5452 157 5468 173 sw
tri 5512 157 5528 173 se
rect 5528 157 5558 258
rect 5616 165 5646 266
tri 5646 250 5662 266 nw
tri 5706 250 5722 266 ne
tri 5646 165 5662 181 sw
tri 5706 165 5722 181 se
rect 5722 165 5752 266
tri 5422 127 5452 157 ne
rect 5452 127 5528 157
tri 5528 127 5558 157 nw
tri 5616 135 5646 165 ne
rect 5646 135 5722 165
tri 5722 135 5752 165 nw
rect 6088 288 6118 349
tri 6118 288 6134 304 sw
rect 6282 296 6312 349
tri 6312 296 6328 312 sw
rect 6088 258 6194 288
tri 6194 258 6224 288 sw
rect 6282 266 6388 296
tri 6388 266 6418 296 sw
rect 6088 157 6118 258
tri 6118 242 6134 258 nw
tri 6178 242 6194 258 ne
tri 6118 157 6134 173 sw
tri 6178 157 6194 173 se
rect 6194 157 6224 258
rect 6282 165 6312 266
tri 6312 250 6328 266 nw
tri 6372 250 6388 266 ne
tri 6312 165 6328 181 sw
tri 6372 165 6388 181 se
rect 6388 165 6418 266
tri 6088 127 6118 157 ne
rect 6118 127 6194 157
tri 6194 127 6224 157 nw
tri 6282 135 6312 165 ne
rect 6312 135 6388 165
tri 6388 135 6418 165 nw
rect 6754 288 6784 349
tri 6784 288 6800 304 sw
rect 6948 296 6978 349
tri 6978 296 6994 312 sw
rect 6754 258 6860 288
tri 6860 258 6890 288 sw
rect 6948 266 7054 296
tri 7054 266 7084 296 sw
rect 6754 157 6784 258
tri 6784 242 6800 258 nw
tri 6844 242 6860 258 ne
tri 6784 157 6800 173 sw
tri 6844 157 6860 173 se
rect 6860 157 6890 258
rect 6948 165 6978 266
tri 6978 250 6994 266 nw
tri 7038 250 7054 266 ne
tri 6978 165 6994 181 sw
tri 7038 165 7054 181 se
rect 7054 165 7084 266
tri 6754 127 6784 157 ne
rect 6784 127 6860 157
tri 6860 127 6890 157 nw
tri 6948 135 6978 165 ne
rect 6978 135 7054 165
tri 7054 135 7084 165 nw
rect 7420 288 7450 349
tri 7450 288 7466 304 sw
rect 7614 296 7644 349
tri 7644 296 7660 312 sw
rect 7420 258 7526 288
tri 7526 258 7556 288 sw
rect 7614 266 7720 296
tri 7720 266 7750 296 sw
rect 7420 157 7450 258
tri 7450 242 7466 258 nw
tri 7510 242 7526 258 ne
tri 7450 157 7466 173 sw
tri 7510 157 7526 173 se
rect 7526 157 7556 258
rect 7614 165 7644 266
tri 7644 250 7660 266 nw
tri 7704 250 7720 266 ne
tri 7644 165 7660 181 sw
tri 7704 165 7720 181 se
rect 7720 165 7750 266
tri 7420 127 7450 157 ne
rect 7450 127 7526 157
tri 7526 127 7556 157 nw
tri 7614 135 7644 165 ne
rect 7644 135 7720 165
tri 7720 135 7750 165 nw
rect 8086 288 8116 349
tri 8116 288 8132 304 sw
rect 8280 296 8310 349
tri 8310 296 8326 312 sw
rect 8086 258 8192 288
tri 8192 258 8222 288 sw
rect 8280 266 8386 296
tri 8386 266 8416 296 sw
rect 8086 157 8116 258
tri 8116 242 8132 258 nw
tri 8176 242 8192 258 ne
tri 8116 157 8132 173 sw
tri 8176 157 8192 173 se
rect 8192 157 8222 258
rect 8280 165 8310 266
tri 8310 250 8326 266 nw
tri 8370 250 8386 266 ne
tri 8310 165 8326 181 sw
tri 8370 165 8386 181 se
rect 8386 165 8416 266
tri 8086 127 8116 157 ne
rect 8116 127 8192 157
tri 8192 127 8222 157 nw
tri 8280 135 8310 165 ne
rect 8310 135 8386 165
tri 8386 135 8416 165 nw
rect 8731 290 8761 351
tri 8761 290 8777 306 sw
rect 9031 290 9061 351
rect 8731 260 8837 290
tri 8837 260 8867 290 sw
rect 8731 159 8761 260
tri 8761 244 8777 260 nw
tri 8821 244 8837 260 ne
tri 8761 159 8777 175 sw
tri 8821 159 8837 175 se
rect 8837 159 8867 260
tri 8926 260 8956 290 se
rect 8956 260 9061 290
rect 8926 166 8956 260
tri 8956 244 8972 260 nw
tri 9015 244 9031 260 ne
tri 8956 166 8972 182 sw
tri 9015 166 9031 182 se
rect 9031 166 9061 260
tri 8731 129 8761 159 ne
rect 8761 129 8837 159
tri 8837 129 8867 159 nw
tri 8926 136 8956 166 ne
rect 8956 136 9031 166
tri 9031 136 9061 166 nw
rect 9233 298 9263 351
tri 9263 298 9279 314 sw
rect 9233 268 9339 298
tri 9339 268 9369 298 sw
rect 9233 167 9263 268
tri 9263 252 9279 268 nw
tri 9323 252 9339 268 ne
tri 9263 167 9279 183 sw
tri 9323 167 9339 183 se
rect 9339 167 9369 268
tri 9233 137 9263 167 ne
rect 9263 137 9339 167
tri 9339 137 9369 167 nw
rect 9714 288 9744 349
tri 9744 288 9760 304 sw
rect 9908 296 9938 349
tri 9938 296 9954 312 sw
rect 9714 258 9820 288
tri 9820 258 9850 288 sw
rect 9908 266 10014 296
tri 10014 266 10044 296 sw
rect 9714 157 9744 258
tri 9744 242 9760 258 nw
tri 9804 242 9820 258 ne
tri 9744 157 9760 173 sw
tri 9804 157 9820 173 se
rect 9820 157 9850 258
rect 9908 165 9938 266
tri 9938 250 9954 266 nw
tri 9998 250 10014 266 ne
tri 9938 165 9954 181 sw
tri 9998 165 10014 181 se
rect 10014 165 10044 266
tri 9714 127 9744 157 ne
rect 9744 127 9820 157
tri 9820 127 9850 157 nw
tri 9908 135 9938 165 ne
rect 9938 135 10014 165
tri 10014 135 10044 165 nw
rect 10380 288 10410 349
tri 10410 288 10426 304 sw
rect 10574 296 10604 349
tri 10604 296 10620 312 sw
rect 10380 258 10486 288
tri 10486 258 10516 288 sw
rect 10574 266 10680 296
tri 10680 266 10710 296 sw
rect 10380 157 10410 258
tri 10410 242 10426 258 nw
tri 10470 242 10486 258 ne
tri 10410 157 10426 173 sw
tri 10470 157 10486 173 se
rect 10486 157 10516 258
rect 10574 165 10604 266
tri 10604 250 10620 266 nw
tri 10664 250 10680 266 ne
tri 10604 165 10620 181 sw
tri 10664 165 10680 181 se
rect 10680 165 10710 266
tri 10380 127 10410 157 ne
rect 10410 127 10486 157
tri 10486 127 10516 157 nw
tri 10574 135 10604 165 ne
rect 10604 135 10680 165
tri 10680 135 10710 165 nw
rect 11046 288 11076 349
tri 11076 288 11092 304 sw
rect 11240 296 11270 349
tri 11270 296 11286 312 sw
rect 11046 258 11152 288
tri 11152 258 11182 288 sw
rect 11240 266 11346 296
tri 11346 266 11376 296 sw
rect 11046 157 11076 258
tri 11076 242 11092 258 nw
tri 11136 242 11152 258 ne
tri 11076 157 11092 173 sw
tri 11136 157 11152 173 se
rect 11152 157 11182 258
rect 11240 165 11270 266
tri 11270 250 11286 266 nw
tri 11330 250 11346 266 ne
tri 11270 165 11286 181 sw
tri 11330 165 11346 181 se
rect 11346 165 11376 266
tri 11046 127 11076 157 ne
rect 11076 127 11152 157
tri 11152 127 11182 157 nw
tri 11240 135 11270 165 ne
rect 11270 135 11346 165
tri 11346 135 11376 165 nw
rect 11712 288 11742 349
tri 11742 288 11758 304 sw
rect 11906 296 11936 349
tri 11936 296 11952 312 sw
rect 11712 258 11818 288
tri 11818 258 11848 288 sw
rect 11906 266 12012 296
tri 12012 266 12042 296 sw
rect 11712 157 11742 258
tri 11742 242 11758 258 nw
tri 11802 242 11818 258 ne
tri 11742 157 11758 173 sw
tri 11802 157 11818 173 se
rect 11818 157 11848 258
rect 11906 165 11936 266
tri 11936 250 11952 266 nw
tri 11996 250 12012 266 ne
tri 11936 165 11952 181 sw
tri 11996 165 12012 181 se
rect 12012 165 12042 266
tri 11712 127 11742 157 ne
rect 11742 127 11818 157
tri 11818 127 11848 157 nw
tri 11906 135 11936 165 ne
rect 11936 135 12012 165
tri 12012 135 12042 165 nw
rect 12378 288 12408 349
tri 12408 288 12424 304 sw
rect 12572 296 12602 349
tri 12602 296 12618 312 sw
rect 12378 258 12484 288
tri 12484 258 12514 288 sw
rect 12572 266 12678 296
tri 12678 266 12708 296 sw
rect 12378 157 12408 258
tri 12408 242 12424 258 nw
tri 12468 242 12484 258 ne
tri 12408 157 12424 173 sw
tri 12468 157 12484 173 se
rect 12484 157 12514 258
rect 12572 165 12602 266
tri 12602 250 12618 266 nw
tri 12662 250 12678 266 ne
tri 12602 165 12618 181 sw
tri 12662 165 12678 181 se
rect 12678 165 12708 266
tri 12378 127 12408 157 ne
rect 12408 127 12484 157
tri 12484 127 12514 157 nw
tri 12572 135 12602 165 ne
rect 12602 135 12678 165
tri 12678 135 12708 165 nw
rect 13044 288 13074 349
tri 13074 288 13090 304 sw
rect 13238 296 13268 349
tri 13268 296 13284 312 sw
rect 13044 258 13150 288
tri 13150 258 13180 288 sw
rect 13238 266 13344 296
tri 13344 266 13374 296 sw
rect 13044 157 13074 258
tri 13074 242 13090 258 nw
tri 13134 242 13150 258 ne
tri 13074 157 13090 173 sw
tri 13134 157 13150 173 se
rect 13150 157 13180 258
rect 13238 165 13268 266
tri 13268 250 13284 266 nw
tri 13328 250 13344 266 ne
tri 13268 165 13284 181 sw
tri 13328 165 13344 181 se
rect 13344 165 13374 266
tri 13044 127 13074 157 ne
rect 13074 127 13150 157
tri 13150 127 13180 157 nw
tri 13238 135 13268 165 ne
rect 13268 135 13344 165
tri 13344 135 13374 165 nw
rect 13710 288 13740 349
tri 13740 288 13756 304 sw
tri 13994 296 14010 312 se
rect 14010 296 14040 349
rect 13710 258 13816 288
tri 13816 258 13846 288 sw
tri 13904 266 13934 296 se
rect 13934 266 14040 296
rect 13710 157 13740 258
tri 13740 242 13756 258 nw
tri 13800 242 13816 258 ne
tri 13740 157 13756 173 sw
tri 13800 157 13816 173 se
rect 13816 157 13846 258
rect 13904 165 13934 266
tri 13934 250 13950 266 nw
tri 13994 250 14010 266 ne
tri 13934 165 13950 181 sw
tri 13994 165 14010 181 se
rect 14010 165 14040 266
tri 13710 127 13740 157 ne
rect 13740 127 13816 157
tri 13816 127 13846 157 nw
tri 13904 135 13934 165 ne
rect 13934 135 14010 165
tri 14010 135 14040 165 nw
rect 14376 288 14406 349
tri 14406 288 14422 304 sw
rect 14570 296 14600 349
tri 14600 296 14616 312 sw
rect 14376 258 14482 288
tri 14482 258 14512 288 sw
rect 14570 266 14676 296
tri 14676 266 14706 296 sw
rect 14376 157 14406 258
tri 14406 242 14422 258 nw
tri 14466 242 14482 258 ne
tri 14406 157 14422 173 sw
tri 14466 157 14482 173 se
rect 14482 157 14512 258
rect 14570 251 14601 266
tri 14601 251 14616 266 nw
tri 14660 251 14675 266 ne
rect 14675 251 14706 266
rect 14570 165 14600 251
tri 14600 165 14616 181 sw
tri 14660 165 14676 181 se
rect 14676 165 14706 251
tri 14376 127 14406 157 ne
rect 14406 127 14482 157
tri 14482 127 14512 157 nw
tri 14570 135 14600 165 ne
rect 14600 135 14676 165
tri 14676 135 14706 165 nw
<< pmos >>
rect 247 1004 277 1404
rect 335 1004 365 1404
rect 423 1004 453 1404
rect 511 1004 541 1404
rect 599 1004 629 1404
rect 687 1004 717 1404
rect 1149 1004 1179 1404
rect 1237 1004 1267 1404
rect 1325 1004 1355 1404
rect 1413 1004 1443 1404
rect 1815 1004 1845 1404
rect 1903 1004 1933 1404
rect 1991 1004 2021 1404
rect 2079 1004 2109 1404
rect 2481 1004 2511 1404
rect 2569 1004 2599 1404
rect 2657 1004 2687 1404
rect 2745 1004 2775 1404
rect 3147 1004 3177 1404
rect 3235 1004 3265 1404
rect 3323 1004 3353 1404
rect 3411 1004 3441 1404
rect 3813 1004 3843 1404
rect 3901 1004 3931 1404
rect 3989 1004 4019 1404
rect 4077 1004 4107 1404
rect 4539 1004 4569 1404
rect 4627 1004 4657 1404
rect 4715 1004 4745 1404
rect 4803 1004 4833 1404
rect 4891 1004 4921 1404
rect 4979 1004 5009 1404
rect 5441 1004 5471 1404
rect 5529 1004 5559 1404
rect 5617 1004 5647 1404
rect 5705 1004 5735 1404
rect 6107 1004 6137 1404
rect 6195 1004 6225 1404
rect 6283 1004 6313 1404
rect 6371 1004 6401 1404
rect 6773 1004 6803 1404
rect 6861 1004 6891 1404
rect 6949 1004 6979 1404
rect 7037 1004 7067 1404
rect 7439 1004 7469 1404
rect 7527 1004 7557 1404
rect 7615 1004 7645 1404
rect 7703 1004 7733 1404
rect 8105 1004 8135 1404
rect 8193 1004 8223 1404
rect 8281 1004 8311 1404
rect 8369 1004 8399 1404
rect 8831 1004 8861 1404
rect 8919 1004 8949 1404
rect 9007 1004 9037 1404
rect 9095 1004 9125 1404
rect 9183 1004 9213 1404
rect 9271 1004 9301 1404
rect 9733 1004 9763 1404
rect 9821 1004 9851 1404
rect 9909 1004 9939 1404
rect 9997 1004 10027 1404
rect 10399 1004 10429 1404
rect 10487 1004 10517 1404
rect 10575 1004 10605 1404
rect 10663 1004 10693 1404
rect 11065 1004 11095 1404
rect 11153 1004 11183 1404
rect 11241 1004 11271 1404
rect 11329 1004 11359 1404
rect 11731 1004 11761 1404
rect 11819 1004 11849 1404
rect 11907 1004 11937 1404
rect 11995 1004 12025 1404
rect 12397 1004 12427 1404
rect 12485 1004 12515 1404
rect 12573 1004 12603 1404
rect 12661 1004 12691 1404
rect 13063 1005 13093 1405
rect 13151 1005 13181 1405
rect 13239 1005 13269 1405
rect 13327 1005 13357 1405
rect 13727 1005 13757 1405
rect 13815 1005 13845 1405
rect 13903 1005 13933 1405
rect 13991 1005 14021 1405
rect 14395 1005 14425 1405
rect 14483 1005 14513 1405
rect 14571 1005 14601 1405
rect 14659 1005 14689 1405
<< ndiff >>
rect 91 335 147 351
rect 91 301 101 335
rect 135 301 147 335
rect 91 263 147 301
rect 177 335 447 351
rect 177 306 198 335
tri 177 290 193 306 ne
rect 193 301 198 306
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 447 335
rect 193 290 447 301
rect 477 335 533 351
rect 477 301 489 335
rect 523 301 533 335
rect 91 229 101 263
rect 135 229 147 263
tri 253 260 283 290 ne
rect 283 263 342 290
rect 91 195 147 229
rect 91 161 101 195
rect 135 161 147 195
rect 91 129 147 161
tri 177 244 193 260 se
rect 193 244 237 260
tri 237 244 253 260 sw
rect 177 210 253 244
rect 177 176 198 210
rect 232 176 253 210
rect 177 175 253 176
tri 177 159 193 175 ne
rect 193 159 237 175
tri 237 159 253 175 nw
rect 283 229 295 263
rect 329 229 342 263
tri 342 260 372 290 nw
rect 283 195 342 229
rect 283 161 295 195
rect 329 161 342 195
tri 372 244 388 260 se
rect 388 244 431 260
tri 431 244 447 260 sw
rect 372 216 447 244
rect 372 182 393 216
rect 427 182 447 216
tri 372 166 388 182 ne
rect 388 166 431 182
tri 431 166 447 182 nw
tri 147 129 177 159 sw
tri 253 129 283 159 se
rect 283 136 342 161
tri 342 136 372 166 sw
tri 447 136 477 166 se
rect 477 136 533 301
rect 283 129 533 136
rect 91 125 533 129
rect 91 91 101 125
rect 135 91 295 125
rect 329 91 392 125
rect 426 91 489 125
rect 523 91 533 125
rect 91 75 533 91
rect 593 335 649 351
rect 593 301 603 335
rect 637 301 649 335
rect 593 263 649 301
rect 679 314 841 351
tri 679 298 695 314 ne
rect 695 298 841 314
tri 755 268 785 298 ne
rect 593 229 603 263
rect 637 229 649 263
rect 593 195 649 229
rect 593 161 603 195
rect 637 161 649 195
tri 679 252 695 268 se
rect 695 252 739 268
tri 739 252 755 268 sw
rect 679 219 755 252
rect 679 185 700 219
rect 734 185 755 219
rect 679 183 755 185
tri 679 167 695 183 ne
rect 695 167 739 183
tri 739 167 755 183 nw
rect 785 263 841 298
rect 785 229 797 263
rect 831 229 841 263
rect 785 195 841 229
rect 593 137 649 161
tri 649 137 679 167 sw
tri 755 137 785 167 se
rect 785 161 797 195
rect 831 161 841 195
rect 785 137 841 161
rect 593 125 841 137
rect 593 91 603 125
rect 637 91 700 125
rect 734 91 797 125
rect 831 91 841 125
rect 593 75 841 91
rect 1074 333 1130 349
rect 1074 299 1084 333
rect 1118 299 1130 333
rect 1074 261 1130 299
rect 1160 333 1324 349
rect 1160 304 1181 333
tri 1160 288 1176 304 ne
rect 1176 299 1181 304
rect 1215 299 1278 333
rect 1312 299 1324 333
rect 1176 288 1324 299
rect 1354 312 1516 349
tri 1354 296 1370 312 ne
rect 1370 296 1516 312
rect 1074 227 1084 261
rect 1118 227 1130 261
tri 1236 258 1266 288 ne
rect 1266 261 1324 288
tri 1430 266 1460 296 ne
rect 1074 193 1130 227
rect 1074 159 1084 193
rect 1118 159 1130 193
rect 1074 127 1130 159
tri 1160 242 1176 258 se
rect 1176 242 1220 258
tri 1220 242 1236 258 sw
rect 1160 208 1236 242
rect 1160 174 1181 208
rect 1215 174 1236 208
rect 1160 173 1236 174
tri 1160 157 1176 173 ne
rect 1176 157 1220 173
tri 1220 157 1236 173 nw
rect 1266 227 1278 261
rect 1312 227 1324 261
rect 1266 193 1324 227
rect 1266 159 1278 193
rect 1312 159 1324 193
tri 1354 250 1370 266 se
rect 1370 250 1414 266
tri 1414 250 1430 266 sw
rect 1354 217 1430 250
rect 1354 183 1375 217
rect 1409 183 1430 217
rect 1354 181 1430 183
tri 1354 165 1370 181 ne
rect 1370 165 1414 181
tri 1414 165 1430 181 nw
rect 1460 261 1516 296
rect 1460 227 1472 261
rect 1506 227 1516 261
rect 1460 193 1516 227
tri 1130 127 1160 157 sw
tri 1236 127 1266 157 se
rect 1266 135 1324 159
tri 1324 135 1354 165 sw
tri 1430 135 1460 165 se
rect 1460 159 1472 193
rect 1506 159 1516 193
rect 1460 135 1516 159
rect 1266 127 1516 135
rect 1074 123 1516 127
rect 1074 89 1084 123
rect 1118 89 1278 123
rect 1312 89 1375 123
rect 1409 89 1472 123
rect 1506 89 1516 123
rect 1074 73 1516 89
rect 1740 333 1796 349
rect 1740 299 1750 333
rect 1784 299 1796 333
rect 1740 261 1796 299
rect 1826 333 1990 349
rect 1826 304 1847 333
tri 1826 288 1842 304 ne
rect 1842 299 1847 304
rect 1881 299 1944 333
rect 1978 299 1990 333
rect 1842 288 1990 299
rect 2020 312 2182 349
tri 2020 296 2036 312 ne
rect 2036 296 2182 312
rect 1740 227 1750 261
rect 1784 227 1796 261
tri 1902 258 1932 288 ne
rect 1932 261 1990 288
tri 2096 266 2126 296 ne
rect 1740 193 1796 227
rect 1740 159 1750 193
rect 1784 159 1796 193
rect 1740 127 1796 159
tri 1826 242 1842 258 se
rect 1842 242 1886 258
tri 1886 242 1902 258 sw
rect 1826 208 1902 242
rect 1826 174 1847 208
rect 1881 174 1902 208
rect 1826 173 1902 174
tri 1826 157 1842 173 ne
rect 1842 157 1886 173
tri 1886 157 1902 173 nw
rect 1932 227 1944 261
rect 1978 227 1990 261
rect 1932 193 1990 227
rect 1932 159 1944 193
rect 1978 159 1990 193
tri 2020 250 2036 266 se
rect 2036 250 2080 266
tri 2080 250 2096 266 sw
rect 2020 217 2096 250
rect 2020 183 2041 217
rect 2075 183 2096 217
rect 2020 181 2096 183
tri 2020 165 2036 181 ne
rect 2036 165 2080 181
tri 2080 165 2096 181 nw
rect 2126 261 2182 296
rect 2126 227 2138 261
rect 2172 227 2182 261
rect 2126 193 2182 227
tri 1796 127 1826 157 sw
tri 1902 127 1932 157 se
rect 1932 135 1990 159
tri 1990 135 2020 165 sw
tri 2096 135 2126 165 se
rect 2126 159 2138 193
rect 2172 159 2182 193
rect 2126 135 2182 159
rect 1932 127 2182 135
rect 1740 123 2182 127
rect 1740 89 1750 123
rect 1784 89 1944 123
rect 1978 89 2041 123
rect 2075 89 2138 123
rect 2172 89 2182 123
rect 1740 73 2182 89
rect 2406 333 2462 349
rect 2406 299 2416 333
rect 2450 299 2462 333
rect 2406 261 2462 299
rect 2492 333 2656 349
rect 2492 304 2513 333
tri 2492 288 2508 304 ne
rect 2508 299 2513 304
rect 2547 299 2610 333
rect 2644 299 2656 333
rect 2508 288 2656 299
rect 2686 312 2848 349
tri 2686 296 2702 312 ne
rect 2702 296 2848 312
rect 2406 227 2416 261
rect 2450 227 2462 261
tri 2568 258 2598 288 ne
rect 2598 261 2656 288
tri 2762 266 2792 296 ne
rect 2406 193 2462 227
rect 2406 159 2416 193
rect 2450 159 2462 193
rect 2406 127 2462 159
tri 2492 242 2508 258 se
rect 2508 242 2552 258
tri 2552 242 2568 258 sw
rect 2492 208 2568 242
rect 2492 174 2513 208
rect 2547 174 2568 208
rect 2492 173 2568 174
tri 2492 157 2508 173 ne
rect 2508 157 2552 173
tri 2552 157 2568 173 nw
rect 2598 227 2610 261
rect 2644 227 2656 261
rect 2598 193 2656 227
rect 2598 159 2610 193
rect 2644 159 2656 193
tri 2686 250 2702 266 se
rect 2702 250 2746 266
tri 2746 250 2762 266 sw
rect 2686 217 2762 250
rect 2686 183 2707 217
rect 2741 183 2762 217
rect 2686 181 2762 183
tri 2686 165 2702 181 ne
rect 2702 165 2746 181
tri 2746 165 2762 181 nw
rect 2792 261 2848 296
rect 2792 227 2804 261
rect 2838 227 2848 261
rect 2792 193 2848 227
tri 2462 127 2492 157 sw
tri 2568 127 2598 157 se
rect 2598 135 2656 159
tri 2656 135 2686 165 sw
tri 2762 135 2792 165 se
rect 2792 159 2804 193
rect 2838 159 2848 193
rect 2792 135 2848 159
rect 2598 127 2848 135
rect 2406 123 2848 127
rect 2406 89 2416 123
rect 2450 89 2610 123
rect 2644 89 2707 123
rect 2741 89 2804 123
rect 2838 89 2848 123
rect 2406 73 2848 89
rect 3072 333 3128 349
rect 3072 299 3082 333
rect 3116 299 3128 333
rect 3072 261 3128 299
rect 3158 333 3322 349
rect 3158 304 3179 333
tri 3158 288 3174 304 ne
rect 3174 299 3179 304
rect 3213 299 3276 333
rect 3310 299 3322 333
rect 3174 288 3322 299
rect 3352 312 3514 349
tri 3352 296 3368 312 ne
rect 3368 296 3514 312
rect 3072 227 3082 261
rect 3116 227 3128 261
tri 3234 258 3264 288 ne
rect 3264 261 3322 288
tri 3428 266 3458 296 ne
rect 3072 193 3128 227
rect 3072 159 3082 193
rect 3116 159 3128 193
rect 3072 127 3128 159
tri 3158 242 3174 258 se
rect 3174 242 3218 258
tri 3218 242 3234 258 sw
rect 3158 208 3234 242
rect 3158 174 3179 208
rect 3213 174 3234 208
rect 3158 173 3234 174
tri 3158 157 3174 173 ne
rect 3174 157 3218 173
tri 3218 157 3234 173 nw
rect 3264 227 3276 261
rect 3310 227 3322 261
rect 3264 193 3322 227
rect 3264 159 3276 193
rect 3310 159 3322 193
tri 3352 250 3368 266 se
rect 3368 250 3412 266
tri 3412 250 3428 266 sw
rect 3352 217 3428 250
rect 3352 183 3373 217
rect 3407 183 3428 217
rect 3352 181 3428 183
tri 3352 165 3368 181 ne
rect 3368 165 3412 181
tri 3412 165 3428 181 nw
rect 3458 261 3514 296
rect 3458 227 3470 261
rect 3504 227 3514 261
rect 3458 193 3514 227
tri 3128 127 3158 157 sw
tri 3234 127 3264 157 se
rect 3264 135 3322 159
tri 3322 135 3352 165 sw
tri 3428 135 3458 165 se
rect 3458 159 3470 193
rect 3504 159 3514 193
rect 3458 135 3514 159
rect 3264 127 3514 135
rect 3072 123 3514 127
rect 3072 89 3082 123
rect 3116 89 3276 123
rect 3310 89 3373 123
rect 3407 89 3470 123
rect 3504 89 3514 123
rect 3072 73 3514 89
rect 3738 333 3794 349
rect 3738 299 3748 333
rect 3782 299 3794 333
rect 3738 261 3794 299
rect 3824 333 3988 349
rect 3824 304 3845 333
tri 3824 288 3840 304 ne
rect 3840 299 3845 304
rect 3879 299 3942 333
rect 3976 299 3988 333
rect 3840 288 3988 299
rect 4018 312 4180 349
tri 4018 296 4034 312 ne
rect 4034 296 4180 312
rect 3738 227 3748 261
rect 3782 227 3794 261
tri 3900 258 3930 288 ne
rect 3930 261 3988 288
tri 4094 266 4124 296 ne
rect 3738 193 3794 227
rect 3738 159 3748 193
rect 3782 159 3794 193
rect 3738 127 3794 159
tri 3824 242 3840 258 se
rect 3840 242 3884 258
tri 3884 242 3900 258 sw
rect 3824 208 3900 242
rect 3824 174 3845 208
rect 3879 174 3900 208
rect 3824 173 3900 174
tri 3824 157 3840 173 ne
rect 3840 157 3884 173
tri 3884 157 3900 173 nw
rect 3930 227 3942 261
rect 3976 227 3988 261
rect 3930 193 3988 227
rect 3930 159 3942 193
rect 3976 159 3988 193
tri 4018 250 4034 266 se
rect 4034 250 4078 266
tri 4078 250 4094 266 sw
rect 4018 217 4094 250
rect 4018 183 4039 217
rect 4073 183 4094 217
rect 4018 181 4094 183
tri 4018 165 4034 181 ne
rect 4034 165 4078 181
tri 4078 165 4094 181 nw
rect 4124 261 4180 296
rect 4124 227 4136 261
rect 4170 227 4180 261
rect 4124 193 4180 227
tri 3794 127 3824 157 sw
tri 3900 127 3930 157 se
rect 3930 135 3988 159
tri 3988 135 4018 165 sw
tri 4094 135 4124 165 se
rect 4124 159 4136 193
rect 4170 159 4180 193
rect 4124 135 4180 159
rect 3930 127 4180 135
rect 3738 123 4180 127
rect 3738 89 3748 123
rect 3782 89 3942 123
rect 3976 89 4039 123
rect 4073 89 4136 123
rect 4170 89 4180 123
rect 3738 73 4180 89
rect 4383 335 4439 351
rect 4383 301 4393 335
rect 4427 301 4439 335
rect 4383 263 4439 301
rect 4469 335 4739 351
rect 4469 306 4490 335
tri 4469 290 4485 306 ne
rect 4485 301 4490 306
rect 4524 301 4587 335
rect 4621 301 4684 335
rect 4718 301 4739 335
rect 4485 290 4739 301
rect 4769 335 4825 351
rect 4769 301 4781 335
rect 4815 301 4825 335
rect 4383 229 4393 263
rect 4427 229 4439 263
tri 4545 260 4575 290 ne
rect 4575 263 4634 290
rect 4383 195 4439 229
rect 4383 161 4393 195
rect 4427 161 4439 195
rect 4383 129 4439 161
tri 4469 244 4485 260 se
rect 4485 244 4529 260
tri 4529 244 4545 260 sw
rect 4469 210 4545 244
rect 4469 176 4490 210
rect 4524 176 4545 210
rect 4469 175 4545 176
tri 4469 159 4485 175 ne
rect 4485 159 4529 175
tri 4529 159 4545 175 nw
rect 4575 229 4587 263
rect 4621 229 4634 263
tri 4634 260 4664 290 nw
rect 4575 195 4634 229
rect 4575 161 4587 195
rect 4621 161 4634 195
tri 4664 244 4680 260 se
rect 4680 244 4723 260
tri 4723 244 4739 260 sw
rect 4664 216 4739 244
rect 4664 182 4685 216
rect 4719 182 4739 216
tri 4664 166 4680 182 ne
rect 4680 166 4723 182
tri 4723 166 4739 182 nw
tri 4439 129 4469 159 sw
tri 4545 129 4575 159 se
rect 4575 136 4634 161
tri 4634 136 4664 166 sw
tri 4739 136 4769 166 se
rect 4769 136 4825 301
rect 4575 129 4825 136
rect 4383 125 4825 129
rect 4383 91 4393 125
rect 4427 91 4587 125
rect 4621 91 4684 125
rect 4718 91 4781 125
rect 4815 91 4825 125
rect 4383 75 4825 91
rect 4885 335 4941 351
rect 4885 301 4895 335
rect 4929 301 4941 335
rect 4885 263 4941 301
rect 4971 314 5133 351
tri 4971 298 4987 314 ne
rect 4987 298 5133 314
tri 5047 268 5077 298 ne
rect 4885 229 4895 263
rect 4929 229 4941 263
rect 4885 195 4941 229
rect 4885 161 4895 195
rect 4929 161 4941 195
tri 4971 252 4987 268 se
rect 4987 252 5031 268
tri 5031 252 5047 268 sw
rect 4971 219 5047 252
rect 4971 185 4992 219
rect 5026 185 5047 219
rect 4971 183 5047 185
tri 4971 167 4987 183 ne
rect 4987 167 5031 183
tri 5031 167 5047 183 nw
rect 5077 263 5133 298
rect 5077 229 5089 263
rect 5123 229 5133 263
rect 5077 195 5133 229
rect 4885 137 4941 161
tri 4941 137 4971 167 sw
tri 5047 137 5077 167 se
rect 5077 161 5089 195
rect 5123 161 5133 195
rect 5077 137 5133 161
rect 4885 125 5133 137
rect 4885 91 4895 125
rect 4929 91 4992 125
rect 5026 91 5089 125
rect 5123 91 5133 125
rect 4885 75 5133 91
rect 5366 333 5422 349
rect 5366 299 5376 333
rect 5410 299 5422 333
rect 5366 261 5422 299
rect 5452 333 5616 349
rect 5452 304 5473 333
tri 5452 288 5468 304 ne
rect 5468 299 5473 304
rect 5507 299 5570 333
rect 5604 299 5616 333
rect 5468 288 5616 299
rect 5646 312 5808 349
tri 5646 296 5662 312 ne
rect 5662 296 5808 312
rect 5366 227 5376 261
rect 5410 227 5422 261
tri 5528 258 5558 288 ne
rect 5558 261 5616 288
tri 5722 266 5752 296 ne
rect 5366 193 5422 227
rect 5366 159 5376 193
rect 5410 159 5422 193
rect 5366 127 5422 159
tri 5452 242 5468 258 se
rect 5468 242 5512 258
tri 5512 242 5528 258 sw
rect 5452 208 5528 242
rect 5452 174 5473 208
rect 5507 174 5528 208
rect 5452 173 5528 174
tri 5452 157 5468 173 ne
rect 5468 157 5512 173
tri 5512 157 5528 173 nw
rect 5558 227 5570 261
rect 5604 227 5616 261
rect 5558 193 5616 227
rect 5558 159 5570 193
rect 5604 159 5616 193
tri 5646 250 5662 266 se
rect 5662 250 5706 266
tri 5706 250 5722 266 sw
rect 5646 217 5722 250
rect 5646 183 5667 217
rect 5701 183 5722 217
rect 5646 181 5722 183
tri 5646 165 5662 181 ne
rect 5662 165 5706 181
tri 5706 165 5722 181 nw
rect 5752 261 5808 296
rect 5752 227 5764 261
rect 5798 227 5808 261
rect 5752 193 5808 227
tri 5422 127 5452 157 sw
tri 5528 127 5558 157 se
rect 5558 135 5616 159
tri 5616 135 5646 165 sw
tri 5722 135 5752 165 se
rect 5752 159 5764 193
rect 5798 159 5808 193
rect 5752 135 5808 159
rect 5558 127 5808 135
rect 5366 123 5808 127
rect 5366 89 5376 123
rect 5410 89 5570 123
rect 5604 89 5667 123
rect 5701 89 5764 123
rect 5798 89 5808 123
rect 5366 73 5808 89
rect 6032 333 6088 349
rect 6032 299 6042 333
rect 6076 299 6088 333
rect 6032 261 6088 299
rect 6118 333 6282 349
rect 6118 304 6139 333
tri 6118 288 6134 304 ne
rect 6134 299 6139 304
rect 6173 299 6236 333
rect 6270 299 6282 333
rect 6134 288 6282 299
rect 6312 312 6474 349
tri 6312 296 6328 312 ne
rect 6328 296 6474 312
rect 6032 227 6042 261
rect 6076 227 6088 261
tri 6194 258 6224 288 ne
rect 6224 261 6282 288
tri 6388 266 6418 296 ne
rect 6032 193 6088 227
rect 6032 159 6042 193
rect 6076 159 6088 193
rect 6032 127 6088 159
tri 6118 242 6134 258 se
rect 6134 242 6178 258
tri 6178 242 6194 258 sw
rect 6118 208 6194 242
rect 6118 174 6139 208
rect 6173 174 6194 208
rect 6118 173 6194 174
tri 6118 157 6134 173 ne
rect 6134 157 6178 173
tri 6178 157 6194 173 nw
rect 6224 227 6236 261
rect 6270 227 6282 261
rect 6224 193 6282 227
rect 6224 159 6236 193
rect 6270 159 6282 193
tri 6312 250 6328 266 se
rect 6328 250 6372 266
tri 6372 250 6388 266 sw
rect 6312 217 6388 250
rect 6312 183 6333 217
rect 6367 183 6388 217
rect 6312 181 6388 183
tri 6312 165 6328 181 ne
rect 6328 165 6372 181
tri 6372 165 6388 181 nw
rect 6418 261 6474 296
rect 6418 227 6430 261
rect 6464 227 6474 261
rect 6418 193 6474 227
tri 6088 127 6118 157 sw
tri 6194 127 6224 157 se
rect 6224 135 6282 159
tri 6282 135 6312 165 sw
tri 6388 135 6418 165 se
rect 6418 159 6430 193
rect 6464 159 6474 193
rect 6418 135 6474 159
rect 6224 127 6474 135
rect 6032 123 6474 127
rect 6032 89 6042 123
rect 6076 89 6236 123
rect 6270 89 6333 123
rect 6367 89 6430 123
rect 6464 89 6474 123
rect 6032 73 6474 89
rect 6698 333 6754 349
rect 6698 299 6708 333
rect 6742 299 6754 333
rect 6698 261 6754 299
rect 6784 333 6948 349
rect 6784 304 6805 333
tri 6784 288 6800 304 ne
rect 6800 299 6805 304
rect 6839 299 6902 333
rect 6936 299 6948 333
rect 6800 288 6948 299
rect 6978 312 7140 349
tri 6978 296 6994 312 ne
rect 6994 296 7140 312
rect 6698 227 6708 261
rect 6742 227 6754 261
tri 6860 258 6890 288 ne
rect 6890 261 6948 288
tri 7054 266 7084 296 ne
rect 6698 193 6754 227
rect 6698 159 6708 193
rect 6742 159 6754 193
rect 6698 127 6754 159
tri 6784 242 6800 258 se
rect 6800 242 6844 258
tri 6844 242 6860 258 sw
rect 6784 208 6860 242
rect 6784 174 6805 208
rect 6839 174 6860 208
rect 6784 173 6860 174
tri 6784 157 6800 173 ne
rect 6800 157 6844 173
tri 6844 157 6860 173 nw
rect 6890 227 6902 261
rect 6936 227 6948 261
rect 6890 193 6948 227
rect 6890 159 6902 193
rect 6936 159 6948 193
tri 6978 250 6994 266 se
rect 6994 250 7038 266
tri 7038 250 7054 266 sw
rect 6978 217 7054 250
rect 6978 183 6999 217
rect 7033 183 7054 217
rect 6978 181 7054 183
tri 6978 165 6994 181 ne
rect 6994 165 7038 181
tri 7038 165 7054 181 nw
rect 7084 261 7140 296
rect 7084 227 7096 261
rect 7130 227 7140 261
rect 7084 193 7140 227
tri 6754 127 6784 157 sw
tri 6860 127 6890 157 se
rect 6890 135 6948 159
tri 6948 135 6978 165 sw
tri 7054 135 7084 165 se
rect 7084 159 7096 193
rect 7130 159 7140 193
rect 7084 135 7140 159
rect 6890 127 7140 135
rect 6698 123 7140 127
rect 6698 89 6708 123
rect 6742 89 6902 123
rect 6936 89 6999 123
rect 7033 89 7096 123
rect 7130 89 7140 123
rect 6698 73 7140 89
rect 7364 333 7420 349
rect 7364 299 7374 333
rect 7408 299 7420 333
rect 7364 261 7420 299
rect 7450 333 7614 349
rect 7450 304 7471 333
tri 7450 288 7466 304 ne
rect 7466 299 7471 304
rect 7505 299 7568 333
rect 7602 299 7614 333
rect 7466 288 7614 299
rect 7644 312 7806 349
tri 7644 296 7660 312 ne
rect 7660 296 7806 312
rect 7364 227 7374 261
rect 7408 227 7420 261
tri 7526 258 7556 288 ne
rect 7556 261 7614 288
tri 7720 266 7750 296 ne
rect 7364 193 7420 227
rect 7364 159 7374 193
rect 7408 159 7420 193
rect 7364 127 7420 159
tri 7450 242 7466 258 se
rect 7466 242 7510 258
tri 7510 242 7526 258 sw
rect 7450 208 7526 242
rect 7450 174 7471 208
rect 7505 174 7526 208
rect 7450 173 7526 174
tri 7450 157 7466 173 ne
rect 7466 157 7510 173
tri 7510 157 7526 173 nw
rect 7556 227 7568 261
rect 7602 227 7614 261
rect 7556 193 7614 227
rect 7556 159 7568 193
rect 7602 159 7614 193
tri 7644 250 7660 266 se
rect 7660 250 7704 266
tri 7704 250 7720 266 sw
rect 7644 217 7720 250
rect 7644 183 7665 217
rect 7699 183 7720 217
rect 7644 181 7720 183
tri 7644 165 7660 181 ne
rect 7660 165 7704 181
tri 7704 165 7720 181 nw
rect 7750 261 7806 296
rect 7750 227 7762 261
rect 7796 227 7806 261
rect 7750 193 7806 227
tri 7420 127 7450 157 sw
tri 7526 127 7556 157 se
rect 7556 135 7614 159
tri 7614 135 7644 165 sw
tri 7720 135 7750 165 se
rect 7750 159 7762 193
rect 7796 159 7806 193
rect 7750 135 7806 159
rect 7556 127 7806 135
rect 7364 123 7806 127
rect 7364 89 7374 123
rect 7408 89 7568 123
rect 7602 89 7665 123
rect 7699 89 7762 123
rect 7796 89 7806 123
rect 7364 73 7806 89
rect 8030 333 8086 349
rect 8030 299 8040 333
rect 8074 299 8086 333
rect 8030 261 8086 299
rect 8116 333 8280 349
rect 8116 304 8137 333
tri 8116 288 8132 304 ne
rect 8132 299 8137 304
rect 8171 299 8234 333
rect 8268 299 8280 333
rect 8132 288 8280 299
rect 8310 312 8472 349
tri 8310 296 8326 312 ne
rect 8326 296 8472 312
rect 8030 227 8040 261
rect 8074 227 8086 261
tri 8192 258 8222 288 ne
rect 8222 261 8280 288
tri 8386 266 8416 296 ne
rect 8030 193 8086 227
rect 8030 159 8040 193
rect 8074 159 8086 193
rect 8030 127 8086 159
tri 8116 242 8132 258 se
rect 8132 242 8176 258
tri 8176 242 8192 258 sw
rect 8116 208 8192 242
rect 8116 174 8137 208
rect 8171 174 8192 208
rect 8116 173 8192 174
tri 8116 157 8132 173 ne
rect 8132 157 8176 173
tri 8176 157 8192 173 nw
rect 8222 227 8234 261
rect 8268 227 8280 261
rect 8222 193 8280 227
rect 8222 159 8234 193
rect 8268 159 8280 193
tri 8310 250 8326 266 se
rect 8326 250 8370 266
tri 8370 250 8386 266 sw
rect 8310 217 8386 250
rect 8310 183 8331 217
rect 8365 183 8386 217
rect 8310 181 8386 183
tri 8310 165 8326 181 ne
rect 8326 165 8370 181
tri 8370 165 8386 181 nw
rect 8416 261 8472 296
rect 8416 227 8428 261
rect 8462 227 8472 261
rect 8416 193 8472 227
tri 8086 127 8116 157 sw
tri 8192 127 8222 157 se
rect 8222 135 8280 159
tri 8280 135 8310 165 sw
tri 8386 135 8416 165 se
rect 8416 159 8428 193
rect 8462 159 8472 193
rect 8416 135 8472 159
rect 8222 127 8472 135
rect 8030 123 8472 127
rect 8030 89 8040 123
rect 8074 89 8234 123
rect 8268 89 8331 123
rect 8365 89 8428 123
rect 8462 89 8472 123
rect 8030 73 8472 89
rect 8675 335 8731 351
rect 8675 301 8685 335
rect 8719 301 8731 335
rect 8675 263 8731 301
rect 8761 335 9031 351
rect 8761 306 8782 335
tri 8761 290 8777 306 ne
rect 8777 301 8782 306
rect 8816 301 8879 335
rect 8913 301 8976 335
rect 9010 301 9031 335
rect 8777 290 9031 301
rect 9061 335 9117 351
rect 9061 301 9073 335
rect 9107 301 9117 335
rect 8675 229 8685 263
rect 8719 229 8731 263
tri 8837 260 8867 290 ne
rect 8867 263 8926 290
rect 8675 195 8731 229
rect 8675 161 8685 195
rect 8719 161 8731 195
rect 8675 129 8731 161
tri 8761 244 8777 260 se
rect 8777 244 8821 260
tri 8821 244 8837 260 sw
rect 8761 210 8837 244
rect 8761 176 8782 210
rect 8816 176 8837 210
rect 8761 175 8837 176
tri 8761 159 8777 175 ne
rect 8777 159 8821 175
tri 8821 159 8837 175 nw
rect 8867 229 8879 263
rect 8913 229 8926 263
tri 8926 260 8956 290 nw
rect 8867 195 8926 229
rect 8867 161 8879 195
rect 8913 161 8926 195
tri 8956 244 8972 260 se
rect 8972 244 9015 260
tri 9015 244 9031 260 sw
rect 8956 216 9031 244
rect 8956 182 8977 216
rect 9011 182 9031 216
tri 8956 166 8972 182 ne
rect 8972 166 9015 182
tri 9015 166 9031 182 nw
tri 8731 129 8761 159 sw
tri 8837 129 8867 159 se
rect 8867 136 8926 161
tri 8926 136 8956 166 sw
tri 9031 136 9061 166 se
rect 9061 136 9117 301
rect 8867 129 9117 136
rect 8675 125 9117 129
rect 8675 91 8685 125
rect 8719 91 8879 125
rect 8913 91 8976 125
rect 9010 91 9073 125
rect 9107 91 9117 125
rect 8675 75 9117 91
rect 9177 335 9233 351
rect 9177 301 9187 335
rect 9221 301 9233 335
rect 9177 263 9233 301
rect 9263 314 9425 351
tri 9263 298 9279 314 ne
rect 9279 298 9425 314
tri 9339 268 9369 298 ne
rect 9177 229 9187 263
rect 9221 229 9233 263
rect 9177 195 9233 229
rect 9177 161 9187 195
rect 9221 161 9233 195
tri 9263 252 9279 268 se
rect 9279 252 9323 268
tri 9323 252 9339 268 sw
rect 9263 219 9339 252
rect 9263 185 9284 219
rect 9318 185 9339 219
rect 9263 183 9339 185
tri 9263 167 9279 183 ne
rect 9279 167 9323 183
tri 9323 167 9339 183 nw
rect 9369 263 9425 298
rect 9369 229 9381 263
rect 9415 229 9425 263
rect 9369 195 9425 229
rect 9177 137 9233 161
tri 9233 137 9263 167 sw
tri 9339 137 9369 167 se
rect 9369 161 9381 195
rect 9415 161 9425 195
rect 9369 137 9425 161
rect 9177 125 9425 137
rect 9177 91 9187 125
rect 9221 91 9284 125
rect 9318 91 9381 125
rect 9415 91 9425 125
rect 9177 75 9425 91
rect 9658 333 9714 349
rect 9658 299 9668 333
rect 9702 299 9714 333
rect 9658 261 9714 299
rect 9744 333 9908 349
rect 9744 304 9765 333
tri 9744 288 9760 304 ne
rect 9760 299 9765 304
rect 9799 299 9862 333
rect 9896 299 9908 333
rect 9760 288 9908 299
rect 9938 312 10100 349
tri 9938 296 9954 312 ne
rect 9954 296 10100 312
rect 9658 227 9668 261
rect 9702 227 9714 261
tri 9820 258 9850 288 ne
rect 9850 261 9908 288
tri 10014 266 10044 296 ne
rect 9658 193 9714 227
rect 9658 159 9668 193
rect 9702 159 9714 193
rect 9658 127 9714 159
tri 9744 242 9760 258 se
rect 9760 242 9804 258
tri 9804 242 9820 258 sw
rect 9744 208 9820 242
rect 9744 174 9765 208
rect 9799 174 9820 208
rect 9744 173 9820 174
tri 9744 157 9760 173 ne
rect 9760 157 9804 173
tri 9804 157 9820 173 nw
rect 9850 227 9862 261
rect 9896 227 9908 261
rect 9850 193 9908 227
rect 9850 159 9862 193
rect 9896 159 9908 193
tri 9938 250 9954 266 se
rect 9954 250 9998 266
tri 9998 250 10014 266 sw
rect 9938 217 10014 250
rect 9938 183 9959 217
rect 9993 183 10014 217
rect 9938 181 10014 183
tri 9938 165 9954 181 ne
rect 9954 165 9998 181
tri 9998 165 10014 181 nw
rect 10044 261 10100 296
rect 10044 227 10056 261
rect 10090 227 10100 261
rect 10044 193 10100 227
tri 9714 127 9744 157 sw
tri 9820 127 9850 157 se
rect 9850 135 9908 159
tri 9908 135 9938 165 sw
tri 10014 135 10044 165 se
rect 10044 159 10056 193
rect 10090 159 10100 193
rect 10044 135 10100 159
rect 9850 127 10100 135
rect 9658 123 10100 127
rect 9658 89 9668 123
rect 9702 89 9862 123
rect 9896 89 9959 123
rect 9993 89 10056 123
rect 10090 89 10100 123
rect 9658 73 10100 89
rect 10324 333 10380 349
rect 10324 299 10334 333
rect 10368 299 10380 333
rect 10324 261 10380 299
rect 10410 333 10574 349
rect 10410 304 10431 333
tri 10410 288 10426 304 ne
rect 10426 299 10431 304
rect 10465 299 10528 333
rect 10562 299 10574 333
rect 10426 288 10574 299
rect 10604 312 10766 349
tri 10604 296 10620 312 ne
rect 10620 296 10766 312
rect 10324 227 10334 261
rect 10368 227 10380 261
tri 10486 258 10516 288 ne
rect 10516 261 10574 288
tri 10680 266 10710 296 ne
rect 10324 193 10380 227
rect 10324 159 10334 193
rect 10368 159 10380 193
rect 10324 127 10380 159
tri 10410 242 10426 258 se
rect 10426 242 10470 258
tri 10470 242 10486 258 sw
rect 10410 208 10486 242
rect 10410 174 10431 208
rect 10465 174 10486 208
rect 10410 173 10486 174
tri 10410 157 10426 173 ne
rect 10426 157 10470 173
tri 10470 157 10486 173 nw
rect 10516 227 10528 261
rect 10562 227 10574 261
rect 10516 193 10574 227
rect 10516 159 10528 193
rect 10562 159 10574 193
tri 10604 250 10620 266 se
rect 10620 250 10664 266
tri 10664 250 10680 266 sw
rect 10604 217 10680 250
rect 10604 183 10625 217
rect 10659 183 10680 217
rect 10604 181 10680 183
tri 10604 165 10620 181 ne
rect 10620 165 10664 181
tri 10664 165 10680 181 nw
rect 10710 261 10766 296
rect 10710 227 10722 261
rect 10756 227 10766 261
rect 10710 193 10766 227
tri 10380 127 10410 157 sw
tri 10486 127 10516 157 se
rect 10516 135 10574 159
tri 10574 135 10604 165 sw
tri 10680 135 10710 165 se
rect 10710 159 10722 193
rect 10756 159 10766 193
rect 10710 135 10766 159
rect 10516 127 10766 135
rect 10324 123 10766 127
rect 10324 89 10334 123
rect 10368 89 10528 123
rect 10562 89 10625 123
rect 10659 89 10722 123
rect 10756 89 10766 123
rect 10324 73 10766 89
rect 10990 333 11046 349
rect 10990 299 11000 333
rect 11034 299 11046 333
rect 10990 261 11046 299
rect 11076 333 11240 349
rect 11076 304 11097 333
tri 11076 288 11092 304 ne
rect 11092 299 11097 304
rect 11131 299 11194 333
rect 11228 299 11240 333
rect 11092 288 11240 299
rect 11270 312 11432 349
tri 11270 296 11286 312 ne
rect 11286 296 11432 312
rect 10990 227 11000 261
rect 11034 227 11046 261
tri 11152 258 11182 288 ne
rect 11182 261 11240 288
tri 11346 266 11376 296 ne
rect 10990 193 11046 227
rect 10990 159 11000 193
rect 11034 159 11046 193
rect 10990 127 11046 159
tri 11076 242 11092 258 se
rect 11092 242 11136 258
tri 11136 242 11152 258 sw
rect 11076 208 11152 242
rect 11076 174 11097 208
rect 11131 174 11152 208
rect 11076 173 11152 174
tri 11076 157 11092 173 ne
rect 11092 157 11136 173
tri 11136 157 11152 173 nw
rect 11182 227 11194 261
rect 11228 227 11240 261
rect 11182 193 11240 227
rect 11182 159 11194 193
rect 11228 159 11240 193
tri 11270 250 11286 266 se
rect 11286 250 11330 266
tri 11330 250 11346 266 sw
rect 11270 217 11346 250
rect 11270 183 11291 217
rect 11325 183 11346 217
rect 11270 181 11346 183
tri 11270 165 11286 181 ne
rect 11286 165 11330 181
tri 11330 165 11346 181 nw
rect 11376 261 11432 296
rect 11376 227 11388 261
rect 11422 227 11432 261
rect 11376 193 11432 227
tri 11046 127 11076 157 sw
tri 11152 127 11182 157 se
rect 11182 135 11240 159
tri 11240 135 11270 165 sw
tri 11346 135 11376 165 se
rect 11376 159 11388 193
rect 11422 159 11432 193
rect 11376 135 11432 159
rect 11182 127 11432 135
rect 10990 123 11432 127
rect 10990 89 11000 123
rect 11034 89 11194 123
rect 11228 89 11291 123
rect 11325 89 11388 123
rect 11422 89 11432 123
rect 10990 73 11432 89
rect 11656 333 11712 349
rect 11656 299 11666 333
rect 11700 299 11712 333
rect 11656 261 11712 299
rect 11742 333 11906 349
rect 11742 304 11763 333
tri 11742 288 11758 304 ne
rect 11758 299 11763 304
rect 11797 299 11860 333
rect 11894 299 11906 333
rect 11758 288 11906 299
rect 11936 312 12098 349
tri 11936 296 11952 312 ne
rect 11952 296 12098 312
rect 11656 227 11666 261
rect 11700 227 11712 261
tri 11818 258 11848 288 ne
rect 11848 261 11906 288
tri 12012 266 12042 296 ne
rect 11656 193 11712 227
rect 11656 159 11666 193
rect 11700 159 11712 193
rect 11656 127 11712 159
tri 11742 242 11758 258 se
rect 11758 242 11802 258
tri 11802 242 11818 258 sw
rect 11742 208 11818 242
rect 11742 174 11763 208
rect 11797 174 11818 208
rect 11742 173 11818 174
tri 11742 157 11758 173 ne
rect 11758 157 11802 173
tri 11802 157 11818 173 nw
rect 11848 227 11860 261
rect 11894 227 11906 261
rect 11848 193 11906 227
rect 11848 159 11860 193
rect 11894 159 11906 193
tri 11936 250 11952 266 se
rect 11952 250 11996 266
tri 11996 250 12012 266 sw
rect 11936 217 12012 250
rect 11936 183 11957 217
rect 11991 183 12012 217
rect 11936 181 12012 183
tri 11936 165 11952 181 ne
rect 11952 165 11996 181
tri 11996 165 12012 181 nw
rect 12042 261 12098 296
rect 12042 227 12054 261
rect 12088 227 12098 261
rect 12042 193 12098 227
tri 11712 127 11742 157 sw
tri 11818 127 11848 157 se
rect 11848 135 11906 159
tri 11906 135 11936 165 sw
tri 12012 135 12042 165 se
rect 12042 159 12054 193
rect 12088 159 12098 193
rect 12042 135 12098 159
rect 11848 127 12098 135
rect 11656 123 12098 127
rect 11656 89 11666 123
rect 11700 89 11860 123
rect 11894 89 11957 123
rect 11991 89 12054 123
rect 12088 89 12098 123
rect 11656 73 12098 89
rect 12322 333 12378 349
rect 12322 299 12332 333
rect 12366 299 12378 333
rect 12322 261 12378 299
rect 12408 333 12572 349
rect 12408 304 12429 333
tri 12408 288 12424 304 ne
rect 12424 299 12429 304
rect 12463 299 12526 333
rect 12560 299 12572 333
rect 12424 288 12572 299
rect 12602 312 12764 349
tri 12602 296 12618 312 ne
rect 12618 296 12764 312
rect 12322 227 12332 261
rect 12366 227 12378 261
tri 12484 258 12514 288 ne
rect 12514 261 12572 288
tri 12678 266 12708 296 ne
rect 12322 193 12378 227
rect 12322 159 12332 193
rect 12366 159 12378 193
rect 12322 127 12378 159
tri 12408 242 12424 258 se
rect 12424 242 12468 258
tri 12468 242 12484 258 sw
rect 12408 208 12484 242
rect 12408 174 12429 208
rect 12463 174 12484 208
rect 12408 173 12484 174
tri 12408 157 12424 173 ne
rect 12424 157 12468 173
tri 12468 157 12484 173 nw
rect 12514 227 12526 261
rect 12560 227 12572 261
rect 12514 193 12572 227
rect 12514 159 12526 193
rect 12560 159 12572 193
tri 12602 250 12618 266 se
rect 12618 250 12662 266
tri 12662 250 12678 266 sw
rect 12602 217 12678 250
rect 12602 183 12623 217
rect 12657 183 12678 217
rect 12602 181 12678 183
tri 12602 165 12618 181 ne
rect 12618 165 12662 181
tri 12662 165 12678 181 nw
rect 12708 261 12764 296
rect 12708 227 12720 261
rect 12754 227 12764 261
rect 12708 193 12764 227
tri 12378 127 12408 157 sw
tri 12484 127 12514 157 se
rect 12514 135 12572 159
tri 12572 135 12602 165 sw
tri 12678 135 12708 165 se
rect 12708 159 12720 193
rect 12754 159 12764 193
rect 12708 135 12764 159
rect 12514 127 12764 135
rect 12322 123 12764 127
rect 12322 89 12332 123
rect 12366 89 12526 123
rect 12560 89 12623 123
rect 12657 89 12720 123
rect 12754 89 12764 123
rect 12322 73 12764 89
rect 12988 333 13044 349
rect 12988 299 12998 333
rect 13032 299 13044 333
rect 12988 261 13044 299
rect 13074 333 13238 349
rect 13074 304 13095 333
tri 13074 288 13090 304 ne
rect 13090 299 13095 304
rect 13129 299 13192 333
rect 13226 299 13238 333
rect 13090 288 13238 299
rect 13268 333 13428 349
rect 13268 312 13386 333
tri 13268 296 13284 312 ne
rect 13284 299 13386 312
rect 13420 299 13428 333
rect 13284 296 13428 299
rect 12988 227 12998 261
rect 13032 227 13044 261
tri 13150 258 13180 288 ne
rect 13180 261 13238 288
tri 13344 266 13374 296 ne
rect 12988 193 13044 227
rect 12988 159 12998 193
rect 13032 159 13044 193
rect 12988 127 13044 159
tri 13074 242 13090 258 se
rect 13090 242 13134 258
tri 13134 242 13150 258 sw
rect 13074 208 13150 242
rect 13074 174 13095 208
rect 13129 174 13150 208
rect 13074 173 13150 174
tri 13074 157 13090 173 ne
rect 13090 157 13134 173
tri 13134 157 13150 173 nw
rect 13180 227 13192 261
rect 13226 227 13238 261
rect 13180 193 13238 227
rect 13180 159 13192 193
rect 13226 159 13238 193
tri 13268 250 13284 266 se
rect 13284 250 13328 266
tri 13328 250 13344 266 sw
rect 13268 217 13344 250
rect 13268 183 13288 217
rect 13322 183 13344 217
rect 13268 181 13344 183
tri 13268 165 13284 181 ne
rect 13284 165 13328 181
tri 13328 165 13344 181 nw
rect 13374 261 13428 296
rect 13374 227 13386 261
rect 13420 227 13428 261
rect 13374 193 13428 227
tri 13044 127 13074 157 sw
tri 13150 127 13180 157 se
rect 13180 135 13238 159
tri 13238 135 13268 165 sw
tri 13344 135 13374 165 se
rect 13374 159 13386 193
rect 13420 159 13428 193
rect 13374 135 13428 159
rect 13180 127 13428 135
rect 12988 123 13428 127
rect 12988 89 12998 123
rect 13032 89 13192 123
rect 13226 89 13288 123
rect 13322 89 13386 123
rect 13420 89 13428 123
rect 12988 73 13428 89
rect 13654 333 13710 349
rect 13654 299 13664 333
rect 13698 299 13710 333
rect 13654 261 13710 299
rect 13740 333 14010 349
rect 13740 304 13761 333
tri 13740 288 13756 304 ne
rect 13756 299 13761 304
rect 13795 299 13858 333
rect 13892 312 14010 333
rect 13892 299 13994 312
rect 13756 296 13994 299
tri 13994 296 14010 312 nw
rect 14040 333 14096 349
rect 14040 299 14052 333
rect 14086 299 14096 333
rect 13756 288 13904 296
rect 13654 227 13664 261
rect 13698 227 13710 261
tri 13816 258 13846 288 ne
rect 13846 261 13904 288
tri 13904 266 13934 296 nw
rect 13654 193 13710 227
rect 13654 159 13664 193
rect 13698 159 13710 193
rect 13654 127 13710 159
tri 13740 242 13756 258 se
rect 13756 242 13800 258
tri 13800 242 13816 258 sw
rect 13740 208 13816 242
rect 13740 174 13761 208
rect 13795 174 13816 208
rect 13740 173 13816 174
tri 13740 157 13756 173 ne
rect 13756 157 13800 173
tri 13800 157 13816 173 nw
rect 13846 227 13858 261
rect 13892 227 13904 261
rect 13846 193 13904 227
rect 13846 159 13858 193
rect 13892 159 13904 193
tri 13934 250 13950 266 se
rect 13950 250 13994 266
tri 13994 250 14010 266 sw
rect 13934 217 14010 250
rect 13934 183 13955 217
rect 13989 183 14010 217
rect 13934 181 14010 183
tri 13934 165 13950 181 ne
rect 13950 165 13994 181
tri 13994 165 14010 181 nw
rect 14040 261 14096 299
rect 14040 227 14052 261
rect 14086 227 14096 261
rect 14040 193 14096 227
tri 13710 127 13740 157 sw
tri 13816 127 13846 157 se
rect 13846 135 13904 159
tri 13904 135 13934 165 sw
tri 14010 135 14040 165 se
rect 14040 159 14052 193
rect 14086 159 14096 193
rect 14040 135 14096 159
rect 13846 127 14096 135
rect 13654 123 14096 127
rect 13654 89 13664 123
rect 13698 89 13858 123
rect 13892 89 13955 123
rect 13989 89 14052 123
rect 14086 89 14096 123
rect 13654 73 14096 89
rect 14320 333 14376 349
rect 14320 299 14330 333
rect 14364 299 14376 333
rect 14320 261 14376 299
rect 14406 333 14570 349
rect 14406 304 14427 333
tri 14406 288 14422 304 ne
rect 14422 299 14427 304
rect 14461 299 14524 333
rect 14558 299 14570 333
rect 14422 288 14570 299
rect 14600 312 14762 349
tri 14600 296 14616 312 ne
rect 14616 296 14762 312
rect 14320 227 14330 261
rect 14364 227 14376 261
tri 14482 258 14512 288 ne
rect 14512 261 14570 288
tri 14676 266 14706 296 ne
rect 14320 193 14376 227
rect 14320 159 14330 193
rect 14364 159 14376 193
rect 14320 127 14376 159
tri 14406 242 14422 258 se
rect 14422 242 14466 258
tri 14466 242 14482 258 sw
rect 14406 208 14482 242
rect 14406 174 14427 208
rect 14461 174 14482 208
rect 14406 173 14482 174
tri 14406 157 14422 173 ne
rect 14422 157 14466 173
tri 14466 157 14482 173 nw
rect 14512 227 14524 261
rect 14558 227 14570 261
tri 14601 251 14616 266 se
rect 14616 251 14660 266
tri 14660 251 14675 266 sw
rect 14706 261 14762 296
rect 14512 193 14570 227
rect 14512 159 14524 193
rect 14558 159 14570 193
rect 14600 217 14676 251
rect 14600 183 14621 217
rect 14655 183 14676 217
rect 14600 181 14676 183
tri 14600 165 14616 181 ne
rect 14616 165 14660 181
tri 14660 165 14676 181 nw
rect 14706 227 14718 261
rect 14752 227 14762 261
rect 14706 193 14762 227
tri 14376 127 14406 157 sw
tri 14482 127 14512 157 se
rect 14512 135 14570 159
tri 14570 135 14600 165 sw
tri 14676 135 14706 165 se
rect 14706 159 14718 193
rect 14752 159 14762 193
rect 14706 135 14762 159
rect 14512 127 14762 135
rect 14320 123 14762 127
rect 14320 89 14330 123
rect 14364 89 14524 123
rect 14558 89 14621 123
rect 14655 89 14718 123
rect 14752 89 14762 123
rect 14320 73 14762 89
<< pdiff >>
rect 191 1366 247 1404
rect 191 1332 201 1366
rect 235 1332 247 1366
rect 191 1298 247 1332
rect 191 1264 201 1298
rect 235 1264 247 1298
rect 191 1230 247 1264
rect 191 1196 201 1230
rect 235 1196 247 1230
rect 191 1162 247 1196
rect 191 1128 201 1162
rect 235 1128 247 1162
rect 191 1093 247 1128
rect 191 1059 201 1093
rect 235 1059 247 1093
rect 191 1004 247 1059
rect 277 1366 335 1404
rect 277 1332 289 1366
rect 323 1332 335 1366
rect 277 1298 335 1332
rect 277 1264 289 1298
rect 323 1264 335 1298
rect 277 1230 335 1264
rect 277 1196 289 1230
rect 323 1196 335 1230
rect 277 1162 335 1196
rect 277 1128 289 1162
rect 323 1128 335 1162
rect 277 1093 335 1128
rect 277 1059 289 1093
rect 323 1059 335 1093
rect 277 1004 335 1059
rect 365 1366 423 1404
rect 365 1332 377 1366
rect 411 1332 423 1366
rect 365 1298 423 1332
rect 365 1264 377 1298
rect 411 1264 423 1298
rect 365 1230 423 1264
rect 365 1196 377 1230
rect 411 1196 423 1230
rect 365 1162 423 1196
rect 365 1128 377 1162
rect 411 1128 423 1162
rect 365 1004 423 1128
rect 453 1366 511 1404
rect 453 1332 465 1366
rect 499 1332 511 1366
rect 453 1298 511 1332
rect 453 1264 465 1298
rect 499 1264 511 1298
rect 453 1230 511 1264
rect 453 1196 465 1230
rect 499 1196 511 1230
rect 453 1162 511 1196
rect 453 1128 465 1162
rect 499 1128 511 1162
rect 453 1093 511 1128
rect 453 1059 465 1093
rect 499 1059 511 1093
rect 453 1004 511 1059
rect 541 1366 599 1404
rect 541 1332 553 1366
rect 587 1332 599 1366
rect 541 1298 599 1332
rect 541 1264 553 1298
rect 587 1264 599 1298
rect 541 1230 599 1264
rect 541 1196 553 1230
rect 587 1196 599 1230
rect 541 1162 599 1196
rect 541 1128 553 1162
rect 587 1128 599 1162
rect 541 1004 599 1128
rect 629 1366 687 1404
rect 629 1332 641 1366
rect 675 1332 687 1366
rect 629 1298 687 1332
rect 629 1264 641 1298
rect 675 1264 687 1298
rect 629 1230 687 1264
rect 629 1196 641 1230
rect 675 1196 687 1230
rect 629 1162 687 1196
rect 629 1128 641 1162
rect 675 1128 687 1162
rect 629 1093 687 1128
rect 629 1059 641 1093
rect 675 1059 687 1093
rect 629 1004 687 1059
rect 717 1366 771 1404
rect 717 1332 729 1366
rect 763 1332 771 1366
rect 717 1298 771 1332
rect 717 1264 729 1298
rect 763 1264 771 1298
rect 717 1230 771 1264
rect 717 1196 729 1230
rect 763 1196 771 1230
rect 717 1162 771 1196
rect 717 1128 729 1162
rect 763 1128 771 1162
rect 717 1004 771 1128
rect 1093 1366 1149 1404
rect 1093 1332 1103 1366
rect 1137 1332 1149 1366
rect 1093 1298 1149 1332
rect 1093 1264 1103 1298
rect 1137 1264 1149 1298
rect 1093 1230 1149 1264
rect 1093 1196 1103 1230
rect 1137 1196 1149 1230
rect 1093 1162 1149 1196
rect 1093 1128 1103 1162
rect 1137 1128 1149 1162
rect 1093 1093 1149 1128
rect 1093 1059 1103 1093
rect 1137 1059 1149 1093
rect 1093 1004 1149 1059
rect 1179 1366 1237 1404
rect 1179 1332 1191 1366
rect 1225 1332 1237 1366
rect 1179 1298 1237 1332
rect 1179 1264 1191 1298
rect 1225 1264 1237 1298
rect 1179 1230 1237 1264
rect 1179 1196 1191 1230
rect 1225 1196 1237 1230
rect 1179 1162 1237 1196
rect 1179 1128 1191 1162
rect 1225 1128 1237 1162
rect 1179 1093 1237 1128
rect 1179 1059 1191 1093
rect 1225 1059 1237 1093
rect 1179 1004 1237 1059
rect 1267 1366 1325 1404
rect 1267 1332 1279 1366
rect 1313 1332 1325 1366
rect 1267 1298 1325 1332
rect 1267 1264 1279 1298
rect 1313 1264 1325 1298
rect 1267 1230 1325 1264
rect 1267 1196 1279 1230
rect 1313 1196 1325 1230
rect 1267 1162 1325 1196
rect 1267 1128 1279 1162
rect 1313 1128 1325 1162
rect 1267 1004 1325 1128
rect 1355 1366 1413 1404
rect 1355 1332 1367 1366
rect 1401 1332 1413 1366
rect 1355 1298 1413 1332
rect 1355 1264 1367 1298
rect 1401 1264 1413 1298
rect 1355 1230 1413 1264
rect 1355 1196 1367 1230
rect 1401 1196 1413 1230
rect 1355 1162 1413 1196
rect 1355 1128 1367 1162
rect 1401 1128 1413 1162
rect 1355 1093 1413 1128
rect 1355 1059 1367 1093
rect 1401 1059 1413 1093
rect 1355 1004 1413 1059
rect 1443 1366 1497 1404
rect 1443 1332 1455 1366
rect 1489 1332 1497 1366
rect 1443 1298 1497 1332
rect 1443 1264 1455 1298
rect 1489 1264 1497 1298
rect 1443 1230 1497 1264
rect 1443 1196 1455 1230
rect 1489 1196 1497 1230
rect 1443 1162 1497 1196
rect 1443 1128 1455 1162
rect 1489 1128 1497 1162
rect 1443 1004 1497 1128
rect 1759 1366 1815 1404
rect 1759 1332 1769 1366
rect 1803 1332 1815 1366
rect 1759 1298 1815 1332
rect 1759 1264 1769 1298
rect 1803 1264 1815 1298
rect 1759 1230 1815 1264
rect 1759 1196 1769 1230
rect 1803 1196 1815 1230
rect 1759 1162 1815 1196
rect 1759 1128 1769 1162
rect 1803 1128 1815 1162
rect 1759 1093 1815 1128
rect 1759 1059 1769 1093
rect 1803 1059 1815 1093
rect 1759 1004 1815 1059
rect 1845 1366 1903 1404
rect 1845 1332 1857 1366
rect 1891 1332 1903 1366
rect 1845 1298 1903 1332
rect 1845 1264 1857 1298
rect 1891 1264 1903 1298
rect 1845 1230 1903 1264
rect 1845 1196 1857 1230
rect 1891 1196 1903 1230
rect 1845 1162 1903 1196
rect 1845 1128 1857 1162
rect 1891 1128 1903 1162
rect 1845 1093 1903 1128
rect 1845 1059 1857 1093
rect 1891 1059 1903 1093
rect 1845 1004 1903 1059
rect 1933 1366 1991 1404
rect 1933 1332 1945 1366
rect 1979 1332 1991 1366
rect 1933 1298 1991 1332
rect 1933 1264 1945 1298
rect 1979 1264 1991 1298
rect 1933 1230 1991 1264
rect 1933 1196 1945 1230
rect 1979 1196 1991 1230
rect 1933 1162 1991 1196
rect 1933 1128 1945 1162
rect 1979 1128 1991 1162
rect 1933 1004 1991 1128
rect 2021 1366 2079 1404
rect 2021 1332 2033 1366
rect 2067 1332 2079 1366
rect 2021 1298 2079 1332
rect 2021 1264 2033 1298
rect 2067 1264 2079 1298
rect 2021 1230 2079 1264
rect 2021 1196 2033 1230
rect 2067 1196 2079 1230
rect 2021 1162 2079 1196
rect 2021 1128 2033 1162
rect 2067 1128 2079 1162
rect 2021 1093 2079 1128
rect 2021 1059 2033 1093
rect 2067 1059 2079 1093
rect 2021 1004 2079 1059
rect 2109 1366 2163 1404
rect 2109 1332 2121 1366
rect 2155 1332 2163 1366
rect 2109 1298 2163 1332
rect 2109 1264 2121 1298
rect 2155 1264 2163 1298
rect 2109 1230 2163 1264
rect 2109 1196 2121 1230
rect 2155 1196 2163 1230
rect 2109 1162 2163 1196
rect 2109 1128 2121 1162
rect 2155 1128 2163 1162
rect 2109 1004 2163 1128
rect 2425 1366 2481 1404
rect 2425 1332 2435 1366
rect 2469 1332 2481 1366
rect 2425 1298 2481 1332
rect 2425 1264 2435 1298
rect 2469 1264 2481 1298
rect 2425 1230 2481 1264
rect 2425 1196 2435 1230
rect 2469 1196 2481 1230
rect 2425 1162 2481 1196
rect 2425 1128 2435 1162
rect 2469 1128 2481 1162
rect 2425 1093 2481 1128
rect 2425 1059 2435 1093
rect 2469 1059 2481 1093
rect 2425 1004 2481 1059
rect 2511 1366 2569 1404
rect 2511 1332 2523 1366
rect 2557 1332 2569 1366
rect 2511 1298 2569 1332
rect 2511 1264 2523 1298
rect 2557 1264 2569 1298
rect 2511 1230 2569 1264
rect 2511 1196 2523 1230
rect 2557 1196 2569 1230
rect 2511 1162 2569 1196
rect 2511 1128 2523 1162
rect 2557 1128 2569 1162
rect 2511 1093 2569 1128
rect 2511 1059 2523 1093
rect 2557 1059 2569 1093
rect 2511 1004 2569 1059
rect 2599 1366 2657 1404
rect 2599 1332 2611 1366
rect 2645 1332 2657 1366
rect 2599 1298 2657 1332
rect 2599 1264 2611 1298
rect 2645 1264 2657 1298
rect 2599 1230 2657 1264
rect 2599 1196 2611 1230
rect 2645 1196 2657 1230
rect 2599 1162 2657 1196
rect 2599 1128 2611 1162
rect 2645 1128 2657 1162
rect 2599 1004 2657 1128
rect 2687 1366 2745 1404
rect 2687 1332 2699 1366
rect 2733 1332 2745 1366
rect 2687 1298 2745 1332
rect 2687 1264 2699 1298
rect 2733 1264 2745 1298
rect 2687 1230 2745 1264
rect 2687 1196 2699 1230
rect 2733 1196 2745 1230
rect 2687 1162 2745 1196
rect 2687 1128 2699 1162
rect 2733 1128 2745 1162
rect 2687 1093 2745 1128
rect 2687 1059 2699 1093
rect 2733 1059 2745 1093
rect 2687 1004 2745 1059
rect 2775 1366 2829 1404
rect 2775 1332 2787 1366
rect 2821 1332 2829 1366
rect 2775 1298 2829 1332
rect 2775 1264 2787 1298
rect 2821 1264 2829 1298
rect 2775 1230 2829 1264
rect 2775 1196 2787 1230
rect 2821 1196 2829 1230
rect 2775 1162 2829 1196
rect 2775 1128 2787 1162
rect 2821 1128 2829 1162
rect 2775 1004 2829 1128
rect 3091 1366 3147 1404
rect 3091 1332 3101 1366
rect 3135 1332 3147 1366
rect 3091 1298 3147 1332
rect 3091 1264 3101 1298
rect 3135 1264 3147 1298
rect 3091 1230 3147 1264
rect 3091 1196 3101 1230
rect 3135 1196 3147 1230
rect 3091 1162 3147 1196
rect 3091 1128 3101 1162
rect 3135 1128 3147 1162
rect 3091 1093 3147 1128
rect 3091 1059 3101 1093
rect 3135 1059 3147 1093
rect 3091 1004 3147 1059
rect 3177 1366 3235 1404
rect 3177 1332 3189 1366
rect 3223 1332 3235 1366
rect 3177 1298 3235 1332
rect 3177 1264 3189 1298
rect 3223 1264 3235 1298
rect 3177 1230 3235 1264
rect 3177 1196 3189 1230
rect 3223 1196 3235 1230
rect 3177 1162 3235 1196
rect 3177 1128 3189 1162
rect 3223 1128 3235 1162
rect 3177 1093 3235 1128
rect 3177 1059 3189 1093
rect 3223 1059 3235 1093
rect 3177 1004 3235 1059
rect 3265 1366 3323 1404
rect 3265 1332 3277 1366
rect 3311 1332 3323 1366
rect 3265 1298 3323 1332
rect 3265 1264 3277 1298
rect 3311 1264 3323 1298
rect 3265 1230 3323 1264
rect 3265 1196 3277 1230
rect 3311 1196 3323 1230
rect 3265 1162 3323 1196
rect 3265 1128 3277 1162
rect 3311 1128 3323 1162
rect 3265 1004 3323 1128
rect 3353 1366 3411 1404
rect 3353 1332 3365 1366
rect 3399 1332 3411 1366
rect 3353 1298 3411 1332
rect 3353 1264 3365 1298
rect 3399 1264 3411 1298
rect 3353 1230 3411 1264
rect 3353 1196 3365 1230
rect 3399 1196 3411 1230
rect 3353 1162 3411 1196
rect 3353 1128 3365 1162
rect 3399 1128 3411 1162
rect 3353 1093 3411 1128
rect 3353 1059 3365 1093
rect 3399 1059 3411 1093
rect 3353 1004 3411 1059
rect 3441 1366 3495 1404
rect 3441 1332 3453 1366
rect 3487 1332 3495 1366
rect 3441 1298 3495 1332
rect 3441 1264 3453 1298
rect 3487 1264 3495 1298
rect 3441 1230 3495 1264
rect 3441 1196 3453 1230
rect 3487 1196 3495 1230
rect 3441 1162 3495 1196
rect 3441 1128 3453 1162
rect 3487 1128 3495 1162
rect 3441 1004 3495 1128
rect 3757 1366 3813 1404
rect 3757 1332 3767 1366
rect 3801 1332 3813 1366
rect 3757 1298 3813 1332
rect 3757 1264 3767 1298
rect 3801 1264 3813 1298
rect 3757 1230 3813 1264
rect 3757 1196 3767 1230
rect 3801 1196 3813 1230
rect 3757 1162 3813 1196
rect 3757 1128 3767 1162
rect 3801 1128 3813 1162
rect 3757 1093 3813 1128
rect 3757 1059 3767 1093
rect 3801 1059 3813 1093
rect 3757 1004 3813 1059
rect 3843 1366 3901 1404
rect 3843 1332 3855 1366
rect 3889 1332 3901 1366
rect 3843 1298 3901 1332
rect 3843 1264 3855 1298
rect 3889 1264 3901 1298
rect 3843 1230 3901 1264
rect 3843 1196 3855 1230
rect 3889 1196 3901 1230
rect 3843 1162 3901 1196
rect 3843 1128 3855 1162
rect 3889 1128 3901 1162
rect 3843 1093 3901 1128
rect 3843 1059 3855 1093
rect 3889 1059 3901 1093
rect 3843 1004 3901 1059
rect 3931 1366 3989 1404
rect 3931 1332 3943 1366
rect 3977 1332 3989 1366
rect 3931 1298 3989 1332
rect 3931 1264 3943 1298
rect 3977 1264 3989 1298
rect 3931 1230 3989 1264
rect 3931 1196 3943 1230
rect 3977 1196 3989 1230
rect 3931 1162 3989 1196
rect 3931 1128 3943 1162
rect 3977 1128 3989 1162
rect 3931 1004 3989 1128
rect 4019 1366 4077 1404
rect 4019 1332 4031 1366
rect 4065 1332 4077 1366
rect 4019 1298 4077 1332
rect 4019 1264 4031 1298
rect 4065 1264 4077 1298
rect 4019 1230 4077 1264
rect 4019 1196 4031 1230
rect 4065 1196 4077 1230
rect 4019 1162 4077 1196
rect 4019 1128 4031 1162
rect 4065 1128 4077 1162
rect 4019 1093 4077 1128
rect 4019 1059 4031 1093
rect 4065 1059 4077 1093
rect 4019 1004 4077 1059
rect 4107 1366 4161 1404
rect 4107 1332 4119 1366
rect 4153 1332 4161 1366
rect 4107 1298 4161 1332
rect 4107 1264 4119 1298
rect 4153 1264 4161 1298
rect 4107 1230 4161 1264
rect 4107 1196 4119 1230
rect 4153 1196 4161 1230
rect 4107 1162 4161 1196
rect 4107 1128 4119 1162
rect 4153 1128 4161 1162
rect 4107 1004 4161 1128
rect 4483 1366 4539 1404
rect 4483 1332 4493 1366
rect 4527 1332 4539 1366
rect 4483 1298 4539 1332
rect 4483 1264 4493 1298
rect 4527 1264 4539 1298
rect 4483 1230 4539 1264
rect 4483 1196 4493 1230
rect 4527 1196 4539 1230
rect 4483 1162 4539 1196
rect 4483 1128 4493 1162
rect 4527 1128 4539 1162
rect 4483 1093 4539 1128
rect 4483 1059 4493 1093
rect 4527 1059 4539 1093
rect 4483 1004 4539 1059
rect 4569 1366 4627 1404
rect 4569 1332 4581 1366
rect 4615 1332 4627 1366
rect 4569 1298 4627 1332
rect 4569 1264 4581 1298
rect 4615 1264 4627 1298
rect 4569 1230 4627 1264
rect 4569 1196 4581 1230
rect 4615 1196 4627 1230
rect 4569 1162 4627 1196
rect 4569 1128 4581 1162
rect 4615 1128 4627 1162
rect 4569 1093 4627 1128
rect 4569 1059 4581 1093
rect 4615 1059 4627 1093
rect 4569 1004 4627 1059
rect 4657 1366 4715 1404
rect 4657 1332 4669 1366
rect 4703 1332 4715 1366
rect 4657 1298 4715 1332
rect 4657 1264 4669 1298
rect 4703 1264 4715 1298
rect 4657 1230 4715 1264
rect 4657 1196 4669 1230
rect 4703 1196 4715 1230
rect 4657 1162 4715 1196
rect 4657 1128 4669 1162
rect 4703 1128 4715 1162
rect 4657 1004 4715 1128
rect 4745 1366 4803 1404
rect 4745 1332 4757 1366
rect 4791 1332 4803 1366
rect 4745 1298 4803 1332
rect 4745 1264 4757 1298
rect 4791 1264 4803 1298
rect 4745 1230 4803 1264
rect 4745 1196 4757 1230
rect 4791 1196 4803 1230
rect 4745 1162 4803 1196
rect 4745 1128 4757 1162
rect 4791 1128 4803 1162
rect 4745 1093 4803 1128
rect 4745 1059 4757 1093
rect 4791 1059 4803 1093
rect 4745 1004 4803 1059
rect 4833 1366 4891 1404
rect 4833 1332 4845 1366
rect 4879 1332 4891 1366
rect 4833 1298 4891 1332
rect 4833 1264 4845 1298
rect 4879 1264 4891 1298
rect 4833 1230 4891 1264
rect 4833 1196 4845 1230
rect 4879 1196 4891 1230
rect 4833 1162 4891 1196
rect 4833 1128 4845 1162
rect 4879 1128 4891 1162
rect 4833 1004 4891 1128
rect 4921 1366 4979 1404
rect 4921 1332 4933 1366
rect 4967 1332 4979 1366
rect 4921 1298 4979 1332
rect 4921 1264 4933 1298
rect 4967 1264 4979 1298
rect 4921 1230 4979 1264
rect 4921 1196 4933 1230
rect 4967 1196 4979 1230
rect 4921 1162 4979 1196
rect 4921 1128 4933 1162
rect 4967 1128 4979 1162
rect 4921 1093 4979 1128
rect 4921 1059 4933 1093
rect 4967 1059 4979 1093
rect 4921 1004 4979 1059
rect 5009 1366 5063 1404
rect 5009 1332 5021 1366
rect 5055 1332 5063 1366
rect 5009 1298 5063 1332
rect 5009 1264 5021 1298
rect 5055 1264 5063 1298
rect 5009 1230 5063 1264
rect 5009 1196 5021 1230
rect 5055 1196 5063 1230
rect 5009 1162 5063 1196
rect 5009 1128 5021 1162
rect 5055 1128 5063 1162
rect 5009 1004 5063 1128
rect 5385 1366 5441 1404
rect 5385 1332 5395 1366
rect 5429 1332 5441 1366
rect 5385 1298 5441 1332
rect 5385 1264 5395 1298
rect 5429 1264 5441 1298
rect 5385 1230 5441 1264
rect 5385 1196 5395 1230
rect 5429 1196 5441 1230
rect 5385 1162 5441 1196
rect 5385 1128 5395 1162
rect 5429 1128 5441 1162
rect 5385 1093 5441 1128
rect 5385 1059 5395 1093
rect 5429 1059 5441 1093
rect 5385 1004 5441 1059
rect 5471 1366 5529 1404
rect 5471 1332 5483 1366
rect 5517 1332 5529 1366
rect 5471 1298 5529 1332
rect 5471 1264 5483 1298
rect 5517 1264 5529 1298
rect 5471 1230 5529 1264
rect 5471 1196 5483 1230
rect 5517 1196 5529 1230
rect 5471 1162 5529 1196
rect 5471 1128 5483 1162
rect 5517 1128 5529 1162
rect 5471 1093 5529 1128
rect 5471 1059 5483 1093
rect 5517 1059 5529 1093
rect 5471 1004 5529 1059
rect 5559 1366 5617 1404
rect 5559 1332 5571 1366
rect 5605 1332 5617 1366
rect 5559 1298 5617 1332
rect 5559 1264 5571 1298
rect 5605 1264 5617 1298
rect 5559 1230 5617 1264
rect 5559 1196 5571 1230
rect 5605 1196 5617 1230
rect 5559 1162 5617 1196
rect 5559 1128 5571 1162
rect 5605 1128 5617 1162
rect 5559 1004 5617 1128
rect 5647 1366 5705 1404
rect 5647 1332 5659 1366
rect 5693 1332 5705 1366
rect 5647 1298 5705 1332
rect 5647 1264 5659 1298
rect 5693 1264 5705 1298
rect 5647 1230 5705 1264
rect 5647 1196 5659 1230
rect 5693 1196 5705 1230
rect 5647 1162 5705 1196
rect 5647 1128 5659 1162
rect 5693 1128 5705 1162
rect 5647 1093 5705 1128
rect 5647 1059 5659 1093
rect 5693 1059 5705 1093
rect 5647 1004 5705 1059
rect 5735 1366 5789 1404
rect 5735 1332 5747 1366
rect 5781 1332 5789 1366
rect 5735 1298 5789 1332
rect 5735 1264 5747 1298
rect 5781 1264 5789 1298
rect 5735 1230 5789 1264
rect 5735 1196 5747 1230
rect 5781 1196 5789 1230
rect 5735 1162 5789 1196
rect 5735 1128 5747 1162
rect 5781 1128 5789 1162
rect 5735 1004 5789 1128
rect 6051 1366 6107 1404
rect 6051 1332 6061 1366
rect 6095 1332 6107 1366
rect 6051 1298 6107 1332
rect 6051 1264 6061 1298
rect 6095 1264 6107 1298
rect 6051 1230 6107 1264
rect 6051 1196 6061 1230
rect 6095 1196 6107 1230
rect 6051 1162 6107 1196
rect 6051 1128 6061 1162
rect 6095 1128 6107 1162
rect 6051 1093 6107 1128
rect 6051 1059 6061 1093
rect 6095 1059 6107 1093
rect 6051 1004 6107 1059
rect 6137 1366 6195 1404
rect 6137 1332 6149 1366
rect 6183 1332 6195 1366
rect 6137 1298 6195 1332
rect 6137 1264 6149 1298
rect 6183 1264 6195 1298
rect 6137 1230 6195 1264
rect 6137 1196 6149 1230
rect 6183 1196 6195 1230
rect 6137 1162 6195 1196
rect 6137 1128 6149 1162
rect 6183 1128 6195 1162
rect 6137 1093 6195 1128
rect 6137 1059 6149 1093
rect 6183 1059 6195 1093
rect 6137 1004 6195 1059
rect 6225 1366 6283 1404
rect 6225 1332 6237 1366
rect 6271 1332 6283 1366
rect 6225 1298 6283 1332
rect 6225 1264 6237 1298
rect 6271 1264 6283 1298
rect 6225 1230 6283 1264
rect 6225 1196 6237 1230
rect 6271 1196 6283 1230
rect 6225 1162 6283 1196
rect 6225 1128 6237 1162
rect 6271 1128 6283 1162
rect 6225 1004 6283 1128
rect 6313 1366 6371 1404
rect 6313 1332 6325 1366
rect 6359 1332 6371 1366
rect 6313 1298 6371 1332
rect 6313 1264 6325 1298
rect 6359 1264 6371 1298
rect 6313 1230 6371 1264
rect 6313 1196 6325 1230
rect 6359 1196 6371 1230
rect 6313 1162 6371 1196
rect 6313 1128 6325 1162
rect 6359 1128 6371 1162
rect 6313 1093 6371 1128
rect 6313 1059 6325 1093
rect 6359 1059 6371 1093
rect 6313 1004 6371 1059
rect 6401 1366 6455 1404
rect 6401 1332 6413 1366
rect 6447 1332 6455 1366
rect 6401 1298 6455 1332
rect 6401 1264 6413 1298
rect 6447 1264 6455 1298
rect 6401 1230 6455 1264
rect 6401 1196 6413 1230
rect 6447 1196 6455 1230
rect 6401 1162 6455 1196
rect 6401 1128 6413 1162
rect 6447 1128 6455 1162
rect 6401 1004 6455 1128
rect 6717 1366 6773 1404
rect 6717 1332 6727 1366
rect 6761 1332 6773 1366
rect 6717 1298 6773 1332
rect 6717 1264 6727 1298
rect 6761 1264 6773 1298
rect 6717 1230 6773 1264
rect 6717 1196 6727 1230
rect 6761 1196 6773 1230
rect 6717 1162 6773 1196
rect 6717 1128 6727 1162
rect 6761 1128 6773 1162
rect 6717 1093 6773 1128
rect 6717 1059 6727 1093
rect 6761 1059 6773 1093
rect 6717 1004 6773 1059
rect 6803 1366 6861 1404
rect 6803 1332 6815 1366
rect 6849 1332 6861 1366
rect 6803 1298 6861 1332
rect 6803 1264 6815 1298
rect 6849 1264 6861 1298
rect 6803 1230 6861 1264
rect 6803 1196 6815 1230
rect 6849 1196 6861 1230
rect 6803 1162 6861 1196
rect 6803 1128 6815 1162
rect 6849 1128 6861 1162
rect 6803 1093 6861 1128
rect 6803 1059 6815 1093
rect 6849 1059 6861 1093
rect 6803 1004 6861 1059
rect 6891 1366 6949 1404
rect 6891 1332 6903 1366
rect 6937 1332 6949 1366
rect 6891 1298 6949 1332
rect 6891 1264 6903 1298
rect 6937 1264 6949 1298
rect 6891 1230 6949 1264
rect 6891 1196 6903 1230
rect 6937 1196 6949 1230
rect 6891 1162 6949 1196
rect 6891 1128 6903 1162
rect 6937 1128 6949 1162
rect 6891 1004 6949 1128
rect 6979 1366 7037 1404
rect 6979 1332 6991 1366
rect 7025 1332 7037 1366
rect 6979 1298 7037 1332
rect 6979 1264 6991 1298
rect 7025 1264 7037 1298
rect 6979 1230 7037 1264
rect 6979 1196 6991 1230
rect 7025 1196 7037 1230
rect 6979 1162 7037 1196
rect 6979 1128 6991 1162
rect 7025 1128 7037 1162
rect 6979 1093 7037 1128
rect 6979 1059 6991 1093
rect 7025 1059 7037 1093
rect 6979 1004 7037 1059
rect 7067 1366 7121 1404
rect 7067 1332 7079 1366
rect 7113 1332 7121 1366
rect 7067 1298 7121 1332
rect 7067 1264 7079 1298
rect 7113 1264 7121 1298
rect 7067 1230 7121 1264
rect 7067 1196 7079 1230
rect 7113 1196 7121 1230
rect 7067 1162 7121 1196
rect 7067 1128 7079 1162
rect 7113 1128 7121 1162
rect 7067 1004 7121 1128
rect 7383 1366 7439 1404
rect 7383 1332 7393 1366
rect 7427 1332 7439 1366
rect 7383 1298 7439 1332
rect 7383 1264 7393 1298
rect 7427 1264 7439 1298
rect 7383 1230 7439 1264
rect 7383 1196 7393 1230
rect 7427 1196 7439 1230
rect 7383 1162 7439 1196
rect 7383 1128 7393 1162
rect 7427 1128 7439 1162
rect 7383 1093 7439 1128
rect 7383 1059 7393 1093
rect 7427 1059 7439 1093
rect 7383 1004 7439 1059
rect 7469 1366 7527 1404
rect 7469 1332 7481 1366
rect 7515 1332 7527 1366
rect 7469 1298 7527 1332
rect 7469 1264 7481 1298
rect 7515 1264 7527 1298
rect 7469 1230 7527 1264
rect 7469 1196 7481 1230
rect 7515 1196 7527 1230
rect 7469 1162 7527 1196
rect 7469 1128 7481 1162
rect 7515 1128 7527 1162
rect 7469 1093 7527 1128
rect 7469 1059 7481 1093
rect 7515 1059 7527 1093
rect 7469 1004 7527 1059
rect 7557 1366 7615 1404
rect 7557 1332 7569 1366
rect 7603 1332 7615 1366
rect 7557 1298 7615 1332
rect 7557 1264 7569 1298
rect 7603 1264 7615 1298
rect 7557 1230 7615 1264
rect 7557 1196 7569 1230
rect 7603 1196 7615 1230
rect 7557 1162 7615 1196
rect 7557 1128 7569 1162
rect 7603 1128 7615 1162
rect 7557 1004 7615 1128
rect 7645 1366 7703 1404
rect 7645 1332 7657 1366
rect 7691 1332 7703 1366
rect 7645 1298 7703 1332
rect 7645 1264 7657 1298
rect 7691 1264 7703 1298
rect 7645 1230 7703 1264
rect 7645 1196 7657 1230
rect 7691 1196 7703 1230
rect 7645 1162 7703 1196
rect 7645 1128 7657 1162
rect 7691 1128 7703 1162
rect 7645 1093 7703 1128
rect 7645 1059 7657 1093
rect 7691 1059 7703 1093
rect 7645 1004 7703 1059
rect 7733 1366 7787 1404
rect 7733 1332 7745 1366
rect 7779 1332 7787 1366
rect 7733 1298 7787 1332
rect 7733 1264 7745 1298
rect 7779 1264 7787 1298
rect 7733 1230 7787 1264
rect 7733 1196 7745 1230
rect 7779 1196 7787 1230
rect 7733 1162 7787 1196
rect 7733 1128 7745 1162
rect 7779 1128 7787 1162
rect 7733 1004 7787 1128
rect 8049 1366 8105 1404
rect 8049 1332 8059 1366
rect 8093 1332 8105 1366
rect 8049 1298 8105 1332
rect 8049 1264 8059 1298
rect 8093 1264 8105 1298
rect 8049 1230 8105 1264
rect 8049 1196 8059 1230
rect 8093 1196 8105 1230
rect 8049 1162 8105 1196
rect 8049 1128 8059 1162
rect 8093 1128 8105 1162
rect 8049 1093 8105 1128
rect 8049 1059 8059 1093
rect 8093 1059 8105 1093
rect 8049 1004 8105 1059
rect 8135 1366 8193 1404
rect 8135 1332 8147 1366
rect 8181 1332 8193 1366
rect 8135 1298 8193 1332
rect 8135 1264 8147 1298
rect 8181 1264 8193 1298
rect 8135 1230 8193 1264
rect 8135 1196 8147 1230
rect 8181 1196 8193 1230
rect 8135 1162 8193 1196
rect 8135 1128 8147 1162
rect 8181 1128 8193 1162
rect 8135 1093 8193 1128
rect 8135 1059 8147 1093
rect 8181 1059 8193 1093
rect 8135 1004 8193 1059
rect 8223 1366 8281 1404
rect 8223 1332 8235 1366
rect 8269 1332 8281 1366
rect 8223 1298 8281 1332
rect 8223 1264 8235 1298
rect 8269 1264 8281 1298
rect 8223 1230 8281 1264
rect 8223 1196 8235 1230
rect 8269 1196 8281 1230
rect 8223 1162 8281 1196
rect 8223 1128 8235 1162
rect 8269 1128 8281 1162
rect 8223 1004 8281 1128
rect 8311 1366 8369 1404
rect 8311 1332 8323 1366
rect 8357 1332 8369 1366
rect 8311 1298 8369 1332
rect 8311 1264 8323 1298
rect 8357 1264 8369 1298
rect 8311 1230 8369 1264
rect 8311 1196 8323 1230
rect 8357 1196 8369 1230
rect 8311 1162 8369 1196
rect 8311 1128 8323 1162
rect 8357 1128 8369 1162
rect 8311 1093 8369 1128
rect 8311 1059 8323 1093
rect 8357 1059 8369 1093
rect 8311 1004 8369 1059
rect 8399 1366 8453 1404
rect 8399 1332 8411 1366
rect 8445 1332 8453 1366
rect 8399 1298 8453 1332
rect 8399 1264 8411 1298
rect 8445 1264 8453 1298
rect 8399 1230 8453 1264
rect 8399 1196 8411 1230
rect 8445 1196 8453 1230
rect 8399 1162 8453 1196
rect 8399 1128 8411 1162
rect 8445 1128 8453 1162
rect 8399 1004 8453 1128
rect 8775 1366 8831 1404
rect 8775 1332 8785 1366
rect 8819 1332 8831 1366
rect 8775 1298 8831 1332
rect 8775 1264 8785 1298
rect 8819 1264 8831 1298
rect 8775 1230 8831 1264
rect 8775 1196 8785 1230
rect 8819 1196 8831 1230
rect 8775 1162 8831 1196
rect 8775 1128 8785 1162
rect 8819 1128 8831 1162
rect 8775 1093 8831 1128
rect 8775 1059 8785 1093
rect 8819 1059 8831 1093
rect 8775 1004 8831 1059
rect 8861 1366 8919 1404
rect 8861 1332 8873 1366
rect 8907 1332 8919 1366
rect 8861 1298 8919 1332
rect 8861 1264 8873 1298
rect 8907 1264 8919 1298
rect 8861 1230 8919 1264
rect 8861 1196 8873 1230
rect 8907 1196 8919 1230
rect 8861 1162 8919 1196
rect 8861 1128 8873 1162
rect 8907 1128 8919 1162
rect 8861 1093 8919 1128
rect 8861 1059 8873 1093
rect 8907 1059 8919 1093
rect 8861 1004 8919 1059
rect 8949 1366 9007 1404
rect 8949 1332 8961 1366
rect 8995 1332 9007 1366
rect 8949 1298 9007 1332
rect 8949 1264 8961 1298
rect 8995 1264 9007 1298
rect 8949 1230 9007 1264
rect 8949 1196 8961 1230
rect 8995 1196 9007 1230
rect 8949 1162 9007 1196
rect 8949 1128 8961 1162
rect 8995 1128 9007 1162
rect 8949 1004 9007 1128
rect 9037 1366 9095 1404
rect 9037 1332 9049 1366
rect 9083 1332 9095 1366
rect 9037 1298 9095 1332
rect 9037 1264 9049 1298
rect 9083 1264 9095 1298
rect 9037 1230 9095 1264
rect 9037 1196 9049 1230
rect 9083 1196 9095 1230
rect 9037 1162 9095 1196
rect 9037 1128 9049 1162
rect 9083 1128 9095 1162
rect 9037 1093 9095 1128
rect 9037 1059 9049 1093
rect 9083 1059 9095 1093
rect 9037 1004 9095 1059
rect 9125 1366 9183 1404
rect 9125 1332 9137 1366
rect 9171 1332 9183 1366
rect 9125 1298 9183 1332
rect 9125 1264 9137 1298
rect 9171 1264 9183 1298
rect 9125 1230 9183 1264
rect 9125 1196 9137 1230
rect 9171 1196 9183 1230
rect 9125 1162 9183 1196
rect 9125 1128 9137 1162
rect 9171 1128 9183 1162
rect 9125 1004 9183 1128
rect 9213 1366 9271 1404
rect 9213 1332 9225 1366
rect 9259 1332 9271 1366
rect 9213 1298 9271 1332
rect 9213 1264 9225 1298
rect 9259 1264 9271 1298
rect 9213 1230 9271 1264
rect 9213 1196 9225 1230
rect 9259 1196 9271 1230
rect 9213 1162 9271 1196
rect 9213 1128 9225 1162
rect 9259 1128 9271 1162
rect 9213 1093 9271 1128
rect 9213 1059 9225 1093
rect 9259 1059 9271 1093
rect 9213 1004 9271 1059
rect 9301 1366 9355 1404
rect 9301 1332 9313 1366
rect 9347 1332 9355 1366
rect 9301 1298 9355 1332
rect 9301 1264 9313 1298
rect 9347 1264 9355 1298
rect 9301 1230 9355 1264
rect 9301 1196 9313 1230
rect 9347 1196 9355 1230
rect 9301 1162 9355 1196
rect 9301 1128 9313 1162
rect 9347 1128 9355 1162
rect 9301 1004 9355 1128
rect 9677 1366 9733 1404
rect 9677 1332 9687 1366
rect 9721 1332 9733 1366
rect 9677 1298 9733 1332
rect 9677 1264 9687 1298
rect 9721 1264 9733 1298
rect 9677 1230 9733 1264
rect 9677 1196 9687 1230
rect 9721 1196 9733 1230
rect 9677 1162 9733 1196
rect 9677 1128 9687 1162
rect 9721 1128 9733 1162
rect 9677 1093 9733 1128
rect 9677 1059 9687 1093
rect 9721 1059 9733 1093
rect 9677 1004 9733 1059
rect 9763 1366 9821 1404
rect 9763 1332 9775 1366
rect 9809 1332 9821 1366
rect 9763 1298 9821 1332
rect 9763 1264 9775 1298
rect 9809 1264 9821 1298
rect 9763 1230 9821 1264
rect 9763 1196 9775 1230
rect 9809 1196 9821 1230
rect 9763 1162 9821 1196
rect 9763 1128 9775 1162
rect 9809 1128 9821 1162
rect 9763 1093 9821 1128
rect 9763 1059 9775 1093
rect 9809 1059 9821 1093
rect 9763 1004 9821 1059
rect 9851 1366 9909 1404
rect 9851 1332 9863 1366
rect 9897 1332 9909 1366
rect 9851 1298 9909 1332
rect 9851 1264 9863 1298
rect 9897 1264 9909 1298
rect 9851 1230 9909 1264
rect 9851 1196 9863 1230
rect 9897 1196 9909 1230
rect 9851 1162 9909 1196
rect 9851 1128 9863 1162
rect 9897 1128 9909 1162
rect 9851 1004 9909 1128
rect 9939 1366 9997 1404
rect 9939 1332 9951 1366
rect 9985 1332 9997 1366
rect 9939 1298 9997 1332
rect 9939 1264 9951 1298
rect 9985 1264 9997 1298
rect 9939 1230 9997 1264
rect 9939 1196 9951 1230
rect 9985 1196 9997 1230
rect 9939 1162 9997 1196
rect 9939 1128 9951 1162
rect 9985 1128 9997 1162
rect 9939 1093 9997 1128
rect 9939 1059 9951 1093
rect 9985 1059 9997 1093
rect 9939 1004 9997 1059
rect 10027 1366 10081 1404
rect 10027 1332 10039 1366
rect 10073 1332 10081 1366
rect 10027 1298 10081 1332
rect 10027 1264 10039 1298
rect 10073 1264 10081 1298
rect 10027 1230 10081 1264
rect 10027 1196 10039 1230
rect 10073 1196 10081 1230
rect 10027 1162 10081 1196
rect 10027 1128 10039 1162
rect 10073 1128 10081 1162
rect 10027 1004 10081 1128
rect 10343 1366 10399 1404
rect 10343 1332 10353 1366
rect 10387 1332 10399 1366
rect 10343 1298 10399 1332
rect 10343 1264 10353 1298
rect 10387 1264 10399 1298
rect 10343 1230 10399 1264
rect 10343 1196 10353 1230
rect 10387 1196 10399 1230
rect 10343 1162 10399 1196
rect 10343 1128 10353 1162
rect 10387 1128 10399 1162
rect 10343 1093 10399 1128
rect 10343 1059 10353 1093
rect 10387 1059 10399 1093
rect 10343 1004 10399 1059
rect 10429 1366 10487 1404
rect 10429 1332 10441 1366
rect 10475 1332 10487 1366
rect 10429 1298 10487 1332
rect 10429 1264 10441 1298
rect 10475 1264 10487 1298
rect 10429 1230 10487 1264
rect 10429 1196 10441 1230
rect 10475 1196 10487 1230
rect 10429 1162 10487 1196
rect 10429 1128 10441 1162
rect 10475 1128 10487 1162
rect 10429 1093 10487 1128
rect 10429 1059 10441 1093
rect 10475 1059 10487 1093
rect 10429 1004 10487 1059
rect 10517 1366 10575 1404
rect 10517 1332 10529 1366
rect 10563 1332 10575 1366
rect 10517 1298 10575 1332
rect 10517 1264 10529 1298
rect 10563 1264 10575 1298
rect 10517 1230 10575 1264
rect 10517 1196 10529 1230
rect 10563 1196 10575 1230
rect 10517 1162 10575 1196
rect 10517 1128 10529 1162
rect 10563 1128 10575 1162
rect 10517 1004 10575 1128
rect 10605 1366 10663 1404
rect 10605 1332 10617 1366
rect 10651 1332 10663 1366
rect 10605 1298 10663 1332
rect 10605 1264 10617 1298
rect 10651 1264 10663 1298
rect 10605 1230 10663 1264
rect 10605 1196 10617 1230
rect 10651 1196 10663 1230
rect 10605 1162 10663 1196
rect 10605 1128 10617 1162
rect 10651 1128 10663 1162
rect 10605 1093 10663 1128
rect 10605 1059 10617 1093
rect 10651 1059 10663 1093
rect 10605 1004 10663 1059
rect 10693 1366 10747 1404
rect 10693 1332 10705 1366
rect 10739 1332 10747 1366
rect 10693 1298 10747 1332
rect 10693 1264 10705 1298
rect 10739 1264 10747 1298
rect 10693 1230 10747 1264
rect 10693 1196 10705 1230
rect 10739 1196 10747 1230
rect 10693 1162 10747 1196
rect 10693 1128 10705 1162
rect 10739 1128 10747 1162
rect 10693 1004 10747 1128
rect 11009 1366 11065 1404
rect 11009 1332 11019 1366
rect 11053 1332 11065 1366
rect 11009 1298 11065 1332
rect 11009 1264 11019 1298
rect 11053 1264 11065 1298
rect 11009 1230 11065 1264
rect 11009 1196 11019 1230
rect 11053 1196 11065 1230
rect 11009 1162 11065 1196
rect 11009 1128 11019 1162
rect 11053 1128 11065 1162
rect 11009 1093 11065 1128
rect 11009 1059 11019 1093
rect 11053 1059 11065 1093
rect 11009 1004 11065 1059
rect 11095 1366 11153 1404
rect 11095 1332 11107 1366
rect 11141 1332 11153 1366
rect 11095 1298 11153 1332
rect 11095 1264 11107 1298
rect 11141 1264 11153 1298
rect 11095 1230 11153 1264
rect 11095 1196 11107 1230
rect 11141 1196 11153 1230
rect 11095 1162 11153 1196
rect 11095 1128 11107 1162
rect 11141 1128 11153 1162
rect 11095 1093 11153 1128
rect 11095 1059 11107 1093
rect 11141 1059 11153 1093
rect 11095 1004 11153 1059
rect 11183 1366 11241 1404
rect 11183 1332 11195 1366
rect 11229 1332 11241 1366
rect 11183 1298 11241 1332
rect 11183 1264 11195 1298
rect 11229 1264 11241 1298
rect 11183 1230 11241 1264
rect 11183 1196 11195 1230
rect 11229 1196 11241 1230
rect 11183 1162 11241 1196
rect 11183 1128 11195 1162
rect 11229 1128 11241 1162
rect 11183 1004 11241 1128
rect 11271 1366 11329 1404
rect 11271 1332 11283 1366
rect 11317 1332 11329 1366
rect 11271 1298 11329 1332
rect 11271 1264 11283 1298
rect 11317 1264 11329 1298
rect 11271 1230 11329 1264
rect 11271 1196 11283 1230
rect 11317 1196 11329 1230
rect 11271 1162 11329 1196
rect 11271 1128 11283 1162
rect 11317 1128 11329 1162
rect 11271 1093 11329 1128
rect 11271 1059 11283 1093
rect 11317 1059 11329 1093
rect 11271 1004 11329 1059
rect 11359 1366 11413 1404
rect 11359 1332 11371 1366
rect 11405 1332 11413 1366
rect 11359 1298 11413 1332
rect 11359 1264 11371 1298
rect 11405 1264 11413 1298
rect 11359 1230 11413 1264
rect 11359 1196 11371 1230
rect 11405 1196 11413 1230
rect 11359 1162 11413 1196
rect 11359 1128 11371 1162
rect 11405 1128 11413 1162
rect 11359 1004 11413 1128
rect 11675 1366 11731 1404
rect 11675 1332 11685 1366
rect 11719 1332 11731 1366
rect 11675 1298 11731 1332
rect 11675 1264 11685 1298
rect 11719 1264 11731 1298
rect 11675 1230 11731 1264
rect 11675 1196 11685 1230
rect 11719 1196 11731 1230
rect 11675 1162 11731 1196
rect 11675 1128 11685 1162
rect 11719 1128 11731 1162
rect 11675 1093 11731 1128
rect 11675 1059 11685 1093
rect 11719 1059 11731 1093
rect 11675 1004 11731 1059
rect 11761 1366 11819 1404
rect 11761 1332 11773 1366
rect 11807 1332 11819 1366
rect 11761 1298 11819 1332
rect 11761 1264 11773 1298
rect 11807 1264 11819 1298
rect 11761 1230 11819 1264
rect 11761 1196 11773 1230
rect 11807 1196 11819 1230
rect 11761 1162 11819 1196
rect 11761 1128 11773 1162
rect 11807 1128 11819 1162
rect 11761 1093 11819 1128
rect 11761 1059 11773 1093
rect 11807 1059 11819 1093
rect 11761 1004 11819 1059
rect 11849 1366 11907 1404
rect 11849 1332 11861 1366
rect 11895 1332 11907 1366
rect 11849 1298 11907 1332
rect 11849 1264 11861 1298
rect 11895 1264 11907 1298
rect 11849 1230 11907 1264
rect 11849 1196 11861 1230
rect 11895 1196 11907 1230
rect 11849 1162 11907 1196
rect 11849 1128 11861 1162
rect 11895 1128 11907 1162
rect 11849 1004 11907 1128
rect 11937 1366 11995 1404
rect 11937 1332 11949 1366
rect 11983 1332 11995 1366
rect 11937 1298 11995 1332
rect 11937 1264 11949 1298
rect 11983 1264 11995 1298
rect 11937 1230 11995 1264
rect 11937 1196 11949 1230
rect 11983 1196 11995 1230
rect 11937 1162 11995 1196
rect 11937 1128 11949 1162
rect 11983 1128 11995 1162
rect 11937 1093 11995 1128
rect 11937 1059 11949 1093
rect 11983 1059 11995 1093
rect 11937 1004 11995 1059
rect 12025 1366 12079 1404
rect 12025 1332 12037 1366
rect 12071 1332 12079 1366
rect 12025 1298 12079 1332
rect 12025 1264 12037 1298
rect 12071 1264 12079 1298
rect 12025 1230 12079 1264
rect 12025 1196 12037 1230
rect 12071 1196 12079 1230
rect 12025 1162 12079 1196
rect 12025 1128 12037 1162
rect 12071 1128 12079 1162
rect 12025 1004 12079 1128
rect 12341 1366 12397 1404
rect 12341 1332 12351 1366
rect 12385 1332 12397 1366
rect 12341 1298 12397 1332
rect 12341 1264 12351 1298
rect 12385 1264 12397 1298
rect 12341 1230 12397 1264
rect 12341 1196 12351 1230
rect 12385 1196 12397 1230
rect 12341 1162 12397 1196
rect 12341 1128 12351 1162
rect 12385 1128 12397 1162
rect 12341 1093 12397 1128
rect 12341 1059 12351 1093
rect 12385 1059 12397 1093
rect 12341 1004 12397 1059
rect 12427 1366 12485 1404
rect 12427 1332 12439 1366
rect 12473 1332 12485 1366
rect 12427 1298 12485 1332
rect 12427 1264 12439 1298
rect 12473 1264 12485 1298
rect 12427 1230 12485 1264
rect 12427 1196 12439 1230
rect 12473 1196 12485 1230
rect 12427 1162 12485 1196
rect 12427 1128 12439 1162
rect 12473 1128 12485 1162
rect 12427 1093 12485 1128
rect 12427 1059 12439 1093
rect 12473 1059 12485 1093
rect 12427 1004 12485 1059
rect 12515 1366 12573 1404
rect 12515 1332 12527 1366
rect 12561 1332 12573 1366
rect 12515 1298 12573 1332
rect 12515 1264 12527 1298
rect 12561 1264 12573 1298
rect 12515 1230 12573 1264
rect 12515 1196 12527 1230
rect 12561 1196 12573 1230
rect 12515 1162 12573 1196
rect 12515 1128 12527 1162
rect 12561 1128 12573 1162
rect 12515 1004 12573 1128
rect 12603 1366 12661 1404
rect 12603 1332 12615 1366
rect 12649 1332 12661 1366
rect 12603 1298 12661 1332
rect 12603 1264 12615 1298
rect 12649 1264 12661 1298
rect 12603 1230 12661 1264
rect 12603 1196 12615 1230
rect 12649 1196 12661 1230
rect 12603 1162 12661 1196
rect 12603 1128 12615 1162
rect 12649 1128 12661 1162
rect 12603 1093 12661 1128
rect 12603 1059 12615 1093
rect 12649 1059 12661 1093
rect 12603 1004 12661 1059
rect 12691 1366 12745 1404
rect 12691 1332 12703 1366
rect 12737 1332 12745 1366
rect 12691 1298 12745 1332
rect 12691 1264 12703 1298
rect 12737 1264 12745 1298
rect 12691 1230 12745 1264
rect 12691 1196 12703 1230
rect 12737 1196 12745 1230
rect 12691 1162 12745 1196
rect 12691 1128 12703 1162
rect 12737 1128 12745 1162
rect 12691 1004 12745 1128
rect 13007 1365 13063 1405
rect 13007 1331 13017 1365
rect 13051 1331 13063 1365
rect 13007 1297 13063 1331
rect 13007 1263 13017 1297
rect 13051 1263 13063 1297
rect 13007 1229 13063 1263
rect 13007 1195 13017 1229
rect 13051 1195 13063 1229
rect 13007 1161 13063 1195
rect 13007 1127 13017 1161
rect 13051 1127 13063 1161
rect 13007 1093 13063 1127
rect 13007 1059 13017 1093
rect 13051 1059 13063 1093
rect 13007 1005 13063 1059
rect 13093 1365 13151 1405
rect 13093 1331 13105 1365
rect 13139 1331 13151 1365
rect 13093 1297 13151 1331
rect 13093 1263 13105 1297
rect 13139 1263 13151 1297
rect 13093 1229 13151 1263
rect 13093 1195 13105 1229
rect 13139 1195 13151 1229
rect 13093 1161 13151 1195
rect 13093 1127 13105 1161
rect 13139 1127 13151 1161
rect 13093 1093 13151 1127
rect 13093 1059 13105 1093
rect 13139 1059 13151 1093
rect 13093 1005 13151 1059
rect 13181 1365 13239 1405
rect 13181 1331 13193 1365
rect 13227 1331 13239 1365
rect 13181 1297 13239 1331
rect 13181 1263 13193 1297
rect 13227 1263 13239 1297
rect 13181 1229 13239 1263
rect 13181 1195 13193 1229
rect 13227 1195 13239 1229
rect 13181 1161 13239 1195
rect 13181 1127 13193 1161
rect 13227 1127 13239 1161
rect 13181 1005 13239 1127
rect 13269 1365 13327 1405
rect 13269 1331 13281 1365
rect 13315 1331 13327 1365
rect 13269 1297 13327 1331
rect 13269 1263 13281 1297
rect 13315 1263 13327 1297
rect 13269 1229 13327 1263
rect 13269 1195 13281 1229
rect 13315 1195 13327 1229
rect 13269 1161 13327 1195
rect 13269 1127 13281 1161
rect 13315 1127 13327 1161
rect 13269 1005 13327 1127
rect 13357 1365 13411 1405
rect 13357 1331 13369 1365
rect 13403 1331 13411 1365
rect 13357 1297 13411 1331
rect 13357 1263 13369 1297
rect 13403 1263 13411 1297
rect 13357 1229 13411 1263
rect 13357 1195 13369 1229
rect 13403 1195 13411 1229
rect 13357 1161 13411 1195
rect 13357 1127 13369 1161
rect 13403 1127 13411 1161
rect 13357 1093 13411 1127
rect 13357 1059 13369 1093
rect 13403 1059 13411 1093
rect 13357 1005 13411 1059
rect 13673 1365 13727 1405
rect 13673 1331 13681 1365
rect 13715 1331 13727 1365
rect 13673 1297 13727 1331
rect 13673 1263 13681 1297
rect 13715 1263 13727 1297
rect 13673 1229 13727 1263
rect 13673 1195 13681 1229
rect 13715 1195 13727 1229
rect 13673 1161 13727 1195
rect 13673 1127 13681 1161
rect 13715 1127 13727 1161
rect 13673 1005 13727 1127
rect 13757 1297 13815 1405
rect 13757 1263 13769 1297
rect 13803 1263 13815 1297
rect 13757 1229 13815 1263
rect 13757 1195 13769 1229
rect 13803 1195 13815 1229
rect 13757 1161 13815 1195
rect 13757 1127 13769 1161
rect 13803 1127 13815 1161
rect 13757 1093 13815 1127
rect 13757 1059 13769 1093
rect 13803 1059 13815 1093
rect 13757 1005 13815 1059
rect 13845 1365 13903 1405
rect 13845 1331 13857 1365
rect 13891 1331 13903 1365
rect 13845 1297 13903 1331
rect 13845 1263 13857 1297
rect 13891 1263 13903 1297
rect 13845 1229 13903 1263
rect 13845 1195 13857 1229
rect 13891 1195 13903 1229
rect 13845 1161 13903 1195
rect 13845 1127 13857 1161
rect 13891 1127 13903 1161
rect 13845 1005 13903 1127
rect 13933 1297 13991 1405
rect 13933 1263 13945 1297
rect 13979 1263 13991 1297
rect 13933 1229 13991 1263
rect 13933 1195 13945 1229
rect 13979 1195 13991 1229
rect 13933 1161 13991 1195
rect 13933 1127 13945 1161
rect 13979 1127 13991 1161
rect 13933 1005 13991 1127
rect 14021 1365 14077 1405
rect 14021 1331 14033 1365
rect 14067 1331 14077 1365
rect 14021 1297 14077 1331
rect 14021 1263 14033 1297
rect 14067 1263 14077 1297
rect 14021 1229 14077 1263
rect 14021 1195 14033 1229
rect 14067 1195 14077 1229
rect 14021 1161 14077 1195
rect 14021 1127 14033 1161
rect 14067 1127 14077 1161
rect 14021 1005 14077 1127
rect 14339 1365 14395 1405
rect 14339 1331 14349 1365
rect 14383 1331 14395 1365
rect 14339 1297 14395 1331
rect 14339 1263 14349 1297
rect 14383 1263 14395 1297
rect 14339 1229 14395 1263
rect 14339 1195 14349 1229
rect 14383 1195 14395 1229
rect 14339 1161 14395 1195
rect 14339 1127 14349 1161
rect 14383 1127 14395 1161
rect 14339 1005 14395 1127
rect 14425 1297 14483 1405
rect 14425 1263 14437 1297
rect 14471 1263 14483 1297
rect 14425 1229 14483 1263
rect 14425 1195 14437 1229
rect 14471 1195 14483 1229
rect 14425 1161 14483 1195
rect 14425 1127 14437 1161
rect 14471 1127 14483 1161
rect 14425 1093 14483 1127
rect 14425 1059 14437 1093
rect 14471 1059 14483 1093
rect 14425 1005 14483 1059
rect 14513 1365 14571 1405
rect 14513 1331 14525 1365
rect 14559 1331 14571 1365
rect 14513 1297 14571 1331
rect 14513 1263 14525 1297
rect 14559 1263 14571 1297
rect 14513 1229 14571 1263
rect 14513 1195 14525 1229
rect 14559 1195 14571 1229
rect 14513 1161 14571 1195
rect 14513 1127 14525 1161
rect 14559 1127 14571 1161
rect 14513 1005 14571 1127
rect 14601 1297 14659 1405
rect 14601 1263 14613 1297
rect 14647 1263 14659 1297
rect 14601 1229 14659 1263
rect 14601 1195 14613 1229
rect 14647 1195 14659 1229
rect 14601 1161 14659 1195
rect 14601 1127 14613 1161
rect 14647 1127 14659 1161
rect 14601 1093 14659 1127
rect 14601 1059 14613 1093
rect 14647 1059 14659 1093
rect 14601 1005 14659 1059
rect 14689 1365 14743 1405
rect 14689 1331 14701 1365
rect 14735 1331 14743 1365
rect 14689 1297 14743 1331
rect 14689 1263 14701 1297
rect 14735 1263 14743 1297
rect 14689 1229 14743 1263
rect 14689 1195 14701 1229
rect 14735 1195 14743 1229
rect 14689 1161 14743 1195
rect 14689 1127 14701 1161
rect 14735 1127 14743 1161
rect 14689 1005 14743 1127
<< ndiffc >>
rect 101 301 135 335
rect 198 301 232 335
rect 295 301 329 335
rect 392 301 426 335
rect 489 301 523 335
rect 101 229 135 263
rect 101 161 135 195
rect 198 176 232 210
rect 295 229 329 263
rect 295 161 329 195
rect 393 182 427 216
rect 101 91 135 125
rect 295 91 329 125
rect 392 91 426 125
rect 489 91 523 125
rect 603 301 637 335
rect 603 229 637 263
rect 603 161 637 195
rect 700 185 734 219
rect 797 229 831 263
rect 797 161 831 195
rect 603 91 637 125
rect 700 91 734 125
rect 797 91 831 125
rect 1084 299 1118 333
rect 1181 299 1215 333
rect 1278 299 1312 333
rect 1084 227 1118 261
rect 1084 159 1118 193
rect 1181 174 1215 208
rect 1278 227 1312 261
rect 1278 159 1312 193
rect 1375 183 1409 217
rect 1472 227 1506 261
rect 1472 159 1506 193
rect 1084 89 1118 123
rect 1278 89 1312 123
rect 1375 89 1409 123
rect 1472 89 1506 123
rect 1750 299 1784 333
rect 1847 299 1881 333
rect 1944 299 1978 333
rect 1750 227 1784 261
rect 1750 159 1784 193
rect 1847 174 1881 208
rect 1944 227 1978 261
rect 1944 159 1978 193
rect 2041 183 2075 217
rect 2138 227 2172 261
rect 2138 159 2172 193
rect 1750 89 1784 123
rect 1944 89 1978 123
rect 2041 89 2075 123
rect 2138 89 2172 123
rect 2416 299 2450 333
rect 2513 299 2547 333
rect 2610 299 2644 333
rect 2416 227 2450 261
rect 2416 159 2450 193
rect 2513 174 2547 208
rect 2610 227 2644 261
rect 2610 159 2644 193
rect 2707 183 2741 217
rect 2804 227 2838 261
rect 2804 159 2838 193
rect 2416 89 2450 123
rect 2610 89 2644 123
rect 2707 89 2741 123
rect 2804 89 2838 123
rect 3082 299 3116 333
rect 3179 299 3213 333
rect 3276 299 3310 333
rect 3082 227 3116 261
rect 3082 159 3116 193
rect 3179 174 3213 208
rect 3276 227 3310 261
rect 3276 159 3310 193
rect 3373 183 3407 217
rect 3470 227 3504 261
rect 3470 159 3504 193
rect 3082 89 3116 123
rect 3276 89 3310 123
rect 3373 89 3407 123
rect 3470 89 3504 123
rect 3748 299 3782 333
rect 3845 299 3879 333
rect 3942 299 3976 333
rect 3748 227 3782 261
rect 3748 159 3782 193
rect 3845 174 3879 208
rect 3942 227 3976 261
rect 3942 159 3976 193
rect 4039 183 4073 217
rect 4136 227 4170 261
rect 4136 159 4170 193
rect 3748 89 3782 123
rect 3942 89 3976 123
rect 4039 89 4073 123
rect 4136 89 4170 123
rect 4393 301 4427 335
rect 4490 301 4524 335
rect 4587 301 4621 335
rect 4684 301 4718 335
rect 4781 301 4815 335
rect 4393 229 4427 263
rect 4393 161 4427 195
rect 4490 176 4524 210
rect 4587 229 4621 263
rect 4587 161 4621 195
rect 4685 182 4719 216
rect 4393 91 4427 125
rect 4587 91 4621 125
rect 4684 91 4718 125
rect 4781 91 4815 125
rect 4895 301 4929 335
rect 4895 229 4929 263
rect 4895 161 4929 195
rect 4992 185 5026 219
rect 5089 229 5123 263
rect 5089 161 5123 195
rect 4895 91 4929 125
rect 4992 91 5026 125
rect 5089 91 5123 125
rect 5376 299 5410 333
rect 5473 299 5507 333
rect 5570 299 5604 333
rect 5376 227 5410 261
rect 5376 159 5410 193
rect 5473 174 5507 208
rect 5570 227 5604 261
rect 5570 159 5604 193
rect 5667 183 5701 217
rect 5764 227 5798 261
rect 5764 159 5798 193
rect 5376 89 5410 123
rect 5570 89 5604 123
rect 5667 89 5701 123
rect 5764 89 5798 123
rect 6042 299 6076 333
rect 6139 299 6173 333
rect 6236 299 6270 333
rect 6042 227 6076 261
rect 6042 159 6076 193
rect 6139 174 6173 208
rect 6236 227 6270 261
rect 6236 159 6270 193
rect 6333 183 6367 217
rect 6430 227 6464 261
rect 6430 159 6464 193
rect 6042 89 6076 123
rect 6236 89 6270 123
rect 6333 89 6367 123
rect 6430 89 6464 123
rect 6708 299 6742 333
rect 6805 299 6839 333
rect 6902 299 6936 333
rect 6708 227 6742 261
rect 6708 159 6742 193
rect 6805 174 6839 208
rect 6902 227 6936 261
rect 6902 159 6936 193
rect 6999 183 7033 217
rect 7096 227 7130 261
rect 7096 159 7130 193
rect 6708 89 6742 123
rect 6902 89 6936 123
rect 6999 89 7033 123
rect 7096 89 7130 123
rect 7374 299 7408 333
rect 7471 299 7505 333
rect 7568 299 7602 333
rect 7374 227 7408 261
rect 7374 159 7408 193
rect 7471 174 7505 208
rect 7568 227 7602 261
rect 7568 159 7602 193
rect 7665 183 7699 217
rect 7762 227 7796 261
rect 7762 159 7796 193
rect 7374 89 7408 123
rect 7568 89 7602 123
rect 7665 89 7699 123
rect 7762 89 7796 123
rect 8040 299 8074 333
rect 8137 299 8171 333
rect 8234 299 8268 333
rect 8040 227 8074 261
rect 8040 159 8074 193
rect 8137 174 8171 208
rect 8234 227 8268 261
rect 8234 159 8268 193
rect 8331 183 8365 217
rect 8428 227 8462 261
rect 8428 159 8462 193
rect 8040 89 8074 123
rect 8234 89 8268 123
rect 8331 89 8365 123
rect 8428 89 8462 123
rect 8685 301 8719 335
rect 8782 301 8816 335
rect 8879 301 8913 335
rect 8976 301 9010 335
rect 9073 301 9107 335
rect 8685 229 8719 263
rect 8685 161 8719 195
rect 8782 176 8816 210
rect 8879 229 8913 263
rect 8879 161 8913 195
rect 8977 182 9011 216
rect 8685 91 8719 125
rect 8879 91 8913 125
rect 8976 91 9010 125
rect 9073 91 9107 125
rect 9187 301 9221 335
rect 9187 229 9221 263
rect 9187 161 9221 195
rect 9284 185 9318 219
rect 9381 229 9415 263
rect 9381 161 9415 195
rect 9187 91 9221 125
rect 9284 91 9318 125
rect 9381 91 9415 125
rect 9668 299 9702 333
rect 9765 299 9799 333
rect 9862 299 9896 333
rect 9668 227 9702 261
rect 9668 159 9702 193
rect 9765 174 9799 208
rect 9862 227 9896 261
rect 9862 159 9896 193
rect 9959 183 9993 217
rect 10056 227 10090 261
rect 10056 159 10090 193
rect 9668 89 9702 123
rect 9862 89 9896 123
rect 9959 89 9993 123
rect 10056 89 10090 123
rect 10334 299 10368 333
rect 10431 299 10465 333
rect 10528 299 10562 333
rect 10334 227 10368 261
rect 10334 159 10368 193
rect 10431 174 10465 208
rect 10528 227 10562 261
rect 10528 159 10562 193
rect 10625 183 10659 217
rect 10722 227 10756 261
rect 10722 159 10756 193
rect 10334 89 10368 123
rect 10528 89 10562 123
rect 10625 89 10659 123
rect 10722 89 10756 123
rect 11000 299 11034 333
rect 11097 299 11131 333
rect 11194 299 11228 333
rect 11000 227 11034 261
rect 11000 159 11034 193
rect 11097 174 11131 208
rect 11194 227 11228 261
rect 11194 159 11228 193
rect 11291 183 11325 217
rect 11388 227 11422 261
rect 11388 159 11422 193
rect 11000 89 11034 123
rect 11194 89 11228 123
rect 11291 89 11325 123
rect 11388 89 11422 123
rect 11666 299 11700 333
rect 11763 299 11797 333
rect 11860 299 11894 333
rect 11666 227 11700 261
rect 11666 159 11700 193
rect 11763 174 11797 208
rect 11860 227 11894 261
rect 11860 159 11894 193
rect 11957 183 11991 217
rect 12054 227 12088 261
rect 12054 159 12088 193
rect 11666 89 11700 123
rect 11860 89 11894 123
rect 11957 89 11991 123
rect 12054 89 12088 123
rect 12332 299 12366 333
rect 12429 299 12463 333
rect 12526 299 12560 333
rect 12332 227 12366 261
rect 12332 159 12366 193
rect 12429 174 12463 208
rect 12526 227 12560 261
rect 12526 159 12560 193
rect 12623 183 12657 217
rect 12720 227 12754 261
rect 12720 159 12754 193
rect 12332 89 12366 123
rect 12526 89 12560 123
rect 12623 89 12657 123
rect 12720 89 12754 123
rect 12998 299 13032 333
rect 13095 299 13129 333
rect 13192 299 13226 333
rect 13386 299 13420 333
rect 12998 227 13032 261
rect 12998 159 13032 193
rect 13095 174 13129 208
rect 13192 227 13226 261
rect 13192 159 13226 193
rect 13288 183 13322 217
rect 13386 227 13420 261
rect 13386 159 13420 193
rect 12998 89 13032 123
rect 13192 89 13226 123
rect 13288 89 13322 123
rect 13386 89 13420 123
rect 13664 299 13698 333
rect 13761 299 13795 333
rect 13858 299 13892 333
rect 14052 299 14086 333
rect 13664 227 13698 261
rect 13664 159 13698 193
rect 13761 174 13795 208
rect 13858 227 13892 261
rect 13858 159 13892 193
rect 13955 183 13989 217
rect 14052 227 14086 261
rect 14052 159 14086 193
rect 13664 89 13698 123
rect 13858 89 13892 123
rect 13955 89 13989 123
rect 14052 89 14086 123
rect 14330 299 14364 333
rect 14427 299 14461 333
rect 14524 299 14558 333
rect 14330 227 14364 261
rect 14330 159 14364 193
rect 14427 174 14461 208
rect 14524 227 14558 261
rect 14524 159 14558 193
rect 14621 183 14655 217
rect 14718 227 14752 261
rect 14718 159 14752 193
rect 14330 89 14364 123
rect 14524 89 14558 123
rect 14621 89 14655 123
rect 14718 89 14752 123
<< pdiffc >>
rect 201 1332 235 1366
rect 201 1264 235 1298
rect 201 1196 235 1230
rect 201 1128 235 1162
rect 201 1059 235 1093
rect 289 1332 323 1366
rect 289 1264 323 1298
rect 289 1196 323 1230
rect 289 1128 323 1162
rect 289 1059 323 1093
rect 377 1332 411 1366
rect 377 1264 411 1298
rect 377 1196 411 1230
rect 377 1128 411 1162
rect 465 1332 499 1366
rect 465 1264 499 1298
rect 465 1196 499 1230
rect 465 1128 499 1162
rect 465 1059 499 1093
rect 553 1332 587 1366
rect 553 1264 587 1298
rect 553 1196 587 1230
rect 553 1128 587 1162
rect 641 1332 675 1366
rect 641 1264 675 1298
rect 641 1196 675 1230
rect 641 1128 675 1162
rect 641 1059 675 1093
rect 729 1332 763 1366
rect 729 1264 763 1298
rect 729 1196 763 1230
rect 729 1128 763 1162
rect 1103 1332 1137 1366
rect 1103 1264 1137 1298
rect 1103 1196 1137 1230
rect 1103 1128 1137 1162
rect 1103 1059 1137 1093
rect 1191 1332 1225 1366
rect 1191 1264 1225 1298
rect 1191 1196 1225 1230
rect 1191 1128 1225 1162
rect 1191 1059 1225 1093
rect 1279 1332 1313 1366
rect 1279 1264 1313 1298
rect 1279 1196 1313 1230
rect 1279 1128 1313 1162
rect 1367 1332 1401 1366
rect 1367 1264 1401 1298
rect 1367 1196 1401 1230
rect 1367 1128 1401 1162
rect 1367 1059 1401 1093
rect 1455 1332 1489 1366
rect 1455 1264 1489 1298
rect 1455 1196 1489 1230
rect 1455 1128 1489 1162
rect 1769 1332 1803 1366
rect 1769 1264 1803 1298
rect 1769 1196 1803 1230
rect 1769 1128 1803 1162
rect 1769 1059 1803 1093
rect 1857 1332 1891 1366
rect 1857 1264 1891 1298
rect 1857 1196 1891 1230
rect 1857 1128 1891 1162
rect 1857 1059 1891 1093
rect 1945 1332 1979 1366
rect 1945 1264 1979 1298
rect 1945 1196 1979 1230
rect 1945 1128 1979 1162
rect 2033 1332 2067 1366
rect 2033 1264 2067 1298
rect 2033 1196 2067 1230
rect 2033 1128 2067 1162
rect 2033 1059 2067 1093
rect 2121 1332 2155 1366
rect 2121 1264 2155 1298
rect 2121 1196 2155 1230
rect 2121 1128 2155 1162
rect 2435 1332 2469 1366
rect 2435 1264 2469 1298
rect 2435 1196 2469 1230
rect 2435 1128 2469 1162
rect 2435 1059 2469 1093
rect 2523 1332 2557 1366
rect 2523 1264 2557 1298
rect 2523 1196 2557 1230
rect 2523 1128 2557 1162
rect 2523 1059 2557 1093
rect 2611 1332 2645 1366
rect 2611 1264 2645 1298
rect 2611 1196 2645 1230
rect 2611 1128 2645 1162
rect 2699 1332 2733 1366
rect 2699 1264 2733 1298
rect 2699 1196 2733 1230
rect 2699 1128 2733 1162
rect 2699 1059 2733 1093
rect 2787 1332 2821 1366
rect 2787 1264 2821 1298
rect 2787 1196 2821 1230
rect 2787 1128 2821 1162
rect 3101 1332 3135 1366
rect 3101 1264 3135 1298
rect 3101 1196 3135 1230
rect 3101 1128 3135 1162
rect 3101 1059 3135 1093
rect 3189 1332 3223 1366
rect 3189 1264 3223 1298
rect 3189 1196 3223 1230
rect 3189 1128 3223 1162
rect 3189 1059 3223 1093
rect 3277 1332 3311 1366
rect 3277 1264 3311 1298
rect 3277 1196 3311 1230
rect 3277 1128 3311 1162
rect 3365 1332 3399 1366
rect 3365 1264 3399 1298
rect 3365 1196 3399 1230
rect 3365 1128 3399 1162
rect 3365 1059 3399 1093
rect 3453 1332 3487 1366
rect 3453 1264 3487 1298
rect 3453 1196 3487 1230
rect 3453 1128 3487 1162
rect 3767 1332 3801 1366
rect 3767 1264 3801 1298
rect 3767 1196 3801 1230
rect 3767 1128 3801 1162
rect 3767 1059 3801 1093
rect 3855 1332 3889 1366
rect 3855 1264 3889 1298
rect 3855 1196 3889 1230
rect 3855 1128 3889 1162
rect 3855 1059 3889 1093
rect 3943 1332 3977 1366
rect 3943 1264 3977 1298
rect 3943 1196 3977 1230
rect 3943 1128 3977 1162
rect 4031 1332 4065 1366
rect 4031 1264 4065 1298
rect 4031 1196 4065 1230
rect 4031 1128 4065 1162
rect 4031 1059 4065 1093
rect 4119 1332 4153 1366
rect 4119 1264 4153 1298
rect 4119 1196 4153 1230
rect 4119 1128 4153 1162
rect 4493 1332 4527 1366
rect 4493 1264 4527 1298
rect 4493 1196 4527 1230
rect 4493 1128 4527 1162
rect 4493 1059 4527 1093
rect 4581 1332 4615 1366
rect 4581 1264 4615 1298
rect 4581 1196 4615 1230
rect 4581 1128 4615 1162
rect 4581 1059 4615 1093
rect 4669 1332 4703 1366
rect 4669 1264 4703 1298
rect 4669 1196 4703 1230
rect 4669 1128 4703 1162
rect 4757 1332 4791 1366
rect 4757 1264 4791 1298
rect 4757 1196 4791 1230
rect 4757 1128 4791 1162
rect 4757 1059 4791 1093
rect 4845 1332 4879 1366
rect 4845 1264 4879 1298
rect 4845 1196 4879 1230
rect 4845 1128 4879 1162
rect 4933 1332 4967 1366
rect 4933 1264 4967 1298
rect 4933 1196 4967 1230
rect 4933 1128 4967 1162
rect 4933 1059 4967 1093
rect 5021 1332 5055 1366
rect 5021 1264 5055 1298
rect 5021 1196 5055 1230
rect 5021 1128 5055 1162
rect 5395 1332 5429 1366
rect 5395 1264 5429 1298
rect 5395 1196 5429 1230
rect 5395 1128 5429 1162
rect 5395 1059 5429 1093
rect 5483 1332 5517 1366
rect 5483 1264 5517 1298
rect 5483 1196 5517 1230
rect 5483 1128 5517 1162
rect 5483 1059 5517 1093
rect 5571 1332 5605 1366
rect 5571 1264 5605 1298
rect 5571 1196 5605 1230
rect 5571 1128 5605 1162
rect 5659 1332 5693 1366
rect 5659 1264 5693 1298
rect 5659 1196 5693 1230
rect 5659 1128 5693 1162
rect 5659 1059 5693 1093
rect 5747 1332 5781 1366
rect 5747 1264 5781 1298
rect 5747 1196 5781 1230
rect 5747 1128 5781 1162
rect 6061 1332 6095 1366
rect 6061 1264 6095 1298
rect 6061 1196 6095 1230
rect 6061 1128 6095 1162
rect 6061 1059 6095 1093
rect 6149 1332 6183 1366
rect 6149 1264 6183 1298
rect 6149 1196 6183 1230
rect 6149 1128 6183 1162
rect 6149 1059 6183 1093
rect 6237 1332 6271 1366
rect 6237 1264 6271 1298
rect 6237 1196 6271 1230
rect 6237 1128 6271 1162
rect 6325 1332 6359 1366
rect 6325 1264 6359 1298
rect 6325 1196 6359 1230
rect 6325 1128 6359 1162
rect 6325 1059 6359 1093
rect 6413 1332 6447 1366
rect 6413 1264 6447 1298
rect 6413 1196 6447 1230
rect 6413 1128 6447 1162
rect 6727 1332 6761 1366
rect 6727 1264 6761 1298
rect 6727 1196 6761 1230
rect 6727 1128 6761 1162
rect 6727 1059 6761 1093
rect 6815 1332 6849 1366
rect 6815 1264 6849 1298
rect 6815 1196 6849 1230
rect 6815 1128 6849 1162
rect 6815 1059 6849 1093
rect 6903 1332 6937 1366
rect 6903 1264 6937 1298
rect 6903 1196 6937 1230
rect 6903 1128 6937 1162
rect 6991 1332 7025 1366
rect 6991 1264 7025 1298
rect 6991 1196 7025 1230
rect 6991 1128 7025 1162
rect 6991 1059 7025 1093
rect 7079 1332 7113 1366
rect 7079 1264 7113 1298
rect 7079 1196 7113 1230
rect 7079 1128 7113 1162
rect 7393 1332 7427 1366
rect 7393 1264 7427 1298
rect 7393 1196 7427 1230
rect 7393 1128 7427 1162
rect 7393 1059 7427 1093
rect 7481 1332 7515 1366
rect 7481 1264 7515 1298
rect 7481 1196 7515 1230
rect 7481 1128 7515 1162
rect 7481 1059 7515 1093
rect 7569 1332 7603 1366
rect 7569 1264 7603 1298
rect 7569 1196 7603 1230
rect 7569 1128 7603 1162
rect 7657 1332 7691 1366
rect 7657 1264 7691 1298
rect 7657 1196 7691 1230
rect 7657 1128 7691 1162
rect 7657 1059 7691 1093
rect 7745 1332 7779 1366
rect 7745 1264 7779 1298
rect 7745 1196 7779 1230
rect 7745 1128 7779 1162
rect 8059 1332 8093 1366
rect 8059 1264 8093 1298
rect 8059 1196 8093 1230
rect 8059 1128 8093 1162
rect 8059 1059 8093 1093
rect 8147 1332 8181 1366
rect 8147 1264 8181 1298
rect 8147 1196 8181 1230
rect 8147 1128 8181 1162
rect 8147 1059 8181 1093
rect 8235 1332 8269 1366
rect 8235 1264 8269 1298
rect 8235 1196 8269 1230
rect 8235 1128 8269 1162
rect 8323 1332 8357 1366
rect 8323 1264 8357 1298
rect 8323 1196 8357 1230
rect 8323 1128 8357 1162
rect 8323 1059 8357 1093
rect 8411 1332 8445 1366
rect 8411 1264 8445 1298
rect 8411 1196 8445 1230
rect 8411 1128 8445 1162
rect 8785 1332 8819 1366
rect 8785 1264 8819 1298
rect 8785 1196 8819 1230
rect 8785 1128 8819 1162
rect 8785 1059 8819 1093
rect 8873 1332 8907 1366
rect 8873 1264 8907 1298
rect 8873 1196 8907 1230
rect 8873 1128 8907 1162
rect 8873 1059 8907 1093
rect 8961 1332 8995 1366
rect 8961 1264 8995 1298
rect 8961 1196 8995 1230
rect 8961 1128 8995 1162
rect 9049 1332 9083 1366
rect 9049 1264 9083 1298
rect 9049 1196 9083 1230
rect 9049 1128 9083 1162
rect 9049 1059 9083 1093
rect 9137 1332 9171 1366
rect 9137 1264 9171 1298
rect 9137 1196 9171 1230
rect 9137 1128 9171 1162
rect 9225 1332 9259 1366
rect 9225 1264 9259 1298
rect 9225 1196 9259 1230
rect 9225 1128 9259 1162
rect 9225 1059 9259 1093
rect 9313 1332 9347 1366
rect 9313 1264 9347 1298
rect 9313 1196 9347 1230
rect 9313 1128 9347 1162
rect 9687 1332 9721 1366
rect 9687 1264 9721 1298
rect 9687 1196 9721 1230
rect 9687 1128 9721 1162
rect 9687 1059 9721 1093
rect 9775 1332 9809 1366
rect 9775 1264 9809 1298
rect 9775 1196 9809 1230
rect 9775 1128 9809 1162
rect 9775 1059 9809 1093
rect 9863 1332 9897 1366
rect 9863 1264 9897 1298
rect 9863 1196 9897 1230
rect 9863 1128 9897 1162
rect 9951 1332 9985 1366
rect 9951 1264 9985 1298
rect 9951 1196 9985 1230
rect 9951 1128 9985 1162
rect 9951 1059 9985 1093
rect 10039 1332 10073 1366
rect 10039 1264 10073 1298
rect 10039 1196 10073 1230
rect 10039 1128 10073 1162
rect 10353 1332 10387 1366
rect 10353 1264 10387 1298
rect 10353 1196 10387 1230
rect 10353 1128 10387 1162
rect 10353 1059 10387 1093
rect 10441 1332 10475 1366
rect 10441 1264 10475 1298
rect 10441 1196 10475 1230
rect 10441 1128 10475 1162
rect 10441 1059 10475 1093
rect 10529 1332 10563 1366
rect 10529 1264 10563 1298
rect 10529 1196 10563 1230
rect 10529 1128 10563 1162
rect 10617 1332 10651 1366
rect 10617 1264 10651 1298
rect 10617 1196 10651 1230
rect 10617 1128 10651 1162
rect 10617 1059 10651 1093
rect 10705 1332 10739 1366
rect 10705 1264 10739 1298
rect 10705 1196 10739 1230
rect 10705 1128 10739 1162
rect 11019 1332 11053 1366
rect 11019 1264 11053 1298
rect 11019 1196 11053 1230
rect 11019 1128 11053 1162
rect 11019 1059 11053 1093
rect 11107 1332 11141 1366
rect 11107 1264 11141 1298
rect 11107 1196 11141 1230
rect 11107 1128 11141 1162
rect 11107 1059 11141 1093
rect 11195 1332 11229 1366
rect 11195 1264 11229 1298
rect 11195 1196 11229 1230
rect 11195 1128 11229 1162
rect 11283 1332 11317 1366
rect 11283 1264 11317 1298
rect 11283 1196 11317 1230
rect 11283 1128 11317 1162
rect 11283 1059 11317 1093
rect 11371 1332 11405 1366
rect 11371 1264 11405 1298
rect 11371 1196 11405 1230
rect 11371 1128 11405 1162
rect 11685 1332 11719 1366
rect 11685 1264 11719 1298
rect 11685 1196 11719 1230
rect 11685 1128 11719 1162
rect 11685 1059 11719 1093
rect 11773 1332 11807 1366
rect 11773 1264 11807 1298
rect 11773 1196 11807 1230
rect 11773 1128 11807 1162
rect 11773 1059 11807 1093
rect 11861 1332 11895 1366
rect 11861 1264 11895 1298
rect 11861 1196 11895 1230
rect 11861 1128 11895 1162
rect 11949 1332 11983 1366
rect 11949 1264 11983 1298
rect 11949 1196 11983 1230
rect 11949 1128 11983 1162
rect 11949 1059 11983 1093
rect 12037 1332 12071 1366
rect 12037 1264 12071 1298
rect 12037 1196 12071 1230
rect 12037 1128 12071 1162
rect 12351 1332 12385 1366
rect 12351 1264 12385 1298
rect 12351 1196 12385 1230
rect 12351 1128 12385 1162
rect 12351 1059 12385 1093
rect 12439 1332 12473 1366
rect 12439 1264 12473 1298
rect 12439 1196 12473 1230
rect 12439 1128 12473 1162
rect 12439 1059 12473 1093
rect 12527 1332 12561 1366
rect 12527 1264 12561 1298
rect 12527 1196 12561 1230
rect 12527 1128 12561 1162
rect 12615 1332 12649 1366
rect 12615 1264 12649 1298
rect 12615 1196 12649 1230
rect 12615 1128 12649 1162
rect 12615 1059 12649 1093
rect 12703 1332 12737 1366
rect 12703 1264 12737 1298
rect 12703 1196 12737 1230
rect 12703 1128 12737 1162
rect 13017 1331 13051 1365
rect 13017 1263 13051 1297
rect 13017 1195 13051 1229
rect 13017 1127 13051 1161
rect 13017 1059 13051 1093
rect 13105 1331 13139 1365
rect 13105 1263 13139 1297
rect 13105 1195 13139 1229
rect 13105 1127 13139 1161
rect 13105 1059 13139 1093
rect 13193 1331 13227 1365
rect 13193 1263 13227 1297
rect 13193 1195 13227 1229
rect 13193 1127 13227 1161
rect 13281 1331 13315 1365
rect 13281 1263 13315 1297
rect 13281 1195 13315 1229
rect 13281 1127 13315 1161
rect 13369 1331 13403 1365
rect 13369 1263 13403 1297
rect 13369 1195 13403 1229
rect 13369 1127 13403 1161
rect 13369 1059 13403 1093
rect 13681 1331 13715 1365
rect 13681 1263 13715 1297
rect 13681 1195 13715 1229
rect 13681 1127 13715 1161
rect 13769 1263 13803 1297
rect 13769 1195 13803 1229
rect 13769 1127 13803 1161
rect 13769 1059 13803 1093
rect 13857 1331 13891 1365
rect 13857 1263 13891 1297
rect 13857 1195 13891 1229
rect 13857 1127 13891 1161
rect 13945 1263 13979 1297
rect 13945 1195 13979 1229
rect 13945 1127 13979 1161
rect 14033 1331 14067 1365
rect 14033 1263 14067 1297
rect 14033 1195 14067 1229
rect 14033 1127 14067 1161
rect 14349 1331 14383 1365
rect 14349 1263 14383 1297
rect 14349 1195 14383 1229
rect 14349 1127 14383 1161
rect 14437 1263 14471 1297
rect 14437 1195 14471 1229
rect 14437 1127 14471 1161
rect 14437 1059 14471 1093
rect 14525 1331 14559 1365
rect 14525 1263 14559 1297
rect 14525 1195 14559 1229
rect 14525 1127 14559 1161
rect 14613 1263 14647 1297
rect 14613 1195 14647 1229
rect 14613 1127 14647 1161
rect 14613 1059 14647 1093
rect 14701 1331 14735 1365
rect 14701 1263 14735 1297
rect 14701 1195 14735 1229
rect 14701 1127 14735 1161
<< psubdiff >>
rect -34 482 14908 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 928 461 996 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 928 427 945 461
rect 979 427 996 461
rect 1594 461 1662 482
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 928 313 996 353
rect 1594 427 1611 461
rect 1645 427 1662 461
rect 2260 461 2328 482
rect 1594 387 1662 427
rect 1594 353 1611 387
rect 1645 353 1662 387
rect 928 279 945 313
rect 979 279 996 313
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect -34 17 34 57
rect 928 57 945 91
rect 979 57 996 91
rect 1594 313 1662 353
rect 2260 427 2277 461
rect 2311 427 2328 461
rect 2926 461 2994 482
rect 2260 387 2328 427
rect 2260 353 2277 387
rect 2311 353 2328 387
rect 1594 279 1611 313
rect 1645 279 1662 313
rect 1594 239 1662 279
rect 1594 205 1611 239
rect 1645 205 1662 239
rect 1594 165 1662 205
rect 1594 131 1611 165
rect 1645 131 1662 165
rect 1594 91 1662 131
rect 928 17 996 57
rect 1594 57 1611 91
rect 1645 57 1662 91
rect 2260 313 2328 353
rect 2926 427 2943 461
rect 2977 427 2994 461
rect 3592 461 3660 482
rect 2926 387 2994 427
rect 2926 353 2943 387
rect 2977 353 2994 387
rect 2260 279 2277 313
rect 2311 279 2328 313
rect 2260 239 2328 279
rect 2260 205 2277 239
rect 2311 205 2328 239
rect 2260 165 2328 205
rect 2260 131 2277 165
rect 2311 131 2328 165
rect 2260 91 2328 131
rect 1594 17 1662 57
rect 2260 57 2277 91
rect 2311 57 2328 91
rect 2926 313 2994 353
rect 3592 427 3609 461
rect 3643 427 3660 461
rect 4258 461 4326 482
rect 3592 387 3660 427
rect 3592 353 3609 387
rect 3643 353 3660 387
rect 2926 279 2943 313
rect 2977 279 2994 313
rect 2926 239 2994 279
rect 2926 205 2943 239
rect 2977 205 2994 239
rect 2926 165 2994 205
rect 2926 131 2943 165
rect 2977 131 2994 165
rect 2926 91 2994 131
rect 2260 17 2328 57
rect 2926 57 2943 91
rect 2977 57 2994 91
rect 3592 313 3660 353
rect 4258 427 4275 461
rect 4309 427 4326 461
rect 5220 461 5288 482
rect 4258 387 4326 427
rect 4258 353 4275 387
rect 4309 353 4326 387
rect 3592 279 3609 313
rect 3643 279 3660 313
rect 3592 239 3660 279
rect 3592 205 3609 239
rect 3643 205 3660 239
rect 3592 165 3660 205
rect 3592 131 3609 165
rect 3643 131 3660 165
rect 3592 91 3660 131
rect 2926 17 2994 57
rect 3592 57 3609 91
rect 3643 57 3660 91
rect 4258 313 4326 353
rect 5220 427 5237 461
rect 5271 427 5288 461
rect 5886 461 5954 482
rect 5220 387 5288 427
rect 5220 353 5237 387
rect 5271 353 5288 387
rect 4258 279 4275 313
rect 4309 279 4326 313
rect 4258 239 4326 279
rect 4258 205 4275 239
rect 4309 205 4326 239
rect 4258 165 4326 205
rect 4258 131 4275 165
rect 4309 131 4326 165
rect 4258 91 4326 131
rect 3592 17 3660 57
rect 4258 57 4275 91
rect 4309 57 4326 91
rect 5220 313 5288 353
rect 5886 427 5903 461
rect 5937 427 5954 461
rect 6552 461 6620 482
rect 5886 387 5954 427
rect 5886 353 5903 387
rect 5937 353 5954 387
rect 5220 279 5237 313
rect 5271 279 5288 313
rect 5220 239 5288 279
rect 5220 205 5237 239
rect 5271 205 5288 239
rect 5220 165 5288 205
rect 5220 131 5237 165
rect 5271 131 5288 165
rect 5220 91 5288 131
rect 4258 17 4326 57
rect 5220 57 5237 91
rect 5271 57 5288 91
rect 5886 313 5954 353
rect 6552 427 6569 461
rect 6603 427 6620 461
rect 7218 461 7286 482
rect 6552 387 6620 427
rect 6552 353 6569 387
rect 6603 353 6620 387
rect 5886 279 5903 313
rect 5937 279 5954 313
rect 5886 239 5954 279
rect 5886 205 5903 239
rect 5937 205 5954 239
rect 5886 165 5954 205
rect 5886 131 5903 165
rect 5937 131 5954 165
rect 5886 91 5954 131
rect 5220 17 5288 57
rect 5886 57 5903 91
rect 5937 57 5954 91
rect 6552 313 6620 353
rect 7218 427 7235 461
rect 7269 427 7286 461
rect 7884 461 7952 482
rect 7218 387 7286 427
rect 7218 353 7235 387
rect 7269 353 7286 387
rect 6552 279 6569 313
rect 6603 279 6620 313
rect 6552 239 6620 279
rect 6552 205 6569 239
rect 6603 205 6620 239
rect 6552 165 6620 205
rect 6552 131 6569 165
rect 6603 131 6620 165
rect 6552 91 6620 131
rect 5886 17 5954 57
rect 6552 57 6569 91
rect 6603 57 6620 91
rect 7218 313 7286 353
rect 7884 427 7901 461
rect 7935 427 7952 461
rect 8550 461 8618 482
rect 7884 387 7952 427
rect 7884 353 7901 387
rect 7935 353 7952 387
rect 7218 279 7235 313
rect 7269 279 7286 313
rect 7218 239 7286 279
rect 7218 205 7235 239
rect 7269 205 7286 239
rect 7218 165 7286 205
rect 7218 131 7235 165
rect 7269 131 7286 165
rect 7218 91 7286 131
rect 6552 17 6620 57
rect 7218 57 7235 91
rect 7269 57 7286 91
rect 7884 313 7952 353
rect 8550 427 8567 461
rect 8601 427 8618 461
rect 9512 461 9580 482
rect 8550 387 8618 427
rect 8550 353 8567 387
rect 8601 353 8618 387
rect 7884 279 7901 313
rect 7935 279 7952 313
rect 7884 239 7952 279
rect 7884 205 7901 239
rect 7935 205 7952 239
rect 7884 165 7952 205
rect 7884 131 7901 165
rect 7935 131 7952 165
rect 7884 91 7952 131
rect 7218 17 7286 57
rect 7884 57 7901 91
rect 7935 57 7952 91
rect 8550 313 8618 353
rect 9512 427 9529 461
rect 9563 427 9580 461
rect 10178 461 10246 482
rect 9512 387 9580 427
rect 9512 353 9529 387
rect 9563 353 9580 387
rect 8550 279 8567 313
rect 8601 279 8618 313
rect 8550 239 8618 279
rect 8550 205 8567 239
rect 8601 205 8618 239
rect 8550 165 8618 205
rect 8550 131 8567 165
rect 8601 131 8618 165
rect 8550 91 8618 131
rect 7884 17 7952 57
rect 8550 57 8567 91
rect 8601 57 8618 91
rect 9512 313 9580 353
rect 10178 427 10195 461
rect 10229 427 10246 461
rect 10844 461 10912 482
rect 10178 387 10246 427
rect 10178 353 10195 387
rect 10229 353 10246 387
rect 9512 279 9529 313
rect 9563 279 9580 313
rect 9512 239 9580 279
rect 9512 205 9529 239
rect 9563 205 9580 239
rect 9512 165 9580 205
rect 9512 131 9529 165
rect 9563 131 9580 165
rect 9512 91 9580 131
rect 8550 17 8618 57
rect 9512 57 9529 91
rect 9563 57 9580 91
rect 10178 313 10246 353
rect 10844 427 10861 461
rect 10895 427 10912 461
rect 11510 461 11578 482
rect 10844 387 10912 427
rect 10844 353 10861 387
rect 10895 353 10912 387
rect 10178 279 10195 313
rect 10229 279 10246 313
rect 10178 239 10246 279
rect 10178 205 10195 239
rect 10229 205 10246 239
rect 10178 165 10246 205
rect 10178 131 10195 165
rect 10229 131 10246 165
rect 10178 91 10246 131
rect 9512 17 9580 57
rect 10178 57 10195 91
rect 10229 57 10246 91
rect 10844 313 10912 353
rect 11510 427 11527 461
rect 11561 427 11578 461
rect 12176 461 12244 482
rect 11510 387 11578 427
rect 11510 353 11527 387
rect 11561 353 11578 387
rect 10844 279 10861 313
rect 10895 279 10912 313
rect 10844 239 10912 279
rect 10844 205 10861 239
rect 10895 205 10912 239
rect 10844 165 10912 205
rect 10844 131 10861 165
rect 10895 131 10912 165
rect 10844 91 10912 131
rect 10178 17 10246 57
rect 10844 57 10861 91
rect 10895 57 10912 91
rect 11510 313 11578 353
rect 12176 427 12193 461
rect 12227 427 12244 461
rect 12842 461 12910 482
rect 12176 387 12244 427
rect 12176 353 12193 387
rect 12227 353 12244 387
rect 11510 279 11527 313
rect 11561 279 11578 313
rect 11510 239 11578 279
rect 11510 205 11527 239
rect 11561 205 11578 239
rect 11510 165 11578 205
rect 11510 131 11527 165
rect 11561 131 11578 165
rect 11510 91 11578 131
rect 10844 17 10912 57
rect 11510 57 11527 91
rect 11561 57 11578 91
rect 12176 313 12244 353
rect 12842 427 12859 461
rect 12893 427 12910 461
rect 13508 461 13576 482
rect 12842 387 12910 427
rect 12842 353 12859 387
rect 12893 353 12910 387
rect 13508 427 13525 461
rect 13559 427 13576 461
rect 14174 461 14242 482
rect 13508 387 13576 427
rect 12176 279 12193 313
rect 12227 279 12244 313
rect 12176 239 12244 279
rect 12176 205 12193 239
rect 12227 205 12244 239
rect 12176 165 12244 205
rect 12176 131 12193 165
rect 12227 131 12244 165
rect 12176 91 12244 131
rect 11510 17 11578 57
rect 12176 57 12193 91
rect 12227 57 12244 91
rect 12842 313 12910 353
rect 13508 353 13525 387
rect 13559 353 13576 387
rect 12842 279 12859 313
rect 12893 279 12910 313
rect 12842 239 12910 279
rect 12842 205 12859 239
rect 12893 205 12910 239
rect 12842 165 12910 205
rect 12842 131 12859 165
rect 12893 131 12910 165
rect 12842 91 12910 131
rect 12176 17 12244 57
rect 12842 57 12859 91
rect 12893 57 12910 91
rect 13508 313 13576 353
rect 14174 427 14191 461
rect 14225 427 14242 461
rect 14840 461 14908 482
rect 14174 387 14242 427
rect 14174 353 14191 387
rect 14225 353 14242 387
rect 14840 427 14857 461
rect 14891 427 14908 461
rect 14840 387 14908 427
rect 13508 279 13525 313
rect 13559 279 13576 313
rect 13508 239 13576 279
rect 13508 205 13525 239
rect 13559 205 13576 239
rect 13508 165 13576 205
rect 13508 131 13525 165
rect 13559 131 13576 165
rect 13508 91 13576 131
rect 12842 17 12910 57
rect 13508 57 13525 91
rect 13559 57 13576 91
rect 14174 313 14242 353
rect 14840 353 14857 387
rect 14891 353 14908 387
rect 14174 279 14191 313
rect 14225 279 14242 313
rect 14174 239 14242 279
rect 14174 205 14191 239
rect 14225 205 14242 239
rect 14174 165 14242 205
rect 14174 131 14191 165
rect 14225 131 14242 165
rect 14174 91 14242 131
rect 13508 17 13576 57
rect 14174 57 14191 91
rect 14225 57 14242 91
rect 14840 313 14908 353
rect 14840 279 14857 313
rect 14891 279 14908 313
rect 14840 239 14908 279
rect 14840 205 14857 239
rect 14891 205 14908 239
rect 14840 165 14908 205
rect 14840 131 14857 165
rect 14891 131 14908 165
rect 14840 91 14908 131
rect 14174 17 14242 57
rect 14840 57 14857 91
rect 14891 57 14908 91
rect 14840 17 14908 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5163 17
rect 5197 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5533 17
rect 5567 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5755 17
rect 5789 -17 5829 17
rect 5863 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6125 17
rect 6159 -17 6199 17
rect 6233 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6495 17
rect 6529 -17 6643 17
rect 6677 -17 6717 17
rect 6751 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7087 17
rect 7121 -17 7161 17
rect 7195 -17 7309 17
rect 7343 -17 7383 17
rect 7417 -17 7457 17
rect 7491 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7679 17
rect 7713 -17 7753 17
rect 7787 -17 7827 17
rect 7861 -17 7975 17
rect 8009 -17 8049 17
rect 8083 -17 8123 17
rect 8157 -17 8197 17
rect 8231 -17 8271 17
rect 8305 -17 8345 17
rect 8379 -17 8419 17
rect 8453 -17 8493 17
rect 8527 -17 8641 17
rect 8675 -17 8715 17
rect 8749 -17 8789 17
rect 8823 -17 8863 17
rect 8897 -17 8937 17
rect 8971 -17 9011 17
rect 9045 -17 9085 17
rect 9119 -17 9159 17
rect 9193 -17 9233 17
rect 9267 -17 9307 17
rect 9341 -17 9381 17
rect 9415 -17 9455 17
rect 9489 -17 9603 17
rect 9637 -17 9677 17
rect 9711 -17 9751 17
rect 9785 -17 9825 17
rect 9859 -17 9899 17
rect 9933 -17 9973 17
rect 10007 -17 10047 17
rect 10081 -17 10121 17
rect 10155 -17 10269 17
rect 10303 -17 10343 17
rect 10377 -17 10417 17
rect 10451 -17 10491 17
rect 10525 -17 10565 17
rect 10599 -17 10639 17
rect 10673 -17 10713 17
rect 10747 -17 10787 17
rect 10821 -17 10935 17
rect 10969 -17 11009 17
rect 11043 -17 11083 17
rect 11117 -17 11157 17
rect 11191 -17 11231 17
rect 11265 -17 11305 17
rect 11339 -17 11379 17
rect 11413 -17 11453 17
rect 11487 -17 11601 17
rect 11635 -17 11675 17
rect 11709 -17 11749 17
rect 11783 -17 11823 17
rect 11857 -17 11897 17
rect 11931 -17 11971 17
rect 12005 -17 12045 17
rect 12079 -17 12119 17
rect 12153 -17 12267 17
rect 12301 -17 12341 17
rect 12375 -17 12415 17
rect 12449 -17 12489 17
rect 12523 -17 12563 17
rect 12597 -17 12637 17
rect 12671 -17 12711 17
rect 12745 -17 12785 17
rect 12819 -17 12933 17
rect 12967 -17 13007 17
rect 13041 -17 13081 17
rect 13115 -17 13155 17
rect 13189 -17 13229 17
rect 13263 -17 13303 17
rect 13337 -17 13377 17
rect 13411 -17 13451 17
rect 13485 -17 13599 17
rect 13633 -17 13673 17
rect 13707 -17 13747 17
rect 13781 -17 13821 17
rect 13855 -17 13895 17
rect 13929 -17 13969 17
rect 14003 -17 14043 17
rect 14077 -17 14117 17
rect 14151 -17 14265 17
rect 14299 -17 14339 17
rect 14373 -17 14413 17
rect 14447 -17 14487 17
rect 14521 -17 14561 17
rect 14595 -17 14635 17
rect 14669 -17 14709 17
rect 14743 -17 14783 17
rect 14817 -17 14908 17
rect -34 -34 14908 -17
<< nsubdiff >>
rect -34 1497 14908 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5163 1497
rect 5197 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5533 1497
rect 5567 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5755 1497
rect 5789 1463 5829 1497
rect 5863 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6125 1497
rect 6159 1463 6199 1497
rect 6233 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6495 1497
rect 6529 1463 6643 1497
rect 6677 1463 6717 1497
rect 6751 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7087 1497
rect 7121 1463 7161 1497
rect 7195 1463 7309 1497
rect 7343 1463 7383 1497
rect 7417 1463 7457 1497
rect 7491 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7679 1497
rect 7713 1463 7753 1497
rect 7787 1463 7827 1497
rect 7861 1463 7975 1497
rect 8009 1463 8049 1497
rect 8083 1463 8123 1497
rect 8157 1463 8197 1497
rect 8231 1463 8271 1497
rect 8305 1463 8345 1497
rect 8379 1463 8419 1497
rect 8453 1463 8493 1497
rect 8527 1463 8641 1497
rect 8675 1463 8715 1497
rect 8749 1463 8789 1497
rect 8823 1463 8863 1497
rect 8897 1463 8937 1497
rect 8971 1463 9011 1497
rect 9045 1463 9085 1497
rect 9119 1463 9159 1497
rect 9193 1463 9233 1497
rect 9267 1463 9307 1497
rect 9341 1463 9381 1497
rect 9415 1463 9455 1497
rect 9489 1463 9603 1497
rect 9637 1463 9677 1497
rect 9711 1463 9751 1497
rect 9785 1463 9825 1497
rect 9859 1463 9899 1497
rect 9933 1463 9973 1497
rect 10007 1463 10047 1497
rect 10081 1463 10121 1497
rect 10155 1463 10269 1497
rect 10303 1463 10343 1497
rect 10377 1463 10417 1497
rect 10451 1463 10491 1497
rect 10525 1463 10565 1497
rect 10599 1463 10639 1497
rect 10673 1463 10713 1497
rect 10747 1463 10787 1497
rect 10821 1463 10935 1497
rect 10969 1463 11009 1497
rect 11043 1463 11083 1497
rect 11117 1463 11157 1497
rect 11191 1463 11231 1497
rect 11265 1463 11305 1497
rect 11339 1463 11379 1497
rect 11413 1463 11453 1497
rect 11487 1463 11601 1497
rect 11635 1463 11675 1497
rect 11709 1463 11749 1497
rect 11783 1463 11823 1497
rect 11857 1463 11897 1497
rect 11931 1463 11971 1497
rect 12005 1463 12045 1497
rect 12079 1463 12119 1497
rect 12153 1463 12267 1497
rect 12301 1463 12341 1497
rect 12375 1463 12415 1497
rect 12449 1463 12489 1497
rect 12523 1463 12563 1497
rect 12597 1463 12637 1497
rect 12671 1463 12711 1497
rect 12745 1463 12785 1497
rect 12819 1463 12933 1497
rect 12967 1463 13007 1497
rect 13041 1463 13081 1497
rect 13115 1463 13155 1497
rect 13189 1463 13229 1497
rect 13263 1463 13303 1497
rect 13337 1463 13377 1497
rect 13411 1463 13451 1497
rect 13485 1463 13599 1497
rect 13633 1463 13673 1497
rect 13707 1463 13747 1497
rect 13781 1463 13821 1497
rect 13855 1463 13895 1497
rect 13929 1463 13969 1497
rect 14003 1463 14043 1497
rect 14077 1463 14117 1497
rect 14151 1463 14265 1497
rect 14299 1463 14339 1497
rect 14373 1463 14413 1497
rect 14447 1463 14487 1497
rect 14521 1463 14561 1497
rect 14595 1463 14635 1497
rect 14669 1463 14709 1497
rect 14743 1463 14783 1497
rect 14817 1463 14908 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 928 1423 996 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 1594 1423 1662 1463
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect 928 1019 945 1053
rect 979 1019 996 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 928 979 996 1019
rect 1594 1389 1611 1423
rect 1645 1389 1662 1423
rect 2260 1423 2328 1463
rect 1594 1349 1662 1389
rect 1594 1315 1611 1349
rect 1645 1315 1662 1349
rect 1594 1275 1662 1315
rect 1594 1241 1611 1275
rect 1645 1241 1662 1275
rect 1594 1201 1662 1241
rect 1594 1167 1611 1201
rect 1645 1167 1662 1201
rect 1594 1127 1662 1167
rect 1594 1093 1611 1127
rect 1645 1093 1662 1127
rect 1594 1053 1662 1093
rect 1594 1019 1611 1053
rect 1645 1019 1662 1053
rect 928 945 945 979
rect 979 945 996 979
rect -34 871 -17 905
rect 17 884 34 905
rect 928 905 996 945
rect 1594 979 1662 1019
rect 2260 1389 2277 1423
rect 2311 1389 2328 1423
rect 2926 1423 2994 1463
rect 2260 1349 2328 1389
rect 2260 1315 2277 1349
rect 2311 1315 2328 1349
rect 2260 1275 2328 1315
rect 2260 1241 2277 1275
rect 2311 1241 2328 1275
rect 2260 1201 2328 1241
rect 2260 1167 2277 1201
rect 2311 1167 2328 1201
rect 2260 1127 2328 1167
rect 2260 1093 2277 1127
rect 2311 1093 2328 1127
rect 2260 1053 2328 1093
rect 2260 1019 2277 1053
rect 2311 1019 2328 1053
rect 1594 945 1611 979
rect 1645 945 1662 979
rect 928 884 945 905
rect 17 871 945 884
rect 979 884 996 905
rect 1594 905 1662 945
rect 2260 979 2328 1019
rect 2926 1389 2943 1423
rect 2977 1389 2994 1423
rect 3592 1423 3660 1463
rect 2926 1349 2994 1389
rect 2926 1315 2943 1349
rect 2977 1315 2994 1349
rect 2926 1275 2994 1315
rect 2926 1241 2943 1275
rect 2977 1241 2994 1275
rect 2926 1201 2994 1241
rect 2926 1167 2943 1201
rect 2977 1167 2994 1201
rect 2926 1127 2994 1167
rect 2926 1093 2943 1127
rect 2977 1093 2994 1127
rect 2926 1053 2994 1093
rect 2926 1019 2943 1053
rect 2977 1019 2994 1053
rect 2260 945 2277 979
rect 2311 945 2328 979
rect 1594 884 1611 905
rect 979 871 1611 884
rect 1645 884 1662 905
rect 2260 905 2328 945
rect 2926 979 2994 1019
rect 3592 1389 3609 1423
rect 3643 1389 3660 1423
rect 4258 1423 4326 1463
rect 3592 1349 3660 1389
rect 3592 1315 3609 1349
rect 3643 1315 3660 1349
rect 3592 1275 3660 1315
rect 3592 1241 3609 1275
rect 3643 1241 3660 1275
rect 3592 1201 3660 1241
rect 3592 1167 3609 1201
rect 3643 1167 3660 1201
rect 3592 1127 3660 1167
rect 3592 1093 3609 1127
rect 3643 1093 3660 1127
rect 3592 1053 3660 1093
rect 3592 1019 3609 1053
rect 3643 1019 3660 1053
rect 2926 945 2943 979
rect 2977 945 2994 979
rect 2260 884 2277 905
rect 1645 871 2277 884
rect 2311 884 2328 905
rect 2926 905 2994 945
rect 3592 979 3660 1019
rect 4258 1389 4275 1423
rect 4309 1389 4326 1423
rect 5220 1423 5288 1463
rect 4258 1349 4326 1389
rect 4258 1315 4275 1349
rect 4309 1315 4326 1349
rect 4258 1275 4326 1315
rect 4258 1241 4275 1275
rect 4309 1241 4326 1275
rect 4258 1201 4326 1241
rect 4258 1167 4275 1201
rect 4309 1167 4326 1201
rect 4258 1127 4326 1167
rect 4258 1093 4275 1127
rect 4309 1093 4326 1127
rect 4258 1053 4326 1093
rect 4258 1019 4275 1053
rect 4309 1019 4326 1053
rect 3592 945 3609 979
rect 3643 945 3660 979
rect 2926 884 2943 905
rect 2311 871 2943 884
rect 2977 884 2994 905
rect 3592 905 3660 945
rect 4258 979 4326 1019
rect 5220 1389 5237 1423
rect 5271 1389 5288 1423
rect 5886 1423 5954 1463
rect 5220 1349 5288 1389
rect 5220 1315 5237 1349
rect 5271 1315 5288 1349
rect 5220 1275 5288 1315
rect 5220 1241 5237 1275
rect 5271 1241 5288 1275
rect 5220 1201 5288 1241
rect 5220 1167 5237 1201
rect 5271 1167 5288 1201
rect 5220 1127 5288 1167
rect 5220 1093 5237 1127
rect 5271 1093 5288 1127
rect 5220 1053 5288 1093
rect 5220 1019 5237 1053
rect 5271 1019 5288 1053
rect 4258 945 4275 979
rect 4309 945 4326 979
rect 3592 884 3609 905
rect 2977 871 3609 884
rect 3643 884 3660 905
rect 4258 905 4326 945
rect 5220 979 5288 1019
rect 5886 1389 5903 1423
rect 5937 1389 5954 1423
rect 6552 1423 6620 1463
rect 5886 1349 5954 1389
rect 5886 1315 5903 1349
rect 5937 1315 5954 1349
rect 5886 1275 5954 1315
rect 5886 1241 5903 1275
rect 5937 1241 5954 1275
rect 5886 1201 5954 1241
rect 5886 1167 5903 1201
rect 5937 1167 5954 1201
rect 5886 1127 5954 1167
rect 5886 1093 5903 1127
rect 5937 1093 5954 1127
rect 5886 1053 5954 1093
rect 5886 1019 5903 1053
rect 5937 1019 5954 1053
rect 5220 945 5237 979
rect 5271 945 5288 979
rect 4258 884 4275 905
rect 3643 871 4275 884
rect 4309 884 4326 905
rect 5220 905 5288 945
rect 5886 979 5954 1019
rect 6552 1389 6569 1423
rect 6603 1389 6620 1423
rect 7218 1423 7286 1463
rect 6552 1349 6620 1389
rect 6552 1315 6569 1349
rect 6603 1315 6620 1349
rect 6552 1275 6620 1315
rect 6552 1241 6569 1275
rect 6603 1241 6620 1275
rect 6552 1201 6620 1241
rect 6552 1167 6569 1201
rect 6603 1167 6620 1201
rect 6552 1127 6620 1167
rect 6552 1093 6569 1127
rect 6603 1093 6620 1127
rect 6552 1053 6620 1093
rect 6552 1019 6569 1053
rect 6603 1019 6620 1053
rect 5886 945 5903 979
rect 5937 945 5954 979
rect 5220 884 5237 905
rect 4309 871 5237 884
rect 5271 884 5288 905
rect 5886 905 5954 945
rect 6552 979 6620 1019
rect 7218 1389 7235 1423
rect 7269 1389 7286 1423
rect 7884 1423 7952 1463
rect 7218 1349 7286 1389
rect 7218 1315 7235 1349
rect 7269 1315 7286 1349
rect 7218 1275 7286 1315
rect 7218 1241 7235 1275
rect 7269 1241 7286 1275
rect 7218 1201 7286 1241
rect 7218 1167 7235 1201
rect 7269 1167 7286 1201
rect 7218 1127 7286 1167
rect 7218 1093 7235 1127
rect 7269 1093 7286 1127
rect 7218 1053 7286 1093
rect 7218 1019 7235 1053
rect 7269 1019 7286 1053
rect 6552 945 6569 979
rect 6603 945 6620 979
rect 5886 884 5903 905
rect 5271 871 5903 884
rect 5937 884 5954 905
rect 6552 905 6620 945
rect 7218 979 7286 1019
rect 7884 1389 7901 1423
rect 7935 1389 7952 1423
rect 8550 1423 8618 1463
rect 7884 1349 7952 1389
rect 7884 1315 7901 1349
rect 7935 1315 7952 1349
rect 7884 1275 7952 1315
rect 7884 1241 7901 1275
rect 7935 1241 7952 1275
rect 7884 1201 7952 1241
rect 7884 1167 7901 1201
rect 7935 1167 7952 1201
rect 7884 1127 7952 1167
rect 7884 1093 7901 1127
rect 7935 1093 7952 1127
rect 7884 1053 7952 1093
rect 7884 1019 7901 1053
rect 7935 1019 7952 1053
rect 7218 945 7235 979
rect 7269 945 7286 979
rect 6552 884 6569 905
rect 5937 871 6569 884
rect 6603 884 6620 905
rect 7218 905 7286 945
rect 7884 979 7952 1019
rect 8550 1389 8567 1423
rect 8601 1389 8618 1423
rect 9512 1423 9580 1463
rect 8550 1349 8618 1389
rect 8550 1315 8567 1349
rect 8601 1315 8618 1349
rect 8550 1275 8618 1315
rect 8550 1241 8567 1275
rect 8601 1241 8618 1275
rect 8550 1201 8618 1241
rect 8550 1167 8567 1201
rect 8601 1167 8618 1201
rect 8550 1127 8618 1167
rect 8550 1093 8567 1127
rect 8601 1093 8618 1127
rect 8550 1053 8618 1093
rect 8550 1019 8567 1053
rect 8601 1019 8618 1053
rect 7884 945 7901 979
rect 7935 945 7952 979
rect 7218 884 7235 905
rect 6603 871 7235 884
rect 7269 884 7286 905
rect 7884 905 7952 945
rect 8550 979 8618 1019
rect 9512 1389 9529 1423
rect 9563 1389 9580 1423
rect 10178 1423 10246 1463
rect 9512 1349 9580 1389
rect 9512 1315 9529 1349
rect 9563 1315 9580 1349
rect 9512 1275 9580 1315
rect 9512 1241 9529 1275
rect 9563 1241 9580 1275
rect 9512 1201 9580 1241
rect 9512 1167 9529 1201
rect 9563 1167 9580 1201
rect 9512 1127 9580 1167
rect 9512 1093 9529 1127
rect 9563 1093 9580 1127
rect 9512 1053 9580 1093
rect 9512 1019 9529 1053
rect 9563 1019 9580 1053
rect 8550 945 8567 979
rect 8601 945 8618 979
rect 7884 884 7901 905
rect 7269 871 7901 884
rect 7935 884 7952 905
rect 8550 905 8618 945
rect 9512 979 9580 1019
rect 10178 1389 10195 1423
rect 10229 1389 10246 1423
rect 10844 1423 10912 1463
rect 10178 1349 10246 1389
rect 10178 1315 10195 1349
rect 10229 1315 10246 1349
rect 10178 1275 10246 1315
rect 10178 1241 10195 1275
rect 10229 1241 10246 1275
rect 10178 1201 10246 1241
rect 10178 1167 10195 1201
rect 10229 1167 10246 1201
rect 10178 1127 10246 1167
rect 10178 1093 10195 1127
rect 10229 1093 10246 1127
rect 10178 1053 10246 1093
rect 10178 1019 10195 1053
rect 10229 1019 10246 1053
rect 9512 945 9529 979
rect 9563 945 9580 979
rect 8550 884 8567 905
rect 7935 871 8567 884
rect 8601 884 8618 905
rect 9512 905 9580 945
rect 10178 979 10246 1019
rect 10844 1389 10861 1423
rect 10895 1389 10912 1423
rect 11510 1423 11578 1463
rect 10844 1349 10912 1389
rect 10844 1315 10861 1349
rect 10895 1315 10912 1349
rect 10844 1275 10912 1315
rect 10844 1241 10861 1275
rect 10895 1241 10912 1275
rect 10844 1201 10912 1241
rect 10844 1167 10861 1201
rect 10895 1167 10912 1201
rect 10844 1127 10912 1167
rect 10844 1093 10861 1127
rect 10895 1093 10912 1127
rect 10844 1053 10912 1093
rect 10844 1019 10861 1053
rect 10895 1019 10912 1053
rect 10178 945 10195 979
rect 10229 945 10246 979
rect 9512 884 9529 905
rect 8601 871 9529 884
rect 9563 884 9580 905
rect 10178 905 10246 945
rect 10844 979 10912 1019
rect 11510 1389 11527 1423
rect 11561 1389 11578 1423
rect 12176 1423 12244 1463
rect 11510 1349 11578 1389
rect 11510 1315 11527 1349
rect 11561 1315 11578 1349
rect 11510 1275 11578 1315
rect 11510 1241 11527 1275
rect 11561 1241 11578 1275
rect 11510 1201 11578 1241
rect 11510 1167 11527 1201
rect 11561 1167 11578 1201
rect 11510 1127 11578 1167
rect 11510 1093 11527 1127
rect 11561 1093 11578 1127
rect 11510 1053 11578 1093
rect 11510 1019 11527 1053
rect 11561 1019 11578 1053
rect 10844 945 10861 979
rect 10895 945 10912 979
rect 10178 884 10195 905
rect 9563 871 10195 884
rect 10229 884 10246 905
rect 10844 905 10912 945
rect 11510 979 11578 1019
rect 12176 1389 12193 1423
rect 12227 1389 12244 1423
rect 12842 1423 12910 1463
rect 12176 1349 12244 1389
rect 12176 1315 12193 1349
rect 12227 1315 12244 1349
rect 12176 1275 12244 1315
rect 12176 1241 12193 1275
rect 12227 1241 12244 1275
rect 12176 1201 12244 1241
rect 12176 1167 12193 1201
rect 12227 1167 12244 1201
rect 12176 1127 12244 1167
rect 12176 1093 12193 1127
rect 12227 1093 12244 1127
rect 12176 1053 12244 1093
rect 12176 1019 12193 1053
rect 12227 1019 12244 1053
rect 11510 945 11527 979
rect 11561 945 11578 979
rect 10844 884 10861 905
rect 10229 871 10861 884
rect 10895 884 10912 905
rect 11510 905 11578 945
rect 12176 979 12244 1019
rect 12842 1389 12859 1423
rect 12893 1389 12910 1423
rect 13508 1423 13576 1463
rect 12842 1349 12910 1389
rect 12842 1315 12859 1349
rect 12893 1315 12910 1349
rect 12842 1275 12910 1315
rect 12842 1241 12859 1275
rect 12893 1241 12910 1275
rect 12842 1201 12910 1241
rect 12842 1167 12859 1201
rect 12893 1167 12910 1201
rect 12842 1127 12910 1167
rect 12842 1093 12859 1127
rect 12893 1093 12910 1127
rect 12842 1053 12910 1093
rect 12842 1019 12859 1053
rect 12893 1019 12910 1053
rect 12176 945 12193 979
rect 12227 945 12244 979
rect 11510 884 11527 905
rect 10895 871 11527 884
rect 11561 884 11578 905
rect 12176 905 12244 945
rect 12842 979 12910 1019
rect 13508 1389 13525 1423
rect 13559 1389 13576 1423
rect 14174 1423 14242 1463
rect 14822 1459 14908 1463
rect 13508 1349 13576 1389
rect 13508 1315 13525 1349
rect 13559 1315 13576 1349
rect 13508 1275 13576 1315
rect 13508 1241 13525 1275
rect 13559 1241 13576 1275
rect 13508 1201 13576 1241
rect 13508 1167 13525 1201
rect 13559 1167 13576 1201
rect 13508 1127 13576 1167
rect 13508 1093 13525 1127
rect 13559 1093 13576 1127
rect 13508 1053 13576 1093
rect 13508 1019 13525 1053
rect 13559 1019 13576 1053
rect 12842 945 12859 979
rect 12893 945 12910 979
rect 12176 884 12193 905
rect 11561 871 12193 884
rect 12227 884 12244 905
rect 12842 905 12910 945
rect 13508 979 13576 1019
rect 14174 1389 14191 1423
rect 14225 1389 14242 1423
rect 14840 1423 14908 1459
rect 14174 1349 14242 1389
rect 14174 1315 14191 1349
rect 14225 1315 14242 1349
rect 14174 1275 14242 1315
rect 14174 1241 14191 1275
rect 14225 1241 14242 1275
rect 14174 1201 14242 1241
rect 14174 1167 14191 1201
rect 14225 1167 14242 1201
rect 14174 1127 14242 1167
rect 14174 1093 14191 1127
rect 14225 1093 14242 1127
rect 14174 1053 14242 1093
rect 14174 1019 14191 1053
rect 14225 1019 14242 1053
rect 13508 945 13525 979
rect 13559 945 13576 979
rect 12842 884 12859 905
rect 12227 871 12859 884
rect 12893 884 12910 905
rect 13508 905 13576 945
rect 14174 979 14242 1019
rect 14840 1389 14857 1423
rect 14891 1389 14908 1423
rect 14840 1349 14908 1389
rect 14840 1315 14857 1349
rect 14891 1315 14908 1349
rect 14840 1275 14908 1315
rect 14840 1241 14857 1275
rect 14891 1241 14908 1275
rect 14840 1201 14908 1241
rect 14840 1167 14857 1201
rect 14891 1167 14908 1201
rect 14840 1127 14908 1167
rect 14840 1093 14857 1127
rect 14891 1093 14908 1127
rect 14840 1053 14908 1093
rect 14840 1019 14857 1053
rect 14891 1019 14908 1053
rect 14174 945 14191 979
rect 14225 945 14242 979
rect 13508 884 13525 905
rect 12893 871 13525 884
rect 13559 884 13576 905
rect 14174 905 14242 945
rect 14840 979 14908 1019
rect 14840 945 14857 979
rect 14891 945 14908 979
rect 14174 884 14191 905
rect 13559 871 14191 884
rect 14225 884 14242 905
rect 14840 905 14908 945
rect 14840 884 14857 905
rect 14225 871 14857 884
rect 14891 871 14908 905
rect -34 822 14908 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 945 427 979 461
rect 945 353 979 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1611 427 1645 461
rect 1611 353 1645 387
rect 945 279 979 313
rect 945 205 979 239
rect 945 131 979 165
rect 945 57 979 91
rect 2277 427 2311 461
rect 2277 353 2311 387
rect 1611 279 1645 313
rect 1611 205 1645 239
rect 1611 131 1645 165
rect 1611 57 1645 91
rect 2943 427 2977 461
rect 2943 353 2977 387
rect 2277 279 2311 313
rect 2277 205 2311 239
rect 2277 131 2311 165
rect 2277 57 2311 91
rect 3609 427 3643 461
rect 3609 353 3643 387
rect 2943 279 2977 313
rect 2943 205 2977 239
rect 2943 131 2977 165
rect 2943 57 2977 91
rect 4275 427 4309 461
rect 4275 353 4309 387
rect 3609 279 3643 313
rect 3609 205 3643 239
rect 3609 131 3643 165
rect 3609 57 3643 91
rect 5237 427 5271 461
rect 5237 353 5271 387
rect 4275 279 4309 313
rect 4275 205 4309 239
rect 4275 131 4309 165
rect 4275 57 4309 91
rect 5903 427 5937 461
rect 5903 353 5937 387
rect 5237 279 5271 313
rect 5237 205 5271 239
rect 5237 131 5271 165
rect 5237 57 5271 91
rect 6569 427 6603 461
rect 6569 353 6603 387
rect 5903 279 5937 313
rect 5903 205 5937 239
rect 5903 131 5937 165
rect 5903 57 5937 91
rect 7235 427 7269 461
rect 7235 353 7269 387
rect 6569 279 6603 313
rect 6569 205 6603 239
rect 6569 131 6603 165
rect 6569 57 6603 91
rect 7901 427 7935 461
rect 7901 353 7935 387
rect 7235 279 7269 313
rect 7235 205 7269 239
rect 7235 131 7269 165
rect 7235 57 7269 91
rect 8567 427 8601 461
rect 8567 353 8601 387
rect 7901 279 7935 313
rect 7901 205 7935 239
rect 7901 131 7935 165
rect 7901 57 7935 91
rect 9529 427 9563 461
rect 9529 353 9563 387
rect 8567 279 8601 313
rect 8567 205 8601 239
rect 8567 131 8601 165
rect 8567 57 8601 91
rect 10195 427 10229 461
rect 10195 353 10229 387
rect 9529 279 9563 313
rect 9529 205 9563 239
rect 9529 131 9563 165
rect 9529 57 9563 91
rect 10861 427 10895 461
rect 10861 353 10895 387
rect 10195 279 10229 313
rect 10195 205 10229 239
rect 10195 131 10229 165
rect 10195 57 10229 91
rect 11527 427 11561 461
rect 11527 353 11561 387
rect 10861 279 10895 313
rect 10861 205 10895 239
rect 10861 131 10895 165
rect 10861 57 10895 91
rect 12193 427 12227 461
rect 12193 353 12227 387
rect 11527 279 11561 313
rect 11527 205 11561 239
rect 11527 131 11561 165
rect 11527 57 11561 91
rect 12859 427 12893 461
rect 12859 353 12893 387
rect 13525 427 13559 461
rect 12193 279 12227 313
rect 12193 205 12227 239
rect 12193 131 12227 165
rect 12193 57 12227 91
rect 13525 353 13559 387
rect 12859 279 12893 313
rect 12859 205 12893 239
rect 12859 131 12893 165
rect 12859 57 12893 91
rect 14191 427 14225 461
rect 14191 353 14225 387
rect 14857 427 14891 461
rect 13525 279 13559 313
rect 13525 205 13559 239
rect 13525 131 13559 165
rect 13525 57 13559 91
rect 14857 353 14891 387
rect 14191 279 14225 313
rect 14191 205 14225 239
rect 14191 131 14225 165
rect 14191 57 14225 91
rect 14857 279 14891 313
rect 14857 205 14891 239
rect 14857 131 14891 165
rect 14857 57 14891 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4497 -17 4531 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4793 -17 4827 17
rect 4867 -17 4901 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5089 -17 5123 17
rect 5163 -17 5197 17
rect 5311 -17 5345 17
rect 5385 -17 5419 17
rect 5459 -17 5493 17
rect 5533 -17 5567 17
rect 5607 -17 5641 17
rect 5681 -17 5715 17
rect 5755 -17 5789 17
rect 5829 -17 5863 17
rect 5977 -17 6011 17
rect 6051 -17 6085 17
rect 6125 -17 6159 17
rect 6199 -17 6233 17
rect 6273 -17 6307 17
rect 6347 -17 6381 17
rect 6421 -17 6455 17
rect 6495 -17 6529 17
rect 6643 -17 6677 17
rect 6717 -17 6751 17
rect 6791 -17 6825 17
rect 6865 -17 6899 17
rect 6939 -17 6973 17
rect 7013 -17 7047 17
rect 7087 -17 7121 17
rect 7161 -17 7195 17
rect 7309 -17 7343 17
rect 7383 -17 7417 17
rect 7457 -17 7491 17
rect 7531 -17 7565 17
rect 7605 -17 7639 17
rect 7679 -17 7713 17
rect 7753 -17 7787 17
rect 7827 -17 7861 17
rect 7975 -17 8009 17
rect 8049 -17 8083 17
rect 8123 -17 8157 17
rect 8197 -17 8231 17
rect 8271 -17 8305 17
rect 8345 -17 8379 17
rect 8419 -17 8453 17
rect 8493 -17 8527 17
rect 8641 -17 8675 17
rect 8715 -17 8749 17
rect 8789 -17 8823 17
rect 8863 -17 8897 17
rect 8937 -17 8971 17
rect 9011 -17 9045 17
rect 9085 -17 9119 17
rect 9159 -17 9193 17
rect 9233 -17 9267 17
rect 9307 -17 9341 17
rect 9381 -17 9415 17
rect 9455 -17 9489 17
rect 9603 -17 9637 17
rect 9677 -17 9711 17
rect 9751 -17 9785 17
rect 9825 -17 9859 17
rect 9899 -17 9933 17
rect 9973 -17 10007 17
rect 10047 -17 10081 17
rect 10121 -17 10155 17
rect 10269 -17 10303 17
rect 10343 -17 10377 17
rect 10417 -17 10451 17
rect 10491 -17 10525 17
rect 10565 -17 10599 17
rect 10639 -17 10673 17
rect 10713 -17 10747 17
rect 10787 -17 10821 17
rect 10935 -17 10969 17
rect 11009 -17 11043 17
rect 11083 -17 11117 17
rect 11157 -17 11191 17
rect 11231 -17 11265 17
rect 11305 -17 11339 17
rect 11379 -17 11413 17
rect 11453 -17 11487 17
rect 11601 -17 11635 17
rect 11675 -17 11709 17
rect 11749 -17 11783 17
rect 11823 -17 11857 17
rect 11897 -17 11931 17
rect 11971 -17 12005 17
rect 12045 -17 12079 17
rect 12119 -17 12153 17
rect 12267 -17 12301 17
rect 12341 -17 12375 17
rect 12415 -17 12449 17
rect 12489 -17 12523 17
rect 12563 -17 12597 17
rect 12637 -17 12671 17
rect 12711 -17 12745 17
rect 12785 -17 12819 17
rect 12933 -17 12967 17
rect 13007 -17 13041 17
rect 13081 -17 13115 17
rect 13155 -17 13189 17
rect 13229 -17 13263 17
rect 13303 -17 13337 17
rect 13377 -17 13411 17
rect 13451 -17 13485 17
rect 13599 -17 13633 17
rect 13673 -17 13707 17
rect 13747 -17 13781 17
rect 13821 -17 13855 17
rect 13895 -17 13929 17
rect 13969 -17 14003 17
rect 14043 -17 14077 17
rect 14117 -17 14151 17
rect 14265 -17 14299 17
rect 14339 -17 14373 17
rect 14413 -17 14447 17
rect 14487 -17 14521 17
rect 14561 -17 14595 17
rect 14635 -17 14669 17
rect 14709 -17 14743 17
rect 14783 -17 14817 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4497 1463 4531 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4793 1463 4827 1497
rect 4867 1463 4901 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5089 1463 5123 1497
rect 5163 1463 5197 1497
rect 5311 1463 5345 1497
rect 5385 1463 5419 1497
rect 5459 1463 5493 1497
rect 5533 1463 5567 1497
rect 5607 1463 5641 1497
rect 5681 1463 5715 1497
rect 5755 1463 5789 1497
rect 5829 1463 5863 1497
rect 5977 1463 6011 1497
rect 6051 1463 6085 1497
rect 6125 1463 6159 1497
rect 6199 1463 6233 1497
rect 6273 1463 6307 1497
rect 6347 1463 6381 1497
rect 6421 1463 6455 1497
rect 6495 1463 6529 1497
rect 6643 1463 6677 1497
rect 6717 1463 6751 1497
rect 6791 1463 6825 1497
rect 6865 1463 6899 1497
rect 6939 1463 6973 1497
rect 7013 1463 7047 1497
rect 7087 1463 7121 1497
rect 7161 1463 7195 1497
rect 7309 1463 7343 1497
rect 7383 1463 7417 1497
rect 7457 1463 7491 1497
rect 7531 1463 7565 1497
rect 7605 1463 7639 1497
rect 7679 1463 7713 1497
rect 7753 1463 7787 1497
rect 7827 1463 7861 1497
rect 7975 1463 8009 1497
rect 8049 1463 8083 1497
rect 8123 1463 8157 1497
rect 8197 1463 8231 1497
rect 8271 1463 8305 1497
rect 8345 1463 8379 1497
rect 8419 1463 8453 1497
rect 8493 1463 8527 1497
rect 8641 1463 8675 1497
rect 8715 1463 8749 1497
rect 8789 1463 8823 1497
rect 8863 1463 8897 1497
rect 8937 1463 8971 1497
rect 9011 1463 9045 1497
rect 9085 1463 9119 1497
rect 9159 1463 9193 1497
rect 9233 1463 9267 1497
rect 9307 1463 9341 1497
rect 9381 1463 9415 1497
rect 9455 1463 9489 1497
rect 9603 1463 9637 1497
rect 9677 1463 9711 1497
rect 9751 1463 9785 1497
rect 9825 1463 9859 1497
rect 9899 1463 9933 1497
rect 9973 1463 10007 1497
rect 10047 1463 10081 1497
rect 10121 1463 10155 1497
rect 10269 1463 10303 1497
rect 10343 1463 10377 1497
rect 10417 1463 10451 1497
rect 10491 1463 10525 1497
rect 10565 1463 10599 1497
rect 10639 1463 10673 1497
rect 10713 1463 10747 1497
rect 10787 1463 10821 1497
rect 10935 1463 10969 1497
rect 11009 1463 11043 1497
rect 11083 1463 11117 1497
rect 11157 1463 11191 1497
rect 11231 1463 11265 1497
rect 11305 1463 11339 1497
rect 11379 1463 11413 1497
rect 11453 1463 11487 1497
rect 11601 1463 11635 1497
rect 11675 1463 11709 1497
rect 11749 1463 11783 1497
rect 11823 1463 11857 1497
rect 11897 1463 11931 1497
rect 11971 1463 12005 1497
rect 12045 1463 12079 1497
rect 12119 1463 12153 1497
rect 12267 1463 12301 1497
rect 12341 1463 12375 1497
rect 12415 1463 12449 1497
rect 12489 1463 12523 1497
rect 12563 1463 12597 1497
rect 12637 1463 12671 1497
rect 12711 1463 12745 1497
rect 12785 1463 12819 1497
rect 12933 1463 12967 1497
rect 13007 1463 13041 1497
rect 13081 1463 13115 1497
rect 13155 1463 13189 1497
rect 13229 1463 13263 1497
rect 13303 1463 13337 1497
rect 13377 1463 13411 1497
rect 13451 1463 13485 1497
rect 13599 1463 13633 1497
rect 13673 1463 13707 1497
rect 13747 1463 13781 1497
rect 13821 1463 13855 1497
rect 13895 1463 13929 1497
rect 13969 1463 14003 1497
rect 14043 1463 14077 1497
rect 14117 1463 14151 1497
rect 14265 1463 14299 1497
rect 14339 1463 14373 1497
rect 14413 1463 14447 1497
rect 14487 1463 14521 1497
rect 14561 1463 14595 1497
rect 14635 1463 14669 1497
rect 14709 1463 14743 1497
rect 14783 1463 14817 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 945 1389 979 1423
rect 945 1315 979 1349
rect 945 1241 979 1275
rect 945 1167 979 1201
rect 945 1093 979 1127
rect 945 1019 979 1053
rect -17 945 17 979
rect 1611 1389 1645 1423
rect 1611 1315 1645 1349
rect 1611 1241 1645 1275
rect 1611 1167 1645 1201
rect 1611 1093 1645 1127
rect 1611 1019 1645 1053
rect 945 945 979 979
rect -17 871 17 905
rect 2277 1389 2311 1423
rect 2277 1315 2311 1349
rect 2277 1241 2311 1275
rect 2277 1167 2311 1201
rect 2277 1093 2311 1127
rect 2277 1019 2311 1053
rect 1611 945 1645 979
rect 945 871 979 905
rect 2943 1389 2977 1423
rect 2943 1315 2977 1349
rect 2943 1241 2977 1275
rect 2943 1167 2977 1201
rect 2943 1093 2977 1127
rect 2943 1019 2977 1053
rect 2277 945 2311 979
rect 1611 871 1645 905
rect 3609 1389 3643 1423
rect 3609 1315 3643 1349
rect 3609 1241 3643 1275
rect 3609 1167 3643 1201
rect 3609 1093 3643 1127
rect 3609 1019 3643 1053
rect 2943 945 2977 979
rect 2277 871 2311 905
rect 4275 1389 4309 1423
rect 4275 1315 4309 1349
rect 4275 1241 4309 1275
rect 4275 1167 4309 1201
rect 4275 1093 4309 1127
rect 4275 1019 4309 1053
rect 3609 945 3643 979
rect 2943 871 2977 905
rect 5237 1389 5271 1423
rect 5237 1315 5271 1349
rect 5237 1241 5271 1275
rect 5237 1167 5271 1201
rect 5237 1093 5271 1127
rect 5237 1019 5271 1053
rect 4275 945 4309 979
rect 3609 871 3643 905
rect 5903 1389 5937 1423
rect 5903 1315 5937 1349
rect 5903 1241 5937 1275
rect 5903 1167 5937 1201
rect 5903 1093 5937 1127
rect 5903 1019 5937 1053
rect 5237 945 5271 979
rect 4275 871 4309 905
rect 6569 1389 6603 1423
rect 6569 1315 6603 1349
rect 6569 1241 6603 1275
rect 6569 1167 6603 1201
rect 6569 1093 6603 1127
rect 6569 1019 6603 1053
rect 5903 945 5937 979
rect 5237 871 5271 905
rect 7235 1389 7269 1423
rect 7235 1315 7269 1349
rect 7235 1241 7269 1275
rect 7235 1167 7269 1201
rect 7235 1093 7269 1127
rect 7235 1019 7269 1053
rect 6569 945 6603 979
rect 5903 871 5937 905
rect 7901 1389 7935 1423
rect 7901 1315 7935 1349
rect 7901 1241 7935 1275
rect 7901 1167 7935 1201
rect 7901 1093 7935 1127
rect 7901 1019 7935 1053
rect 7235 945 7269 979
rect 6569 871 6603 905
rect 8567 1389 8601 1423
rect 8567 1315 8601 1349
rect 8567 1241 8601 1275
rect 8567 1167 8601 1201
rect 8567 1093 8601 1127
rect 8567 1019 8601 1053
rect 7901 945 7935 979
rect 7235 871 7269 905
rect 9529 1389 9563 1423
rect 9529 1315 9563 1349
rect 9529 1241 9563 1275
rect 9529 1167 9563 1201
rect 9529 1093 9563 1127
rect 9529 1019 9563 1053
rect 8567 945 8601 979
rect 7901 871 7935 905
rect 10195 1389 10229 1423
rect 10195 1315 10229 1349
rect 10195 1241 10229 1275
rect 10195 1167 10229 1201
rect 10195 1093 10229 1127
rect 10195 1019 10229 1053
rect 9529 945 9563 979
rect 8567 871 8601 905
rect 10861 1389 10895 1423
rect 10861 1315 10895 1349
rect 10861 1241 10895 1275
rect 10861 1167 10895 1201
rect 10861 1093 10895 1127
rect 10861 1019 10895 1053
rect 10195 945 10229 979
rect 9529 871 9563 905
rect 11527 1389 11561 1423
rect 11527 1315 11561 1349
rect 11527 1241 11561 1275
rect 11527 1167 11561 1201
rect 11527 1093 11561 1127
rect 11527 1019 11561 1053
rect 10861 945 10895 979
rect 10195 871 10229 905
rect 12193 1389 12227 1423
rect 12193 1315 12227 1349
rect 12193 1241 12227 1275
rect 12193 1167 12227 1201
rect 12193 1093 12227 1127
rect 12193 1019 12227 1053
rect 11527 945 11561 979
rect 10861 871 10895 905
rect 12859 1389 12893 1423
rect 12859 1315 12893 1349
rect 12859 1241 12893 1275
rect 12859 1167 12893 1201
rect 12859 1093 12893 1127
rect 12859 1019 12893 1053
rect 12193 945 12227 979
rect 11527 871 11561 905
rect 13525 1389 13559 1423
rect 13525 1315 13559 1349
rect 13525 1241 13559 1275
rect 13525 1167 13559 1201
rect 13525 1093 13559 1127
rect 13525 1019 13559 1053
rect 12859 945 12893 979
rect 12193 871 12227 905
rect 14191 1389 14225 1423
rect 14191 1315 14225 1349
rect 14191 1241 14225 1275
rect 14191 1167 14225 1201
rect 14191 1093 14225 1127
rect 14191 1019 14225 1053
rect 13525 945 13559 979
rect 12859 871 12893 905
rect 14857 1389 14891 1423
rect 14857 1315 14891 1349
rect 14857 1241 14891 1275
rect 14857 1167 14891 1201
rect 14857 1093 14891 1127
rect 14857 1019 14891 1053
rect 14191 945 14225 979
rect 13525 871 13559 905
rect 14857 945 14891 979
rect 14191 871 14225 905
rect 14857 871 14891 905
<< poly >>
rect 247 1404 277 1430
rect 335 1404 365 1430
rect 423 1404 453 1430
rect 511 1404 541 1430
rect 599 1404 629 1430
rect 687 1404 717 1430
rect 1149 1404 1179 1430
rect 1237 1404 1267 1430
rect 1325 1404 1355 1430
rect 1413 1404 1443 1430
rect 247 973 277 1004
rect 335 973 365 1004
rect 423 973 453 1004
rect 511 973 541 1004
rect 195 957 365 973
rect 195 923 205 957
rect 239 943 365 957
rect 417 957 541 973
rect 239 923 249 943
rect 195 907 249 923
rect 417 923 427 957
rect 461 943 541 957
rect 599 973 629 1004
rect 687 973 717 1004
rect 599 957 717 973
rect 599 943 649 957
rect 461 923 471 943
rect 417 907 471 923
rect 639 923 649 943
rect 683 943 717 957
rect 1815 1404 1845 1430
rect 1903 1404 1933 1430
rect 1991 1404 2021 1430
rect 2079 1404 2109 1430
rect 683 923 693 943
rect 639 907 693 923
rect 1149 973 1179 1004
rect 1237 973 1267 1004
rect 1325 973 1355 1004
rect 1413 973 1443 1004
rect 1149 957 1267 973
rect 1149 943 1167 957
rect 1157 923 1167 943
rect 1201 943 1267 957
rect 1311 957 1443 973
rect 1201 923 1211 943
rect 1157 907 1211 923
rect 1311 923 1321 957
rect 1355 943 1443 957
rect 2481 1404 2511 1430
rect 2569 1404 2599 1430
rect 2657 1404 2687 1430
rect 2745 1404 2775 1430
rect 1355 923 1365 943
rect 1311 907 1365 923
rect 1815 973 1845 1004
rect 1903 973 1933 1004
rect 1991 973 2021 1004
rect 2079 973 2109 1004
rect 1815 957 1933 973
rect 1815 943 1833 957
rect 1823 923 1833 943
rect 1867 943 1933 957
rect 1977 957 2109 973
rect 1867 923 1877 943
rect 1823 907 1877 923
rect 1977 923 1987 957
rect 2021 943 2109 957
rect 3147 1404 3177 1430
rect 3235 1404 3265 1430
rect 3323 1404 3353 1430
rect 3411 1404 3441 1430
rect 2021 923 2031 943
rect 1977 907 2031 923
rect 2481 973 2511 1004
rect 2569 973 2599 1004
rect 2657 973 2687 1004
rect 2745 973 2775 1004
rect 2481 957 2599 973
rect 2481 943 2499 957
rect 2489 923 2499 943
rect 2533 943 2599 957
rect 2643 957 2775 973
rect 2533 923 2543 943
rect 2489 907 2543 923
rect 2643 923 2653 957
rect 2687 943 2775 957
rect 3813 1404 3843 1430
rect 3901 1404 3931 1430
rect 3989 1404 4019 1430
rect 4077 1404 4107 1430
rect 2687 923 2697 943
rect 2643 907 2697 923
rect 3147 973 3177 1004
rect 3235 973 3265 1004
rect 3323 973 3353 1004
rect 3411 973 3441 1004
rect 3147 957 3265 973
rect 3147 943 3165 957
rect 3155 923 3165 943
rect 3199 943 3265 957
rect 3309 957 3441 973
rect 3199 923 3209 943
rect 3155 907 3209 923
rect 3309 923 3319 957
rect 3353 943 3441 957
rect 4539 1404 4569 1430
rect 4627 1404 4657 1430
rect 4715 1404 4745 1430
rect 4803 1404 4833 1430
rect 4891 1404 4921 1430
rect 4979 1404 5009 1430
rect 3353 923 3363 943
rect 3309 907 3363 923
rect 3813 973 3843 1004
rect 3901 973 3931 1004
rect 3989 973 4019 1004
rect 4077 973 4107 1004
rect 3813 957 3931 973
rect 3813 943 3831 957
rect 3821 923 3831 943
rect 3865 943 3931 957
rect 3975 957 4107 973
rect 3865 923 3875 943
rect 3821 907 3875 923
rect 3975 923 3985 957
rect 4019 943 4107 957
rect 5441 1404 5471 1430
rect 5529 1404 5559 1430
rect 5617 1404 5647 1430
rect 5705 1404 5735 1430
rect 4539 973 4569 1004
rect 4627 973 4657 1004
rect 4715 973 4745 1004
rect 4803 973 4833 1004
rect 4019 923 4029 943
rect 3975 907 4029 923
rect 4487 957 4657 973
rect 4487 923 4497 957
rect 4531 943 4657 957
rect 4709 957 4833 973
rect 4531 923 4541 943
rect 4487 907 4541 923
rect 4709 923 4719 957
rect 4753 943 4833 957
rect 4891 973 4921 1004
rect 4979 973 5009 1004
rect 4891 957 5009 973
rect 4891 943 4941 957
rect 4753 923 4763 943
rect 4709 907 4763 923
rect 4931 923 4941 943
rect 4975 943 5009 957
rect 6107 1404 6137 1430
rect 6195 1404 6225 1430
rect 6283 1404 6313 1430
rect 6371 1404 6401 1430
rect 4975 923 4985 943
rect 4931 907 4985 923
rect 5441 973 5471 1004
rect 5529 973 5559 1004
rect 5617 973 5647 1004
rect 5705 973 5735 1004
rect 5441 957 5559 973
rect 5441 943 5459 957
rect 5449 923 5459 943
rect 5493 943 5559 957
rect 5603 957 5735 973
rect 5493 923 5503 943
rect 5449 907 5503 923
rect 5603 923 5613 957
rect 5647 943 5735 957
rect 6773 1404 6803 1430
rect 6861 1404 6891 1430
rect 6949 1404 6979 1430
rect 7037 1404 7067 1430
rect 5647 923 5657 943
rect 5603 907 5657 923
rect 6107 973 6137 1004
rect 6195 973 6225 1004
rect 6283 973 6313 1004
rect 6371 973 6401 1004
rect 6107 957 6225 973
rect 6107 943 6125 957
rect 6115 923 6125 943
rect 6159 943 6225 957
rect 6269 957 6401 973
rect 6159 923 6169 943
rect 6115 907 6169 923
rect 6269 923 6279 957
rect 6313 943 6401 957
rect 7439 1404 7469 1430
rect 7527 1404 7557 1430
rect 7615 1404 7645 1430
rect 7703 1404 7733 1430
rect 6313 923 6323 943
rect 6269 907 6323 923
rect 6773 973 6803 1004
rect 6861 973 6891 1004
rect 6949 973 6979 1004
rect 7037 973 7067 1004
rect 6773 957 6891 973
rect 6773 943 6791 957
rect 6781 923 6791 943
rect 6825 943 6891 957
rect 6935 957 7067 973
rect 6825 923 6835 943
rect 6781 907 6835 923
rect 6935 923 6945 957
rect 6979 943 7067 957
rect 8105 1404 8135 1430
rect 8193 1404 8223 1430
rect 8281 1404 8311 1430
rect 8369 1404 8399 1430
rect 6979 923 6989 943
rect 6935 907 6989 923
rect 7439 973 7469 1004
rect 7527 973 7557 1004
rect 7615 973 7645 1004
rect 7703 973 7733 1004
rect 7439 957 7557 973
rect 7439 943 7457 957
rect 7447 923 7457 943
rect 7491 943 7557 957
rect 7601 957 7733 973
rect 7491 923 7501 943
rect 7447 907 7501 923
rect 7601 923 7611 957
rect 7645 943 7733 957
rect 8831 1404 8861 1430
rect 8919 1404 8949 1430
rect 9007 1404 9037 1430
rect 9095 1404 9125 1430
rect 9183 1404 9213 1430
rect 9271 1404 9301 1430
rect 7645 923 7655 943
rect 7601 907 7655 923
rect 8105 973 8135 1004
rect 8193 973 8223 1004
rect 8281 973 8311 1004
rect 8369 973 8399 1004
rect 8105 957 8223 973
rect 8105 943 8123 957
rect 8113 923 8123 943
rect 8157 943 8223 957
rect 8267 957 8399 973
rect 8157 923 8167 943
rect 8113 907 8167 923
rect 8267 923 8277 957
rect 8311 943 8399 957
rect 9733 1404 9763 1430
rect 9821 1404 9851 1430
rect 9909 1404 9939 1430
rect 9997 1404 10027 1430
rect 8831 973 8861 1004
rect 8919 973 8949 1004
rect 9007 973 9037 1004
rect 9095 973 9125 1004
rect 8311 923 8321 943
rect 8267 907 8321 923
rect 8779 957 8949 973
rect 8779 923 8789 957
rect 8823 943 8949 957
rect 9001 957 9125 973
rect 8823 923 8833 943
rect 8779 907 8833 923
rect 9001 923 9011 957
rect 9045 943 9125 957
rect 9183 973 9213 1004
rect 9271 973 9301 1004
rect 9183 957 9301 973
rect 9183 943 9233 957
rect 9045 923 9055 943
rect 9001 907 9055 923
rect 9223 923 9233 943
rect 9267 943 9301 957
rect 10399 1404 10429 1430
rect 10487 1404 10517 1430
rect 10575 1404 10605 1430
rect 10663 1404 10693 1430
rect 9267 923 9277 943
rect 9223 907 9277 923
rect 9733 973 9763 1004
rect 9821 973 9851 1004
rect 9909 973 9939 1004
rect 9997 973 10027 1004
rect 9733 957 9851 973
rect 9733 943 9751 957
rect 9741 923 9751 943
rect 9785 943 9851 957
rect 9895 957 10027 973
rect 9785 923 9795 943
rect 9741 907 9795 923
rect 9895 923 9905 957
rect 9939 943 10027 957
rect 11065 1404 11095 1430
rect 11153 1404 11183 1430
rect 11241 1404 11271 1430
rect 11329 1404 11359 1430
rect 9939 923 9949 943
rect 9895 907 9949 923
rect 10399 973 10429 1004
rect 10487 973 10517 1004
rect 10575 973 10605 1004
rect 10663 973 10693 1004
rect 10399 957 10517 973
rect 10399 943 10417 957
rect 10407 923 10417 943
rect 10451 943 10517 957
rect 10561 957 10693 973
rect 10451 923 10461 943
rect 10407 907 10461 923
rect 10561 923 10571 957
rect 10605 943 10693 957
rect 11731 1404 11761 1430
rect 11819 1404 11849 1430
rect 11907 1404 11937 1430
rect 11995 1404 12025 1430
rect 10605 923 10615 943
rect 10561 907 10615 923
rect 11065 973 11095 1004
rect 11153 973 11183 1004
rect 11241 973 11271 1004
rect 11329 973 11359 1004
rect 11065 957 11183 973
rect 11065 943 11083 957
rect 11073 923 11083 943
rect 11117 943 11183 957
rect 11227 957 11359 973
rect 11117 923 11127 943
rect 11073 907 11127 923
rect 11227 923 11237 957
rect 11271 943 11359 957
rect 12397 1404 12427 1430
rect 12485 1404 12515 1430
rect 12573 1404 12603 1430
rect 12661 1404 12691 1430
rect 11271 923 11281 943
rect 11227 907 11281 923
rect 11731 973 11761 1004
rect 11819 973 11849 1004
rect 11907 973 11937 1004
rect 11995 973 12025 1004
rect 11731 957 11849 973
rect 11731 943 11749 957
rect 11739 923 11749 943
rect 11783 943 11849 957
rect 11893 957 12025 973
rect 11783 923 11793 943
rect 11739 907 11793 923
rect 11893 923 11903 957
rect 11937 943 12025 957
rect 13063 1405 13093 1431
rect 13151 1405 13181 1431
rect 13239 1405 13269 1431
rect 13327 1405 13357 1431
rect 11937 923 11947 943
rect 11893 907 11947 923
rect 12397 973 12427 1004
rect 12485 973 12515 1004
rect 12573 973 12603 1004
rect 12661 973 12691 1004
rect 12397 957 12515 973
rect 12397 943 12415 957
rect 12405 923 12415 943
rect 12449 943 12515 957
rect 12559 957 12691 973
rect 12449 923 12459 943
rect 12405 907 12459 923
rect 12559 923 12569 957
rect 12603 943 12691 957
rect 13727 1405 13757 1431
rect 13815 1405 13845 1431
rect 13903 1405 13933 1431
rect 13991 1405 14021 1431
rect 13063 974 13093 1005
rect 13151 974 13181 1005
rect 13239 974 13269 1005
rect 13327 974 13357 1005
rect 12603 923 12613 943
rect 12559 907 12613 923
rect 12997 958 13181 974
rect 12997 924 13007 958
rect 13041 944 13181 958
rect 13227 958 13357 974
rect 13041 924 13051 944
rect 12997 908 13051 924
rect 13227 924 13237 958
rect 13271 944 13357 958
rect 14395 1405 14425 1431
rect 14483 1405 14513 1431
rect 14571 1405 14601 1431
rect 14659 1405 14689 1431
rect 13271 924 13281 944
rect 13227 908 13281 924
rect 13727 974 13757 1005
rect 13815 974 13845 1005
rect 13727 958 13845 974
rect 13727 944 13747 958
rect 13737 924 13747 944
rect 13781 944 13845 958
rect 13903 974 13933 1005
rect 13991 974 14021 1005
rect 13903 958 14087 974
rect 13903 944 14043 958
rect 13781 924 13791 944
rect 13737 908 13791 924
rect 14033 924 14043 944
rect 14077 924 14087 958
rect 14033 908 14087 924
rect 14395 974 14425 1005
rect 14483 974 14513 1005
rect 14571 974 14601 1005
rect 14659 974 14689 1005
rect 14329 958 14513 974
rect 14329 924 14339 958
rect 14373 944 14513 958
rect 14555 958 14689 974
rect 14373 924 14383 944
rect 14329 908 14383 924
rect 14555 924 14565 958
rect 14599 944 14689 958
rect 14599 924 14609 944
rect 14555 908 14609 924
rect 195 433 249 449
rect 195 413 205 433
rect 147 399 205 413
rect 239 399 249 433
rect 147 383 249 399
rect 417 433 471 449
rect 417 399 427 433
rect 461 413 471 433
rect 639 433 693 449
rect 461 399 477 413
rect 417 383 477 399
rect 639 399 649 433
rect 683 399 693 433
rect 639 383 693 399
rect 1157 433 1211 449
rect 1157 413 1167 433
rect 147 351 177 383
rect 447 351 477 383
rect 649 351 679 383
rect 1130 399 1167 413
rect 1201 399 1211 433
rect 1130 383 1211 399
rect 1305 433 1359 449
rect 1305 399 1315 433
rect 1349 399 1359 433
rect 1305 383 1359 399
rect 1823 433 1877 449
rect 1823 413 1833 433
rect 1130 349 1160 383
rect 1324 349 1354 383
rect 1796 399 1833 413
rect 1867 399 1877 433
rect 1796 383 1877 399
rect 1971 433 2025 449
rect 1971 399 1981 433
rect 2015 399 2025 433
rect 1971 383 2025 399
rect 2489 433 2543 449
rect 2489 413 2499 433
rect 1796 349 1826 383
rect 1990 349 2020 383
rect 2462 399 2499 413
rect 2533 399 2543 433
rect 2462 383 2543 399
rect 2637 433 2691 449
rect 2637 399 2647 433
rect 2681 399 2691 433
rect 2637 383 2691 399
rect 3155 433 3209 449
rect 3155 413 3165 433
rect 2462 349 2492 383
rect 2656 349 2686 383
rect 3128 399 3165 413
rect 3199 399 3209 433
rect 3128 383 3209 399
rect 3303 433 3357 449
rect 3303 399 3313 433
rect 3347 399 3357 433
rect 3303 383 3357 399
rect 3821 433 3875 449
rect 3821 413 3831 433
rect 3128 349 3158 383
rect 3322 349 3352 383
rect 3794 399 3831 413
rect 3865 399 3875 433
rect 3794 383 3875 399
rect 3969 433 4023 449
rect 3969 399 3979 433
rect 4013 399 4023 433
rect 3969 383 4023 399
rect 4487 433 4541 449
rect 4487 413 4497 433
rect 3794 349 3824 383
rect 3988 349 4018 383
rect 4439 399 4497 413
rect 4531 399 4541 433
rect 4439 383 4541 399
rect 4709 433 4763 449
rect 4709 399 4719 433
rect 4753 413 4763 433
rect 4931 433 4985 449
rect 4753 399 4769 413
rect 4709 383 4769 399
rect 4931 399 4941 433
rect 4975 399 4985 433
rect 4931 383 4985 399
rect 5449 433 5503 449
rect 5449 413 5459 433
rect 4439 351 4469 383
rect 4739 351 4769 383
rect 4941 351 4971 383
rect 5422 399 5459 413
rect 5493 399 5503 433
rect 5422 383 5503 399
rect 5597 433 5651 449
rect 5597 399 5607 433
rect 5641 399 5651 433
rect 5597 383 5651 399
rect 6115 433 6169 449
rect 6115 413 6125 433
rect 5422 349 5452 383
rect 5616 349 5646 383
rect 6088 399 6125 413
rect 6159 399 6169 433
rect 6088 383 6169 399
rect 6263 433 6317 449
rect 6263 399 6273 433
rect 6307 399 6317 433
rect 6263 383 6317 399
rect 6781 433 6835 449
rect 6781 413 6791 433
rect 6088 349 6118 383
rect 6282 349 6312 383
rect 6754 399 6791 413
rect 6825 399 6835 433
rect 6754 383 6835 399
rect 6929 433 6983 449
rect 6929 399 6939 433
rect 6973 399 6983 433
rect 6929 383 6983 399
rect 7447 433 7501 449
rect 7447 413 7457 433
rect 6754 349 6784 383
rect 6948 349 6978 383
rect 7420 399 7457 413
rect 7491 399 7501 433
rect 7420 383 7501 399
rect 7595 433 7649 449
rect 7595 399 7605 433
rect 7639 399 7649 433
rect 7595 383 7649 399
rect 8113 433 8167 449
rect 8113 413 8123 433
rect 7420 349 7450 383
rect 7614 349 7644 383
rect 8086 399 8123 413
rect 8157 399 8167 433
rect 8086 383 8167 399
rect 8261 433 8315 449
rect 8261 399 8271 433
rect 8305 399 8315 433
rect 8261 383 8315 399
rect 8779 433 8833 449
rect 8779 413 8789 433
rect 8086 349 8116 383
rect 8280 349 8310 383
rect 8731 399 8789 413
rect 8823 399 8833 433
rect 8731 383 8833 399
rect 9001 433 9055 449
rect 9001 399 9011 433
rect 9045 413 9055 433
rect 9223 433 9277 449
rect 9045 399 9061 413
rect 9001 383 9061 399
rect 9223 399 9233 433
rect 9267 399 9277 433
rect 9223 383 9277 399
rect 9741 433 9795 449
rect 9741 413 9751 433
rect 8731 351 8761 383
rect 9031 351 9061 383
rect 9233 351 9263 383
rect 9714 399 9751 413
rect 9785 399 9795 433
rect 9714 383 9795 399
rect 9889 433 9943 449
rect 9889 399 9899 433
rect 9933 399 9943 433
rect 9889 383 9943 399
rect 10407 433 10461 449
rect 10407 413 10417 433
rect 9714 349 9744 383
rect 9908 349 9938 383
rect 10380 399 10417 413
rect 10451 399 10461 433
rect 10380 383 10461 399
rect 10555 433 10609 449
rect 10555 399 10565 433
rect 10599 399 10609 433
rect 10555 383 10609 399
rect 11073 433 11127 449
rect 11073 413 11083 433
rect 10380 349 10410 383
rect 10574 349 10604 383
rect 11046 399 11083 413
rect 11117 399 11127 433
rect 11046 383 11127 399
rect 11221 433 11275 449
rect 11221 399 11231 433
rect 11265 399 11275 433
rect 11221 383 11275 399
rect 11739 433 11793 449
rect 11739 413 11749 433
rect 11046 349 11076 383
rect 11240 349 11270 383
rect 11712 399 11749 413
rect 11783 399 11793 433
rect 11712 383 11793 399
rect 11887 433 11941 449
rect 11887 399 11897 433
rect 11931 399 11941 433
rect 11887 383 11941 399
rect 12405 433 12459 449
rect 12405 413 12415 433
rect 11712 349 11742 383
rect 11906 349 11936 383
rect 12378 399 12415 413
rect 12449 399 12459 433
rect 12378 383 12459 399
rect 12553 433 12607 449
rect 12553 399 12563 433
rect 12597 399 12607 433
rect 12553 383 12607 399
rect 12378 349 12408 383
rect 12572 349 12602 383
rect 12997 433 13051 449
rect 12997 399 13007 433
rect 13041 413 13051 433
rect 13219 433 13273 449
rect 13041 399 13074 413
rect 12997 383 13074 399
rect 13219 399 13229 433
rect 13263 399 13273 433
rect 13219 383 13273 399
rect 13737 433 13791 449
rect 13737 413 13747 433
rect 13044 349 13074 383
rect 13238 349 13268 383
rect 13710 399 13747 413
rect 13781 399 13791 433
rect 14033 433 14087 449
rect 14033 413 14043 433
rect 13710 383 13791 399
rect 14010 399 14043 413
rect 14077 399 14087 433
rect 14010 383 14087 399
rect 13710 349 13740 383
rect 14010 349 14040 383
rect 14329 433 14383 449
rect 14329 399 14339 433
rect 14373 413 14383 433
rect 14551 433 14605 449
rect 14373 399 14406 413
rect 14329 383 14406 399
rect 14551 399 14561 433
rect 14595 399 14605 433
rect 14551 383 14605 399
rect 14376 349 14406 383
rect 14570 349 14600 383
<< polycont >>
rect 205 923 239 957
rect 427 923 461 957
rect 649 923 683 957
rect 1167 923 1201 957
rect 1321 923 1355 957
rect 1833 923 1867 957
rect 1987 923 2021 957
rect 2499 923 2533 957
rect 2653 923 2687 957
rect 3165 923 3199 957
rect 3319 923 3353 957
rect 3831 923 3865 957
rect 3985 923 4019 957
rect 4497 923 4531 957
rect 4719 923 4753 957
rect 4941 923 4975 957
rect 5459 923 5493 957
rect 5613 923 5647 957
rect 6125 923 6159 957
rect 6279 923 6313 957
rect 6791 923 6825 957
rect 6945 923 6979 957
rect 7457 923 7491 957
rect 7611 923 7645 957
rect 8123 923 8157 957
rect 8277 923 8311 957
rect 8789 923 8823 957
rect 9011 923 9045 957
rect 9233 923 9267 957
rect 9751 923 9785 957
rect 9905 923 9939 957
rect 10417 923 10451 957
rect 10571 923 10605 957
rect 11083 923 11117 957
rect 11237 923 11271 957
rect 11749 923 11783 957
rect 11903 923 11937 957
rect 12415 923 12449 957
rect 12569 923 12603 957
rect 13007 924 13041 958
rect 13237 924 13271 958
rect 13747 924 13781 958
rect 14043 924 14077 958
rect 14339 924 14373 958
rect 14565 924 14599 958
rect 205 399 239 433
rect 427 399 461 433
rect 649 399 683 433
rect 1167 399 1201 433
rect 1315 399 1349 433
rect 1833 399 1867 433
rect 1981 399 2015 433
rect 2499 399 2533 433
rect 2647 399 2681 433
rect 3165 399 3199 433
rect 3313 399 3347 433
rect 3831 399 3865 433
rect 3979 399 4013 433
rect 4497 399 4531 433
rect 4719 399 4753 433
rect 4941 399 4975 433
rect 5459 399 5493 433
rect 5607 399 5641 433
rect 6125 399 6159 433
rect 6273 399 6307 433
rect 6791 399 6825 433
rect 6939 399 6973 433
rect 7457 399 7491 433
rect 7605 399 7639 433
rect 8123 399 8157 433
rect 8271 399 8305 433
rect 8789 399 8823 433
rect 9011 399 9045 433
rect 9233 399 9267 433
rect 9751 399 9785 433
rect 9899 399 9933 433
rect 10417 399 10451 433
rect 10565 399 10599 433
rect 11083 399 11117 433
rect 11231 399 11265 433
rect 11749 399 11783 433
rect 11897 399 11931 433
rect 12415 399 12449 433
rect 12563 399 12597 433
rect 13007 399 13041 433
rect 13229 399 13263 433
rect 13747 399 13781 433
rect 14043 399 14077 433
rect 14339 399 14373 433
rect 14561 399 14595 433
<< locali >>
rect -34 1497 14908 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5163 1497
rect 5197 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5533 1497
rect 5567 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5755 1497
rect 5789 1463 5829 1497
rect 5863 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6125 1497
rect 6159 1463 6199 1497
rect 6233 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6495 1497
rect 6529 1463 6643 1497
rect 6677 1463 6717 1497
rect 6751 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7087 1497
rect 7121 1463 7161 1497
rect 7195 1463 7309 1497
rect 7343 1463 7383 1497
rect 7417 1463 7457 1497
rect 7491 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7679 1497
rect 7713 1463 7753 1497
rect 7787 1463 7827 1497
rect 7861 1463 7975 1497
rect 8009 1463 8049 1497
rect 8083 1463 8123 1497
rect 8157 1463 8197 1497
rect 8231 1463 8271 1497
rect 8305 1463 8345 1497
rect 8379 1463 8419 1497
rect 8453 1463 8493 1497
rect 8527 1463 8641 1497
rect 8675 1463 8715 1497
rect 8749 1463 8789 1497
rect 8823 1463 8863 1497
rect 8897 1463 8937 1497
rect 8971 1463 9011 1497
rect 9045 1463 9085 1497
rect 9119 1463 9159 1497
rect 9193 1463 9233 1497
rect 9267 1463 9307 1497
rect 9341 1463 9381 1497
rect 9415 1463 9455 1497
rect 9489 1463 9603 1497
rect 9637 1463 9677 1497
rect 9711 1463 9751 1497
rect 9785 1463 9825 1497
rect 9859 1463 9899 1497
rect 9933 1463 9973 1497
rect 10007 1463 10047 1497
rect 10081 1463 10121 1497
rect 10155 1463 10269 1497
rect 10303 1463 10343 1497
rect 10377 1463 10417 1497
rect 10451 1463 10491 1497
rect 10525 1463 10565 1497
rect 10599 1463 10639 1497
rect 10673 1463 10713 1497
rect 10747 1463 10787 1497
rect 10821 1463 10935 1497
rect 10969 1463 11009 1497
rect 11043 1463 11083 1497
rect 11117 1463 11157 1497
rect 11191 1463 11231 1497
rect 11265 1463 11305 1497
rect 11339 1463 11379 1497
rect 11413 1463 11453 1497
rect 11487 1463 11601 1497
rect 11635 1463 11675 1497
rect 11709 1463 11749 1497
rect 11783 1463 11823 1497
rect 11857 1463 11897 1497
rect 11931 1463 11971 1497
rect 12005 1463 12045 1497
rect 12079 1463 12119 1497
rect 12153 1463 12267 1497
rect 12301 1463 12341 1497
rect 12375 1463 12415 1497
rect 12449 1463 12489 1497
rect 12523 1463 12563 1497
rect 12597 1463 12637 1497
rect 12671 1463 12711 1497
rect 12745 1463 12785 1497
rect 12819 1463 12933 1497
rect 12967 1463 13007 1497
rect 13041 1463 13081 1497
rect 13115 1463 13155 1497
rect 13189 1463 13229 1497
rect 13263 1463 13303 1497
rect 13337 1463 13377 1497
rect 13411 1463 13451 1497
rect 13485 1463 13599 1497
rect 13633 1463 13673 1497
rect 13707 1463 13747 1497
rect 13781 1463 13821 1497
rect 13855 1463 13895 1497
rect 13929 1463 13969 1497
rect 14003 1463 14043 1497
rect 14077 1463 14117 1497
rect 14151 1463 14265 1497
rect 14299 1463 14339 1497
rect 14373 1463 14413 1497
rect 14447 1463 14487 1497
rect 14521 1463 14561 1497
rect 14595 1463 14635 1497
rect 14669 1463 14709 1497
rect 14743 1463 14783 1497
rect 14817 1463 14908 1497
rect -34 1446 14908 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 201 1366 235 1446
rect 201 1298 235 1332
rect 201 1230 235 1264
rect 201 1162 235 1196
rect 201 1093 235 1128
rect 201 1043 235 1059
rect 289 1366 323 1404
rect 289 1298 323 1332
rect 289 1230 323 1264
rect 289 1162 323 1196
rect 289 1093 323 1128
rect 377 1366 411 1446
rect 377 1298 411 1332
rect 377 1230 411 1264
rect 377 1162 411 1196
rect 377 1111 411 1128
rect 465 1366 499 1404
rect 465 1298 499 1332
rect 465 1230 499 1264
rect 465 1162 499 1196
rect 289 1048 323 1059
rect 465 1093 499 1128
rect 553 1366 587 1446
rect 553 1298 587 1332
rect 553 1230 587 1264
rect 553 1162 587 1196
rect 553 1111 587 1128
rect 641 1366 675 1404
rect 641 1298 675 1332
rect 641 1230 675 1264
rect 641 1162 675 1196
rect 465 1048 499 1059
rect 641 1093 675 1128
rect 729 1366 763 1446
rect 729 1298 763 1332
rect 729 1230 763 1264
rect 729 1162 763 1196
rect 729 1111 763 1128
rect 928 1423 996 1446
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 641 1048 675 1059
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect -34 979 34 1019
rect 289 1014 831 1048
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect 205 831 239 923
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 797
rect 205 383 239 399
rect 427 957 461 973
rect 427 905 461 923
rect 427 433 461 871
rect 427 383 461 399
rect 649 957 683 973
rect 649 683 683 923
rect 649 433 683 649
rect 649 383 683 399
rect 797 757 831 1014
rect 928 1019 945 1053
rect 979 1019 996 1053
rect 1103 1366 1137 1446
rect 1103 1298 1137 1332
rect 1103 1230 1137 1264
rect 1103 1162 1137 1196
rect 1103 1093 1137 1128
rect 1103 1027 1137 1059
rect 1191 1366 1225 1404
rect 1191 1298 1225 1332
rect 1191 1230 1225 1264
rect 1191 1162 1225 1196
rect 1191 1093 1225 1128
rect 1279 1366 1313 1446
rect 1279 1298 1313 1332
rect 1279 1230 1313 1264
rect 1279 1162 1313 1196
rect 1279 1111 1313 1128
rect 1367 1366 1401 1404
rect 1367 1298 1401 1332
rect 1367 1230 1401 1264
rect 1367 1162 1401 1196
rect 1191 1057 1225 1059
rect 1367 1093 1401 1128
rect 1455 1366 1489 1446
rect 1455 1298 1489 1332
rect 1455 1230 1489 1264
rect 1455 1162 1489 1196
rect 1455 1111 1489 1128
rect 1594 1423 1662 1446
rect 1594 1389 1611 1423
rect 1645 1389 1662 1423
rect 1594 1349 1662 1389
rect 1594 1315 1611 1349
rect 1645 1315 1662 1349
rect 1594 1275 1662 1315
rect 1594 1241 1611 1275
rect 1645 1241 1662 1275
rect 1594 1201 1662 1241
rect 1594 1167 1611 1201
rect 1645 1167 1662 1201
rect 1594 1127 1662 1167
rect 1367 1057 1401 1059
rect 1594 1093 1611 1127
rect 1645 1093 1662 1127
rect 1191 1023 1497 1057
rect 928 979 996 1019
rect 928 945 945 979
rect 979 945 996 979
rect 928 905 996 945
rect 928 871 945 905
rect 979 871 996 905
rect 928 822 996 871
rect 1167 957 1201 973
rect 1321 957 1355 973
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 101 335 135 351
rect 295 335 329 351
rect 489 335 523 351
rect 135 301 198 335
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 489 335
rect 101 263 135 301
rect 101 195 135 229
rect 295 263 329 301
rect 489 285 523 301
rect 603 335 637 351
rect 797 350 831 723
rect 1167 757 1201 923
rect 603 263 637 301
rect 101 125 135 161
rect 101 75 135 91
rect 198 210 232 226
rect -34 34 34 57
rect 198 34 232 176
rect 295 195 329 229
rect 393 216 427 232
rect 603 216 637 229
rect 427 195 637 216
rect 427 182 603 195
rect 393 166 427 182
rect 295 125 329 161
rect 700 316 831 350
rect 928 461 996 544
rect 928 427 945 461
rect 979 427 996 461
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect 1167 433 1201 723
rect 1167 383 1201 399
rect 1315 923 1321 942
rect 1315 907 1355 923
rect 1315 535 1349 907
rect 1315 433 1349 501
rect 1315 383 1349 399
rect 1463 683 1497 1023
rect 1594 1053 1662 1093
rect 1594 1019 1611 1053
rect 1645 1019 1662 1053
rect 1769 1366 1803 1446
rect 1769 1298 1803 1332
rect 1769 1230 1803 1264
rect 1769 1162 1803 1196
rect 1769 1093 1803 1128
rect 1769 1027 1803 1059
rect 1857 1366 1891 1404
rect 1857 1298 1891 1332
rect 1857 1230 1891 1264
rect 1857 1162 1891 1196
rect 1857 1093 1891 1128
rect 1945 1366 1979 1446
rect 1945 1298 1979 1332
rect 1945 1230 1979 1264
rect 1945 1162 1979 1196
rect 1945 1111 1979 1128
rect 2033 1366 2067 1404
rect 2033 1298 2067 1332
rect 2033 1230 2067 1264
rect 2033 1162 2067 1196
rect 1857 1057 1891 1059
rect 2033 1093 2067 1128
rect 2121 1366 2155 1446
rect 2121 1298 2155 1332
rect 2121 1230 2155 1264
rect 2121 1162 2155 1196
rect 2121 1111 2155 1128
rect 2260 1423 2328 1446
rect 2260 1389 2277 1423
rect 2311 1389 2328 1423
rect 2260 1349 2328 1389
rect 2260 1315 2277 1349
rect 2311 1315 2328 1349
rect 2260 1275 2328 1315
rect 2260 1241 2277 1275
rect 2311 1241 2328 1275
rect 2260 1201 2328 1241
rect 2260 1167 2277 1201
rect 2311 1167 2328 1201
rect 2260 1127 2328 1167
rect 2033 1057 2067 1059
rect 2260 1093 2277 1127
rect 2311 1093 2328 1127
rect 1857 1023 2163 1057
rect 1594 979 1662 1019
rect 1594 945 1611 979
rect 1645 945 1662 979
rect 1594 905 1662 945
rect 1594 871 1611 905
rect 1645 871 1662 905
rect 1594 822 1662 871
rect 1833 957 1867 973
rect 1987 957 2021 973
rect 700 219 734 316
rect 928 313 996 353
rect 928 279 945 313
rect 979 279 996 313
rect 700 169 734 185
rect 797 263 831 279
rect 797 195 831 229
rect 489 125 523 141
rect 329 91 392 125
rect 426 91 489 125
rect 295 75 329 91
rect 489 75 523 91
rect 603 125 637 161
rect 797 125 831 161
rect 637 91 700 125
rect 734 91 797 125
rect 603 75 637 91
rect 797 75 831 91
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect 928 57 945 91
rect 979 57 996 91
rect 1084 333 1118 349
rect 1278 333 1312 349
rect 1463 348 1497 649
rect 1833 683 1867 923
rect 1118 299 1181 333
rect 1215 299 1278 333
rect 1084 261 1118 299
rect 1084 193 1118 227
rect 1278 261 1312 299
rect 1084 123 1118 159
rect 1084 73 1118 89
rect 1181 208 1215 224
rect 928 34 996 57
rect 1181 34 1215 174
rect 1278 193 1312 227
rect 1375 314 1497 348
rect 1594 461 1662 544
rect 1594 427 1611 461
rect 1645 427 1662 461
rect 1594 387 1662 427
rect 1594 353 1611 387
rect 1645 353 1662 387
rect 1833 433 1867 649
rect 1833 383 1867 399
rect 1981 923 1987 942
rect 1981 907 2021 923
rect 1981 831 2015 907
rect 1981 433 2015 797
rect 1981 383 2015 399
rect 2129 683 2163 1023
rect 2260 1053 2328 1093
rect 2260 1019 2277 1053
rect 2311 1019 2328 1053
rect 2435 1366 2469 1446
rect 2435 1298 2469 1332
rect 2435 1230 2469 1264
rect 2435 1162 2469 1196
rect 2435 1093 2469 1128
rect 2435 1027 2469 1059
rect 2523 1366 2557 1404
rect 2523 1298 2557 1332
rect 2523 1230 2557 1264
rect 2523 1162 2557 1196
rect 2523 1093 2557 1128
rect 2611 1366 2645 1446
rect 2611 1298 2645 1332
rect 2611 1230 2645 1264
rect 2611 1162 2645 1196
rect 2611 1111 2645 1128
rect 2699 1366 2733 1404
rect 2699 1298 2733 1332
rect 2699 1230 2733 1264
rect 2699 1162 2733 1196
rect 2523 1057 2557 1059
rect 2699 1093 2733 1128
rect 2787 1366 2821 1446
rect 2787 1298 2821 1332
rect 2787 1230 2821 1264
rect 2787 1162 2821 1196
rect 2787 1111 2821 1128
rect 2926 1423 2994 1446
rect 2926 1389 2943 1423
rect 2977 1389 2994 1423
rect 2926 1349 2994 1389
rect 2926 1315 2943 1349
rect 2977 1315 2994 1349
rect 2926 1275 2994 1315
rect 2926 1241 2943 1275
rect 2977 1241 2994 1275
rect 2926 1201 2994 1241
rect 2926 1167 2943 1201
rect 2977 1167 2994 1201
rect 2926 1127 2994 1167
rect 2699 1057 2733 1059
rect 2926 1093 2943 1127
rect 2977 1093 2994 1127
rect 2523 1023 2829 1057
rect 2260 979 2328 1019
rect 2260 945 2277 979
rect 2311 945 2328 979
rect 2260 905 2328 945
rect 2260 871 2277 905
rect 2311 871 2328 905
rect 2260 822 2328 871
rect 2499 957 2533 973
rect 2653 957 2687 973
rect 1375 217 1409 314
rect 1594 313 1662 353
rect 1594 279 1611 313
rect 1645 279 1662 313
rect 1375 167 1409 183
rect 1472 261 1506 277
rect 1472 193 1506 227
rect 1278 123 1312 159
rect 1472 123 1506 159
rect 1312 89 1375 123
rect 1409 89 1472 123
rect 1278 73 1312 89
rect 1472 73 1506 89
rect 1594 239 1662 279
rect 1594 205 1611 239
rect 1645 205 1662 239
rect 1594 165 1662 205
rect 1594 131 1611 165
rect 1645 131 1662 165
rect 1594 91 1662 131
rect 1594 57 1611 91
rect 1645 57 1662 91
rect 1750 333 1784 349
rect 1944 333 1978 349
rect 2129 348 2163 649
rect 2499 683 2533 923
rect 1784 299 1847 333
rect 1881 299 1944 333
rect 1750 261 1784 299
rect 1750 193 1784 227
rect 1944 261 1978 299
rect 1750 123 1784 159
rect 1750 73 1784 89
rect 1847 208 1881 224
rect 1594 34 1662 57
rect 1847 34 1881 174
rect 1944 193 1978 227
rect 2041 314 2163 348
rect 2260 461 2328 544
rect 2260 427 2277 461
rect 2311 427 2328 461
rect 2260 387 2328 427
rect 2260 353 2277 387
rect 2311 353 2328 387
rect 2499 433 2533 649
rect 2499 383 2533 399
rect 2647 923 2653 942
rect 2647 907 2687 923
rect 2647 905 2681 907
rect 2647 433 2681 871
rect 2647 383 2681 399
rect 2795 831 2829 1023
rect 2926 1053 2994 1093
rect 2926 1019 2943 1053
rect 2977 1019 2994 1053
rect 3101 1366 3135 1446
rect 3101 1298 3135 1332
rect 3101 1230 3135 1264
rect 3101 1162 3135 1196
rect 3101 1093 3135 1128
rect 3101 1027 3135 1059
rect 3189 1366 3223 1404
rect 3189 1298 3223 1332
rect 3189 1230 3223 1264
rect 3189 1162 3223 1196
rect 3189 1093 3223 1128
rect 3277 1366 3311 1446
rect 3277 1298 3311 1332
rect 3277 1230 3311 1264
rect 3277 1162 3311 1196
rect 3277 1111 3311 1128
rect 3365 1366 3399 1404
rect 3365 1298 3399 1332
rect 3365 1230 3399 1264
rect 3365 1162 3399 1196
rect 3189 1057 3223 1059
rect 3365 1093 3399 1128
rect 3453 1366 3487 1446
rect 3453 1298 3487 1332
rect 3453 1230 3487 1264
rect 3453 1162 3487 1196
rect 3453 1111 3487 1128
rect 3592 1423 3660 1446
rect 3592 1389 3609 1423
rect 3643 1389 3660 1423
rect 3592 1349 3660 1389
rect 3592 1315 3609 1349
rect 3643 1315 3660 1349
rect 3592 1275 3660 1315
rect 3592 1241 3609 1275
rect 3643 1241 3660 1275
rect 3592 1201 3660 1241
rect 3592 1167 3609 1201
rect 3643 1167 3660 1201
rect 3592 1127 3660 1167
rect 3365 1057 3399 1059
rect 3592 1093 3609 1127
rect 3643 1093 3660 1127
rect 3189 1023 3495 1057
rect 2926 979 2994 1019
rect 2926 945 2943 979
rect 2977 945 2994 979
rect 2926 905 2994 945
rect 2926 871 2943 905
rect 2977 871 2994 905
rect 2926 822 2994 871
rect 3165 957 3199 973
rect 3319 957 3353 973
rect 2041 217 2075 314
rect 2260 313 2328 353
rect 2260 279 2277 313
rect 2311 279 2328 313
rect 2041 167 2075 183
rect 2138 261 2172 277
rect 2138 193 2172 227
rect 1944 123 1978 159
rect 2138 123 2172 159
rect 1978 89 2041 123
rect 2075 89 2138 123
rect 1944 73 1978 89
rect 2138 73 2172 89
rect 2260 239 2328 279
rect 2260 205 2277 239
rect 2311 205 2328 239
rect 2260 165 2328 205
rect 2260 131 2277 165
rect 2311 131 2328 165
rect 2260 91 2328 131
rect 2260 57 2277 91
rect 2311 57 2328 91
rect 2416 333 2450 349
rect 2610 333 2644 349
rect 2795 348 2829 797
rect 3165 757 3199 923
rect 2450 299 2513 333
rect 2547 299 2610 333
rect 2416 261 2450 299
rect 2416 193 2450 227
rect 2610 261 2644 299
rect 2416 123 2450 159
rect 2416 73 2450 89
rect 2513 208 2547 224
rect 2260 34 2328 57
rect 2513 34 2547 174
rect 2610 193 2644 227
rect 2707 314 2829 348
rect 2926 461 2994 544
rect 2926 427 2943 461
rect 2977 427 2994 461
rect 2926 387 2994 427
rect 2926 353 2943 387
rect 2977 353 2994 387
rect 3165 433 3199 723
rect 3165 383 3199 399
rect 3313 923 3319 942
rect 3313 907 3353 923
rect 3313 609 3347 907
rect 3313 433 3347 575
rect 3313 383 3347 399
rect 3461 757 3495 1023
rect 3592 1053 3660 1093
rect 3592 1019 3609 1053
rect 3643 1019 3660 1053
rect 3767 1366 3801 1446
rect 3767 1298 3801 1332
rect 3767 1230 3801 1264
rect 3767 1162 3801 1196
rect 3767 1093 3801 1128
rect 3767 1027 3801 1059
rect 3855 1366 3889 1404
rect 3855 1298 3889 1332
rect 3855 1230 3889 1264
rect 3855 1162 3889 1196
rect 3855 1093 3889 1128
rect 3943 1366 3977 1446
rect 3943 1298 3977 1332
rect 3943 1230 3977 1264
rect 3943 1162 3977 1196
rect 3943 1111 3977 1128
rect 4031 1366 4065 1404
rect 4031 1298 4065 1332
rect 4031 1230 4065 1264
rect 4031 1162 4065 1196
rect 3855 1057 3889 1059
rect 4031 1093 4065 1128
rect 4119 1366 4153 1446
rect 4119 1298 4153 1332
rect 4119 1230 4153 1264
rect 4119 1162 4153 1196
rect 4119 1111 4153 1128
rect 4258 1423 4326 1446
rect 4258 1389 4275 1423
rect 4309 1389 4326 1423
rect 4258 1349 4326 1389
rect 4258 1315 4275 1349
rect 4309 1315 4326 1349
rect 4258 1275 4326 1315
rect 4258 1241 4275 1275
rect 4309 1241 4326 1275
rect 4258 1201 4326 1241
rect 4258 1167 4275 1201
rect 4309 1167 4326 1201
rect 4258 1127 4326 1167
rect 4031 1057 4065 1059
rect 4258 1093 4275 1127
rect 4309 1093 4326 1127
rect 3855 1023 4161 1057
rect 3592 979 3660 1019
rect 3592 945 3609 979
rect 3643 945 3660 979
rect 3592 905 3660 945
rect 3592 871 3609 905
rect 3643 871 3660 905
rect 3592 822 3660 871
rect 3831 957 3865 973
rect 3985 957 4019 973
rect 2707 217 2741 314
rect 2926 313 2994 353
rect 2926 279 2943 313
rect 2977 279 2994 313
rect 2707 167 2741 183
rect 2804 261 2838 277
rect 2804 193 2838 227
rect 2610 123 2644 159
rect 2804 123 2838 159
rect 2644 89 2707 123
rect 2741 89 2804 123
rect 2610 73 2644 89
rect 2804 73 2838 89
rect 2926 239 2994 279
rect 2926 205 2943 239
rect 2977 205 2994 239
rect 2926 165 2994 205
rect 2926 131 2943 165
rect 2977 131 2994 165
rect 2926 91 2994 131
rect 2926 57 2943 91
rect 2977 57 2994 91
rect 3082 333 3116 349
rect 3276 333 3310 349
rect 3461 348 3495 723
rect 3831 757 3865 923
rect 3116 299 3179 333
rect 3213 299 3276 333
rect 3082 261 3116 299
rect 3082 193 3116 227
rect 3276 261 3310 299
rect 3082 123 3116 159
rect 3082 73 3116 89
rect 3179 208 3213 224
rect 2926 34 2994 57
rect 3179 34 3213 174
rect 3276 193 3310 227
rect 3373 314 3495 348
rect 3592 461 3660 544
rect 3592 427 3609 461
rect 3643 427 3660 461
rect 3592 387 3660 427
rect 3592 353 3609 387
rect 3643 353 3660 387
rect 3831 433 3865 723
rect 3831 383 3865 399
rect 3979 923 3985 942
rect 3979 907 4019 923
rect 3979 831 4013 907
rect 3979 433 4013 797
rect 3979 383 4013 399
rect 4127 609 4161 1023
rect 4258 1053 4326 1093
rect 4258 1019 4275 1053
rect 4309 1019 4326 1053
rect 4493 1366 4527 1446
rect 4493 1298 4527 1332
rect 4493 1230 4527 1264
rect 4493 1162 4527 1196
rect 4493 1093 4527 1128
rect 4493 1043 4527 1059
rect 4581 1366 4615 1404
rect 4581 1298 4615 1332
rect 4581 1230 4615 1264
rect 4581 1162 4615 1196
rect 4581 1093 4615 1128
rect 4669 1366 4703 1446
rect 4669 1298 4703 1332
rect 4669 1230 4703 1264
rect 4669 1162 4703 1196
rect 4669 1111 4703 1128
rect 4757 1366 4791 1404
rect 4757 1298 4791 1332
rect 4757 1230 4791 1264
rect 4757 1162 4791 1196
rect 4581 1048 4615 1059
rect 4757 1093 4791 1128
rect 4845 1366 4879 1446
rect 4845 1298 4879 1332
rect 4845 1230 4879 1264
rect 4845 1162 4879 1196
rect 4845 1111 4879 1128
rect 4933 1366 4967 1404
rect 4933 1298 4967 1332
rect 4933 1230 4967 1264
rect 4933 1162 4967 1196
rect 4757 1048 4791 1059
rect 4933 1093 4967 1128
rect 5021 1366 5055 1446
rect 5021 1298 5055 1332
rect 5021 1230 5055 1264
rect 5021 1162 5055 1196
rect 5021 1111 5055 1128
rect 5220 1423 5288 1446
rect 5220 1389 5237 1423
rect 5271 1389 5288 1423
rect 5220 1349 5288 1389
rect 5220 1315 5237 1349
rect 5271 1315 5288 1349
rect 5220 1275 5288 1315
rect 5220 1241 5237 1275
rect 5271 1241 5288 1275
rect 5220 1201 5288 1241
rect 5220 1167 5237 1201
rect 5271 1167 5288 1201
rect 5220 1127 5288 1167
rect 4933 1048 4967 1059
rect 5220 1093 5237 1127
rect 5271 1093 5288 1127
rect 5220 1053 5288 1093
rect 4258 979 4326 1019
rect 4581 1014 5123 1048
rect 4258 945 4275 979
rect 4309 945 4326 979
rect 4258 905 4326 945
rect 4258 871 4275 905
rect 4309 871 4326 905
rect 4258 822 4326 871
rect 4497 957 4531 973
rect 4497 831 4531 923
rect 3373 217 3407 314
rect 3592 313 3660 353
rect 3592 279 3609 313
rect 3643 279 3660 313
rect 3373 167 3407 183
rect 3470 261 3504 277
rect 3470 193 3504 227
rect 3276 123 3310 159
rect 3470 123 3504 159
rect 3310 89 3373 123
rect 3407 89 3470 123
rect 3276 73 3310 89
rect 3470 73 3504 89
rect 3592 239 3660 279
rect 3592 205 3609 239
rect 3643 205 3660 239
rect 3592 165 3660 205
rect 3592 131 3609 165
rect 3643 131 3660 165
rect 3592 91 3660 131
rect 3592 57 3609 91
rect 3643 57 3660 91
rect 3748 333 3782 349
rect 3942 333 3976 349
rect 4127 348 4161 575
rect 3782 299 3845 333
rect 3879 299 3942 333
rect 3748 261 3782 299
rect 3748 193 3782 227
rect 3942 261 3976 299
rect 3748 123 3782 159
rect 3748 73 3782 89
rect 3845 208 3879 224
rect 3592 34 3660 57
rect 3845 34 3879 174
rect 3942 193 3976 227
rect 4039 314 4161 348
rect 4258 461 4326 544
rect 4258 427 4275 461
rect 4309 427 4326 461
rect 4258 387 4326 427
rect 4258 353 4275 387
rect 4309 353 4326 387
rect 4497 433 4531 797
rect 4497 383 4531 399
rect 4719 957 4753 973
rect 4719 905 4753 923
rect 4719 433 4753 871
rect 4719 383 4753 399
rect 4941 957 4975 973
rect 4941 683 4975 923
rect 4941 433 4975 649
rect 4941 383 4975 399
rect 5089 757 5123 1014
rect 5220 1019 5237 1053
rect 5271 1019 5288 1053
rect 5395 1366 5429 1446
rect 5395 1298 5429 1332
rect 5395 1230 5429 1264
rect 5395 1162 5429 1196
rect 5395 1093 5429 1128
rect 5395 1027 5429 1059
rect 5483 1366 5517 1404
rect 5483 1298 5517 1332
rect 5483 1230 5517 1264
rect 5483 1162 5517 1196
rect 5483 1093 5517 1128
rect 5571 1366 5605 1446
rect 5571 1298 5605 1332
rect 5571 1230 5605 1264
rect 5571 1162 5605 1196
rect 5571 1111 5605 1128
rect 5659 1366 5693 1404
rect 5659 1298 5693 1332
rect 5659 1230 5693 1264
rect 5659 1162 5693 1196
rect 5483 1057 5517 1059
rect 5659 1093 5693 1128
rect 5747 1366 5781 1446
rect 5747 1298 5781 1332
rect 5747 1230 5781 1264
rect 5747 1162 5781 1196
rect 5747 1111 5781 1128
rect 5886 1423 5954 1446
rect 5886 1389 5903 1423
rect 5937 1389 5954 1423
rect 5886 1349 5954 1389
rect 5886 1315 5903 1349
rect 5937 1315 5954 1349
rect 5886 1275 5954 1315
rect 5886 1241 5903 1275
rect 5937 1241 5954 1275
rect 5886 1201 5954 1241
rect 5886 1167 5903 1201
rect 5937 1167 5954 1201
rect 5886 1127 5954 1167
rect 5659 1057 5693 1059
rect 5886 1093 5903 1127
rect 5937 1093 5954 1127
rect 5483 1023 5789 1057
rect 5220 979 5288 1019
rect 5220 945 5237 979
rect 5271 945 5288 979
rect 5220 905 5288 945
rect 5220 871 5237 905
rect 5271 871 5288 905
rect 5220 822 5288 871
rect 5459 957 5493 973
rect 5613 957 5647 973
rect 4039 217 4073 314
rect 4258 313 4326 353
rect 4258 279 4275 313
rect 4309 279 4326 313
rect 4039 167 4073 183
rect 4136 261 4170 277
rect 4136 193 4170 227
rect 3942 123 3976 159
rect 4136 123 4170 159
rect 3976 89 4039 123
rect 4073 89 4136 123
rect 3942 73 3976 89
rect 4136 73 4170 89
rect 4258 239 4326 279
rect 4258 205 4275 239
rect 4309 205 4326 239
rect 4258 165 4326 205
rect 4258 131 4275 165
rect 4309 131 4326 165
rect 4258 91 4326 131
rect 4258 57 4275 91
rect 4309 57 4326 91
rect 4393 335 4427 351
rect 4587 335 4621 351
rect 4781 335 4815 351
rect 4427 301 4490 335
rect 4524 301 4587 335
rect 4621 301 4684 335
rect 4718 301 4781 335
rect 4393 263 4427 301
rect 4393 195 4427 229
rect 4587 263 4621 301
rect 4781 285 4815 301
rect 4895 335 4929 351
rect 5089 350 5123 723
rect 5459 757 5493 923
rect 4895 263 4929 301
rect 4393 125 4427 161
rect 4393 75 4427 91
rect 4490 210 4524 226
rect 4258 34 4326 57
rect 4490 34 4524 176
rect 4587 195 4621 229
rect 4685 216 4719 232
rect 4895 216 4929 229
rect 4719 195 4929 216
rect 4719 182 4895 195
rect 4685 166 4719 182
rect 4587 125 4621 161
rect 4992 316 5123 350
rect 5220 461 5288 544
rect 5220 427 5237 461
rect 5271 427 5288 461
rect 5220 387 5288 427
rect 5220 353 5237 387
rect 5271 353 5288 387
rect 5459 433 5493 723
rect 5459 383 5493 399
rect 5607 923 5613 942
rect 5607 907 5647 923
rect 5607 535 5641 907
rect 5607 433 5641 501
rect 5607 383 5641 399
rect 5755 683 5789 1023
rect 5886 1053 5954 1093
rect 5886 1019 5903 1053
rect 5937 1019 5954 1053
rect 6061 1366 6095 1446
rect 6061 1298 6095 1332
rect 6061 1230 6095 1264
rect 6061 1162 6095 1196
rect 6061 1093 6095 1128
rect 6061 1027 6095 1059
rect 6149 1366 6183 1404
rect 6149 1298 6183 1332
rect 6149 1230 6183 1264
rect 6149 1162 6183 1196
rect 6149 1093 6183 1128
rect 6237 1366 6271 1446
rect 6237 1298 6271 1332
rect 6237 1230 6271 1264
rect 6237 1162 6271 1196
rect 6237 1111 6271 1128
rect 6325 1366 6359 1404
rect 6325 1298 6359 1332
rect 6325 1230 6359 1264
rect 6325 1162 6359 1196
rect 6149 1057 6183 1059
rect 6325 1093 6359 1128
rect 6413 1366 6447 1446
rect 6413 1298 6447 1332
rect 6413 1230 6447 1264
rect 6413 1162 6447 1196
rect 6413 1111 6447 1128
rect 6552 1423 6620 1446
rect 6552 1389 6569 1423
rect 6603 1389 6620 1423
rect 6552 1349 6620 1389
rect 6552 1315 6569 1349
rect 6603 1315 6620 1349
rect 6552 1275 6620 1315
rect 6552 1241 6569 1275
rect 6603 1241 6620 1275
rect 6552 1201 6620 1241
rect 6552 1167 6569 1201
rect 6603 1167 6620 1201
rect 6552 1127 6620 1167
rect 6325 1057 6359 1059
rect 6552 1093 6569 1127
rect 6603 1093 6620 1127
rect 6149 1023 6455 1057
rect 5886 979 5954 1019
rect 5886 945 5903 979
rect 5937 945 5954 979
rect 5886 905 5954 945
rect 5886 871 5903 905
rect 5937 871 5954 905
rect 5886 822 5954 871
rect 6125 957 6159 973
rect 6279 957 6313 973
rect 4992 219 5026 316
rect 5220 313 5288 353
rect 5220 279 5237 313
rect 5271 279 5288 313
rect 4992 169 5026 185
rect 5089 263 5123 279
rect 5089 195 5123 229
rect 4781 125 4815 141
rect 4621 91 4684 125
rect 4718 91 4781 125
rect 4587 75 4621 91
rect 4781 75 4815 91
rect 4895 125 4929 161
rect 5089 125 5123 161
rect 4929 91 4992 125
rect 5026 91 5089 125
rect 4895 75 4929 91
rect 5089 75 5123 91
rect 5220 239 5288 279
rect 5220 205 5237 239
rect 5271 205 5288 239
rect 5220 165 5288 205
rect 5220 131 5237 165
rect 5271 131 5288 165
rect 5220 91 5288 131
rect 5220 57 5237 91
rect 5271 57 5288 91
rect 5376 333 5410 349
rect 5570 333 5604 349
rect 5755 348 5789 649
rect 6125 683 6159 923
rect 5410 299 5473 333
rect 5507 299 5570 333
rect 5376 261 5410 299
rect 5376 193 5410 227
rect 5570 261 5604 299
rect 5376 123 5410 159
rect 5376 73 5410 89
rect 5473 208 5507 224
rect 5220 34 5288 57
rect 5473 34 5507 174
rect 5570 193 5604 227
rect 5667 314 5789 348
rect 5886 461 5954 544
rect 5886 427 5903 461
rect 5937 427 5954 461
rect 5886 387 5954 427
rect 5886 353 5903 387
rect 5937 353 5954 387
rect 6125 433 6159 649
rect 6125 383 6159 399
rect 6273 923 6279 942
rect 6273 907 6313 923
rect 6273 831 6307 907
rect 6273 433 6307 797
rect 6273 383 6307 399
rect 6421 683 6455 1023
rect 6552 1053 6620 1093
rect 6552 1019 6569 1053
rect 6603 1019 6620 1053
rect 6727 1366 6761 1446
rect 6727 1298 6761 1332
rect 6727 1230 6761 1264
rect 6727 1162 6761 1196
rect 6727 1093 6761 1128
rect 6727 1027 6761 1059
rect 6815 1366 6849 1404
rect 6815 1298 6849 1332
rect 6815 1230 6849 1264
rect 6815 1162 6849 1196
rect 6815 1093 6849 1128
rect 6903 1366 6937 1446
rect 6903 1298 6937 1332
rect 6903 1230 6937 1264
rect 6903 1162 6937 1196
rect 6903 1111 6937 1128
rect 6991 1366 7025 1404
rect 6991 1298 7025 1332
rect 6991 1230 7025 1264
rect 6991 1162 7025 1196
rect 6815 1057 6849 1059
rect 6991 1093 7025 1128
rect 7079 1366 7113 1446
rect 7079 1298 7113 1332
rect 7079 1230 7113 1264
rect 7079 1162 7113 1196
rect 7079 1111 7113 1128
rect 7218 1423 7286 1446
rect 7218 1389 7235 1423
rect 7269 1389 7286 1423
rect 7218 1349 7286 1389
rect 7218 1315 7235 1349
rect 7269 1315 7286 1349
rect 7218 1275 7286 1315
rect 7218 1241 7235 1275
rect 7269 1241 7286 1275
rect 7218 1201 7286 1241
rect 7218 1167 7235 1201
rect 7269 1167 7286 1201
rect 7218 1127 7286 1167
rect 6991 1057 7025 1059
rect 7218 1093 7235 1127
rect 7269 1093 7286 1127
rect 6815 1023 7121 1057
rect 6552 979 6620 1019
rect 6552 945 6569 979
rect 6603 945 6620 979
rect 6552 905 6620 945
rect 6552 871 6569 905
rect 6603 871 6620 905
rect 6552 822 6620 871
rect 6791 957 6825 973
rect 6945 957 6979 973
rect 5667 217 5701 314
rect 5886 313 5954 353
rect 5886 279 5903 313
rect 5937 279 5954 313
rect 5667 167 5701 183
rect 5764 261 5798 277
rect 5764 193 5798 227
rect 5570 123 5604 159
rect 5764 123 5798 159
rect 5604 89 5667 123
rect 5701 89 5764 123
rect 5570 73 5604 89
rect 5764 73 5798 89
rect 5886 239 5954 279
rect 5886 205 5903 239
rect 5937 205 5954 239
rect 5886 165 5954 205
rect 5886 131 5903 165
rect 5937 131 5954 165
rect 5886 91 5954 131
rect 5886 57 5903 91
rect 5937 57 5954 91
rect 6042 333 6076 349
rect 6236 333 6270 349
rect 6421 348 6455 649
rect 6791 683 6825 923
rect 6076 299 6139 333
rect 6173 299 6236 333
rect 6042 261 6076 299
rect 6042 193 6076 227
rect 6236 261 6270 299
rect 6042 123 6076 159
rect 6042 73 6076 89
rect 6139 208 6173 224
rect 5886 34 5954 57
rect 6139 34 6173 174
rect 6236 193 6270 227
rect 6333 314 6455 348
rect 6552 461 6620 544
rect 6552 427 6569 461
rect 6603 427 6620 461
rect 6552 387 6620 427
rect 6552 353 6569 387
rect 6603 353 6620 387
rect 6791 433 6825 649
rect 6791 383 6825 399
rect 6939 923 6945 942
rect 6939 907 6979 923
rect 6939 905 6973 907
rect 6939 433 6973 871
rect 6939 383 6973 399
rect 7087 831 7121 1023
rect 7218 1053 7286 1093
rect 7218 1019 7235 1053
rect 7269 1019 7286 1053
rect 7393 1366 7427 1446
rect 7393 1298 7427 1332
rect 7393 1230 7427 1264
rect 7393 1162 7427 1196
rect 7393 1093 7427 1128
rect 7393 1027 7427 1059
rect 7481 1366 7515 1404
rect 7481 1298 7515 1332
rect 7481 1230 7515 1264
rect 7481 1162 7515 1196
rect 7481 1093 7515 1128
rect 7569 1366 7603 1446
rect 7569 1298 7603 1332
rect 7569 1230 7603 1264
rect 7569 1162 7603 1196
rect 7569 1111 7603 1128
rect 7657 1366 7691 1404
rect 7657 1298 7691 1332
rect 7657 1230 7691 1264
rect 7657 1162 7691 1196
rect 7481 1057 7515 1059
rect 7657 1093 7691 1128
rect 7745 1366 7779 1446
rect 7745 1298 7779 1332
rect 7745 1230 7779 1264
rect 7745 1162 7779 1196
rect 7745 1111 7779 1128
rect 7884 1423 7952 1446
rect 7884 1389 7901 1423
rect 7935 1389 7952 1423
rect 7884 1349 7952 1389
rect 7884 1315 7901 1349
rect 7935 1315 7952 1349
rect 7884 1275 7952 1315
rect 7884 1241 7901 1275
rect 7935 1241 7952 1275
rect 7884 1201 7952 1241
rect 7884 1167 7901 1201
rect 7935 1167 7952 1201
rect 7884 1127 7952 1167
rect 7657 1057 7691 1059
rect 7884 1093 7901 1127
rect 7935 1093 7952 1127
rect 7481 1023 7787 1057
rect 7218 979 7286 1019
rect 7218 945 7235 979
rect 7269 945 7286 979
rect 7218 905 7286 945
rect 7218 871 7235 905
rect 7269 871 7286 905
rect 7218 822 7286 871
rect 7457 957 7491 973
rect 7611 957 7645 973
rect 6333 217 6367 314
rect 6552 313 6620 353
rect 6552 279 6569 313
rect 6603 279 6620 313
rect 6333 167 6367 183
rect 6430 261 6464 277
rect 6430 193 6464 227
rect 6236 123 6270 159
rect 6430 123 6464 159
rect 6270 89 6333 123
rect 6367 89 6430 123
rect 6236 73 6270 89
rect 6430 73 6464 89
rect 6552 239 6620 279
rect 6552 205 6569 239
rect 6603 205 6620 239
rect 6552 165 6620 205
rect 6552 131 6569 165
rect 6603 131 6620 165
rect 6552 91 6620 131
rect 6552 57 6569 91
rect 6603 57 6620 91
rect 6708 333 6742 349
rect 6902 333 6936 349
rect 7087 348 7121 797
rect 7457 757 7491 923
rect 6742 299 6805 333
rect 6839 299 6902 333
rect 6708 261 6742 299
rect 6708 193 6742 227
rect 6902 261 6936 299
rect 6708 123 6742 159
rect 6708 73 6742 89
rect 6805 208 6839 224
rect 6552 34 6620 57
rect 6805 34 6839 174
rect 6902 193 6936 227
rect 6999 314 7121 348
rect 7218 461 7286 544
rect 7218 427 7235 461
rect 7269 427 7286 461
rect 7218 387 7286 427
rect 7218 353 7235 387
rect 7269 353 7286 387
rect 7457 433 7491 723
rect 7457 383 7491 399
rect 7605 923 7611 942
rect 7605 907 7645 923
rect 7605 461 7639 907
rect 7605 383 7639 399
rect 7753 757 7787 1023
rect 7884 1053 7952 1093
rect 7884 1019 7901 1053
rect 7935 1019 7952 1053
rect 8059 1366 8093 1446
rect 8059 1298 8093 1332
rect 8059 1230 8093 1264
rect 8059 1162 8093 1196
rect 8059 1093 8093 1128
rect 8059 1027 8093 1059
rect 8147 1366 8181 1404
rect 8147 1298 8181 1332
rect 8147 1230 8181 1264
rect 8147 1162 8181 1196
rect 8147 1093 8181 1128
rect 8235 1366 8269 1446
rect 8235 1298 8269 1332
rect 8235 1230 8269 1264
rect 8235 1162 8269 1196
rect 8235 1111 8269 1128
rect 8323 1366 8357 1404
rect 8323 1298 8357 1332
rect 8323 1230 8357 1264
rect 8323 1162 8357 1196
rect 8147 1057 8181 1059
rect 8323 1093 8357 1128
rect 8411 1366 8445 1446
rect 8411 1298 8445 1332
rect 8411 1230 8445 1264
rect 8411 1162 8445 1196
rect 8411 1111 8445 1128
rect 8550 1423 8618 1446
rect 8550 1389 8567 1423
rect 8601 1389 8618 1423
rect 8550 1349 8618 1389
rect 8550 1315 8567 1349
rect 8601 1315 8618 1349
rect 8550 1275 8618 1315
rect 8550 1241 8567 1275
rect 8601 1241 8618 1275
rect 8550 1201 8618 1241
rect 8550 1167 8567 1201
rect 8601 1167 8618 1201
rect 8550 1127 8618 1167
rect 8323 1057 8357 1059
rect 8550 1093 8567 1127
rect 8601 1093 8618 1127
rect 8147 1023 8453 1057
rect 7884 979 7952 1019
rect 7884 945 7901 979
rect 7935 945 7952 979
rect 7884 905 7952 945
rect 7884 871 7901 905
rect 7935 871 7952 905
rect 7884 822 7952 871
rect 8123 957 8157 973
rect 8277 957 8311 973
rect 6999 217 7033 314
rect 7218 313 7286 353
rect 7218 279 7235 313
rect 7269 279 7286 313
rect 6999 167 7033 183
rect 7096 261 7130 277
rect 7096 193 7130 227
rect 6902 123 6936 159
rect 7096 123 7130 159
rect 6936 89 6999 123
rect 7033 89 7096 123
rect 6902 73 6936 89
rect 7096 73 7130 89
rect 7218 239 7286 279
rect 7218 205 7235 239
rect 7269 205 7286 239
rect 7218 165 7286 205
rect 7218 131 7235 165
rect 7269 131 7286 165
rect 7218 91 7286 131
rect 7218 57 7235 91
rect 7269 57 7286 91
rect 7374 333 7408 349
rect 7568 333 7602 349
rect 7753 348 7787 723
rect 8123 757 8157 923
rect 7408 299 7471 333
rect 7505 299 7568 333
rect 7374 261 7408 299
rect 7374 193 7408 227
rect 7568 261 7602 299
rect 7374 123 7408 159
rect 7374 73 7408 89
rect 7471 208 7505 224
rect 7218 34 7286 57
rect 7471 34 7505 174
rect 7568 193 7602 227
rect 7665 314 7787 348
rect 7884 461 7952 544
rect 7884 427 7901 461
rect 7935 427 7952 461
rect 7884 387 7952 427
rect 7884 353 7901 387
rect 7935 353 7952 387
rect 8123 433 8157 723
rect 8123 383 8157 399
rect 8271 923 8277 942
rect 8271 907 8311 923
rect 8271 831 8305 907
rect 8271 433 8305 797
rect 8271 383 8305 399
rect 8419 461 8453 1023
rect 8550 1053 8618 1093
rect 8550 1019 8567 1053
rect 8601 1019 8618 1053
rect 8785 1366 8819 1446
rect 8785 1298 8819 1332
rect 8785 1230 8819 1264
rect 8785 1162 8819 1196
rect 8785 1093 8819 1128
rect 8785 1043 8819 1059
rect 8873 1366 8907 1404
rect 8873 1298 8907 1332
rect 8873 1230 8907 1264
rect 8873 1162 8907 1196
rect 8873 1093 8907 1128
rect 8961 1366 8995 1446
rect 8961 1298 8995 1332
rect 8961 1230 8995 1264
rect 8961 1162 8995 1196
rect 8961 1111 8995 1128
rect 9049 1366 9083 1404
rect 9049 1298 9083 1332
rect 9049 1230 9083 1264
rect 9049 1162 9083 1196
rect 8873 1048 8907 1059
rect 9049 1093 9083 1128
rect 9137 1366 9171 1446
rect 9137 1298 9171 1332
rect 9137 1230 9171 1264
rect 9137 1162 9171 1196
rect 9137 1111 9171 1128
rect 9225 1366 9259 1404
rect 9225 1298 9259 1332
rect 9225 1230 9259 1264
rect 9225 1162 9259 1196
rect 9049 1048 9083 1059
rect 9225 1093 9259 1128
rect 9313 1366 9347 1446
rect 9313 1298 9347 1332
rect 9313 1230 9347 1264
rect 9313 1162 9347 1196
rect 9313 1111 9347 1128
rect 9512 1423 9580 1446
rect 9512 1389 9529 1423
rect 9563 1389 9580 1423
rect 9512 1349 9580 1389
rect 9512 1315 9529 1349
rect 9563 1315 9580 1349
rect 9512 1275 9580 1315
rect 9512 1241 9529 1275
rect 9563 1241 9580 1275
rect 9512 1201 9580 1241
rect 9512 1167 9529 1201
rect 9563 1167 9580 1201
rect 9512 1127 9580 1167
rect 9225 1048 9259 1059
rect 9512 1093 9529 1127
rect 9563 1093 9580 1127
rect 9512 1053 9580 1093
rect 8550 979 8618 1019
rect 8873 1014 9415 1048
rect 8550 945 8567 979
rect 8601 945 8618 979
rect 8550 905 8618 945
rect 8550 871 8567 905
rect 8601 871 8618 905
rect 8550 822 8618 871
rect 8789 957 8823 973
rect 8789 831 8823 923
rect 7665 217 7699 314
rect 7884 313 7952 353
rect 7884 279 7901 313
rect 7935 279 7952 313
rect 7665 167 7699 183
rect 7762 261 7796 277
rect 7762 193 7796 227
rect 7568 123 7602 159
rect 7762 123 7796 159
rect 7602 89 7665 123
rect 7699 89 7762 123
rect 7568 73 7602 89
rect 7762 73 7796 89
rect 7884 239 7952 279
rect 7884 205 7901 239
rect 7935 205 7952 239
rect 7884 165 7952 205
rect 7884 131 7901 165
rect 7935 131 7952 165
rect 7884 91 7952 131
rect 7884 57 7901 91
rect 7935 57 7952 91
rect 8040 333 8074 349
rect 8234 333 8268 349
rect 8419 348 8453 427
rect 8074 299 8137 333
rect 8171 299 8234 333
rect 8040 261 8074 299
rect 8040 193 8074 227
rect 8234 261 8268 299
rect 8040 123 8074 159
rect 8040 73 8074 89
rect 8137 208 8171 224
rect 7884 34 7952 57
rect 8137 34 8171 174
rect 8234 193 8268 227
rect 8331 314 8453 348
rect 8550 461 8618 544
rect 8550 427 8567 461
rect 8601 427 8618 461
rect 8550 387 8618 427
rect 8550 353 8567 387
rect 8601 353 8618 387
rect 8789 433 8823 797
rect 8789 383 8823 399
rect 9011 957 9045 973
rect 9011 905 9045 923
rect 9011 433 9045 871
rect 9011 383 9045 399
rect 9233 957 9267 973
rect 9233 683 9267 923
rect 9233 433 9267 649
rect 9233 383 9267 399
rect 9381 757 9415 1014
rect 9512 1019 9529 1053
rect 9563 1019 9580 1053
rect 9687 1366 9721 1446
rect 9687 1298 9721 1332
rect 9687 1230 9721 1264
rect 9687 1162 9721 1196
rect 9687 1093 9721 1128
rect 9687 1027 9721 1059
rect 9775 1366 9809 1404
rect 9775 1298 9809 1332
rect 9775 1230 9809 1264
rect 9775 1162 9809 1196
rect 9775 1093 9809 1128
rect 9863 1366 9897 1446
rect 9863 1298 9897 1332
rect 9863 1230 9897 1264
rect 9863 1162 9897 1196
rect 9863 1111 9897 1128
rect 9951 1366 9985 1404
rect 9951 1298 9985 1332
rect 9951 1230 9985 1264
rect 9951 1162 9985 1196
rect 9775 1057 9809 1059
rect 9951 1093 9985 1128
rect 10039 1366 10073 1446
rect 10039 1298 10073 1332
rect 10039 1230 10073 1264
rect 10039 1162 10073 1196
rect 10039 1111 10073 1128
rect 10178 1423 10246 1446
rect 10178 1389 10195 1423
rect 10229 1389 10246 1423
rect 10178 1349 10246 1389
rect 10178 1315 10195 1349
rect 10229 1315 10246 1349
rect 10178 1275 10246 1315
rect 10178 1241 10195 1275
rect 10229 1241 10246 1275
rect 10178 1201 10246 1241
rect 10178 1167 10195 1201
rect 10229 1167 10246 1201
rect 10178 1127 10246 1167
rect 9951 1057 9985 1059
rect 10178 1093 10195 1127
rect 10229 1093 10246 1127
rect 9775 1023 10081 1057
rect 9512 979 9580 1019
rect 9512 945 9529 979
rect 9563 945 9580 979
rect 9512 905 9580 945
rect 9512 871 9529 905
rect 9563 871 9580 905
rect 9512 822 9580 871
rect 9751 957 9785 973
rect 9905 957 9939 973
rect 8331 217 8365 314
rect 8550 313 8618 353
rect 8550 279 8567 313
rect 8601 279 8618 313
rect 8331 167 8365 183
rect 8428 261 8462 277
rect 8428 193 8462 227
rect 8234 123 8268 159
rect 8428 123 8462 159
rect 8268 89 8331 123
rect 8365 89 8428 123
rect 8234 73 8268 89
rect 8428 73 8462 89
rect 8550 239 8618 279
rect 8550 205 8567 239
rect 8601 205 8618 239
rect 8550 165 8618 205
rect 8550 131 8567 165
rect 8601 131 8618 165
rect 8550 91 8618 131
rect 8550 57 8567 91
rect 8601 57 8618 91
rect 8685 335 8719 351
rect 8879 335 8913 351
rect 9073 335 9107 351
rect 8719 301 8782 335
rect 8816 301 8879 335
rect 8913 301 8976 335
rect 9010 301 9073 335
rect 8685 263 8719 301
rect 8685 195 8719 229
rect 8879 263 8913 301
rect 9073 285 9107 301
rect 9187 335 9221 351
rect 9381 350 9415 723
rect 9751 757 9785 923
rect 9187 263 9221 301
rect 8685 125 8719 161
rect 8685 75 8719 91
rect 8782 210 8816 226
rect 8550 34 8618 57
rect 8782 34 8816 176
rect 8879 195 8913 229
rect 8977 216 9011 232
rect 9187 216 9221 229
rect 9011 195 9221 216
rect 9011 182 9187 195
rect 8977 166 9011 182
rect 8879 125 8913 161
rect 9284 316 9415 350
rect 9512 461 9580 544
rect 9512 427 9529 461
rect 9563 427 9580 461
rect 9512 387 9580 427
rect 9512 353 9529 387
rect 9563 353 9580 387
rect 9751 433 9785 723
rect 9751 383 9785 399
rect 9899 923 9905 942
rect 9899 907 9939 923
rect 9899 535 9933 907
rect 9899 433 9933 501
rect 9899 383 9933 399
rect 10047 683 10081 1023
rect 10178 1053 10246 1093
rect 10178 1019 10195 1053
rect 10229 1019 10246 1053
rect 10353 1366 10387 1446
rect 10353 1298 10387 1332
rect 10353 1230 10387 1264
rect 10353 1162 10387 1196
rect 10353 1093 10387 1128
rect 10353 1027 10387 1059
rect 10441 1366 10475 1404
rect 10441 1298 10475 1332
rect 10441 1230 10475 1264
rect 10441 1162 10475 1196
rect 10441 1093 10475 1128
rect 10529 1366 10563 1446
rect 10529 1298 10563 1332
rect 10529 1230 10563 1264
rect 10529 1162 10563 1196
rect 10529 1111 10563 1128
rect 10617 1366 10651 1404
rect 10617 1298 10651 1332
rect 10617 1230 10651 1264
rect 10617 1162 10651 1196
rect 10441 1057 10475 1059
rect 10617 1093 10651 1128
rect 10705 1366 10739 1446
rect 10705 1298 10739 1332
rect 10705 1230 10739 1264
rect 10705 1162 10739 1196
rect 10705 1111 10739 1128
rect 10844 1423 10912 1446
rect 10844 1389 10861 1423
rect 10895 1389 10912 1423
rect 10844 1349 10912 1389
rect 10844 1315 10861 1349
rect 10895 1315 10912 1349
rect 10844 1275 10912 1315
rect 10844 1241 10861 1275
rect 10895 1241 10912 1275
rect 10844 1201 10912 1241
rect 10844 1167 10861 1201
rect 10895 1167 10912 1201
rect 10844 1127 10912 1167
rect 10617 1057 10651 1059
rect 10844 1093 10861 1127
rect 10895 1093 10912 1127
rect 10441 1023 10747 1057
rect 10178 979 10246 1019
rect 10178 945 10195 979
rect 10229 945 10246 979
rect 10178 905 10246 945
rect 10178 871 10195 905
rect 10229 871 10246 905
rect 10178 822 10246 871
rect 10417 957 10451 973
rect 10571 957 10605 973
rect 9284 219 9318 316
rect 9512 313 9580 353
rect 9512 279 9529 313
rect 9563 279 9580 313
rect 9284 169 9318 185
rect 9381 263 9415 279
rect 9381 195 9415 229
rect 9073 125 9107 141
rect 8913 91 8976 125
rect 9010 91 9073 125
rect 8879 75 8913 91
rect 9073 75 9107 91
rect 9187 125 9221 161
rect 9381 125 9415 161
rect 9221 91 9284 125
rect 9318 91 9381 125
rect 9187 75 9221 91
rect 9381 75 9415 91
rect 9512 239 9580 279
rect 9512 205 9529 239
rect 9563 205 9580 239
rect 9512 165 9580 205
rect 9512 131 9529 165
rect 9563 131 9580 165
rect 9512 91 9580 131
rect 9512 57 9529 91
rect 9563 57 9580 91
rect 9668 333 9702 349
rect 9862 333 9896 349
rect 10047 348 10081 649
rect 10417 683 10451 923
rect 9702 299 9765 333
rect 9799 299 9862 333
rect 9668 261 9702 299
rect 9668 193 9702 227
rect 9862 261 9896 299
rect 9668 123 9702 159
rect 9668 73 9702 89
rect 9765 208 9799 224
rect 9512 34 9580 57
rect 9765 34 9799 174
rect 9862 193 9896 227
rect 9959 314 10081 348
rect 10178 461 10246 544
rect 10178 427 10195 461
rect 10229 427 10246 461
rect 10178 387 10246 427
rect 10178 353 10195 387
rect 10229 353 10246 387
rect 10417 433 10451 649
rect 10417 383 10451 399
rect 10565 923 10571 942
rect 10565 907 10605 923
rect 10565 831 10599 907
rect 10565 433 10599 797
rect 10565 383 10599 399
rect 10713 683 10747 1023
rect 10844 1053 10912 1093
rect 10844 1019 10861 1053
rect 10895 1019 10912 1053
rect 11019 1366 11053 1446
rect 11019 1298 11053 1332
rect 11019 1230 11053 1264
rect 11019 1162 11053 1196
rect 11019 1093 11053 1128
rect 11019 1027 11053 1059
rect 11107 1366 11141 1404
rect 11107 1298 11141 1332
rect 11107 1230 11141 1264
rect 11107 1162 11141 1196
rect 11107 1093 11141 1128
rect 11195 1366 11229 1446
rect 11195 1298 11229 1332
rect 11195 1230 11229 1264
rect 11195 1162 11229 1196
rect 11195 1111 11229 1128
rect 11283 1366 11317 1404
rect 11283 1298 11317 1332
rect 11283 1230 11317 1264
rect 11283 1162 11317 1196
rect 11107 1057 11141 1059
rect 11283 1093 11317 1128
rect 11371 1366 11405 1446
rect 11371 1298 11405 1332
rect 11371 1230 11405 1264
rect 11371 1162 11405 1196
rect 11371 1111 11405 1128
rect 11510 1423 11578 1446
rect 11510 1389 11527 1423
rect 11561 1389 11578 1423
rect 11510 1349 11578 1389
rect 11510 1315 11527 1349
rect 11561 1315 11578 1349
rect 11510 1275 11578 1315
rect 11510 1241 11527 1275
rect 11561 1241 11578 1275
rect 11510 1201 11578 1241
rect 11510 1167 11527 1201
rect 11561 1167 11578 1201
rect 11510 1127 11578 1167
rect 11283 1057 11317 1059
rect 11510 1093 11527 1127
rect 11561 1093 11578 1127
rect 11107 1023 11413 1057
rect 10844 979 10912 1019
rect 10844 945 10861 979
rect 10895 945 10912 979
rect 10844 905 10912 945
rect 10844 871 10861 905
rect 10895 871 10912 905
rect 10844 822 10912 871
rect 11083 957 11117 973
rect 11237 957 11271 973
rect 9959 217 9993 314
rect 10178 313 10246 353
rect 10178 279 10195 313
rect 10229 279 10246 313
rect 9959 167 9993 183
rect 10056 261 10090 277
rect 10056 193 10090 227
rect 9862 123 9896 159
rect 10056 123 10090 159
rect 9896 89 9959 123
rect 9993 89 10056 123
rect 9862 73 9896 89
rect 10056 73 10090 89
rect 10178 239 10246 279
rect 10178 205 10195 239
rect 10229 205 10246 239
rect 10178 165 10246 205
rect 10178 131 10195 165
rect 10229 131 10246 165
rect 10178 91 10246 131
rect 10178 57 10195 91
rect 10229 57 10246 91
rect 10334 333 10368 349
rect 10528 333 10562 349
rect 10713 348 10747 649
rect 11083 683 11117 923
rect 10368 299 10431 333
rect 10465 299 10528 333
rect 10334 261 10368 299
rect 10334 193 10368 227
rect 10528 261 10562 299
rect 10334 123 10368 159
rect 10334 73 10368 89
rect 10431 208 10465 224
rect 10178 34 10246 57
rect 10431 34 10465 174
rect 10528 193 10562 227
rect 10625 314 10747 348
rect 10844 461 10912 544
rect 10844 427 10861 461
rect 10895 427 10912 461
rect 10844 387 10912 427
rect 10844 353 10861 387
rect 10895 353 10912 387
rect 11083 433 11117 649
rect 11083 383 11117 399
rect 11231 923 11237 942
rect 11231 907 11271 923
rect 11231 905 11265 907
rect 11231 433 11265 871
rect 11231 383 11265 399
rect 11379 831 11413 1023
rect 11510 1053 11578 1093
rect 11510 1019 11527 1053
rect 11561 1019 11578 1053
rect 11685 1366 11719 1446
rect 11685 1298 11719 1332
rect 11685 1230 11719 1264
rect 11685 1162 11719 1196
rect 11685 1093 11719 1128
rect 11685 1027 11719 1059
rect 11773 1366 11807 1404
rect 11773 1298 11807 1332
rect 11773 1230 11807 1264
rect 11773 1162 11807 1196
rect 11773 1093 11807 1128
rect 11861 1366 11895 1446
rect 11861 1298 11895 1332
rect 11861 1230 11895 1264
rect 11861 1162 11895 1196
rect 11861 1111 11895 1128
rect 11949 1366 11983 1404
rect 11949 1298 11983 1332
rect 11949 1230 11983 1264
rect 11949 1162 11983 1196
rect 11773 1057 11807 1059
rect 11949 1093 11983 1128
rect 12037 1366 12071 1446
rect 12037 1298 12071 1332
rect 12037 1230 12071 1264
rect 12037 1162 12071 1196
rect 12037 1111 12071 1128
rect 12176 1423 12244 1446
rect 12176 1389 12193 1423
rect 12227 1389 12244 1423
rect 12176 1349 12244 1389
rect 12176 1315 12193 1349
rect 12227 1315 12244 1349
rect 12176 1275 12244 1315
rect 12176 1241 12193 1275
rect 12227 1241 12244 1275
rect 12176 1201 12244 1241
rect 12176 1167 12193 1201
rect 12227 1167 12244 1201
rect 12176 1127 12244 1167
rect 11949 1057 11983 1059
rect 12176 1093 12193 1127
rect 12227 1093 12244 1127
rect 11773 1023 12079 1057
rect 11510 979 11578 1019
rect 11510 945 11527 979
rect 11561 945 11578 979
rect 11510 905 11578 945
rect 11510 871 11527 905
rect 11561 871 11578 905
rect 11510 822 11578 871
rect 11749 957 11783 973
rect 11903 957 11937 973
rect 10625 217 10659 314
rect 10844 313 10912 353
rect 10844 279 10861 313
rect 10895 279 10912 313
rect 10625 167 10659 183
rect 10722 261 10756 277
rect 10722 193 10756 227
rect 10528 123 10562 159
rect 10722 123 10756 159
rect 10562 89 10625 123
rect 10659 89 10722 123
rect 10528 73 10562 89
rect 10722 73 10756 89
rect 10844 239 10912 279
rect 10844 205 10861 239
rect 10895 205 10912 239
rect 10844 165 10912 205
rect 10844 131 10861 165
rect 10895 131 10912 165
rect 10844 91 10912 131
rect 10844 57 10861 91
rect 10895 57 10912 91
rect 11000 333 11034 349
rect 11194 333 11228 349
rect 11379 348 11413 797
rect 11749 757 11783 923
rect 11034 299 11097 333
rect 11131 299 11194 333
rect 11000 261 11034 299
rect 11000 193 11034 227
rect 11194 261 11228 299
rect 11000 123 11034 159
rect 11000 73 11034 89
rect 11097 208 11131 224
rect 10844 34 10912 57
rect 11097 34 11131 174
rect 11194 193 11228 227
rect 11291 314 11413 348
rect 11510 461 11578 544
rect 11510 427 11527 461
rect 11561 427 11578 461
rect 11510 387 11578 427
rect 11510 353 11527 387
rect 11561 353 11578 387
rect 11749 433 11783 723
rect 11749 383 11783 399
rect 11897 923 11903 942
rect 11897 907 11937 923
rect 11897 757 11931 907
rect 11897 433 11931 723
rect 11897 383 11931 399
rect 12045 905 12079 1023
rect 11291 217 11325 314
rect 11510 313 11578 353
rect 11510 279 11527 313
rect 11561 279 11578 313
rect 11291 167 11325 183
rect 11388 261 11422 277
rect 11388 193 11422 227
rect 11194 123 11228 159
rect 11388 123 11422 159
rect 11228 89 11291 123
rect 11325 89 11388 123
rect 11194 73 11228 89
rect 11388 73 11422 89
rect 11510 239 11578 279
rect 11510 205 11527 239
rect 11561 205 11578 239
rect 11510 165 11578 205
rect 11510 131 11527 165
rect 11561 131 11578 165
rect 11510 91 11578 131
rect 11510 57 11527 91
rect 11561 57 11578 91
rect 11666 333 11700 349
rect 11860 333 11894 349
rect 12045 348 12079 871
rect 12176 1053 12244 1093
rect 12176 1019 12193 1053
rect 12227 1019 12244 1053
rect 12351 1366 12385 1446
rect 12351 1298 12385 1332
rect 12351 1230 12385 1264
rect 12351 1162 12385 1196
rect 12351 1093 12385 1128
rect 12351 1027 12385 1059
rect 12439 1366 12473 1404
rect 12439 1298 12473 1332
rect 12439 1230 12473 1264
rect 12439 1162 12473 1196
rect 12439 1093 12473 1128
rect 12527 1366 12561 1446
rect 12527 1298 12561 1332
rect 12527 1230 12561 1264
rect 12527 1162 12561 1196
rect 12527 1111 12561 1128
rect 12615 1366 12649 1404
rect 12615 1298 12649 1332
rect 12615 1230 12649 1264
rect 12615 1162 12649 1196
rect 12439 1057 12473 1059
rect 12615 1093 12649 1128
rect 12703 1366 12737 1446
rect 12703 1298 12737 1332
rect 12703 1230 12737 1264
rect 12703 1162 12737 1196
rect 12703 1111 12737 1128
rect 12842 1423 12910 1446
rect 12842 1389 12859 1423
rect 12893 1389 12910 1423
rect 12842 1349 12910 1389
rect 12842 1315 12859 1349
rect 12893 1315 12910 1349
rect 12842 1275 12910 1315
rect 12842 1241 12859 1275
rect 12893 1241 12910 1275
rect 12842 1201 12910 1241
rect 12842 1167 12859 1201
rect 12893 1167 12910 1201
rect 12842 1127 12910 1167
rect 12615 1057 12649 1059
rect 12842 1093 12859 1127
rect 12893 1093 12910 1127
rect 12439 1023 12745 1057
rect 12176 979 12244 1019
rect 12176 945 12193 979
rect 12227 945 12244 979
rect 12176 905 12244 945
rect 12176 871 12193 905
rect 12227 871 12244 905
rect 12176 822 12244 871
rect 12415 957 12449 973
rect 12569 957 12603 973
rect 12415 905 12449 923
rect 11700 299 11763 333
rect 11797 299 11860 333
rect 11666 261 11700 299
rect 11666 193 11700 227
rect 11860 261 11894 299
rect 11666 123 11700 159
rect 11666 73 11700 89
rect 11763 208 11797 224
rect 11510 34 11578 57
rect 11763 34 11797 174
rect 11860 193 11894 227
rect 11957 314 12079 348
rect 12176 461 12244 544
rect 12176 427 12193 461
rect 12227 427 12244 461
rect 12176 387 12244 427
rect 12176 353 12193 387
rect 12227 353 12244 387
rect 12415 433 12449 871
rect 12415 383 12449 399
rect 12563 923 12569 942
rect 12563 907 12603 923
rect 12563 831 12597 907
rect 12563 433 12597 797
rect 12563 383 12597 399
rect 12711 757 12745 1023
rect 12842 1053 12910 1093
rect 12842 1019 12859 1053
rect 12893 1019 12910 1053
rect 13017 1365 13051 1446
rect 13017 1297 13051 1331
rect 13017 1229 13051 1263
rect 13017 1161 13051 1195
rect 13017 1093 13051 1127
rect 13017 1025 13051 1059
rect 13105 1365 13141 1399
rect 13193 1365 13227 1446
rect 13105 1297 13139 1331
rect 13105 1229 13139 1263
rect 13105 1161 13139 1195
rect 13105 1093 13139 1127
rect 13193 1297 13227 1331
rect 13193 1229 13227 1263
rect 13193 1161 13227 1195
rect 13193 1111 13227 1127
rect 13281 1365 13315 1399
rect 13281 1297 13315 1331
rect 13281 1229 13315 1263
rect 13281 1161 13315 1195
rect 13281 1059 13315 1127
rect 13105 1025 13281 1059
rect 13369 1365 13403 1446
rect 13369 1297 13403 1331
rect 13369 1229 13403 1263
rect 13369 1161 13403 1195
rect 13369 1093 13403 1127
rect 13369 1025 13403 1059
rect 13508 1423 13576 1446
rect 13508 1389 13525 1423
rect 13559 1389 13576 1423
rect 14174 1423 14242 1446
rect 13508 1349 13576 1389
rect 13508 1315 13525 1349
rect 13559 1315 13576 1349
rect 13508 1275 13576 1315
rect 13508 1241 13525 1275
rect 13559 1241 13576 1275
rect 13508 1201 13576 1241
rect 13508 1167 13525 1201
rect 13559 1167 13576 1201
rect 13508 1127 13576 1167
rect 13508 1093 13525 1127
rect 13559 1093 13576 1127
rect 13508 1053 13576 1093
rect 12842 979 12910 1019
rect 13281 1009 13315 1025
rect 13508 1019 13525 1053
rect 13559 1019 13576 1053
rect 12842 945 12859 979
rect 12893 945 12910 979
rect 13508 979 13576 1019
rect 13681 1365 14067 1399
rect 13681 1297 13715 1331
rect 13681 1229 13715 1263
rect 13681 1161 13715 1195
rect 13681 1059 13715 1127
rect 13769 1297 13803 1313
rect 13769 1229 13803 1263
rect 13769 1161 13803 1195
rect 13769 1093 13803 1127
rect 13857 1297 13891 1331
rect 13857 1229 13891 1263
rect 13857 1161 13891 1195
rect 13857 1111 13891 1127
rect 13945 1297 13979 1313
rect 13945 1229 13979 1263
rect 13945 1161 13979 1195
rect 13945 1059 13979 1127
rect 14033 1297 14067 1331
rect 14033 1229 14067 1263
rect 14033 1161 14067 1195
rect 14033 1075 14067 1127
rect 14174 1389 14191 1423
rect 14225 1389 14242 1423
rect 14840 1423 14908 1446
rect 14174 1349 14242 1389
rect 14174 1315 14191 1349
rect 14225 1315 14242 1349
rect 14174 1275 14242 1315
rect 14174 1241 14191 1275
rect 14225 1241 14242 1275
rect 14174 1201 14242 1241
rect 14174 1167 14191 1201
rect 14225 1167 14242 1201
rect 14174 1127 14242 1167
rect 14174 1093 14191 1127
rect 14225 1093 14242 1127
rect 13769 1025 13945 1059
rect 13681 1009 13715 1025
rect 13945 1009 13979 1025
rect 14174 1053 14242 1093
rect 14174 1019 14191 1053
rect 14225 1019 14242 1053
rect 12842 905 12910 945
rect 12842 871 12859 905
rect 12893 871 12910 905
rect 12842 822 12910 871
rect 13007 958 13041 974
rect 13237 958 13271 974
rect 13007 905 13041 924
rect 11957 217 11991 314
rect 12176 313 12244 353
rect 12176 279 12193 313
rect 12227 279 12244 313
rect 11957 167 11991 183
rect 12054 261 12088 277
rect 12054 193 12088 227
rect 11860 123 11894 159
rect 12054 123 12088 159
rect 11894 89 11957 123
rect 11991 89 12054 123
rect 11860 73 11894 89
rect 12054 73 12088 89
rect 12176 239 12244 279
rect 12176 205 12193 239
rect 12227 205 12244 239
rect 12176 165 12244 205
rect 12176 131 12193 165
rect 12227 131 12244 165
rect 12176 91 12244 131
rect 12176 57 12193 91
rect 12227 57 12244 91
rect 12332 333 12366 349
rect 12526 333 12560 349
rect 12711 348 12745 723
rect 13007 757 13041 871
rect 12366 299 12429 333
rect 12463 299 12526 333
rect 12332 261 12366 299
rect 12332 193 12366 227
rect 12526 261 12560 299
rect 12332 123 12366 159
rect 12332 73 12366 89
rect 12429 208 12463 224
rect 12176 34 12244 57
rect 12429 34 12463 174
rect 12526 193 12560 227
rect 12623 314 12745 348
rect 12842 461 12910 544
rect 12842 427 12859 461
rect 12893 427 12910 461
rect 12842 387 12910 427
rect 12842 353 12859 387
rect 12893 353 12910 387
rect 13007 433 13041 723
rect 13007 383 13041 399
rect 13229 924 13237 942
rect 13229 908 13271 924
rect 13508 945 13525 979
rect 13559 945 13576 979
rect 14174 979 14242 1019
rect 14349 1365 14735 1399
rect 14349 1297 14383 1331
rect 14349 1229 14383 1263
rect 14349 1161 14383 1195
rect 14349 1059 14383 1127
rect 14437 1297 14471 1313
rect 14437 1229 14471 1263
rect 14437 1161 14471 1195
rect 14437 1093 14471 1127
rect 14525 1297 14559 1331
rect 14525 1229 14559 1263
rect 14525 1161 14559 1195
rect 14525 1111 14559 1127
rect 14613 1297 14647 1313
rect 14613 1229 14647 1263
rect 14613 1161 14647 1195
rect 14613 1093 14647 1127
rect 14701 1297 14735 1331
rect 14701 1229 14735 1263
rect 14701 1161 14735 1195
rect 14701 1111 14735 1127
rect 14840 1389 14857 1423
rect 14891 1389 14908 1423
rect 14840 1349 14908 1389
rect 14840 1315 14857 1349
rect 14891 1315 14908 1349
rect 14840 1275 14908 1315
rect 14840 1241 14857 1275
rect 14891 1241 14908 1275
rect 14840 1201 14908 1241
rect 14840 1167 14857 1201
rect 14891 1167 14908 1201
rect 14840 1127 14908 1167
rect 14840 1093 14857 1127
rect 14891 1093 14908 1127
rect 14437 1025 14743 1059
rect 14349 1009 14383 1025
rect 13229 831 13263 908
rect 13508 905 13576 945
rect 13508 871 13525 905
rect 13559 871 13576 905
rect 13508 822 13576 871
rect 13747 958 13781 974
rect 13747 905 13781 924
rect 13229 461 13263 797
rect 13229 383 13263 399
rect 13508 461 13576 544
rect 13508 427 13525 461
rect 13559 427 13576 461
rect 13508 387 13576 427
rect 12623 217 12657 314
rect 12842 313 12910 353
rect 13508 353 13525 387
rect 13559 353 13576 387
rect 13747 433 13781 871
rect 13747 383 13781 399
rect 14043 958 14077 974
rect 14043 609 14077 924
rect 14174 945 14191 979
rect 14225 945 14242 979
rect 14174 905 14242 945
rect 14174 871 14191 905
rect 14225 871 14242 905
rect 14174 822 14242 871
rect 14339 958 14373 974
rect 14043 433 14077 575
rect 14043 383 14077 399
rect 14174 461 14242 544
rect 14174 427 14191 461
rect 14225 427 14242 461
rect 14174 387 14242 427
rect 12842 279 12859 313
rect 12893 279 12910 313
rect 12623 167 12657 183
rect 12720 261 12754 277
rect 12720 193 12754 227
rect 12526 123 12560 159
rect 12720 123 12754 159
rect 12560 89 12623 123
rect 12657 89 12720 123
rect 12526 73 12560 89
rect 12720 73 12754 89
rect 12842 239 12910 279
rect 12842 205 12859 239
rect 12893 205 12910 239
rect 12842 165 12910 205
rect 12842 131 12859 165
rect 12893 131 12910 165
rect 12842 91 12910 131
rect 12842 57 12859 91
rect 12893 57 12910 91
rect 12998 333 13032 349
rect 13192 333 13226 349
rect 13032 299 13095 333
rect 13129 299 13192 333
rect 12998 261 13032 299
rect 12998 193 13032 227
rect 13192 261 13226 299
rect 13386 333 13420 349
rect 13289 253 13323 269
rect 12998 123 13032 159
rect 12998 73 13032 89
rect 13095 208 13129 224
rect 12842 34 12910 57
rect 13095 34 13129 174
rect 13192 193 13226 227
rect 13288 219 13289 234
rect 13288 217 13323 219
rect 13322 203 13323 217
rect 13386 261 13420 299
rect 13288 167 13322 183
rect 13386 193 13420 227
rect 13192 123 13226 159
rect 13386 123 13420 159
rect 13226 89 13288 123
rect 13322 89 13386 123
rect 13192 73 13226 89
rect 13386 73 13420 89
rect 13508 313 13576 353
rect 14174 353 14191 387
rect 14225 353 14242 387
rect 14339 433 14373 924
rect 14339 383 14373 399
rect 14561 958 14599 974
rect 14561 924 14565 958
rect 14561 908 14599 924
rect 14561 831 14595 908
rect 14561 433 14595 797
rect 14561 383 14595 399
rect 13508 279 13525 313
rect 13559 279 13576 313
rect 13508 239 13576 279
rect 13508 205 13525 239
rect 13559 205 13576 239
rect 13508 165 13576 205
rect 13508 131 13525 165
rect 13559 131 13576 165
rect 13508 91 13576 131
rect 13508 57 13525 91
rect 13559 57 13576 91
rect 13664 333 13698 349
rect 13858 333 13892 349
rect 13698 299 13761 333
rect 13795 299 13858 333
rect 13664 261 13698 299
rect 13664 193 13698 227
rect 13858 261 13892 299
rect 14052 333 14086 349
rect 13664 123 13698 159
rect 13664 73 13698 89
rect 13761 208 13795 224
rect 13508 34 13576 57
rect 13761 34 13795 174
rect 13858 193 13892 227
rect 13955 253 13989 269
rect 13955 217 13989 219
rect 13955 167 13989 183
rect 14052 261 14086 299
rect 14052 193 14086 227
rect 13858 123 13892 159
rect 14052 123 14086 159
rect 13892 89 13955 123
rect 13989 89 14052 123
rect 13858 73 13892 89
rect 14052 73 14086 89
rect 14174 313 14242 353
rect 14174 279 14191 313
rect 14225 279 14242 313
rect 14174 239 14242 279
rect 14174 205 14191 239
rect 14225 205 14242 239
rect 14174 165 14242 205
rect 14174 131 14191 165
rect 14225 131 14242 165
rect 14174 91 14242 131
rect 14174 57 14191 91
rect 14225 57 14242 91
rect 14330 333 14364 349
rect 14524 333 14558 349
rect 14709 346 14743 1025
rect 14840 1053 14908 1093
rect 14840 1019 14857 1053
rect 14891 1019 14908 1053
rect 14840 979 14908 1019
rect 14840 945 14857 979
rect 14891 945 14908 979
rect 14840 905 14908 945
rect 14840 871 14857 905
rect 14891 871 14908 905
rect 14840 822 14908 871
rect 14364 299 14427 333
rect 14461 299 14524 333
rect 14330 261 14364 299
rect 14330 193 14364 227
rect 14524 261 14558 299
rect 14330 123 14364 159
rect 14330 73 14364 89
rect 14427 208 14461 224
rect 14174 34 14242 57
rect 14427 34 14461 174
rect 14524 193 14558 227
rect 14621 312 14743 346
rect 14840 461 14908 544
rect 14840 427 14857 461
rect 14891 427 14908 461
rect 14840 387 14908 427
rect 14840 353 14857 387
rect 14891 353 14908 387
rect 14840 313 14908 353
rect 14621 253 14655 312
rect 14840 279 14857 313
rect 14891 279 14908 313
rect 14621 217 14655 219
rect 14621 167 14655 183
rect 14718 261 14752 278
rect 14718 193 14752 227
rect 14524 123 14558 159
rect 14718 123 14752 159
rect 14558 89 14621 123
rect 14655 89 14718 123
rect 14524 73 14558 89
rect 14718 73 14752 89
rect 14840 239 14908 279
rect 14840 205 14857 239
rect 14891 205 14908 239
rect 14840 165 14908 205
rect 14840 131 14857 165
rect 14891 131 14908 165
rect 14840 91 14908 131
rect 14840 57 14857 91
rect 14891 57 14908 91
rect 14840 34 14908 57
rect -34 17 14908 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5163 17
rect 5197 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5533 17
rect 5567 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5755 17
rect 5789 -17 5829 17
rect 5863 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6125 17
rect 6159 -17 6199 17
rect 6233 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6495 17
rect 6529 -17 6643 17
rect 6677 -17 6717 17
rect 6751 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7087 17
rect 7121 -17 7161 17
rect 7195 -17 7309 17
rect 7343 -17 7383 17
rect 7417 -17 7457 17
rect 7491 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7679 17
rect 7713 -17 7753 17
rect 7787 -17 7827 17
rect 7861 -17 7975 17
rect 8009 -17 8049 17
rect 8083 -17 8123 17
rect 8157 -17 8197 17
rect 8231 -17 8271 17
rect 8305 -17 8345 17
rect 8379 -17 8419 17
rect 8453 -17 8493 17
rect 8527 -17 8641 17
rect 8675 -17 8715 17
rect 8749 -17 8789 17
rect 8823 -17 8863 17
rect 8897 -17 8937 17
rect 8971 -17 9011 17
rect 9045 -17 9085 17
rect 9119 -17 9159 17
rect 9193 -17 9233 17
rect 9267 -17 9307 17
rect 9341 -17 9381 17
rect 9415 -17 9455 17
rect 9489 -17 9603 17
rect 9637 -17 9677 17
rect 9711 -17 9751 17
rect 9785 -17 9825 17
rect 9859 -17 9899 17
rect 9933 -17 9973 17
rect 10007 -17 10047 17
rect 10081 -17 10121 17
rect 10155 -17 10269 17
rect 10303 -17 10343 17
rect 10377 -17 10417 17
rect 10451 -17 10491 17
rect 10525 -17 10565 17
rect 10599 -17 10639 17
rect 10673 -17 10713 17
rect 10747 -17 10787 17
rect 10821 -17 10935 17
rect 10969 -17 11009 17
rect 11043 -17 11083 17
rect 11117 -17 11157 17
rect 11191 -17 11231 17
rect 11265 -17 11305 17
rect 11339 -17 11379 17
rect 11413 -17 11453 17
rect 11487 -17 11601 17
rect 11635 -17 11675 17
rect 11709 -17 11749 17
rect 11783 -17 11823 17
rect 11857 -17 11897 17
rect 11931 -17 11971 17
rect 12005 -17 12045 17
rect 12079 -17 12119 17
rect 12153 -17 12267 17
rect 12301 -17 12341 17
rect 12375 -17 12415 17
rect 12449 -17 12489 17
rect 12523 -17 12563 17
rect 12597 -17 12637 17
rect 12671 -17 12711 17
rect 12745 -17 12785 17
rect 12819 -17 12933 17
rect 12967 -17 13007 17
rect 13041 -17 13081 17
rect 13115 -17 13155 17
rect 13189 -17 13229 17
rect 13263 -17 13303 17
rect 13337 -17 13377 17
rect 13411 -17 13451 17
rect 13485 -17 13599 17
rect 13633 -17 13673 17
rect 13707 -17 13747 17
rect 13781 -17 13821 17
rect 13855 -17 13895 17
rect 13929 -17 13969 17
rect 14003 -17 14043 17
rect 14077 -17 14117 17
rect 14151 -17 14265 17
rect 14299 -17 14339 17
rect 14373 -17 14413 17
rect 14447 -17 14487 17
rect 14521 -17 14561 17
rect 14595 -17 14635 17
rect 14669 -17 14709 17
rect 14743 -17 14783 17
rect 14817 -17 14908 17
rect -34 -34 14908 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4497 1463 4531 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4793 1463 4827 1497
rect 4867 1463 4901 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5089 1463 5123 1497
rect 5163 1463 5197 1497
rect 5311 1463 5345 1497
rect 5385 1463 5419 1497
rect 5459 1463 5493 1497
rect 5533 1463 5567 1497
rect 5607 1463 5641 1497
rect 5681 1463 5715 1497
rect 5755 1463 5789 1497
rect 5829 1463 5863 1497
rect 5977 1463 6011 1497
rect 6051 1463 6085 1497
rect 6125 1463 6159 1497
rect 6199 1463 6233 1497
rect 6273 1463 6307 1497
rect 6347 1463 6381 1497
rect 6421 1463 6455 1497
rect 6495 1463 6529 1497
rect 6643 1463 6677 1497
rect 6717 1463 6751 1497
rect 6791 1463 6825 1497
rect 6865 1463 6899 1497
rect 6939 1463 6973 1497
rect 7013 1463 7047 1497
rect 7087 1463 7121 1497
rect 7161 1463 7195 1497
rect 7309 1463 7343 1497
rect 7383 1463 7417 1497
rect 7457 1463 7491 1497
rect 7531 1463 7565 1497
rect 7605 1463 7639 1497
rect 7679 1463 7713 1497
rect 7753 1463 7787 1497
rect 7827 1463 7861 1497
rect 7975 1463 8009 1497
rect 8049 1463 8083 1497
rect 8123 1463 8157 1497
rect 8197 1463 8231 1497
rect 8271 1463 8305 1497
rect 8345 1463 8379 1497
rect 8419 1463 8453 1497
rect 8493 1463 8527 1497
rect 8641 1463 8675 1497
rect 8715 1463 8749 1497
rect 8789 1463 8823 1497
rect 8863 1463 8897 1497
rect 8937 1463 8971 1497
rect 9011 1463 9045 1497
rect 9085 1463 9119 1497
rect 9159 1463 9193 1497
rect 9233 1463 9267 1497
rect 9307 1463 9341 1497
rect 9381 1463 9415 1497
rect 9455 1463 9489 1497
rect 9603 1463 9637 1497
rect 9677 1463 9711 1497
rect 9751 1463 9785 1497
rect 9825 1463 9859 1497
rect 9899 1463 9933 1497
rect 9973 1463 10007 1497
rect 10047 1463 10081 1497
rect 10121 1463 10155 1497
rect 10269 1463 10303 1497
rect 10343 1463 10377 1497
rect 10417 1463 10451 1497
rect 10491 1463 10525 1497
rect 10565 1463 10599 1497
rect 10639 1463 10673 1497
rect 10713 1463 10747 1497
rect 10787 1463 10821 1497
rect 10935 1463 10969 1497
rect 11009 1463 11043 1497
rect 11083 1463 11117 1497
rect 11157 1463 11191 1497
rect 11231 1463 11265 1497
rect 11305 1463 11339 1497
rect 11379 1463 11413 1497
rect 11453 1463 11487 1497
rect 11601 1463 11635 1497
rect 11675 1463 11709 1497
rect 11749 1463 11783 1497
rect 11823 1463 11857 1497
rect 11897 1463 11931 1497
rect 11971 1463 12005 1497
rect 12045 1463 12079 1497
rect 12119 1463 12153 1497
rect 12267 1463 12301 1497
rect 12341 1463 12375 1497
rect 12415 1463 12449 1497
rect 12489 1463 12523 1497
rect 12563 1463 12597 1497
rect 12637 1463 12671 1497
rect 12711 1463 12745 1497
rect 12785 1463 12819 1497
rect 12933 1463 12967 1497
rect 13007 1463 13041 1497
rect 13081 1463 13115 1497
rect 13155 1463 13189 1497
rect 13229 1463 13263 1497
rect 13303 1463 13337 1497
rect 13377 1463 13411 1497
rect 13451 1463 13485 1497
rect 13599 1463 13633 1497
rect 13673 1463 13707 1497
rect 13747 1463 13781 1497
rect 13821 1463 13855 1497
rect 13895 1463 13929 1497
rect 13969 1463 14003 1497
rect 14043 1463 14077 1497
rect 14117 1463 14151 1497
rect 14265 1463 14299 1497
rect 14339 1463 14373 1497
rect 14413 1463 14447 1497
rect 14487 1463 14521 1497
rect 14561 1463 14595 1497
rect 14635 1463 14669 1497
rect 14709 1463 14743 1497
rect 14783 1463 14817 1497
rect 205 797 239 831
rect 427 871 461 905
rect 649 649 683 683
rect 797 723 831 757
rect 1167 723 1201 757
rect 1315 501 1349 535
rect 1463 649 1497 683
rect 1833 649 1867 683
rect 1981 797 2015 831
rect 2129 649 2163 683
rect 2499 649 2533 683
rect 2647 871 2681 905
rect 2795 797 2829 831
rect 3165 723 3199 757
rect 3313 575 3347 609
rect 3461 723 3495 757
rect 3831 723 3865 757
rect 3979 797 4013 831
rect 4127 575 4161 609
rect 4497 797 4531 831
rect 4719 871 4753 905
rect 4941 649 4975 683
rect 5089 723 5123 757
rect 5459 723 5493 757
rect 5607 501 5641 535
rect 5755 649 5789 683
rect 6125 649 6159 683
rect 6273 797 6307 831
rect 6421 649 6455 683
rect 6791 649 6825 683
rect 6939 871 6973 905
rect 7087 797 7121 831
rect 7457 723 7491 757
rect 7605 433 7639 461
rect 7605 427 7639 433
rect 7753 723 7787 757
rect 8123 723 8157 757
rect 8271 797 8305 831
rect 8789 797 8823 831
rect 8419 427 8453 461
rect 9011 871 9045 905
rect 9233 649 9267 683
rect 9381 723 9415 757
rect 9751 723 9785 757
rect 9899 501 9933 535
rect 10047 649 10081 683
rect 10417 649 10451 683
rect 10565 797 10599 831
rect 10713 649 10747 683
rect 11083 649 11117 683
rect 11231 871 11265 905
rect 11379 797 11413 831
rect 11749 723 11783 757
rect 11897 723 11931 757
rect 12045 871 12079 905
rect 12415 871 12449 905
rect 12563 797 12597 831
rect 13281 1025 13315 1059
rect 13681 1025 13715 1059
rect 13945 1025 13979 1059
rect 13007 871 13041 905
rect 12711 723 12745 757
rect 13007 723 13041 757
rect 14349 1025 14383 1059
rect 13229 797 13263 831
rect 13747 871 13781 905
rect 13229 433 13263 461
rect 13229 427 13263 433
rect 14043 575 14077 609
rect 14043 399 14077 433
rect 13289 219 13323 253
rect 14339 399 14373 433
rect 14561 797 14595 831
rect 13955 219 13989 253
rect 14621 219 14655 253
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4497 -17 4531 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4793 -17 4827 17
rect 4867 -17 4901 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5089 -17 5123 17
rect 5163 -17 5197 17
rect 5311 -17 5345 17
rect 5385 -17 5419 17
rect 5459 -17 5493 17
rect 5533 -17 5567 17
rect 5607 -17 5641 17
rect 5681 -17 5715 17
rect 5755 -17 5789 17
rect 5829 -17 5863 17
rect 5977 -17 6011 17
rect 6051 -17 6085 17
rect 6125 -17 6159 17
rect 6199 -17 6233 17
rect 6273 -17 6307 17
rect 6347 -17 6381 17
rect 6421 -17 6455 17
rect 6495 -17 6529 17
rect 6643 -17 6677 17
rect 6717 -17 6751 17
rect 6791 -17 6825 17
rect 6865 -17 6899 17
rect 6939 -17 6973 17
rect 7013 -17 7047 17
rect 7087 -17 7121 17
rect 7161 -17 7195 17
rect 7309 -17 7343 17
rect 7383 -17 7417 17
rect 7457 -17 7491 17
rect 7531 -17 7565 17
rect 7605 -17 7639 17
rect 7679 -17 7713 17
rect 7753 -17 7787 17
rect 7827 -17 7861 17
rect 7975 -17 8009 17
rect 8049 -17 8083 17
rect 8123 -17 8157 17
rect 8197 -17 8231 17
rect 8271 -17 8305 17
rect 8345 -17 8379 17
rect 8419 -17 8453 17
rect 8493 -17 8527 17
rect 8641 -17 8675 17
rect 8715 -17 8749 17
rect 8789 -17 8823 17
rect 8863 -17 8897 17
rect 8937 -17 8971 17
rect 9011 -17 9045 17
rect 9085 -17 9119 17
rect 9159 -17 9193 17
rect 9233 -17 9267 17
rect 9307 -17 9341 17
rect 9381 -17 9415 17
rect 9455 -17 9489 17
rect 9603 -17 9637 17
rect 9677 -17 9711 17
rect 9751 -17 9785 17
rect 9825 -17 9859 17
rect 9899 -17 9933 17
rect 9973 -17 10007 17
rect 10047 -17 10081 17
rect 10121 -17 10155 17
rect 10269 -17 10303 17
rect 10343 -17 10377 17
rect 10417 -17 10451 17
rect 10491 -17 10525 17
rect 10565 -17 10599 17
rect 10639 -17 10673 17
rect 10713 -17 10747 17
rect 10787 -17 10821 17
rect 10935 -17 10969 17
rect 11009 -17 11043 17
rect 11083 -17 11117 17
rect 11157 -17 11191 17
rect 11231 -17 11265 17
rect 11305 -17 11339 17
rect 11379 -17 11413 17
rect 11453 -17 11487 17
rect 11601 -17 11635 17
rect 11675 -17 11709 17
rect 11749 -17 11783 17
rect 11823 -17 11857 17
rect 11897 -17 11931 17
rect 11971 -17 12005 17
rect 12045 -17 12079 17
rect 12119 -17 12153 17
rect 12267 -17 12301 17
rect 12341 -17 12375 17
rect 12415 -17 12449 17
rect 12489 -17 12523 17
rect 12563 -17 12597 17
rect 12637 -17 12671 17
rect 12711 -17 12745 17
rect 12785 -17 12819 17
rect 12933 -17 12967 17
rect 13007 -17 13041 17
rect 13081 -17 13115 17
rect 13155 -17 13189 17
rect 13229 -17 13263 17
rect 13303 -17 13337 17
rect 13377 -17 13411 17
rect 13451 -17 13485 17
rect 13599 -17 13633 17
rect 13673 -17 13707 17
rect 13747 -17 13781 17
rect 13821 -17 13855 17
rect 13895 -17 13929 17
rect 13969 -17 14003 17
rect 14043 -17 14077 17
rect 14117 -17 14151 17
rect 14265 -17 14299 17
rect 14339 -17 14373 17
rect 14413 -17 14447 17
rect 14487 -17 14521 17
rect 14561 -17 14595 17
rect 14635 -17 14669 17
rect 14709 -17 14743 17
rect 14783 -17 14817 17
<< metal1 >>
rect -34 1497 14908 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5163 1497
rect 5197 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5533 1497
rect 5567 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5755 1497
rect 5789 1463 5829 1497
rect 5863 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6125 1497
rect 6159 1463 6199 1497
rect 6233 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6495 1497
rect 6529 1463 6643 1497
rect 6677 1463 6717 1497
rect 6751 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7087 1497
rect 7121 1463 7161 1497
rect 7195 1463 7309 1497
rect 7343 1463 7383 1497
rect 7417 1463 7457 1497
rect 7491 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7679 1497
rect 7713 1463 7753 1497
rect 7787 1463 7827 1497
rect 7861 1463 7975 1497
rect 8009 1463 8049 1497
rect 8083 1463 8123 1497
rect 8157 1463 8197 1497
rect 8231 1463 8271 1497
rect 8305 1463 8345 1497
rect 8379 1463 8419 1497
rect 8453 1463 8493 1497
rect 8527 1463 8641 1497
rect 8675 1463 8715 1497
rect 8749 1463 8789 1497
rect 8823 1463 8863 1497
rect 8897 1463 8937 1497
rect 8971 1463 9011 1497
rect 9045 1463 9085 1497
rect 9119 1463 9159 1497
rect 9193 1463 9233 1497
rect 9267 1463 9307 1497
rect 9341 1463 9381 1497
rect 9415 1463 9455 1497
rect 9489 1463 9603 1497
rect 9637 1463 9677 1497
rect 9711 1463 9751 1497
rect 9785 1463 9825 1497
rect 9859 1463 9899 1497
rect 9933 1463 9973 1497
rect 10007 1463 10047 1497
rect 10081 1463 10121 1497
rect 10155 1463 10269 1497
rect 10303 1463 10343 1497
rect 10377 1463 10417 1497
rect 10451 1463 10491 1497
rect 10525 1463 10565 1497
rect 10599 1463 10639 1497
rect 10673 1463 10713 1497
rect 10747 1463 10787 1497
rect 10821 1463 10935 1497
rect 10969 1463 11009 1497
rect 11043 1463 11083 1497
rect 11117 1463 11157 1497
rect 11191 1463 11231 1497
rect 11265 1463 11305 1497
rect 11339 1463 11379 1497
rect 11413 1463 11453 1497
rect 11487 1463 11601 1497
rect 11635 1463 11675 1497
rect 11709 1463 11749 1497
rect 11783 1463 11823 1497
rect 11857 1463 11897 1497
rect 11931 1463 11971 1497
rect 12005 1463 12045 1497
rect 12079 1463 12119 1497
rect 12153 1463 12267 1497
rect 12301 1463 12341 1497
rect 12375 1463 12415 1497
rect 12449 1463 12489 1497
rect 12523 1463 12563 1497
rect 12597 1463 12637 1497
rect 12671 1463 12711 1497
rect 12745 1463 12785 1497
rect 12819 1463 12933 1497
rect 12967 1463 13007 1497
rect 13041 1463 13081 1497
rect 13115 1463 13155 1497
rect 13189 1463 13229 1497
rect 13263 1463 13303 1497
rect 13337 1463 13377 1497
rect 13411 1463 13451 1497
rect 13485 1463 13599 1497
rect 13633 1463 13673 1497
rect 13707 1463 13747 1497
rect 13781 1463 13821 1497
rect 13855 1463 13895 1497
rect 13929 1463 13969 1497
rect 14003 1463 14043 1497
rect 14077 1463 14117 1497
rect 14151 1463 14265 1497
rect 14299 1463 14339 1497
rect 14373 1463 14413 1497
rect 14447 1463 14487 1497
rect 14521 1463 14561 1497
rect 14595 1463 14635 1497
rect 14669 1463 14709 1497
rect 14743 1463 14783 1497
rect 14817 1463 14908 1497
rect -34 1446 14908 1463
rect 13275 1059 13321 1065
rect 13675 1059 13721 1065
rect 13939 1059 13985 1065
rect 14343 1059 14389 1065
rect 13269 1025 13281 1059
rect 13315 1025 13681 1059
rect 13715 1025 13727 1059
rect 13933 1025 13945 1059
rect 13979 1025 14349 1059
rect 14383 1025 14395 1059
rect 13275 1019 13321 1025
rect 13675 1019 13721 1025
rect 13939 1019 13985 1025
rect 14343 1019 14389 1025
rect 421 905 467 911
rect 2641 905 2687 911
rect 4713 905 4759 911
rect 6933 905 6979 911
rect 9005 905 9051 911
rect 11225 905 11271 911
rect 12039 905 12085 911
rect 12409 905 12455 911
rect 13001 905 13047 911
rect 13741 905 13787 911
rect 415 871 427 905
rect 461 871 2647 905
rect 2681 904 2693 905
rect 3349 904 4719 905
rect 2681 873 4719 904
rect 2681 871 2693 873
rect 3349 871 4719 873
rect 4753 871 6939 905
rect 6973 871 9011 905
rect 9045 871 11231 905
rect 11265 871 11277 905
rect 12033 871 12045 905
rect 12079 871 12415 905
rect 12449 871 12461 905
rect 12995 871 13007 905
rect 13041 871 13747 905
rect 13781 871 13793 905
rect 421 865 467 871
rect 2641 865 2687 871
rect 4713 865 4759 871
rect 6933 865 6979 871
rect 9005 865 9051 871
rect 11225 865 11271 871
rect 12039 865 12085 871
rect 12409 865 12455 871
rect 13001 865 13047 871
rect 13741 865 13787 871
rect 199 831 245 837
rect 1975 831 2021 837
rect 2789 831 2835 837
rect 3973 831 4019 837
rect 4491 831 4537 837
rect 6267 831 6313 837
rect 7081 831 7127 837
rect 8265 831 8311 837
rect 8783 831 8829 837
rect 10559 831 10605 837
rect 11373 831 11419 837
rect 12557 831 12603 837
rect 13223 831 13269 837
rect 14555 831 14601 837
rect 193 797 205 831
rect 239 797 1981 831
rect 2015 797 2795 831
rect 2829 797 3979 831
rect 4013 797 4025 831
rect 4485 797 4497 831
rect 4531 797 6273 831
rect 6307 797 7087 831
rect 7121 797 8271 831
rect 8305 797 8317 831
rect 8777 797 8789 831
rect 8823 797 10565 831
rect 10599 797 11379 831
rect 11413 797 12563 831
rect 12597 797 12609 831
rect 13217 797 13229 831
rect 13263 797 14561 831
rect 14595 797 14607 831
rect 199 791 245 797
rect 1975 791 2021 797
rect 2789 791 2835 797
rect 3973 791 4019 797
rect 4491 791 4537 797
rect 6267 791 6313 797
rect 7081 791 7127 797
rect 8265 791 8311 797
rect 8783 791 8829 797
rect 10559 791 10605 797
rect 11373 791 11419 797
rect 12557 791 12603 797
rect 13223 791 13269 797
rect 14555 791 14601 797
rect 791 757 837 763
rect 1161 757 1207 763
rect 3159 757 3205 763
rect 3455 757 3501 763
rect 3825 757 3871 763
rect 5083 757 5129 763
rect 5453 757 5499 763
rect 7451 757 7497 763
rect 7747 757 7793 763
rect 8117 757 8163 763
rect 9375 757 9421 763
rect 9745 757 9791 763
rect 11743 757 11789 763
rect 11891 757 11937 763
rect 12705 757 12751 763
rect 13001 757 13047 763
rect 785 723 797 757
rect 831 723 1167 757
rect 1201 723 3165 757
rect 3199 723 3211 757
rect 3449 723 3461 757
rect 3495 723 3831 757
rect 3865 723 3877 757
rect 5077 723 5089 757
rect 5123 723 5459 757
rect 5493 723 7457 757
rect 7491 723 7503 757
rect 7741 723 7753 757
rect 7787 723 8123 757
rect 8157 723 8169 757
rect 9369 723 9381 757
rect 9415 723 9751 757
rect 9785 723 11749 757
rect 11783 723 11795 757
rect 11885 723 11897 757
rect 11931 723 12711 757
rect 12745 723 13007 757
rect 13041 723 13053 757
rect 791 717 837 723
rect 1161 717 1207 723
rect 3159 717 3205 723
rect 3455 717 3501 723
rect 3825 717 3871 723
rect 5083 717 5129 723
rect 5453 717 5499 723
rect 7451 717 7497 723
rect 7747 717 7793 723
rect 8117 717 8163 723
rect 9375 717 9421 723
rect 9745 717 9791 723
rect 11743 717 11789 723
rect 11891 717 11937 723
rect 12705 717 12751 723
rect 13001 717 13047 723
rect 643 683 689 689
rect 1457 683 1503 689
rect 1827 683 1873 689
rect 2123 683 2169 689
rect 2493 683 2539 689
rect 4935 683 4981 689
rect 5749 683 5795 689
rect 6119 683 6165 689
rect 6415 683 6461 689
rect 6785 683 6831 689
rect 9227 683 9273 689
rect 10041 683 10087 689
rect 10411 683 10457 689
rect 10707 683 10753 689
rect 11077 683 11123 689
rect 637 649 649 683
rect 683 649 1463 683
rect 1497 649 1833 683
rect 1867 649 1879 683
rect 2117 649 2129 683
rect 2163 649 2499 683
rect 2533 649 2545 683
rect 4929 649 4941 683
rect 4975 649 5755 683
rect 5789 649 6125 683
rect 6159 649 6171 683
rect 6409 649 6421 683
rect 6455 649 6791 683
rect 6825 649 6837 683
rect 9221 649 9233 683
rect 9267 649 10047 683
rect 10081 649 10417 683
rect 10451 649 10463 683
rect 10701 649 10713 683
rect 10747 649 11083 683
rect 11117 649 11129 683
rect 643 643 689 649
rect 1457 643 1503 649
rect 1827 643 1873 649
rect 2123 643 2169 649
rect 2493 643 2539 649
rect 4935 643 4981 649
rect 5749 643 5795 649
rect 6119 643 6165 649
rect 6415 643 6461 649
rect 6785 643 6831 649
rect 9227 643 9273 649
rect 10041 643 10087 649
rect 10411 643 10457 649
rect 10707 643 10753 649
rect 11077 643 11123 649
rect 3307 609 3353 615
rect 4121 609 4167 615
rect 14037 609 14083 615
rect 3301 575 3313 609
rect 3347 575 4127 609
rect 4161 575 14043 609
rect 14077 575 14089 609
rect 3307 569 3353 575
rect 4121 569 4167 575
rect 14037 569 14083 575
rect 1309 535 1355 541
rect 5601 535 5647 541
rect 9893 535 9939 541
rect 1303 501 1315 535
rect 1349 501 5607 535
rect 5641 501 9899 535
rect 9933 501 9945 535
rect 1309 495 1355 501
rect 5601 495 5647 501
rect 9893 495 9939 501
rect 7599 461 7645 467
rect 8413 461 8459 467
rect 13223 461 13269 467
rect 7593 427 7605 461
rect 7639 427 8419 461
rect 8453 427 13229 461
rect 13263 427 13275 461
rect 14037 433 14083 439
rect 14333 433 14379 439
rect 7599 421 7645 427
rect 8413 421 8459 427
rect 13223 421 13269 427
rect 14031 399 14043 433
rect 14077 399 14339 433
rect 14373 399 14385 433
rect 14037 393 14083 399
rect 14333 393 14379 399
rect 13283 253 13329 259
rect 13949 253 13995 259
rect 14615 253 14661 259
rect 13277 219 13289 253
rect 13323 219 13955 253
rect 13989 219 14621 253
rect 14655 219 14667 253
rect 13283 213 13329 219
rect 13949 213 13995 219
rect 14615 213 14661 219
rect -34 17 14908 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5163 17
rect 5197 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5533 17
rect 5567 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5755 17
rect 5789 -17 5829 17
rect 5863 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6125 17
rect 6159 -17 6199 17
rect 6233 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6495 17
rect 6529 -17 6643 17
rect 6677 -17 6717 17
rect 6751 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7087 17
rect 7121 -17 7161 17
rect 7195 -17 7309 17
rect 7343 -17 7383 17
rect 7417 -17 7457 17
rect 7491 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7679 17
rect 7713 -17 7753 17
rect 7787 -17 7827 17
rect 7861 -17 7975 17
rect 8009 -17 8049 17
rect 8083 -17 8123 17
rect 8157 -17 8197 17
rect 8231 -17 8271 17
rect 8305 -17 8345 17
rect 8379 -17 8419 17
rect 8453 -17 8493 17
rect 8527 -17 8641 17
rect 8675 -17 8715 17
rect 8749 -17 8789 17
rect 8823 -17 8863 17
rect 8897 -17 8937 17
rect 8971 -17 9011 17
rect 9045 -17 9085 17
rect 9119 -17 9159 17
rect 9193 -17 9233 17
rect 9267 -17 9307 17
rect 9341 -17 9381 17
rect 9415 -17 9455 17
rect 9489 -17 9603 17
rect 9637 -17 9677 17
rect 9711 -17 9751 17
rect 9785 -17 9825 17
rect 9859 -17 9899 17
rect 9933 -17 9973 17
rect 10007 -17 10047 17
rect 10081 -17 10121 17
rect 10155 -17 10269 17
rect 10303 -17 10343 17
rect 10377 -17 10417 17
rect 10451 -17 10491 17
rect 10525 -17 10565 17
rect 10599 -17 10639 17
rect 10673 -17 10713 17
rect 10747 -17 10787 17
rect 10821 -17 10935 17
rect 10969 -17 11009 17
rect 11043 -17 11083 17
rect 11117 -17 11157 17
rect 11191 -17 11231 17
rect 11265 -17 11305 17
rect 11339 -17 11379 17
rect 11413 -17 11453 17
rect 11487 -17 11601 17
rect 11635 -17 11675 17
rect 11709 -17 11749 17
rect 11783 -17 11823 17
rect 11857 -17 11897 17
rect 11931 -17 11971 17
rect 12005 -17 12045 17
rect 12079 -17 12119 17
rect 12153 -17 12267 17
rect 12301 -17 12341 17
rect 12375 -17 12415 17
rect 12449 -17 12489 17
rect 12523 -17 12563 17
rect 12597 -17 12637 17
rect 12671 -17 12711 17
rect 12745 -17 12785 17
rect 12819 -17 12933 17
rect 12967 -17 13007 17
rect 13041 -17 13081 17
rect 13115 -17 13155 17
rect 13189 -17 13229 17
rect 13263 -17 13303 17
rect 13337 -17 13377 17
rect 13411 -17 13451 17
rect 13485 -17 13599 17
rect 13633 -17 13673 17
rect 13707 -17 13747 17
rect 13781 -17 13821 17
rect 13855 -17 13895 17
rect 13929 -17 13969 17
rect 14003 -17 14043 17
rect 14077 -17 14117 17
rect 14151 -17 14265 17
rect 14299 -17 14339 17
rect 14373 -17 14413 17
rect 14447 -17 14487 17
rect 14521 -17 14561 17
rect 14595 -17 14635 17
rect 14669 -17 14709 17
rect 14743 -17 14783 17
rect 14817 -17 14908 17
rect -34 -34 14908 -17
<< labels >>
rlabel locali 14709 723 14743 757 1 QN
port 1 nsew signal output
rlabel locali 14709 797 14743 831 1 QN
port 1 nsew signal output
rlabel locali 14709 871 14743 905 1 QN
port 1 nsew signal output
rlabel locali 14709 945 14743 979 1 QN
port 1 nsew signal output
rlabel locali 14709 649 14743 683 1 QN
port 1 nsew signal output
rlabel locali 14709 575 14743 609 1 QN
port 1 nsew signal output
rlabel locali 14709 501 14743 535 1 QN
port 1 nsew signal output
rlabel locali 14709 427 14743 461 1 QN
port 1 nsew signal output
rlabel locali 1315 501 1349 535 1 D
port 2 nsew signal input
rlabel locali 5607 501 5641 535 1 D
port 2 nsew signal input
rlabel locali 9899 501 9933 535 1 D
port 2 nsew signal input
rlabel locali 1315 575 1349 609 1 D
port 2 nsew signal input
rlabel locali 427 871 461 905 1 CLK
port 3 nsew signal input
rlabel locali 427 723 461 757 1 CLK
port 3 nsew signal input
rlabel locali 427 649 461 683 1 CLK
port 3 nsew signal input
rlabel locali 427 575 461 609 1 CLK
port 3 nsew signal input
rlabel locali 427 501 461 535 1 CLK
port 3 nsew signal input
rlabel locali 4719 649 4753 683 1 CLK
port 3 nsew signal input
rlabel locali 4719 723 4753 757 1 CLK
port 3 nsew signal input
rlabel locali 2647 649 2681 683 1 CLK
port 3 nsew signal input
rlabel locali 2647 575 2681 609 1 CLK
port 3 nsew signal input
rlabel locali 6939 649 6973 683 1 CLK
port 3 nsew signal input
rlabel locali 9011 649 9045 683 1 CLK
port 3 nsew signal input
rlabel locali 9011 723 9045 757 1 CLK
port 3 nsew signal input
rlabel locali 11231 649 11265 683 1 CLK
port 3 nsew signal input
rlabel locali 2647 871 2681 905 1 CLK
port 3 nsew signal input
rlabel locali 4719 871 4753 905 1 CLK
port 3 nsew signal input
rlabel locali 6939 871 6973 905 1 CLK
port 3 nsew signal input
rlabel locali 9011 871 9045 905 1 CLK
port 3 nsew signal input
rlabel locali 11231 501 11265 535 1 CLK
port 3 nsew signal input
rlabel locali 11231 871 11265 905 1 CLK
port 3 nsew signal input
rlabel metal1 -34 1446 14908 1514 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 -34 -34 14908 34 1 GND
port 5 nsew power bidirectional abutment
<< end >>
