* SPICE3 file created from OR2X1.ext - technology: sky130A

.subckt OR2X1 Y A B VDD GND
M1000 a_198_209.t3 B.t0 a_131_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 Y.t0 a_198_209.t5 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_131_1051.t0 A.t1 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_131_1051.t2 B.t2 a_198_209.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VDD.t2 a_198_209.t6 Y.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y a_198_209.t4 GND.t2 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1006 VDD.t1 A.t2 a_131_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VDD A 0.08fF
C1 Y VDD 0.76fF
C2 B A 0.26fF
C3 B VDD 0.07fF
R0 a_198_209.n2 a_198_209.t6 512.525
R1 a_198_209.n2 a_198_209.t5 371.139
R2 a_198_209.n3 a_198_209.t4 210.434
R3 a_198_209.n4 a_198_209.n1 191.889
R4 a_198_209.n3 a_198_209.n2 173.2
R5 a_198_209.n4 a_198_209.n3 153.043
R6 a_198_209.n9 a_198_209.n4 135.634
R7 a_198_209.n9 a_198_209.n8 118.016
R8 a_198_209.n12 a_198_209.n0 55.263
R9 a_198_209.n11 a_198_209.n9 48.405
R10 a_198_209.n8 a_198_209.n7 30
R11 a_198_209.n11 a_198_209.n10 30
R12 a_198_209.n12 a_198_209.n11 25.263
R13 a_198_209.n6 a_198_209.n5 24.383
R14 a_198_209.n8 a_198_209.n6 23.684
R15 a_198_209.n1 a_198_209.t2 14.282
R16 a_198_209.n1 a_198_209.t3 14.282
R17 GND.n32 GND.n31 219.745
R18 GND.n32 GND.n30 85.529
R19 GND.n9 GND.n1 76.145
R20 GND.n39 GND.n38 76
R21 GND.n9 GND.n8 76
R22 GND.n17 GND.n16 76
R23 GND.n26 GND.n25 76
R24 GND.n29 GND.n28 76
R25 GND.n36 GND.n35 76
R26 GND.n73 GND.n72 76
R27 GND.n66 GND.n65 76
R28 GND.n60 GND.n59 76
R29 GND.n54 GND.n53 76
R30 GND.n51 GND.n50 76
R31 GND.n46 GND.n45 76
R32 GND.n22 GND.t2 39.412
R33 GND.n5 GND.n4 35.01
R34 GND.n6 GND.n5 19.735
R35 GND.n14 GND.n13 19.735
R36 GND.n24 GND.n23 19.735
R37 GND.n48 GND.n47 19.735
R38 GND.n58 GND.n57 19.735
R39 GND.n64 GND.n63 19.735
R40 GND.n70 GND.n69 19.735
R41 GND.n44 GND.n43 19.735
R42 GND.n63 GND.t1 19.724
R43 GND.n47 GND.t0 19.724
R44 GND.n5 GND.n3 19.017
R45 GND.n22 GND.n21 17.185
R46 GND.n35 GND.n33 14.167
R47 GND.n45 GND.n40 13.653
R48 GND.n50 GND.n49 13.653
R49 GND.n53 GND.n52 13.653
R50 GND.n59 GND.n55 13.653
R51 GND.n65 GND.n61 13.653
R52 GND.n72 GND.n71 13.653
R53 GND.n35 GND.n34 13.653
R54 GND.n28 GND.n27 13.653
R55 GND.n25 GND.n18 13.653
R56 GND.n16 GND.n15 13.653
R57 GND.n8 GND.n7 13.653
R58 GND.n43 GND.n42 12.837
R59 GND.n69 GND.n68 11.605
R60 GND.n68 GND.n67 9.809
R61 GND.n59 GND.n58 8.854
R62 GND.n42 GND.n41 7.566
R63 GND.n3 GND.n2 7.5
R64 GND.n12 GND.n11 7.5
R65 GND.n33 GND.n32 7.312
R66 GND.t1 GND.n62 7.04
R67 GND.n23 GND.n22 6.139
R68 GND.n57 GND.n56 5.774
R69 GND.n20 GND.n19 4.551
R70 GND.n8 GND.n6 3.935
R71 GND.n65 GND.n64 3.935
R72 GND.n50 GND.n48 3.935
R73 GND.n25 GND.n24 3.541
R74 GND.t2 GND.n20 2.238
R75 GND.n11 GND.n10 1.935
R76 GND.n72 GND.n70 0.983
R77 GND.n45 GND.n44 0.983
R78 GND.n1 GND.n0 0.596
R79 GND.n38 GND.n37 0.596
R80 GND.n13 GND.n12 0.358
R81 GND.n36 GND.n29 0.29
R82 GND.n39 GND 0.207
R83 GND.n16 GND.n14 0.196
R84 GND.n60 GND.n54 0.181
R85 GND.n17 GND.n9 0.157
R86 GND.n26 GND.n17 0.157
R87 GND.n29 GND.n26 0.145
R88 GND.n73 GND.n66 0.145
R89 GND.n66 GND.n60 0.145
R90 GND.n54 GND.n51 0.145
R91 GND.n51 GND.n46 0.145
R92 GND.n46 GND.n39 0.145
R93 GND GND.n36 0.078
R94 GND GND.n73 0.066
R95 Y.n2 Y.n1 200.754
R96 Y.n2 Y.n0 184.007
R97 Y Y.n2 76
R98 Y.n0 Y.t1 14.282
R99 Y.n0 Y.t0 14.282
R100 B.n0 B.t2 470.752
R101 B.n0 B.t0 384.527
R102 B.n1 B.t1 241.172
R103 B.n1 B.n0 110.173
R104 B B.n1 76
R105 a_131_1051.t2 a_131_1051.n0 101.663
R106 a_131_1051.n0 a_131_1051.t1 101.661
R107 a_131_1051.n0 a_131_1051.t3 14.294
R108 a_131_1051.n0 a_131_1051.t0 14.282
R109 VDD.n68 VDD.n66 144.705
R110 VDD.n26 VDD.n25 77.792
R111 VDD.n35 VDD.n34 77.792
R112 VDD.n29 VDD.n23 76.145
R113 VDD.n29 VDD.n28 76
R114 VDD.n33 VDD.n32 76
R115 VDD.n39 VDD.n38 76
R116 VDD.n43 VDD.n42 76
R117 VDD.n70 VDD.n69 76
R118 VDD.n121 VDD.n120 76
R119 VDD.n117 VDD.n116 76
R120 VDD.n113 VDD.n112 76
R121 VDD.n109 VDD.n108 76
R122 VDD.n104 VDD.n103 76
R123 VDD.n97 VDD.n96 76
R124 VDD.n93 VDD.n92 76
R125 VDD.n37 VDD.t3 55.106
R126 VDD.n24 VDD.t2 55.106
R127 VDD.n99 VDD.n98 41.183
R128 VDD.n59 VDD.n58 36.774
R129 VDD.n101 VDD.n100 32.032
R130 VDD.n92 VDD.n89 21.841
R131 VDD.n23 VDD.n20 21.841
R132 VDD.n98 VDD.t0 14.282
R133 VDD.n98 VDD.t1 14.282
R134 VDD.n89 VDD.n72 14.167
R135 VDD.n72 VDD.n71 14.167
R136 VDD.n64 VDD.n45 14.167
R137 VDD.n45 VDD.n44 14.167
R138 VDD.n20 VDD.n19 14.167
R139 VDD.n19 VDD.n17 14.167
R140 VDD.n69 VDD.n65 14.167
R141 VDD.n23 VDD.n22 13.653
R142 VDD.n22 VDD.n21 13.653
R143 VDD.n28 VDD.n27 13.653
R144 VDD.n27 VDD.n26 13.653
R145 VDD.n32 VDD.n31 13.653
R146 VDD.n31 VDD.n30 13.653
R147 VDD.n38 VDD.n36 13.653
R148 VDD.n36 VDD.n35 13.653
R149 VDD.n42 VDD.n41 13.653
R150 VDD.n41 VDD.n40 13.653
R151 VDD.n69 VDD.n68 13.653
R152 VDD.n68 VDD.n67 13.653
R153 VDD.n120 VDD.n119 13.653
R154 VDD.n119 VDD.n118 13.653
R155 VDD.n116 VDD.n115 13.653
R156 VDD.n115 VDD.n114 13.653
R157 VDD.n112 VDD.n111 13.653
R158 VDD.n111 VDD.n110 13.653
R159 VDD.n108 VDD.n107 13.653
R160 VDD.n107 VDD.n106 13.653
R161 VDD.n103 VDD.n102 13.653
R162 VDD.n102 VDD.n101 13.653
R163 VDD.n96 VDD.n95 13.653
R164 VDD.n95 VDD.n94 13.653
R165 VDD.n92 VDD.n91 13.653
R166 VDD.n91 VDD.n90 13.653
R167 VDD.n4 VDD.n2 12.915
R168 VDD.n4 VDD.n3 12.66
R169 VDD.n13 VDD.n12 12.343
R170 VDD.n10 VDD.n9 12.343
R171 VDD.n7 VDD.n6 12.343
R172 VDD.n65 VDD.n64 7.674
R173 VDD.n49 VDD.n48 7.5
R174 VDD.n52 VDD.n51 7.5
R175 VDD.n54 VDD.n53 7.5
R176 VDD.n57 VDD.n56 7.5
R177 VDD.n64 VDD.n63 7.5
R178 VDD.n84 VDD.n83 7.5
R179 VDD.n78 VDD.n77 7.5
R180 VDD.n80 VDD.n79 7.5
R181 VDD.n86 VDD.n76 7.5
R182 VDD.n86 VDD.n74 7.5
R183 VDD.n89 VDD.n88 7.5
R184 VDD.n20 VDD.n16 7.5
R185 VDD.n2 VDD.n1 7.5
R186 VDD.n6 VDD.n5 7.5
R187 VDD.n9 VDD.n8 7.5
R188 VDD.n19 VDD.n18 7.5
R189 VDD.n14 VDD.n0 7.5
R190 VDD.n87 VDD.n73 6.772
R191 VDD.n85 VDD.n82 6.772
R192 VDD.n81 VDD.n78 6.772
R193 VDD.n81 VDD.n80 6.772
R194 VDD.n85 VDD.n84 6.772
R195 VDD.n88 VDD.n87 6.772
R196 VDD.n63 VDD.n62 6.772
R197 VDD.n50 VDD.n47 6.772
R198 VDD.n55 VDD.n52 6.772
R199 VDD.n60 VDD.n57 6.772
R200 VDD.n60 VDD.n59 6.772
R201 VDD.n55 VDD.n54 6.772
R202 VDD.n50 VDD.n49 6.772
R203 VDD.n62 VDD.n46 6.772
R204 VDD.n16 VDD.n15 6.458
R205 VDD.n76 VDD.n75 6.202
R206 VDD.n103 VDD.n99 5.903
R207 VDD.n106 VDD.n105 4.576
R208 VDD.n28 VDD.n24 1.967
R209 VDD.n38 VDD.n37 1.967
R210 VDD.n14 VDD.n7 1.329
R211 VDD.n14 VDD.n10 1.329
R212 VDD.n14 VDD.n11 1.329
R213 VDD.n14 VDD.n13 1.329
R214 VDD.n15 VDD.n14 0.696
R215 VDD.n14 VDD.n4 0.696
R216 VDD.n86 VDD.n85 0.365
R217 VDD.n86 VDD.n81 0.365
R218 VDD.n87 VDD.n86 0.365
R219 VDD.n61 VDD.n60 0.365
R220 VDD.n61 VDD.n55 0.365
R221 VDD.n61 VDD.n50 0.365
R222 VDD.n62 VDD.n61 0.365
R223 VDD.n70 VDD.n43 0.29
R224 VDD.n93 VDD 0.207
R225 VDD.n113 VDD.n109 0.181
R226 VDD.n33 VDD.n29 0.157
R227 VDD.n39 VDD.n33 0.157
R228 VDD.n43 VDD.n39 0.145
R229 VDD.n121 VDD.n117 0.145
R230 VDD.n117 VDD.n113 0.145
R231 VDD.n109 VDD.n104 0.145
R232 VDD.n104 VDD.n97 0.145
R233 VDD.n97 VDD.n93 0.145
R234 VDD VDD.n70 0.078
R235 VDD VDD.n121 0.066
R236 A.n0 A.t1 486.819
R237 A.n0 A.t2 384.527
R238 A.n1 A.t0 303.607
R239 A.n1 A.n0 79.994
R240 A A.n1 76
C4 VDD GND 4.98fF
C5 VDD.n0 GND 0.11fF
C6 VDD.n1 GND 0.02fF
C7 VDD.n2 GND 0.02fF
C8 VDD.n3 GND 0.04fF
C9 VDD.n4 GND 0.01fF
C10 VDD.n5 GND 0.02fF
C11 VDD.n6 GND 0.02fF
C12 VDD.n8 GND 0.02fF
C13 VDD.n9 GND 0.02fF
C14 VDD.n12 GND 0.02fF
C15 VDD.n14 GND 0.42fF
C16 VDD.n16 GND 0.03fF
C17 VDD.n17 GND 0.02fF
C18 VDD.n18 GND 0.02fF
C19 VDD.n19 GND 0.02fF
C20 VDD.n20 GND 0.03fF
C21 VDD.n21 GND 0.25fF
C22 VDD.n22 GND 0.02fF
C23 VDD.n23 GND 0.03fF
C24 VDD.n24 GND 0.05fF
C25 VDD.n25 GND 0.14fF
C26 VDD.n26 GND 0.19fF
C27 VDD.n27 GND 0.01fF
C28 VDD.n28 GND 0.01fF
C29 VDD.n29 GND 0.06fF
C30 VDD.n30 GND 0.15fF
C31 VDD.n31 GND 0.01fF
C32 VDD.n32 GND 0.02fF
C33 VDD.n33 GND 0.02fF
C34 VDD.n34 GND 0.14fF
C35 VDD.n35 GND 0.19fF
C36 VDD.n36 GND 0.01fF
C37 VDD.n37 GND 0.06fF
C38 VDD.n38 GND 0.01fF
C39 VDD.n39 GND 0.02fF
C40 VDD.n40 GND 0.25fF
C41 VDD.n41 GND 0.01fF
C42 VDD.n42 GND 0.02fF
C43 VDD.n43 GND 0.03fF
C44 VDD.n44 GND 0.02fF
C45 VDD.n45 GND 0.02fF
C46 VDD.n46 GND 0.02fF
C47 VDD.n47 GND 0.02fF
C48 VDD.n48 GND 0.02fF
C49 VDD.n49 GND 0.02fF
C50 VDD.n51 GND 0.02fF
C51 VDD.n52 GND 0.02fF
C52 VDD.n53 GND 0.02fF
C53 VDD.n54 GND 0.02fF
C54 VDD.n56 GND 0.03fF
C55 VDD.n57 GND 0.02fF
C56 VDD.n58 GND 0.17fF
C57 VDD.n59 GND 0.04fF
C58 VDD.n61 GND 0.25fF
C59 VDD.n63 GND 0.02fF
C60 VDD.n64 GND 0.02fF
C61 VDD.n65 GND 0.03fF
C62 VDD.n66 GND 0.02fF
C63 VDD.n67 GND 0.25fF
C64 VDD.n68 GND 0.01fF
C65 VDD.n69 GND 0.02fF
C66 VDD.n70 GND 0.03fF
C67 VDD.n71 GND 0.02fF
C68 VDD.n72 GND 0.02fF
C69 VDD.n73 GND 0.02fF
C70 VDD.n74 GND 0.14fF
C71 VDD.n75 GND 0.03fF
C72 VDD.n76 GND 0.02fF
C73 VDD.n77 GND 0.02fF
C74 VDD.n78 GND 0.02fF
C75 VDD.n79 GND 0.02fF
C76 VDD.n80 GND 0.02fF
C77 VDD.n82 GND 0.02fF
C78 VDD.n83 GND 0.02fF
C79 VDD.n84 GND 0.02fF
C80 VDD.n86 GND 0.42fF
C81 VDD.n88 GND 0.03fF
C82 VDD.n89 GND 0.03fF
C83 VDD.n90 GND 0.25fF
C84 VDD.n91 GND 0.02fF
C85 VDD.n92 GND 0.03fF
C86 VDD.n93 GND 0.03fF
C87 VDD.n94 GND 0.23fF
C88 VDD.n95 GND 0.01fF
C89 VDD.n96 GND 0.02fF
C90 VDD.n97 GND 0.02fF
C91 VDD.n98 GND 0.10fF
C92 VDD.n99 GND 0.02fF
C93 VDD.n100 GND 0.13fF
C94 VDD.n101 GND 0.15fF
C95 VDD.n102 GND 0.01fF
C96 VDD.n103 GND 0.01fF
C97 VDD.n104 GND 0.02fF
C98 VDD.n105 GND 0.16fF
C99 VDD.n106 GND 0.13fF
C100 VDD.n107 GND 0.01fF
C101 VDD.n108 GND 0.02fF
C102 VDD.n109 GND 0.02fF
C103 VDD.n110 GND 0.28fF
C104 VDD.n111 GND 0.01fF
C105 VDD.n112 GND 0.02fF
C106 VDD.n113 GND 0.02fF
C107 VDD.n114 GND 0.25fF
C108 VDD.n115 GND 0.01fF
C109 VDD.n116 GND 0.02fF
C110 VDD.n117 GND 0.02fF
C111 VDD.n118 GND 0.25fF
C112 VDD.n119 GND 0.01fF
C113 VDD.n120 GND 0.02fF
C114 VDD.n121 GND 0.02fF
C115 a_131_1051.n0 GND 0.52fF
C116 Y.n0 GND 0.82fF
C117 Y.n1 GND 0.38fF
C118 Y.n2 GND 0.51fF
C119 a_198_209.n0 GND 0.04fF
C120 a_198_209.n1 GND 0.58fF
C121 a_198_209.n2 GND 0.31fF
C122 a_198_209.n3 GND 0.48fF
C123 a_198_209.n4 GND 0.44fF
C124 a_198_209.n5 GND 0.03fF
C125 a_198_209.n6 GND 0.04fF
C126 a_198_209.n7 GND 0.03fF
C127 a_198_209.n8 GND 0.15fF
C128 a_198_209.n9 GND 0.30fF
C129 a_198_209.n10 GND 0.03fF
C130 a_198_209.n11 GND 0.08fF
C131 a_198_209.n12 GND 0.04fF
.ends
