* SPICE3 file created from AOA4X1.ext - technology: sky130A

.subckt AOA4X1 Y A B C D VDD GND
X0 Y aoa4x1_pcell_0/m1_1869_501# GND GND nshort w=3 l=0.15
X1 VDD aoa4x1_pcell_0/m1_1869_501# Y VDD pshort w=2 l=0.15
X2 VDD aoa4x1_pcell_0/aoai4x1_pcell_0/m1_537_501# aoa4x1_pcell_0/aoai4x1_pcell_0/nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X3 aoa4x1_pcell_0/aoai4x1_pcell_0/m1_1203_501# C aoa4x1_pcell_0/aoai4x1_pcell_0/nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X4 aoa4x1_pcell_0/aoai4x1_pcell_0/m1_1203_501# aoa4x1_pcell_0/aoai4x1_pcell_0/m1_537_501# GND GND nshort w=3 l=0.15
X5 aoa4x1_pcell_0/aoai4x1_pcell_0/m1_1203_501# C GND GND nshort w=3 l=0.15
X6 GND A aoa4x1_pcell_0/aoai4x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X7 aoa4x1_pcell_0/aoai4x1_pcell_0/m1_537_501# B aoa4x1_pcell_0/aoai4x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X8 VDD A aoa4x1_pcell_0/aoai4x1_pcell_0/m1_537_501# VDD pshort w=2 l=0.15
X9 VDD B aoa4x1_pcell_0/aoai4x1_pcell_0/m1_537_501# VDD pshort w=2 l=0.15
X10 GND aoa4x1_pcell_0/aoai4x1_pcell_0/m1_1203_501# aoa4x1_pcell_0/aoai4x1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X11 aoa4x1_pcell_0/m1_1869_501# D aoa4x1_pcell_0/aoai4x1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X12 VDD aoa4x1_pcell_0/aoai4x1_pcell_0/m1_1203_501# aoa4x1_pcell_0/m1_1869_501# VDD pshort w=2 l=0.15
X13 VDD D aoa4x1_pcell_0/m1_1869_501# VDD pshort w=2 l=0.15
C0 VDD GND 3.00fF
.ends
