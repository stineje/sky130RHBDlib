* SPICE3 file created from NOR2X1.ext - technology: sky130A

.subckt NOR2X1 Y A B VDD GND
X0 Y A GND GND nshort w=3 l=0.15
X1 a_131_1005 A VDD VDD pshort w=2 l=0.15 M=2
X2 a_131_1005 B Y VDD pshort w=2 l=0.15 M=2
X3 Y B GND GND nshort w=3 l=0.15
.ends
