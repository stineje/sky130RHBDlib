magic
tech sky130A
magscale 1 2
timestamp 1669507662
<< nwell >>
rect -87 786 2085 1550
<< pwell >>
rect -34 -34 2032 544
<< nmos >>
rect 168 288 198 349
tri 198 288 214 304 sw
rect 362 296 392 349
tri 392 296 408 312 sw
rect 168 258 274 288
tri 274 258 304 288 sw
rect 362 266 468 296
tri 468 266 498 296 sw
rect 168 157 198 258
tri 198 242 214 258 nw
tri 258 242 274 258 ne
tri 198 157 214 173 sw
tri 258 157 274 173 se
rect 274 157 304 258
rect 362 165 392 266
tri 392 250 408 266 nw
tri 452 250 468 266 ne
tri 392 165 408 181 sw
tri 452 165 468 181 se
rect 468 165 498 266
tri 168 127 198 157 ne
rect 198 127 274 157
tri 274 127 304 157 nw
tri 362 135 392 165 ne
rect 392 135 468 165
tri 468 135 498 165 nw
rect 834 288 864 349
tri 864 288 880 304 sw
tri 1118 296 1134 312 se
rect 1134 296 1164 349
rect 834 258 940 288
tri 940 258 970 288 sw
tri 1028 266 1058 296 se
rect 1058 266 1164 296
rect 834 157 864 258
tri 864 242 880 258 nw
tri 924 242 940 258 ne
tri 864 157 880 173 sw
tri 924 157 940 173 se
rect 940 157 970 258
rect 1028 165 1058 266
tri 1058 250 1074 266 nw
tri 1118 250 1134 266 ne
tri 1058 165 1074 181 sw
tri 1118 165 1134 181 se
rect 1134 165 1164 266
tri 834 127 864 157 ne
rect 864 127 940 157
tri 940 127 970 157 nw
tri 1028 135 1058 165 ne
rect 1058 135 1134 165
tri 1134 135 1164 165 nw
rect 1500 288 1530 349
tri 1530 288 1546 304 sw
rect 1694 296 1724 349
tri 1724 296 1740 312 sw
rect 1500 258 1606 288
tri 1606 258 1636 288 sw
rect 1694 266 1800 296
tri 1800 266 1830 296 sw
rect 1500 157 1530 258
tri 1530 242 1546 258 nw
tri 1590 242 1606 258 ne
tri 1530 157 1546 173 sw
tri 1590 157 1606 173 se
rect 1606 157 1636 258
rect 1694 251 1725 266
tri 1725 251 1740 266 nw
tri 1784 251 1799 266 ne
rect 1799 251 1830 266
rect 1694 165 1724 251
tri 1724 165 1740 181 sw
tri 1784 165 1800 181 se
rect 1800 165 1830 251
tri 1500 127 1530 157 ne
rect 1530 127 1606 157
tri 1606 127 1636 157 nw
tri 1694 135 1724 165 ne
rect 1724 135 1800 165
tri 1800 135 1830 165 nw
<< pmos >>
rect 187 1005 217 1405
rect 275 1005 305 1405
rect 363 1005 393 1405
rect 451 1005 481 1405
rect 851 1005 881 1405
rect 939 1005 969 1405
rect 1027 1005 1057 1405
rect 1115 1005 1145 1405
rect 1519 1005 1549 1405
rect 1607 1005 1637 1405
rect 1695 1005 1725 1405
rect 1783 1005 1813 1405
<< ndiff >>
rect 112 333 168 349
rect 112 299 122 333
rect 156 299 168 333
rect 112 261 168 299
rect 198 333 362 349
rect 198 304 219 333
tri 198 288 214 304 ne
rect 214 299 219 304
rect 253 299 316 333
rect 350 299 362 333
rect 214 288 362 299
rect 392 333 552 349
rect 392 312 510 333
tri 392 296 408 312 ne
rect 408 299 510 312
rect 544 299 552 333
rect 408 296 552 299
rect 112 227 122 261
rect 156 227 168 261
tri 274 258 304 288 ne
rect 304 261 362 288
tri 468 266 498 296 ne
rect 112 193 168 227
rect 112 159 122 193
rect 156 159 168 193
rect 112 127 168 159
tri 198 242 214 258 se
rect 214 242 258 258
tri 258 242 274 258 sw
rect 198 208 274 242
rect 198 174 219 208
rect 253 174 274 208
rect 198 173 274 174
tri 198 157 214 173 ne
rect 214 157 258 173
tri 258 157 274 173 nw
rect 304 227 316 261
rect 350 227 362 261
rect 304 193 362 227
rect 304 159 316 193
rect 350 159 362 193
tri 392 250 408 266 se
rect 408 250 452 266
tri 452 250 468 266 sw
rect 392 217 468 250
rect 392 183 412 217
rect 446 183 468 217
rect 392 181 468 183
tri 392 165 408 181 ne
rect 408 165 452 181
tri 452 165 468 181 nw
rect 498 261 552 296
rect 498 227 510 261
rect 544 227 552 261
rect 498 193 552 227
tri 168 127 198 157 sw
tri 274 127 304 157 se
rect 304 135 362 159
tri 362 135 392 165 sw
tri 468 135 498 165 se
rect 498 159 510 193
rect 544 159 552 193
rect 498 135 552 159
rect 304 127 552 135
rect 112 123 552 127
rect 112 89 122 123
rect 156 89 316 123
rect 350 89 412 123
rect 446 89 510 123
rect 544 89 552 123
rect 112 73 552 89
rect 778 333 834 349
rect 778 299 788 333
rect 822 299 834 333
rect 778 261 834 299
rect 864 333 1134 349
rect 864 304 885 333
tri 864 288 880 304 ne
rect 880 299 885 304
rect 919 299 982 333
rect 1016 312 1134 333
rect 1016 299 1118 312
rect 880 296 1118 299
tri 1118 296 1134 312 nw
rect 1164 333 1220 349
rect 1164 299 1176 333
rect 1210 299 1220 333
rect 880 288 1028 296
rect 778 227 788 261
rect 822 227 834 261
tri 940 258 970 288 ne
rect 970 261 1028 288
tri 1028 266 1058 296 nw
rect 778 193 834 227
rect 778 159 788 193
rect 822 159 834 193
rect 778 127 834 159
tri 864 242 880 258 se
rect 880 242 924 258
tri 924 242 940 258 sw
rect 864 208 940 242
rect 864 174 885 208
rect 919 174 940 208
rect 864 173 940 174
tri 864 157 880 173 ne
rect 880 157 924 173
tri 924 157 940 173 nw
rect 970 227 982 261
rect 1016 227 1028 261
rect 970 193 1028 227
rect 970 159 982 193
rect 1016 159 1028 193
tri 1058 250 1074 266 se
rect 1074 250 1118 266
tri 1118 250 1134 266 sw
rect 1058 217 1134 250
rect 1058 183 1079 217
rect 1113 183 1134 217
rect 1058 181 1134 183
tri 1058 165 1074 181 ne
rect 1074 165 1118 181
tri 1118 165 1134 181 nw
rect 1164 261 1220 299
rect 1164 227 1176 261
rect 1210 227 1220 261
rect 1164 193 1220 227
tri 834 127 864 157 sw
tri 940 127 970 157 se
rect 970 135 1028 159
tri 1028 135 1058 165 sw
tri 1134 135 1164 165 se
rect 1164 159 1176 193
rect 1210 159 1220 193
rect 1164 135 1220 159
rect 970 127 1220 135
rect 778 123 1220 127
rect 778 89 788 123
rect 822 89 982 123
rect 1016 89 1079 123
rect 1113 89 1176 123
rect 1210 89 1220 123
rect 778 73 1220 89
rect 1444 333 1500 349
rect 1444 299 1454 333
rect 1488 299 1500 333
rect 1444 261 1500 299
rect 1530 333 1694 349
rect 1530 304 1551 333
tri 1530 288 1546 304 ne
rect 1546 299 1551 304
rect 1585 299 1648 333
rect 1682 299 1694 333
rect 1546 288 1694 299
rect 1724 312 1886 349
tri 1724 296 1740 312 ne
rect 1740 296 1886 312
rect 1444 227 1454 261
rect 1488 227 1500 261
tri 1606 258 1636 288 ne
rect 1636 261 1694 288
tri 1800 266 1830 296 ne
rect 1444 193 1500 227
rect 1444 159 1454 193
rect 1488 159 1500 193
rect 1444 127 1500 159
tri 1530 242 1546 258 se
rect 1546 242 1590 258
tri 1590 242 1606 258 sw
rect 1530 208 1606 242
rect 1530 174 1551 208
rect 1585 174 1606 208
rect 1530 173 1606 174
tri 1530 157 1546 173 ne
rect 1546 157 1590 173
tri 1590 157 1606 173 nw
rect 1636 227 1648 261
rect 1682 227 1694 261
tri 1725 251 1740 266 se
rect 1740 251 1784 266
tri 1784 251 1799 266 sw
rect 1830 261 1886 296
rect 1636 193 1694 227
rect 1636 159 1648 193
rect 1682 159 1694 193
rect 1724 217 1800 251
rect 1724 183 1745 217
rect 1779 183 1800 217
rect 1724 181 1800 183
tri 1724 165 1740 181 ne
rect 1740 165 1784 181
tri 1784 165 1800 181 nw
rect 1830 227 1842 261
rect 1876 227 1886 261
rect 1830 193 1886 227
tri 1500 127 1530 157 sw
tri 1606 127 1636 157 se
rect 1636 135 1694 159
tri 1694 135 1724 165 sw
tri 1800 135 1830 165 se
rect 1830 159 1842 193
rect 1876 159 1886 193
rect 1830 135 1886 159
rect 1636 127 1886 135
rect 1444 123 1886 127
rect 1444 89 1454 123
rect 1488 89 1648 123
rect 1682 89 1745 123
rect 1779 89 1842 123
rect 1876 89 1886 123
rect 1444 73 1886 89
<< pdiff >>
rect 131 1365 187 1405
rect 131 1331 141 1365
rect 175 1331 187 1365
rect 131 1297 187 1331
rect 131 1263 141 1297
rect 175 1263 187 1297
rect 131 1229 187 1263
rect 131 1195 141 1229
rect 175 1195 187 1229
rect 131 1161 187 1195
rect 131 1127 141 1161
rect 175 1127 187 1161
rect 131 1093 187 1127
rect 131 1059 141 1093
rect 175 1059 187 1093
rect 131 1005 187 1059
rect 217 1365 275 1405
rect 217 1331 229 1365
rect 263 1331 275 1365
rect 217 1297 275 1331
rect 217 1263 229 1297
rect 263 1263 275 1297
rect 217 1229 275 1263
rect 217 1195 229 1229
rect 263 1195 275 1229
rect 217 1161 275 1195
rect 217 1127 229 1161
rect 263 1127 275 1161
rect 217 1093 275 1127
rect 217 1059 229 1093
rect 263 1059 275 1093
rect 217 1005 275 1059
rect 305 1365 363 1405
rect 305 1331 317 1365
rect 351 1331 363 1365
rect 305 1297 363 1331
rect 305 1263 317 1297
rect 351 1263 363 1297
rect 305 1229 363 1263
rect 305 1195 317 1229
rect 351 1195 363 1229
rect 305 1161 363 1195
rect 305 1127 317 1161
rect 351 1127 363 1161
rect 305 1005 363 1127
rect 393 1365 451 1405
rect 393 1331 405 1365
rect 439 1331 451 1365
rect 393 1297 451 1331
rect 393 1263 405 1297
rect 439 1263 451 1297
rect 393 1229 451 1263
rect 393 1195 405 1229
rect 439 1195 451 1229
rect 393 1161 451 1195
rect 393 1127 405 1161
rect 439 1127 451 1161
rect 393 1005 451 1127
rect 481 1365 535 1405
rect 481 1331 493 1365
rect 527 1331 535 1365
rect 481 1297 535 1331
rect 481 1263 493 1297
rect 527 1263 535 1297
rect 481 1229 535 1263
rect 481 1195 493 1229
rect 527 1195 535 1229
rect 481 1161 535 1195
rect 481 1127 493 1161
rect 527 1127 535 1161
rect 481 1093 535 1127
rect 481 1059 493 1093
rect 527 1059 535 1093
rect 481 1005 535 1059
rect 797 1365 851 1405
rect 797 1331 805 1365
rect 839 1331 851 1365
rect 797 1297 851 1331
rect 797 1263 805 1297
rect 839 1263 851 1297
rect 797 1229 851 1263
rect 797 1195 805 1229
rect 839 1195 851 1229
rect 797 1161 851 1195
rect 797 1127 805 1161
rect 839 1127 851 1161
rect 797 1005 851 1127
rect 881 1297 939 1405
rect 881 1263 893 1297
rect 927 1263 939 1297
rect 881 1229 939 1263
rect 881 1195 893 1229
rect 927 1195 939 1229
rect 881 1161 939 1195
rect 881 1127 893 1161
rect 927 1127 939 1161
rect 881 1093 939 1127
rect 881 1059 893 1093
rect 927 1059 939 1093
rect 881 1005 939 1059
rect 969 1365 1027 1405
rect 969 1331 981 1365
rect 1015 1331 1027 1365
rect 969 1297 1027 1331
rect 969 1263 981 1297
rect 1015 1263 1027 1297
rect 969 1229 1027 1263
rect 969 1195 981 1229
rect 1015 1195 1027 1229
rect 969 1161 1027 1195
rect 969 1127 981 1161
rect 1015 1127 1027 1161
rect 969 1005 1027 1127
rect 1057 1297 1115 1405
rect 1057 1263 1069 1297
rect 1103 1263 1115 1297
rect 1057 1229 1115 1263
rect 1057 1195 1069 1229
rect 1103 1195 1115 1229
rect 1057 1161 1115 1195
rect 1057 1127 1069 1161
rect 1103 1127 1115 1161
rect 1057 1005 1115 1127
rect 1145 1365 1201 1405
rect 1145 1331 1157 1365
rect 1191 1331 1201 1365
rect 1145 1297 1201 1331
rect 1145 1263 1157 1297
rect 1191 1263 1201 1297
rect 1145 1229 1201 1263
rect 1145 1195 1157 1229
rect 1191 1195 1201 1229
rect 1145 1161 1201 1195
rect 1145 1127 1157 1161
rect 1191 1127 1201 1161
rect 1145 1005 1201 1127
rect 1463 1365 1519 1405
rect 1463 1331 1473 1365
rect 1507 1331 1519 1365
rect 1463 1297 1519 1331
rect 1463 1263 1473 1297
rect 1507 1263 1519 1297
rect 1463 1229 1519 1263
rect 1463 1195 1473 1229
rect 1507 1195 1519 1229
rect 1463 1161 1519 1195
rect 1463 1127 1473 1161
rect 1507 1127 1519 1161
rect 1463 1005 1519 1127
rect 1549 1297 1607 1405
rect 1549 1263 1561 1297
rect 1595 1263 1607 1297
rect 1549 1229 1607 1263
rect 1549 1195 1561 1229
rect 1595 1195 1607 1229
rect 1549 1161 1607 1195
rect 1549 1127 1561 1161
rect 1595 1127 1607 1161
rect 1549 1093 1607 1127
rect 1549 1059 1561 1093
rect 1595 1059 1607 1093
rect 1549 1005 1607 1059
rect 1637 1365 1695 1405
rect 1637 1331 1649 1365
rect 1683 1331 1695 1365
rect 1637 1297 1695 1331
rect 1637 1263 1649 1297
rect 1683 1263 1695 1297
rect 1637 1229 1695 1263
rect 1637 1195 1649 1229
rect 1683 1195 1695 1229
rect 1637 1161 1695 1195
rect 1637 1127 1649 1161
rect 1683 1127 1695 1161
rect 1637 1005 1695 1127
rect 1725 1297 1783 1405
rect 1725 1263 1737 1297
rect 1771 1263 1783 1297
rect 1725 1229 1783 1263
rect 1725 1195 1737 1229
rect 1771 1195 1783 1229
rect 1725 1161 1783 1195
rect 1725 1127 1737 1161
rect 1771 1127 1783 1161
rect 1725 1093 1783 1127
rect 1725 1059 1737 1093
rect 1771 1059 1783 1093
rect 1725 1005 1783 1059
rect 1813 1365 1867 1405
rect 1813 1331 1825 1365
rect 1859 1331 1867 1365
rect 1813 1297 1867 1331
rect 1813 1263 1825 1297
rect 1859 1263 1867 1297
rect 1813 1229 1867 1263
rect 1813 1195 1825 1229
rect 1859 1195 1867 1229
rect 1813 1161 1867 1195
rect 1813 1127 1825 1161
rect 1859 1127 1867 1161
rect 1813 1005 1867 1127
<< ndiffc >>
rect 122 299 156 333
rect 219 299 253 333
rect 316 299 350 333
rect 510 299 544 333
rect 122 227 156 261
rect 122 159 156 193
rect 219 174 253 208
rect 316 227 350 261
rect 316 159 350 193
rect 412 183 446 217
rect 510 227 544 261
rect 510 159 544 193
rect 122 89 156 123
rect 316 89 350 123
rect 412 89 446 123
rect 510 89 544 123
rect 788 299 822 333
rect 885 299 919 333
rect 982 299 1016 333
rect 1176 299 1210 333
rect 788 227 822 261
rect 788 159 822 193
rect 885 174 919 208
rect 982 227 1016 261
rect 982 159 1016 193
rect 1079 183 1113 217
rect 1176 227 1210 261
rect 1176 159 1210 193
rect 788 89 822 123
rect 982 89 1016 123
rect 1079 89 1113 123
rect 1176 89 1210 123
rect 1454 299 1488 333
rect 1551 299 1585 333
rect 1648 299 1682 333
rect 1454 227 1488 261
rect 1454 159 1488 193
rect 1551 174 1585 208
rect 1648 227 1682 261
rect 1648 159 1682 193
rect 1745 183 1779 217
rect 1842 227 1876 261
rect 1842 159 1876 193
rect 1454 89 1488 123
rect 1648 89 1682 123
rect 1745 89 1779 123
rect 1842 89 1876 123
<< pdiffc >>
rect 141 1331 175 1365
rect 141 1263 175 1297
rect 141 1195 175 1229
rect 141 1127 175 1161
rect 141 1059 175 1093
rect 229 1331 263 1365
rect 229 1263 263 1297
rect 229 1195 263 1229
rect 229 1127 263 1161
rect 229 1059 263 1093
rect 317 1331 351 1365
rect 317 1263 351 1297
rect 317 1195 351 1229
rect 317 1127 351 1161
rect 405 1331 439 1365
rect 405 1263 439 1297
rect 405 1195 439 1229
rect 405 1127 439 1161
rect 493 1331 527 1365
rect 493 1263 527 1297
rect 493 1195 527 1229
rect 493 1127 527 1161
rect 493 1059 527 1093
rect 805 1331 839 1365
rect 805 1263 839 1297
rect 805 1195 839 1229
rect 805 1127 839 1161
rect 893 1263 927 1297
rect 893 1195 927 1229
rect 893 1127 927 1161
rect 893 1059 927 1093
rect 981 1331 1015 1365
rect 981 1263 1015 1297
rect 981 1195 1015 1229
rect 981 1127 1015 1161
rect 1069 1263 1103 1297
rect 1069 1195 1103 1229
rect 1069 1127 1103 1161
rect 1157 1331 1191 1365
rect 1157 1263 1191 1297
rect 1157 1195 1191 1229
rect 1157 1127 1191 1161
rect 1473 1331 1507 1365
rect 1473 1263 1507 1297
rect 1473 1195 1507 1229
rect 1473 1127 1507 1161
rect 1561 1263 1595 1297
rect 1561 1195 1595 1229
rect 1561 1127 1595 1161
rect 1561 1059 1595 1093
rect 1649 1331 1683 1365
rect 1649 1263 1683 1297
rect 1649 1195 1683 1229
rect 1649 1127 1683 1161
rect 1737 1263 1771 1297
rect 1737 1195 1771 1229
rect 1737 1127 1771 1161
rect 1737 1059 1771 1093
rect 1825 1331 1859 1365
rect 1825 1263 1859 1297
rect 1825 1195 1859 1229
rect 1825 1127 1859 1161
<< psubdiff >>
rect -34 482 2032 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 632 461 700 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 632 427 649 461
rect 683 427 700 461
rect 1298 461 1366 482
rect 632 387 700 427
rect -34 313 34 353
rect 632 353 649 387
rect 683 353 700 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 632 313 700 353
rect 1298 427 1315 461
rect 1349 427 1366 461
rect 1964 461 2032 482
rect 1298 387 1366 427
rect 1298 353 1315 387
rect 1349 353 1366 387
rect 1964 427 1981 461
rect 2015 427 2032 461
rect 1964 387 2032 427
rect 632 279 649 313
rect 683 279 700 313
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect -34 17 34 57
rect 632 57 649 91
rect 683 57 700 91
rect 1298 313 1366 353
rect 1964 353 1981 387
rect 2015 353 2032 387
rect 1298 279 1315 313
rect 1349 279 1366 313
rect 1298 239 1366 279
rect 1298 205 1315 239
rect 1349 205 1366 239
rect 1298 165 1366 205
rect 1298 131 1315 165
rect 1349 131 1366 165
rect 1298 91 1366 131
rect 632 17 700 57
rect 1298 57 1315 91
rect 1349 57 1366 91
rect 1964 313 2032 353
rect 1964 279 1981 313
rect 2015 279 2032 313
rect 1964 239 2032 279
rect 1964 205 1981 239
rect 2015 205 2032 239
rect 1964 165 2032 205
rect 1964 131 1981 165
rect 2015 131 2032 165
rect 1964 91 2032 131
rect 1298 17 1366 57
rect 1964 57 1981 91
rect 2015 57 2032 91
rect 1964 17 2032 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 2032 17
rect -34 -34 2032 -17
<< nsubdiff >>
rect -34 1497 2032 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 2032 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 632 1423 700 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 1298 1423 1366 1463
rect 1946 1459 2032 1463
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 632 979 700 1019
rect 1298 1389 1315 1423
rect 1349 1389 1366 1423
rect 1964 1423 2032 1459
rect 1298 1349 1366 1389
rect 1298 1315 1315 1349
rect 1349 1315 1366 1349
rect 1298 1275 1366 1315
rect 1298 1241 1315 1275
rect 1349 1241 1366 1275
rect 1298 1201 1366 1241
rect 1298 1167 1315 1201
rect 1349 1167 1366 1201
rect 1298 1127 1366 1167
rect 1298 1093 1315 1127
rect 1349 1093 1366 1127
rect 1298 1053 1366 1093
rect 1298 1019 1315 1053
rect 1349 1019 1366 1053
rect 632 945 649 979
rect 683 945 700 979
rect -34 871 -17 905
rect 17 884 34 905
rect 632 905 700 945
rect 1298 979 1366 1019
rect 1964 1389 1981 1423
rect 2015 1389 2032 1423
rect 1964 1349 2032 1389
rect 1964 1315 1981 1349
rect 2015 1315 2032 1349
rect 1964 1275 2032 1315
rect 1964 1241 1981 1275
rect 2015 1241 2032 1275
rect 1964 1201 2032 1241
rect 1964 1167 1981 1201
rect 2015 1167 2032 1201
rect 1964 1127 2032 1167
rect 1964 1093 1981 1127
rect 2015 1093 2032 1127
rect 1964 1053 2032 1093
rect 1964 1019 1981 1053
rect 2015 1019 2032 1053
rect 1298 945 1315 979
rect 1349 945 1366 979
rect 632 884 649 905
rect 17 871 649 884
rect 683 884 700 905
rect 1298 905 1366 945
rect 1964 979 2032 1019
rect 1964 945 1981 979
rect 2015 945 2032 979
rect 1298 884 1315 905
rect 683 871 1315 884
rect 1349 884 1366 905
rect 1964 905 2032 945
rect 1964 884 1981 905
rect 1349 871 1981 884
rect 2015 871 2032 905
rect -34 822 2032 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 649 427 683 461
rect 649 353 683 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1315 427 1349 461
rect 1315 353 1349 387
rect 1981 427 2015 461
rect 649 279 683 313
rect 649 205 683 239
rect 649 131 683 165
rect 649 57 683 91
rect 1981 353 2015 387
rect 1315 279 1349 313
rect 1315 205 1349 239
rect 1315 131 1349 165
rect 1315 57 1349 91
rect 1981 279 2015 313
rect 1981 205 2015 239
rect 1981 131 2015 165
rect 1981 57 2015 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 649 1389 683 1423
rect 649 1315 683 1349
rect 649 1241 683 1275
rect 649 1167 683 1201
rect 649 1093 683 1127
rect 649 1019 683 1053
rect -17 945 17 979
rect 1315 1389 1349 1423
rect 1315 1315 1349 1349
rect 1315 1241 1349 1275
rect 1315 1167 1349 1201
rect 1315 1093 1349 1127
rect 1315 1019 1349 1053
rect 649 945 683 979
rect -17 871 17 905
rect 1981 1389 2015 1423
rect 1981 1315 2015 1349
rect 1981 1241 2015 1275
rect 1981 1167 2015 1201
rect 1981 1093 2015 1127
rect 1981 1019 2015 1053
rect 1315 945 1349 979
rect 649 871 683 905
rect 1981 945 2015 979
rect 1315 871 1349 905
rect 1981 871 2015 905
<< poly >>
rect 187 1405 217 1431
rect 275 1405 305 1431
rect 363 1405 393 1431
rect 451 1405 481 1431
rect 851 1405 881 1431
rect 939 1405 969 1431
rect 1027 1405 1057 1431
rect 1115 1405 1145 1431
rect 187 974 217 1005
rect 275 974 305 1005
rect 363 974 393 1005
rect 451 974 481 1005
rect 121 958 305 974
rect 121 924 131 958
rect 165 944 305 958
rect 351 958 481 974
rect 165 924 175 944
rect 121 908 175 924
rect 351 924 361 958
rect 395 944 481 958
rect 1519 1405 1549 1431
rect 1607 1405 1637 1431
rect 1695 1405 1725 1431
rect 1783 1405 1813 1431
rect 395 924 405 944
rect 351 908 405 924
rect 851 974 881 1005
rect 939 974 969 1005
rect 851 958 969 974
rect 851 944 871 958
rect 861 924 871 944
rect 905 944 969 958
rect 1027 974 1057 1005
rect 1115 974 1145 1005
rect 1027 958 1211 974
rect 1027 944 1167 958
rect 905 924 915 944
rect 861 908 915 924
rect 1157 924 1167 944
rect 1201 924 1211 958
rect 1157 908 1211 924
rect 1519 974 1549 1005
rect 1607 974 1637 1005
rect 1695 974 1725 1005
rect 1783 974 1813 1005
rect 1453 958 1637 974
rect 1453 924 1463 958
rect 1497 944 1637 958
rect 1679 958 1813 974
rect 1497 924 1507 944
rect 1453 908 1507 924
rect 1679 924 1689 958
rect 1723 944 1813 958
rect 1723 924 1733 944
rect 1679 908 1733 924
rect 121 433 175 449
rect 121 399 131 433
rect 165 413 175 433
rect 343 433 397 449
rect 165 399 198 413
rect 121 383 198 399
rect 343 399 353 433
rect 387 399 397 433
rect 343 383 397 399
rect 861 433 915 449
rect 861 413 871 433
rect 168 349 198 383
rect 362 349 392 383
rect 834 399 871 413
rect 905 399 915 433
rect 1157 433 1211 449
rect 1157 413 1167 433
rect 834 383 915 399
rect 1134 399 1167 413
rect 1201 399 1211 433
rect 1134 383 1211 399
rect 834 349 864 383
rect 1134 349 1164 383
rect 1453 433 1507 449
rect 1453 399 1463 433
rect 1497 413 1507 433
rect 1675 433 1729 449
rect 1497 399 1530 413
rect 1453 383 1530 399
rect 1675 399 1685 433
rect 1719 399 1729 433
rect 1675 383 1729 399
rect 1500 349 1530 383
rect 1694 349 1724 383
<< polycont >>
rect 131 924 165 958
rect 361 924 395 958
rect 871 924 905 958
rect 1167 924 1201 958
rect 1463 924 1497 958
rect 1689 924 1723 958
rect 131 399 165 433
rect 353 399 387 433
rect 871 399 905 433
rect 1167 399 1201 433
rect 1463 399 1497 433
rect 1685 399 1719 433
<< locali >>
rect -34 1497 2032 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 2032 1497
rect -34 1446 2032 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 141 1365 175 1446
rect 141 1297 175 1331
rect 141 1229 175 1263
rect 141 1161 175 1195
rect 141 1093 175 1127
rect 141 1025 175 1059
rect 229 1365 265 1399
rect 317 1365 351 1446
rect 229 1297 263 1331
rect 229 1229 263 1263
rect 229 1161 263 1195
rect 229 1093 263 1127
rect 317 1297 351 1331
rect 317 1229 351 1263
rect 317 1161 351 1195
rect 317 1111 351 1127
rect 405 1365 439 1399
rect 405 1297 439 1331
rect 405 1229 439 1263
rect 405 1161 439 1195
rect 405 1059 439 1127
rect 229 1025 405 1059
rect 493 1365 527 1446
rect 493 1297 527 1331
rect 493 1229 527 1263
rect 493 1161 527 1195
rect 493 1093 527 1127
rect 493 1025 527 1059
rect 632 1423 700 1446
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 1298 1423 1366 1446
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 632 1053 700 1093
rect -34 979 34 1019
rect 405 1009 439 1025
rect 632 1019 649 1053
rect 683 1019 700 1053
rect -34 945 -17 979
rect 17 945 34 979
rect 632 979 700 1019
rect 805 1365 1191 1399
rect 805 1297 839 1331
rect 805 1229 839 1263
rect 805 1161 839 1195
rect 805 1059 839 1127
rect 893 1297 927 1313
rect 893 1229 927 1263
rect 893 1161 927 1195
rect 893 1093 927 1127
rect 981 1297 1015 1331
rect 981 1229 1015 1263
rect 981 1161 1015 1195
rect 981 1111 1015 1127
rect 1069 1297 1103 1313
rect 1069 1229 1103 1263
rect 1069 1161 1103 1195
rect 1069 1059 1103 1127
rect 1157 1297 1191 1331
rect 1157 1229 1191 1263
rect 1157 1161 1191 1195
rect 1157 1075 1191 1127
rect 1298 1389 1315 1423
rect 1349 1389 1366 1423
rect 1964 1423 2032 1446
rect 1298 1349 1366 1389
rect 1298 1315 1315 1349
rect 1349 1315 1366 1349
rect 1298 1275 1366 1315
rect 1298 1241 1315 1275
rect 1349 1241 1366 1275
rect 1298 1201 1366 1241
rect 1298 1167 1315 1201
rect 1349 1167 1366 1201
rect 1298 1127 1366 1167
rect 1298 1093 1315 1127
rect 1349 1093 1366 1127
rect 893 1025 1069 1059
rect 805 1009 839 1025
rect 1069 1009 1103 1025
rect 1298 1053 1366 1093
rect 1298 1019 1315 1053
rect 1349 1019 1366 1053
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 131 958 165 974
rect 361 958 395 974
rect 131 905 165 924
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 131 433 165 871
rect 131 383 165 399
rect 353 924 361 942
rect 353 908 395 924
rect 632 945 649 979
rect 683 945 700 979
rect 1298 979 1366 1019
rect 1473 1365 1859 1399
rect 1473 1297 1507 1331
rect 1473 1229 1507 1263
rect 1473 1161 1507 1195
rect 1473 1059 1507 1127
rect 1561 1297 1595 1313
rect 1561 1229 1595 1263
rect 1561 1161 1595 1195
rect 1561 1093 1595 1127
rect 1649 1297 1683 1331
rect 1649 1229 1683 1263
rect 1649 1161 1683 1195
rect 1649 1111 1683 1127
rect 1737 1297 1771 1313
rect 1737 1229 1771 1263
rect 1737 1161 1771 1195
rect 1737 1093 1771 1127
rect 1825 1297 1859 1331
rect 1825 1229 1859 1263
rect 1825 1161 1859 1195
rect 1825 1111 1859 1127
rect 1964 1389 1981 1423
rect 2015 1389 2032 1423
rect 1964 1349 2032 1389
rect 1964 1315 1981 1349
rect 2015 1315 2032 1349
rect 1964 1275 2032 1315
rect 1964 1241 1981 1275
rect 2015 1241 2032 1275
rect 1964 1201 2032 1241
rect 1964 1167 1981 1201
rect 2015 1167 2032 1201
rect 1964 1127 2032 1167
rect 1964 1093 1981 1127
rect 2015 1093 2032 1127
rect 1561 1025 1867 1059
rect 1473 1009 1507 1025
rect 353 831 387 908
rect 632 905 700 945
rect 632 871 649 905
rect 683 871 700 905
rect 632 822 700 871
rect 871 958 905 974
rect 871 905 905 924
rect 353 433 387 797
rect 353 383 387 399
rect 632 461 700 544
rect 632 427 649 461
rect 683 427 700 461
rect 632 387 700 427
rect -34 313 34 353
rect 632 353 649 387
rect 683 353 700 387
rect 871 433 905 871
rect 871 383 905 399
rect 1167 958 1201 974
rect 1167 433 1201 924
rect 1298 945 1315 979
rect 1349 945 1366 979
rect 1298 905 1366 945
rect 1298 871 1315 905
rect 1349 871 1366 905
rect 1298 822 1366 871
rect 1463 958 1497 974
rect 1167 383 1201 399
rect 1298 461 1366 544
rect 1298 427 1315 461
rect 1349 427 1366 461
rect 1298 387 1366 427
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 122 333 156 349
rect 316 333 350 349
rect 156 299 219 333
rect 253 299 316 333
rect 122 261 156 299
rect 122 193 156 227
rect 316 261 350 299
rect 510 333 544 349
rect 413 253 447 269
rect 122 123 156 159
rect 122 73 156 89
rect 219 208 253 224
rect -34 34 34 57
rect 219 34 253 174
rect 316 193 350 227
rect 412 219 413 234
rect 412 217 447 219
rect 446 203 447 217
rect 510 261 544 299
rect 412 167 446 183
rect 510 193 544 227
rect 316 123 350 159
rect 510 123 544 159
rect 350 89 412 123
rect 446 89 510 123
rect 316 73 350 89
rect 510 73 544 89
rect 632 313 700 353
rect 1298 353 1315 387
rect 1349 353 1366 387
rect 1463 433 1497 924
rect 1463 383 1497 399
rect 1685 958 1723 974
rect 1685 924 1689 958
rect 1685 908 1723 924
rect 1685 831 1719 908
rect 1685 433 1719 797
rect 1685 383 1719 399
rect 632 279 649 313
rect 683 279 700 313
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect 632 57 649 91
rect 683 57 700 91
rect 788 333 822 349
rect 982 333 1016 349
rect 822 299 885 333
rect 919 299 982 333
rect 788 261 822 299
rect 788 193 822 227
rect 982 261 1016 299
rect 1176 333 1210 349
rect 788 123 822 159
rect 788 73 822 89
rect 885 208 919 224
rect 632 34 700 57
rect 885 34 919 174
rect 982 193 1016 227
rect 1079 253 1113 269
rect 1079 217 1113 219
rect 1079 167 1113 183
rect 1176 261 1210 299
rect 1176 193 1210 227
rect 982 123 1016 159
rect 1176 123 1210 159
rect 1016 89 1079 123
rect 1113 89 1176 123
rect 982 73 1016 89
rect 1176 73 1210 89
rect 1298 313 1366 353
rect 1298 279 1315 313
rect 1349 279 1366 313
rect 1298 239 1366 279
rect 1298 205 1315 239
rect 1349 205 1366 239
rect 1298 165 1366 205
rect 1298 131 1315 165
rect 1349 131 1366 165
rect 1298 91 1366 131
rect 1298 57 1315 91
rect 1349 57 1366 91
rect 1454 333 1488 349
rect 1648 333 1682 349
rect 1833 346 1867 1025
rect 1964 1053 2032 1093
rect 1964 1019 1981 1053
rect 2015 1019 2032 1053
rect 1964 979 2032 1019
rect 1964 945 1981 979
rect 2015 945 2032 979
rect 1964 905 2032 945
rect 1964 871 1981 905
rect 2015 871 2032 905
rect 1964 822 2032 871
rect 1488 299 1551 333
rect 1585 299 1648 333
rect 1454 261 1488 299
rect 1454 193 1488 227
rect 1648 261 1682 299
rect 1454 123 1488 159
rect 1454 73 1488 89
rect 1551 208 1585 224
rect 1298 34 1366 57
rect 1551 34 1585 174
rect 1648 193 1682 227
rect 1745 312 1867 346
rect 1964 461 2032 544
rect 1964 427 1981 461
rect 2015 427 2032 461
rect 1964 387 2032 427
rect 1964 353 1981 387
rect 2015 353 2032 387
rect 1964 313 2032 353
rect 1745 253 1779 312
rect 1964 279 1981 313
rect 2015 279 2032 313
rect 1745 217 1779 219
rect 1745 167 1779 183
rect 1842 261 1876 278
rect 1842 193 1876 227
rect 1648 123 1682 159
rect 1842 123 1876 159
rect 1682 89 1745 123
rect 1779 89 1842 123
rect 1648 73 1682 89
rect 1842 73 1876 89
rect 1964 239 2032 279
rect 1964 205 1981 239
rect 2015 205 2032 239
rect 1964 165 2032 205
rect 1964 131 1981 165
rect 2015 131 2032 165
rect 1964 91 2032 131
rect 1964 57 1981 91
rect 2015 57 2032 91
rect 1964 34 2032 57
rect -34 17 2032 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 2032 17
rect -34 -34 2032 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 405 1025 439 1059
rect 805 1025 839 1059
rect 1069 1025 1103 1059
rect 131 871 165 905
rect 1473 1025 1507 1059
rect 353 797 387 831
rect 871 871 905 905
rect 1167 399 1201 433
rect 413 219 447 253
rect 1463 399 1497 433
rect 1685 797 1719 831
rect 1079 219 1113 253
rect 1745 219 1779 253
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
<< metal1 >>
rect -34 1497 2032 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 2032 1497
rect -34 1446 2032 1463
rect 399 1059 445 1065
rect 799 1059 845 1065
rect 1063 1059 1109 1065
rect 1467 1059 1513 1065
rect 393 1025 405 1059
rect 439 1025 805 1059
rect 839 1025 851 1059
rect 1057 1025 1069 1059
rect 1103 1025 1473 1059
rect 1507 1025 1519 1059
rect 399 1019 445 1025
rect 799 1019 845 1025
rect 1063 1019 1109 1025
rect 1467 1019 1513 1025
rect 125 905 171 911
rect 865 905 911 911
rect 119 871 131 905
rect 165 871 871 905
rect 905 871 917 905
rect 125 865 171 871
rect 865 865 911 871
rect 347 831 393 837
rect 1679 831 1725 837
rect 341 797 353 831
rect 387 797 1685 831
rect 1719 797 1731 831
rect 347 791 393 797
rect 1679 791 1725 797
rect 1161 433 1207 439
rect 1457 433 1503 439
rect 1155 399 1167 433
rect 1201 399 1463 433
rect 1497 399 1509 433
rect 1161 393 1207 399
rect 1457 393 1503 399
rect 407 253 453 259
rect 1073 253 1119 259
rect 1739 253 1785 259
rect 401 219 413 253
rect 447 219 1079 253
rect 1113 219 1745 253
rect 1779 219 1791 253
rect 407 213 453 219
rect 1073 213 1119 219
rect 1739 213 1785 219
rect -34 17 2032 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 2032 17
rect -34 -34 2032 -17
<< labels >>
rlabel metal1 1833 649 1867 683 1 YN
port 1 n
rlabel metal1 1833 723 1867 757 1 YN
port 2 n
rlabel metal1 1833 797 1867 831 1 YN
port 3 n
rlabel metal1 1833 871 1867 905 1 YN
port 4 n
rlabel metal1 1833 945 1867 979 1 YN
port 5 n
rlabel metal1 1833 575 1867 609 1 YN
port 6 n
rlabel metal1 1833 501 1867 535 1 YN
port 7 n
rlabel metal1 1833 427 1867 461 1 YN
port 8 n
rlabel metal1 353 723 387 757 1 A
port 9 n
rlabel metal1 353 797 387 831 1 A
port 10 n
rlabel metal1 353 649 387 683 1 A
port 11 n
rlabel metal1 353 575 387 609 1 A
port 12 n
rlabel metal1 353 501 387 535 1 A
port 13 n
rlabel metal1 1685 501 1719 535 1 A
port 14 n
rlabel metal1 1685 575 1719 609 1 A
port 15 n
rlabel metal1 1685 649 1719 683 1 A
port 16 n
rlabel metal1 1685 723 1719 757 1 A
port 17 n
rlabel metal1 1685 797 1719 831 1 A
port 18 n
rlabel metal1 1685 871 1719 905 1 A
port 19 n
rlabel metal1 131 797 165 831 1 B
port 20 n
rlabel metal1 131 723 165 757 1 B
port 21 n
rlabel metal1 131 649 165 683 1 B
port 22 n
rlabel metal1 131 575 165 609 1 B
port 23 n
rlabel metal1 131 501 165 535 1 B
port 24 n
rlabel metal1 871 723 905 757 1 B
port 25 n
rlabel metal1 871 649 905 683 1 B
port 26 n
rlabel metal1 871 575 905 609 1 B
port 27 n
rlabel metal1 871 501 905 535 1 B
port 28 n
rlabel metal1 131 871 165 905 1 B
port 29 n
rlabel metal1 871 871 905 905 1 B
port 30 n
rlabel metal1 1167 501 1201 535 1 C
port 31 n
rlabel metal1 1167 575 1201 609 1 C
port 32 n
rlabel metal1 1167 649 1201 683 1 C
port 33 n
rlabel metal1 1167 723 1201 757 1 C
port 34 n
rlabel metal1 1167 871 1201 905 1 C
port 35 n
rlabel metal1 1463 723 1497 757 1 C
port 36 n
rlabel metal1 1463 649 1497 683 1 C
port 37 n
rlabel metal1 1463 575 1497 609 1 C
port 38 n
rlabel metal1 1463 501 1497 535 1 C
port 39 n
rlabel metal1 1463 871 1497 905 1 C
port 40 n
rlabel metal1 -34 1446 2032 1514 1 VPWR
port 41 n
rlabel metal1 -34 -34 2032 34 1 VGND
port 42 n
rlabel nwell 55 1463 89 1497 1 VPB
port 43 n
rlabel pwell 57 -17 91 17 1 VNB
port 44 n
<< end >>
