* SPICE3 file created from MUX2X1.ext - technology: sky130A

.subckt MUX2X1 Y A0 A1 S VDD GND
X0 GND mux2x1_pcell_0/m1_981_575# mux2x1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X1 Y mux2x1_pcell_0/m1_1647_649# mux2x1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X2 VDD mux2x1_pcell_0/m1_981_575# Y VDD pshort w=2 l=0.15
X3 VDD mux2x1_pcell_0/m1_1647_649# Y VDD pshort w=2 l=0.15
X4 mux2x1_pcell_0/m1_315_649# S GND GND nshort w=3 l=0.15
X5 VDD S mux2x1_pcell_0/m1_315_649# VDD pshort w=2 l=0.15
X6 GND S mux2x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X7 mux2x1_pcell_0/m1_981_575# A0 mux2x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X8 VDD S mux2x1_pcell_0/m1_981_575# VDD pshort w=2 l=0.15
X9 VDD A0 mux2x1_pcell_0/m1_981_575# VDD pshort w=2 l=0.15
X10 GND mux2x1_pcell_0/m1_315_649# mux2x1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X11 mux2x1_pcell_0/m1_1647_649# A1 mux2x1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X12 VDD mux2x1_pcell_0/m1_315_649# mux2x1_pcell_0/m1_1647_649# VDD pshort w=2 l=0.15
X13 VDD A1 mux2x1_pcell_0/m1_1647_649# VDD pshort w=2 l=0.15
C0 VDD GND 3.24fF
.ends
