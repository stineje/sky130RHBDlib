* SPICE3 file created from AO3X1.ext - technology: sky130A

.subckt AO3X1 Y A B C VPB VNB
M1000 VNB a_168_157# a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=3.2565p pd=22.61u as=0p ps=0u
M1001 VPB.t5 a_168_157# a_217_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPB.t3 a_217_1004.t5 a_797_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t1 a_343_383# a_217_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1517_182.t2 a_864_181.t4 VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_797_1005.t3 a_1009_383# a_864_181.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_217_1004.t3 a_168_157# VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_217_1004.t2 a_343_383# VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_797_1005.t0 a_217_1004.t6 VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPB.t7 a_864_181.t6 a_1517_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_864_181.t1 a_1009_383# a_797_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 a_168_157# a_343_383# 0.26fF
C1 VPB a_168_157# 0.08fF
C2 VPB a_343_383# 0.07fF
C3 VPB a_1009_383# 0.07fF
R0 a_217_1004.n4 a_217_1004.t6 486.819
R1 a_217_1004.n4 a_217_1004.t5 384.527
R2 a_217_1004.n6 a_217_1004.n3 215.652
R3 a_217_1004.n5 a_217_1004.t7 207.443
R4 a_217_1004.n5 a_217_1004.n4 169.7
R5 a_217_1004.n6 a_217_1004.n5 153.315
R6 a_217_1004.n8 a_217_1004.n6 140.981
R7 a_217_1004.n3 a_217_1004.n2 76.002
R8 a_217_1004.n8 a_217_1004.n7 30
R9 a_217_1004.n9 a_217_1004.n0 24.383
R10 a_217_1004.n9 a_217_1004.n8 23.684
R11 a_217_1004.n1 a_217_1004.t1 14.282
R12 a_217_1004.n1 a_217_1004.t2 14.282
R13 a_217_1004.n2 a_217_1004.t4 14.282
R14 a_217_1004.n2 a_217_1004.t3 14.282
R15 a_217_1004.n3 a_217_1004.n1 12.85
R16 VPB VPB.n184 126.832
R17 VPB.n153 VPB.n151 94.117
R18 VPB.n91 VPB.n89 94.117
R19 VPB.n166 VPB.n165 76
R20 VPB.n105 VPB.n25 76
R21 VPB.n177 VPB.n176 76
R22 VPB.n81 VPB.n80 68.979
R23 VPB.n74 VPB.n73 64.528
R24 VPB.n113 VPB.n112 61.764
R25 VPB.n33 VPB.n32 61.764
R26 VPB.n129 VPB.t4 55.106
R27 VPB.n84 VPB.t6 55.106
R28 VPB.n72 VPB.t7 55.106
R29 VPB.n147 VPB.t1 55.106
R30 VPB.n144 VPB.n143 48.952
R31 VPB.n163 VPB.n162 44.502
R32 VPB.n131 VPB.n130 44.502
R33 VPB.n106 VPB.n26 41.183
R34 VPB.n138 VPB.n128 40.824
R35 VPB.n181 VPB.n177 20.452
R36 VPB.n71 VPB.n68 20.452
R37 VPB.n140 VPB.n139 17.801
R38 VPB.n128 VPB.t0 14.282
R39 VPB.n128 VPB.t5 14.282
R40 VPB.n26 VPB.t2 14.282
R41 VPB.n26 VPB.t3 14.282
R42 VPB.n71 VPB.n70 13.653
R43 VPB.n70 VPB.n69 13.653
R44 VPB.n76 VPB.n75 13.653
R45 VPB.n75 VPB.n74 13.653
R46 VPB.n79 VPB.n78 13.653
R47 VPB.n78 VPB.n77 13.653
R48 VPB.n83 VPB.n82 13.653
R49 VPB.n82 VPB.n81 13.653
R50 VPB.n87 VPB.n86 13.653
R51 VPB.n86 VPB.n85 13.653
R52 VPB.n92 VPB.n91 13.653
R53 VPB.n91 VPB.n90 13.653
R54 VPB.n95 VPB.n94 13.653
R55 VPB.n94 VPB.n93 13.653
R56 VPB.n98 VPB.n97 13.653
R57 VPB.n97 VPB.n96 13.653
R58 VPB.n101 VPB.n100 13.653
R59 VPB.n100 VPB.n99 13.653
R60 VPB.n105 VPB.n104 13.653
R61 VPB.n104 VPB.n103 13.653
R62 VPB.n165 VPB.n164 13.653
R63 VPB.n164 VPB.n163 13.653
R64 VPB.n161 VPB.n160 13.653
R65 VPB.n160 VPB.n159 13.653
R66 VPB.n158 VPB.n157 13.653
R67 VPB.n157 VPB.n156 13.653
R68 VPB.n154 VPB.n153 13.653
R69 VPB.n153 VPB.n152 13.653
R70 VPB.n150 VPB.n149 13.653
R71 VPB.n149 VPB.n148 13.653
R72 VPB.n146 VPB.n145 13.653
R73 VPB.n145 VPB.n144 13.653
R74 VPB.n142 VPB.n141 13.653
R75 VPB.n141 VPB.n140 13.653
R76 VPB.n137 VPB.n136 13.653
R77 VPB.n136 VPB.n135 13.653
R78 VPB.n133 VPB.n132 13.653
R79 VPB.n132 VPB.n131 13.653
R80 VPB.n16 VPB.n15 13.653
R81 VPB.n15 VPB.n14 13.653
R82 VPB.n177 VPB.n0 13.653
R83 VPB VPB.n0 13.653
R84 VPB.n103 VPB.n102 13.35
R85 VPB.n135 VPB.n134 13.35
R86 VPB.n181 VPB.n180 13.276
R87 VPB.n180 VPB.n178 13.276
R88 VPB.n127 VPB.n109 13.276
R89 VPB.n109 VPB.n107 13.276
R90 VPB.n47 VPB.n29 13.276
R91 VPB.n29 VPB.n27 13.276
R92 VPB.n79 VPB.n76 13.276
R93 VPB.n83 VPB.n79 13.276
R94 VPB.n88 VPB.n87 13.276
R95 VPB.n92 VPB.n88 13.276
R96 VPB.n95 VPB.n92 13.276
R97 VPB.n98 VPB.n95 13.276
R98 VPB.n101 VPB.n98 13.276
R99 VPB.n105 VPB.n101 13.276
R100 VPB.n165 VPB.n161 13.276
R101 VPB.n161 VPB.n158 13.276
R102 VPB.n158 VPB.n155 13.276
R103 VPB.n155 VPB.n154 13.276
R104 VPB.n154 VPB.n150 13.276
R105 VPB.n146 VPB.n142 13.276
R106 VPB.n137 VPB.n133 13.276
R107 VPB.n177 VPB.n16 13.276
R108 VPB.n68 VPB.n50 13.276
R109 VPB.n50 VPB.n48 13.276
R110 VPB.n55 VPB.n53 12.796
R111 VPB.n55 VPB.n54 12.564
R112 VPB.n63 VPB.n62 12.198
R113 VPB.n63 VPB.n60 12.198
R114 VPB.n58 VPB.n57 12.198
R115 VPB.n147 VPB.n146 11.841
R116 VPB.n133 VPB.n129 11.482
R117 VPB.n87 VPB.n84 10.944
R118 VPB.n72 VPB.n71 10.585
R119 VPB.n106 VPB.n105 8.97
R120 VPB.n68 VPB.n67 7.5
R121 VPB.n53 VPB.n52 7.5
R122 VPB.n57 VPB.n56 7.5
R123 VPB.n62 VPB.n61 7.5
R124 VPB.n50 VPB.n49 7.5
R125 VPB.n65 VPB.n51 7.5
R126 VPB.n29 VPB.n28 7.5
R127 VPB.n42 VPB.n41 7.5
R128 VPB.n36 VPB.n35 7.5
R129 VPB.n38 VPB.n37 7.5
R130 VPB.n31 VPB.n30 7.5
R131 VPB.n47 VPB.n46 7.5
R132 VPB.n109 VPB.n108 7.5
R133 VPB.n122 VPB.n121 7.5
R134 VPB.n116 VPB.n115 7.5
R135 VPB.n118 VPB.n117 7.5
R136 VPB.n111 VPB.n110 7.5
R137 VPB.n127 VPB.n126 7.5
R138 VPB.n180 VPB.n179 7.5
R139 VPB.n12 VPB.n11 7.5
R140 VPB.n6 VPB.n5 7.5
R141 VPB.n8 VPB.n7 7.5
R142 VPB.n2 VPB.n1 7.5
R143 VPB.n182 VPB.n181 7.5
R144 VPB.n155 VPB.n127 7.176
R145 VPB.n88 VPB.n47 7.176
R146 VPB.n138 VPB.n137 6.817
R147 VPB.n43 VPB.n40 6.729
R148 VPB.n39 VPB.n36 6.729
R149 VPB.n34 VPB.n31 6.729
R150 VPB.n123 VPB.n120 6.729
R151 VPB.n119 VPB.n116 6.729
R152 VPB.n114 VPB.n111 6.729
R153 VPB.n13 VPB.n10 6.729
R154 VPB.n9 VPB.n6 6.729
R155 VPB.n4 VPB.n2 6.729
R156 VPB.n34 VPB.n33 6.728
R157 VPB.n39 VPB.n38 6.728
R158 VPB.n43 VPB.n42 6.728
R159 VPB.n46 VPB.n45 6.728
R160 VPB.n114 VPB.n113 6.728
R161 VPB.n119 VPB.n118 6.728
R162 VPB.n123 VPB.n122 6.728
R163 VPB.n126 VPB.n125 6.728
R164 VPB.n4 VPB.n3 6.728
R165 VPB.n9 VPB.n8 6.728
R166 VPB.n13 VPB.n12 6.728
R167 VPB.n183 VPB.n182 6.728
R168 VPB.n142 VPB.n138 6.458
R169 VPB.n67 VPB.n66 6.398
R170 VPB.n165 VPB.n106 4.305
R171 VPB.n76 VPB.n72 2.691
R172 VPB.n84 VPB.n83 2.332
R173 VPB.n129 VPB.n16 1.794
R174 VPB.n150 VPB.n147 1.435
R175 VPB.n65 VPB.n58 1.402
R176 VPB.n65 VPB.n59 1.402
R177 VPB.n65 VPB.n63 1.402
R178 VPB.n65 VPB.n64 1.402
R179 VPB.n66 VPB.n65 0.735
R180 VPB.n65 VPB.n55 0.735
R181 VPB.n44 VPB.n43 0.387
R182 VPB.n44 VPB.n39 0.387
R183 VPB.n44 VPB.n34 0.387
R184 VPB.n45 VPB.n44 0.387
R185 VPB.n124 VPB.n123 0.387
R186 VPB.n124 VPB.n119 0.387
R187 VPB.n124 VPB.n114 0.387
R188 VPB.n125 VPB.n124 0.387
R189 VPB.n184 VPB.n13 0.387
R190 VPB.n184 VPB.n9 0.387
R191 VPB.n184 VPB.n4 0.387
R192 VPB.n184 VPB.n183 0.387
R193 VPB.n21 VPB.n20 0.272
R194 VPB.n169 VPB.n168 0.272
R195 VPB.n176 VPB 0.198
R196 VPB.n18 VPB.n17 0.136
R197 VPB.n19 VPB.n18 0.136
R198 VPB.n20 VPB.n19 0.136
R199 VPB.n22 VPB.n21 0.136
R200 VPB.n23 VPB.n22 0.136
R201 VPB.n24 VPB.n23 0.136
R202 VPB.n25 VPB.n24 0.136
R203 VPB.n166 VPB.n25 0.136
R204 VPB.n167 VPB.n166 0.136
R205 VPB.n168 VPB.n167 0.136
R206 VPB.n170 VPB.n169 0.136
R207 VPB.n171 VPB.n170 0.136
R208 VPB.n172 VPB.n171 0.136
R209 VPB.n173 VPB.n172 0.136
R210 VPB.n174 VPB.n173 0.136
R211 VPB.n175 VPB.n174 0.136
R212 VPB.n176 VPB.n175 0.136
R213 a_797_1005.t1 a_797_1005.n0 101.66
R214 a_797_1005.n0 a_797_1005.t3 101.659
R215 a_797_1005.n0 a_797_1005.t2 14.294
R216 a_797_1005.n0 a_797_1005.t0 14.282
R217 a_112_73.t0 a_112_73.n1 93.333
R218 a_112_73.n4 a_112_73.n2 55.07
R219 a_112_73.t0 a_112_73.n0 8.137
R220 a_112_73.n4 a_112_73.n3 4.619
R221 a_112_73.t0 a_112_73.n4 0.071
R222 a_864_181.n2 a_864_181.t6 512.525
R223 a_864_181.n2 a_864_181.t4 371.139
R224 a_864_181.n4 a_864_181.n1 228.489
R225 a_864_181.n3 a_864_181.n2 211.406
R226 a_864_181.n3 a_864_181.t5 167.157
R227 a_864_181.n4 a_864_181.n3 153.043
R228 a_864_181.n9 a_864_181.n8 118.016
R229 a_864_181.n9 a_864_181.n4 92.576
R230 a_864_181.n12 a_864_181.n0 55.263
R231 a_864_181.n11 a_864_181.n9 48.405
R232 a_864_181.n8 a_864_181.n7 30
R233 a_864_181.n11 a_864_181.n10 30
R234 a_864_181.n12 a_864_181.n11 25.263
R235 a_864_181.n6 a_864_181.n5 24.383
R236 a_864_181.n8 a_864_181.n6 23.684
R237 a_864_181.n1 a_864_181.t2 14.282
R238 a_864_181.n1 a_864_181.t1 14.282
R239 a_1517_182.n3 a_1517_182.n1 355.848
R240 a_1517_182.n3 a_1517_182.n2 30
R241 a_1517_182.n4 a_1517_182.n0 24.383
R242 a_1517_182.n4 a_1517_182.n3 23.684
R243 a_1517_182.n1 a_1517_182.t1 14.282
R244 a_1517_182.n1 a_1517_182.t2 14.282
R245 VNB VNB.n180 300.778
R246 VNB.n34 VNB.n33 199.897
R247 VNB.n118 VNB.n117 199.897
R248 VNB.n87 VNB.n85 154.509
R249 VNB.n143 VNB.n141 154.509
R250 VNB.n128 VNB.n124 84.842
R251 VNB.n156 VNB.n155 76
R252 VNB.n167 VNB.n166 76
R253 VNB.n103 VNB.n15 76
R254 VNB.n154 VNB.n153 62.533
R255 VNB.n75 VNB.n74 49.896
R256 VNB.n126 VNB.n125 36.678
R257 VNB.n94 VNB.n93 36.267
R258 VNB.n50 VNB.n49 35.01
R259 VNB.t2 VNB.n42 32.601
R260 VNB.n68 VNB.n65 20.452
R261 VNB.n168 VNB.n167 20.452
R262 VNB.n69 VNB.n50 20.094
R263 VNB.n73 VNB.n47 20.094
R264 VNB.n80 VNB.n45 20.094
R265 VNB.n104 VNB.n16 19.735
R266 VNB.n100 VNB.n19 19.735
R267 VNB.n96 VNB.n20 19.735
R268 VNB.n89 VNB.n23 19.735
R269 VNB.n149 VNB.n107 19.735
R270 VNB.n50 VNB.n48 19.017
R271 VNB.n44 VNB.t2 17.353
R272 VNB.n106 VNB.t0 17.353
R273 VNB.n18 VNB.t3 13.654
R274 VNB.n72 VNB.n71 13.653
R275 VNB.n71 VNB.n70 13.653
R276 VNB.n76 VNB.n75 13.653
R277 VNB.n79 VNB.n78 13.653
R278 VNB.n78 VNB.n77 13.653
R279 VNB.n83 VNB.n82 13.653
R280 VNB.n82 VNB.n81 13.653
R281 VNB.n88 VNB.n87 13.653
R282 VNB.n87 VNB.n86 13.653
R283 VNB.n92 VNB.n91 13.653
R284 VNB.n91 VNB.n90 13.653
R285 VNB.n95 VNB.n94 13.653
R286 VNB.n99 VNB.n98 13.653
R287 VNB.n98 VNB.n97 13.653
R288 VNB.n103 VNB.n102 13.653
R289 VNB.n102 VNB.n101 13.653
R290 VNB.n155 VNB.n154 13.653
R291 VNB.n152 VNB.n151 13.653
R292 VNB.n151 VNB.n150 13.653
R293 VNB.n148 VNB.n147 13.653
R294 VNB.n147 VNB.n146 13.653
R295 VNB.n144 VNB.n143 13.653
R296 VNB.n143 VNB.n142 13.653
R297 VNB.n140 VNB.n139 13.653
R298 VNB.n139 VNB.n138 13.653
R299 VNB.n137 VNB.n136 13.653
R300 VNB.n136 VNB.n135 13.653
R301 VNB.n134 VNB.n133 13.653
R302 VNB.n133 VNB.n132 13.653
R303 VNB.n131 VNB.n130 13.653
R304 VNB.n130 VNB.n129 13.653
R305 VNB.n127 VNB.n126 13.653
R306 VNB.n6 VNB.n5 13.653
R307 VNB.n5 VNB.n4 13.653
R308 VNB.n167 VNB.n0 13.653
R309 VNB VNB.n0 13.653
R310 VNB.n68 VNB.n67 13.653
R311 VNB.n67 VNB.n66 13.653
R312 VNB.n175 VNB.n172 13.577
R313 VNB.n53 VNB.n51 13.276
R314 VNB.n65 VNB.n53 13.276
R315 VNB.n26 VNB.n24 13.276
R316 VNB.n39 VNB.n26 13.276
R317 VNB.n110 VNB.n108 13.276
R318 VNB.n123 VNB.n110 13.276
R319 VNB.n79 VNB.n76 13.276
R320 VNB.n84 VNB.n83 13.276
R321 VNB.n88 VNB.n84 13.276
R322 VNB.n95 VNB.n92 13.276
R323 VNB.n155 VNB.n152 13.276
R324 VNB.n148 VNB.n145 13.276
R325 VNB.n145 VNB.n144 13.276
R326 VNB.n144 VNB.n140 13.276
R327 VNB.n140 VNB.n137 13.276
R328 VNB.n137 VNB.n134 13.276
R329 VNB.n134 VNB.n131 13.276
R330 VNB.n127 VNB.n6 13.276
R331 VNB.n167 VNB.n6 13.276
R332 VNB.n3 VNB.n1 13.276
R333 VNB.n168 VNB.n3 13.276
R334 VNB.n73 VNB.n72 13.097
R335 VNB.n45 VNB.n44 12.837
R336 VNB.n107 VNB.n106 12.837
R337 VNB.n89 VNB.n88 11.661
R338 VNB.n149 VNB.n148 11.661
R339 VNB.n23 VNB.n22 11.605
R340 VNB.n99 VNB.n96 10.764
R341 VNB.n104 VNB.n103 10.764
R342 VNB.n131 VNB.n128 10.764
R343 VNB.n22 VNB.n21 9.809
R344 VNB.n83 VNB.n80 9.329
R345 VNB.n69 VNB.n68 8.97
R346 VNB.n44 VNB.n43 7.566
R347 VNB.n106 VNB.n105 7.566
R348 VNB.n177 VNB.n176 7.5
R349 VNB.n32 VNB.n31 7.5
R350 VNB.n28 VNB.n27 7.5
R351 VNB.n26 VNB.n25 7.5
R352 VNB.n39 VNB.n38 7.5
R353 VNB.n116 VNB.n115 7.5
R354 VNB.n112 VNB.n111 7.5
R355 VNB.n110 VNB.n109 7.5
R356 VNB.n123 VNB.n122 7.5
R357 VNB.n169 VNB.n168 7.5
R358 VNB.n3 VNB.n2 7.5
R359 VNB.n174 VNB.n173 7.5
R360 VNB.n59 VNB.n58 7.5
R361 VNB.n55 VNB.n54 7.5
R362 VNB.n53 VNB.n52 7.5
R363 VNB.n65 VNB.n64 7.5
R364 VNB.n84 VNB.n39 7.176
R365 VNB.n145 VNB.n123 7.176
R366 VNB.t3 VNB.n17 7.04
R367 VNB.n179 VNB.n177 7.011
R368 VNB.n35 VNB.n32 7.011
R369 VNB.n30 VNB.n28 7.011
R370 VNB.n119 VNB.n116 7.011
R371 VNB.n114 VNB.n112 7.011
R372 VNB.n61 VNB.n59 7.011
R373 VNB.n57 VNB.n55 7.011
R374 VNB.n38 VNB.n37 7.01
R375 VNB.n30 VNB.n29 7.01
R376 VNB.n35 VNB.n34 7.01
R377 VNB.n122 VNB.n121 7.01
R378 VNB.n114 VNB.n113 7.01
R379 VNB.n119 VNB.n118 7.01
R380 VNB.n64 VNB.n63 7.01
R381 VNB.n57 VNB.n56 7.01
R382 VNB.n61 VNB.n60 7.01
R383 VNB.n179 VNB.n178 7.01
R384 VNB.n175 VNB.n174 6.788
R385 VNB.n170 VNB.n169 6.788
R386 VNB.n100 VNB.n99 6.638
R387 VNB.n103 VNB.n100 6.638
R388 VNB.n19 VNB.n18 5.774
R389 VNB.n41 VNB.n40 4.551
R390 VNB.n72 VNB.n69 4.305
R391 VNB.n80 VNB.n79 3.947
R392 VNB.n96 VNB.n95 2.511
R393 VNB.n155 VNB.n104 2.511
R394 VNB.n128 VNB.n127 2.511
R395 VNB.t2 VNB.n41 2.238
R396 VNB.n92 VNB.n89 1.614
R397 VNB.n152 VNB.n149 1.614
R398 VNB.n180 VNB.n171 0.921
R399 VNB.n180 VNB.n175 0.476
R400 VNB.n180 VNB.n170 0.475
R401 VNB.n47 VNB.n46 0.358
R402 VNB.n11 VNB.n10 0.272
R403 VNB.n159 VNB.n158 0.272
R404 VNB.n36 VNB.n30 0.246
R405 VNB.n37 VNB.n36 0.246
R406 VNB.n36 VNB.n35 0.246
R407 VNB.n120 VNB.n114 0.246
R408 VNB.n121 VNB.n120 0.246
R409 VNB.n120 VNB.n119 0.246
R410 VNB.n62 VNB.n57 0.246
R411 VNB.n63 VNB.n62 0.246
R412 VNB.n62 VNB.n61 0.246
R413 VNB.n180 VNB.n179 0.246
R414 VNB.n166 VNB 0.198
R415 VNB.n76 VNB.n73 0.179
R416 VNB.n8 VNB.n7 0.136
R417 VNB.n9 VNB.n8 0.136
R418 VNB.n10 VNB.n9 0.136
R419 VNB.n12 VNB.n11 0.136
R420 VNB.n13 VNB.n12 0.136
R421 VNB.n14 VNB.n13 0.136
R422 VNB.n15 VNB.n14 0.136
R423 VNB.n156 VNB.n15 0.136
R424 VNB.n157 VNB.n156 0.136
R425 VNB.n158 VNB.n157 0.136
R426 VNB.n160 VNB.n159 0.136
R427 VNB.n161 VNB.n160 0.136
R428 VNB.n162 VNB.n161 0.136
R429 VNB.n163 VNB.n162 0.136
R430 VNB.n164 VNB.n163 0.136
R431 VNB.n165 VNB.n164 0.136
R432 VNB.n166 VNB.n165 0.136
C4 VPB VNB 7.90fF
C5 a_1517_182.n0 VNB 0.04fF
C6 a_1517_182.n1 VNB 1.02fF
C7 a_1517_182.n2 VNB 0.04fF
C8 a_1517_182.n3 VNB 0.50fF
C9 a_1517_182.n4 VNB 0.06fF
C10 a_864_181.n0 VNB 0.04fF
C11 a_864_181.n1 VNB 0.62fF
C12 a_864_181.n2 VNB 0.35fF
C13 a_864_181.t5 VNB 0.39fF
C14 a_864_181.n3 VNB 0.48fF
C15 a_864_181.n4 VNB 0.44fF
C16 a_864_181.n5 VNB 0.03fF
C17 a_864_181.n6 VNB 0.05fF
C18 a_864_181.n7 VNB 0.03fF
C19 a_864_181.n8 VNB 0.15fF
C20 a_864_181.n9 VNB 0.26fF
C21 a_864_181.n10 VNB 0.03fF
C22 a_864_181.n11 VNB 0.08fF
C23 a_864_181.n12 VNB 0.04fF
C24 a_112_73.n0 VNB 0.05fF
C25 a_112_73.n1 VNB 0.02fF
C26 a_112_73.n2 VNB 0.12fF
C27 a_112_73.n3 VNB 0.04fF
C28 a_112_73.n4 VNB 0.16fF
C29 a_797_1005.n0 VNB 0.55fF
C30 VPB.n0 VNB 0.03fF
C31 VPB.n1 VNB 0.03fF
C32 VPB.n2 VNB 0.02fF
C33 VPB.n3 VNB 0.13fF
C34 VPB.n5 VNB 0.02fF
C35 VPB.n6 VNB 0.02fF
C36 VPB.n7 VNB 0.02fF
C37 VPB.n8 VNB 0.02fF
C38 VPB.n10 VNB 0.02fF
C39 VPB.n11 VNB 0.02fF
C40 VPB.n12 VNB 0.02fF
C41 VPB.n14 VNB 0.22fF
C42 VPB.n15 VNB 0.02fF
C43 VPB.n16 VNB 0.01fF
C44 VPB.n17 VNB 0.07fF
C45 VPB.n18 VNB 0.02fF
C46 VPB.n19 VNB 0.02fF
C47 VPB.n20 VNB 0.03fF
C48 VPB.n21 VNB 0.03fF
C49 VPB.n22 VNB 0.02fF
C50 VPB.n23 VNB 0.02fF
C51 VPB.n24 VNB 0.02fF
C52 VPB.n25 VNB 0.02fF
C53 VPB.n26 VNB 0.10fF
C54 VPB.n27 VNB 0.02fF
C55 VPB.n28 VNB 0.02fF
C56 VPB.n29 VNB 0.02fF
C57 VPB.n30 VNB 0.03fF
C58 VPB.n31 VNB 0.02fF
C59 VPB.n32 VNB 0.16fF
C60 VPB.n33 VNB 0.04fF
C61 VPB.n35 VNB 0.02fF
C62 VPB.n36 VNB 0.02fF
C63 VPB.n37 VNB 0.02fF
C64 VPB.n38 VNB 0.02fF
C65 VPB.n40 VNB 0.02fF
C66 VPB.n41 VNB 0.02fF
C67 VPB.n42 VNB 0.02fF
C68 VPB.n44 VNB 0.26fF
C69 VPB.n46 VNB 0.02fF
C70 VPB.n47 VNB 0.02fF
C71 VPB.n48 VNB 0.02fF
C72 VPB.n49 VNB 0.02fF
C73 VPB.n50 VNB 0.02fF
C74 VPB.n51 VNB 0.10fF
C75 VPB.n52 VNB 0.03fF
C76 VPB.n53 VNB 0.02fF
C77 VPB.n54 VNB 0.04fF
C78 VPB.n55 VNB 0.01fF
C79 VPB.n56 VNB 0.02fF
C80 VPB.n57 VNB 0.02fF
C81 VPB.n60 VNB 0.02fF
C82 VPB.n61 VNB 0.02fF
C83 VPB.n62 VNB 0.02fF
C84 VPB.n65 VNB 0.43fF
C85 VPB.n67 VNB 0.03fF
C86 VPB.n68 VNB 0.04fF
C87 VPB.n69 VNB 0.26fF
C88 VPB.n70 VNB 0.03fF
C89 VPB.n71 VNB 0.03fF
C90 VPB.n72 VNB 0.05fF
C91 VPB.n73 VNB 0.13fF
C92 VPB.n74 VNB 0.18fF
C93 VPB.n75 VNB 0.02fF
C94 VPB.n76 VNB 0.01fF
C95 VPB.n77 VNB 0.15fF
C96 VPB.n78 VNB 0.02fF
C97 VPB.n79 VNB 0.02fF
C98 VPB.n80 VNB 0.13fF
C99 VPB.n81 VNB 0.18fF
C100 VPB.n82 VNB 0.02fF
C101 VPB.n83 VNB 0.01fF
C102 VPB.n84 VNB 0.05fF
C103 VPB.n85 VNB 0.26fF
C104 VPB.n86 VNB 0.01fF
C105 VPB.n87 VNB 0.02fF
C106 VPB.n88 VNB 0.03fF
C107 VPB.n89 VNB 0.03fF
C108 VPB.n90 VNB 0.26fF
C109 VPB.n91 VNB 0.01fF
C110 VPB.n92 VNB 0.02fF
C111 VPB.n93 VNB 0.26fF
C112 VPB.n94 VNB 0.02fF
C113 VPB.n95 VNB 0.02fF
C114 VPB.n96 VNB 0.26fF
C115 VPB.n97 VNB 0.02fF
C116 VPB.n98 VNB 0.02fF
C117 VPB.n99 VNB 0.26fF
C118 VPB.n100 VNB 0.02fF
C119 VPB.n101 VNB 0.02fF
C120 VPB.n102 VNB 0.13fF
C121 VPB.n103 VNB 0.14fF
C122 VPB.n104 VNB 0.02fF
C123 VPB.n105 VNB 0.02fF
C124 VPB.n106 VNB 0.02fF
C125 VPB.n107 VNB 0.02fF
C126 VPB.n108 VNB 0.02fF
C127 VPB.n109 VNB 0.02fF
C128 VPB.n110 VNB 0.03fF
C129 VPB.n111 VNB 0.02fF
C130 VPB.n112 VNB 0.19fF
C131 VPB.n113 VNB 0.04fF
C132 VPB.n115 VNB 0.02fF
C133 VPB.n116 VNB 0.02fF
C134 VPB.n117 VNB 0.02fF
C135 VPB.n118 VNB 0.02fF
C136 VPB.n120 VNB 0.02fF
C137 VPB.n121 VNB 0.02fF
C138 VPB.n122 VNB 0.02fF
C139 VPB.n124 VNB 0.26fF
C140 VPB.n126 VNB 0.02fF
C141 VPB.n127 VNB 0.02fF
C142 VPB.n128 VNB 0.10fF
C143 VPB.n129 VNB 0.06fF
C144 VPB.n130 VNB 0.13fF
C145 VPB.n131 VNB 0.15fF
C146 VPB.n132 VNB 0.02fF
C147 VPB.n133 VNB 0.02fF
C148 VPB.n134 VNB 0.13fF
C149 VPB.n135 VNB 0.14fF
C150 VPB.n136 VNB 0.02fF
C151 VPB.n137 VNB 0.02fF
C152 VPB.n138 VNB 0.02fF
C153 VPB.n139 VNB 0.13fF
C154 VPB.n140 VNB 0.14fF
C155 VPB.n141 VNB 0.02fF
C156 VPB.n142 VNB 0.02fF
C157 VPB.n143 VNB 0.13fF
C158 VPB.n144 VNB 0.15fF
C159 VPB.n145 VNB 0.02fF
C160 VPB.n146 VNB 0.02fF
C161 VPB.n147 VNB 0.05fF
C162 VPB.n148 VNB 0.22fF
C163 VPB.n149 VNB 0.02fF
C164 VPB.n150 VNB 0.01fF
C165 VPB.n151 VNB 0.03fF
C166 VPB.n152 VNB 0.26fF
C167 VPB.n153 VNB 0.01fF
C168 VPB.n154 VNB 0.02fF
C169 VPB.n155 VNB 0.03fF
C170 VPB.n156 VNB 0.26fF
C171 VPB.n157 VNB 0.01fF
C172 VPB.n158 VNB 0.02fF
C173 VPB.n159 VNB 0.22fF
C174 VPB.n160 VNB 0.02fF
C175 VPB.n161 VNB 0.02fF
C176 VPB.n162 VNB 0.13fF
C177 VPB.n163 VNB 0.15fF
C178 VPB.n164 VNB 0.02fF
C179 VPB.n165 VNB 0.02fF
C180 VPB.n166 VNB 0.02fF
C181 VPB.n167 VNB 0.02fF
C182 VPB.n168 VNB 0.03fF
C183 VPB.n169 VNB 0.03fF
C184 VPB.n170 VNB 0.02fF
C185 VPB.n171 VNB 0.02fF
C186 VPB.n172 VNB 0.02fF
C187 VPB.n173 VNB 0.02fF
C188 VPB.n174 VNB 0.02fF
C189 VPB.n175 VNB 0.02fF
C190 VPB.n176 VNB 0.03fF
C191 VPB.n177 VNB 0.03fF
C192 VPB.n178 VNB 0.02fF
C193 VPB.n179 VNB 0.02fF
C194 VPB.n180 VNB 0.02fF
C195 VPB.n181 VNB 0.04fF
C196 VPB.n182 VNB 0.03fF
C197 VPB.n184 VNB 0.40fF
C198 a_217_1004.n0 VNB 0.03fF
C199 a_217_1004.n1 VNB 0.43fF
C200 a_217_1004.n2 VNB 0.51fF
C201 a_217_1004.n3 VNB 0.31fF
C202 a_217_1004.n4 VNB 0.35fF
C203 a_217_1004.t7 VNB 0.38fF
C204 a_217_1004.n5 VNB 0.45fF
C205 a_217_1004.n6 VNB 0.49fF
C206 a_217_1004.n7 VNB 0.03fF
C207 a_217_1004.n8 VNB 0.17fF
C208 a_217_1004.n9 VNB 0.04fF
.ends
