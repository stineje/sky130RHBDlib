* SPICE3 file created from DFFSNX1.ext - technology: sky130A

.subckt DFFSNX1 Q QN D CLK SN VDD GND
X0 GND dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X1 QN Q dffsnx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X2 VDD dffsnx1_pcell_0/m1_406_797# QN VDD pshort w=2 l=0.15
X3 VDD Q QN VDD pshort w=2 l=0.15
X4 GND D dffsnx1_pcell_0/nand2x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X5 dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/nand2x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X6 VDD D dffsnx1_pcell_0/m1_537_501# VDD pshort w=2 l=0.15
X7 VDD dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/m1_537_501# VDD pshort w=2 l=0.15
X8 GND dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X9 dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X10 dffsnx1_pcell_0/nand3x1_pcell_0/li_393_182# CLK dffsnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X11 VDD dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/m1_406_797# VDD pshort w=2 l=0.15
X12 VDD CLK dffsnx1_pcell_0/m1_406_797# VDD pshort w=2 l=0.15
X13 VDD dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/m1_406_797# VDD pshort w=2 l=0.15
X14 GND QN dffsnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X15 Q dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X16 dffsnx1_pcell_0/nand3x1_pcell_1/li_393_182# SN dffsnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X17 VDD QN Q VDD pshort w=2 l=0.15
X18 VDD SN Q VDD pshort w=2 l=0.15
X19 VDD dffsnx1_pcell_0/m1_1351_723# Q VDD pshort w=2 l=0.15
X20 GND dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X21 dffsnx1_pcell_0/m1_2461_501# dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/nand3x1_pcell_2/li_393_182# GND nshort w=3 l=0.15
X22 dffsnx1_pcell_0/nand3x1_pcell_2/li_393_182# SN dffsnx1_pcell_0/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X23 VDD dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/m1_2461_501# VDD pshort w=2 l=0.15
X24 VDD SN dffsnx1_pcell_0/m1_2461_501# VDD pshort w=2 l=0.15
X25 VDD dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/m1_2461_501# VDD pshort w=2 l=0.15
X26 GND dffsnx1_pcell_0/m1_2461_501# dffsnx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X27 dffsnx1_pcell_0/m1_1351_723# CLK dffsnx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X28 VDD dffsnx1_pcell_0/m1_2461_501# dffsnx1_pcell_0/m1_1351_723# VDD pshort w=2 l=0.15
X29 VDD CLK dffsnx1_pcell_0/m1_1351_723# VDD pshort w=2 l=0.15
C0 dffsnx1_pcell_0/m1_406_797# CLK 2.36fF
C1 dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/m1_1351_723# 2.89fF
C2 dffsnx1_pcell_0/m1_406_797# VDD 2.24fF
.ends
