magic
tech sky130A
magscale 1 2
timestamp 1654964392
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 5607 945 5641 979
rect 205 871 239 905
rect 427 871 461 905
rect 3535 871 3569 905
rect 4275 871 4309 905
rect 4497 871 4531 905
rect 4645 871 4679 905
rect 5015 871 5049 905
rect 5237 871 5271 905
rect 5607 871 5641 905
rect 205 797 239 831
rect 427 797 461 831
rect 1389 797 1423 831
rect 5607 797 5641 831
rect 205 723 239 757
rect 427 723 461 757
rect 4275 723 4309 757
rect 4497 723 4531 757
rect 5607 723 5641 757
rect 205 649 239 683
rect 427 649 461 683
rect 1389 649 1423 683
rect 3313 649 3347 683
rect 3535 649 3569 683
rect 4275 649 4309 683
rect 4497 649 4531 683
rect 4645 649 4679 683
rect 5015 649 5049 683
rect 5237 649 5271 683
rect 5607 649 5641 683
rect 205 575 239 609
rect 427 575 461 609
rect 2351 575 2385 609
rect 3313 575 3347 609
rect 3535 575 3569 609
rect 4275 575 4309 609
rect 4497 575 4531 609
rect 4645 575 4679 609
rect 5015 575 5049 609
rect 5237 575 5271 609
rect 5607 575 5641 609
rect 205 501 239 535
rect 427 501 461 535
rect 1389 501 1423 535
rect 2351 501 2385 535
rect 5237 501 5271 535
rect 5607 501 5641 535
rect 4497 427 4531 461
rect 4645 427 4679 461
rect 5015 427 5049 461
rect 5607 427 5641 461
<< metal1 >>
rect -34 1446 5806 1514
rect 497 871 3523 905
rect 3605 871 4239 905
rect 1660 797 5490 831
rect 716 723 4024 757
rect 4531 723 5571 757
rect 1459 649 3291 683
rect 4715 649 4989 683
rect 831 576 2174 610
rect 2757 575 3055 609
rect 2421 501 5210 535
rect -34 -34 5806 34
use li1_M1_contact  li1_M1_contact_1 pcells
timestamp 1648061256
transform -1 0 666 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform -1 0 444 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 814 0 -1 593
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_1 pcells
timestamp 1652319931
transform 1 0 962 0 1 0
box -87 -34 1049 1550
use nand3x1_pcell  nand3x1_pcell_0
timestamp 1652319931
transform 1 0 0 0 1 0
box -87 -34 1049 1550
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform -1 0 1627 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform -1 0 1406 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 1184 0 -1 593
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 2146 0 1 593
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform -1 0 1776 0 -1 740
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_2
timestamp 1652319931
transform 1 0 1924 0 1 0
box -87 -34 1049 1550
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform -1 0 2368 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_17
timestamp 1648061256
transform 1 0 3108 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform 1 0 2590 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform 1 0 3330 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform -1 0 2738 0 -1 592
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_3
timestamp 1652319931
transform 1 0 2886 0 1 0
box -87 -34 1049 1550
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform -1 0 3552 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_19
timestamp 1648061256
transform 1 0 4070 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_18
timestamp 1648061256
transform 1 0 4292 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform -1 0 3700 0 -1 814
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_4
timestamp 1652319931
transform 1 0 3848 0 1 0
box -87 -34 1049 1550
use li1_M1_contact  li1_M1_contact_20
timestamp 1648061256
transform 1 0 5476 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_21
timestamp 1648061256
transform 1 0 5032 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_22
timestamp 1648061256
transform 1 0 5254 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform -1 0 4662 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_14
timestamp 1648061256
transform -1 0 4514 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_23
timestamp 1648061256
transform 1 0 5624 0 1 740
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_5
timestamp 1652319931
transform 1 0 4810 0 1 0
box -87 -34 1049 1550
<< labels >>
rlabel locali 5607 723 5641 757 1 Q
port 1 nsew signal output
rlabel locali 5607 797 5641 831 1 Q
port 1 nsew signal output
rlabel locali 5607 871 5641 905 1 Q
port 1 nsew signal output
rlabel locali 5607 945 5641 979 1 Q
port 1 nsew signal output
rlabel locali 5607 649 5641 683 1 Q
port 1 nsew signal output
rlabel locali 5607 575 5641 609 1 Q
port 1 nsew signal output
rlabel locali 5607 501 5641 535 1 Q
port 1 nsew signal output
rlabel locali 5607 427 5641 461 1 Q
port 1 nsew signal output
rlabel locali 4497 427 4531 461 1 Q
port 1 nsew signal output
rlabel locali 4497 575 4531 609 1 Q
port 1 nsew signal output
rlabel locali 4497 649 4531 683 1 Q
port 1 nsew signal output
rlabel locali 4497 723 4531 757 1 Q
port 1 nsew signal output
rlabel locali 4497 871 4531 905 1 Q
port 1 nsew signal output
rlabel locali 4645 649 4679 683 1 QN
port 2 nsew signal output
rlabel locali 4645 871 4679 905 1 QN
port 2 nsew signal output
rlabel locali 4645 575 4679 609 1 QN
port 2 nsew signal output
rlabel locali 4645 427 4679 461 1 QN
port 2 nsew signal output
rlabel locali 5015 427 5049 461 1 QN
port 2 nsew signal output
rlabel locali 5015 575 5049 609 1 QN
port 2 nsew signal output
rlabel locali 5015 649 5049 683 1 QN
port 2 nsew signal output
rlabel locali 5015 871 5049 905 1 QN
port 2 nsew signal output
rlabel locali 205 575 239 609 1 D
port 3 nsew signal input
rlabel locali 205 501 239 535 1 D
port 3 nsew signal input
rlabel locali 205 649 239 683 1 D
port 3 nsew signal input
rlabel locali 205 723 239 757 1 D
port 3 nsew signal input
rlabel locali 205 797 239 831 1 D
port 3 nsew signal input
rlabel locali 205 871 239 905 1 D
port 3 nsew signal input
rlabel locali 1389 649 1423 683 1 CLK
port 4 nsew signal input
rlabel locali 1389 797 1423 831 1 CLK
port 4 nsew signal input
rlabel locali 1389 501 1423 535 1 CLK
port 4 nsew signal input
rlabel locali 3313 575 3347 609 1 CLK
port 4 nsew signal input
rlabel locali 3313 649 3347 683 1 CLK
port 4 nsew signal input
rlabel locali 2351 501 2385 535 1 SN
port 5 nsew signal input
rlabel locali 2351 575 2385 609 1 SN
port 5 nsew signal input
rlabel locali 5237 575 5271 609 1 SN
port 5 nsew signal input
rlabel locali 5237 649 5271 683 1 SN
port 5 nsew signal input
rlabel locali 5237 871 5271 905 1 SN
port 5 nsew signal input
rlabel locali 5237 501 5271 535 1 SN
port 5 nsew signal input
rlabel locali 427 871 461 905 1 RN
port 6 nsew signal input
rlabel locali 427 797 461 831 1 RN
port 6 nsew signal input
rlabel locali 427 723 461 757 1 RN
port 6 nsew signal input
rlabel locali 427 649 461 683 1 RN
port 6 nsew signal input
rlabel locali 427 575 461 609 1 RN
port 6 nsew signal input
rlabel locali 427 501 461 535 1 RN
port 6 nsew signal input
rlabel locali 3535 871 3569 905 1 RN
port 6 nsew signal input
rlabel locali 3535 649 3569 683 1 RN
port 6 nsew signal input
rlabel locali 3535 575 3569 609 1 RN
port 6 nsew signal input
rlabel locali 4275 871 4309 905 1 RN
port 6 nsew signal input
rlabel locali 4275 723 4309 757 1 RN
port 6 nsew signal input
rlabel locali 4275 649 4309 683 1 RN
port 6 nsew signal input
rlabel locali 4275 575 4309 609 1 RN
port 6 nsew signal input
rlabel metal1 -34 1446 5806 1514 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 -34 -34 5806 34 1 GND
port 8 nsew ground bidirectional abutment


<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 5772 1480
string LEFsymmetry X Y R90
<< end >>
