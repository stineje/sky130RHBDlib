// File: or2x1_pcell.spi.pex
// Created: Tue Oct 15 15:59:49 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_OR2X1_PCELL\%noxref_1 ( 11 23 27 35 39 47 53 61 65 76 79 98 110 111 )
c74 ( 111 0 ) capacitor c=0.0600324f //x=3.825 //y=0.37
c75 ( 110 0 ) capacitor c=0.0737024f //x=0.56 //y=0.365
c76 ( 98 0 ) capacitor c=0.0992376f //x=3.33 //y=0
c77 ( 79 0 ) capacitor c=0.202778f //x=0.695 //y=0
c78 ( 76 0 ) capacitor c=0.198211f //x=5.18 //y=0
c79 ( 74 0 ) capacitor c=0.0360689f //x=5.015 //y=0
c80 ( 68 0 ) capacitor c=0.00587411f //x=4.93 //y=0.45
c81 ( 65 0 ) capacitor c=0.00542558f //x=4.845 //y=0.535
c82 ( 64 0 ) capacitor c=0.00479856f //x=4.445 //y=0.45
c83 ( 61 0 ) capacitor c=0.0068422f //x=4.36 //y=0.535
c84 ( 56 0 ) capacitor c=0.00592191f //x=3.96 //y=0.45
c85 ( 53 0 ) capacitor c=0.0164879f //x=3.875 //y=0
c86 ( 48 0 ) capacitor c=0.0659516f //x=2.72 //y=0
c87 ( 47 0 ) capacitor c=0.0195795f //x=3.16 //y=0
c88 ( 42 0 ) capacitor c=0.00609805f //x=2.635 //y=0.445
c89 ( 39 0 ) capacitor c=0.00508468f //x=2.55 //y=0.53
c90 ( 38 0 ) capacitor c=0.00468234f //x=2.15 //y=0.445
c91 ( 35 0 ) capacitor c=0.00556167f //x=2.065 //y=0.53
c92 ( 30 0 ) capacitor c=0.00468234f //x=1.665 //y=0.445
c93 ( 27 0 ) capacitor c=0.00556167f //x=1.58 //y=0.53
c94 ( 26 0 ) capacitor c=0.00468234f //x=1.18 //y=0.445
c95 ( 23 0 ) capacitor c=0.00709092f //x=1.095 //y=0.53
c96 ( 18 0 ) capacitor c=0.00609805f //x=0.695 //y=0.445
c97 ( 11 0 ) capacitor c=0.224767f //x=5.18 //y=0
r98 (  102 103 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.445 //y=0 //x2=4.93 //y2=0
r99 (  101 102 ) resistor r=0.179272 //w=0.357 //l=0.005 //layer=li \
 //thickness=0.1 //x=4.44 //y=0 //x2=4.445 //y2=0
r100 (  99 101 ) resistor r=17.2101 //w=0.357 //l=0.48 //layer=li \
 //thickness=0.1 //x=3.96 //y=0 //x2=4.44 //y2=0
r101 (  86 87 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.15 //y=0 //x2=2.635 //y2=0
r102 (  85 86 ) resistor r=10.7563 //w=0.357 //l=0.3 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.15 //y2=0
r103 (  83 85 ) resistor r=6.63305 //w=0.357 //l=0.185 //layer=li \
 //thickness=0.1 //x=1.665 //y=0 //x2=1.85 //y2=0
r104 (  82 83 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.18 //y=0 //x2=1.665 //y2=0
r105 (  81 82 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.18 //y2=0
r106 (  79 81 ) resistor r=1.61345 //w=0.357 //l=0.045 //layer=li \
 //thickness=0.1 //x=0.695 //y=0 //x2=0.74 //y2=0
r107 (  74 103 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.015 //y=0 //x2=4.93 //y2=0
r108 (  74 76 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=5.015 //y=0 //x2=5.18 //y2=0
r109 (  69 111 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.62 //x2=4.93 //y2=0.535
r110 (  69 111 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.62 //x2=4.93 //y2=1.225
r111 (  68 111 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.45 //x2=4.93 //y2=0.535
r112 (  67 103 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.17 //x2=4.93 //y2=0
r113 (  67 68 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.17 //x2=4.93 //y2=0.45
r114 (  66 111 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.53 //y=0.535 //x2=4.445 //y2=0.535
r115 (  65 111 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.845 //y=0.535 //x2=4.93 //y2=0.535
r116 (  65 66 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=4.845 //y=0.535 //x2=4.53 //y2=0.535
r117 (  64 111 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.445 //y=0.45 //x2=4.445 //y2=0.535
r118 (  63 102 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.445 //y=0.17 //x2=4.445 //y2=0
r119 (  63 64 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=4.445 //y=0.17 //x2=4.445 //y2=0.45
r120 (  62 111 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.045 //y=0.535 //x2=3.96 //y2=0.535
r121 (  61 111 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.36 //y=0.535 //x2=4.445 //y2=0.535
r122 (  61 62 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=4.36 //y=0.535 //x2=4.045 //y2=0.535
r123 (  57 111 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.62 //x2=3.96 //y2=0.535
r124 (  57 111 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.62 //x2=3.96 //y2=1.225
r125 (  56 111 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.45 //x2=3.96 //y2=0.535
r126 (  55 99 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.17 //x2=3.96 //y2=0
r127 (  55 56 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.17 //x2=3.96 //y2=0.45
r128 (  54 98 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.5 //y=0 //x2=3.33 //y2=0
r129 (  53 99 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.875 //y=0 //x2=3.96 //y2=0
r130 (  53 54 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=3.875 //y=0 //x2=3.5 //y2=0
r131 (  48 87 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.72 //y=0 //x2=2.635 //y2=0
r132 (  48 50 ) resistor r=8.60504 //w=0.357 //l=0.24 //layer=li \
 //thickness=0.1 //x=2.72 //y=0 //x2=2.96 //y2=0
r133 (  47 98 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.16 //y=0 //x2=3.33 //y2=0
r134 (  47 50 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=2.96 //y2=0
r135 (  43 110 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.53
r136 (  43 110 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r137 (  42 110 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.445 //x2=2.635 //y2=0.53
r138 (  41 87 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.17 //x2=2.635 //y2=0
r139 (  41 42 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.17 //x2=2.635 //y2=0.445
r140 (  40 110 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.235 //y=0.53 //x2=2.15 //y2=0.53
r141 (  39 110 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.53
r142 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.235 //y2=0.53
r143 (  38 110 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.445 //x2=2.15 //y2=0.53
r144 (  37 86 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.17 //x2=2.15 //y2=0
r145 (  37 38 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.17 //x2=2.15 //y2=0.445
r146 (  36 110 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=1.665 //y2=0.53
r147 (  35 110 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.065 //y=0.53 //x2=2.15 //y2=0.53
r148 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=2.065 //y=0.53 //x2=1.75 //y2=0.53
r149 (  31 110 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.53
r150 (  31 110 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r151 (  30 110 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.445 //x2=1.665 //y2=0.53
r152 (  29 83 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.17 //x2=1.665 //y2=0
r153 (  29 30 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.17 //x2=1.665 //y2=0.445
r154 (  28 110 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0.53 //x2=1.18 //y2=0.53
r155 (  27 110 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.58 //y=0.53 //x2=1.665 //y2=0.53
r156 (  27 28 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.58 //y=0.53 //x2=1.265 //y2=0.53
r157 (  26 110 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.445 //x2=1.18 //y2=0.53
r158 (  25 82 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r159 (  25 26 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.445
r160 (  24 110 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.78 //y=0.53 //x2=0.695 //y2=0.53
r161 (  23 110 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0.53 //x2=1.18 //y2=0.53
r162 (  23 24 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.095 //y=0.53 //x2=0.78 //y2=0.53
r163 (  19 110 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.615 //x2=0.695 //y2=0.53
r164 (  19 110 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.615 //x2=0.695 //y2=1.22
r165 (  18 110 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.445 //x2=0.695 //y2=0.53
r166 (  17 79 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.17 //x2=0.695 //y2=0
r167 (  17 18 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.17 //x2=0.695 //y2=0.445
r168 (  11 76 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.18 //y=0 //x2=5.18 //y2=0
r169 (  9 101 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r170 (  9 11 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.18 //y2=0
r171 (  7 50 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r172 (  7 9 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.44 //y2=0
r173 (  5 85 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r174 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r175 (  2 81 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r176 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
ends PM_OR2X1_PCELL\%noxref_1

subckt PM_OR2X1_PCELL\%noxref_2 ( 11 15 18 25 41 54 58 61 62 63 )
c72 ( 63 0 ) capacitor c=0.0451925f //x=4.74 //y=5.02
c73 ( 62 0 ) capacitor c=0.0423715f //x=3.87 //y=5.02
c74 ( 61 0 ) capacitor c=0.0256796f //x=1.085 //y=5.025
c75 ( 60 0 ) capacitor c=0.00591168f //x=4.885 //y=7.4
c76 ( 59 0 ) capacitor c=0.00591168f //x=4.005 //y=7.4
c77 ( 58 0 ) capacitor c=0.109776f //x=3.33 //y=7.4
c78 ( 57 0 ) capacitor c=0.00591168f //x=1.23 //y=7.4
c79 ( 54 0 ) capacitor c=0.228884f //x=5.18 //y=7.4
c80 ( 41 0 ) capacitor c=0.0287207f //x=4.8 //y=7.4
c81 ( 33 0 ) capacitor c=0.0216067f //x=3.92 //y=7.4
c82 ( 25 0 ) capacitor c=0.0778183f //x=3.16 //y=7.4
c83 ( 18 0 ) capacitor c=0.210107f //x=0.74 //y=7.4
c84 ( 15 0 ) capacitor c=0.0465804f //x=1.145 //y=7.4
c85 ( 11 0 ) capacitor c=0.22902f //x=5.18 //y=7.4
r86 (  52 60 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.97 //y=7.4 //x2=4.885 //y2=7.4
r87 (  52 54 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=4.97 //y=7.4 //x2=5.18 //y2=7.4
r88 (  45 60 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=4.885 //y=7.23 //x2=4.885 //y2=7.4
r89 (  45 63 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=4.885 //y=7.23 //x2=4.885 //y2=6.405
r90 (  42 59 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.09 //y=7.4 //x2=4.005 //y2=7.4
r91 (  42 44 ) resistor r=12.549 //w=0.357 //l=0.35 //layer=li //thickness=0.1 \
 //x=4.09 //y=7.4 //x2=4.44 //y2=7.4
r92 (  41 60 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.8 //y=7.4 //x2=4.885 //y2=7.4
r93 (  41 44 ) resistor r=12.9076 //w=0.357 //l=0.36 //layer=li \
 //thickness=0.1 //x=4.8 //y=7.4 //x2=4.44 //y2=7.4
r94 (  35 59 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=4.005 //y=7.23 //x2=4.005 //y2=7.4
r95 (  35 62 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=4.005 //y=7.23 //x2=4.005 //y2=6.405
r96 (  34 58 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.5 //y=7.4 //x2=3.33 //y2=7.4
r97 (  33 59 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.92 //y=7.4 //x2=4.005 //y2=7.4
r98 (  33 34 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=3.92 //y=7.4 //x2=3.5 //y2=7.4
r99 (  28 30 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r100 (  26 57 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.315 //y=7.4 //x2=1.23 //y2=7.4
r101 (  26 28 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=1.315 //y=7.4 //x2=1.85 //y2=7.4
r102 (  25 58 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.16 //y=7.4 //x2=3.33 //y2=7.4
r103 (  25 30 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=2.96 //y2=7.4
r104 (  19 57 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.23 //y=7.23 //x2=1.23 //y2=7.4
r105 (  19 61 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=1.23 //y=7.23 //x2=1.23 //y2=6.74
r106 (  15 57 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.145 //y=7.4 //x2=1.23 //y2=7.4
r107 (  15 18 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=1.145 //y=7.4 //x2=0.74 //y2=7.4
r108 (  11 54 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.18 //y=7.4 //x2=5.18 //y2=7.4
r109 (  9 44 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r110 (  9 11 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.18 //y2=7.4
r111 (  7 30 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r112 (  7 9 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.44 //y2=7.4
r113 (  5 28 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r114 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r115 (  2 18 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r116 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_OR2X1_PCELL\%noxref_2

subckt PM_OR2X1_PCELL\%noxref_3 ( 1 2 11 12 23 24 25 30 32 40 41 42 43 44 45 \
 46 50 51 52 54 60 61 63 71 72 75 )
c136 ( 75 0 ) capacitor c=0.0159573f //x=1.965 //y=5.025
c137 ( 72 0 ) capacitor c=0.00905936f //x=1.96 //y=0.905
c138 ( 71 0 ) capacitor c=0.007684f //x=0.99 //y=0.905
c139 ( 63 0 ) capacitor c=0.0528806f //x=4.07 //y=2.085
c140 ( 61 0 ) capacitor c=0.0435629f //x=4.71 //y=1.255
c141 ( 60 0 ) capacitor c=0.0200386f //x=4.71 //y=0.91
c142 ( 54 0 ) capacitor c=0.0152946f //x=4.555 //y=1.41
c143 ( 52 0 ) capacitor c=0.0157804f //x=4.555 //y=0.755
c144 ( 51 0 ) capacitor c=0.0524991f //x=4.3 //y=4.79
c145 ( 50 0 ) capacitor c=0.0322983f //x=4.59 //y=4.79
c146 ( 46 0 ) capacitor c=0.0290017f //x=4.18 //y=1.92
c147 ( 45 0 ) capacitor c=0.0250027f //x=4.18 //y=1.565
c148 ( 44 0 ) capacitor c=0.0234316f //x=4.18 //y=1.255
c149 ( 43 0 ) capacitor c=0.0200596f //x=4.18 //y=0.91
c150 ( 42 0 ) capacitor c=0.154218f //x=4.665 //y=6.02
c151 ( 41 0 ) capacitor c=0.154243f //x=4.225 //y=6.02
c152 ( 39 0 ) capacitor c=0.00710337f //x=2.15 //y=1.655
c153 ( 32 0 ) capacitor c=0.0944546f //x=4.07 //y=2.085
c154 ( 30 0 ) capacitor c=0.112871f //x=2.59 //y=3.33
c155 ( 25 0 ) capacitor c=0.0162468f //x=2.505 //y=1.655
c156 ( 24 0 ) capacitor c=0.00499395f //x=2.195 //y=5.21
c157 ( 23 0 ) capacitor c=0.0155365f //x=2.505 //y=5.21
c158 ( 12 0 ) capacitor c=0.00277607f //x=1.265 //y=1.655
c159 ( 11 0 ) capacitor c=0.0280953f //x=2.065 //y=1.655
c160 ( 2 0 ) capacitor c=0.0155913f //x=2.705 //y=3.33
c161 ( 1 0 ) capacitor c=0.0801529f //x=3.955 //y=3.33
r162 (  63 64 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.07 //y=2.085 //x2=4.18 //y2=2.085
r163 (  61 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.71 //y=1.255 //x2=4.67 //y2=1.41
r164 (  60 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.71 //y=0.91 //x2=4.67 //y2=0.755
r165 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.71 //y=0.91 //x2=4.71 //y2=1.255
r166 (  55 68 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.335 //y=1.41 //x2=4.22 //y2=1.41
r167 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.555 //y=1.41 //x2=4.67 //y2=1.41
r168 (  53 67 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.335 //y=0.755 //x2=4.22 //y2=0.755
r169 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.555 //y=0.755 //x2=4.67 //y2=0.755
r170 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.555 //y=0.755 //x2=4.335 //y2=0.755
r171 (  50 57 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.59 //y=4.79 //x2=4.665 //y2=4.865
r172 (  50 51 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=4.59 //y=4.79 //x2=4.3 //y2=4.79
r173 (  47 51 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.225 //y=4.865 //x2=4.3 //y2=4.79
r174 (  47 66 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=4.225 //y=4.865 //x2=4.07 //y2=4.7
r175 (  46 64 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.92 //x2=4.18 //y2=2.085
r176 (  45 68 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.565 //x2=4.22 //y2=1.41
r177 (  45 46 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.565 //x2=4.18 //y2=1.92
r178 (  44 68 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.255 //x2=4.22 //y2=1.41
r179 (  43 67 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.18 //y=0.91 //x2=4.22 //y2=0.755
r180 (  43 44 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.18 //y=0.91 //x2=4.18 //y2=1.255
r181 (  42 57 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.665 //y=6.02 //x2=4.665 //y2=4.865
r182 (  41 47 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.225 //y=6.02 //x2=4.225 //y2=4.865
r183 (  40 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.445 //y=1.41 //x2=4.555 //y2=1.41
r184 (  40 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.445 //y=1.41 //x2=4.335 //y2=1.41
r185 (  37 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.07 //y=4.7 //x2=4.07 //y2=4.7
r186 (  35 37 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=4.07 //y=3.33 //x2=4.07 //y2=4.7
r187 (  32 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.07 //y=2.085 //x2=4.07 //y2=2.085
r188 (  32 35 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=4.07 //y=2.085 //x2=4.07 //y2=3.33
r189 (  28 30 ) resistor r=122.866 //w=0.187 //l=1.795 //layer=li \
 //thickness=0.1 //x=2.59 //y=5.125 //x2=2.59 //y2=3.33
r190 (  27 30 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=2.59 //y=1.74 //x2=2.59 //y2=3.33
r191 (  26 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.235 //y=1.655 //x2=2.15 //y2=1.655
r192 (  25 27 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.59 //y2=1.74
r193 (  25 26 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.235 //y2=1.655
r194 (  23 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.21 //x2=2.59 //y2=5.125
r195 (  23 24 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.21 //x2=2.195 //y2=5.21
r196 (  19 39 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1.655
r197 (  19 72 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r198 (  13 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.295 //x2=2.195 //y2=5.21
r199 (  13 75 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.295 //x2=2.11 //y2=5.72
r200 (  11 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.065 //y=1.655 //x2=2.15 //y2=1.655
r201 (  11 12 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li \
 //thickness=0.1 //x=2.065 //y=1.655 //x2=1.265 //y2=1.655
r202 (  7 12 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.18 //y=1.57 //x2=1.265 //y2=1.655
r203 (  7 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=1.18 //y=1.57 //x2=1.18 //y2=1
r204 (  6 35 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=3.33 //x2=4.07 //y2=3.33
r205 (  4 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.59 //y=3.33 //x2=2.59 //y2=3.33
r206 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.705 //y=3.33 //x2=2.59 //y2=3.33
r207 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.955 //y=3.33 //x2=4.07 //y2=3.33
r208 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=3.955 //y=3.33 //x2=2.705 //y2=3.33
ends PM_OR2X1_PCELL\%noxref_3

subckt PM_OR2X1_PCELL\%noxref_4 ( 3 6 8 9 10 11 12 13 14 18 20 23 25 26 31 )
c66 ( 31 0 ) capacitor c=0.04214f //x=0.955 //y=4.705
c67 ( 26 0 ) capacitor c=0.0321911f //x=1.445 //y=1.25
c68 ( 25 0 ) capacitor c=0.0185201f //x=1.445 //y=0.905
c69 ( 23 0 ) capacitor c=0.0344254f //x=1.375 //y=4.795
c70 ( 20 0 ) capacitor c=0.0133656f //x=1.29 //y=1.405
c71 ( 18 0 ) capacitor c=0.0157804f //x=1.29 //y=0.75
c72 ( 14 0 ) capacitor c=0.0828832f //x=0.915 //y=1.915
c73 ( 13 0 ) capacitor c=0.022867f //x=0.915 //y=1.56
c74 ( 12 0 ) capacitor c=0.0234318f //x=0.915 //y=1.25
c75 ( 11 0 ) capacitor c=0.0192004f //x=0.915 //y=0.905
c76 ( 10 0 ) capacitor c=0.110795f //x=1.45 //y=6.025
c77 ( 9 0 ) capacitor c=0.153847f //x=1.01 //y=6.025
c78 ( 6 0 ) capacitor c=0.00993392f //x=0.955 //y=4.705
c79 ( 3 0 ) capacitor c=0.112424f //x=1.11 //y=2.08
r80 (  33 34 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=0.955 //y=4.795 //x2=0.955 //y2=4.87
r81 (  31 33 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=0.955 //y=4.705 //x2=0.955 //y2=4.795
r82 (  26 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.25 //x2=1.405 //y2=1.405
r83 (  25 39 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.905 //x2=1.405 //y2=0.75
r84 (  25 26 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.905 //x2=1.445 //y2=1.25
r85 (  24 33 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=1.09 //y=4.795 //x2=0.955 //y2=4.795
r86 (  23 27 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.375 //y=4.795 //x2=1.45 //y2=4.87
r87 (  23 24 ) resistor r=146.138 //w=0.094 //l=0.285 //layer=ply \
 //thickness=0.18 //x=1.375 //y=4.795 //x2=1.09 //y2=4.795
r88 (  21 38 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.405 //x2=0.955 //y2=1.405
r89 (  20 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.405 //x2=1.405 //y2=1.405
r90 (  19 37 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.75 //x2=0.955 //y2=0.75
r91 (  18 39 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.75 //x2=1.405 //y2=0.75
r92 (  18 19 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.75 //x2=1.07 //y2=0.75
r93 (  14 36 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r94 (  13 38 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.56 //x2=0.955 //y2=1.405
r95 (  13 14 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.56 //x2=0.915 //y2=1.915
r96 (  12 38 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.25 //x2=0.955 //y2=1.405
r97 (  11 37 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.905 //x2=0.955 //y2=0.75
r98 (  11 12 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.905 //x2=0.915 //y2=1.25
r99 (  10 27 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.025 //x2=1.45 //y2=4.87
r100 (  9 34 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.025 //x2=1.01 //y2=4.87
r101 (  8 20 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.405 //x2=1.29 //y2=1.405
r102 (  8 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.405 //x2=1.07 //y2=1.405
r103 (  6 31 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.955 //y=4.705 //x2=0.955 //y2=4.705
r104 (  6 7 ) resistor r=7.81102 //w=0.254 //l=0.155 //layer=li \
 //thickness=0.1 //x=0.955 //y=4.705 //x2=1.11 //y2=4.705
r105 (  3 36 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r106 (  1 7 ) resistor r=3.23951 //w=0.254 //l=0.165 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.54 //x2=1.11 //y2=4.705
r107 (  1 3 ) resistor r=168.385 //w=0.187 //l=2.46 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.54 //x2=1.11 //y2=2.08
ends PM_OR2X1_PCELL\%noxref_4

subckt PM_OR2X1_PCELL\%noxref_5 ( 1 3 7 8 9 10 11 12 17 19 21 27 28 30 31 34 )
c69 ( 34 0 ) capacitor c=0.0369822f //x=1.885 //y=4.705
c70 ( 31 0 ) capacitor c=0.0279572f //x=1.85 //y=1.915
c71 ( 30 0 ) capacitor c=0.0422144f //x=1.85 //y=2.08
c72 ( 28 0 ) capacitor c=0.0237734f //x=2.415 //y=1.255
c73 ( 27 0 ) capacitor c=0.0191782f //x=2.415 //y=0.905
c74 ( 21 0 ) capacitor c=0.0346941f //x=2.26 //y=1.405
c75 ( 19 0 ) capacitor c=0.0157803f //x=2.26 //y=0.75
c76 ( 17 0 ) capacitor c=0.0360787f //x=2.255 //y=4.795
c77 ( 12 0 ) capacitor c=0.0199921f //x=1.885 //y=1.56
c78 ( 11 0 ) capacitor c=0.0169608f //x=1.885 //y=1.255
c79 ( 10 0 ) capacitor c=0.0185462f //x=1.885 //y=0.905
c80 ( 9 0 ) capacitor c=0.15325f //x=2.33 //y=6.025
c81 ( 8 0 ) capacitor c=0.110232f //x=1.89 //y=6.025
c82 ( 3 0 ) capacitor c=0.0809838f //x=1.85 //y=2.08
c83 ( 1 0 ) capacitor c=0.00521267f //x=1.85 //y=4.54
r84 (  36 37 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.885 //y=4.795 //x2=1.885 //y2=4.87
r85 (  34 36 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.885 //y=4.705 //x2=1.885 //y2=4.795
r86 (  30 31 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r87 (  28 41 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.255 //x2=2.415 //y2=1.367
r88 (  27 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r89 (  27 28 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.255
r90 (  22 39 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r91 (  21 41 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.415 //y2=1.367
r92 (  20 38 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r93 (  19 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r94 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r95 (  18 36 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.02 //y=4.795 //x2=1.885 //y2=4.795
r96 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.795 //x2=2.33 //y2=4.87
r97 (  17 18 ) resistor r=120.5 //w=0.094 //l=0.235 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.795 //x2=2.02 //y2=4.795
r98 (  12 39 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r99 (  12 31 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r100 (  11 39 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.255 //x2=1.925 //y2=1.405
r101 (  10 38 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r102 (  10 11 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.255
r103 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.025 //x2=2.33 //y2=4.87
r104 (  8 37 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.025 //x2=1.89 //y2=4.87
r105 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r106 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r107 (  6 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.885 //y=4.705 //x2=1.885 //y2=4.705
r108 (  3 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r109 (  1 6 ) resistor r=11.332 //w=0.189 //l=0.173292 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.54 //x2=1.867 //y2=4.705
r110 (  1 3 ) resistor r=168.385 //w=0.187 //l=2.46 //layer=li //thickness=0.1 \
 //x=1.85 //y=4.54 //x2=1.85 //y2=2.08
ends PM_OR2X1_PCELL\%noxref_5

subckt PM_OR2X1_PCELL\%noxref_6 ( 7 8 15 16 23 24 25 )
c41 ( 25 0 ) capacitor c=0.030764f //x=2.405 //y=5.025
c42 ( 24 0 ) capacitor c=0.0185379f //x=1.525 //y=5.025
c43 ( 23 0 ) capacitor c=0.0409962f //x=0.655 //y=5.025
c44 ( 16 0 ) capacitor c=0.00193672f //x=1.755 //y=6.91
c45 ( 15 0 ) capacitor c=0.01354f //x=2.465 //y=6.91
c46 ( 8 0 ) capacitor c=0.00844339f //x=0.875 //y=5.21
c47 ( 7 0 ) capacitor c=0.0240359f //x=1.585 //y=5.21
r48 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.55 //y=6.825 //x2=2.55 //y2=6.74
r49 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.465 //y=6.91 //x2=2.55 //y2=6.825
r50 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.465 //y=6.91 //x2=1.755 //y2=6.91
r51 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.67 //y=6.825 //x2=1.755 //y2=6.91
r52 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.67 //y=6.825 //x2=1.67 //y2=6.4
r53 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.67 //y=5.295 //x2=1.67 //y2=5.72
r54 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.585 //y=5.21 //x2=1.67 //y2=5.295
r55 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=1.585 //y=5.21 //x2=0.875 //y2=5.21
r56 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=0.79 //y=5.295 //x2=0.875 //y2=5.21
r57 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=0.79 //y=5.295 //x2=0.79 //y2=5.72
ends PM_OR2X1_PCELL\%noxref_6

subckt PM_OR2X1_PCELL\%noxref_7 ( 11 12 13 14 16 17 19 )
c44 ( 19 0 ) capacitor c=0.028734f //x=4.3 //y=5.02
c45 ( 17 0 ) capacitor c=0.0173218f //x=4.255 //y=0.91
c46 ( 16 0 ) capacitor c=0.105613f //x=4.81 //y=4.495
c47 ( 14 0 ) capacitor c=0.00575887f //x=4.53 //y=4.58
c48 ( 13 0 ) capacitor c=0.0136889f //x=4.725 //y=4.58
c49 ( 12 0 ) capacitor c=0.00636159f //x=4.525 //y=2.08
c50 ( 11 0 ) capacitor c=0.0140707f //x=4.725 //y=2.08
r51 (  15 16 ) resistor r=159.487 //w=0.187 //l=2.33 //layer=li \
 //thickness=0.1 //x=4.81 //y=2.165 //x2=4.81 //y2=4.495
r52 (  13 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=4.58 //x2=4.81 //y2=4.495
r53 (  13 14 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=4.725 //y=4.58 //x2=4.53 //y2=4.58
r54 (  11 15 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=2.08 //x2=4.81 //y2=2.165
r55 (  11 12 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=4.725 //y=2.08 //x2=4.525 //y2=2.08
r56 (  5 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.445 //y=4.665 //x2=4.53 //y2=4.58
r57 (  5 19 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li //thickness=0.1 \
 //x=4.445 //y=4.665 //x2=4.445 //y2=5.725
r58 (  1 12 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.44 //y=1.995 //x2=4.525 //y2=2.08
r59 (  1 17 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=4.44 //y=1.995 //x2=4.44 //y2=1.005
ends PM_OR2X1_PCELL\%noxref_7

