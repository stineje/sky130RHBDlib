magic
tech sky130A
magscale 1 2
timestamp 1652471870
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 3461 945 3495 979
rect 427 871 461 905
rect 2647 871 2681 905
rect 3461 871 3495 905
rect 3831 871 3865 905
rect 427 723 461 757
rect 427 649 461 683
rect 2647 649 2681 683
rect 3461 649 3495 683
rect 3831 649 3865 683
rect 427 575 461 609
rect 1315 575 1349 609
rect 2647 575 2681 609
rect 3461 575 3495 609
rect 3831 575 3865 609
rect 427 501 461 535
rect 1315 501 1349 535
rect 2647 501 2681 535
rect 3461 501 3495 535
rect 3831 501 3865 535
rect 3461 427 3495 461
<< metal1 >>
rect -34 1446 4326 1514
rect 3383 723 4091 757
rect 3531 649 3795 683
rect -34 -34 4326 34
use li1_M1_contact  li1_M1_contact_15 pcells
timestamp 1648061256
transform 1 0 4144 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 3848 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 3478 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform -1 0 3330 0 -1 740
box -53 -33 29 33
use dffx1_pcell  dffx1_pcell_0 pcells
timestamp 1652395794
transform 1 0 0 0 1 0
box -87 -34 4379 1550
<< labels >>
rlabel locali 3831 649 3865 683 1 QN
port 1 nsew signal output
rlabel locali 3831 575 3865 609 1 QN
port 1 nsew signal output
rlabel locali 3831 501 3865 535 1 QN
port 1 nsew signal output
rlabel locali 3831 871 3865 905 1 QN
port 1 nsew signal output
rlabel locali 3461 649 3495 683 1 QN
port 1 nsew signal output
rlabel locali 3461 575 3495 609 1 QN
port 1 nsew signal output
rlabel locali 3461 501 3495 535 1 QN
port 1 nsew signal output
rlabel locali 3461 427 3495 461 1 QN
port 1 nsew signal output
rlabel locali 3461 871 3495 905 1 QN
port 1 nsew signal output
rlabel locali 3461 945 3495 979 1 QN
port 1 nsew signal output
rlabel locali 1315 575 1349 609 1 D
port 2 nsew signal input
rlabel locali 1315 501 1349 535 1 D
port 2 nsew signal input
rlabel locali 427 871 461 905 1 CLK
port 3 nsew signal input
rlabel locali 427 723 461 757 1 CLK
port 3 nsew signal input
rlabel locali 427 649 461 683 1 CLK
port 3 nsew signal input
rlabel locali 427 575 461 609 1 CLK
port 3 nsew signal input
rlabel locali 427 501 461 535 1 CLK
port 3 nsew signal input
rlabel locali 2647 501 2681 535 1 CLK
port 3 nsew signal input
rlabel locali 2647 575 2681 609 1 CLK
port 3 nsew signal input
rlabel locali 2647 649 2681 683 1 CLK
port 3 nsew signal input
rlabel locali 2647 871 2681 905 1 CLK
port 3 nsew signal input
rlabel metal1 -34 1446 4326 1514 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 -34 -34 4326 34 1 GND
port 5 nsew ground bidirectional abutment
<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 4292 1480
string LEFsymmetry X Y R90
<< end >>
