* SPICE3 file created from OR2X1.ext - technology: sky130A

.subckt OR2X1 Y A B VDD GND
X0 a_198_181 A GND GND nshort w=3 l=0.15
X1 Y a_198_181 GND GND nshort w=3 l=0.15
X2 VDD a_198_181 Y VDD pshort w=2 l=0.15 M=2
X3 a_131_1005 A VDD VDD pshort w=2 l=0.15 M=2
X4 a_131_1005 B a_198_181 VDD pshort w=2 l=0.15 M=2
X5 a_198_181 B GND GND nshort w=3 l=0.15
C0 VDD GND 3.03fF
.ends
