* SPICE3 file created from NOR2X1.ext - technology: sky130A

.subckt NOR2X1 Y A B VDD GND
M1000 Y.t3 B.t0 a_131_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 Y A.t0 GND.t0 nshort w=-1.605u l=1.765u
+  ad=0.3582p pd=3.15u as=0p ps=0u
M1002 Y A GND GND nshort w=3u l=0.15u
+  ad=0p pd=0u as=1.9366p ps=12.94u
M1003 Y B.t1 GND.t1 nshort w=-1.83u l=2.06u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_131_1051.t1 A.t1 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B GND GND nshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_131_1051.t2 B.t2 Y.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VDD.t0 A.t2 a_131_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 B VDD 0.07fF
C1 Y VDD 0.25fF
C2 B A 0.26fF
C3 Y A 0.11fF
C4 Y B 0.29fF
C5 A VDD 0.08fF
R0 B.n0 B.t2 470.752
R1 B.n0 B.t0 384.527
R2 B.n1 B.t1 241.172
R3 B.n1 B.n0 110.173
R4 B.n2 B.n1 76
R5 B.n2 B 0.046
R6 a_131_1051.t0 a_131_1051.n0 101.66
R7 a_131_1051.n0 a_131_1051.t2 101.659
R8 a_131_1051.n0 a_131_1051.t3 14.294
R9 a_131_1051.n0 a_131_1051.t1 14.282
R10 Y.n8 Y.n0 164.997
R11 Y.n8 Y.n7 161.848
R12 Y.n7 Y.n6 133.539
R13 Y.n3 Y.n1 80.526
R14 Y.n9 Y.n8 76
R15 Y.n7 Y.n3 48.405
R16 Y.n3 Y.n2 30
R17 Y.n6 Y.n5 22.578
R18 Y.n0 Y.t2 14.282
R19 Y.n0 Y.t3 14.282
R20 Y.n6 Y.n4 8.58
R21 Y.n9 Y 0.046
R22 A.n0 A.t1 486.819
R23 A.n0 A.t2 384.527
R24 A.n1 A.t0 303.607
R25 A.n1 A.n0 79.994
R26 A.n2 A.n1 76
R27 A.n2 A 0.046
R28 GND.n8 GND.n1 76.145
R29 GND.n20 GND.n19 76
R30 GND.n8 GND.n7 76
R31 GND.n14 GND.n13 76
R32 GND.n17 GND.n16 76
R33 GND.n38 GND.n37 76
R34 GND.n32 GND.n31 76
R35 GND.n27 GND.n26 76
R36 GND.n29 GND.n28 19.735
R37 GND.n35 GND.n34 19.735
R38 GND.n12 GND.n11 19.735
R39 GND.n5 GND.n4 19.735
R40 GND.n25 GND.n24 19.735
R41 GND.n11 GND.t1 19.724
R42 GND.n28 GND.t0 19.724
R43 GND.n26 GND.n21 13.653
R44 GND.n31 GND.n30 13.653
R45 GND.n37 GND.n36 13.653
R46 GND.n16 GND.n15 13.653
R47 GND.n13 GND.n9 13.653
R48 GND.n7 GND.n6 13.653
R49 GND.n24 GND.n23 12.837
R50 GND.n4 GND.n3 11.605
R51 GND.n3 GND.n2 9.809
R52 GND.n37 GND.n35 8.854
R53 GND.n23 GND.n22 7.566
R54 GND.t1 GND.n10 7.04
R55 GND.n34 GND.n33 5.774
R56 GND.n13 GND.n12 3.935
R57 GND.n31 GND.n29 3.935
R58 GND.n7 GND.n5 0.983
R59 GND.n26 GND.n25 0.983
R60 GND.n1 GND.n0 0.596
R61 GND.n19 GND.n18 0.596
R62 GND.n20 GND 0.207
R63 GND.n14 GND.n8 0.145
R64 GND.n17 GND.n14 0.145
R65 GND.n38 GND.n32 0.145
R66 GND.n32 GND.n27 0.145
R67 GND.n27 GND.n20 0.145
R68 GND GND.n17 0.09
R69 GND GND.n38 0.09
R70 VDD.n75 VDD.n74 76
R71 VDD.n70 VDD.n69 76
R72 VDD.n63 VDD.n62 76
R73 VDD.n59 VDD.n58 76
R74 VDD.n65 VDD.n64 41.183
R75 VDD.n34 VDD.n33 34.942
R76 VDD.n67 VDD.n66 32.032
R77 VDD.n58 VDD.n55 21.841
R78 VDD.n23 VDD.n20 21.841
R79 VDD.n64 VDD.t1 14.282
R80 VDD.n64 VDD.t0 14.282
R81 VDD.n55 VDD.n37 14.167
R82 VDD.n37 VDD.n36 14.167
R83 VDD.n20 VDD.n19 14.167
R84 VDD.n19 VDD.n17 14.167
R85 VDD.n32 VDD.n29 14.167
R86 VDD.n29 VDD.n28 14.167
R87 VDD.n23 VDD.n22 13.653
R88 VDD.n22 VDD.n21 13.653
R89 VDD.n32 VDD.n31 13.653
R90 VDD.n31 VDD.n30 13.653
R91 VDD.n29 VDD.n25 13.653
R92 VDD.n25 VDD.n24 13.653
R93 VDD.n28 VDD.n27 13.653
R94 VDD.n27 VDD.n26 13.653
R95 VDD.n74 VDD.n73 13.653
R96 VDD.n73 VDD.n72 13.653
R97 VDD.n69 VDD.n68 13.653
R98 VDD.n68 VDD.n67 13.653
R99 VDD.n62 VDD.n61 13.653
R100 VDD.n61 VDD.n60 13.653
R101 VDD.n58 VDD.n57 13.653
R102 VDD.n57 VDD.n56 13.653
R103 VDD.n4 VDD.n2 12.915
R104 VDD.n4 VDD.n3 12.66
R105 VDD.n13 VDD.n12 12.343
R106 VDD.n11 VDD.n10 12.343
R107 VDD.n8 VDD.n7 12.343
R108 VDD.n41 VDD.n40 7.5
R109 VDD.n44 VDD.n43 7.5
R110 VDD.n46 VDD.n45 7.5
R111 VDD.n49 VDD.n48 7.5
R112 VDD.n55 VDD.n54 7.5
R113 VDD.n20 VDD.n16 7.5
R114 VDD.n2 VDD.n1 7.5
R115 VDD.n7 VDD.n6 7.5
R116 VDD.n10 VDD.n9 7.5
R117 VDD.n19 VDD.n18 7.5
R118 VDD.n14 VDD.n0 7.5
R119 VDD.n54 VDD.n53 6.772
R120 VDD.n42 VDD.n39 6.772
R121 VDD.n47 VDD.n44 6.772
R122 VDD.n51 VDD.n49 6.772
R123 VDD.n51 VDD.n50 6.772
R124 VDD.n47 VDD.n46 6.772
R125 VDD.n42 VDD.n41 6.772
R126 VDD.n53 VDD.n38 6.772
R127 VDD.n33 VDD.n23 6.487
R128 VDD.n33 VDD.n32 6.475
R129 VDD.n16 VDD.n15 6.458
R130 VDD.n69 VDD.n65 5.903
R131 VDD.n72 VDD.n71 4.576
R132 VDD.n14 VDD.n5 1.329
R133 VDD.n14 VDD.n8 1.329
R134 VDD.n14 VDD.n11 1.329
R135 VDD.n14 VDD.n13 1.329
R136 VDD.n15 VDD.n14 0.696
R137 VDD.n14 VDD.n4 0.696
R138 VDD.n52 VDD.n51 0.365
R139 VDD.n52 VDD.n47 0.365
R140 VDD.n52 VDD.n42 0.365
R141 VDD.n53 VDD.n52 0.365
R142 VDD.n59 VDD 0.207
R143 VDD.n35 VDD.n34 0.145
R144 VDD.n75 VDD.n70 0.145
R145 VDD.n70 VDD.n63 0.145
R146 VDD.n63 VDD.n59 0.145
R147 VDD VDD.n35 0.09
R148 VDD VDD.n75 0.09
C6 VDD GND 3.27fF
C7 VDD.n0 GND 0.15fF
C8 VDD.n1 GND 0.02fF
C9 VDD.n2 GND 0.02fF
C10 VDD.n3 GND 0.04fF
C11 VDD.n4 GND 0.01fF
C12 VDD.n6 GND 0.02fF
C13 VDD.n7 GND 0.02fF
C14 VDD.n9 GND 0.02fF
C15 VDD.n10 GND 0.02fF
C16 VDD.n12 GND 0.02fF
C17 VDD.n14 GND 0.42fF
C18 VDD.n16 GND 0.03fF
C19 VDD.n17 GND 0.02fF
C20 VDD.n18 GND 0.02fF
C21 VDD.n19 GND 0.02fF
C22 VDD.n20 GND 0.03fF
C23 VDD.n21 GND 0.25fF
C24 VDD.n22 GND 0.02fF
C25 VDD.n23 GND 0.03fF
C26 VDD.n24 GND 0.25fF
C27 VDD.n25 GND 0.01fF
C28 VDD.n26 GND 0.28fF
C29 VDD.n27 GND 0.01fF
C30 VDD.n28 GND 0.02fF
C31 VDD.n29 GND 0.02fF
C32 VDD.n30 GND 0.25fF
C33 VDD.n31 GND 0.01fF
C34 VDD.n32 GND 0.02fF
C35 VDD.n33 GND 0.00fF
C36 VDD.n34 GND 0.08fF
C37 VDD.n35 GND 0.02fF
C38 VDD.n36 GND 0.02fF
C39 VDD.n37 GND 0.02fF
C40 VDD.n38 GND 0.02fF
C41 VDD.n39 GND 0.02fF
C42 VDD.n40 GND 0.02fF
C43 VDD.n41 GND 0.02fF
C44 VDD.n43 GND 0.02fF
C45 VDD.n44 GND 0.02fF
C46 VDD.n45 GND 0.02fF
C47 VDD.n46 GND 0.02fF
C48 VDD.n48 GND 0.03fF
C49 VDD.n49 GND 0.02fF
C50 VDD.n50 GND 0.15fF
C51 VDD.n52 GND 0.42fF
C52 VDD.n54 GND 0.03fF
C53 VDD.n55 GND 0.03fF
C54 VDD.n56 GND 0.25fF
C55 VDD.n57 GND 0.02fF
C56 VDD.n58 GND 0.03fF
C57 VDD.n59 GND 0.03fF
C58 VDD.n60 GND 0.23fF
C59 VDD.n61 GND 0.01fF
C60 VDD.n62 GND 0.02fF
C61 VDD.n63 GND 0.02fF
C62 VDD.n64 GND 0.10fF
C63 VDD.n65 GND 0.02fF
C64 VDD.n66 GND 0.13fF
C65 VDD.n67 GND 0.15fF
C66 VDD.n68 GND 0.01fF
C67 VDD.n69 GND 0.01fF
C68 VDD.n70 GND 0.02fF
C69 VDD.n71 GND 0.16fF
C70 VDD.n72 GND 0.13fF
C71 VDD.n73 GND 0.01fF
C72 VDD.n74 GND 0.02fF
C73 VDD.n75 GND 0.02fF
C74 Y.n0 GND 0.68fF
C75 Y.n1 GND 0.06fF
C76 Y.n2 GND 0.03fF
C77 Y.n3 GND 0.13fF
C78 Y.n4 GND 0.04fF
C79 Y.n5 GND 0.05fF
C80 Y.n6 GND 0.19fF
C81 Y.n7 GND 0.42fF
C82 Y.n8 GND 0.39fF
C83 Y.n9 GND 0.01fF
C84 a_131_1051.n0 GND 0.50fF
.ends
