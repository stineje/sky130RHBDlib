// File: votern3x1_pcell.spi.pex
// Created: Tue Oct 15 16:01:02 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_VOTERN3X1_PCELL\%noxref_1 ( 17 21 24 29 37 43 49 62 66 69 71 72 73 )
c138 ( 73 0 ) capacitor c=0.021507f //x=7.65 //y=0.865
c139 ( 72 0 ) capacitor c=0.021507f //x=4.32 //y=0.865
c140 ( 71 0 ) capacitor c=0.0208055f //x=0.99 //y=0.865
c141 ( 70 0 ) capacitor c=0.00440095f //x=7.84 //y=0
c142 ( 69 0 ) capacitor c=0.101477f //x=6.66 //y=0
c143 ( 68 0 ) capacitor c=0.00440095f //x=4.44 //y=0
c144 ( 66 0 ) capacitor c=0.118054f //x=3.33 //y=0
c145 ( 65 0 ) capacitor c=0.00440095f //x=1.18 //y=0
c146 ( 62 0 ) capacitor c=0.259174f //x=9.25 //y=0
c147 ( 49 0 ) capacitor c=0.0389876f //x=7.755 //y=0
c148 ( 43 0 ) capacitor c=0.0716428f //x=6.49 //y=0
c149 ( 37 0 ) capacitor c=0.0388276f //x=4.425 //y=0
c150 ( 29 0 ) capacitor c=0.0717807f //x=3.16 //y=0
c151 ( 24 0 ) capacitor c=0.177035f //x=0.74 //y=0
c152 ( 21 0 ) capacitor c=0.0422406f //x=1.095 //y=0
c153 ( 17 0 ) capacitor c=0.338433f //x=9.25 //y=0
r154 (  60 62 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=8.14 //y=0 //x2=9.25 //y2=0
r155 (  58 70 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.925 //y=0 //x2=7.84 //y2=0
r156 (  58 60 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=7.925 //y=0 //x2=8.14 //y2=0
r157 (  53 70 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.84 //y=0.17 //x2=7.84 //y2=0
r158 (  53 73 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=7.84 //y=0.17 //x2=7.84 //y2=0.955
r159 (  50 69 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=6.83 //y=0 //x2=6.66 //y2=0
r160 (  50 52 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=6.83 //y=0 //x2=7.03 //y2=0
r161 (  49 70 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.755 //y=0 //x2=7.84 //y2=0
r162 (  49 52 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=7.755 //y=0 //x2=7.03 //y2=0
r163 (  44 68 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.595 //y=0 //x2=4.51 //y2=0
r164 (  44 46 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=4.595 //y=0 //x2=5.55 //y2=0
r165 (  43 69 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=6.49 //y=0 //x2=6.66 //y2=0
r166 (  43 46 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=6.49 //y=0 //x2=5.55 //y2=0
r167 (  39 68 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.51 //y=0.17 //x2=4.51 //y2=0
r168 (  39 72 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=4.51 //y=0.17 //x2=4.51 //y2=0.955
r169 (  38 66 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.5 //y=0 //x2=3.33 //y2=0
r170 (  37 68 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.425 //y=0 //x2=4.51 //y2=0
r171 (  37 38 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=4.425 //y=0 //x2=3.5 //y2=0
r172 (  32 34 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r173 (  30 65 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.18 //y2=0
r174 (  30 32 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.85 //y2=0
r175 (  29 66 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.16 //y=0 //x2=3.33 //y2=0
r176 (  29 34 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=2.96 //y2=0
r177 (  25 65 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r178 (  25 71 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.955
r179 (  21 65 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=1.18 //y2=0
r180 (  21 24 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=0.74 //y2=0
r181 (  17 62 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=0 //x2=9.25 //y2=0
r182 (  15 60 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.14 //y=0 //x2=8.14 //y2=0
r183 (  15 17 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=8.14 //y=0 //x2=9.25 //y2=0
r184 (  13 52 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=0 //x2=7.03 //y2=0
r185 (  13 15 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=0 //x2=8.14 //y2=0
r186 (  11 46 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r187 (  11 13 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=7.03 //y2=0
r188 (  9 68 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r189 (  9 11 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.55 //y2=0
r190 (  7 34 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r191 (  7 9 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.44 //y2=0
r192 (  5 32 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r193 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r194 (  2 24 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r195 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
ends PM_VOTERN3X1_PCELL\%noxref_1

subckt PM_VOTERN3X1_PCELL\%noxref_2 ( 17 29 37 53 68 72 75 76 77 78 79 )
c106 ( 79 0 ) capacitor c=0.0476806f //x=2.405 //y=5.025
c107 ( 78 0 ) capacitor c=0.0241714f //x=1.525 //y=5.025
c108 ( 77 0 ) capacitor c=0.0467094f //x=0.655 //y=5.025
c109 ( 76 0 ) capacitor c=0.11314f //x=6.66 //y=7.4
c110 ( 75 0 ) capacitor c=0.121063f //x=3.33 //y=7.4
c111 ( 74 0 ) capacitor c=0.00591168f //x=2.55 //y=7.4
c112 ( 73 0 ) capacitor c=0.00591168f //x=1.67 //y=7.4
c113 ( 72 0 ) capacitor c=0.245236f //x=0.74 //y=7.4
c114 ( 68 0 ) capacitor c=0.336964f //x=9.25 //y=7.4
c115 ( 53 0 ) capacitor c=0.1275f //x=6.49 //y=7.4
c116 ( 47 0 ) capacitor c=0.0275781f //x=3.16 //y=7.4
c117 ( 37 0 ) capacitor c=0.0292737f //x=2.465 //y=7.4
c118 ( 29 0 ) capacitor c=0.0290962f //x=1.585 //y=7.4
c119 ( 17 0 ) capacitor c=0.382468f //x=9.25 //y=7.4
r120 (  66 68 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=8.14 //y=7.4 //x2=9.25 //y2=7.4
r121 (  64 66 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=7.03 //y=7.4 //x2=8.14 //y2=7.4
r122 (  62 76 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=6.83 //y=7.4 //x2=6.66 //y2=7.4
r123 (  62 64 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=6.83 //y=7.4 //x2=7.03 //y2=7.4
r124 (  56 58 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=4.44 //y=7.4 //x2=5.55 //y2=7.4
r125 (  54 75 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.5 //y=7.4 //x2=3.33 //y2=7.4
r126 (  54 56 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=3.5 //y=7.4 //x2=4.44 //y2=7.4
r127 (  53 76 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=6.49 //y=7.4 //x2=6.66 //y2=7.4
r128 (  53 58 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=6.49 //y=7.4 //x2=5.55 //y2=7.4
r129 (  48 74 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.55 //y2=7.4
r130 (  48 50 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.96 //y2=7.4
r131 (  47 75 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.16 //y=7.4 //x2=3.33 //y2=7.4
r132 (  47 50 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=2.96 //y2=7.4
r133 (  41 74 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=7.4
r134 (  41 79 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=6.4
r135 (  38 73 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.67 //y2=7.4
r136 (  38 40 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.85 //y2=7.4
r137 (  37 74 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=2.55 //y2=7.4
r138 (  37 40 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=1.85 //y2=7.4
r139 (  31 73 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=7.4
r140 (  31 78 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=6.74
r141 (  30 72 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.875 //y=7.4 //x2=0.79 //y2=7.4
r142 (  29 73 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=1.67 //y2=7.4
r143 (  29 30 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=0.875 //y2=7.4
r144 (  23 72 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=7.4
r145 (  23 77 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=6.4
r146 (  17 68 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=7.4 //x2=9.25 //y2=7.4
r147 (  15 66 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.14 //y=7.4 //x2=8.14 //y2=7.4
r148 (  15 17 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=8.14 //y=7.4 //x2=9.25 //y2=7.4
r149 (  13 64 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=7.4 //x2=7.03 //y2=7.4
r150 (  13 15 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=7.4 //x2=8.14 //y2=7.4
r151 (  11 58 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r152 (  11 13 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=7.03 //y2=7.4
r153 (  9 56 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r154 (  9 11 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.55 //y2=7.4
r155 (  7 50 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r156 (  7 9 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.44 //y2=7.4
r157 (  5 40 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r158 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r159 (  2 72 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r160 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_VOTERN3X1_PCELL\%noxref_2

subckt PM_VOTERN3X1_PCELL\%noxref_3 ( 1 2 13 14 15 23 29 30 37 49 50 51 52 53 \
 54 )
c91 ( 54 0 ) capacitor c=0.034295f //x=5.725 //y=5.025
c92 ( 53 0 ) capacitor c=0.0174957f //x=4.845 //y=5.025
c93 ( 51 0 ) capacitor c=0.0214849f //x=1.965 //y=5.025
c94 ( 50 0 ) capacitor c=0.0218033f //x=1.085 //y=5.025
c95 ( 49 0 ) capacitor c=0.00115294f //x=4.99 //y=6.91
c96 ( 37 0 ) capacitor c=0.0131338f //x=5.785 //y=6.91
c97 ( 30 0 ) capacitor c=0.00386507f //x=4.195 //y=6.91
c98 ( 29 0 ) capacitor c=0.0100992f //x=4.905 //y=6.91
c99 ( 23 0 ) capacitor c=0.0453878f //x=4.11 //y=5.21
c100 ( 15 0 ) capacitor c=0.00855201f //x=2.11 //y=5.295
c101 ( 14 0 ) capacitor c=0.00290434f //x=1.315 //y=5.21
c102 ( 13 0 ) capacitor c=0.0150963f //x=2.025 //y=5.21
c103 ( 2 0 ) capacitor c=0.0111402f //x=2.225 //y=5.21
c104 ( 1 0 ) capacitor c=0.0706872f //x=3.995 //y=5.21
r105 (  39 54 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.87 //y=6.825 //x2=5.87 //y2=6.74
r106 (  38 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.075 //y=6.91 //x2=4.99 //y2=6.91
r107 (  37 39 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5.785 //y=6.91 //x2=5.87 //y2=6.825
r108 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=5.785 //y=6.91 //x2=5.075 //y2=6.91
r109 (  31 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.99 //y=6.825 //x2=4.99 //y2=6.91
r110 (  31 53 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.99 //y=6.825 //x2=4.99 //y2=6.74
r111 (  29 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.905 //y=6.91 //x2=4.99 //y2=6.91
r112 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=4.905 //y=6.91 //x2=4.195 //y2=6.91
r113 (  23 52 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=4.11 //y=5.21 //x2=4.11 //y2=6.06
r114 (  21 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.11 //y=6.825 //x2=4.195 //y2=6.91
r115 (  21 52 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.11 //y=6.825 //x2=4.11 //y2=6.74
r116 (  15 48 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.295 //x2=2.11 //y2=5.17
r117 (  15 51 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.295 //x2=2.11 //y2=6.06
r118 (  13 48 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.21 //x2=2.11 //y2=5.17
r119 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.21 //x2=1.315 //y2=5.21
r120 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.295 //x2=1.315 //y2=5.21
r121 (  7 50 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.295 //x2=1.23 //y2=5.72
r122 (  6 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.11 //y=5.21 //x2=4.11 //y2=5.21
r123 (  4 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.11 //y=5.21 //x2=2.11 //y2=5.21
r124 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.225 //y=5.21 //x2=2.11 //y2=5.21
r125 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.995 //y=5.21 //x2=4.11 //y2=5.21
r126 (  1 2 ) resistor r=1.68893 //w=0.131 //l=1.77 //layer=m1 \
 //thickness=0.36 //x=3.995 //y=5.21 //x2=2.225 //y2=5.21
ends PM_VOTERN3X1_PCELL\%noxref_3

subckt PM_VOTERN3X1_PCELL\%noxref_4 ( 1 2 8 16 23 24 25 26 27 28 29 30 31 32 \
 36 38 41 42 43 44 48 49 50 51 55 57 63 64 66 79 )
c153 ( 79 0 ) capacitor c=0.0655948f //x=4.44 //y=4.705
c154 ( 66 0 ) capacitor c=0.0582862f //x=0.74 //y=2.08
c155 ( 64 0 ) capacitor c=0.0342409f //x=4.775 //y=1.21
c156 ( 63 0 ) capacitor c=0.0187384f //x=4.775 //y=0.865
c157 ( 57 0 ) capacitor c=0.0141797f //x=4.62 //y=1.365
c158 ( 55 0 ) capacitor c=0.0149844f //x=4.62 //y=0.71
c159 ( 51 0 ) capacitor c=0.10193f //x=4.245 //y=1.915
c160 ( 50 0 ) capacitor c=0.0225105f //x=4.245 //y=1.52
c161 ( 49 0 ) capacitor c=0.0234376f //x=4.245 //y=1.21
c162 ( 48 0 ) capacitor c=0.0199343f //x=4.245 //y=0.865
c163 ( 44 0 ) capacitor c=0.0318948f //x=1.445 //y=1.21
c164 ( 43 0 ) capacitor c=0.0187384f //x=1.445 //y=0.865
c165 ( 42 0 ) capacitor c=0.0607141f //x=1.085 //y=4.795
c166 ( 41 0 ) capacitor c=0.0292043f //x=1.375 //y=4.795
c167 ( 38 0 ) capacitor c=0.0157913f //x=1.29 //y=1.365
c168 ( 36 0 ) capacitor c=0.0149844f //x=1.29 //y=0.71
c169 ( 32 0 ) capacitor c=0.0302441f //x=0.915 //y=1.915
c170 ( 31 0 ) capacitor c=0.0238107f //x=0.915 //y=1.52
c171 ( 30 0 ) capacitor c=0.0234352f //x=0.915 //y=1.21
c172 ( 29 0 ) capacitor c=0.0199931f //x=0.915 //y=0.865
c173 ( 28 0 ) capacitor c=0.110336f //x=4.77 //y=6.025
c174 ( 27 0 ) capacitor c=0.154049f //x=4.33 //y=6.025
c175 ( 26 0 ) capacitor c=0.110003f //x=1.45 //y=6.025
c176 ( 25 0 ) capacitor c=0.15424f //x=1.01 //y=6.025
c177 ( 16 0 ) capacitor c=0.122411f //x=4.44 //y=2.08
c178 ( 8 0 ) capacitor c=0.12196f //x=0.74 //y=2.08
c179 ( 2 0 ) capacitor c=0.0208472f //x=0.855 //y=4.44
c180 ( 1 0 ) capacitor c=0.119494f //x=4.325 //y=4.44
r181 (  77 79 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.33 //y=4.705 //x2=4.44 //y2=4.705
r182 (  64 81 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.775 //y=1.21 //x2=4.735 //y2=1.365
r183 (  63 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.775 //y=0.865 //x2=4.735 //y2=0.71
r184 (  63 64 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.775 //y=0.865 //x2=4.775 //y2=1.21
r185 (  60 79 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=4.77 //y=4.87 //x2=4.44 //y2=4.705
r186 (  58 76 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.4 //y=1.365 //x2=4.285 //y2=1.365
r187 (  57 81 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.62 //y=1.365 //x2=4.735 //y2=1.365
r188 (  56 75 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.4 //y=0.71 //x2=4.285 //y2=0.71
r189 (  55 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.62 //y=0.71 //x2=4.735 //y2=0.71
r190 (  55 56 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.62 //y=0.71 //x2=4.4 //y2=0.71
r191 (  52 77 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=4.33 //y=4.87 //x2=4.33 //y2=4.705
r192 (  51 74 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=4.245 //y=1.915 //x2=4.44 //y2=2.08
r193 (  50 76 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.245 //y=1.52 //x2=4.285 //y2=1.365
r194 (  50 51 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=4.245 //y=1.52 //x2=4.245 //y2=1.915
r195 (  49 76 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.245 //y=1.21 //x2=4.285 //y2=1.365
r196 (  48 75 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.245 //y=0.865 //x2=4.285 //y2=0.71
r197 (  48 49 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.245 //y=0.865 //x2=4.245 //y2=1.21
r198 (  44 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.21 //x2=1.405 //y2=1.365
r199 (  43 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.405 //y2=0.71
r200 (  43 44 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.445 //y2=1.21
r201 (  41 45 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.375 //y=4.795 //x2=1.45 //y2=4.87
r202 (  41 42 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.375 //y=4.795 //x2=1.085 //y2=4.795
r203 (  39 70 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.365 //x2=0.955 //y2=1.365
r204 (  38 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.365 //x2=1.405 //y2=1.365
r205 (  37 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.71 //x2=0.955 //y2=0.71
r206 (  36 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.405 //y2=0.71
r207 (  36 37 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.07 //y2=0.71
r208 (  33 42 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.87 //x2=1.085 //y2=4.795
r209 (  33 68 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.87 //x2=0.74 //y2=4.705
r210 (  32 66 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=0.74 //y2=2.08
r211 (  31 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.955 //y2=1.365
r212 (  31 32 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.915 //y2=1.915
r213 (  30 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.21 //x2=0.955 //y2=1.365
r214 (  29 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.955 //y2=0.71
r215 (  29 30 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.915 //y2=1.21
r216 (  28 60 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.77 //y=6.025 //x2=4.77 //y2=4.87
r217 (  27 52 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.33 //y=6.025 //x2=4.33 //y2=4.87
r218 (  26 45 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.025 //x2=1.45 //y2=4.87
r219 (  25 33 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.025 //x2=1.01 //y2=4.87
r220 (  24 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.51 //y=1.365 //x2=4.62 //y2=1.365
r221 (  24 58 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.51 //y=1.365 //x2=4.4 //y2=1.365
r222 (  23 38 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.29 //y2=1.365
r223 (  23 39 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.07 //y2=1.365
r224 (  21 79 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=4.705 //x2=4.44 //y2=4.705
r225 (  19 21 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.44 //y=4.44 //x2=4.44 //y2=4.705
r226 (  16 74 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=2.08 //x2=4.44 //y2=2.08
r227 (  16 19 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.08 //x2=4.44 //y2=4.44
r228 (  13 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=4.705 //x2=0.74 //y2=4.705
r229 (  11 13 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=0.74 //y=4.44 //x2=0.74 //y2=4.705
r230 (  8 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=2.08 //x2=0.74 //y2=2.08
r231 (  8 11 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.08 //x2=0.74 //y2=4.44
r232 (  6 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.44 //y=4.44 //x2=4.44 //y2=4.44
r233 (  4 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=0.74 //y=4.44 //x2=0.74 //y2=4.44
r234 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=0.855 //y=4.44 //x2=0.74 //y2=4.44
r235 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.325 //y=4.44 //x2=4.44 //y2=4.44
r236 (  1 2 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=4.325 //y=4.44 //x2=0.855 //y2=4.44
ends PM_VOTERN3X1_PCELL\%noxref_4

subckt PM_VOTERN3X1_PCELL\%noxref_5 ( 1 2 8 15 21 22 23 24 25 26 30 31 32 33 \
 34 36 39 42 43 44 45 46 47 48 49 53 55 58 59 60 61 74 )
c165 ( 74 0 ) capacitor c=0.0583848f //x=7.4 //y=2.08
c166 ( 61 0 ) capacitor c=0.0316774f //x=8.105 //y=1.21
c167 ( 60 0 ) capacitor c=0.0187384f //x=8.105 //y=0.865
c168 ( 59 0 ) capacitor c=0.0590362f //x=7.745 //y=4.795
c169 ( 58 0 ) capacitor c=0.0296075f //x=8.035 //y=4.795
c170 ( 55 0 ) capacitor c=0.0157912f //x=7.95 //y=1.365
c171 ( 53 0 ) capacitor c=0.0149844f //x=7.95 //y=0.71
c172 ( 49 0 ) capacitor c=0.0302441f //x=7.575 //y=1.915
c173 ( 48 0 ) capacitor c=0.0234157f //x=7.575 //y=1.52
c174 ( 47 0 ) capacitor c=0.0234376f //x=7.575 //y=1.21
c175 ( 46 0 ) capacitor c=0.0199931f //x=7.575 //y=0.865
c176 ( 45 0 ) capacitor c=0.0970773f //x=5.745 //y=1.915
c177 ( 44 0 ) capacitor c=0.0249466f //x=5.745 //y=1.56
c178 ( 43 0 ) capacitor c=0.0234397f //x=5.745 //y=1.25
c179 ( 42 0 ) capacitor c=0.0193195f //x=5.745 //y=0.905
c180 ( 39 0 ) capacitor c=0.0631944f //x=5.65 //y=4.87
c181 ( 36 0 ) capacitor c=0.0187941f //x=5.59 //y=1.405
c182 ( 34 0 ) capacitor c=0.0157803f //x=5.59 //y=0.75
c183 ( 33 0 ) capacitor c=0.010629f //x=5.285 //y=4.795
c184 ( 32 0 ) capacitor c=0.0194269f //x=5.575 //y=4.795
c185 ( 31 0 ) capacitor c=0.0365717f //x=5.215 //y=1.25
c186 ( 30 0 ) capacitor c=0.0175988f //x=5.215 //y=0.905
c187 ( 26 0 ) capacitor c=0.110622f //x=8.11 //y=6.025
c188 ( 25 0 ) capacitor c=0.154068f //x=7.67 //y=6.025
c189 ( 24 0 ) capacitor c=0.154291f //x=5.65 //y=6.025
c190 ( 23 0 ) capacitor c=0.110404f //x=5.21 //y=6.025
c191 ( 15 0 ) capacitor c=0.100999f //x=7.4 //y=2.08
c192 ( 8 0 ) capacitor c=0.109253f //x=5.92 //y=2.08
c193 ( 2 0 ) capacitor c=0.011507f //x=6.035 //y=2.08
c194 ( 1 0 ) capacitor c=0.0463146f //x=7.285 //y=2.08
r195 (  61 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.105 //y=1.21 //x2=8.065 //y2=1.365
r196 (  60 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.105 //y=0.865 //x2=8.065 //y2=0.71
r197 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.105 //y=0.865 //x2=8.105 //y2=1.21
r198 (  58 62 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=8.035 //y=4.795 //x2=8.11 //y2=4.87
r199 (  58 59 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=8.035 //y=4.795 //x2=7.745 //y2=4.795
r200 (  56 78 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.73 //y=1.365 //x2=7.615 //y2=1.365
r201 (  55 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.95 //y=1.365 //x2=8.065 //y2=1.365
r202 (  54 77 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.73 //y=0.71 //x2=7.615 //y2=0.71
r203 (  53 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.95 //y=0.71 //x2=8.065 //y2=0.71
r204 (  53 54 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.95 //y=0.71 //x2=7.73 //y2=0.71
r205 (  50 59 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.67 //y=4.87 //x2=7.745 //y2=4.795
r206 (  50 76 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=7.67 //y=4.87 //x2=7.4 //y2=4.705
r207 (  49 74 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=7.575 //y=1.915 //x2=7.4 //y2=2.08
r208 (  48 78 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.575 //y=1.52 //x2=7.615 //y2=1.365
r209 (  48 49 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=7.575 //y=1.52 //x2=7.575 //y2=1.915
r210 (  47 78 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.575 //y=1.21 //x2=7.615 //y2=1.365
r211 (  46 77 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.575 //y=0.865 //x2=7.615 //y2=0.71
r212 (  46 47 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.575 //y=0.865 //x2=7.575 //y2=1.21
r213 (  45 70 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=5.745 //y=1.915 //x2=5.92 //y2=2.08
r214 (  44 68 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.745 //y=1.56 //x2=5.705 //y2=1.405
r215 (  44 45 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=5.745 //y=1.56 //x2=5.745 //y2=1.915
r216 (  43 68 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.745 //y=1.25 //x2=5.705 //y2=1.405
r217 (  42 67 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.745 //y=0.905 //x2=5.705 //y2=0.75
r218 (  42 43 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.745 //y=0.905 //x2=5.745 //y2=1.25
r219 (  39 72 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=5.65 //y=4.87 //x2=5.92 //y2=4.705
r220 (  37 66 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.37 //y=1.405 //x2=5.255 //y2=1.405
r221 (  36 68 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.59 //y=1.405 //x2=5.705 //y2=1.405
r222 (  35 65 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.37 //y=0.75 //x2=5.255 //y2=0.75
r223 (  34 67 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.59 //y=0.75 //x2=5.705 //y2=0.75
r224 (  34 35 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=5.59 //y=0.75 //x2=5.37 //y2=0.75
r225 (  32 39 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.575 //y=4.795 //x2=5.65 //y2=4.87
r226 (  32 33 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=5.575 //y=4.795 //x2=5.285 //y2=4.795
r227 (  31 66 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.215 //y=1.25 //x2=5.255 //y2=1.405
r228 (  30 65 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.215 //y=0.905 //x2=5.255 //y2=0.75
r229 (  30 31 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.215 //y=0.905 //x2=5.215 //y2=1.25
r230 (  27 33 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.21 //y=4.87 //x2=5.285 //y2=4.795
r231 (  26 62 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.11 //y=6.025 //x2=8.11 //y2=4.87
r232 (  25 50 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.67 //y=6.025 //x2=7.67 //y2=4.87
r233 (  24 39 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.65 //y=6.025 //x2=5.65 //y2=4.87
r234 (  23 27 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.21 //y=6.025 //x2=5.21 //y2=4.87
r235 (  22 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.84 //y=1.365 //x2=7.95 //y2=1.365
r236 (  22 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.84 //y=1.365 //x2=7.73 //y2=1.365
r237 (  21 36 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.48 //y=1.405 //x2=5.59 //y2=1.405
r238 (  21 37 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.48 //y=1.405 //x2=5.37 //y2=1.405
r239 (  19 76 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.4 //y=4.705 //x2=7.4 //y2=4.705
r240 (  15 74 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.4 //y=2.08 //x2=7.4 //y2=2.08
r241 (  15 19 ) resistor r=179.679 //w=0.187 //l=2.625 //layer=li \
 //thickness=0.1 //x=7.4 //y=2.08 //x2=7.4 //y2=4.705
r242 (  12 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=4.705 //x2=5.92 //y2=4.705
r243 (  8 70 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=2.08 //x2=5.92 //y2=2.08
r244 (  8 12 ) resistor r=179.679 //w=0.187 //l=2.625 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.08 //x2=5.92 //y2=4.705
r245 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=7.4 \
 //y=2.08 //x2=7.4 //y2=2.08
r246 (  4 8 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=5.92 \
 //y=2.08 //x2=5.92 //y2=2.08
r247 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.035 //y=2.08 //x2=5.92 //y2=2.08
r248 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.285 //y=2.08 //x2=7.4 //y2=2.08
r249 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=7.285 //y=2.08 //x2=6.035 //y2=2.08
ends PM_VOTERN3X1_PCELL\%noxref_5

subckt PM_VOTERN3X1_PCELL\%noxref_6 ( 1 2 13 14 15 21 27 28 35 45 46 47 48 49 \
 50 )
c86 ( 50 0 ) capacitor c=0.0308836f //x=9.065 //y=5.025
c87 ( 49 0 ) capacitor c=0.0173945f //x=8.185 //y=5.025
c88 ( 47 0 ) capacitor c=0.0169278f //x=5.285 //y=5.025
c89 ( 46 0 ) capacitor c=0.0166762f //x=4.405 //y=5.025
c90 ( 45 0 ) capacitor c=0.00115294f //x=8.33 //y=6.91
c91 ( 35 0 ) capacitor c=0.0134683f //x=9.125 //y=6.91
c92 ( 28 0 ) capacitor c=0.00388794f //x=7.535 //y=6.91
c93 ( 27 0 ) capacitor c=0.0107731f //x=8.245 //y=6.91
c94 ( 21 0 ) capacitor c=0.0442221f //x=7.45 //y=5.21
c95 ( 15 0 ) capacitor c=0.0103611f //x=5.43 //y=5.295
c96 ( 14 0 ) capacitor c=0.00227812f //x=4.635 //y=5.21
c97 ( 13 0 ) capacitor c=0.0177888f //x=5.345 //y=5.21
c98 ( 2 0 ) capacitor c=0.00818801f //x=5.545 //y=5.21
c99 ( 1 0 ) capacitor c=0.0820623f //x=7.335 //y=5.21
r100 (  37 50 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.21 //y=6.825 //x2=9.21 //y2=6.74
r101 (  36 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.415 //y=6.91 //x2=8.33 //y2=6.91
r102 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.125 //y=6.91 //x2=9.21 //y2=6.825
r103 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=9.125 //y=6.91 //x2=8.415 //y2=6.91
r104 (  29 45 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.33 //y=6.825 //x2=8.33 //y2=6.91
r105 (  29 49 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.33 //y=6.825 //x2=8.33 //y2=6.74
r106 (  27 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.245 //y=6.91 //x2=8.33 //y2=6.91
r107 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.245 //y=6.91 //x2=7.535 //y2=6.91
r108 (  21 48 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=7.45 //y=5.21 //x2=7.45 //y2=6.06
r109 (  19 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.45 //y=6.825 //x2=7.535 //y2=6.91
r110 (  19 48 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.45 //y=6.825 //x2=7.45 //y2=6.74
r111 (  15 44 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=5.43 //y=5.295 //x2=5.43 //y2=5.17
r112 (  15 47 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=5.43 //y=5.295 //x2=5.43 //y2=6.06
r113 (  13 44 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.345 //y=5.21 //x2=5.43 //y2=5.17
r114 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=5.345 //y=5.21 //x2=4.635 //y2=5.21
r115 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.55 //y=5.295 //x2=4.635 //y2=5.21
r116 (  7 46 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=4.55 //y=5.295 //x2=4.55 //y2=5.72
r117 (  6 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.45 //y=5.21 //x2=7.45 //y2=5.21
r118 (  4 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.43 //y=5.21 //x2=5.43 //y2=5.21
r119 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.545 //y=5.21 //x2=5.43 //y2=5.21
r120 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.335 //y=5.21 //x2=7.45 //y2=5.21
r121 (  1 2 ) resistor r=1.70802 //w=0.131 //l=1.79 //layer=m1 \
 //thickness=0.36 //x=7.335 //y=5.21 //x2=5.545 //y2=5.21
ends PM_VOTERN3X1_PCELL\%noxref_6

subckt PM_VOTERN3X1_PCELL\%noxref_7 ( 1 2 7 9 15 22 25 26 27 28 29 30 31 32 33 \
 38 40 42 48 49 50 51 52 57 59 61 67 68 70 71 74 82 83 86 )
c180 ( 86 0 ) capacitor c=0.0352016f //x=8.53 //y=4.705
c181 ( 83 0 ) capacitor c=0.0279733f //x=8.51 //y=1.915
c182 ( 82 0 ) capacitor c=0.0467621f //x=8.51 //y=2.08
c183 ( 74 0 ) capacitor c=0.0384604f //x=1.89 //y=4.705
c184 ( 71 0 ) capacitor c=0.0300885f //x=1.85 //y=1.915
c185 ( 70 0 ) capacitor c=0.053505f //x=1.85 //y=2.08
c186 ( 68 0 ) capacitor c=0.0237734f //x=9.075 //y=1.255
c187 ( 67 0 ) capacitor c=0.0191782f //x=9.075 //y=0.905
c188 ( 61 0 ) capacitor c=0.0351663f //x=8.92 //y=1.405
c189 ( 59 0 ) capacitor c=0.0157803f //x=8.92 //y=0.75
c190 ( 57 0 ) capacitor c=0.0373879f //x=8.915 //y=4.795
c191 ( 52 0 ) capacitor c=0.0200628f //x=8.545 //y=1.56
c192 ( 51 0 ) capacitor c=0.0168575f //x=8.545 //y=1.255
c193 ( 50 0 ) capacitor c=0.0174993f //x=8.545 //y=0.905
c194 ( 49 0 ) capacitor c=0.0447087f //x=2.415 //y=1.25
c195 ( 48 0 ) capacitor c=0.019286f //x=2.415 //y=0.905
c196 ( 42 0 ) capacitor c=0.0187932f //x=2.26 //y=1.405
c197 ( 40 0 ) capacitor c=0.0157795f //x=2.26 //y=0.75
c198 ( 38 0 ) capacitor c=0.029531f //x=2.255 //y=4.795
c199 ( 33 0 ) capacitor c=0.0206178f //x=1.885 //y=1.56
c200 ( 32 0 ) capacitor c=0.016848f //x=1.885 //y=1.25
c201 ( 31 0 ) capacitor c=0.0174777f //x=1.885 //y=0.905
c202 ( 30 0 ) capacitor c=0.15325f //x=8.99 //y=6.025
c203 ( 29 0 ) capacitor c=0.110411f //x=8.55 //y=6.025
c204 ( 28 0 ) capacitor c=0.154236f //x=2.33 //y=6.025
c205 ( 27 0 ) capacitor c=0.110294f //x=1.89 //y=6.025
c206 ( 22 0 ) capacitor c=0.00501304f //x=8.53 //y=4.705
c207 ( 15 0 ) capacitor c=0.0902071f //x=8.51 //y=2.08
c208 ( 9 0 ) capacitor c=0.11342f //x=1.85 //y=2.08
c209 ( 7 0 ) capacitor c=0.00669947f //x=1.85 //y=4.54
c210 ( 2 0 ) capacitor c=0.0161064f //x=1.965 //y=4.07
c211 ( 1 0 ) capacitor c=0.304963f //x=8.395 //y=4.07
r212 (  88 89 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=8.53 //y=4.795 //x2=8.53 //y2=4.87
r213 (  86 88 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=8.53 //y=4.705 //x2=8.53 //y2=4.795
r214 (  82 83 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=8.51 //y=2.08 //x2=8.51 //y2=1.915
r215 (  74 76 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.89 //y=4.705 //x2=1.89 //y2=4.795
r216 (  70 71 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r217 (  68 93 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=9.075 //y=1.255 //x2=9.075 //y2=1.367
r218 (  67 92 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.075 //y=0.905 //x2=9.035 //y2=0.75
r219 (  67 68 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=9.075 //y=0.905 //x2=9.075 //y2=1.255
r220 (  62 91 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.7 //y=1.405 //x2=8.585 //y2=1.405
r221 (  61 93 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=8.92 //y=1.405 //x2=9.075 //y2=1.367
r222 (  60 90 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.7 //y=0.75 //x2=8.585 //y2=0.75
r223 (  59 92 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.92 //y=0.75 //x2=9.035 //y2=0.75
r224 (  59 60 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=8.92 //y=0.75 //x2=8.7 //y2=0.75
r225 (  58 88 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=8.665 //y=4.795 //x2=8.53 //y2=4.795
r226 (  57 64 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=8.915 //y=4.795 //x2=8.99 //y2=4.87
r227 (  57 58 ) resistor r=128.191 //w=0.094 //l=0.25 //layer=ply \
 //thickness=0.18 //x=8.915 //y=4.795 //x2=8.665 //y2=4.795
r228 (  52 91 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.545 //y=1.56 //x2=8.585 //y2=1.405
r229 (  52 83 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=8.545 //y=1.56 //x2=8.545 //y2=1.915
r230 (  51 91 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=8.545 //y=1.255 //x2=8.585 //y2=1.405
r231 (  50 90 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.545 //y=0.905 //x2=8.585 //y2=0.75
r232 (  50 51 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=8.545 //y=0.905 //x2=8.545 //y2=1.255
r233 (  49 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.25 //x2=2.375 //y2=1.405
r234 (  48 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r235 (  48 49 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.25
r236 (  43 78 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r237 (  42 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.375 //y2=1.405
r238 (  41 77 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r239 (  40 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r240 (  40 41 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r241 (  39 76 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.025 //y=4.795 //x2=1.89 //y2=4.795
r242 (  38 45 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.795 //x2=2.33 //y2=4.87
r243 (  38 39 ) resistor r=117.936 //w=0.094 //l=0.23 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.795 //x2=2.025 //y2=4.795
r244 (  35 76 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.89 //y=4.87 //x2=1.89 //y2=4.795
r245 (  33 78 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r246 (  33 71 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r247 (  32 78 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.25 //x2=1.925 //y2=1.405
r248 (  31 77 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r249 (  31 32 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.25
r250 (  30 64 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.99 //y=6.025 //x2=8.99 //y2=4.87
r251 (  29 89 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.55 //y=6.025 //x2=8.55 //y2=4.87
r252 (  28 45 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.025 //x2=2.33 //y2=4.87
r253 (  27 35 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.025 //x2=1.89 //y2=4.87
r254 (  26 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.81 //y=1.405 //x2=8.92 //y2=1.405
r255 (  26 62 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.81 //y=1.405 //x2=8.7 //y2=1.405
r256 (  25 42 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r257 (  25 43 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r258 (  22 86 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.53 //y=4.705 //x2=8.53 //y2=4.705
r259 (  22 23 ) resistor r=10.3507 //w=0.207 //l=0.165 //layer=li \
 //thickness=0.1 //x=8.52 //y=4.705 //x2=8.52 //y2=4.54
r260 (  20 74 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.89 //y=4.705 //x2=1.89 //y2=4.705
r261 (  18 23 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=8.51 //y=4.07 //x2=8.51 //y2=4.54
r262 (  15 82 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.51 //y=2.08 //x2=8.51 //y2=2.08
r263 (  15 18 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=8.51 //y=2.08 //x2=8.51 //y2=4.07
r264 (  9 70 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r265 (  9 12 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=1.85 //y=2.08 //x2=1.85 //y2=4.07
r266 (  7 20 ) resistor r=11.2426 //w=0.191 //l=0.174714 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.54 //x2=1.87 //y2=4.705
r267 (  7 12 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.54 //x2=1.85 //y2=4.07
r268 (  6 18 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.51 //y=4.07 //x2=8.51 //y2=4.07
r269 (  4 12 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.85 //y=4.07 //x2=1.85 //y2=4.07
r270 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.965 //y=4.07 //x2=1.85 //y2=4.07
r271 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.395 //y=4.07 //x2=8.51 //y2=4.07
r272 (  1 2 ) resistor r=6.1355 //w=0.131 //l=6.43 //layer=m1 //thickness=0.36 \
 //x=8.395 //y=4.07 //x2=1.965 //y2=4.07
ends PM_VOTERN3X1_PCELL\%noxref_7

subckt PM_VOTERN3X1_PCELL\%noxref_8 ( 1 2 3 4 23 24 37 39 40 42 47 48 49 50 54 \
 55 )
c158 ( 55 0 ) capacitor c=0.0167617f //x=8.625 //y=5.025
c159 ( 54 0 ) capacitor c=0.0164812f //x=7.745 //y=5.025
c160 ( 50 0 ) capacitor c=0.0108176f //x=8.62 //y=0.905
c161 ( 49 0 ) capacitor c=0.0131637f //x=5.29 //y=0.905
c162 ( 48 0 ) capacitor c=0.0131367f //x=1.96 //y=0.905
c163 ( 47 0 ) capacitor c=0.00421476f //x=8.77 //y=5.21
c164 ( 42 0 ) capacitor c=0.133261f //x=9.25 //y=5.125
c165 ( 40 0 ) capacitor c=0.00775877f //x=8.895 //y=1.645
c166 ( 39 0 ) capacitor c=0.0165978f //x=9.165 //y=1.645
c167 ( 37 0 ) capacitor c=0.0164794f //x=9.165 //y=5.21
c168 ( 24 0 ) capacitor c=0.0029383f //x=7.975 //y=5.21
c169 ( 23 0 ) capacitor c=0.0159694f //x=8.685 //y=5.21
c170 ( 4 0 ) capacitor c=0.0117447f //x=5.595 //y=1.18
c171 ( 3 0 ) capacitor c=0.0835197f //x=8.695 //y=1.18
c172 ( 2 0 ) capacitor c=0.0203114f //x=2.265 //y=1.18
c173 ( 1 0 ) capacitor c=0.0989941f //x=5.365 //y=1.18
r174 (  46 48 ) resistor r=13.3953 //w=0.172 //l=0.18 //layer=li \
 //thickness=0.1 //x=2.147 //y=1.18 //x2=2.147 //y2=1
r175 (  41 42 ) resistor r=232.385 //w=0.187 //l=3.395 //layer=li \
 //thickness=0.1 //x=9.25 //y=1.73 //x2=9.25 //y2=5.125
r176 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.165 //y=1.645 //x2=9.25 //y2=1.73
r177 (  39 40 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=9.165 //y=1.645 //x2=8.895 //y2=1.645
r178 (  38 47 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.855 //y=5.21 //x2=8.77 //y2=5.21
r179 (  37 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.165 //y=5.21 //x2=9.25 //y2=5.125
r180 (  37 38 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=9.165 //y=5.21 //x2=8.855 //y2=5.21
r181 (  36 50 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=8.81 //y=1.18 //x2=8.81 //y2=1
r182 (  31 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.81 //y=1.56 //x2=8.895 //y2=1.645
r183 (  31 36 ) resistor r=26.0107 //w=0.187 //l=0.38 //layer=li \
 //thickness=0.1 //x=8.81 //y=1.56 //x2=8.81 //y2=1.18
r184 (  25 47 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.77 //y=5.295 //x2=8.77 //y2=5.21
r185 (  25 55 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=8.77 //y=5.295 //x2=8.77 //y2=5.72
r186 (  23 47 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.685 //y=5.21 //x2=8.77 //y2=5.21
r187 (  23 24 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.685 //y=5.21 //x2=7.975 //y2=5.21
r188 (  17 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.89 //y=5.295 //x2=7.975 //y2=5.21
r189 (  17 54 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=7.89 //y=5.295 //x2=7.89 //y2=5.72
r190 (  15 49 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=5.48 //y=1.18 //x2=5.48 //y2=1
r191 (  10 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.81 //y=1.18 //x2=8.81 //y2=1.18
r192 (  8 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.48 //y=1.18 //x2=5.48 //y2=1.18
r193 (  6 46 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.15 //y=1.18 //x2=2.15 //y2=1.18
r194 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.595 //y=1.18 //x2=5.48 //y2=1.18
r195 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.695 //y=1.18 //x2=8.81 //y2=1.18
r196 (  3 4 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=8.695 //y=1.18 //x2=5.595 //y2=1.18
r197 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.265 //y=1.18 //x2=2.15 //y2=1.18
r198 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.365 //y=1.18 //x2=5.48 //y2=1.18
r199 (  1 2 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=5.365 //y=1.18 //x2=2.265 //y2=1.18
ends PM_VOTERN3X1_PCELL\%noxref_8

subckt PM_VOTERN3X1_PCELL\%noxref_9 ( 1 5 9 10 13 17 29 )
c54 ( 29 0 ) capacitor c=0.0790202f //x=0.56 //y=0.365
c55 ( 17 0 ) capacitor c=0.0072249f //x=2.635 //y=0.615
c56 ( 13 0 ) capacitor c=0.0156987f //x=2.55 //y=0.53
c57 ( 10 0 ) capacitor c=0.0104129f //x=1.665 //y=1.495
c58 ( 9 0 ) capacitor c=0.006761f //x=1.665 //y=0.615
c59 ( 5 0 ) capacitor c=0.029726f //x=1.58 //y=1.58
c60 ( 1 0 ) capacitor c=0.00522395f //x=0.695 //y=1.495
r61 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.49
r62 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=1.22
r63 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.75 //y=0.53 //x2=1.665 //y2=0.49
r64 (  14 29 ) resistor r=27.0374 //w=0.187 //l=0.395 //layer=li \
 //thickness=0.1 //x=1.75 //y=0.53 //x2=2.145 //y2=0.53
r65 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.49
r66 (  13 29 ) resistor r=27.7219 //w=0.187 //l=0.405 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.145 //y2=0.53
r67 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=1.62
r68 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=0.88
r69 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.49
r70 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r71 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.78 //y=1.58 //x2=0.695 //y2=1.62
r72 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.78 //y=1.58 //x2=1.18 //y2=1.58
r73 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.58 //y=1.58 //x2=1.665 //y2=1.62
r74 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.58 //y=1.58 //x2=1.18 //y2=1.58
r75 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.695 //y=1.495 //x2=0.695 //y2=1.62
r76 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.695 //y=1.495 //x2=0.695 //y2=0.88
ends PM_VOTERN3X1_PCELL\%noxref_9

subckt PM_VOTERN3X1_PCELL\%noxref_10 ( 1 5 9 10 13 17 29 )
c56 ( 29 0 ) capacitor c=0.0723467f //x=3.89 //y=0.365
c57 ( 17 0 ) capacitor c=0.0072249f //x=5.965 //y=0.615
c58 ( 13 0 ) capacitor c=0.0155051f //x=5.88 //y=0.53
c59 ( 10 0 ) capacitor c=0.0121386f //x=4.995 //y=1.495
c60 ( 9 0 ) capacitor c=0.006761f //x=4.995 //y=0.615
c61 ( 5 0 ) capacitor c=0.0249342f //x=4.91 //y=1.58
c62 ( 1 0 ) capacitor c=0.0107269f //x=4.025 //y=1.495
r63 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=5.965 //y=0.615 //x2=5.965 //y2=0.49
r64 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=5.965 //y=0.615 //x2=5.965 //y2=1.22
r65 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.08 //y=0.53 //x2=4.995 //y2=0.49
r66 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.08 //y=0.53 //x2=5.48 //y2=0.53
r67 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.88 //y=0.53 //x2=5.965 //y2=0.49
r68 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.88 //y=0.53 //x2=5.48 //y2=0.53
r69 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.995 //y=1.495 //x2=4.995 //y2=1.62
r70 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=4.995 //y=1.495 //x2=4.995 //y2=0.88
r71 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=4.995 //y=0.615 //x2=4.995 //y2=0.49
r72 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=4.995 //y=0.615 //x2=4.995 //y2=0.88
r73 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.11 //y=1.58 //x2=4.025 //y2=1.62
r74 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.11 //y=1.58 //x2=4.51 //y2=1.58
r75 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.91 //y=1.58 //x2=4.995 //y2=1.62
r76 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.91 //y=1.58 //x2=4.51 //y2=1.58
r77 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=4.025 //y=1.495 //x2=4.025 //y2=1.62
r78 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=4.025 //y=1.495 //x2=4.025 //y2=0.88
ends PM_VOTERN3X1_PCELL\%noxref_10

subckt PM_VOTERN3X1_PCELL\%noxref_11 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0643762f //x=7.22 //y=0.365
c52 ( 17 0 ) capacitor c=0.00722228f //x=9.295 //y=0.615
c53 ( 13 0 ) capacitor c=0.0141607f //x=9.21 //y=0.53
c54 ( 10 0 ) capacitor c=0.00928228f //x=8.325 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=8.325 //y=0.615
c56 ( 5 0 ) capacitor c=0.0289528f //x=8.24 //y=1.58
c57 ( 1 0 ) capacitor c=0.00481264f //x=7.355 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=9.295 //y=0.615 //x2=9.295 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=9.295 //y=0.615 //x2=9.295 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.41 //y=0.53 //x2=8.325 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.41 //y=0.53 //x2=8.81 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.21 //y=0.53 //x2=9.295 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.21 //y=0.53 //x2=8.81 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=8.325 //y=1.495 //x2=8.325 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=8.325 //y=1.495 //x2=8.325 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=8.325 //y=0.615 //x2=8.325 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=8.325 //y=0.615 //x2=8.325 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.44 //y=1.58 //x2=7.355 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.44 //y=1.58 //x2=7.84 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.24 //y=1.58 //x2=8.325 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.24 //y=1.58 //x2=7.84 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=7.355 //y=1.495 //x2=7.355 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=7.355 //y=1.495 //x2=7.355 //y2=0.88
ends PM_VOTERN3X1_PCELL\%noxref_11

