magic
tech sky130A
magscale 1 2
timestamp 1670281630
<< nwell >>
rect -87 786 975 1550
<< pwell >>
rect -34 -34 922 544
<< nmos >>
rect 155 297 185 350
tri 185 297 201 313 sw
rect 155 267 261 297
tri 261 267 291 297 sw
rect 155 166 185 267
tri 185 251 201 267 nw
tri 245 251 261 267 ne
tri 185 166 201 182 sw
tri 245 166 261 182 se
rect 261 166 291 267
tri 155 136 185 166 ne
rect 185 136 261 166
tri 261 136 291 166 nw
rect 599 297 629 350
tri 629 297 645 313 sw
rect 599 267 705 297
tri 705 267 735 297 sw
rect 599 166 629 267
tri 629 251 645 267 nw
tri 689 251 705 267 ne
tri 629 166 645 182 sw
tri 689 166 705 182 se
rect 705 166 735 267
tri 599 136 629 166 ne
rect 629 136 705 166
tri 705 136 735 166 nw
<< pmos >>
rect 164 1004 194 1404
rect 252 1004 282 1404
rect 608 1004 638 1404
rect 696 1004 726 1404
<< ndiff >>
rect 99 334 155 350
rect 99 300 109 334
rect 143 300 155 334
rect 99 262 155 300
rect 185 334 345 350
rect 185 313 303 334
tri 185 297 201 313 ne
rect 201 300 303 313
rect 337 300 345 334
rect 201 297 345 300
tri 261 267 291 297 ne
rect 99 228 109 262
rect 143 228 155 262
rect 99 194 155 228
rect 99 160 109 194
rect 143 160 155 194
tri 185 251 201 267 se
rect 201 251 245 267
tri 245 251 261 267 sw
rect 185 218 261 251
rect 185 184 205 218
rect 239 184 261 218
rect 185 182 261 184
tri 185 166 201 182 ne
rect 201 166 245 182
tri 245 166 261 182 nw
rect 291 262 345 297
rect 291 228 303 262
rect 337 228 345 262
rect 291 194 345 228
rect 99 136 155 160
tri 155 136 185 166 sw
tri 261 136 291 166 se
rect 291 160 303 194
rect 337 160 345 194
rect 291 136 345 160
rect 99 124 345 136
rect 99 90 109 124
rect 143 90 205 124
rect 239 90 303 124
rect 337 90 345 124
rect 99 74 345 90
rect 543 334 599 350
rect 543 300 553 334
rect 587 300 599 334
rect 543 262 599 300
rect 629 334 789 350
rect 629 313 747 334
tri 629 297 645 313 ne
rect 645 300 747 313
rect 781 300 789 334
rect 645 297 789 300
tri 705 267 735 297 ne
rect 543 228 553 262
rect 587 228 599 262
rect 543 194 599 228
rect 543 160 553 194
rect 587 160 599 194
tri 629 251 645 267 se
rect 645 251 689 267
tri 689 251 705 267 sw
rect 629 218 705 251
rect 629 184 649 218
rect 683 184 705 218
rect 629 182 705 184
tri 629 166 645 182 ne
rect 645 166 689 182
tri 689 166 705 182 nw
rect 735 262 789 297
rect 735 228 747 262
rect 781 228 789 262
rect 735 194 789 228
rect 543 136 599 160
tri 599 136 629 166 sw
tri 705 136 735 166 se
rect 735 160 747 194
rect 781 160 789 194
rect 735 136 789 160
rect 543 124 789 136
rect 543 90 553 124
rect 587 90 649 124
rect 683 90 747 124
rect 781 90 789 124
rect 543 74 789 90
<< pdiff >>
rect 108 1366 164 1404
rect 108 1332 118 1366
rect 152 1332 164 1366
rect 108 1298 164 1332
rect 108 1264 118 1298
rect 152 1264 164 1298
rect 108 1230 164 1264
rect 108 1196 118 1230
rect 152 1196 164 1230
rect 108 1162 164 1196
rect 108 1128 118 1162
rect 152 1128 164 1162
rect 108 1093 164 1128
rect 108 1059 118 1093
rect 152 1059 164 1093
rect 108 1004 164 1059
rect 194 1366 252 1404
rect 194 1332 206 1366
rect 240 1332 252 1366
rect 194 1298 252 1332
rect 194 1264 206 1298
rect 240 1264 252 1298
rect 194 1230 252 1264
rect 194 1196 206 1230
rect 240 1196 252 1230
rect 194 1162 252 1196
rect 194 1128 206 1162
rect 240 1128 252 1162
rect 194 1093 252 1128
rect 194 1059 206 1093
rect 240 1059 252 1093
rect 194 1004 252 1059
rect 282 1366 336 1404
rect 282 1332 294 1366
rect 328 1332 336 1366
rect 282 1298 336 1332
rect 282 1264 294 1298
rect 328 1264 336 1298
rect 282 1230 336 1264
rect 282 1196 294 1230
rect 328 1196 336 1230
rect 282 1162 336 1196
rect 282 1128 294 1162
rect 328 1128 336 1162
rect 282 1093 336 1128
rect 282 1059 294 1093
rect 328 1059 336 1093
rect 282 1004 336 1059
rect 552 1366 608 1404
rect 552 1332 562 1366
rect 596 1332 608 1366
rect 552 1298 608 1332
rect 552 1264 562 1298
rect 596 1264 608 1298
rect 552 1230 608 1264
rect 552 1196 562 1230
rect 596 1196 608 1230
rect 552 1162 608 1196
rect 552 1128 562 1162
rect 596 1128 608 1162
rect 552 1093 608 1128
rect 552 1059 562 1093
rect 596 1059 608 1093
rect 552 1004 608 1059
rect 638 1366 696 1404
rect 638 1332 650 1366
rect 684 1332 696 1366
rect 638 1298 696 1332
rect 638 1264 650 1298
rect 684 1264 696 1298
rect 638 1230 696 1264
rect 638 1196 650 1230
rect 684 1196 696 1230
rect 638 1162 696 1196
rect 638 1128 650 1162
rect 684 1128 696 1162
rect 638 1093 696 1128
rect 638 1059 650 1093
rect 684 1059 696 1093
rect 638 1004 696 1059
rect 726 1366 780 1404
rect 726 1332 738 1366
rect 772 1332 780 1366
rect 726 1298 780 1332
rect 726 1264 738 1298
rect 772 1264 780 1298
rect 726 1230 780 1264
rect 726 1196 738 1230
rect 772 1196 780 1230
rect 726 1162 780 1196
rect 726 1128 738 1162
rect 772 1128 780 1162
rect 726 1093 780 1128
rect 726 1059 738 1093
rect 772 1059 780 1093
rect 726 1004 780 1059
<< ndiffc >>
rect 109 300 143 334
rect 303 300 337 334
rect 109 228 143 262
rect 109 160 143 194
rect 205 184 239 218
rect 303 228 337 262
rect 303 160 337 194
rect 109 90 143 124
rect 205 90 239 124
rect 303 90 337 124
rect 553 300 587 334
rect 747 300 781 334
rect 553 228 587 262
rect 553 160 587 194
rect 649 184 683 218
rect 747 228 781 262
rect 747 160 781 194
rect 553 90 587 124
rect 649 90 683 124
rect 747 90 781 124
<< pdiffc >>
rect 118 1332 152 1366
rect 118 1264 152 1298
rect 118 1196 152 1230
rect 118 1128 152 1162
rect 118 1059 152 1093
rect 206 1332 240 1366
rect 206 1264 240 1298
rect 206 1196 240 1230
rect 206 1128 240 1162
rect 206 1059 240 1093
rect 294 1332 328 1366
rect 294 1264 328 1298
rect 294 1196 328 1230
rect 294 1128 328 1162
rect 294 1059 328 1093
rect 562 1332 596 1366
rect 562 1264 596 1298
rect 562 1196 596 1230
rect 562 1128 596 1162
rect 562 1059 596 1093
rect 650 1332 684 1366
rect 650 1264 684 1298
rect 650 1196 684 1230
rect 650 1128 684 1162
rect 650 1059 684 1093
rect 738 1332 772 1366
rect 738 1264 772 1298
rect 738 1196 772 1230
rect 738 1128 772 1162
rect 738 1059 772 1093
<< psubdiff >>
rect -34 482 922 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 410 461 478 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 410 427 427 461
rect 461 427 478 461
rect 854 461 922 482
rect -34 313 34 353
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect 854 427 871 461
rect 905 427 922 461
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 410 313 478 353
rect 854 387 922 427
rect 854 353 871 387
rect 905 353 922 387
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect -34 17 34 57
rect 410 57 427 91
rect 461 57 478 91
rect 854 313 922 353
rect 854 279 871 313
rect 905 279 922 313
rect 854 239 922 279
rect 854 205 871 239
rect 905 205 922 239
rect 854 165 922 205
rect 854 131 871 165
rect 905 131 922 165
rect 854 91 922 131
rect 410 17 478 57
rect 854 57 871 91
rect 905 57 922 91
rect 854 17 922 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 922 17
rect -34 -34 922 -17
<< nsubdiff >>
rect -34 1497 922 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 922 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 410 1423 478 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 854 1423 922 1463
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 410 979 478 1019
rect 854 1389 871 1423
rect 905 1389 922 1423
rect 854 1349 922 1389
rect 854 1315 871 1349
rect 905 1315 922 1349
rect 854 1275 922 1315
rect 854 1241 871 1275
rect 905 1241 922 1275
rect 854 1201 922 1241
rect 854 1167 871 1201
rect 905 1167 922 1201
rect 854 1127 922 1167
rect 854 1093 871 1127
rect 905 1093 922 1127
rect 854 1053 922 1093
rect 854 1019 871 1053
rect 905 1019 922 1053
rect 410 945 427 979
rect 461 945 478 979
rect -34 871 -17 905
rect 17 884 34 905
rect 410 905 478 945
rect 854 979 922 1019
rect 854 945 871 979
rect 905 945 922 979
rect 410 884 427 905
rect 17 871 427 884
rect 461 884 478 905
rect 854 905 922 945
rect 854 884 871 905
rect 461 871 871 884
rect 905 871 922 905
rect -34 822 922 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 427 427 461 461
rect 427 353 461 387
rect 871 427 905 461
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 871 353 905 387
rect 427 279 461 313
rect 427 205 461 239
rect 427 131 461 165
rect 427 57 461 91
rect 871 279 905 313
rect 871 205 905 239
rect 871 131 905 165
rect 871 57 905 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 427 1389 461 1423
rect 427 1315 461 1349
rect 427 1241 461 1275
rect 427 1167 461 1201
rect 427 1093 461 1127
rect 427 1019 461 1053
rect -17 945 17 979
rect 871 1389 905 1423
rect 871 1315 905 1349
rect 871 1241 905 1275
rect 871 1167 905 1201
rect 871 1093 905 1127
rect 871 1019 905 1053
rect 427 945 461 979
rect -17 871 17 905
rect 871 945 905 979
rect 427 871 461 905
rect 871 871 905 905
<< poly >>
rect 164 1404 194 1430
rect 252 1404 282 1430
rect 608 1404 638 1430
rect 696 1404 726 1430
rect 164 973 194 1004
rect 252 973 282 1004
rect 121 957 282 973
rect 121 923 131 957
rect 165 943 282 957
rect 608 973 638 1004
rect 696 973 726 1004
rect 165 923 175 943
rect 121 907 175 923
rect 565 957 726 973
rect 565 923 575 957
rect 609 943 726 957
rect 609 923 619 943
rect 565 907 619 923
rect 121 434 175 450
rect 121 400 131 434
rect 165 413 175 434
rect 165 400 185 413
rect 121 384 185 400
rect 155 350 185 384
rect 565 434 619 450
rect 565 400 575 434
rect 609 413 619 434
rect 609 400 629 413
rect 565 384 629 400
rect 599 350 629 384
<< polycont >>
rect 131 923 165 957
rect 575 923 609 957
rect 131 400 165 434
rect 575 400 609 434
<< locali >>
rect -34 1497 922 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 922 1497
rect -34 1446 922 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 118 1366 152 1446
rect 118 1298 152 1332
rect 118 1230 152 1264
rect 118 1162 152 1196
rect 118 1093 152 1128
rect 118 1037 152 1059
rect 206 1366 240 1404
rect 206 1298 240 1332
rect 206 1230 240 1264
rect 206 1162 240 1196
rect 206 1093 240 1128
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 131 957 165 973
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 131 434 165 923
rect 206 933 240 1059
rect 294 1366 328 1446
rect 294 1298 328 1332
rect 294 1230 328 1264
rect 294 1162 328 1196
rect 294 1093 328 1128
rect 294 1037 328 1059
rect 410 1423 478 1446
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect 562 1366 596 1446
rect 562 1298 596 1332
rect 562 1230 596 1264
rect 562 1162 596 1196
rect 562 1093 596 1128
rect 562 1037 596 1059
rect 650 1366 684 1404
rect 650 1298 684 1332
rect 650 1230 684 1264
rect 650 1162 684 1196
rect 650 1093 684 1128
rect 410 979 478 1019
rect 410 945 427 979
rect 461 945 478 979
rect 206 899 313 933
rect 279 535 313 899
rect 410 905 478 945
rect 410 871 427 905
rect 461 871 478 905
rect 410 822 478 871
rect 575 957 609 973
rect 279 433 313 501
rect 131 384 165 400
rect 205 399 313 433
rect 410 461 478 544
rect 410 427 427 461
rect 461 427 478 461
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect -34 34 34 57
rect 109 334 143 350
rect 109 262 143 300
rect 109 194 143 228
rect 205 218 239 399
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect 575 535 609 923
rect 650 933 684 1059
rect 738 1366 772 1446
rect 738 1298 772 1332
rect 738 1230 772 1264
rect 738 1162 772 1196
rect 738 1093 772 1128
rect 738 1037 772 1059
rect 854 1423 922 1446
rect 854 1389 871 1423
rect 905 1389 922 1423
rect 854 1349 922 1389
rect 854 1315 871 1349
rect 905 1315 922 1349
rect 854 1275 922 1315
rect 854 1241 871 1275
rect 905 1241 922 1275
rect 854 1201 922 1241
rect 854 1167 871 1201
rect 905 1167 922 1201
rect 854 1127 922 1167
rect 854 1093 871 1127
rect 905 1093 922 1127
rect 854 1053 922 1093
rect 854 1019 871 1053
rect 905 1019 922 1053
rect 854 979 922 1019
rect 854 945 871 979
rect 905 945 922 979
rect 650 899 757 933
rect 575 434 609 501
rect 723 433 757 899
rect 854 905 922 945
rect 854 871 871 905
rect 905 871 922 905
rect 854 822 922 871
rect 575 384 609 400
rect 649 399 757 433
rect 854 461 922 544
rect 854 427 871 461
rect 905 427 922 461
rect 205 168 239 184
rect 303 334 337 350
rect 303 262 337 300
rect 303 194 337 228
rect 109 124 143 160
rect 303 124 337 160
rect 143 90 205 124
rect 239 90 303 124
rect 109 34 143 90
rect 206 34 240 90
rect 303 34 337 90
rect 410 313 478 353
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect 410 57 427 91
rect 461 57 478 91
rect 410 34 478 57
rect 553 334 587 350
rect 553 262 587 300
rect 553 194 587 228
rect 649 218 683 399
rect 854 387 922 427
rect 854 353 871 387
rect 905 353 922 387
rect 649 168 683 184
rect 747 334 781 350
rect 747 262 781 300
rect 747 194 781 228
rect 553 124 587 160
rect 747 124 781 160
rect 587 90 649 124
rect 683 90 747 124
rect 553 34 587 90
rect 650 34 684 90
rect 747 34 781 90
rect 854 313 922 353
rect 854 279 871 313
rect 905 279 922 313
rect 854 239 922 279
rect 854 205 871 239
rect 905 205 922 239
rect 854 165 922 205
rect 854 131 871 165
rect 905 131 922 165
rect 854 91 922 131
rect 854 57 871 91
rect 905 57 922 91
rect 854 34 922 57
rect -34 17 922 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 922 17
rect -34 -34 922 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 279 501 313 535
rect 575 501 609 535
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
<< metal1 >>
rect -34 1497 922 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 922 1497
rect -34 1446 922 1463
rect 273 535 319 541
rect 569 535 615 541
rect 267 501 279 535
rect 313 501 575 535
rect 609 501 621 535
rect 273 495 319 501
rect 569 495 615 501
rect -34 17 922 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 922 17
rect -34 -34 922 -17
<< labels >>
rlabel locali 723 427 757 461 1 Y
port 1 nsew signal output
rlabel locali 723 501 757 535 1 Y
port 1 nsew signal output
rlabel locali 723 575 757 609 1 Y
port 1 nsew signal output
rlabel locali 723 649 757 683 1 Y
port 1 nsew signal output
rlabel locali 723 723 757 757 1 Y
port 1 nsew signal output
rlabel locali 723 797 757 831 1 Y
port 1 nsew signal output
rlabel locali 723 871 757 905 1 Y
port 1 nsew signal output
rlabel locali 131 427 165 461 1 A
port 2 nsew signal input
rlabel locali 131 501 165 535 1 A
port 2 nsew signal input
rlabel locali 131 575 165 609 1 A
port 2 nsew signal input
rlabel locali 131 649 165 683 1 A
port 2 nsew signal input
rlabel locali 131 723 165 757 1 A
port 2 nsew signal input
rlabel locali 131 797 165 831 1 A
port 2 nsew signal input
rlabel locali 131 871 165 905 1 A
port 2 nsew signal input
rlabel metal1 -34 1446 922 1514 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 -34 -34 922 34 1 GND
port 4 nsew ground bidirectional abutment
<< end >>
