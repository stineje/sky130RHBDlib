// File: TMRDFFSNQX1.spi.TMRDFFSNQX1.pxi
// Created: Tue Oct 15 15:52:45 2024
// 
simulator lang=spectre
x_PM_TMRDFFSNQX1\%GND ( GND N_GND_c_24_p N_GND_c_249_p N_GND_c_1_p \
 N_GND_c_25_p N_GND_c_26_p N_GND_c_31_p N_GND_c_32_p N_GND_c_58_p N_GND_c_69_p \
 N_GND_c_76_p N_GND_c_84_p N_GND_c_91_p N_GND_c_98_p N_GND_c_105_p \
 N_GND_c_259_p N_GND_c_266_p N_GND_c_128_p N_GND_c_135_p N_GND_c_138_p \
 N_GND_c_145_p N_GND_c_156_p N_GND_c_163_p N_GND_c_171_p N_GND_c_178_p \
 N_GND_c_188_p N_GND_c_195_p N_GND_c_269_p N_GND_c_276_p N_GND_c_288_p \
 N_GND_c_295_p N_GND_c_298_p N_GND_c_305_p N_GND_c_316_p N_GND_c_323_p \
 N_GND_c_340_p N_GND_c_347_p N_GND_c_354_p N_GND_c_212_p N_GND_c_213_p \
 N_GND_c_451_p N_GND_c_454_p N_GND_c_460_p N_GND_c_476_p N_GND_c_482_p \
 N_GND_c_995_p N_GND_c_511_p N_GND_c_519_p N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p \
 N_GND_c_5_p N_GND_c_6_p N_GND_c_7_p N_GND_c_8_p N_GND_c_9_p N_GND_c_10_p \
 N_GND_c_11_p N_GND_c_12_p N_GND_c_13_p N_GND_c_14_p N_GND_c_15_p N_GND_c_16_p \
 N_GND_c_17_p N_GND_c_18_p N_GND_c_19_p N_GND_c_20_p N_GND_c_21_p N_GND_c_22_p \
 N_GND_c_23_p N_GND_M0_noxref_d N_GND_M2_noxref_d N_GND_M5_noxref_d \
 N_GND_M8_noxref_d N_GND_M10_noxref_d N_GND_M12_noxref_d N_GND_M15_noxref_d \
 N_GND_M17_noxref_d N_GND_M20_noxref_d N_GND_M23_noxref_d N_GND_M25_noxref_d \
 N_GND_M27_noxref_d N_GND_M30_noxref_d N_GND_M32_noxref_d N_GND_M35_noxref_d \
 N_GND_M38_noxref_d N_GND_M40_noxref_d N_GND_M42_noxref_d N_GND_M45_noxref_d \
 N_GND_M47_noxref_d N_GND_M49_noxref_d N_GND_M51_noxref_s )  PM_TMRDFFSNQX1\%GND
x_PM_TMRDFFSNQX1\%VDD ( VDD N_VDD_c_1035_p N_VDD_c_1036_p N_VDD_c_1037_p \
 N_VDD_c_1114_p N_VDD_c_1115_p N_VDD_c_1052_p N_VDD_c_1129_p N_VDD_c_1135_p \
 N_VDD_c_1139_p N_VDD_c_1602_p N_VDD_c_1056_p N_VDD_c_1077_p N_VDD_c_1083_p \
 N_VDD_c_1087_p N_VDD_c_1605_p N_VDD_c_1091_p N_VDD_c_1207_p N_VDD_c_1613_p \
 N_VDD_c_1614_p N_VDD_c_1142_p N_VDD_c_1174_p N_VDD_c_1616_p N_VDD_c_1617_p \
 N_VDD_c_1186_p N_VDD_c_1839_p N_VDD_c_1226_p N_VDD_c_1619_p N_VDD_c_1620_p \
 N_VDD_c_1242_p N_VDD_c_1243_p N_VDD_c_1622_p N_VDD_c_1623_p N_VDD_c_1258_p \
 N_VDD_c_1328_p N_VDD_c_1334_p N_VDD_c_1338_p N_VDD_c_1639_p N_VDD_c_1262_p \
 N_VDD_c_1283_p N_VDD_c_1289_p N_VDD_c_1293_p N_VDD_c_1642_p N_VDD_c_1297_p \
 N_VDD_c_1404_p N_VDD_c_1650_p N_VDD_c_1651_p N_VDD_c_1341_p N_VDD_c_1371_p \
 N_VDD_c_1653_p N_VDD_c_1654_p N_VDD_c_1383_p N_VDD_c_1449_p N_VDD_c_1423_p \
 N_VDD_c_1459_p N_VDD_c_1657_p N_VDD_c_1505_p N_VDD_c_1524_p N_VDD_c_1659_p \
 N_VDD_c_1660_p N_VDD_c_1539_p N_VDD_c_1716_p N_VDD_c_1746_p N_VDD_c_1675_p \
 N_VDD_c_1676_p N_VDD_c_1543_p N_VDD_c_1564_p N_VDD_c_1570_p N_VDD_c_1574_p \
 N_VDD_c_1679_p N_VDD_c_1578_p N_VDD_c_1720_p N_VDD_c_1727_p N_VDD_c_1728_p \
 N_VDD_c_1729_p N_VDD_c_1793_p N_VDD_c_1782_p N_VDD_c_1783_p N_VDD_c_1784_p \
 N_VDD_c_1855_p N_VDD_c_1884_p N_VDD_c_1939_p N_VDD_c_1940_p N_VDD_c_1911_p \
 N_VDD_c_1472_p N_VDD_c_1901_p N_VDD_c_1902_p N_VDD_c_1441_p N_VDD_c_2078_p \
 N_VDD_c_2079_p N_VDD_c_1012_n N_VDD_c_1013_n N_VDD_c_1014_n N_VDD_c_1015_n \
 N_VDD_c_1016_n N_VDD_c_1017_n N_VDD_c_1018_n N_VDD_c_1019_n N_VDD_c_1020_n \
 N_VDD_c_1021_n N_VDD_c_1022_n N_VDD_c_1023_n N_VDD_c_1024_n N_VDD_c_1025_n \
 N_VDD_c_1026_n N_VDD_c_1027_n N_VDD_c_1028_n N_VDD_c_1029_n N_VDD_c_1030_n \
 N_VDD_c_1031_n N_VDD_c_1032_n N_VDD_c_1033_n N_VDD_c_1034_n \
 N_VDD_M52_noxref_s N_VDD_M53_noxref_d N_VDD_M55_noxref_d N_VDD_M56_noxref_s \
 N_VDD_M57_noxref_d N_VDD_M59_noxref_d N_VDD_M61_noxref_d N_VDD_M62_noxref_s \
 N_VDD_M63_noxref_d N_VDD_M65_noxref_d N_VDD_M67_noxref_d N_VDD_M68_noxref_s \
 N_VDD_M69_noxref_d N_VDD_M71_noxref_d N_VDD_M72_noxref_s N_VDD_M73_noxref_d \
 N_VDD_M75_noxref_d N_VDD_M76_noxref_s N_VDD_M77_noxref_d N_VDD_M79_noxref_d \
 N_VDD_M81_noxref_d N_VDD_M82_noxref_s N_VDD_M83_noxref_d N_VDD_M85_noxref_d \
 N_VDD_M86_noxref_s N_VDD_M87_noxref_d N_VDD_M89_noxref_d N_VDD_M91_noxref_d \
 N_VDD_M92_noxref_s N_VDD_M93_noxref_d N_VDD_M95_noxref_d N_VDD_M97_noxref_d \
 N_VDD_M98_noxref_s N_VDD_M99_noxref_d N_VDD_M101_noxref_d N_VDD_M102_noxref_s \
 N_VDD_M103_noxref_d N_VDD_M105_noxref_d N_VDD_M106_noxref_s \
 N_VDD_M107_noxref_d N_VDD_M109_noxref_d N_VDD_M111_noxref_d \
 N_VDD_M112_noxref_s N_VDD_M113_noxref_d N_VDD_M115_noxref_d \
 N_VDD_M116_noxref_s N_VDD_M117_noxref_d N_VDD_M119_noxref_d \
 N_VDD_M121_noxref_d N_VDD_M122_noxref_s N_VDD_M123_noxref_d \
 N_VDD_M125_noxref_d N_VDD_M127_noxref_d N_VDD_M128_noxref_s \
 N_VDD_M129_noxref_d N_VDD_M131_noxref_d N_VDD_M132_noxref_s \
 N_VDD_M133_noxref_d N_VDD_M135_noxref_d N_VDD_M136_noxref_s \
 N_VDD_M137_noxref_d N_VDD_M139_noxref_d N_VDD_M141_noxref_d \
 N_VDD_M142_noxref_s N_VDD_M143_noxref_d N_VDD_M145_noxref_d \
 N_VDD_M154_noxref_s N_VDD_M155_noxref_d )  PM_TMRDFFSNQX1\%VDD
x_PM_TMRDFFSNQX1\%noxref_3 ( N_noxref_3_c_2117_n N_noxref_3_c_2121_n \
 N_noxref_3_c_2123_n N_noxref_3_c_2127_n N_noxref_3_c_2157_n \
 N_noxref_3_c_2161_n N_noxref_3_c_2163_n N_noxref_3_c_2129_n \
 N_noxref_3_c_2259_p N_noxref_3_c_2130_n N_noxref_3_c_2132_n \
 N_noxref_3_c_2133_n N_noxref_3_c_2233_p N_noxref_3_M2_noxref_g \
 N_noxref_3_M5_noxref_g N_noxref_3_M56_noxref_g N_noxref_3_M57_noxref_g \
 N_noxref_3_M62_noxref_g N_noxref_3_M63_noxref_g N_noxref_3_c_2134_n \
 N_noxref_3_c_2136_n N_noxref_3_c_2137_n N_noxref_3_c_2138_n \
 N_noxref_3_c_2139_n N_noxref_3_c_2140_n N_noxref_3_c_2141_n \
 N_noxref_3_c_2143_n N_noxref_3_c_2221_p N_noxref_3_c_2182_n \
 N_noxref_3_c_2144_n N_noxref_3_c_2146_n N_noxref_3_c_2147_n \
 N_noxref_3_c_2148_n N_noxref_3_c_2149_n N_noxref_3_c_2150_n \
 N_noxref_3_c_2151_n N_noxref_3_c_2153_n N_noxref_3_c_2200_p \
 N_noxref_3_c_2184_n N_noxref_3_M1_noxref_d N_noxref_3_M52_noxref_d \
 N_noxref_3_M54_noxref_d )  PM_TMRDFFSNQX1\%noxref_3
x_PM_TMRDFFSNQX1\%noxref_4 ( N_noxref_4_c_2361_n N_noxref_4_c_2362_n \
 N_noxref_4_c_2377_n N_noxref_4_c_2381_n N_noxref_4_c_2383_n \
 N_noxref_4_c_2387_n N_noxref_4_c_2363_n N_noxref_4_c_2495_p \
 N_noxref_4_c_2364_n N_noxref_4_c_2365_n N_noxref_4_c_2505_p \
 N_noxref_4_c_2431_p N_noxref_4_M8_noxref_g N_noxref_4_M68_noxref_g \
 N_noxref_4_M69_noxref_g N_noxref_4_c_2366_n N_noxref_4_c_2368_n \
 N_noxref_4_c_2369_n N_noxref_4_c_2370_n N_noxref_4_c_2371_n \
 N_noxref_4_c_2372_n N_noxref_4_c_2373_n N_noxref_4_c_2375_n \
 N_noxref_4_c_2399_n N_noxref_4_M7_noxref_d N_noxref_4_M62_noxref_d \
 N_noxref_4_M64_noxref_d N_noxref_4_M66_noxref_d )  PM_TMRDFFSNQX1\%noxref_4
x_PM_TMRDFFSNQX1\%noxref_5 ( N_noxref_5_c_2540_n N_noxref_5_c_2547_n \
 N_noxref_5_c_2548_n N_noxref_5_c_2551_n N_noxref_5_c_2608_n \
 N_noxref_5_c_2525_n N_noxref_5_c_2554_n N_noxref_5_c_2558_n \
 N_noxref_5_c_2560_n N_noxref_5_c_2564_n N_noxref_5_c_2527_n \
 N_noxref_5_c_2617_n N_noxref_5_c_2666_p N_noxref_5_c_2528_n \
 N_noxref_5_c_2728_p N_noxref_5_c_2667_p N_noxref_5_c_2571_n \
 N_noxref_5_c_2618_n N_noxref_5_M1_noxref_g N_noxref_5_M10_noxref_g \
 N_noxref_5_M54_noxref_g N_noxref_5_M55_noxref_g N_noxref_5_M72_noxref_g \
 N_noxref_5_M73_noxref_g N_noxref_5_c_2624_n N_noxref_5_c_2625_n \
 N_noxref_5_c_2626_n N_noxref_5_c_2627_n N_noxref_5_c_2629_n \
 N_noxref_5_c_2630_n N_noxref_5_c_2632_n N_noxref_5_c_2633_n \
 N_noxref_5_c_2529_n N_noxref_5_c_2531_n N_noxref_5_c_2532_n \
 N_noxref_5_c_2533_n N_noxref_5_c_2534_n N_noxref_5_c_2535_n \
 N_noxref_5_c_2536_n N_noxref_5_c_2538_n N_noxref_5_c_2635_n \
 N_noxref_5_c_2636_n N_noxref_5_c_2638_n N_noxref_5_c_2581_n \
 N_noxref_5_M4_noxref_d N_noxref_5_M56_noxref_d N_noxref_5_M58_noxref_d \
 N_noxref_5_M60_noxref_d )  PM_TMRDFFSNQX1\%noxref_5
x_PM_TMRDFFSNQX1\%noxref_6 ( N_noxref_6_c_2819_n N_noxref_6_c_2820_n \
 N_noxref_6_c_2821_n N_noxref_6_c_2825_n N_noxref_6_c_2827_n \
 N_noxref_6_c_2803_n N_noxref_6_c_2874_p N_noxref_6_c_2804_n \
 N_noxref_6_c_2805_n N_noxref_6_c_2924_p N_noxref_6_M12_noxref_g \
 N_noxref_6_M76_noxref_g N_noxref_6_M77_noxref_g N_noxref_6_c_2806_n \
 N_noxref_6_c_2808_n N_noxref_6_c_2809_n N_noxref_6_c_2810_n \
 N_noxref_6_c_2811_n N_noxref_6_c_2812_n N_noxref_6_c_2813_n \
 N_noxref_6_c_2815_n N_noxref_6_c_2884_p N_noxref_6_c_2839_n \
 N_noxref_6_M11_noxref_d N_noxref_6_M72_noxref_d N_noxref_6_M74_noxref_d )  \
 PM_TMRDFFSNQX1\%noxref_6
x_PM_TMRDFFSNQX1\%noxref_7 ( N_noxref_7_c_3001_n N_noxref_7_c_3003_n \
 N_noxref_7_c_3009_n N_noxref_7_c_3013_n N_noxref_7_c_3053_n \
 N_noxref_7_c_3055_n N_noxref_7_c_2955_n N_noxref_7_c_2956_n \
 N_noxref_7_c_2965_n N_noxref_7_c_2969_n N_noxref_7_c_2971_n \
 N_noxref_7_c_2957_n N_noxref_7_c_3170_p N_noxref_7_c_2958_n \
 N_noxref_7_c_2959_n N_noxref_7_c_3150_p N_noxref_7_M4_noxref_g \
 N_noxref_7_M7_noxref_g N_noxref_7_M14_noxref_g N_noxref_7_M60_noxref_g \
 N_noxref_7_M61_noxref_g N_noxref_7_M66_noxref_g N_noxref_7_M67_noxref_g \
 N_noxref_7_M80_noxref_g N_noxref_7_M81_noxref_g N_noxref_7_c_3070_n \
 N_noxref_7_c_3071_n N_noxref_7_c_3072_n N_noxref_7_c_3073_n \
 N_noxref_7_c_3074_n N_noxref_7_c_3076_n N_noxref_7_c_3077_n \
 N_noxref_7_c_3028_n N_noxref_7_c_3029_n N_noxref_7_c_3030_n \
 N_noxref_7_c_3031_n N_noxref_7_c_3032_n N_noxref_7_c_3034_n \
 N_noxref_7_c_3035_n N_noxref_7_c_3204_p N_noxref_7_c_3205_p \
 N_noxref_7_c_3206_p N_noxref_7_c_3236_p N_noxref_7_c_3178_p \
 N_noxref_7_c_3238_p N_noxref_7_c_3225_p N_noxref_7_c_3008_n \
 N_noxref_7_c_3080_n N_noxref_7_c_3082_n N_noxref_7_c_3037_n \
 N_noxref_7_c_3038_n N_noxref_7_c_3040_n N_noxref_7_c_3179_p \
 N_noxref_7_c_3209_p N_noxref_7_c_3118_p N_noxref_7_M9_noxref_d \
 N_noxref_7_M68_noxref_d N_noxref_7_M70_noxref_d )  PM_TMRDFFSNQX1\%noxref_7
x_PM_TMRDFFSNQX1\%noxref_8 ( N_noxref_8_c_3277_n N_noxref_8_c_3278_n \
 N_noxref_8_c_3279_n N_noxref_8_c_3280_n N_noxref_8_c_3309_n \
 N_noxref_8_c_3313_n N_noxref_8_c_3315_n N_noxref_8_c_3281_n \
 N_noxref_8_c_3444_p N_noxref_8_c_3282_n N_noxref_8_c_3284_n \
 N_noxref_8_c_3285_n N_noxref_8_c_3378_p N_noxref_8_M17_noxref_g \
 N_noxref_8_M20_noxref_g N_noxref_8_M86_noxref_g N_noxref_8_M87_noxref_g \
 N_noxref_8_M92_noxref_g N_noxref_8_M93_noxref_g N_noxref_8_c_3286_n \
 N_noxref_8_c_3288_n N_noxref_8_c_3289_n N_noxref_8_c_3290_n \
 N_noxref_8_c_3291_n N_noxref_8_c_3292_n N_noxref_8_c_3293_n \
 N_noxref_8_c_3295_n N_noxref_8_c_3367_p N_noxref_8_c_3334_n \
 N_noxref_8_c_3296_n N_noxref_8_c_3298_n N_noxref_8_c_3299_n \
 N_noxref_8_c_3300_n N_noxref_8_c_3301_n N_noxref_8_c_3302_n \
 N_noxref_8_c_3303_n N_noxref_8_c_3305_n N_noxref_8_c_3352_p \
 N_noxref_8_c_3336_n N_noxref_8_M16_noxref_d N_noxref_8_M82_noxref_d \
 N_noxref_8_M84_noxref_d )  PM_TMRDFFSNQX1\%noxref_8
x_PM_TMRDFFSNQX1\%noxref_9 ( N_noxref_9_c_3509_n N_noxref_9_c_3510_n \
 N_noxref_9_c_3525_n N_noxref_9_c_3529_n N_noxref_9_c_3531_n \
 N_noxref_9_c_3535_n N_noxref_9_c_3511_n N_noxref_9_c_3641_p \
 N_noxref_9_c_3512_n N_noxref_9_c_3513_n N_noxref_9_c_3651_p \
 N_noxref_9_c_3577_p N_noxref_9_M23_noxref_g N_noxref_9_M98_noxref_g \
 N_noxref_9_M99_noxref_g N_noxref_9_c_3514_n N_noxref_9_c_3516_n \
 N_noxref_9_c_3517_n N_noxref_9_c_3518_n N_noxref_9_c_3519_n \
 N_noxref_9_c_3520_n N_noxref_9_c_3521_n N_noxref_9_c_3523_n \
 N_noxref_9_c_3547_n N_noxref_9_M22_noxref_d N_noxref_9_M92_noxref_d \
 N_noxref_9_M94_noxref_d N_noxref_9_M96_noxref_d )  PM_TMRDFFSNQX1\%noxref_9
x_PM_TMRDFFSNQX1\%noxref_10 ( N_noxref_10_c_3690_n N_noxref_10_c_3742_n \
 N_noxref_10_c_3691_n N_noxref_10_c_3694_n N_noxref_10_c_3745_n \
 N_noxref_10_c_3675_n N_noxref_10_c_3697_n N_noxref_10_c_3701_n \
 N_noxref_10_c_3703_n N_noxref_10_c_3707_n N_noxref_10_c_3677_n \
 N_noxref_10_c_3912_p N_noxref_10_c_3801_p N_noxref_10_c_3678_n \
 N_noxref_10_c_3891_p N_noxref_10_c_3802_p N_noxref_10_c_3714_n \
 N_noxref_10_c_3754_n N_noxref_10_M16_noxref_g N_noxref_10_M25_noxref_g \
 N_noxref_10_M84_noxref_g N_noxref_10_M85_noxref_g N_noxref_10_M102_noxref_g \
 N_noxref_10_M103_noxref_g N_noxref_10_c_3760_n N_noxref_10_c_3761_n \
 N_noxref_10_c_3762_n N_noxref_10_c_3763_n N_noxref_10_c_3765_n \
 N_noxref_10_c_3766_n N_noxref_10_c_3768_n N_noxref_10_c_3769_n \
 N_noxref_10_c_3679_n N_noxref_10_c_3681_n N_noxref_10_c_3682_n \
 N_noxref_10_c_3683_n N_noxref_10_c_3684_n N_noxref_10_c_3685_n \
 N_noxref_10_c_3686_n N_noxref_10_c_3688_n N_noxref_10_c_3771_n \
 N_noxref_10_c_3772_n N_noxref_10_c_3774_n N_noxref_10_c_3724_n \
 N_noxref_10_M19_noxref_d N_noxref_10_M86_noxref_d N_noxref_10_M88_noxref_d \
 N_noxref_10_M90_noxref_d )  PM_TMRDFFSNQX1\%noxref_10
x_PM_TMRDFFSNQX1\%noxref_11 ( N_noxref_11_c_3956_n N_noxref_11_c_3957_n \
 N_noxref_11_c_3975_n N_noxref_11_c_3979_n N_noxref_11_c_3981_n \
 N_noxref_11_c_3958_n N_noxref_11_c_4061_p N_noxref_11_c_3959_n \
 N_noxref_11_c_3961_n N_noxref_11_c_4037_p N_noxref_11_M27_noxref_g \
 N_noxref_11_M106_noxref_g N_noxref_11_M107_noxref_g N_noxref_11_c_3962_n \
 N_noxref_11_c_3964_n N_noxref_11_c_3965_n N_noxref_11_c_3966_n \
 N_noxref_11_c_3967_n N_noxref_11_c_3968_n N_noxref_11_c_3969_n \
 N_noxref_11_c_3971_n N_noxref_11_c_4028_p N_noxref_11_c_3993_n \
 N_noxref_11_M26_noxref_d N_noxref_11_M102_noxref_d N_noxref_11_M104_noxref_d ) \
 PM_TMRDFFSNQX1\%noxref_11
x_PM_TMRDFFSNQX1\%noxref_12 ( N_noxref_12_c_4157_n N_noxref_12_c_4200_n \
 N_noxref_12_c_4162_n N_noxref_12_c_4164_n N_noxref_12_c_4204_n \
 N_noxref_12_c_4206_n N_noxref_12_c_4111_n N_noxref_12_c_4112_n \
 N_noxref_12_c_4121_n N_noxref_12_c_4125_n N_noxref_12_c_4127_n \
 N_noxref_12_c_4113_n N_noxref_12_c_4345_p N_noxref_12_c_4114_n \
 N_noxref_12_c_4115_n N_noxref_12_c_4327_p N_noxref_12_M19_noxref_g \
 N_noxref_12_M22_noxref_g N_noxref_12_M29_noxref_g N_noxref_12_M90_noxref_g \
 N_noxref_12_M91_noxref_g N_noxref_12_M96_noxref_g N_noxref_12_M97_noxref_g \
 N_noxref_12_M110_noxref_g N_noxref_12_M111_noxref_g N_noxref_12_c_4221_n \
 N_noxref_12_c_4222_n N_noxref_12_c_4223_n N_noxref_12_c_4224_n \
 N_noxref_12_c_4225_n N_noxref_12_c_4227_n N_noxref_12_c_4228_n \
 N_noxref_12_c_4179_n N_noxref_12_c_4180_n N_noxref_12_c_4181_n \
 N_noxref_12_c_4182_n N_noxref_12_c_4183_n N_noxref_12_c_4185_n \
 N_noxref_12_c_4186_n N_noxref_12_c_4258_p N_noxref_12_c_4259_p \
 N_noxref_12_c_4260_p N_noxref_12_c_4261_p N_noxref_12_c_4249_p \
 N_noxref_12_c_4263_p N_noxref_12_c_4250_p N_noxref_12_c_4230_n \
 N_noxref_12_c_4231_n N_noxref_12_c_4233_n N_noxref_12_c_4188_n \
 N_noxref_12_c_4189_n N_noxref_12_c_4191_n N_noxref_12_c_4253_p \
 N_noxref_12_c_4254_p N_noxref_12_c_4248_p N_noxref_12_M24_noxref_d \
 N_noxref_12_M98_noxref_d N_noxref_12_M100_noxref_d )  PM_TMRDFFSNQX1\%noxref_12
x_PM_TMRDFFSNQX1\%noxref_13 ( N_noxref_13_c_4455_n N_noxref_13_c_4513_n \
 N_noxref_13_c_4433_n N_noxref_13_c_4434_n N_noxref_13_c_4602_p \
 N_noxref_13_c_4435_n N_noxref_13_c_4603_p N_noxref_13_c_4444_n \
 N_noxref_13_c_4461_n N_noxref_13_c_4515_n N_noxref_13_c_4445_n \
 N_noxref_13_c_4464_n N_noxref_13_c_4468_n N_noxref_13_c_4470_n \
 N_noxref_13_c_4474_n N_noxref_13_c_4447_n N_noxref_13_c_4658_p \
 N_noxref_13_c_4448_n N_noxref_13_c_4479_n N_noxref_13_c_4449_n \
 N_noxref_13_c_4451_n N_noxref_13_c_4671_p N_noxref_13_c_4587_n \
 N_noxref_13_c_4772_p N_noxref_13_M26_noxref_g N_noxref_13_M46_noxref_g \
 N_noxref_13_M50_noxref_g N_noxref_13_M104_noxref_g N_noxref_13_M105_noxref_g \
 N_noxref_13_M144_noxref_g N_noxref_13_M145_noxref_g N_noxref_13_M152_noxref_g \
 N_noxref_13_M153_noxref_g N_noxref_13_c_4523_n N_noxref_13_c_4526_n \
 N_noxref_13_c_4528_n N_noxref_13_c_4557_n N_noxref_13_c_4559_n \
 N_noxref_13_c_4560_n N_noxref_13_c_4531_n N_noxref_13_c_4532_n \
 N_noxref_13_c_4725_p N_noxref_13_c_4727_p N_noxref_13_c_4728_p \
 N_noxref_13_c_4496_n N_noxref_13_c_4803_p N_noxref_13_c_4804_p \
 N_noxref_13_c_4735_p N_noxref_13_c_4738_p N_noxref_13_c_4768_p \
 N_noxref_13_c_4779_p N_noxref_13_c_4770_p N_noxref_13_c_4830_p \
 N_noxref_13_c_4811_p N_noxref_13_c_4781_p N_noxref_13_c_4778_p \
 N_noxref_13_c_4782_p N_noxref_13_c_4533_n N_noxref_13_c_4566_n \
 N_noxref_13_c_4535_n N_noxref_13_c_4453_n N_noxref_13_c_4888_p \
 N_noxref_13_c_4497_n N_noxref_13_c_4756_p N_noxref_13_c_4826_p \
 N_noxref_13_c_4762_p N_noxref_13_M29_noxref_d N_noxref_13_M106_noxref_d \
 N_noxref_13_M108_noxref_d N_noxref_13_M110_noxref_d )  \
 PM_TMRDFFSNQX1\%noxref_13
x_PM_TMRDFFSNQX1\%D ( N_D_c_4900_n N_D_c_4908_n N_D_c_4909_n N_D_c_5060_n D D \
 D D D D D D D D D D D N_D_c_4915_n N_D_c_4916_n N_D_c_4917_n N_D_M0_noxref_g \
 N_D_M15_noxref_g N_D_M30_noxref_g N_D_M52_noxref_g N_D_M53_noxref_g \
 N_D_M82_noxref_g N_D_M83_noxref_g N_D_M112_noxref_g N_D_M113_noxref_g \
 N_D_c_4918_n N_D_c_4920_n N_D_c_4921_n N_D_c_4922_n N_D_c_4923_n N_D_c_4924_n \
 N_D_c_4925_n N_D_c_4927_n N_D_c_4928_n N_D_c_4930_n N_D_c_4931_n N_D_c_4932_n \
 N_D_c_4933_n N_D_c_4934_n N_D_c_4935_n N_D_c_4937_n N_D_c_4938_n N_D_c_4940_n \
 N_D_c_4941_n N_D_c_4942_n N_D_c_4943_n N_D_c_4944_n N_D_c_4945_n N_D_c_4947_n \
 N_D_c_4971_n N_D_c_4972_n N_D_c_4973_n )  PM_TMRDFFSNQX1\%D
x_PM_TMRDFFSNQX1\%noxref_15 ( N_noxref_15_c_5221_n N_noxref_15_c_5222_n \
 N_noxref_15_c_5223_n N_noxref_15_c_5224_n N_noxref_15_c_5253_n \
 N_noxref_15_c_5257_n N_noxref_15_c_5259_n N_noxref_15_c_5225_n \
 N_noxref_15_c_5389_p N_noxref_15_c_5226_n N_noxref_15_c_5228_n \
 N_noxref_15_c_5229_n N_noxref_15_c_5372_p N_noxref_15_M32_noxref_g \
 N_noxref_15_M35_noxref_g N_noxref_15_M116_noxref_g N_noxref_15_M117_noxref_g \
 N_noxref_15_M122_noxref_g N_noxref_15_M123_noxref_g N_noxref_15_c_5230_n \
 N_noxref_15_c_5232_n N_noxref_15_c_5233_n N_noxref_15_c_5234_n \
 N_noxref_15_c_5235_n N_noxref_15_c_5236_n N_noxref_15_c_5237_n \
 N_noxref_15_c_5239_n N_noxref_15_c_5330_p N_noxref_15_c_5278_n \
 N_noxref_15_c_5240_n N_noxref_15_c_5242_n N_noxref_15_c_5243_n \
 N_noxref_15_c_5244_n N_noxref_15_c_5245_n N_noxref_15_c_5246_n \
 N_noxref_15_c_5247_n N_noxref_15_c_5249_n N_noxref_15_c_5315_p \
 N_noxref_15_c_5280_n N_noxref_15_M31_noxref_d N_noxref_15_M112_noxref_d \
 N_noxref_15_M114_noxref_d )  PM_TMRDFFSNQX1\%noxref_15
x_PM_TMRDFFSNQX1\%noxref_16 ( N_noxref_16_c_5458_n N_noxref_16_c_5459_n \
 N_noxref_16_c_5474_n N_noxref_16_c_5478_n N_noxref_16_c_5480_n \
 N_noxref_16_c_5484_n N_noxref_16_c_5460_n N_noxref_16_c_5555_p \
 N_noxref_16_c_5461_n N_noxref_16_c_5462_n N_noxref_16_c_5565_p \
 N_noxref_16_c_5573_p N_noxref_16_M38_noxref_g N_noxref_16_M128_noxref_g \
 N_noxref_16_M129_noxref_g N_noxref_16_c_5463_n N_noxref_16_c_5465_n \
 N_noxref_16_c_5466_n N_noxref_16_c_5467_n N_noxref_16_c_5468_n \
 N_noxref_16_c_5469_n N_noxref_16_c_5470_n N_noxref_16_c_5472_n \
 N_noxref_16_c_5496_n N_noxref_16_M37_noxref_d N_noxref_16_M122_noxref_d \
 N_noxref_16_M124_noxref_d N_noxref_16_M126_noxref_d )  \
 PM_TMRDFFSNQX1\%noxref_16
x_PM_TMRDFFSNQX1\%CLK ( N_CLK_c_5631_n N_CLK_c_5642_n N_CLK_c_5643_n \
 N_CLK_c_5667_n N_CLK_c_5668_n N_CLK_c_5679_n N_CLK_c_5680_n N_CLK_c_5704_n \
 N_CLK_c_5705_n N_CLK_c_5716_n CLK CLK CLK CLK CLK CLK CLK CLK CLK CLK CLK CLK \
 CLK CLK CLK N_CLK_c_5622_n N_CLK_c_5791_n N_CLK_c_5623_n N_CLK_c_5625_n \
 N_CLK_c_5947_n N_CLK_c_5626_n N_CLK_c_5628_n N_CLK_c_6133_n N_CLK_c_5629_n \
 N_CLK_M3_noxref_g N_CLK_M9_noxref_g N_CLK_M18_noxref_g N_CLK_M24_noxref_g \
 N_CLK_M33_noxref_g N_CLK_M39_noxref_g N_CLK_M58_noxref_g N_CLK_M59_noxref_g \
 N_CLK_M70_noxref_g N_CLK_M71_noxref_g N_CLK_M88_noxref_g N_CLK_M89_noxref_g \
 N_CLK_M100_noxref_g N_CLK_M101_noxref_g N_CLK_M118_noxref_g \
 N_CLK_M119_noxref_g N_CLK_M130_noxref_g N_CLK_M131_noxref_g N_CLK_c_5769_n \
 N_CLK_c_5772_n N_CLK_c_6298_p N_CLK_c_6305_p N_CLK_c_5774_n N_CLK_c_5775_n \
 N_CLK_c_5776_n N_CLK_c_5777_n N_CLK_c_5837_n N_CLK_c_5800_n N_CLK_c_5803_n \
 N_CLK_c_5805_n N_CLK_c_5893_n N_CLK_c_5895_n N_CLK_c_5896_n N_CLK_c_5808_n \
 N_CLK_c_5809_n N_CLK_c_5926_n N_CLK_c_5929_n N_CLK_c_6327_p N_CLK_c_6334_p \
 N_CLK_c_5931_n N_CLK_c_5932_n N_CLK_c_5933_n N_CLK_c_5934_n N_CLK_c_6000_n \
 N_CLK_c_5956_n N_CLK_c_5959_n N_CLK_c_5961_n N_CLK_c_6054_n N_CLK_c_6056_n \
 N_CLK_c_6057_n N_CLK_c_5964_n N_CLK_c_5965_n N_CLK_c_6114_n N_CLK_c_6117_n \
 N_CLK_c_6356_p N_CLK_c_6363_p N_CLK_c_6119_n N_CLK_c_6120_n N_CLK_c_6121_n \
 N_CLK_c_6122_n N_CLK_c_6179_p N_CLK_c_6142_n N_CLK_c_6145_n N_CLK_c_6147_n \
 N_CLK_c_6163_p N_CLK_c_6261_p N_CLK_c_6197_p N_CLK_c_6150_n N_CLK_c_6151_n \
 N_CLK_c_5780_n N_CLK_c_5810_n N_CLK_c_5904_n N_CLK_c_5812_n N_CLK_c_5936_n \
 N_CLK_c_5966_n N_CLK_c_6065_n N_CLK_c_5968_n N_CLK_c_6124_n N_CLK_c_6152_n \
 N_CLK_c_6241_p N_CLK_c_6154_n )  PM_TMRDFFSNQX1\%CLK
x_PM_TMRDFFSNQX1\%noxref_18 ( N_noxref_18_c_6392_n N_noxref_18_c_6449_n \
 N_noxref_18_c_6393_n N_noxref_18_c_6402_n N_noxref_18_c_6458_n \
 N_noxref_18_c_6377_n N_noxref_18_c_6405_n N_noxref_18_c_6409_n \
 N_noxref_18_c_6411_n N_noxref_18_c_6415_n N_noxref_18_c_6379_n \
 N_noxref_18_c_6558_p N_noxref_18_c_6539_n N_noxref_18_c_6380_n \
 N_noxref_18_c_6542_n N_noxref_18_c_6583_p N_noxref_18_c_6422_n \
 N_noxref_18_c_6456_n N_noxref_18_M31_noxref_g N_noxref_18_M40_noxref_g \
 N_noxref_18_M114_noxref_g N_noxref_18_M115_noxref_g N_noxref_18_M132_noxref_g \
 N_noxref_18_M133_noxref_g N_noxref_18_c_6466_n N_noxref_18_c_6469_n \
 N_noxref_18_c_6471_n N_noxref_18_c_6503_n N_noxref_18_c_6505_n \
 N_noxref_18_c_6506_n N_noxref_18_c_6474_n N_noxref_18_c_6475_n \
 N_noxref_18_c_6381_n N_noxref_18_c_6383_n N_noxref_18_c_6384_n \
 N_noxref_18_c_6385_n N_noxref_18_c_6386_n N_noxref_18_c_6387_n \
 N_noxref_18_c_6388_n N_noxref_18_c_6390_n N_noxref_18_c_6476_n \
 N_noxref_18_c_6512_n N_noxref_18_c_6478_n N_noxref_18_c_6432_n \
 N_noxref_18_M34_noxref_d N_noxref_18_M116_noxref_d N_noxref_18_M118_noxref_d \
 N_noxref_18_M120_noxref_d )  PM_TMRDFFSNQX1\%noxref_18
x_PM_TMRDFFSNQX1\%noxref_19 ( N_noxref_19_c_6684_n N_noxref_19_c_6690_n \
 N_noxref_19_c_6694_n N_noxref_19_c_6698_n N_noxref_19_c_6700_n \
 N_noxref_19_c_6668_n N_noxref_19_c_6735_p N_noxref_19_c_6669_n \
 N_noxref_19_c_6670_n N_noxref_19_c_6799_p N_noxref_19_M42_noxref_g \
 N_noxref_19_M136_noxref_g N_noxref_19_M137_noxref_g N_noxref_19_c_6671_n \
 N_noxref_19_c_6673_n N_noxref_19_c_6674_n N_noxref_19_c_6675_n \
 N_noxref_19_c_6676_n N_noxref_19_c_6677_n N_noxref_19_c_6678_n \
 N_noxref_19_c_6680_n N_noxref_19_c_6743_p N_noxref_19_c_6713_n \
 N_noxref_19_M41_noxref_d N_noxref_19_M132_noxref_d N_noxref_19_M134_noxref_d ) \
 PM_TMRDFFSNQX1\%noxref_19
x_PM_TMRDFFSNQX1\%SN ( N_SN_c_6833_n N_SN_c_6843_n N_SN_c_6844_n N_SN_c_6854_n \
 N_SN_c_6855_n N_SN_c_6865_n N_SN_c_6866_n N_SN_c_6876_n N_SN_c_6877_n \
 N_SN_c_6887_n SN SN SN SN SN SN SN SN SN SN N_SN_c_6888_n N_SN_c_6889_n \
 N_SN_c_6890_n N_SN_c_6891_n N_SN_c_6892_n N_SN_c_6893_n N_SN_M6_noxref_g \
 N_SN_M13_noxref_g N_SN_M21_noxref_g N_SN_M28_noxref_g N_SN_M36_noxref_g \
 N_SN_M43_noxref_g N_SN_M64_noxref_g N_SN_M65_noxref_g N_SN_M78_noxref_g \
 N_SN_M79_noxref_g N_SN_M94_noxref_g N_SN_M95_noxref_g N_SN_M108_noxref_g \
 N_SN_M109_noxref_g N_SN_M124_noxref_g N_SN_M125_noxref_g N_SN_M138_noxref_g \
 N_SN_M139_noxref_g N_SN_c_6940_n N_SN_c_6943_n N_SN_c_7436_p N_SN_c_7444_p \
 N_SN_c_6945_n N_SN_c_6946_n N_SN_c_6947_n N_SN_c_6948_n N_SN_c_6965_n \
 N_SN_c_6986_n N_SN_c_6989_n N_SN_c_7476_p N_SN_c_7484_p N_SN_c_6991_n \
 N_SN_c_6992_n N_SN_c_6993_n N_SN_c_6994_n N_SN_c_7045_n N_SN_c_7070_n \
 N_SN_c_7073_n N_SN_c_7518_p N_SN_c_7526_p N_SN_c_7075_n N_SN_c_7076_n \
 N_SN_c_7077_n N_SN_c_7078_n N_SN_c_7095_n N_SN_c_7123_n N_SN_c_7126_n \
 N_SN_c_7558_p N_SN_c_7566_p N_SN_c_7128_n N_SN_c_7129_n N_SN_c_7130_n \
 N_SN_c_7131_n N_SN_c_7179_n N_SN_c_7244_n N_SN_c_7247_n N_SN_c_7600_p \
 N_SN_c_7608_p N_SN_c_7249_n N_SN_c_7250_n N_SN_c_7251_n N_SN_c_7252_n \
 N_SN_c_7269_n N_SN_c_7321_n N_SN_c_7324_n N_SN_c_7636_p N_SN_c_7643_p \
 N_SN_c_7326_n N_SN_c_7327_n N_SN_c_7328_n N_SN_c_7204_n N_SN_c_7378_p \
 N_SN_c_6950_n N_SN_c_6996_n N_SN_c_7080_n N_SN_c_7133_n N_SN_c_7254_n \
 N_SN_c_7331_n )  PM_TMRDFFSNQX1\%SN
x_PM_TMRDFFSNQX1\%noxref_21 ( N_noxref_21_c_7696_n N_noxref_21_c_7697_n \
 N_noxref_21_c_7698_n N_noxref_21_c_7699_n N_noxref_21_c_7656_n \
 N_noxref_21_c_7701_n N_noxref_21_c_7648_n N_noxref_21_c_7649_n \
 N_noxref_21_c_7660_n N_noxref_21_c_7664_n N_noxref_21_c_7666_n \
 N_noxref_21_c_7650_n N_noxref_21_c_7858_n N_noxref_21_c_7651_n \
 N_noxref_21_c_7652_n N_noxref_21_c_7774_n N_noxref_21_M34_noxref_g \
 N_noxref_21_M37_noxref_g N_noxref_21_M44_noxref_g N_noxref_21_M120_noxref_g \
 N_noxref_21_M121_noxref_g N_noxref_21_M126_noxref_g N_noxref_21_M127_noxref_g \
 N_noxref_21_M140_noxref_g N_noxref_21_M141_noxref_g N_noxref_21_c_7778_n \
 N_noxref_21_c_7779_n N_noxref_21_c_7780_n N_noxref_21_c_7830_n \
 N_noxref_21_c_7831_n N_noxref_21_c_7833_n N_noxref_21_c_7834_n \
 N_noxref_21_c_7729_n N_noxref_21_c_7730_n N_noxref_21_c_7731_n \
 N_noxref_21_c_7732_n N_noxref_21_c_7733_n N_noxref_21_c_7735_n \
 N_noxref_21_c_7736_n N_noxref_21_c_7875_n N_noxref_21_c_7876_n \
 N_noxref_21_c_7877_n N_noxref_21_c_7918_p N_noxref_21_c_7905_p \
 N_noxref_21_c_7920_p N_noxref_21_c_7906_p N_noxref_21_c_7781_n \
 N_noxref_21_c_7783_n N_noxref_21_c_7784_n N_noxref_21_c_7738_n \
 N_noxref_21_c_7739_n N_noxref_21_c_7741_n N_noxref_21_c_7706_n \
 N_noxref_21_c_7890_n N_noxref_21_c_7891_n N_noxref_21_M39_noxref_d \
 N_noxref_21_M128_noxref_d N_noxref_21_M130_noxref_d )  \
 PM_TMRDFFSNQX1\%noxref_21
x_PM_TMRDFFSNQX1\%noxref_22 ( N_noxref_22_c_7969_n N_noxref_22_c_7975_n \
 N_noxref_22_c_7980_n N_noxref_22_c_7984_n N_noxref_22_c_7986_n \
 N_noxref_22_c_7989_n N_noxref_22_c_8022_p N_noxref_22_c_7991_n \
 N_noxref_22_c_8034_p N_noxref_22_M142_noxref_d N_noxref_22_M144_noxref_d \
 N_noxref_22_M146_noxref_s N_noxref_22_M147_noxref_d N_noxref_22_M149_noxref_d \
 )  PM_TMRDFFSNQX1\%noxref_22
x_PM_TMRDFFSNQX1\%noxref_23 ( N_noxref_23_c_8089_n N_noxref_23_c_8092_n \
 N_noxref_23_c_8093_n N_noxref_23_c_8097_n N_noxref_23_c_8100_n \
 N_noxref_23_c_8105_n N_noxref_23_c_8213_n N_noxref_23_c_8060_n \
 N_noxref_23_c_8111_n N_noxref_23_c_8115_n N_noxref_23_c_8117_n \
 N_noxref_23_c_8121_n N_noxref_23_c_8062_n N_noxref_23_c_8177_n \
 N_noxref_23_c_8126_n N_noxref_23_c_8063_n N_noxref_23_c_8066_n \
 N_noxref_23_c_8288_n N_noxref_23_c_8312_n N_noxref_23_M41_noxref_g \
 N_noxref_23_M45_noxref_g N_noxref_23_M47_noxref_g N_noxref_23_M134_noxref_g \
 N_noxref_23_M135_noxref_g N_noxref_23_M142_noxref_g N_noxref_23_M143_noxref_g \
 N_noxref_23_M146_noxref_g N_noxref_23_M147_noxref_g N_noxref_23_c_8221_n \
 N_noxref_23_c_8224_n N_noxref_23_c_8226_n N_noxref_23_c_8263_n \
 N_noxref_23_c_8266_n N_noxref_23_c_8267_n N_noxref_23_c_8229_n \
 N_noxref_23_c_8230_n N_noxref_23_c_8068_n N_noxref_23_c_8070_n \
 N_noxref_23_c_8071_n N_noxref_23_c_8072_n N_noxref_23_c_8073_n \
 N_noxref_23_c_8074_n N_noxref_23_c_8197_n N_noxref_23_c_8146_n \
 N_noxref_23_c_8075_n N_noxref_23_c_8077_n N_noxref_23_c_8078_n \
 N_noxref_23_c_8080_n N_noxref_23_c_8363_p N_noxref_23_c_8081_n \
 N_noxref_23_c_8082_n N_noxref_23_c_8083_n N_noxref_23_c_8084_n \
 N_noxref_23_c_8086_n N_noxref_23_c_8231_n N_noxref_23_c_8273_n \
 N_noxref_23_c_8233_n N_noxref_23_c_8087_n N_noxref_23_c_8148_n \
 N_noxref_23_M44_noxref_d N_noxref_23_M136_noxref_d N_noxref_23_M138_noxref_d \
 N_noxref_23_M140_noxref_d )  PM_TMRDFFSNQX1\%noxref_23
x_PM_TMRDFFSNQX1\%noxref_24 ( N_noxref_24_c_8520_n N_noxref_24_c_8497_n \
 N_noxref_24_c_8424_n N_noxref_24_c_8558_n N_noxref_24_c_8426_n \
 N_noxref_24_c_8427_n N_noxref_24_c_8498_n N_noxref_24_c_8428_n \
 N_noxref_24_c_8451_n N_noxref_24_c_8455_n N_noxref_24_c_8457_n \
 N_noxref_24_c_8461_n N_noxref_24_c_8430_n N_noxref_24_c_8735_n \
 N_noxref_24_c_8465_n N_noxref_24_c_8431_n N_noxref_24_c_8433_n \
 N_noxref_24_c_8738_n N_noxref_24_c_8571_n N_noxref_24_M11_noxref_g \
 N_noxref_24_M48_noxref_g N_noxref_24_M49_noxref_g N_noxref_24_M74_noxref_g \
 N_noxref_24_M75_noxref_g N_noxref_24_M148_noxref_g N_noxref_24_M149_noxref_g \
 N_noxref_24_M150_noxref_g N_noxref_24_M151_noxref_g N_noxref_24_c_8506_n \
 N_noxref_24_c_8509_n N_noxref_24_c_8511_n N_noxref_24_c_8541_n \
 N_noxref_24_c_8543_n N_noxref_24_c_8544_n N_noxref_24_c_8514_n \
 N_noxref_24_c_8515_n N_noxref_24_c_8778_n N_noxref_24_c_8781_n \
 N_noxref_24_c_8805_p N_noxref_24_c_8640_n N_noxref_24_c_8833_p \
 N_noxref_24_c_8834_p N_noxref_24_c_8480_n N_noxref_24_c_8787_n \
 N_noxref_24_c_8788_n N_noxref_24_c_8789_n N_noxref_24_c_8434_n \
 N_noxref_24_c_8435_n N_noxref_24_c_8437_n N_noxref_24_c_8644_n \
 N_noxref_24_c_8438_n N_noxref_24_c_8439_n N_noxref_24_c_8440_n \
 N_noxref_24_c_8646_n N_noxref_24_c_8481_n N_noxref_24_c_8441_n \
 N_noxref_24_c_8443_n N_noxref_24_c_8516_n N_noxref_24_c_8550_n \
 N_noxref_24_c_8518_n N_noxref_24_c_8444_n N_noxref_24_M14_noxref_d \
 N_noxref_24_M76_noxref_d N_noxref_24_M78_noxref_d N_noxref_24_M80_noxref_d )  \
 PM_TMRDFFSNQX1\%noxref_24
x_PM_TMRDFFSNQX1\%noxref_25 ( N_noxref_25_c_8898_n N_noxref_25_c_8902_n \
 N_noxref_25_c_8916_n N_noxref_25_c_8904_n N_noxref_25_c_8905_n \
 N_noxref_25_c_8906_n N_noxref_25_c_8920_n N_noxref_25_c_8908_n \
 N_noxref_25_c_8921_n N_noxref_25_M146_noxref_d N_noxref_25_M148_noxref_d \
 N_noxref_25_M150_noxref_s N_noxref_25_M151_noxref_d N_noxref_25_M153_noxref_d \
 )  PM_TMRDFFSNQX1\%noxref_25
x_PM_TMRDFFSNQX1\%noxref_26 ( N_noxref_26_c_8988_n N_noxref_26_c_8995_n \
 N_noxref_26_c_8996_n N_noxref_26_c_9003_n N_noxref_26_c_9004_n \
 N_noxref_26_c_9007_n N_noxref_26_c_9089_n N_noxref_26_c_9045_n \
 N_noxref_26_c_9046_n N_noxref_26_c_9008_n N_noxref_26_c_9096_n \
 N_noxref_26_c_9010_n N_noxref_26_c_9011_n N_noxref_26_c_9105_n \
 N_noxref_26_M51_noxref_g N_noxref_26_M154_noxref_g N_noxref_26_M155_noxref_g \
 N_noxref_26_c_9016_n N_noxref_26_c_9216_p N_noxref_26_c_9217_p \
 N_noxref_26_c_9018_n N_noxref_26_c_9060_n N_noxref_26_c_9061_n \
 N_noxref_26_c_9019_n N_noxref_26_c_9208_p N_noxref_26_c_9020_n \
 N_noxref_26_c_9022_n N_noxref_26_c_9023_n N_noxref_26_M46_noxref_d \
 N_noxref_26_M48_noxref_d N_noxref_26_M50_noxref_d N_noxref_26_M150_noxref_d \
 N_noxref_26_M152_noxref_d )  PM_TMRDFFSNQX1\%noxref_26
x_PM_TMRDFFSNQX1\%noxref_27 ( N_noxref_27_c_9246_n N_noxref_27_c_9228_n \
 N_noxref_27_c_9232_n N_noxref_27_c_9235_n N_noxref_27_c_9236_n \
 N_noxref_27_c_9238_n N_noxref_27_M0_noxref_s )  PM_TMRDFFSNQX1\%noxref_27
x_PM_TMRDFFSNQX1\%noxref_28 ( N_noxref_28_c_9293_n N_noxref_28_c_9278_n \
 N_noxref_28_c_9282_n N_noxref_28_c_9285_n N_noxref_28_c_9304_n \
 N_noxref_28_M2_noxref_s )  PM_TMRDFFSNQX1\%noxref_28
x_PM_TMRDFFSNQX1\%noxref_29 ( N_noxref_29_c_9329_n N_noxref_29_c_9331_n \
 N_noxref_29_c_9334_n N_noxref_29_c_9336_n N_noxref_29_c_9347_n \
 N_noxref_29_M3_noxref_d N_noxref_29_M4_noxref_s )  PM_TMRDFFSNQX1\%noxref_29
x_PM_TMRDFFSNQX1\%noxref_30 ( N_noxref_30_c_9396_n N_noxref_30_c_9381_n \
 N_noxref_30_c_9385_n N_noxref_30_c_9388_n N_noxref_30_c_9412_n \
 N_noxref_30_M5_noxref_s )  PM_TMRDFFSNQX1\%noxref_30
x_PM_TMRDFFSNQX1\%noxref_31 ( N_noxref_31_c_9434_n N_noxref_31_c_9436_n \
 N_noxref_31_c_9439_n N_noxref_31_c_9441_n N_noxref_31_c_9449_n \
 N_noxref_31_M6_noxref_d N_noxref_31_M7_noxref_s )  PM_TMRDFFSNQX1\%noxref_31
x_PM_TMRDFFSNQX1\%noxref_32 ( N_noxref_32_c_9504_n N_noxref_32_c_9486_n \
 N_noxref_32_c_9490_n N_noxref_32_c_9493_n N_noxref_32_c_9494_n \
 N_noxref_32_c_9496_n N_noxref_32_M8_noxref_s )  PM_TMRDFFSNQX1\%noxref_32
x_PM_TMRDFFSNQX1\%noxref_33 ( N_noxref_33_c_9555_n N_noxref_33_c_9537_n \
 N_noxref_33_c_9541_n N_noxref_33_c_9544_n N_noxref_33_c_9545_n \
 N_noxref_33_c_9547_n N_noxref_33_M10_noxref_s )  PM_TMRDFFSNQX1\%noxref_33
x_PM_TMRDFFSNQX1\%noxref_34 ( N_noxref_34_c_9603_n N_noxref_34_c_9588_n \
 N_noxref_34_c_9592_n N_noxref_34_c_9595_n N_noxref_34_c_9619_n \
 N_noxref_34_M12_noxref_s )  PM_TMRDFFSNQX1\%noxref_34
x_PM_TMRDFFSNQX1\%noxref_35 ( N_noxref_35_c_9640_n N_noxref_35_c_9642_n \
 N_noxref_35_c_9645_n N_noxref_35_c_9647_n N_noxref_35_c_9657_n \
 N_noxref_35_M13_noxref_d N_noxref_35_M14_noxref_s )  PM_TMRDFFSNQX1\%noxref_35
x_PM_TMRDFFSNQX1\%noxref_36 ( N_noxref_36_c_9710_n N_noxref_36_c_9692_n \
 N_noxref_36_c_9696_n N_noxref_36_c_9699_n N_noxref_36_c_9700_n \
 N_noxref_36_c_9702_n N_noxref_36_M15_noxref_s )  PM_TMRDFFSNQX1\%noxref_36
x_PM_TMRDFFSNQX1\%noxref_37 ( N_noxref_37_c_9758_n N_noxref_37_c_9743_n \
 N_noxref_37_c_9747_n N_noxref_37_c_9750_n N_noxref_37_c_9773_n \
 N_noxref_37_M17_noxref_s )  PM_TMRDFFSNQX1\%noxref_37
x_PM_TMRDFFSNQX1\%noxref_38 ( N_noxref_38_c_9792_n N_noxref_38_c_9794_n \
 N_noxref_38_c_9797_n N_noxref_38_c_9799_n N_noxref_38_c_9807_n \
 N_noxref_38_M18_noxref_d N_noxref_38_M19_noxref_s )  PM_TMRDFFSNQX1\%noxref_38
x_PM_TMRDFFSNQX1\%noxref_39 ( N_noxref_39_c_9859_n N_noxref_39_c_9844_n \
 N_noxref_39_c_9848_n N_noxref_39_c_9851_n N_noxref_39_c_9876_n \
 N_noxref_39_M20_noxref_s )  PM_TMRDFFSNQX1\%noxref_39
x_PM_TMRDFFSNQX1\%noxref_40 ( N_noxref_40_c_9896_n N_noxref_40_c_9898_n \
 N_noxref_40_c_9901_n N_noxref_40_c_9903_n N_noxref_40_c_9911_n \
 N_noxref_40_M21_noxref_d N_noxref_40_M22_noxref_s )  PM_TMRDFFSNQX1\%noxref_40
x_PM_TMRDFFSNQX1\%noxref_41 ( N_noxref_41_c_9966_n N_noxref_41_c_9948_n \
 N_noxref_41_c_9952_n N_noxref_41_c_9955_n N_noxref_41_c_9956_n \
 N_noxref_41_c_9958_n N_noxref_41_M23_noxref_s )  PM_TMRDFFSNQX1\%noxref_41
x_PM_TMRDFFSNQX1\%noxref_42 ( N_noxref_42_c_10017_n N_noxref_42_c_9999_n \
 N_noxref_42_c_10003_n N_noxref_42_c_10006_n N_noxref_42_c_10007_n \
 N_noxref_42_c_10009_n N_noxref_42_M25_noxref_s )  PM_TMRDFFSNQX1\%noxref_42
x_PM_TMRDFFSNQX1\%noxref_43 ( N_noxref_43_c_10065_n N_noxref_43_c_10050_n \
 N_noxref_43_c_10054_n N_noxref_43_c_10057_n N_noxref_43_c_10082_n \
 N_noxref_43_M27_noxref_s )  PM_TMRDFFSNQX1\%noxref_43
x_PM_TMRDFFSNQX1\%noxref_44 ( N_noxref_44_c_10102_n N_noxref_44_c_10104_n \
 N_noxref_44_c_10107_n N_noxref_44_c_10109_n N_noxref_44_c_10119_n \
 N_noxref_44_M28_noxref_d N_noxref_44_M29_noxref_s )  PM_TMRDFFSNQX1\%noxref_44
x_PM_TMRDFFSNQX1\%noxref_45 ( N_noxref_45_c_10172_n N_noxref_45_c_10154_n \
 N_noxref_45_c_10158_n N_noxref_45_c_10161_n N_noxref_45_c_10162_n \
 N_noxref_45_c_10164_n N_noxref_45_M30_noxref_s )  PM_TMRDFFSNQX1\%noxref_45
x_PM_TMRDFFSNQX1\%noxref_46 ( N_noxref_46_c_10220_n N_noxref_46_c_10205_n \
 N_noxref_46_c_10209_n N_noxref_46_c_10212_n N_noxref_46_c_10234_n \
 N_noxref_46_M32_noxref_s )  PM_TMRDFFSNQX1\%noxref_46
x_PM_TMRDFFSNQX1\%noxref_47 ( N_noxref_47_c_10254_n N_noxref_47_c_10256_n \
 N_noxref_47_c_10259_n N_noxref_47_c_10261_n N_noxref_47_c_10281_n \
 N_noxref_47_M33_noxref_d N_noxref_47_M34_noxref_s )  PM_TMRDFFSNQX1\%noxref_47
x_PM_TMRDFFSNQX1\%noxref_48 ( N_noxref_48_c_10321_n N_noxref_48_c_10306_n \
 N_noxref_48_c_10310_n N_noxref_48_c_10313_n N_noxref_48_c_10338_n \
 N_noxref_48_M35_noxref_s )  PM_TMRDFFSNQX1\%noxref_48
x_PM_TMRDFFSNQX1\%noxref_49 ( N_noxref_49_c_10358_n N_noxref_49_c_10360_n \
 N_noxref_49_c_10363_n N_noxref_49_c_10365_n N_noxref_49_c_10373_n \
 N_noxref_49_M36_noxref_d N_noxref_49_M37_noxref_s )  PM_TMRDFFSNQX1\%noxref_49
x_PM_TMRDFFSNQX1\%noxref_50 ( N_noxref_50_c_10428_n N_noxref_50_c_10410_n \
 N_noxref_50_c_10414_n N_noxref_50_c_10417_n N_noxref_50_c_10418_n \
 N_noxref_50_c_10420_n N_noxref_50_M38_noxref_s )  PM_TMRDFFSNQX1\%noxref_50
x_PM_TMRDFFSNQX1\%noxref_51 ( N_noxref_51_c_10479_n N_noxref_51_c_10461_n \
 N_noxref_51_c_10465_n N_noxref_51_c_10468_n N_noxref_51_c_10469_n \
 N_noxref_51_c_10471_n N_noxref_51_M40_noxref_s )  PM_TMRDFFSNQX1\%noxref_51
x_PM_TMRDFFSNQX1\%noxref_52 ( N_noxref_52_c_10529_n N_noxref_52_c_10512_n \
 N_noxref_52_c_10516_n N_noxref_52_c_10519_n N_noxref_52_c_10527_n \
 N_noxref_52_M42_noxref_s )  PM_TMRDFFSNQX1\%noxref_52
x_PM_TMRDFFSNQX1\%noxref_53 ( N_noxref_53_c_10563_n N_noxref_53_c_10565_n \
 N_noxref_53_c_10568_n N_noxref_53_c_10570_n N_noxref_53_c_10595_n \
 N_noxref_53_M43_noxref_d N_noxref_53_M44_noxref_s )  PM_TMRDFFSNQX1\%noxref_53
x_PM_TMRDFFSNQX1\%noxref_54 ( N_noxref_54_c_10633_n N_noxref_54_c_10615_n \
 N_noxref_54_c_10619_n N_noxref_54_c_10622_n N_noxref_54_c_10623_n \
 N_noxref_54_c_10625_n N_noxref_54_M45_noxref_s )  PM_TMRDFFSNQX1\%noxref_54
x_PM_TMRDFFSNQX1\%noxref_55 ( N_noxref_55_c_10689_n N_noxref_55_c_10672_n \
 N_noxref_55_c_10675_n N_noxref_55_c_10678_n N_noxref_55_c_10679_n \
 N_noxref_55_c_10681_n N_noxref_55_M47_noxref_s )  PM_TMRDFFSNQX1\%noxref_55
x_PM_TMRDFFSNQX1\%noxref_56 ( N_noxref_56_c_10757_n N_noxref_56_c_10727_n \
 N_noxref_56_c_10730_n N_noxref_56_c_10733_n N_noxref_56_c_10734_n \
 N_noxref_56_c_10736_n N_noxref_56_M49_noxref_s )  PM_TMRDFFSNQX1\%noxref_56
x_PM_TMRDFFSNQX1\%Q ( Q Q Q Q Q Q Q N_Q_c_10784_n N_Q_c_10808_n N_Q_c_10794_n \
 N_Q_c_10797_n N_Q_M51_noxref_d N_Q_M154_noxref_d )  PM_TMRDFFSNQX1\%Q
cc_1 ( N_GND_c_1_p N_VDD_c_1012_n ) capacitor c=0.00989031f //x=0.74 //y=0 \
 //x2=0.74 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_1013_n ) capacitor c=0.00579636f //x=3.33 //y=0 \
 //x2=3.33 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_1014_n ) capacitor c=0.0057235f //x=8.14 //y=0 \
 //x2=8.14 //y2=7.4
cc_4 ( N_GND_c_4_p N_VDD_c_1015_n ) capacitor c=0.0057235f //x=12.95 //y=0 \
 //x2=12.95 //y2=7.4
cc_5 ( N_GND_c_5_p N_VDD_c_1016_n ) capacitor c=0.00474727f //x=16.28 //y=0 \
 //x2=16.28 //y2=7.4
cc_6 ( N_GND_c_6_p N_VDD_c_1017_n ) capacitor c=0.00474727f //x=19.61 //y=0 \
 //x2=19.61 //y2=7.4
cc_7 ( N_GND_c_7_p N_VDD_c_1018_n ) capacitor c=0.00891408f //x=24.42 //y=0 \
 //x2=24.42 //y2=7.4
cc_8 ( N_GND_c_8_p N_VDD_c_1019_n ) capacitor c=0.00576465f //x=27.75 //y=0 \
 //x2=27.75 //y2=7.4
cc_9 ( N_GND_c_9_p N_VDD_c_1020_n ) capacitor c=0.0057235f //x=32.56 //y=0 \
 //x2=32.56 //y2=7.4
cc_10 ( N_GND_c_10_p N_VDD_c_1021_n ) capacitor c=0.0057235f //x=37.37 //y=0 \
 //x2=37.37 //y2=7.4
cc_11 ( N_GND_c_11_p N_VDD_c_1022_n ) capacitor c=0.00474727f //x=40.7 //y=0 \
 //x2=40.7 //y2=7.4
cc_12 ( N_GND_c_12_p N_VDD_c_1023_n ) capacitor c=0.0057235f //x=44.03 //y=0 \
 //x2=44.03 //y2=7.4
cc_13 ( N_GND_c_13_p N_VDD_c_1024_n ) capacitor c=0.00989031f //x=48.84 //y=0 \
 //x2=48.84 //y2=7.4
cc_14 ( N_GND_c_14_p N_VDD_c_1025_n ) capacitor c=0.00576465f //x=52.17 //y=0 \
 //x2=52.17 //y2=7.4
cc_15 ( N_GND_c_15_p N_VDD_c_1026_n ) capacitor c=0.0057235f //x=56.98 //y=0 \
 //x2=56.98 //y2=7.4
cc_16 ( N_GND_c_16_p N_VDD_c_1027_n ) capacitor c=0.0057235f //x=61.79 //y=0 \
 //x2=61.79 //y2=7.4
cc_17 ( N_GND_c_17_p N_VDD_c_1028_n ) capacitor c=0.00474727f //x=65.12 //y=0 \
 //x2=65.12 //y2=7.4
cc_18 ( N_GND_c_18_p N_VDD_c_1029_n ) capacitor c=0.00891408f //x=68.45 //y=0 \
 //x2=68.45 //y2=7.4
cc_19 ( N_GND_c_19_p N_VDD_c_1030_n ) capacitor c=0.00891408f //x=73.26 //y=0 \
 //x2=73.26 //y2=7.4
cc_20 ( N_GND_c_20_p N_VDD_c_1031_n ) capacitor c=0.00504702f //x=76.59 //y=0 \
 //x2=76.59 //y2=7.4
cc_21 ( N_GND_c_21_p N_VDD_c_1032_n ) capacitor c=0.00553669f //x=79.92 //y=0 \
 //x2=79.92 //y2=7.4
cc_22 ( N_GND_c_22_p N_VDD_c_1033_n ) capacitor c=0.0052832f //x=83.25 //y=0 \
 //x2=83.25 //y2=7.4
cc_23 ( N_GND_c_23_p N_VDD_c_1034_n ) capacitor c=0.00989031f //x=84.85 //y=0 \
 //x2=84.73 //y2=7.4
cc_24 ( N_GND_c_24_p N_noxref_3_c_2117_n ) capacitor c=0.0139834f //x=84.73 \
 //y=0 //x2=4.295 //y2=2.59
cc_25 ( N_GND_c_25_p N_noxref_3_c_2117_n ) capacitor c=0.00230866f //x=3.16 \
 //y=0 //x2=4.295 //y2=2.59
cc_26 ( N_GND_c_26_p N_noxref_3_c_2117_n ) capacitor c=0.00221947f //x=4.32 \
 //y=0 //x2=4.295 //y2=2.59
cc_27 ( N_GND_c_2_p N_noxref_3_c_2117_n ) capacitor c=0.0338055f //x=3.33 \
 //y=0 //x2=4.295 //y2=2.59
cc_28 ( N_GND_c_24_p N_noxref_3_c_2121_n ) capacitor c=0.00222479f //x=84.73 \
 //y=0 //x2=2.705 //y2=2.59
cc_29 ( N_GND_c_2_p N_noxref_3_c_2121_n ) capacitor c=0.00111411f //x=3.33 \
 //y=0 //x2=2.705 //y2=2.59
cc_30 ( N_GND_c_24_p N_noxref_3_c_2123_n ) capacitor c=0.0394349f //x=84.73 \
 //y=0 //x2=9.135 //y2=2.59
cc_31 ( N_GND_c_31_p N_noxref_3_c_2123_n ) capacitor c=0.00344363f //x=7.97 \
 //y=0 //x2=9.135 //y2=2.59
cc_32 ( N_GND_c_32_p N_noxref_3_c_2123_n ) capacitor c=0.00221947f //x=9.13 \
 //y=0 //x2=9.135 //y2=2.59
cc_33 ( N_GND_c_3_p N_noxref_3_c_2123_n ) capacitor c=0.035311f //x=8.14 //y=0 \
 //x2=9.135 //y2=2.59
cc_34 ( N_GND_c_24_p N_noxref_3_c_2127_n ) capacitor c=0.0038075f //x=84.73 \
 //y=0 //x2=4.705 //y2=2.59
cc_35 ( N_GND_c_2_p N_noxref_3_c_2127_n ) capacitor c=7.88768e-19 //x=3.33 \
 //y=0 //x2=4.705 //y2=2.59
cc_36 ( N_GND_c_2_p N_noxref_3_c_2129_n ) capacitor c=0.0430571f //x=3.33 \
 //y=0 //x2=2.505 //y2=1.655
cc_37 ( N_GND_c_1_p N_noxref_3_c_2130_n ) capacitor c=0.00101801f //x=0.74 \
 //y=0 //x2=2.59 //y2=2.59
cc_38 ( N_GND_c_2_p N_noxref_3_c_2130_n ) capacitor c=5.56859e-19 //x=3.33 \
 //y=0 //x2=2.59 //y2=2.59
cc_39 ( N_GND_c_2_p N_noxref_3_c_2132_n ) capacitor c=0.0150282f //x=3.33 \
 //y=0 //x2=4.44 //y2=2.08
cc_40 ( N_GND_c_3_p N_noxref_3_c_2133_n ) capacitor c=0.0147449f //x=8.14 \
 //y=0 //x2=9.25 //y2=2.08
cc_41 ( N_GND_c_26_p N_noxref_3_c_2134_n ) capacitor c=0.00132755f //x=4.32 \
 //y=0 //x2=4.14 //y2=0.875
cc_42 ( N_GND_M2_noxref_d N_noxref_3_c_2134_n ) capacitor c=0.00211996f \
 //x=4.215 //y=0.875 //x2=4.14 //y2=0.875
cc_43 ( N_GND_M2_noxref_d N_noxref_3_c_2136_n ) capacitor c=0.00255985f \
 //x=4.215 //y=0.875 //x2=4.14 //y2=1.22
cc_44 ( N_GND_c_2_p N_noxref_3_c_2137_n ) capacitor c=0.00195164f //x=3.33 \
 //y=0 //x2=4.14 //y2=1.53
cc_45 ( N_GND_c_2_p N_noxref_3_c_2138_n ) capacitor c=0.0126573f //x=3.33 \
 //y=0 //x2=4.14 //y2=1.915
cc_46 ( N_GND_M2_noxref_d N_noxref_3_c_2139_n ) capacitor c=0.0131341f \
 //x=4.215 //y=0.875 //x2=4.515 //y2=0.72
cc_47 ( N_GND_M2_noxref_d N_noxref_3_c_2140_n ) capacitor c=0.00193146f \
 //x=4.215 //y=0.875 //x2=4.515 //y2=1.375
cc_48 ( N_GND_c_31_p N_noxref_3_c_2141_n ) capacitor c=0.00129018f //x=7.97 \
 //y=0 //x2=4.67 //y2=0.875
cc_49 ( N_GND_M2_noxref_d N_noxref_3_c_2141_n ) capacitor c=0.00257848f \
 //x=4.215 //y=0.875 //x2=4.67 //y2=0.875
cc_50 ( N_GND_M2_noxref_d N_noxref_3_c_2143_n ) capacitor c=0.00255985f \
 //x=4.215 //y=0.875 //x2=4.67 //y2=1.22
cc_51 ( N_GND_c_32_p N_noxref_3_c_2144_n ) capacitor c=0.00132755f //x=9.13 \
 //y=0 //x2=8.95 //y2=0.875
cc_52 ( N_GND_M5_noxref_d N_noxref_3_c_2144_n ) capacitor c=0.00211996f \
 //x=9.025 //y=0.875 //x2=8.95 //y2=0.875
cc_53 ( N_GND_M5_noxref_d N_noxref_3_c_2146_n ) capacitor c=0.00255985f \
 //x=9.025 //y=0.875 //x2=8.95 //y2=1.22
cc_54 ( N_GND_c_3_p N_noxref_3_c_2147_n ) capacitor c=0.00204716f //x=8.14 \
 //y=0 //x2=8.95 //y2=1.53
cc_55 ( N_GND_c_3_p N_noxref_3_c_2148_n ) capacitor c=0.0118433f //x=8.14 \
 //y=0 //x2=8.95 //y2=1.915
cc_56 ( N_GND_M5_noxref_d N_noxref_3_c_2149_n ) capacitor c=0.0131341f \
 //x=9.025 //y=0.875 //x2=9.325 //y2=0.72
cc_57 ( N_GND_M5_noxref_d N_noxref_3_c_2150_n ) capacitor c=0.00193146f \
 //x=9.025 //y=0.875 //x2=9.325 //y2=1.375
cc_58 ( N_GND_c_58_p N_noxref_3_c_2151_n ) capacitor c=0.00129018f //x=12.78 \
 //y=0 //x2=9.48 //y2=0.875
cc_59 ( N_GND_M5_noxref_d N_noxref_3_c_2151_n ) capacitor c=0.00257848f \
 //x=9.025 //y=0.875 //x2=9.48 //y2=0.875
cc_60 ( N_GND_M5_noxref_d N_noxref_3_c_2153_n ) capacitor c=0.00255985f \
 //x=9.025 //y=0.875 //x2=9.48 //y2=1.22
cc_61 ( N_GND_c_1_p N_noxref_3_M1_noxref_d ) capacitor c=8.58106e-19 //x=0.74 \
 //y=0 //x2=1.96 //y2=0.905
cc_62 ( N_GND_c_2_p N_noxref_3_M1_noxref_d ) capacitor c=0.00616547f //x=3.33 \
 //y=0 //x2=1.96 //y2=0.905
cc_63 ( N_GND_M0_noxref_d N_noxref_3_M1_noxref_d ) capacitor c=0.00143464f \
 //x=0.99 //y=0.865 //x2=1.96 //y2=0.905
cc_64 ( N_GND_c_4_p N_noxref_4_c_2361_n ) capacitor c=0.0222748f //x=12.95 \
 //y=0 //x2=13.945 //y2=2.59
cc_65 ( N_GND_c_4_p N_noxref_4_c_2362_n ) capacitor c=0.00102529f //x=12.95 \
 //y=0 //x2=12.325 //y2=2.59
cc_66 ( N_GND_c_4_p N_noxref_4_c_2363_n ) capacitor c=0.0401238f //x=12.95 \
 //y=0 //x2=12.125 //y2=1.665
cc_67 ( N_GND_c_4_p N_noxref_4_c_2364_n ) capacitor c=5.56859e-19 //x=12.95 \
 //y=0 //x2=12.21 //y2=2.59
cc_68 ( N_GND_c_4_p N_noxref_4_c_2365_n ) capacitor c=0.0128176f //x=12.95 \
 //y=0 //x2=14.06 //y2=2.08
cc_69 ( N_GND_c_69_p N_noxref_4_c_2366_n ) capacitor c=0.00135046f //x=14.045 \
 //y=0 //x2=13.865 //y2=0.865
cc_70 ( N_GND_M8_noxref_d N_noxref_4_c_2366_n ) capacitor c=0.00220047f \
 //x=13.94 //y=0.865 //x2=13.865 //y2=0.865
cc_71 ( N_GND_M8_noxref_d N_noxref_4_c_2368_n ) capacitor c=0.00255985f \
 //x=13.94 //y=0.865 //x2=13.865 //y2=1.21
cc_72 ( N_GND_c_4_p N_noxref_4_c_2369_n ) capacitor c=0.00189421f //x=12.95 \
 //y=0 //x2=13.865 //y2=1.52
cc_73 ( N_GND_c_4_p N_noxref_4_c_2370_n ) capacitor c=0.00992619f //x=12.95 \
 //y=0 //x2=13.865 //y2=1.915
cc_74 ( N_GND_M8_noxref_d N_noxref_4_c_2371_n ) capacitor c=0.0131326f \
 //x=13.94 //y=0.865 //x2=14.24 //y2=0.71
cc_75 ( N_GND_M8_noxref_d N_noxref_4_c_2372_n ) capacitor c=0.00193127f \
 //x=13.94 //y=0.865 //x2=14.24 //y2=1.365
cc_76 ( N_GND_c_76_p N_noxref_4_c_2373_n ) capacitor c=0.00130622f //x=16.11 \
 //y=0 //x2=14.395 //y2=0.865
cc_77 ( N_GND_M8_noxref_d N_noxref_4_c_2373_n ) capacitor c=0.00257848f \
 //x=13.94 //y=0.865 //x2=14.395 //y2=0.865
cc_78 ( N_GND_M8_noxref_d N_noxref_4_c_2375_n ) capacitor c=0.00255985f \
 //x=13.94 //y=0.865 //x2=14.395 //y2=1.21
cc_79 ( N_GND_c_4_p N_noxref_4_M7_noxref_d ) capacitor c=0.00591582f //x=12.95 \
 //y=0 //x2=11.535 //y2=0.915
cc_80 ( N_GND_c_1_p N_noxref_5_c_2525_n ) capacitor c=0.00115206f //x=0.74 \
 //y=0 //x2=1.85 //y2=2.08
cc_81 ( N_GND_c_2_p N_noxref_5_c_2525_n ) capacitor c=0.00110672f //x=3.33 \
 //y=0 //x2=1.85 //y2=2.08
cc_82 ( N_GND_c_3_p N_noxref_5_c_2527_n ) capacitor c=0.0425027f //x=8.14 \
 //y=0 //x2=7.315 //y2=1.665
cc_83 ( N_GND_c_5_p N_noxref_5_c_2528_n ) capacitor c=0.0154414f //x=16.28 \
 //y=0 //x2=17.39 //y2=2.08
cc_84 ( N_GND_c_84_p N_noxref_5_c_2529_n ) capacitor c=0.00135046f //x=17.375 \
 //y=0 //x2=17.195 //y2=0.865
cc_85 ( N_GND_M10_noxref_d N_noxref_5_c_2529_n ) capacitor c=0.00220047f \
 //x=17.27 //y=0.865 //x2=17.195 //y2=0.865
cc_86 ( N_GND_M10_noxref_d N_noxref_5_c_2531_n ) capacitor c=0.00255985f \
 //x=17.27 //y=0.865 //x2=17.195 //y2=1.21
cc_87 ( N_GND_c_5_p N_noxref_5_c_2532_n ) capacitor c=0.0018059f //x=16.28 \
 //y=0 //x2=17.195 //y2=1.52
cc_88 ( N_GND_c_5_p N_noxref_5_c_2533_n ) capacitor c=0.0101006f //x=16.28 \
 //y=0 //x2=17.195 //y2=1.915
cc_89 ( N_GND_M10_noxref_d N_noxref_5_c_2534_n ) capacitor c=0.0131326f \
 //x=17.27 //y=0.865 //x2=17.57 //y2=0.71
cc_90 ( N_GND_M10_noxref_d N_noxref_5_c_2535_n ) capacitor c=0.00193127f \
 //x=17.27 //y=0.865 //x2=17.57 //y2=1.365
cc_91 ( N_GND_c_91_p N_noxref_5_c_2536_n ) capacitor c=0.00130622f //x=19.44 \
 //y=0 //x2=17.725 //y2=0.865
cc_92 ( N_GND_M10_noxref_d N_noxref_5_c_2536_n ) capacitor c=0.00257848f \
 //x=17.27 //y=0.865 //x2=17.725 //y2=0.865
cc_93 ( N_GND_M10_noxref_d N_noxref_5_c_2538_n ) capacitor c=0.00255985f \
 //x=17.27 //y=0.865 //x2=17.725 //y2=1.21
cc_94 ( N_GND_c_3_p N_noxref_5_M4_noxref_d ) capacitor c=0.00591582f //x=8.14 \
 //y=0 //x2=6.725 //y2=0.915
cc_95 ( N_GND_c_6_p N_noxref_6_c_2803_n ) capacitor c=0.0435299f //x=19.61 \
 //y=0 //x2=18.785 //y2=1.655
cc_96 ( N_GND_c_5_p N_noxref_6_c_2804_n ) capacitor c=9.64732e-19 //x=16.28 \
 //y=0 //x2=18.87 //y2=4.07
cc_97 ( N_GND_c_6_p N_noxref_6_c_2805_n ) capacitor c=0.0156304f //x=19.61 \
 //y=0 //x2=20.72 //y2=2.08
cc_98 ( N_GND_c_98_p N_noxref_6_c_2806_n ) capacitor c=0.00132755f //x=20.6 \
 //y=0 //x2=20.42 //y2=0.875
cc_99 ( N_GND_M12_noxref_d N_noxref_6_c_2806_n ) capacitor c=0.00211996f \
 //x=20.495 //y=0.875 //x2=20.42 //y2=0.875
cc_100 ( N_GND_M12_noxref_d N_noxref_6_c_2808_n ) capacitor c=0.00255985f \
 //x=20.495 //y=0.875 //x2=20.42 //y2=1.22
cc_101 ( N_GND_c_6_p N_noxref_6_c_2809_n ) capacitor c=0.00195164f //x=19.61 \
 //y=0 //x2=20.42 //y2=1.53
cc_102 ( N_GND_c_6_p N_noxref_6_c_2810_n ) capacitor c=0.0110952f //x=19.61 \
 //y=0 //x2=20.42 //y2=1.915
cc_103 ( N_GND_M12_noxref_d N_noxref_6_c_2811_n ) capacitor c=0.0131341f \
 //x=20.495 //y=0.875 //x2=20.795 //y2=0.72
cc_104 ( N_GND_M12_noxref_d N_noxref_6_c_2812_n ) capacitor c=0.00193146f \
 //x=20.495 //y=0.875 //x2=20.795 //y2=1.375
cc_105 ( N_GND_c_105_p N_noxref_6_c_2813_n ) capacitor c=0.00129018f //x=24.25 \
 //y=0 //x2=20.95 //y2=0.875
cc_106 ( N_GND_M12_noxref_d N_noxref_6_c_2813_n ) capacitor c=0.00257848f \
 //x=20.495 //y=0.875 //x2=20.95 //y2=0.875
cc_107 ( N_GND_M12_noxref_d N_noxref_6_c_2815_n ) capacitor c=0.00255985f \
 //x=20.495 //y=0.875 //x2=20.95 //y2=1.22
cc_108 ( N_GND_c_5_p N_noxref_6_M11_noxref_d ) capacitor c=8.58106e-19 \
 //x=16.28 //y=0 //x2=18.24 //y2=0.905
cc_109 ( N_GND_c_6_p N_noxref_6_M11_noxref_d ) capacitor c=0.00616547f \
 //x=19.61 //y=0 //x2=18.24 //y2=0.905
cc_110 ( N_GND_M10_noxref_d N_noxref_6_M11_noxref_d ) capacitor c=0.00143464f \
 //x=17.27 //y=0.865 //x2=18.24 //y2=0.905
cc_111 ( N_GND_c_3_p N_noxref_7_c_2955_n ) capacitor c=7.88616e-19 //x=8.14 \
 //y=0 //x2=6.66 //y2=2.08
cc_112 ( N_GND_c_4_p N_noxref_7_c_2956_n ) capacitor c=0.00101012f //x=12.95 \
 //y=0 //x2=11.47 //y2=2.08
cc_113 ( N_GND_c_5_p N_noxref_7_c_2957_n ) capacitor c=0.0432305f //x=16.28 \
 //y=0 //x2=15.455 //y2=1.655
cc_114 ( N_GND_c_4_p N_noxref_7_c_2958_n ) capacitor c=9.64732e-19 //x=12.95 \
 //y=0 //x2=15.54 //y2=3.7
cc_115 ( N_GND_c_7_p N_noxref_7_c_2959_n ) capacitor c=8.62679e-19 //x=24.42 \
 //y=0 //x2=22.94 //y2=2.08
cc_116 ( N_GND_c_4_p N_noxref_7_M9_noxref_d ) capacitor c=8.58106e-19 \
 //x=12.95 //y=0 //x2=14.91 //y2=0.905
cc_117 ( N_GND_c_5_p N_noxref_7_M9_noxref_d ) capacitor c=0.00616547f \
 //x=16.28 //y=0 //x2=14.91 //y2=0.905
cc_118 ( N_GND_M8_noxref_d N_noxref_7_M9_noxref_d ) capacitor c=0.00143464f \
 //x=13.94 //y=0.865 //x2=14.91 //y2=0.905
cc_119 ( N_GND_c_8_p N_noxref_8_c_3277_n ) capacitor c=0.0215583f //x=27.75 \
 //y=0 //x2=28.715 //y2=2.59
cc_120 ( N_GND_c_8_p N_noxref_8_c_3278_n ) capacitor c=0.00111411f //x=27.75 \
 //y=0 //x2=27.125 //y2=2.59
cc_121 ( N_GND_c_9_p N_noxref_8_c_3279_n ) capacitor c=0.0230638f //x=32.56 \
 //y=0 //x2=33.555 //y2=2.59
cc_122 ( N_GND_c_8_p N_noxref_8_c_3280_n ) capacitor c=7.88768e-19 //x=27.75 \
 //y=0 //x2=29.125 //y2=2.59
cc_123 ( N_GND_c_8_p N_noxref_8_c_3281_n ) capacitor c=0.0404448f //x=27.75 \
 //y=0 //x2=26.925 //y2=1.655
cc_124 ( N_GND_c_7_p N_noxref_8_c_3282_n ) capacitor c=9.64732e-19 //x=24.42 \
 //y=0 //x2=27.01 //y2=2.59
cc_125 ( N_GND_c_8_p N_noxref_8_c_3282_n ) capacitor c=5.56859e-19 //x=27.75 \
 //y=0 //x2=27.01 //y2=2.59
cc_126 ( N_GND_c_8_p N_noxref_8_c_3284_n ) capacitor c=0.0127831f //x=27.75 \
 //y=0 //x2=28.86 //y2=2.08
cc_127 ( N_GND_c_9_p N_noxref_8_c_3285_n ) capacitor c=0.012616f //x=32.56 \
 //y=0 //x2=33.67 //y2=2.08
cc_128 ( N_GND_c_128_p N_noxref_8_c_3286_n ) capacitor c=0.00132755f //x=28.74 \
 //y=0 //x2=28.56 //y2=0.875
cc_129 ( N_GND_M17_noxref_d N_noxref_8_c_3286_n ) capacitor c=0.00211996f \
 //x=28.635 //y=0.875 //x2=28.56 //y2=0.875
cc_130 ( N_GND_M17_noxref_d N_noxref_8_c_3288_n ) capacitor c=0.00255985f \
 //x=28.635 //y=0.875 //x2=28.56 //y2=1.22
cc_131 ( N_GND_c_8_p N_noxref_8_c_3289_n ) capacitor c=0.00195164f //x=27.75 \
 //y=0 //x2=28.56 //y2=1.53
cc_132 ( N_GND_c_8_p N_noxref_8_c_3290_n ) capacitor c=0.0112696f //x=27.75 \
 //y=0 //x2=28.56 //y2=1.915
cc_133 ( N_GND_M17_noxref_d N_noxref_8_c_3291_n ) capacitor c=0.0131341f \
 //x=28.635 //y=0.875 //x2=28.935 //y2=0.72
cc_134 ( N_GND_M17_noxref_d N_noxref_8_c_3292_n ) capacitor c=0.00193146f \
 //x=28.635 //y=0.875 //x2=28.935 //y2=1.375
cc_135 ( N_GND_c_135_p N_noxref_8_c_3293_n ) capacitor c=0.00129018f //x=32.39 \
 //y=0 //x2=29.09 //y2=0.875
cc_136 ( N_GND_M17_noxref_d N_noxref_8_c_3293_n ) capacitor c=0.00257848f \
 //x=28.635 //y=0.875 //x2=29.09 //y2=0.875
cc_137 ( N_GND_M17_noxref_d N_noxref_8_c_3295_n ) capacitor c=0.00255985f \
 //x=28.635 //y=0.875 //x2=29.09 //y2=1.22
cc_138 ( N_GND_c_138_p N_noxref_8_c_3296_n ) capacitor c=0.00132755f //x=33.55 \
 //y=0 //x2=33.37 //y2=0.875
cc_139 ( N_GND_M20_noxref_d N_noxref_8_c_3296_n ) capacitor c=0.00211996f \
 //x=33.445 //y=0.875 //x2=33.37 //y2=0.875
cc_140 ( N_GND_M20_noxref_d N_noxref_8_c_3298_n ) capacitor c=0.00255985f \
 //x=33.445 //y=0.875 //x2=33.37 //y2=1.22
cc_141 ( N_GND_c_9_p N_noxref_8_c_3299_n ) capacitor c=0.00204716f //x=32.56 \
 //y=0 //x2=33.37 //y2=1.53
cc_142 ( N_GND_c_9_p N_noxref_8_c_3300_n ) capacitor c=0.0110952f //x=32.56 \
 //y=0 //x2=33.37 //y2=1.915
cc_143 ( N_GND_M20_noxref_d N_noxref_8_c_3301_n ) capacitor c=0.0131341f \
 //x=33.445 //y=0.875 //x2=33.745 //y2=0.72
cc_144 ( N_GND_M20_noxref_d N_noxref_8_c_3302_n ) capacitor c=0.00193146f \
 //x=33.445 //y=0.875 //x2=33.745 //y2=1.375
cc_145 ( N_GND_c_145_p N_noxref_8_c_3303_n ) capacitor c=0.00129018f //x=37.2 \
 //y=0 //x2=33.9 //y2=0.875
cc_146 ( N_GND_M20_noxref_d N_noxref_8_c_3303_n ) capacitor c=0.00257848f \
 //x=33.445 //y=0.875 //x2=33.9 //y2=0.875
cc_147 ( N_GND_M20_noxref_d N_noxref_8_c_3305_n ) capacitor c=0.00255985f \
 //x=33.445 //y=0.875 //x2=33.9 //y2=1.22
cc_148 ( N_GND_c_7_p N_noxref_8_M16_noxref_d ) capacitor c=8.58106e-19 \
 //x=24.42 //y=0 //x2=26.38 //y2=0.905
cc_149 ( N_GND_c_8_p N_noxref_8_M16_noxref_d ) capacitor c=0.00616547f \
 //x=27.75 //y=0 //x2=26.38 //y2=0.905
cc_150 ( N_GND_M15_noxref_d N_noxref_8_M16_noxref_d ) capacitor c=0.00143464f \
 //x=25.41 //y=0.865 //x2=26.38 //y2=0.905
cc_151 ( N_GND_c_10_p N_noxref_9_c_3509_n ) capacitor c=0.0222748f //x=37.37 \
 //y=0 //x2=38.365 //y2=2.59
cc_152 ( N_GND_c_10_p N_noxref_9_c_3510_n ) capacitor c=0.00102529f //x=37.37 \
 //y=0 //x2=36.745 //y2=2.59
cc_153 ( N_GND_c_10_p N_noxref_9_c_3511_n ) capacitor c=0.0401238f //x=37.37 \
 //y=0 //x2=36.545 //y2=1.665
cc_154 ( N_GND_c_10_p N_noxref_9_c_3512_n ) capacitor c=5.56859e-19 //x=37.37 \
 //y=0 //x2=36.63 //y2=2.59
cc_155 ( N_GND_c_10_p N_noxref_9_c_3513_n ) capacitor c=0.0128176f //x=37.37 \
 //y=0 //x2=38.48 //y2=2.08
cc_156 ( N_GND_c_156_p N_noxref_9_c_3514_n ) capacitor c=0.00135046f \
 //x=38.465 //y=0 //x2=38.285 //y2=0.865
cc_157 ( N_GND_M23_noxref_d N_noxref_9_c_3514_n ) capacitor c=0.00220047f \
 //x=38.36 //y=0.865 //x2=38.285 //y2=0.865
cc_158 ( N_GND_M23_noxref_d N_noxref_9_c_3516_n ) capacitor c=0.00255985f \
 //x=38.36 //y=0.865 //x2=38.285 //y2=1.21
cc_159 ( N_GND_c_10_p N_noxref_9_c_3517_n ) capacitor c=0.00189421f //x=37.37 \
 //y=0 //x2=38.285 //y2=1.52
cc_160 ( N_GND_c_10_p N_noxref_9_c_3518_n ) capacitor c=0.00992619f //x=37.37 \
 //y=0 //x2=38.285 //y2=1.915
cc_161 ( N_GND_M23_noxref_d N_noxref_9_c_3519_n ) capacitor c=0.0131326f \
 //x=38.36 //y=0.865 //x2=38.66 //y2=0.71
cc_162 ( N_GND_M23_noxref_d N_noxref_9_c_3520_n ) capacitor c=0.00193127f \
 //x=38.36 //y=0.865 //x2=38.66 //y2=1.365
cc_163 ( N_GND_c_163_p N_noxref_9_c_3521_n ) capacitor c=0.00130622f //x=40.53 \
 //y=0 //x2=38.815 //y2=0.865
cc_164 ( N_GND_M23_noxref_d N_noxref_9_c_3521_n ) capacitor c=0.00257848f \
 //x=38.36 //y=0.865 //x2=38.815 //y2=0.865
cc_165 ( N_GND_M23_noxref_d N_noxref_9_c_3523_n ) capacitor c=0.00255985f \
 //x=38.36 //y=0.865 //x2=38.815 //y2=1.21
cc_166 ( N_GND_c_10_p N_noxref_9_M22_noxref_d ) capacitor c=0.00591582f \
 //x=37.37 //y=0 //x2=35.955 //y2=0.915
cc_167 ( N_GND_c_7_p N_noxref_10_c_3675_n ) capacitor c=9.42296e-19 //x=24.42 \
 //y=0 //x2=26.27 //y2=2.08
cc_168 ( N_GND_c_8_p N_noxref_10_c_3675_n ) capacitor c=9.30131e-19 //x=27.75 \
 //y=0 //x2=26.27 //y2=2.08
cc_169 ( N_GND_c_9_p N_noxref_10_c_3677_n ) capacitor c=0.0401588f //x=32.56 \
 //y=0 //x2=31.735 //y2=1.665
cc_170 ( N_GND_c_11_p N_noxref_10_c_3678_n ) capacitor c=0.0151571f //x=40.7 \
 //y=0 //x2=41.81 //y2=2.08
cc_171 ( N_GND_c_171_p N_noxref_10_c_3679_n ) capacitor c=0.00135046f \
 //x=41.795 //y=0 //x2=41.615 //y2=0.865
cc_172 ( N_GND_M25_noxref_d N_noxref_10_c_3679_n ) capacitor c=0.00220047f \
 //x=41.69 //y=0.865 //x2=41.615 //y2=0.865
cc_173 ( N_GND_M25_noxref_d N_noxref_10_c_3681_n ) capacitor c=0.00255985f \
 //x=41.69 //y=0.865 //x2=41.615 //y2=1.21
cc_174 ( N_GND_c_11_p N_noxref_10_c_3682_n ) capacitor c=0.0018059f //x=40.7 \
 //y=0 //x2=41.615 //y2=1.52
cc_175 ( N_GND_c_11_p N_noxref_10_c_3683_n ) capacitor c=0.0101006f //x=40.7 \
 //y=0 //x2=41.615 //y2=1.915
cc_176 ( N_GND_M25_noxref_d N_noxref_10_c_3684_n ) capacitor c=0.0131326f \
 //x=41.69 //y=0.865 //x2=41.99 //y2=0.71
cc_177 ( N_GND_M25_noxref_d N_noxref_10_c_3685_n ) capacitor c=0.00193127f \
 //x=41.69 //y=0.865 //x2=41.99 //y2=1.365
cc_178 ( N_GND_c_178_p N_noxref_10_c_3686_n ) capacitor c=0.00130622f \
 //x=43.86 //y=0 //x2=42.145 //y2=0.865
cc_179 ( N_GND_M25_noxref_d N_noxref_10_c_3686_n ) capacitor c=0.00257848f \
 //x=41.69 //y=0.865 //x2=42.145 //y2=0.865
cc_180 ( N_GND_M25_noxref_d N_noxref_10_c_3688_n ) capacitor c=0.00255985f \
 //x=41.69 //y=0.865 //x2=42.145 //y2=1.21
cc_181 ( N_GND_c_9_p N_noxref_10_M19_noxref_d ) capacitor c=0.00591582f \
 //x=32.56 //y=0 //x2=31.145 //y2=0.915
cc_182 ( N_GND_c_12_p N_noxref_11_c_3956_n ) capacitor c=0.0222748f //x=44.03 \
 //y=0 //x2=45.025 //y2=2.59
cc_183 ( N_GND_c_12_p N_noxref_11_c_3957_n ) capacitor c=0.00102529f //x=44.03 \
 //y=0 //x2=43.405 //y2=2.59
cc_184 ( N_GND_c_12_p N_noxref_11_c_3958_n ) capacitor c=0.0403754f //x=44.03 \
 //y=0 //x2=43.205 //y2=1.655
cc_185 ( N_GND_c_11_p N_noxref_11_c_3959_n ) capacitor c=9.64732e-19 //x=40.7 \
 //y=0 //x2=43.29 //y2=2.59
cc_186 ( N_GND_c_12_p N_noxref_11_c_3959_n ) capacitor c=5.56859e-19 //x=44.03 \
 //y=0 //x2=43.29 //y2=2.59
cc_187 ( N_GND_c_12_p N_noxref_11_c_3961_n ) capacitor c=0.0127526f //x=44.03 \
 //y=0 //x2=45.14 //y2=2.08
cc_188 ( N_GND_c_188_p N_noxref_11_c_3962_n ) capacitor c=0.00132755f \
 //x=45.02 //y=0 //x2=44.84 //y2=0.875
cc_189 ( N_GND_M27_noxref_d N_noxref_11_c_3962_n ) capacitor c=0.00211996f \
 //x=44.915 //y=0.875 //x2=44.84 //y2=0.875
cc_190 ( N_GND_M27_noxref_d N_noxref_11_c_3964_n ) capacitor c=0.00255985f \
 //x=44.915 //y=0.875 //x2=44.84 //y2=1.22
cc_191 ( N_GND_c_12_p N_noxref_11_c_3965_n ) capacitor c=0.00195164f //x=44.03 \
 //y=0 //x2=44.84 //y2=1.53
cc_192 ( N_GND_c_12_p N_noxref_11_c_3966_n ) capacitor c=0.0110952f //x=44.03 \
 //y=0 //x2=44.84 //y2=1.915
cc_193 ( N_GND_M27_noxref_d N_noxref_11_c_3967_n ) capacitor c=0.0131341f \
 //x=44.915 //y=0.875 //x2=45.215 //y2=0.72
cc_194 ( N_GND_M27_noxref_d N_noxref_11_c_3968_n ) capacitor c=0.00193146f \
 //x=44.915 //y=0.875 //x2=45.215 //y2=1.375
cc_195 ( N_GND_c_195_p N_noxref_11_c_3969_n ) capacitor c=0.00129018f \
 //x=48.67 //y=0 //x2=45.37 //y2=0.875
cc_196 ( N_GND_M27_noxref_d N_noxref_11_c_3969_n ) capacitor c=0.00257848f \
 //x=44.915 //y=0.875 //x2=45.37 //y2=0.875
cc_197 ( N_GND_M27_noxref_d N_noxref_11_c_3971_n ) capacitor c=0.00255985f \
 //x=44.915 //y=0.875 //x2=45.37 //y2=1.22
cc_198 ( N_GND_c_11_p N_noxref_11_M26_noxref_d ) capacitor c=8.58106e-19 \
 //x=40.7 //y=0 //x2=42.66 //y2=0.905
cc_199 ( N_GND_c_12_p N_noxref_11_M26_noxref_d ) capacitor c=0.00616547f \
 //x=44.03 //y=0 //x2=42.66 //y2=0.905
cc_200 ( N_GND_M25_noxref_d N_noxref_11_M26_noxref_d ) capacitor c=0.00143464f \
 //x=41.69 //y=0.865 //x2=42.66 //y2=0.905
cc_201 ( N_GND_c_9_p N_noxref_12_c_4111_n ) capacitor c=6.12031e-19 //x=32.56 \
 //y=0 //x2=31.08 //y2=2.08
cc_202 ( N_GND_c_10_p N_noxref_12_c_4112_n ) capacitor c=0.00101012f //x=37.37 \
 //y=0 //x2=35.89 //y2=2.08
cc_203 ( N_GND_c_11_p N_noxref_12_c_4113_n ) capacitor c=0.042884f //x=40.7 \
 //y=0 //x2=39.875 //y2=1.655
cc_204 ( N_GND_c_10_p N_noxref_12_c_4114_n ) capacitor c=9.64732e-19 //x=37.37 \
 //y=0 //x2=39.96 //y2=3.7
cc_205 ( N_GND_c_13_p N_noxref_12_c_4115_n ) capacitor c=0.00102842f //x=48.84 \
 //y=0 //x2=47.36 //y2=2.08
cc_206 ( N_GND_c_10_p N_noxref_12_M24_noxref_d ) capacitor c=8.58106e-19 \
 //x=37.37 //y=0 //x2=39.33 //y2=0.905
cc_207 ( N_GND_c_11_p N_noxref_12_M24_noxref_d ) capacitor c=0.00616547f \
 //x=40.7 //y=0 //x2=39.33 //y2=0.905
cc_208 ( N_GND_M23_noxref_d N_noxref_12_M24_noxref_d ) capacitor c=0.00143464f \
 //x=38.36 //y=0.865 //x2=39.33 //y2=0.905
cc_209 ( N_GND_c_13_p N_noxref_13_c_4433_n ) capacitor c=0.0215583f //x=48.84 \
 //y=0 //x2=50.605 //y2=2.59
cc_210 ( N_GND_c_13_p N_noxref_13_c_4434_n ) capacitor c=0.00124977f //x=48.84 \
 //y=0 //x2=48.215 //y2=2.59
cc_211 ( N_GND_c_24_p N_noxref_13_c_4435_n ) capacitor c=0.0571584f //x=84.73 \
 //y=0 //x2=74.995 //y2=2.96
cc_212 ( N_GND_c_212_p N_noxref_13_c_4435_n ) capacitor c=0.00282695f \
 //x=73.09 //y=0 //x2=74.995 //y2=2.96
cc_213 ( N_GND_c_213_p N_noxref_13_c_4435_n ) capacitor c=0.0019279f \
 //x=74.355 //y=0 //x2=74.995 //y2=2.96
cc_214 ( N_GND_c_14_p N_noxref_13_c_4435_n ) capacitor c=0.00750857f //x=52.17 \
 //y=0 //x2=74.995 //y2=2.96
cc_215 ( N_GND_c_15_p N_noxref_13_c_4435_n ) capacitor c=0.00750857f //x=56.98 \
 //y=0 //x2=74.995 //y2=2.96
cc_216 ( N_GND_c_16_p N_noxref_13_c_4435_n ) capacitor c=0.00750857f //x=61.79 \
 //y=0 //x2=74.995 //y2=2.96
cc_217 ( N_GND_c_17_p N_noxref_13_c_4435_n ) capacitor c=0.00949826f //x=65.12 \
 //y=0 //x2=74.995 //y2=2.96
cc_218 ( N_GND_c_18_p N_noxref_13_c_4435_n ) capacitor c=0.00949826f //x=68.45 \
 //y=0 //x2=74.995 //y2=2.96
cc_219 ( N_GND_c_19_p N_noxref_13_c_4435_n ) capacitor c=0.0144849f //x=73.26 \
 //y=0 //x2=74.995 //y2=2.96
cc_220 ( N_GND_c_21_p N_noxref_13_c_4444_n ) capacitor c=0.00281233f //x=79.92 \
 //y=0 //x2=81.655 //y2=4.07
cc_221 ( N_GND_c_11_p N_noxref_13_c_4445_n ) capacitor c=9.42296e-19 //x=40.7 \
 //y=0 //x2=42.55 //y2=2.08
cc_222 ( N_GND_c_12_p N_noxref_13_c_4445_n ) capacitor c=9.24123e-19 //x=44.03 \
 //y=0 //x2=42.55 //y2=2.08
cc_223 ( N_GND_c_13_p N_noxref_13_c_4447_n ) capacitor c=0.040141f //x=48.84 \
 //y=0 //x2=48.015 //y2=1.665
cc_224 ( N_GND_c_13_p N_noxref_13_c_4448_n ) capacitor c=5.56859e-19 //x=48.84 \
 //y=0 //x2=48.1 //y2=2.59
cc_225 ( N_GND_c_19_p N_noxref_13_c_4449_n ) capacitor c=0.00123238f //x=73.26 \
 //y=0 //x2=75.11 //y2=2.08
cc_226 ( N_GND_c_20_p N_noxref_13_c_4449_n ) capacitor c=0.0125771f //x=76.59 \
 //y=0 //x2=75.11 //y2=2.08
cc_227 ( N_GND_c_21_p N_noxref_13_c_4451_n ) capacitor c=8.50308e-19 //x=79.92 \
 //y=0 //x2=81.77 //y2=2.08
cc_228 ( N_GND_c_22_p N_noxref_13_c_4451_n ) capacitor c=0.00128267f //x=83.25 \
 //y=0 //x2=81.77 //y2=2.08
cc_229 ( N_GND_c_20_p N_noxref_13_c_4453_n ) capacitor c=2.63786e-19 //x=76.59 \
 //y=0 //x2=75.11 //y2=2.08
cc_230 ( N_GND_c_13_p N_noxref_13_M29_noxref_d ) capacitor c=0.00591582f \
 //x=48.84 //y=0 //x2=47.425 //y2=0.915
cc_231 ( N_GND_c_24_p N_D_c_4900_n ) capacitor c=0.0727405f //x=84.73 //y=0 \
 //x2=25.415 //y2=2.96
cc_232 ( N_GND_c_25_p N_D_c_4900_n ) capacitor c=6.3489e-19 //x=3.16 //y=0 \
 //x2=25.415 //y2=2.96
cc_233 ( N_GND_c_2_p N_D_c_4900_n ) capacitor c=0.00750857f //x=3.33 //y=0 \
 //x2=25.415 //y2=2.96
cc_234 ( N_GND_c_3_p N_D_c_4900_n ) capacitor c=0.00750857f //x=8.14 //y=0 \
 //x2=25.415 //y2=2.96
cc_235 ( N_GND_c_4_p N_D_c_4900_n ) capacitor c=0.00750857f //x=12.95 //y=0 \
 //x2=25.415 //y2=2.96
cc_236 ( N_GND_c_5_p N_D_c_4900_n ) capacitor c=0.00949826f //x=16.28 //y=0 \
 //x2=25.415 //y2=2.96
cc_237 ( N_GND_c_6_p N_D_c_4900_n ) capacitor c=0.00949826f //x=19.61 //y=0 \
 //x2=25.415 //y2=2.96
cc_238 ( N_GND_c_7_p N_D_c_4900_n ) capacitor c=0.00949826f //x=24.42 //y=0 \
 //x2=25.415 //y2=2.96
cc_239 ( N_GND_c_24_p N_D_c_4908_n ) capacitor c=0.00207889f //x=84.73 //y=0 \
 //x2=1.225 //y2=2.96
cc_240 ( N_GND_c_8_p N_D_c_4909_n ) capacitor c=0.00750857f //x=27.75 //y=0 \
 //x2=49.835 //y2=2.96
cc_241 ( N_GND_c_9_p N_D_c_4909_n ) capacitor c=0.00750857f //x=32.56 //y=0 \
 //x2=49.835 //y2=2.96
cc_242 ( N_GND_c_10_p N_D_c_4909_n ) capacitor c=0.00750857f //x=37.37 //y=0 \
 //x2=49.835 //y2=2.96
cc_243 ( N_GND_c_11_p N_D_c_4909_n ) capacitor c=0.00949826f //x=40.7 //y=0 \
 //x2=49.835 //y2=2.96
cc_244 ( N_GND_c_12_p N_D_c_4909_n ) capacitor c=0.00750857f //x=44.03 //y=0 \
 //x2=49.835 //y2=2.96
cc_245 ( N_GND_c_13_p N_D_c_4909_n ) capacitor c=0.00750857f //x=48.84 //y=0 \
 //x2=49.835 //y2=2.96
cc_246 ( N_GND_c_1_p N_D_c_4915_n ) capacitor c=0.0177675f //x=0.74 //y=0 \
 //x2=1.11 //y2=2.08
cc_247 ( N_GND_c_7_p N_D_c_4916_n ) capacitor c=0.0154111f //x=24.42 //y=0 \
 //x2=25.53 //y2=2.08
cc_248 ( N_GND_c_13_p N_D_c_4917_n ) capacitor c=0.012911f //x=48.84 //y=0 \
 //x2=49.95 //y2=2.08
cc_249 ( N_GND_c_249_p N_D_c_4918_n ) capacitor c=0.00135046f //x=1.095 //y=0 \
 //x2=0.915 //y2=0.865
cc_250 ( N_GND_M0_noxref_d N_D_c_4918_n ) capacitor c=0.00220047f //x=0.99 \
 //y=0.865 //x2=0.915 //y2=0.865
cc_251 ( N_GND_M0_noxref_d N_D_c_4920_n ) capacitor c=0.00255985f //x=0.99 \
 //y=0.865 //x2=0.915 //y2=1.21
cc_252 ( N_GND_c_1_p N_D_c_4921_n ) capacitor c=0.00264481f //x=0.74 //y=0 \
 //x2=0.915 //y2=1.52
cc_253 ( N_GND_c_1_p N_D_c_4922_n ) capacitor c=0.0121947f //x=0.74 //y=0 \
 //x2=0.915 //y2=1.915
cc_254 ( N_GND_M0_noxref_d N_D_c_4923_n ) capacitor c=0.0131326f //x=0.99 \
 //y=0.865 //x2=1.29 //y2=0.71
cc_255 ( N_GND_M0_noxref_d N_D_c_4924_n ) capacitor c=0.00193127f //x=0.99 \
 //y=0.865 //x2=1.29 //y2=1.365
cc_256 ( N_GND_c_25_p N_D_c_4925_n ) capacitor c=0.00130622f //x=3.16 //y=0 \
 //x2=1.445 //y2=0.865
cc_257 ( N_GND_M0_noxref_d N_D_c_4925_n ) capacitor c=0.00257848f //x=0.99 \
 //y=0.865 //x2=1.445 //y2=0.865
cc_258 ( N_GND_M0_noxref_d N_D_c_4927_n ) capacitor c=0.00255985f //x=0.99 \
 //y=0.865 //x2=1.445 //y2=1.21
cc_259 ( N_GND_c_259_p N_D_c_4928_n ) capacitor c=0.00135046f //x=25.515 //y=0 \
 //x2=25.335 //y2=0.865
cc_260 ( N_GND_M15_noxref_d N_D_c_4928_n ) capacitor c=0.00220047f //x=25.41 \
 //y=0.865 //x2=25.335 //y2=0.865
cc_261 ( N_GND_M15_noxref_d N_D_c_4930_n ) capacitor c=0.00255985f //x=25.41 \
 //y=0.865 //x2=25.335 //y2=1.21
cc_262 ( N_GND_c_7_p N_D_c_4931_n ) capacitor c=0.00189421f //x=24.42 //y=0 \
 //x2=25.335 //y2=1.52
cc_263 ( N_GND_c_7_p N_D_c_4932_n ) capacitor c=0.00992619f //x=24.42 //y=0 \
 //x2=25.335 //y2=1.915
cc_264 ( N_GND_M15_noxref_d N_D_c_4933_n ) capacitor c=0.0131326f //x=25.41 \
 //y=0.865 //x2=25.71 //y2=0.71
cc_265 ( N_GND_M15_noxref_d N_D_c_4934_n ) capacitor c=0.00193127f //x=25.41 \
 //y=0.865 //x2=25.71 //y2=1.365
cc_266 ( N_GND_c_266_p N_D_c_4935_n ) capacitor c=0.00130622f //x=27.58 //y=0 \
 //x2=25.865 //y2=0.865
cc_267 ( N_GND_M15_noxref_d N_D_c_4935_n ) capacitor c=0.00257848f //x=25.41 \
 //y=0.865 //x2=25.865 //y2=0.865
cc_268 ( N_GND_M15_noxref_d N_D_c_4937_n ) capacitor c=0.00255985f //x=25.41 \
 //y=0.865 //x2=25.865 //y2=1.21
cc_269 ( N_GND_c_269_p N_D_c_4938_n ) capacitor c=0.00135046f //x=49.935 //y=0 \
 //x2=49.755 //y2=0.865
cc_270 ( N_GND_M30_noxref_d N_D_c_4938_n ) capacitor c=0.00220047f //x=49.83 \
 //y=0.865 //x2=49.755 //y2=0.865
cc_271 ( N_GND_M30_noxref_d N_D_c_4940_n ) capacitor c=0.00255985f //x=49.83 \
 //y=0.865 //x2=49.755 //y2=1.21
cc_272 ( N_GND_c_13_p N_D_c_4941_n ) capacitor c=0.00189421f //x=48.84 //y=0 \
 //x2=49.755 //y2=1.52
cc_273 ( N_GND_c_13_p N_D_c_4942_n ) capacitor c=0.00992619f //x=48.84 //y=0 \
 //x2=49.755 //y2=1.915
cc_274 ( N_GND_M30_noxref_d N_D_c_4943_n ) capacitor c=0.0131326f //x=49.83 \
 //y=0.865 //x2=50.13 //y2=0.71
cc_275 ( N_GND_M30_noxref_d N_D_c_4944_n ) capacitor c=0.00193127f //x=49.83 \
 //y=0.865 //x2=50.13 //y2=1.365
cc_276 ( N_GND_c_276_p N_D_c_4945_n ) capacitor c=0.00130622f //x=52 //y=0 \
 //x2=50.285 //y2=0.865
cc_277 ( N_GND_M30_noxref_d N_D_c_4945_n ) capacitor c=0.00257848f //x=49.83 \
 //y=0.865 //x2=50.285 //y2=0.865
cc_278 ( N_GND_M30_noxref_d N_D_c_4947_n ) capacitor c=0.00255985f //x=49.83 \
 //y=0.865 //x2=50.285 //y2=1.21
cc_279 ( N_GND_c_14_p N_noxref_15_c_5221_n ) capacitor c=0.0215583f //x=52.17 \
 //y=0 //x2=53.135 //y2=2.59
cc_280 ( N_GND_c_14_p N_noxref_15_c_5222_n ) capacitor c=0.00106523f //x=52.17 \
 //y=0 //x2=51.545 //y2=2.59
cc_281 ( N_GND_c_15_p N_noxref_15_c_5223_n ) capacitor c=0.0230638f //x=56.98 \
 //y=0 //x2=57.975 //y2=2.59
cc_282 ( N_GND_c_14_p N_noxref_15_c_5224_n ) capacitor c=7.88768e-19 //x=52.17 \
 //y=0 //x2=53.545 //y2=2.59
cc_283 ( N_GND_c_14_p N_noxref_15_c_5225_n ) capacitor c=0.0404062f //x=52.17 \
 //y=0 //x2=51.345 //y2=1.655
cc_284 ( N_GND_c_13_p N_noxref_15_c_5226_n ) capacitor c=9.64732e-19 //x=48.84 \
 //y=0 //x2=51.43 //y2=2.59
cc_285 ( N_GND_c_14_p N_noxref_15_c_5226_n ) capacitor c=5.56859e-19 //x=52.17 \
 //y=0 //x2=51.43 //y2=2.59
cc_286 ( N_GND_c_14_p N_noxref_15_c_5228_n ) capacitor c=0.012765f //x=52.17 \
 //y=0 //x2=53.28 //y2=2.08
cc_287 ( N_GND_c_15_p N_noxref_15_c_5229_n ) capacitor c=0.012616f //x=56.98 \
 //y=0 //x2=58.09 //y2=2.08
cc_288 ( N_GND_c_288_p N_noxref_15_c_5230_n ) capacitor c=0.00132755f \
 //x=53.16 //y=0 //x2=52.98 //y2=0.875
cc_289 ( N_GND_M32_noxref_d N_noxref_15_c_5230_n ) capacitor c=0.00211996f \
 //x=53.055 //y=0.875 //x2=52.98 //y2=0.875
cc_290 ( N_GND_M32_noxref_d N_noxref_15_c_5232_n ) capacitor c=0.00255985f \
 //x=53.055 //y=0.875 //x2=52.98 //y2=1.22
cc_291 ( N_GND_c_14_p N_noxref_15_c_5233_n ) capacitor c=0.00195164f //x=52.17 \
 //y=0 //x2=52.98 //y2=1.53
cc_292 ( N_GND_c_14_p N_noxref_15_c_5234_n ) capacitor c=0.0112696f //x=52.17 \
 //y=0 //x2=52.98 //y2=1.915
cc_293 ( N_GND_M32_noxref_d N_noxref_15_c_5235_n ) capacitor c=0.0131341f \
 //x=53.055 //y=0.875 //x2=53.355 //y2=0.72
cc_294 ( N_GND_M32_noxref_d N_noxref_15_c_5236_n ) capacitor c=0.00193146f \
 //x=53.055 //y=0.875 //x2=53.355 //y2=1.375
cc_295 ( N_GND_c_295_p N_noxref_15_c_5237_n ) capacitor c=0.00129018f \
 //x=56.81 //y=0 //x2=53.51 //y2=0.875
cc_296 ( N_GND_M32_noxref_d N_noxref_15_c_5237_n ) capacitor c=0.00257848f \
 //x=53.055 //y=0.875 //x2=53.51 //y2=0.875
cc_297 ( N_GND_M32_noxref_d N_noxref_15_c_5239_n ) capacitor c=0.00255985f \
 //x=53.055 //y=0.875 //x2=53.51 //y2=1.22
cc_298 ( N_GND_c_298_p N_noxref_15_c_5240_n ) capacitor c=0.00132755f \
 //x=57.97 //y=0 //x2=57.79 //y2=0.875
cc_299 ( N_GND_M35_noxref_d N_noxref_15_c_5240_n ) capacitor c=0.00211996f \
 //x=57.865 //y=0.875 //x2=57.79 //y2=0.875
cc_300 ( N_GND_M35_noxref_d N_noxref_15_c_5242_n ) capacitor c=0.00255985f \
 //x=57.865 //y=0.875 //x2=57.79 //y2=1.22
cc_301 ( N_GND_c_15_p N_noxref_15_c_5243_n ) capacitor c=0.00204716f //x=56.98 \
 //y=0 //x2=57.79 //y2=1.53
cc_302 ( N_GND_c_15_p N_noxref_15_c_5244_n ) capacitor c=0.0110952f //x=56.98 \
 //y=0 //x2=57.79 //y2=1.915
cc_303 ( N_GND_M35_noxref_d N_noxref_15_c_5245_n ) capacitor c=0.0131341f \
 //x=57.865 //y=0.875 //x2=58.165 //y2=0.72
cc_304 ( N_GND_M35_noxref_d N_noxref_15_c_5246_n ) capacitor c=0.00193146f \
 //x=57.865 //y=0.875 //x2=58.165 //y2=1.375
cc_305 ( N_GND_c_305_p N_noxref_15_c_5247_n ) capacitor c=0.00129018f \
 //x=61.62 //y=0 //x2=58.32 //y2=0.875
cc_306 ( N_GND_M35_noxref_d N_noxref_15_c_5247_n ) capacitor c=0.00257848f \
 //x=57.865 //y=0.875 //x2=58.32 //y2=0.875
cc_307 ( N_GND_M35_noxref_d N_noxref_15_c_5249_n ) capacitor c=0.00255985f \
 //x=57.865 //y=0.875 //x2=58.32 //y2=1.22
cc_308 ( N_GND_c_13_p N_noxref_15_M31_noxref_d ) capacitor c=8.58106e-19 \
 //x=48.84 //y=0 //x2=50.8 //y2=0.905
cc_309 ( N_GND_c_14_p N_noxref_15_M31_noxref_d ) capacitor c=0.00616547f \
 //x=52.17 //y=0 //x2=50.8 //y2=0.905
cc_310 ( N_GND_M30_noxref_d N_noxref_15_M31_noxref_d ) capacitor c=0.00143464f \
 //x=49.83 //y=0.865 //x2=50.8 //y2=0.905
cc_311 ( N_GND_c_16_p N_noxref_16_c_5458_n ) capacitor c=0.0222748f //x=61.79 \
 //y=0 //x2=62.785 //y2=2.59
cc_312 ( N_GND_c_16_p N_noxref_16_c_5459_n ) capacitor c=0.00102529f //x=61.79 \
 //y=0 //x2=61.165 //y2=2.59
cc_313 ( N_GND_c_16_p N_noxref_16_c_5460_n ) capacitor c=0.0401238f //x=61.79 \
 //y=0 //x2=60.965 //y2=1.665
cc_314 ( N_GND_c_16_p N_noxref_16_c_5461_n ) capacitor c=5.56859e-19 //x=61.79 \
 //y=0 //x2=61.05 //y2=2.59
cc_315 ( N_GND_c_16_p N_noxref_16_c_5462_n ) capacitor c=0.0128176f //x=61.79 \
 //y=0 //x2=62.9 //y2=2.08
cc_316 ( N_GND_c_316_p N_noxref_16_c_5463_n ) capacitor c=0.00135046f \
 //x=62.885 //y=0 //x2=62.705 //y2=0.865
cc_317 ( N_GND_M38_noxref_d N_noxref_16_c_5463_n ) capacitor c=0.00220047f \
 //x=62.78 //y=0.865 //x2=62.705 //y2=0.865
cc_318 ( N_GND_M38_noxref_d N_noxref_16_c_5465_n ) capacitor c=0.00255985f \
 //x=62.78 //y=0.865 //x2=62.705 //y2=1.21
cc_319 ( N_GND_c_16_p N_noxref_16_c_5466_n ) capacitor c=0.00189421f //x=61.79 \
 //y=0 //x2=62.705 //y2=1.52
cc_320 ( N_GND_c_16_p N_noxref_16_c_5467_n ) capacitor c=0.00992619f //x=61.79 \
 //y=0 //x2=62.705 //y2=1.915
cc_321 ( N_GND_M38_noxref_d N_noxref_16_c_5468_n ) capacitor c=0.0131326f \
 //x=62.78 //y=0.865 //x2=63.08 //y2=0.71
cc_322 ( N_GND_M38_noxref_d N_noxref_16_c_5469_n ) capacitor c=0.00193127f \
 //x=62.78 //y=0.865 //x2=63.08 //y2=1.365
cc_323 ( N_GND_c_323_p N_noxref_16_c_5470_n ) capacitor c=0.00130622f \
 //x=64.95 //y=0 //x2=63.235 //y2=0.865
cc_324 ( N_GND_M38_noxref_d N_noxref_16_c_5470_n ) capacitor c=0.00257848f \
 //x=62.78 //y=0.865 //x2=63.235 //y2=0.865
cc_325 ( N_GND_M38_noxref_d N_noxref_16_c_5472_n ) capacitor c=0.00255985f \
 //x=62.78 //y=0.865 //x2=63.235 //y2=1.21
cc_326 ( N_GND_c_16_p N_noxref_16_M37_noxref_d ) capacitor c=0.00591582f \
 //x=61.79 //y=0 //x2=60.375 //y2=0.915
cc_327 ( N_GND_c_2_p N_CLK_c_5622_n ) capacitor c=7.5188e-19 //x=3.33 //y=0 \
 //x2=5.55 //y2=2.08
cc_328 ( N_GND_c_4_p N_CLK_c_5623_n ) capacitor c=9.18594e-19 //x=12.95 //y=0 \
 //x2=14.8 //y2=2.08
cc_329 ( N_GND_c_5_p N_CLK_c_5623_n ) capacitor c=0.00110048f //x=16.28 //y=0 \
 //x2=14.8 //y2=2.08
cc_330 ( N_GND_c_8_p N_CLK_c_5625_n ) capacitor c=5.62272e-19 //x=27.75 //y=0 \
 //x2=29.97 //y2=2.08
cc_331 ( N_GND_c_10_p N_CLK_c_5626_n ) capacitor c=9.18594e-19 //x=37.37 //y=0 \
 //x2=39.22 //y2=2.08
cc_332 ( N_GND_c_11_p N_CLK_c_5626_n ) capacitor c=0.00110048f //x=40.7 //y=0 \
 //x2=39.22 //y2=2.08
cc_333 ( N_GND_c_14_p N_CLK_c_5628_n ) capacitor c=5.62272e-19 //x=52.17 //y=0 \
 //x2=54.39 //y2=2.08
cc_334 ( N_GND_c_16_p N_CLK_c_5629_n ) capacitor c=9.18594e-19 //x=61.79 //y=0 \
 //x2=63.64 //y2=2.08
cc_335 ( N_GND_c_17_p N_CLK_c_5629_n ) capacitor c=0.00110048f //x=65.12 //y=0 \
 //x2=63.64 //y2=2.08
cc_336 ( N_GND_c_13_p N_noxref_18_c_6377_n ) capacitor c=6.2409e-19 //x=48.84 \
 //y=0 //x2=50.69 //y2=2.08
cc_337 ( N_GND_c_14_p N_noxref_18_c_6377_n ) capacitor c=6.26561e-19 //x=52.17 \
 //y=0 //x2=50.69 //y2=2.08
cc_338 ( N_GND_c_15_p N_noxref_18_c_6379_n ) capacitor c=0.0401588f //x=56.98 \
 //y=0 //x2=56.155 //y2=1.665
cc_339 ( N_GND_c_17_p N_noxref_18_c_6380_n ) capacitor c=0.0154414f //x=65.12 \
 //y=0 //x2=66.23 //y2=2.08
cc_340 ( N_GND_c_340_p N_noxref_18_c_6381_n ) capacitor c=0.00135046f \
 //x=66.215 //y=0 //x2=66.035 //y2=0.865
cc_341 ( N_GND_M40_noxref_d N_noxref_18_c_6381_n ) capacitor c=0.00220047f \
 //x=66.11 //y=0.865 //x2=66.035 //y2=0.865
cc_342 ( N_GND_M40_noxref_d N_noxref_18_c_6383_n ) capacitor c=0.00255985f \
 //x=66.11 //y=0.865 //x2=66.035 //y2=1.21
cc_343 ( N_GND_c_17_p N_noxref_18_c_6384_n ) capacitor c=0.0018059f //x=65.12 \
 //y=0 //x2=66.035 //y2=1.52
cc_344 ( N_GND_c_17_p N_noxref_18_c_6385_n ) capacitor c=0.0101006f //x=65.12 \
 //y=0 //x2=66.035 //y2=1.915
cc_345 ( N_GND_M40_noxref_d N_noxref_18_c_6386_n ) capacitor c=0.0131326f \
 //x=66.11 //y=0.865 //x2=66.41 //y2=0.71
cc_346 ( N_GND_M40_noxref_d N_noxref_18_c_6387_n ) capacitor c=0.00193127f \
 //x=66.11 //y=0.865 //x2=66.41 //y2=1.365
cc_347 ( N_GND_c_347_p N_noxref_18_c_6388_n ) capacitor c=0.00130622f \
 //x=68.28 //y=0 //x2=66.565 //y2=0.865
cc_348 ( N_GND_M40_noxref_d N_noxref_18_c_6388_n ) capacitor c=0.00257848f \
 //x=66.11 //y=0.865 //x2=66.565 //y2=0.865
cc_349 ( N_GND_M40_noxref_d N_noxref_18_c_6390_n ) capacitor c=0.00255985f \
 //x=66.11 //y=0.865 //x2=66.565 //y2=1.21
cc_350 ( N_GND_c_15_p N_noxref_18_M34_noxref_d ) capacitor c=0.00591582f \
 //x=56.98 //y=0 //x2=55.565 //y2=0.915
cc_351 ( N_GND_c_18_p N_noxref_19_c_6668_n ) capacitor c=0.0435299f //x=68.45 \
 //y=0 //x2=67.625 //y2=1.655
cc_352 ( N_GND_c_17_p N_noxref_19_c_6669_n ) capacitor c=9.64732e-19 //x=65.12 \
 //y=0 //x2=67.71 //y2=4.81
cc_353 ( N_GND_c_18_p N_noxref_19_c_6670_n ) capacitor c=0.0156304f //x=68.45 \
 //y=0 //x2=69.56 //y2=2.08
cc_354 ( N_GND_c_354_p N_noxref_19_c_6671_n ) capacitor c=0.00132755f \
 //x=69.44 //y=0 //x2=69.26 //y2=0.875
cc_355 ( N_GND_M42_noxref_d N_noxref_19_c_6671_n ) capacitor c=0.00211996f \
 //x=69.335 //y=0.875 //x2=69.26 //y2=0.875
cc_356 ( N_GND_M42_noxref_d N_noxref_19_c_6673_n ) capacitor c=0.00255985f \
 //x=69.335 //y=0.875 //x2=69.26 //y2=1.22
cc_357 ( N_GND_c_18_p N_noxref_19_c_6674_n ) capacitor c=0.00195164f //x=68.45 \
 //y=0 //x2=69.26 //y2=1.53
cc_358 ( N_GND_c_18_p N_noxref_19_c_6675_n ) capacitor c=0.0110952f //x=68.45 \
 //y=0 //x2=69.26 //y2=1.915
cc_359 ( N_GND_M42_noxref_d N_noxref_19_c_6676_n ) capacitor c=0.0131341f \
 //x=69.335 //y=0.875 //x2=69.635 //y2=0.72
cc_360 ( N_GND_M42_noxref_d N_noxref_19_c_6677_n ) capacitor c=0.00193146f \
 //x=69.335 //y=0.875 //x2=69.635 //y2=1.375
cc_361 ( N_GND_c_212_p N_noxref_19_c_6678_n ) capacitor c=0.00129018f \
 //x=73.09 //y=0 //x2=69.79 //y2=0.875
cc_362 ( N_GND_M42_noxref_d N_noxref_19_c_6678_n ) capacitor c=0.00257848f \
 //x=69.335 //y=0.875 //x2=69.79 //y2=0.875
cc_363 ( N_GND_M42_noxref_d N_noxref_19_c_6680_n ) capacitor c=0.00255985f \
 //x=69.335 //y=0.875 //x2=69.79 //y2=1.22
cc_364 ( N_GND_c_17_p N_noxref_19_M41_noxref_d ) capacitor c=8.58106e-19 \
 //x=65.12 //y=0 //x2=67.08 //y2=0.905
cc_365 ( N_GND_c_18_p N_noxref_19_M41_noxref_d ) capacitor c=0.00616547f \
 //x=68.45 //y=0 //x2=67.08 //y2=0.905
cc_366 ( N_GND_M40_noxref_d N_noxref_19_M41_noxref_d ) capacitor c=0.00143464f \
 //x=66.11 //y=0.865 //x2=67.08 //y2=0.905
cc_367 ( N_GND_c_24_p N_SN_c_6833_n ) capacitor c=0.106954f //x=84.73 //y=0 \
 //x2=21.715 //y2=2.22
cc_368 ( N_GND_c_58_p N_SN_c_6833_n ) capacitor c=0.00447829f //x=12.78 //y=0 \
 //x2=21.715 //y2=2.22
cc_369 ( N_GND_c_69_p N_SN_c_6833_n ) capacitor c=0.00347653f //x=14.045 //y=0 \
 //x2=21.715 //y2=2.22
cc_370 ( N_GND_c_76_p N_SN_c_6833_n ) capacitor c=0.00411932f //x=16.11 //y=0 \
 //x2=21.715 //y2=2.22
cc_371 ( N_GND_c_84_p N_SN_c_6833_n ) capacitor c=0.00347653f //x=17.375 //y=0 \
 //x2=21.715 //y2=2.22
cc_372 ( N_GND_c_91_p N_SN_c_6833_n ) capacitor c=0.00411932f //x=19.44 //y=0 \
 //x2=21.715 //y2=2.22
cc_373 ( N_GND_c_98_p N_SN_c_6833_n ) capacitor c=0.00274252f //x=20.6 //y=0 \
 //x2=21.715 //y2=2.22
cc_374 ( N_GND_c_4_p N_SN_c_6833_n ) capacitor c=0.0379964f //x=12.95 //y=0 \
 //x2=21.715 //y2=2.22
cc_375 ( N_GND_c_5_p N_SN_c_6833_n ) capacitor c=0.0401775f //x=16.28 //y=0 \
 //x2=21.715 //y2=2.22
cc_376 ( N_GND_c_6_p N_SN_c_6833_n ) capacitor c=0.0401775f //x=19.61 //y=0 \
 //x2=21.715 //y2=2.22
cc_377 ( N_GND_c_24_p N_SN_c_6843_n ) capacitor c=0.0019104f //x=84.73 //y=0 \
 //x2=10.475 //y2=2.22
cc_378 ( N_GND_c_24_p N_SN_c_6844_n ) capacitor c=0.121058f //x=84.73 //y=0 \
 //x2=34.665 //y2=2.22
cc_379 ( N_GND_c_105_p N_SN_c_6844_n ) capacitor c=0.00447829f //x=24.25 //y=0 \
 //x2=34.665 //y2=2.22
cc_380 ( N_GND_c_259_p N_SN_c_6844_n ) capacitor c=0.00347653f //x=25.515 \
 //y=0 //x2=34.665 //y2=2.22
cc_381 ( N_GND_c_266_p N_SN_c_6844_n ) capacitor c=0.00411932f //x=27.58 //y=0 \
 //x2=34.665 //y2=2.22
cc_382 ( N_GND_c_128_p N_SN_c_6844_n ) capacitor c=0.00274252f //x=28.74 //y=0 \
 //x2=34.665 //y2=2.22
cc_383 ( N_GND_c_135_p N_SN_c_6844_n ) capacitor c=0.00450506f //x=32.39 //y=0 \
 //x2=34.665 //y2=2.22
cc_384 ( N_GND_c_138_p N_SN_c_6844_n ) capacitor c=0.00274252f //x=33.55 //y=0 \
 //x2=34.665 //y2=2.22
cc_385 ( N_GND_c_7_p N_SN_c_6844_n ) capacitor c=0.0401775f //x=24.42 //y=0 \
 //x2=34.665 //y2=2.22
cc_386 ( N_GND_c_8_p N_SN_c_6844_n ) capacitor c=0.0379964f //x=27.75 //y=0 \
 //x2=34.665 //y2=2.22
cc_387 ( N_GND_c_9_p N_SN_c_6844_n ) capacitor c=0.0379964f //x=32.56 //y=0 \
 //x2=34.665 //y2=2.22
cc_388 ( N_GND_c_24_p N_SN_c_6854_n ) capacitor c=0.00168059f //x=84.73 //y=0 \
 //x2=21.945 //y2=2.22
cc_389 ( N_GND_c_24_p N_SN_c_6855_n ) capacitor c=0.106954f //x=84.73 //y=0 \
 //x2=46.135 //y2=2.22
cc_390 ( N_GND_c_145_p N_SN_c_6855_n ) capacitor c=0.00447829f //x=37.2 //y=0 \
 //x2=46.135 //y2=2.22
cc_391 ( N_GND_c_156_p N_SN_c_6855_n ) capacitor c=0.00347653f //x=38.465 \
 //y=0 //x2=46.135 //y2=2.22
cc_392 ( N_GND_c_163_p N_SN_c_6855_n ) capacitor c=0.00411932f //x=40.53 //y=0 \
 //x2=46.135 //y2=2.22
cc_393 ( N_GND_c_171_p N_SN_c_6855_n ) capacitor c=0.00347653f //x=41.795 \
 //y=0 //x2=46.135 //y2=2.22
cc_394 ( N_GND_c_178_p N_SN_c_6855_n ) capacitor c=0.00411932f //x=43.86 //y=0 \
 //x2=46.135 //y2=2.22
cc_395 ( N_GND_c_188_p N_SN_c_6855_n ) capacitor c=0.00274252f //x=45.02 //y=0 \
 //x2=46.135 //y2=2.22
cc_396 ( N_GND_c_10_p N_SN_c_6855_n ) capacitor c=0.0379964f //x=37.37 //y=0 \
 //x2=46.135 //y2=2.22
cc_397 ( N_GND_c_11_p N_SN_c_6855_n ) capacitor c=0.0401775f //x=40.7 //y=0 \
 //x2=46.135 //y2=2.22
cc_398 ( N_GND_c_12_p N_SN_c_6855_n ) capacitor c=0.0379964f //x=44.03 //y=0 \
 //x2=46.135 //y2=2.22
cc_399 ( N_GND_c_24_p N_SN_c_6865_n ) capacitor c=0.00168059f //x=84.73 //y=0 \
 //x2=34.895 //y2=2.22
cc_400 ( N_GND_c_24_p N_SN_c_6866_n ) capacitor c=0.121058f //x=84.73 //y=0 \
 //x2=59.085 //y2=2.22
cc_401 ( N_GND_c_195_p N_SN_c_6866_n ) capacitor c=0.00447829f //x=48.67 //y=0 \
 //x2=59.085 //y2=2.22
cc_402 ( N_GND_c_269_p N_SN_c_6866_n ) capacitor c=0.00347653f //x=49.935 \
 //y=0 //x2=59.085 //y2=2.22
cc_403 ( N_GND_c_276_p N_SN_c_6866_n ) capacitor c=0.00411932f //x=52 //y=0 \
 //x2=59.085 //y2=2.22
cc_404 ( N_GND_c_288_p N_SN_c_6866_n ) capacitor c=0.00274252f //x=53.16 //y=0 \
 //x2=59.085 //y2=2.22
cc_405 ( N_GND_c_295_p N_SN_c_6866_n ) capacitor c=0.00450506f //x=56.81 //y=0 \
 //x2=59.085 //y2=2.22
cc_406 ( N_GND_c_298_p N_SN_c_6866_n ) capacitor c=0.00274252f //x=57.97 //y=0 \
 //x2=59.085 //y2=2.22
cc_407 ( N_GND_c_13_p N_SN_c_6866_n ) capacitor c=0.0379964f //x=48.84 //y=0 \
 //x2=59.085 //y2=2.22
cc_408 ( N_GND_c_14_p N_SN_c_6866_n ) capacitor c=0.0379964f //x=52.17 //y=0 \
 //x2=59.085 //y2=2.22
cc_409 ( N_GND_c_15_p N_SN_c_6866_n ) capacitor c=0.0379964f //x=56.98 //y=0 \
 //x2=59.085 //y2=2.22
cc_410 ( N_GND_c_24_p N_SN_c_6876_n ) capacitor c=0.00168059f //x=84.73 //y=0 \
 //x2=46.365 //y2=2.22
cc_411 ( N_GND_c_24_p N_SN_c_6877_n ) capacitor c=0.108864f //x=84.73 //y=0 \
 //x2=70.555 //y2=2.22
cc_412 ( N_GND_c_305_p N_SN_c_6877_n ) capacitor c=0.00447829f //x=61.62 //y=0 \
 //x2=70.555 //y2=2.22
cc_413 ( N_GND_c_316_p N_SN_c_6877_n ) capacitor c=0.00347653f //x=62.885 \
 //y=0 //x2=70.555 //y2=2.22
cc_414 ( N_GND_c_323_p N_SN_c_6877_n ) capacitor c=0.00411932f //x=64.95 //y=0 \
 //x2=70.555 //y2=2.22
cc_415 ( N_GND_c_340_p N_SN_c_6877_n ) capacitor c=0.00347653f //x=66.215 \
 //y=0 //x2=70.555 //y2=2.22
cc_416 ( N_GND_c_347_p N_SN_c_6877_n ) capacitor c=0.00411932f //x=68.28 //y=0 \
 //x2=70.555 //y2=2.22
cc_417 ( N_GND_c_354_p N_SN_c_6877_n ) capacitor c=0.00274252f //x=69.44 //y=0 \
 //x2=70.555 //y2=2.22
cc_418 ( N_GND_c_16_p N_SN_c_6877_n ) capacitor c=0.0379964f //x=61.79 //y=0 \
 //x2=70.555 //y2=2.22
cc_419 ( N_GND_c_17_p N_SN_c_6877_n ) capacitor c=0.0401775f //x=65.12 //y=0 \
 //x2=70.555 //y2=2.22
cc_420 ( N_GND_c_18_p N_SN_c_6877_n ) capacitor c=0.0401775f //x=68.45 //y=0 \
 //x2=70.555 //y2=2.22
cc_421 ( N_GND_c_24_p N_SN_c_6887_n ) capacitor c=0.00168059f //x=84.73 //y=0 \
 //x2=59.315 //y2=2.22
cc_422 ( N_GND_c_3_p N_SN_c_6888_n ) capacitor c=9.83618e-19 //x=8.14 //y=0 \
 //x2=10.36 //y2=2.08
cc_423 ( N_GND_c_6_p N_SN_c_6889_n ) capacitor c=5.94159e-19 //x=19.61 //y=0 \
 //x2=21.83 //y2=2.08
cc_424 ( N_GND_c_9_p N_SN_c_6890_n ) capacitor c=7.57155e-19 //x=32.56 //y=0 \
 //x2=34.78 //y2=2.08
cc_425 ( N_GND_c_12_p N_SN_c_6891_n ) capacitor c=7.57155e-19 //x=44.03 //y=0 \
 //x2=46.25 //y2=2.08
cc_426 ( N_GND_c_15_p N_SN_c_6892_n ) capacitor c=7.57155e-19 //x=56.98 //y=0 \
 //x2=59.2 //y2=2.08
cc_427 ( N_GND_c_18_p N_SN_c_6893_n ) capacitor c=5.94159e-19 //x=68.45 //y=0 \
 //x2=70.67 //y2=2.08
cc_428 ( N_GND_c_15_p N_noxref_21_c_7648_n ) capacitor c=6.12031e-19 //x=56.98 \
 //y=0 //x2=55.5 //y2=2.08
cc_429 ( N_GND_c_16_p N_noxref_21_c_7649_n ) capacitor c=0.00101012f //x=61.79 \
 //y=0 //x2=60.31 //y2=2.08
cc_430 ( N_GND_c_17_p N_noxref_21_c_7650_n ) capacitor c=0.0432305f //x=65.12 \
 //y=0 //x2=64.295 //y2=1.655
cc_431 ( N_GND_c_16_p N_noxref_21_c_7651_n ) capacitor c=9.64732e-19 //x=61.79 \
 //y=0 //x2=64.38 //y2=3.7
cc_432 ( N_GND_c_19_p N_noxref_21_c_7652_n ) capacitor c=0.00128267f //x=73.26 \
 //y=0 //x2=71.78 //y2=2.08
cc_433 ( N_GND_c_16_p N_noxref_21_M39_noxref_d ) capacitor c=8.58106e-19 \
 //x=61.79 //y=0 //x2=63.75 //y2=0.905
cc_434 ( N_GND_c_17_p N_noxref_21_M39_noxref_d ) capacitor c=0.00616547f \
 //x=65.12 //y=0 //x2=63.75 //y2=0.905
cc_435 ( N_GND_M38_noxref_d N_noxref_21_M39_noxref_d ) capacitor c=0.00143464f \
 //x=62.78 //y=0.865 //x2=63.75 //y2=0.905
cc_436 ( N_GND_c_17_p N_noxref_23_c_8060_n ) capacitor c=7.1088e-19 //x=65.12 \
 //y=0 //x2=66.97 //y2=2.08
cc_437 ( N_GND_c_18_p N_noxref_23_c_8060_n ) capacitor c=7.76678e-19 //x=68.45 \
 //y=0 //x2=66.97 //y2=2.08
cc_438 ( N_GND_c_19_p N_noxref_23_c_8062_n ) capacitor c=0.0455602f //x=73.26 \
 //y=0 //x2=72.435 //y2=1.665
cc_439 ( N_GND_c_24_p N_noxref_23_c_8063_n ) capacitor c=2.98913e-19 //x=84.73 \
 //y=0 //x2=74 //y2=2.08
cc_440 ( N_GND_c_19_p N_noxref_23_c_8063_n ) capacitor c=0.0291009f //x=73.26 \
 //y=0 //x2=74 //y2=2.08
cc_441 ( N_GND_c_20_p N_noxref_23_c_8063_n ) capacitor c=3.10504e-19 //x=76.59 \
 //y=0 //x2=74 //y2=2.08
cc_442 ( N_GND_c_20_p N_noxref_23_c_8066_n ) capacitor c=0.0178945f //x=76.59 \
 //y=0 //x2=77.7 //y2=2.08
cc_443 ( N_GND_c_21_p N_noxref_23_c_8066_n ) capacitor c=7.87427e-19 //x=79.92 \
 //y=0 //x2=77.7 //y2=2.08
cc_444 ( N_GND_c_213_p N_noxref_23_c_8068_n ) capacitor c=0.0013864f \
 //x=74.355 //y=0 //x2=74.175 //y2=0.865
cc_445 ( N_GND_M45_noxref_d N_noxref_23_c_8068_n ) capacitor c=0.00220047f \
 //x=74.25 //y=0.865 //x2=74.175 //y2=0.865
cc_446 ( N_GND_M45_noxref_d N_noxref_23_c_8070_n ) capacitor c=0.00255985f \
 //x=74.25 //y=0.865 //x2=74.175 //y2=1.21
cc_447 ( N_GND_c_19_p N_noxref_23_c_8071_n ) capacitor c=0.00189421f //x=73.26 \
 //y=0 //x2=74.175 //y2=1.52
cc_448 ( N_GND_c_19_p N_noxref_23_c_8072_n ) capacitor c=0.00369987f //x=73.26 \
 //y=0 //x2=74.175 //y2=1.915
cc_449 ( N_GND_M45_noxref_d N_noxref_23_c_8073_n ) capacitor c=0.0131326f \
 //x=74.25 //y=0.865 //x2=74.55 //y2=0.71
cc_450 ( N_GND_M45_noxref_d N_noxref_23_c_8074_n ) capacitor c=0.00193127f \
 //x=74.25 //y=0.865 //x2=74.55 //y2=1.365
cc_451 ( N_GND_c_451_p N_noxref_23_c_8075_n ) capacitor c=0.00130622f \
 //x=76.42 //y=0 //x2=74.705 //y2=0.865
cc_452 ( N_GND_M45_noxref_d N_noxref_23_c_8075_n ) capacitor c=0.00257848f \
 //x=74.25 //y=0.865 //x2=74.705 //y2=0.865
cc_453 ( N_GND_M45_noxref_d N_noxref_23_c_8077_n ) capacitor c=0.00255985f \
 //x=74.25 //y=0.865 //x2=74.705 //y2=1.21
cc_454 ( N_GND_c_454_p N_noxref_23_c_8078_n ) capacitor c=0.00135046f \
 //x=77.685 //y=0 //x2=77.505 //y2=0.865
cc_455 ( N_GND_M47_noxref_d N_noxref_23_c_8078_n ) capacitor c=0.00220047f \
 //x=77.58 //y=0.865 //x2=77.505 //y2=0.865
cc_456 ( N_GND_M47_noxref_d N_noxref_23_c_8080_n ) capacitor c=0.00272336f \
 //x=77.58 //y=0.865 //x2=77.505 //y2=1.21
cc_457 ( N_GND_c_20_p N_noxref_23_c_8081_n ) capacitor c=0.0100605f //x=76.59 \
 //y=0 //x2=77.505 //y2=1.915
cc_458 ( N_GND_M47_noxref_d N_noxref_23_c_8082_n ) capacitor c=0.0131326f \
 //x=77.58 //y=0.865 //x2=77.88 //y2=0.71
cc_459 ( N_GND_M47_noxref_d N_noxref_23_c_8083_n ) capacitor c=0.00167494f \
 //x=77.58 //y=0.865 //x2=77.88 //y2=1.365
cc_460 ( N_GND_c_460_p N_noxref_23_c_8084_n ) capacitor c=0.00130622f \
 //x=79.75 //y=0 //x2=78.035 //y2=0.865
cc_461 ( N_GND_M47_noxref_d N_noxref_23_c_8084_n ) capacitor c=0.00257848f \
 //x=77.58 //y=0.865 //x2=78.035 //y2=0.865
cc_462 ( N_GND_M47_noxref_d N_noxref_23_c_8086_n ) capacitor c=0.00272336f \
 //x=77.58 //y=0.865 //x2=78.035 //y2=1.21
cc_463 ( N_GND_c_19_p N_noxref_23_c_8087_n ) capacitor c=0.0096025f //x=73.26 \
 //y=0 //x2=74 //y2=2.08
cc_464 ( N_GND_c_19_p N_noxref_23_M44_noxref_d ) capacitor c=0.00591203f \
 //x=73.26 //y=0 //x2=71.845 //y2=0.915
cc_465 ( N_GND_c_24_p N_noxref_24_c_8424_n ) capacitor c=0.0224606f //x=84.73 \
 //y=0 //x2=79.065 //y2=3.33
cc_466 ( N_GND_c_20_p N_noxref_24_c_8424_n ) capacitor c=0.00731853f //x=76.59 \
 //y=0 //x2=79.065 //y2=3.33
cc_467 ( N_GND_c_21_p N_noxref_24_c_8426_n ) capacitor c=0.0396043f //x=79.92 \
 //y=0 //x2=80.545 //y2=2.08
cc_468 ( N_GND_c_21_p N_noxref_24_c_8427_n ) capacitor c=0.00128384f //x=79.92 \
 //y=0 //x2=79.295 //y2=2.08
cc_469 ( N_GND_c_5_p N_noxref_24_c_8428_n ) capacitor c=7.1088e-19 //x=16.28 \
 //y=0 //x2=18.13 //y2=2.08
cc_470 ( N_GND_c_6_p N_noxref_24_c_8428_n ) capacitor c=7.76678e-19 //x=19.61 \
 //y=0 //x2=18.13 //y2=2.08
cc_471 ( N_GND_c_7_p N_noxref_24_c_8430_n ) capacitor c=0.0429319f //x=24.42 \
 //y=0 //x2=23.595 //y2=1.665
cc_472 ( N_GND_c_20_p N_noxref_24_c_8431_n ) capacitor c=6.95291e-19 //x=76.59 \
 //y=0 //x2=79.18 //y2=2.08
cc_473 ( N_GND_c_21_p N_noxref_24_c_8431_n ) capacitor c=0.0266762f //x=79.92 \
 //y=0 //x2=79.18 //y2=2.08
cc_474 ( N_GND_c_21_p N_noxref_24_c_8433_n ) capacitor c=0.0266762f //x=79.92 \
 //y=0 //x2=80.66 //y2=2.08
cc_475 ( N_GND_c_21_p N_noxref_24_c_8434_n ) capacitor c=0.0103285f //x=79.92 \
 //y=0 //x2=79.005 //y2=1.915
cc_476 ( N_GND_c_476_p N_noxref_24_c_8435_n ) capacitor c=0.0013864f \
 //x=81.015 //y=0 //x2=80.835 //y2=0.865
cc_477 ( N_GND_M49_noxref_d N_noxref_24_c_8435_n ) capacitor c=0.00220047f \
 //x=80.91 //y=0.865 //x2=80.835 //y2=0.865
cc_478 ( N_GND_M49_noxref_d N_noxref_24_c_8437_n ) capacitor c=0.00272336f \
 //x=80.91 //y=0.865 //x2=80.835 //y2=1.21
cc_479 ( N_GND_c_21_p N_noxref_24_c_8438_n ) capacitor c=0.00369763f //x=79.92 \
 //y=0 //x2=80.835 //y2=1.915
cc_480 ( N_GND_M49_noxref_d N_noxref_24_c_8439_n ) capacitor c=0.0131326f \
 //x=80.91 //y=0.865 //x2=81.21 //y2=0.71
cc_481 ( N_GND_M49_noxref_d N_noxref_24_c_8440_n ) capacitor c=0.00167494f \
 //x=80.91 //y=0.865 //x2=81.21 //y2=1.365
cc_482 ( N_GND_c_482_p N_noxref_24_c_8441_n ) capacitor c=0.00130622f \
 //x=83.08 //y=0 //x2=81.365 //y2=0.865
cc_483 ( N_GND_M49_noxref_d N_noxref_24_c_8441_n ) capacitor c=0.00257848f \
 //x=80.91 //y=0.865 //x2=81.365 //y2=0.865
cc_484 ( N_GND_M49_noxref_d N_noxref_24_c_8443_n ) capacitor c=0.00272336f \
 //x=80.91 //y=0.865 //x2=81.365 //y2=1.21
cc_485 ( N_GND_c_21_p N_noxref_24_c_8444_n ) capacitor c=0.00662863f //x=79.92 \
 //y=0 //x2=80.66 //y2=2.08
cc_486 ( N_GND_c_7_p N_noxref_24_M14_noxref_d ) capacitor c=0.00591582f \
 //x=24.42 //y=0 //x2=23.005 //y2=0.915
cc_487 ( N_GND_c_24_p N_noxref_26_c_8988_n ) capacitor c=0.0695894f //x=84.73 \
 //y=0 //x2=78.625 //y2=1.18
cc_488 ( N_GND_c_451_p N_noxref_26_c_8988_n ) capacitor c=0.0081414f //x=76.42 \
 //y=0 //x2=78.625 //y2=1.18
cc_489 ( N_GND_c_454_p N_noxref_26_c_8988_n ) capacitor c=0.0101988f \
 //x=77.685 //y=0 //x2=78.625 //y2=1.18
cc_490 ( N_GND_c_460_p N_noxref_26_c_8988_n ) capacitor c=0.00469062f \
 //x=79.75 //y=0 //x2=78.625 //y2=1.18
cc_491 ( N_GND_c_20_p N_noxref_26_c_8988_n ) capacitor c=0.0420176f //x=76.59 \
 //y=0 //x2=78.625 //y2=1.18
cc_492 ( N_GND_c_23_p N_noxref_26_c_8988_n ) capacitor c=0.00131703f //x=84.85 \
 //y=0 //x2=78.625 //y2=1.18
cc_493 ( N_GND_M47_noxref_d N_noxref_26_c_8988_n ) capacitor c=0.00960943f \
 //x=77.58 //y=0.865 //x2=78.625 //y2=1.18
cc_494 ( N_GND_c_24_p N_noxref_26_c_8995_n ) capacitor c=0.00715563f //x=84.73 \
 //y=0 //x2=75.525 //y2=1.18
cc_495 ( N_GND_c_24_p N_noxref_26_c_8996_n ) capacitor c=0.0769193f //x=84.73 \
 //y=0 //x2=81.955 //y2=1.18
cc_496 ( N_GND_c_460_p N_noxref_26_c_8996_n ) capacitor c=0.00788597f \
 //x=79.75 //y=0 //x2=81.955 //y2=1.18
cc_497 ( N_GND_c_476_p N_noxref_26_c_8996_n ) capacitor c=0.00974891f \
 //x=81.015 //y=0 //x2=81.955 //y2=1.18
cc_498 ( N_GND_c_482_p N_noxref_26_c_8996_n ) capacitor c=0.00446008f \
 //x=83.08 //y=0 //x2=81.955 //y2=1.18
cc_499 ( N_GND_c_21_p N_noxref_26_c_8996_n ) capacitor c=0.0384312f //x=79.92 \
 //y=0 //x2=81.955 //y2=1.18
cc_500 ( N_GND_c_23_p N_noxref_26_c_8996_n ) capacitor c=0.00131703f //x=84.85 \
 //y=0 //x2=81.955 //y2=1.18
cc_501 ( N_GND_M49_noxref_d N_noxref_26_c_8996_n ) capacitor c=0.00960943f \
 //x=80.91 //y=0.865 //x2=81.955 //y2=1.18
cc_502 ( N_GND_c_24_p N_noxref_26_c_9003_n ) capacitor c=0.00664346f //x=84.73 \
 //y=0 //x2=78.855 //y2=1.18
cc_503 ( N_GND_c_24_p N_noxref_26_c_9004_n ) capacitor c=0.00899798f //x=84.73 \
 //y=0 //x2=83.875 //y2=4.07
cc_504 ( N_GND_c_22_p N_noxref_26_c_9004_n ) capacitor c=0.00363802f //x=83.25 \
 //y=0 //x2=83.875 //y2=4.07
cc_505 ( N_GND_M51_noxref_s N_noxref_26_c_9004_n ) capacitor c=9.50279e-19 \
 //x=83.745 //y=0.37 //x2=83.875 //y2=4.07
cc_506 ( N_GND_c_24_p N_noxref_26_c_9007_n ) capacitor c=0.00144743f //x=84.73 \
 //y=0 //x2=82.625 //y2=4.07
cc_507 ( N_GND_c_22_p N_noxref_26_c_9008_n ) capacitor c=0.0461307f //x=83.25 \
 //y=0 //x2=82.425 //y2=1.645
cc_508 ( N_GND_M51_noxref_s N_noxref_26_c_9008_n ) capacitor c=3.58337e-19 \
 //x=83.745 //y=0.37 //x2=82.425 //y2=1.645
cc_509 ( N_GND_c_21_p N_noxref_26_c_9010_n ) capacitor c=0.00109945f //x=79.92 \
 //y=0 //x2=82.51 //y2=4.07
cc_510 ( N_GND_c_24_p N_noxref_26_c_9011_n ) capacitor c=0.00187124f //x=84.73 \
 //y=0 //x2=83.99 //y2=2.085
cc_511 ( N_GND_c_511_p N_noxref_26_c_9011_n ) capacitor c=8.01092e-19 \
 //x=84.28 //y=0.535 //x2=83.99 //y2=2.085
cc_512 ( N_GND_c_22_p N_noxref_26_c_9011_n ) capacitor c=0.0290587f //x=83.25 \
 //y=0 //x2=83.99 //y2=2.085
cc_513 ( N_GND_c_23_p N_noxref_26_c_9011_n ) capacitor c=0.00118981f //x=84.85 \
 //y=0 //x2=83.99 //y2=2.085
cc_514 ( N_GND_M51_noxref_s N_noxref_26_c_9011_n ) capacitor c=0.0110172f \
 //x=83.745 //y=0.37 //x2=83.99 //y2=2.085
cc_515 ( N_GND_c_511_p N_noxref_26_c_9016_n ) capacitor c=0.0120496f //x=84.28 \
 //y=0.535 //x2=84.1 //y2=0.91
cc_516 ( N_GND_M51_noxref_s N_noxref_26_c_9016_n ) capacitor c=0.031817f \
 //x=83.745 //y=0.37 //x2=84.1 //y2=0.91
cc_517 ( N_GND_c_22_p N_noxref_26_c_9018_n ) capacitor c=0.00550606f //x=83.25 \
 //y=0 //x2=84.1 //y2=1.92
cc_518 ( N_GND_M51_noxref_s N_noxref_26_c_9019_n ) capacitor c=0.00483274f \
 //x=83.745 //y=0.37 //x2=84.475 //y2=0.755
cc_519 ( N_GND_c_519_p N_noxref_26_c_9020_n ) capacitor c=0.0118602f \
 //x=84.765 //y=0.535 //x2=84.63 //y2=0.91
cc_520 ( N_GND_M51_noxref_s N_noxref_26_c_9020_n ) capacitor c=0.0143355f \
 //x=83.745 //y=0.37 //x2=84.63 //y2=0.91
cc_521 ( N_GND_M51_noxref_s N_noxref_26_c_9022_n ) capacitor c=0.0074042f \
 //x=83.745 //y=0.37 //x2=84.63 //y2=1.255
cc_522 ( N_GND_c_511_p N_noxref_26_c_9023_n ) capacitor c=2.1838e-19 //x=84.28 \
 //y=0.535 //x2=83.99 //y2=2.085
cc_523 ( N_GND_c_22_p N_noxref_26_c_9023_n ) capacitor c=0.00864459f //x=83.25 \
 //y=0 //x2=83.99 //y2=2.085
cc_524 ( N_GND_M51_noxref_s N_noxref_26_c_9023_n ) capacitor c=0.00655738f \
 //x=83.745 //y=0.37 //x2=83.99 //y2=2.085
cc_525 ( N_GND_c_24_p N_noxref_26_M46_noxref_d ) capacitor c=2.00936e-19 \
 //x=84.73 //y=0 //x2=75.22 //y2=0.905
cc_526 ( N_GND_c_20_p N_noxref_26_M46_noxref_d ) capacitor c=0.00141366f \
 //x=76.59 //y=0 //x2=75.22 //y2=0.905
cc_527 ( N_GND_M45_noxref_d N_noxref_26_M46_noxref_d ) capacitor c=0.00128667f \
 //x=74.25 //y=0.865 //x2=75.22 //y2=0.905
cc_528 ( N_GND_c_24_p N_noxref_26_M48_noxref_d ) capacitor c=2.00936e-19 \
 //x=84.73 //y=0 //x2=78.55 //y2=0.905
cc_529 ( N_GND_c_21_p N_noxref_26_M48_noxref_d ) capacitor c=0.0014176f \
 //x=79.92 //y=0 //x2=78.55 //y2=0.905
cc_530 ( N_GND_M47_noxref_d N_noxref_26_M48_noxref_d ) capacitor c=0.0012247f \
 //x=77.58 //y=0.865 //x2=78.55 //y2=0.905
cc_531 ( N_GND_c_24_p N_noxref_26_M50_noxref_d ) capacitor c=2.00936e-19 \
 //x=84.73 //y=0 //x2=81.88 //y2=0.905
cc_532 ( N_GND_c_21_p N_noxref_26_M50_noxref_d ) capacitor c=8.62423e-19 \
 //x=79.92 //y=0 //x2=81.88 //y2=0.905
cc_533 ( N_GND_c_22_p N_noxref_26_M50_noxref_d ) capacitor c=0.00523456f \
 //x=83.25 //y=0 //x2=81.88 //y2=0.905
cc_534 ( N_GND_M49_noxref_d N_noxref_26_M50_noxref_d ) capacitor c=0.0012247f \
 //x=80.91 //y=0.865 //x2=81.88 //y2=0.905
cc_535 ( N_GND_c_24_p N_noxref_27_c_9228_n ) capacitor c=0.00576803f //x=84.73 \
 //y=0 //x2=1.58 //y2=1.58
cc_536 ( N_GND_c_249_p N_noxref_27_c_9228_n ) capacitor c=0.00111428f \
 //x=1.095 //y=0 //x2=1.58 //y2=1.58
cc_537 ( N_GND_c_25_p N_noxref_27_c_9228_n ) capacitor c=0.00182382f //x=3.16 \
 //y=0 //x2=1.58 //y2=1.58
cc_538 ( N_GND_M0_noxref_d N_noxref_27_c_9228_n ) capacitor c=0.00889643f \
 //x=0.99 //y=0.865 //x2=1.58 //y2=1.58
cc_539 ( N_GND_c_24_p N_noxref_27_c_9232_n ) capacitor c=0.00282937f //x=84.73 \
 //y=0 //x2=1.665 //y2=0.615
cc_540 ( N_GND_c_25_p N_noxref_27_c_9232_n ) capacitor c=0.0148639f //x=3.16 \
 //y=0 //x2=1.665 //y2=0.615
cc_541 ( N_GND_M0_noxref_d N_noxref_27_c_9232_n ) capacitor c=0.033812f \
 //x=0.99 //y=0.865 //x2=1.665 //y2=0.615
cc_542 ( N_GND_c_1_p N_noxref_27_c_9235_n ) capacitor c=2.91423e-19 //x=0.74 \
 //y=0 //x2=1.665 //y2=1.495
cc_543 ( N_GND_c_24_p N_noxref_27_c_9236_n ) capacitor c=0.0115707f //x=84.73 \
 //y=0 //x2=2.55 //y2=0.53
cc_544 ( N_GND_c_25_p N_noxref_27_c_9236_n ) capacitor c=0.037494f //x=3.16 \
 //y=0 //x2=2.55 //y2=0.53
cc_545 ( N_GND_c_24_p N_noxref_27_c_9238_n ) capacitor c=0.0027057f //x=84.73 \
 //y=0 //x2=2.635 //y2=0.615
cc_546 ( N_GND_c_25_p N_noxref_27_c_9238_n ) capacitor c=0.0147125f //x=3.16 \
 //y=0 //x2=2.635 //y2=0.615
cc_547 ( N_GND_c_2_p N_noxref_27_c_9238_n ) capacitor c=0.0431718f //x=3.33 \
 //y=0 //x2=2.635 //y2=0.615
cc_548 ( N_GND_c_24_p N_noxref_27_M0_noxref_s ) capacitor c=0.00723598f \
 //x=84.73 //y=0 //x2=0.56 //y2=0.365
cc_549 ( N_GND_c_249_p N_noxref_27_M0_noxref_s ) capacitor c=0.0146208f \
 //x=1.095 //y=0 //x2=0.56 //y2=0.365
cc_550 ( N_GND_c_1_p N_noxref_27_M0_noxref_s ) capacitor c=0.0594057f //x=0.74 \
 //y=0 //x2=0.56 //y2=0.365
cc_551 ( N_GND_c_2_p N_noxref_27_M0_noxref_s ) capacitor c=0.00198098f \
 //x=3.33 //y=0 //x2=0.56 //y2=0.365
cc_552 ( N_GND_M0_noxref_d N_noxref_27_M0_noxref_s ) capacitor c=0.0334197f \
 //x=0.99 //y=0.865 //x2=0.56 //y2=0.365
cc_553 ( N_GND_c_24_p N_noxref_28_c_9278_n ) capacitor c=0.00529429f //x=84.73 \
 //y=0 //x2=4.805 //y2=1.59
cc_554 ( N_GND_c_26_p N_noxref_28_c_9278_n ) capacitor c=0.00111496f //x=4.32 \
 //y=0 //x2=4.805 //y2=1.59
cc_555 ( N_GND_c_31_p N_noxref_28_c_9278_n ) capacitor c=0.0018066f //x=7.97 \
 //y=0 //x2=4.805 //y2=1.59
cc_556 ( N_GND_M2_noxref_d N_noxref_28_c_9278_n ) capacitor c=0.00868399f \
 //x=4.215 //y=0.875 //x2=4.805 //y2=1.59
cc_557 ( N_GND_c_24_p N_noxref_28_c_9282_n ) capacitor c=0.00266608f //x=84.73 \
 //y=0 //x2=4.89 //y2=0.625
cc_558 ( N_GND_c_31_p N_noxref_28_c_9282_n ) capacitor c=0.0141814f //x=7.97 \
 //y=0 //x2=4.89 //y2=0.625
cc_559 ( N_GND_M2_noxref_d N_noxref_28_c_9282_n ) capacitor c=0.033954f \
 //x=4.215 //y=0.875 //x2=4.89 //y2=0.625
cc_560 ( N_GND_c_24_p N_noxref_28_c_9285_n ) capacitor c=0.0109327f //x=84.73 \
 //y=0 //x2=5.775 //y2=0.54
cc_561 ( N_GND_c_31_p N_noxref_28_c_9285_n ) capacitor c=0.0361235f //x=7.97 \
 //y=0 //x2=5.775 //y2=0.54
cc_562 ( N_GND_c_24_p N_noxref_28_M2_noxref_s ) capacitor c=0.00532331f \
 //x=84.73 //y=0 //x2=3.785 //y2=0.375
cc_563 ( N_GND_c_26_p N_noxref_28_M2_noxref_s ) capacitor c=0.0141814f \
 //x=4.32 //y=0 //x2=3.785 //y2=0.375
cc_564 ( N_GND_c_31_p N_noxref_28_M2_noxref_s ) capacitor c=0.0132355f \
 //x=7.97 //y=0 //x2=3.785 //y2=0.375
cc_565 ( N_GND_c_2_p N_noxref_28_M2_noxref_s ) capacitor c=0.0696963f //x=3.33 \
 //y=0 //x2=3.785 //y2=0.375
cc_566 ( N_GND_c_3_p N_noxref_28_M2_noxref_s ) capacitor c=3.31601e-19 \
 //x=8.14 //y=0 //x2=3.785 //y2=0.375
cc_567 ( N_GND_M2_noxref_d N_noxref_28_M2_noxref_s ) capacitor c=0.033718f \
 //x=4.215 //y=0.875 //x2=3.785 //y2=0.375
cc_568 ( N_GND_c_24_p N_noxref_29_c_9329_n ) capacitor c=0.00364762f //x=84.73 \
 //y=0 //x2=6.345 //y2=0.995
cc_569 ( N_GND_c_31_p N_noxref_29_c_9329_n ) capacitor c=0.00940048f //x=7.97 \
 //y=0 //x2=6.345 //y2=0.995
cc_570 ( N_GND_c_24_p N_noxref_29_c_9331_n ) capacitor c=0.00266608f //x=84.73 \
 //y=0 //x2=6.43 //y2=0.625
cc_571 ( N_GND_c_31_p N_noxref_29_c_9331_n ) capacitor c=0.0141814f //x=7.97 \
 //y=0 //x2=6.43 //y2=0.625
cc_572 ( N_GND_M2_noxref_d N_noxref_29_c_9331_n ) capacitor c=6.21394e-19 \
 //x=4.215 //y=0.875 //x2=6.43 //y2=0.625
cc_573 ( N_GND_c_24_p N_noxref_29_c_9334_n ) capacitor c=0.0110095f //x=84.73 \
 //y=0 //x2=7.315 //y2=0.54
cc_574 ( N_GND_c_31_p N_noxref_29_c_9334_n ) capacitor c=0.0365163f //x=7.97 \
 //y=0 //x2=7.315 //y2=0.54
cc_575 ( N_GND_c_24_p N_noxref_29_c_9336_n ) capacitor c=0.00266421f //x=84.73 \
 //y=0 //x2=7.4 //y2=0.625
cc_576 ( N_GND_c_31_p N_noxref_29_c_9336_n ) capacitor c=0.0141195f //x=7.97 \
 //y=0 //x2=7.4 //y2=0.625
cc_577 ( N_GND_c_3_p N_noxref_29_c_9336_n ) capacitor c=0.0404137f //x=8.14 \
 //y=0 //x2=7.4 //y2=0.625
cc_578 ( N_GND_M2_noxref_d N_noxref_29_M3_noxref_d ) capacitor c=0.00162435f \
 //x=4.215 //y=0.875 //x2=5.19 //y2=0.91
cc_579 ( N_GND_c_2_p N_noxref_29_M4_noxref_s ) capacitor c=8.16352e-19 \
 //x=3.33 //y=0 //x2=6.295 //y2=0.375
cc_580 ( N_GND_c_3_p N_noxref_29_M4_noxref_s ) capacitor c=0.00180469f \
 //x=8.14 //y=0 //x2=6.295 //y2=0.375
cc_581 ( N_GND_c_24_p N_noxref_30_c_9381_n ) capacitor c=0.00532237f //x=84.73 \
 //y=0 //x2=9.615 //y2=1.59
cc_582 ( N_GND_c_32_p N_noxref_30_c_9381_n ) capacitor c=0.00111496f //x=9.13 \
 //y=0 //x2=9.615 //y2=1.59
cc_583 ( N_GND_c_58_p N_noxref_30_c_9381_n ) capacitor c=0.00180702f //x=12.78 \
 //y=0 //x2=9.615 //y2=1.59
cc_584 ( N_GND_M5_noxref_d N_noxref_30_c_9381_n ) capacitor c=0.00868586f \
 //x=9.025 //y=0.875 //x2=9.615 //y2=1.59
cc_585 ( N_GND_c_24_p N_noxref_30_c_9385_n ) capacitor c=0.00277579f //x=84.73 \
 //y=0 //x2=9.7 //y2=0.625
cc_586 ( N_GND_c_58_p N_noxref_30_c_9385_n ) capacitor c=0.0142586f //x=12.78 \
 //y=0 //x2=9.7 //y2=0.625
cc_587 ( N_GND_M5_noxref_d N_noxref_30_c_9385_n ) capacitor c=0.033954f \
 //x=9.025 //y=0.875 //x2=9.7 //y2=0.625
cc_588 ( N_GND_c_24_p N_noxref_30_c_9388_n ) capacitor c=0.0109321f //x=84.73 \
 //y=0 //x2=10.585 //y2=0.54
cc_589 ( N_GND_c_58_p N_noxref_30_c_9388_n ) capacitor c=0.0361222f //x=12.78 \
 //y=0 //x2=10.585 //y2=0.54
cc_590 ( N_GND_c_24_p N_noxref_30_M5_noxref_s ) capacitor c=0.00519789f \
 //x=84.73 //y=0 //x2=8.595 //y2=0.375
cc_591 ( N_GND_c_32_p N_noxref_30_M5_noxref_s ) capacitor c=0.0141814f \
 //x=9.13 //y=0 //x2=8.595 //y2=0.375
cc_592 ( N_GND_c_58_p N_noxref_30_M5_noxref_s ) capacitor c=0.0136651f \
 //x=12.78 //y=0 //x2=8.595 //y2=0.375
cc_593 ( N_GND_c_3_p N_noxref_30_M5_noxref_s ) capacitor c=0.0696963f //x=8.14 \
 //y=0 //x2=8.595 //y2=0.375
cc_594 ( N_GND_c_4_p N_noxref_30_M5_noxref_s ) capacitor c=3.31601e-19 \
 //x=12.95 //y=0 //x2=8.595 //y2=0.375
cc_595 ( N_GND_M5_noxref_d N_noxref_30_M5_noxref_s ) capacitor c=0.033718f \
 //x=9.025 //y=0.875 //x2=8.595 //y2=0.375
cc_596 ( N_GND_c_24_p N_noxref_31_c_9434_n ) capacitor c=0.00352952f //x=84.73 \
 //y=0 //x2=11.155 //y2=0.995
cc_597 ( N_GND_c_58_p N_noxref_31_c_9434_n ) capacitor c=0.00934524f //x=12.78 \
 //y=0 //x2=11.155 //y2=0.995
cc_598 ( N_GND_c_24_p N_noxref_31_c_9436_n ) capacitor c=0.00254475f //x=84.73 \
 //y=0 //x2=11.24 //y2=0.625
cc_599 ( N_GND_c_58_p N_noxref_31_c_9436_n ) capacitor c=0.0140928f //x=12.78 \
 //y=0 //x2=11.24 //y2=0.625
cc_600 ( N_GND_M5_noxref_d N_noxref_31_c_9436_n ) capacitor c=6.21394e-19 \
 //x=9.025 //y=0.875 //x2=11.24 //y2=0.625
cc_601 ( N_GND_c_24_p N_noxref_31_c_9439_n ) capacitor c=0.0105317f //x=84.73 \
 //y=0 //x2=12.125 //y2=0.54
cc_602 ( N_GND_c_58_p N_noxref_31_c_9439_n ) capacitor c=0.0364215f //x=12.78 \
 //y=0 //x2=12.125 //y2=0.54
cc_603 ( N_GND_c_24_p N_noxref_31_c_9441_n ) capacitor c=0.00254232f //x=84.73 \
 //y=0 //x2=12.21 //y2=0.625
cc_604 ( N_GND_c_58_p N_noxref_31_c_9441_n ) capacitor c=0.0140304f //x=12.78 \
 //y=0 //x2=12.21 //y2=0.625
cc_605 ( N_GND_c_4_p N_noxref_31_c_9441_n ) capacitor c=0.0404137f //x=12.95 \
 //y=0 //x2=12.21 //y2=0.625
cc_606 ( N_GND_M5_noxref_d N_noxref_31_M6_noxref_d ) capacitor c=0.00162435f \
 //x=9.025 //y=0.875 //x2=10 //y2=0.91
cc_607 ( N_GND_c_3_p N_noxref_31_M7_noxref_s ) capacitor c=8.16352e-19 \
 //x=8.14 //y=0 //x2=11.105 //y2=0.375
cc_608 ( N_GND_c_4_p N_noxref_31_M7_noxref_s ) capacitor c=0.00183576f \
 //x=12.95 //y=0 //x2=11.105 //y2=0.375
cc_609 ( N_GND_c_24_p N_noxref_32_c_9486_n ) capacitor c=0.00517234f //x=84.73 \
 //y=0 //x2=14.53 //y2=1.58
cc_610 ( N_GND_c_69_p N_noxref_32_c_9486_n ) capacitor c=0.00112872f \
 //x=14.045 //y=0 //x2=14.53 //y2=1.58
cc_611 ( N_GND_c_76_p N_noxref_32_c_9486_n ) capacitor c=0.0018229f //x=16.11 \
 //y=0 //x2=14.53 //y2=1.58
cc_612 ( N_GND_M8_noxref_d N_noxref_32_c_9486_n ) capacitor c=0.008625f \
 //x=13.94 //y=0.865 //x2=14.53 //y2=1.58
cc_613 ( N_GND_c_24_p N_noxref_32_c_9490_n ) capacitor c=0.00259029f //x=84.73 \
 //y=0 //x2=14.615 //y2=0.615
cc_614 ( N_GND_c_76_p N_noxref_32_c_9490_n ) capacitor c=0.0146901f //x=16.11 \
 //y=0 //x2=14.615 //y2=0.615
cc_615 ( N_GND_M8_noxref_d N_noxref_32_c_9490_n ) capacitor c=0.033812f \
 //x=13.94 //y=0.865 //x2=14.615 //y2=0.615
cc_616 ( N_GND_c_4_p N_noxref_32_c_9493_n ) capacitor c=2.91423e-19 //x=12.95 \
 //y=0 //x2=14.615 //y2=1.495
cc_617 ( N_GND_c_24_p N_noxref_32_c_9494_n ) capacitor c=0.0106919f //x=84.73 \
 //y=0 //x2=15.5 //y2=0.53
cc_618 ( N_GND_c_76_p N_noxref_32_c_9494_n ) capacitor c=0.0374253f //x=16.11 \
 //y=0 //x2=15.5 //y2=0.53
cc_619 ( N_GND_c_24_p N_noxref_32_c_9496_n ) capacitor c=0.00258845f //x=84.73 \
 //y=0 //x2=15.585 //y2=0.615
cc_620 ( N_GND_c_76_p N_noxref_32_c_9496_n ) capacitor c=0.0146256f //x=16.11 \
 //y=0 //x2=15.585 //y2=0.615
cc_621 ( N_GND_c_5_p N_noxref_32_c_9496_n ) capacitor c=0.0431718f //x=16.28 \
 //y=0 //x2=15.585 //y2=0.615
cc_622 ( N_GND_c_24_p N_noxref_32_M8_noxref_s ) capacitor c=0.00259029f \
 //x=84.73 //y=0 //x2=13.51 //y2=0.365
cc_623 ( N_GND_c_69_p N_noxref_32_M8_noxref_s ) capacitor c=0.0146901f \
 //x=14.045 //y=0 //x2=13.51 //y2=0.365
cc_624 ( N_GND_c_4_p N_noxref_32_M8_noxref_s ) capacitor c=0.0583534f \
 //x=12.95 //y=0 //x2=13.51 //y2=0.365
cc_625 ( N_GND_c_5_p N_noxref_32_M8_noxref_s ) capacitor c=0.00198043f \
 //x=16.28 //y=0 //x2=13.51 //y2=0.365
cc_626 ( N_GND_M8_noxref_d N_noxref_32_M8_noxref_s ) capacitor c=0.0334197f \
 //x=13.94 //y=0.865 //x2=13.51 //y2=0.365
cc_627 ( N_GND_c_24_p N_noxref_33_c_9537_n ) capacitor c=0.00517234f //x=84.73 \
 //y=0 //x2=17.86 //y2=1.58
cc_628 ( N_GND_c_84_p N_noxref_33_c_9537_n ) capacitor c=0.00112872f \
 //x=17.375 //y=0 //x2=17.86 //y2=1.58
cc_629 ( N_GND_c_91_p N_noxref_33_c_9537_n ) capacitor c=0.0018229f //x=19.44 \
 //y=0 //x2=17.86 //y2=1.58
cc_630 ( N_GND_M10_noxref_d N_noxref_33_c_9537_n ) capacitor c=0.008625f \
 //x=17.27 //y=0.865 //x2=17.86 //y2=1.58
cc_631 ( N_GND_c_24_p N_noxref_33_c_9541_n ) capacitor c=0.00259029f //x=84.73 \
 //y=0 //x2=17.945 //y2=0.615
cc_632 ( N_GND_c_91_p N_noxref_33_c_9541_n ) capacitor c=0.0146901f //x=19.44 \
 //y=0 //x2=17.945 //y2=0.615
cc_633 ( N_GND_M10_noxref_d N_noxref_33_c_9541_n ) capacitor c=0.033812f \
 //x=17.27 //y=0.865 //x2=17.945 //y2=0.615
cc_634 ( N_GND_c_5_p N_noxref_33_c_9544_n ) capacitor c=2.91423e-19 //x=16.28 \
 //y=0 //x2=17.945 //y2=1.495
cc_635 ( N_GND_c_24_p N_noxref_33_c_9545_n ) capacitor c=0.0106919f //x=84.73 \
 //y=0 //x2=18.83 //y2=0.53
cc_636 ( N_GND_c_91_p N_noxref_33_c_9545_n ) capacitor c=0.0374253f //x=19.44 \
 //y=0 //x2=18.83 //y2=0.53
cc_637 ( N_GND_c_24_p N_noxref_33_c_9547_n ) capacitor c=0.00258845f //x=84.73 \
 //y=0 //x2=18.915 //y2=0.615
cc_638 ( N_GND_c_91_p N_noxref_33_c_9547_n ) capacitor c=0.0146256f //x=19.44 \
 //y=0 //x2=18.915 //y2=0.615
cc_639 ( N_GND_c_6_p N_noxref_33_c_9547_n ) capacitor c=0.0431718f //x=19.61 \
 //y=0 //x2=18.915 //y2=0.615
cc_640 ( N_GND_c_24_p N_noxref_33_M10_noxref_s ) capacitor c=0.00259029f \
 //x=84.73 //y=0 //x2=16.84 //y2=0.365
cc_641 ( N_GND_c_84_p N_noxref_33_M10_noxref_s ) capacitor c=0.0146901f \
 //x=17.375 //y=0 //x2=16.84 //y2=0.365
cc_642 ( N_GND_c_5_p N_noxref_33_M10_noxref_s ) capacitor c=0.058339f \
 //x=16.28 //y=0 //x2=16.84 //y2=0.365
cc_643 ( N_GND_c_6_p N_noxref_33_M10_noxref_s ) capacitor c=0.00198098f \
 //x=19.61 //y=0 //x2=16.84 //y2=0.365
cc_644 ( N_GND_M10_noxref_d N_noxref_33_M10_noxref_s ) capacitor c=0.0334197f \
 //x=17.27 //y=0.865 //x2=16.84 //y2=0.365
cc_645 ( N_GND_c_24_p N_noxref_34_c_9588_n ) capacitor c=0.00517576f //x=84.73 \
 //y=0 //x2=21.085 //y2=1.59
cc_646 ( N_GND_c_98_p N_noxref_34_c_9588_n ) capacitor c=0.00111448f //x=20.6 \
 //y=0 //x2=21.085 //y2=1.59
cc_647 ( N_GND_c_105_p N_noxref_34_c_9588_n ) capacitor c=0.00180612f \
 //x=24.25 //y=0 //x2=21.085 //y2=1.59
cc_648 ( N_GND_M12_noxref_d N_noxref_34_c_9588_n ) capacitor c=0.00853078f \
 //x=20.495 //y=0.875 //x2=21.085 //y2=1.59
cc_649 ( N_GND_c_24_p N_noxref_34_c_9592_n ) capacitor c=0.00254475f //x=84.73 \
 //y=0 //x2=21.17 //y2=0.625
cc_650 ( N_GND_c_105_p N_noxref_34_c_9592_n ) capacitor c=0.0140928f //x=24.25 \
 //y=0 //x2=21.17 //y2=0.625
cc_651 ( N_GND_M12_noxref_d N_noxref_34_c_9592_n ) capacitor c=0.033954f \
 //x=20.495 //y=0.875 //x2=21.17 //y2=0.625
cc_652 ( N_GND_c_24_p N_noxref_34_c_9595_n ) capacitor c=0.0104386f //x=84.73 \
 //y=0 //x2=22.055 //y2=0.54
cc_653 ( N_GND_c_105_p N_noxref_34_c_9595_n ) capacitor c=0.0360726f //x=24.25 \
 //y=0 //x2=22.055 //y2=0.54
cc_654 ( N_GND_c_24_p N_noxref_34_M12_noxref_s ) capacitor c=0.00507657f \
 //x=84.73 //y=0 //x2=20.065 //y2=0.375
cc_655 ( N_GND_c_98_p N_noxref_34_M12_noxref_s ) capacitor c=0.0140928f \
 //x=20.6 //y=0 //x2=20.065 //y2=0.375
cc_656 ( N_GND_c_105_p N_noxref_34_M12_noxref_s ) capacitor c=0.0131437f \
 //x=24.25 //y=0 //x2=20.065 //y2=0.375
cc_657 ( N_GND_c_6_p N_noxref_34_M12_noxref_s ) capacitor c=0.0696963f \
 //x=19.61 //y=0 //x2=20.065 //y2=0.375
cc_658 ( N_GND_c_7_p N_noxref_34_M12_noxref_s ) capacitor c=3.31601e-19 \
 //x=24.42 //y=0 //x2=20.065 //y2=0.375
cc_659 ( N_GND_M12_noxref_d N_noxref_34_M12_noxref_s ) capacitor c=0.033718f \
 //x=20.495 //y=0.875 //x2=20.065 //y2=0.375
cc_660 ( N_GND_c_24_p N_noxref_35_c_9640_n ) capacitor c=0.00352952f //x=84.73 \
 //y=0 //x2=22.625 //y2=0.995
cc_661 ( N_GND_c_105_p N_noxref_35_c_9640_n ) capacitor c=0.00934524f \
 //x=24.25 //y=0 //x2=22.625 //y2=0.995
cc_662 ( N_GND_c_24_p N_noxref_35_c_9642_n ) capacitor c=0.00254475f //x=84.73 \
 //y=0 //x2=22.71 //y2=0.625
cc_663 ( N_GND_c_105_p N_noxref_35_c_9642_n ) capacitor c=0.0140928f //x=24.25 \
 //y=0 //x2=22.71 //y2=0.625
cc_664 ( N_GND_M12_noxref_d N_noxref_35_c_9642_n ) capacitor c=6.21394e-19 \
 //x=20.495 //y=0.875 //x2=22.71 //y2=0.625
cc_665 ( N_GND_c_24_p N_noxref_35_c_9645_n ) capacitor c=0.0105317f //x=84.73 \
 //y=0 //x2=23.595 //y2=0.54
cc_666 ( N_GND_c_105_p N_noxref_35_c_9645_n ) capacitor c=0.0364215f //x=24.25 \
 //y=0 //x2=23.595 //y2=0.54
cc_667 ( N_GND_c_24_p N_noxref_35_c_9647_n ) capacitor c=0.00254232f //x=84.73 \
 //y=0 //x2=23.68 //y2=0.625
cc_668 ( N_GND_c_105_p N_noxref_35_c_9647_n ) capacitor c=0.0140304f //x=24.25 \
 //y=0 //x2=23.68 //y2=0.625
cc_669 ( N_GND_c_7_p N_noxref_35_c_9647_n ) capacitor c=0.0404137f //x=24.42 \
 //y=0 //x2=23.68 //y2=0.625
cc_670 ( N_GND_M12_noxref_d N_noxref_35_M13_noxref_d ) capacitor c=0.00162435f \
 //x=20.495 //y=0.875 //x2=21.47 //y2=0.91
cc_671 ( N_GND_c_6_p N_noxref_35_M14_noxref_s ) capacitor c=8.16352e-19 \
 //x=19.61 //y=0 //x2=22.575 //y2=0.375
cc_672 ( N_GND_c_7_p N_noxref_35_M14_noxref_s ) capacitor c=0.00183576f \
 //x=24.42 //y=0 //x2=22.575 //y2=0.375
cc_673 ( N_GND_c_24_p N_noxref_36_c_9692_n ) capacitor c=0.00517234f //x=84.73 \
 //y=0 //x2=26 //y2=1.58
cc_674 ( N_GND_c_259_p N_noxref_36_c_9692_n ) capacitor c=0.00112872f \
 //x=25.515 //y=0 //x2=26 //y2=1.58
cc_675 ( N_GND_c_266_p N_noxref_36_c_9692_n ) capacitor c=0.0018229f //x=27.58 \
 //y=0 //x2=26 //y2=1.58
cc_676 ( N_GND_M15_noxref_d N_noxref_36_c_9692_n ) capacitor c=0.008625f \
 //x=25.41 //y=0.865 //x2=26 //y2=1.58
cc_677 ( N_GND_c_24_p N_noxref_36_c_9696_n ) capacitor c=0.00259029f //x=84.73 \
 //y=0 //x2=26.085 //y2=0.615
cc_678 ( N_GND_c_266_p N_noxref_36_c_9696_n ) capacitor c=0.0146901f //x=27.58 \
 //y=0 //x2=26.085 //y2=0.615
cc_679 ( N_GND_M15_noxref_d N_noxref_36_c_9696_n ) capacitor c=0.033812f \
 //x=25.41 //y=0.865 //x2=26.085 //y2=0.615
cc_680 ( N_GND_c_7_p N_noxref_36_c_9699_n ) capacitor c=2.91423e-19 //x=24.42 \
 //y=0 //x2=26.085 //y2=1.495
cc_681 ( N_GND_c_24_p N_noxref_36_c_9700_n ) capacitor c=0.0106919f //x=84.73 \
 //y=0 //x2=26.97 //y2=0.53
cc_682 ( N_GND_c_266_p N_noxref_36_c_9700_n ) capacitor c=0.0374253f //x=27.58 \
 //y=0 //x2=26.97 //y2=0.53
cc_683 ( N_GND_c_24_p N_noxref_36_c_9702_n ) capacitor c=0.00258845f //x=84.73 \
 //y=0 //x2=27.055 //y2=0.615
cc_684 ( N_GND_c_266_p N_noxref_36_c_9702_n ) capacitor c=0.0146256f //x=27.58 \
 //y=0 //x2=27.055 //y2=0.615
cc_685 ( N_GND_c_8_p N_noxref_36_c_9702_n ) capacitor c=0.0431718f //x=27.75 \
 //y=0 //x2=27.055 //y2=0.615
cc_686 ( N_GND_c_24_p N_noxref_36_M15_noxref_s ) capacitor c=0.00259029f \
 //x=84.73 //y=0 //x2=24.98 //y2=0.365
cc_687 ( N_GND_c_259_p N_noxref_36_M15_noxref_s ) capacitor c=0.0146901f \
 //x=25.515 //y=0 //x2=24.98 //y2=0.365
cc_688 ( N_GND_c_7_p N_noxref_36_M15_noxref_s ) capacitor c=0.0583534f \
 //x=24.42 //y=0 //x2=24.98 //y2=0.365
cc_689 ( N_GND_c_8_p N_noxref_36_M15_noxref_s ) capacitor c=0.00198098f \
 //x=27.75 //y=0 //x2=24.98 //y2=0.365
cc_690 ( N_GND_M15_noxref_d N_noxref_36_M15_noxref_s ) capacitor c=0.0334197f \
 //x=25.41 //y=0.865 //x2=24.98 //y2=0.365
cc_691 ( N_GND_c_24_p N_noxref_37_c_9743_n ) capacitor c=0.00517576f //x=84.73 \
 //y=0 //x2=29.225 //y2=1.59
cc_692 ( N_GND_c_128_p N_noxref_37_c_9743_n ) capacitor c=0.00111448f \
 //x=28.74 //y=0 //x2=29.225 //y2=1.59
cc_693 ( N_GND_c_135_p N_noxref_37_c_9743_n ) capacitor c=0.00180612f \
 //x=32.39 //y=0 //x2=29.225 //y2=1.59
cc_694 ( N_GND_M17_noxref_d N_noxref_37_c_9743_n ) capacitor c=0.00853078f \
 //x=28.635 //y=0.875 //x2=29.225 //y2=1.59
cc_695 ( N_GND_c_24_p N_noxref_37_c_9747_n ) capacitor c=0.00254475f //x=84.73 \
 //y=0 //x2=29.31 //y2=0.625
cc_696 ( N_GND_c_135_p N_noxref_37_c_9747_n ) capacitor c=0.0140928f //x=32.39 \
 //y=0 //x2=29.31 //y2=0.625
cc_697 ( N_GND_M17_noxref_d N_noxref_37_c_9747_n ) capacitor c=0.033954f \
 //x=28.635 //y=0.875 //x2=29.31 //y2=0.625
cc_698 ( N_GND_c_24_p N_noxref_37_c_9750_n ) capacitor c=0.0104506f //x=84.73 \
 //y=0 //x2=30.195 //y2=0.54
cc_699 ( N_GND_c_135_p N_noxref_37_c_9750_n ) capacitor c=0.0360726f //x=32.39 \
 //y=0 //x2=30.195 //y2=0.54
cc_700 ( N_GND_c_24_p N_noxref_37_M17_noxref_s ) capacitor c=0.00507657f \
 //x=84.73 //y=0 //x2=28.205 //y2=0.375
cc_701 ( N_GND_c_128_p N_noxref_37_M17_noxref_s ) capacitor c=0.0140928f \
 //x=28.74 //y=0 //x2=28.205 //y2=0.375
cc_702 ( N_GND_c_135_p N_noxref_37_M17_noxref_s ) capacitor c=0.0131437f \
 //x=32.39 //y=0 //x2=28.205 //y2=0.375
cc_703 ( N_GND_c_8_p N_noxref_37_M17_noxref_s ) capacitor c=0.0696963f \
 //x=27.75 //y=0 //x2=28.205 //y2=0.375
cc_704 ( N_GND_c_9_p N_noxref_37_M17_noxref_s ) capacitor c=3.31601e-19 \
 //x=32.56 //y=0 //x2=28.205 //y2=0.375
cc_705 ( N_GND_M17_noxref_d N_noxref_37_M17_noxref_s ) capacitor c=0.033718f \
 //x=28.635 //y=0.875 //x2=28.205 //y2=0.375
cc_706 ( N_GND_c_24_p N_noxref_38_c_9792_n ) capacitor c=0.00352952f //x=84.73 \
 //y=0 //x2=30.765 //y2=0.995
cc_707 ( N_GND_c_135_p N_noxref_38_c_9792_n ) capacitor c=0.00934524f \
 //x=32.39 //y=0 //x2=30.765 //y2=0.995
cc_708 ( N_GND_c_24_p N_noxref_38_c_9794_n ) capacitor c=0.00254475f //x=84.73 \
 //y=0 //x2=30.85 //y2=0.625
cc_709 ( N_GND_c_135_p N_noxref_38_c_9794_n ) capacitor c=0.0140928f //x=32.39 \
 //y=0 //x2=30.85 //y2=0.625
cc_710 ( N_GND_M17_noxref_d N_noxref_38_c_9794_n ) capacitor c=6.21394e-19 \
 //x=28.635 //y=0.875 //x2=30.85 //y2=0.625
cc_711 ( N_GND_c_24_p N_noxref_38_c_9797_n ) capacitor c=0.010529f //x=84.73 \
 //y=0 //x2=31.735 //y2=0.54
cc_712 ( N_GND_c_135_p N_noxref_38_c_9797_n ) capacitor c=0.0364674f //x=32.39 \
 //y=0 //x2=31.735 //y2=0.54
cc_713 ( N_GND_c_24_p N_noxref_38_c_9799_n ) capacitor c=0.00254232f //x=84.73 \
 //y=0 //x2=31.82 //y2=0.625
cc_714 ( N_GND_c_135_p N_noxref_38_c_9799_n ) capacitor c=0.0140304f //x=32.39 \
 //y=0 //x2=31.82 //y2=0.625
cc_715 ( N_GND_c_9_p N_noxref_38_c_9799_n ) capacitor c=0.0404137f //x=32.56 \
 //y=0 //x2=31.82 //y2=0.625
cc_716 ( N_GND_M17_noxref_d N_noxref_38_M18_noxref_d ) capacitor c=0.00162435f \
 //x=28.635 //y=0.875 //x2=29.61 //y2=0.91
cc_717 ( N_GND_c_8_p N_noxref_38_M19_noxref_s ) capacitor c=8.16352e-19 \
 //x=27.75 //y=0 //x2=30.715 //y2=0.375
cc_718 ( N_GND_c_9_p N_noxref_38_M19_noxref_s ) capacitor c=0.00180469f \
 //x=32.56 //y=0 //x2=30.715 //y2=0.375
cc_719 ( N_GND_c_24_p N_noxref_39_c_9844_n ) capacitor c=0.00517576f //x=84.73 \
 //y=0 //x2=34.035 //y2=1.59
cc_720 ( N_GND_c_138_p N_noxref_39_c_9844_n ) capacitor c=0.00111448f \
 //x=33.55 //y=0 //x2=34.035 //y2=1.59
cc_721 ( N_GND_c_145_p N_noxref_39_c_9844_n ) capacitor c=0.00180612f //x=37.2 \
 //y=0 //x2=34.035 //y2=1.59
cc_722 ( N_GND_M20_noxref_d N_noxref_39_c_9844_n ) capacitor c=0.00853078f \
 //x=33.445 //y=0.875 //x2=34.035 //y2=1.59
cc_723 ( N_GND_c_24_p N_noxref_39_c_9848_n ) capacitor c=0.00254475f //x=84.73 \
 //y=0 //x2=34.12 //y2=0.625
cc_724 ( N_GND_c_145_p N_noxref_39_c_9848_n ) capacitor c=0.0140928f //x=37.2 \
 //y=0 //x2=34.12 //y2=0.625
cc_725 ( N_GND_M20_noxref_d N_noxref_39_c_9848_n ) capacitor c=0.033954f \
 //x=33.445 //y=0.875 //x2=34.12 //y2=0.625
cc_726 ( N_GND_c_24_p N_noxref_39_c_9851_n ) capacitor c=0.0104386f //x=84.73 \
 //y=0 //x2=35.005 //y2=0.54
cc_727 ( N_GND_c_145_p N_noxref_39_c_9851_n ) capacitor c=0.0360726f //x=37.2 \
 //y=0 //x2=35.005 //y2=0.54
cc_728 ( N_GND_c_24_p N_noxref_39_M20_noxref_s ) capacitor c=0.00507657f \
 //x=84.73 //y=0 //x2=33.015 //y2=0.375
cc_729 ( N_GND_c_138_p N_noxref_39_M20_noxref_s ) capacitor c=0.0140928f \
 //x=33.55 //y=0 //x2=33.015 //y2=0.375
cc_730 ( N_GND_c_145_p N_noxref_39_M20_noxref_s ) capacitor c=0.0131437f \
 //x=37.2 //y=0 //x2=33.015 //y2=0.375
cc_731 ( N_GND_c_9_p N_noxref_39_M20_noxref_s ) capacitor c=0.0696963f \
 //x=32.56 //y=0 //x2=33.015 //y2=0.375
cc_732 ( N_GND_c_10_p N_noxref_39_M20_noxref_s ) capacitor c=3.31601e-19 \
 //x=37.37 //y=0 //x2=33.015 //y2=0.375
cc_733 ( N_GND_M20_noxref_d N_noxref_39_M20_noxref_s ) capacitor c=0.033718f \
 //x=33.445 //y=0.875 //x2=33.015 //y2=0.375
cc_734 ( N_GND_c_24_p N_noxref_40_c_9896_n ) capacitor c=0.00352952f //x=84.73 \
 //y=0 //x2=35.575 //y2=0.995
cc_735 ( N_GND_c_145_p N_noxref_40_c_9896_n ) capacitor c=0.00934524f //x=37.2 \
 //y=0 //x2=35.575 //y2=0.995
cc_736 ( N_GND_c_24_p N_noxref_40_c_9898_n ) capacitor c=0.00254475f //x=84.73 \
 //y=0 //x2=35.66 //y2=0.625
cc_737 ( N_GND_c_145_p N_noxref_40_c_9898_n ) capacitor c=0.0140928f //x=37.2 \
 //y=0 //x2=35.66 //y2=0.625
cc_738 ( N_GND_M20_noxref_d N_noxref_40_c_9898_n ) capacitor c=6.21394e-19 \
 //x=33.445 //y=0.875 //x2=35.66 //y2=0.625
cc_739 ( N_GND_c_24_p N_noxref_40_c_9901_n ) capacitor c=0.0105317f //x=84.73 \
 //y=0 //x2=36.545 //y2=0.54
cc_740 ( N_GND_c_145_p N_noxref_40_c_9901_n ) capacitor c=0.0364215f //x=37.2 \
 //y=0 //x2=36.545 //y2=0.54
cc_741 ( N_GND_c_24_p N_noxref_40_c_9903_n ) capacitor c=0.00254232f //x=84.73 \
 //y=0 //x2=36.63 //y2=0.625
cc_742 ( N_GND_c_145_p N_noxref_40_c_9903_n ) capacitor c=0.0140304f //x=37.2 \
 //y=0 //x2=36.63 //y2=0.625
cc_743 ( N_GND_c_10_p N_noxref_40_c_9903_n ) capacitor c=0.0404137f //x=37.37 \
 //y=0 //x2=36.63 //y2=0.625
cc_744 ( N_GND_M20_noxref_d N_noxref_40_M21_noxref_d ) capacitor c=0.00162435f \
 //x=33.445 //y=0.875 //x2=34.42 //y2=0.91
cc_745 ( N_GND_c_9_p N_noxref_40_M22_noxref_s ) capacitor c=8.16352e-19 \
 //x=32.56 //y=0 //x2=35.525 //y2=0.375
cc_746 ( N_GND_c_10_p N_noxref_40_M22_noxref_s ) capacitor c=0.00183576f \
 //x=37.37 //y=0 //x2=35.525 //y2=0.375
cc_747 ( N_GND_c_24_p N_noxref_41_c_9948_n ) capacitor c=0.00517234f //x=84.73 \
 //y=0 //x2=38.95 //y2=1.58
cc_748 ( N_GND_c_156_p N_noxref_41_c_9948_n ) capacitor c=0.00112872f \
 //x=38.465 //y=0 //x2=38.95 //y2=1.58
cc_749 ( N_GND_c_163_p N_noxref_41_c_9948_n ) capacitor c=0.0018229f //x=40.53 \
 //y=0 //x2=38.95 //y2=1.58
cc_750 ( N_GND_M23_noxref_d N_noxref_41_c_9948_n ) capacitor c=0.008625f \
 //x=38.36 //y=0.865 //x2=38.95 //y2=1.58
cc_751 ( N_GND_c_24_p N_noxref_41_c_9952_n ) capacitor c=0.00259029f //x=84.73 \
 //y=0 //x2=39.035 //y2=0.615
cc_752 ( N_GND_c_163_p N_noxref_41_c_9952_n ) capacitor c=0.0146901f //x=40.53 \
 //y=0 //x2=39.035 //y2=0.615
cc_753 ( N_GND_M23_noxref_d N_noxref_41_c_9952_n ) capacitor c=0.033812f \
 //x=38.36 //y=0.865 //x2=39.035 //y2=0.615
cc_754 ( N_GND_c_10_p N_noxref_41_c_9955_n ) capacitor c=2.91423e-19 //x=37.37 \
 //y=0 //x2=39.035 //y2=1.495
cc_755 ( N_GND_c_24_p N_noxref_41_c_9956_n ) capacitor c=0.0106919f //x=84.73 \
 //y=0 //x2=39.92 //y2=0.53
cc_756 ( N_GND_c_163_p N_noxref_41_c_9956_n ) capacitor c=0.0374253f //x=40.53 \
 //y=0 //x2=39.92 //y2=0.53
cc_757 ( N_GND_c_24_p N_noxref_41_c_9958_n ) capacitor c=0.00258845f //x=84.73 \
 //y=0 //x2=40.005 //y2=0.615
cc_758 ( N_GND_c_163_p N_noxref_41_c_9958_n ) capacitor c=0.0146256f //x=40.53 \
 //y=0 //x2=40.005 //y2=0.615
cc_759 ( N_GND_c_11_p N_noxref_41_c_9958_n ) capacitor c=0.0431718f //x=40.7 \
 //y=0 //x2=40.005 //y2=0.615
cc_760 ( N_GND_c_24_p N_noxref_41_M23_noxref_s ) capacitor c=0.00259029f \
 //x=84.73 //y=0 //x2=37.93 //y2=0.365
cc_761 ( N_GND_c_156_p N_noxref_41_M23_noxref_s ) capacitor c=0.0146901f \
 //x=38.465 //y=0 //x2=37.93 //y2=0.365
cc_762 ( N_GND_c_10_p N_noxref_41_M23_noxref_s ) capacitor c=0.0583534f \
 //x=37.37 //y=0 //x2=37.93 //y2=0.365
cc_763 ( N_GND_c_11_p N_noxref_41_M23_noxref_s ) capacitor c=0.00198043f \
 //x=40.7 //y=0 //x2=37.93 //y2=0.365
cc_764 ( N_GND_M23_noxref_d N_noxref_41_M23_noxref_s ) capacitor c=0.0334197f \
 //x=38.36 //y=0.865 //x2=37.93 //y2=0.365
cc_765 ( N_GND_c_24_p N_noxref_42_c_9999_n ) capacitor c=0.00517234f //x=84.73 \
 //y=0 //x2=42.28 //y2=1.58
cc_766 ( N_GND_c_171_p N_noxref_42_c_9999_n ) capacitor c=0.00112872f \
 //x=41.795 //y=0 //x2=42.28 //y2=1.58
cc_767 ( N_GND_c_178_p N_noxref_42_c_9999_n ) capacitor c=0.0018229f //x=43.86 \
 //y=0 //x2=42.28 //y2=1.58
cc_768 ( N_GND_M25_noxref_d N_noxref_42_c_9999_n ) capacitor c=0.008625f \
 //x=41.69 //y=0.865 //x2=42.28 //y2=1.58
cc_769 ( N_GND_c_24_p N_noxref_42_c_10003_n ) capacitor c=0.00259029f \
 //x=84.73 //y=0 //x2=42.365 //y2=0.615
cc_770 ( N_GND_c_178_p N_noxref_42_c_10003_n ) capacitor c=0.0146901f \
 //x=43.86 //y=0 //x2=42.365 //y2=0.615
cc_771 ( N_GND_M25_noxref_d N_noxref_42_c_10003_n ) capacitor c=0.033812f \
 //x=41.69 //y=0.865 //x2=42.365 //y2=0.615
cc_772 ( N_GND_c_11_p N_noxref_42_c_10006_n ) capacitor c=2.91423e-19 //x=40.7 \
 //y=0 //x2=42.365 //y2=1.495
cc_773 ( N_GND_c_24_p N_noxref_42_c_10007_n ) capacitor c=0.0106919f //x=84.73 \
 //y=0 //x2=43.25 //y2=0.53
cc_774 ( N_GND_c_178_p N_noxref_42_c_10007_n ) capacitor c=0.0374253f \
 //x=43.86 //y=0 //x2=43.25 //y2=0.53
cc_775 ( N_GND_c_24_p N_noxref_42_c_10009_n ) capacitor c=0.00258845f \
 //x=84.73 //y=0 //x2=43.335 //y2=0.615
cc_776 ( N_GND_c_178_p N_noxref_42_c_10009_n ) capacitor c=0.0146256f \
 //x=43.86 //y=0 //x2=43.335 //y2=0.615
cc_777 ( N_GND_c_12_p N_noxref_42_c_10009_n ) capacitor c=0.0431718f //x=44.03 \
 //y=0 //x2=43.335 //y2=0.615
cc_778 ( N_GND_c_24_p N_noxref_42_M25_noxref_s ) capacitor c=0.00259029f \
 //x=84.73 //y=0 //x2=41.26 //y2=0.365
cc_779 ( N_GND_c_171_p N_noxref_42_M25_noxref_s ) capacitor c=0.0146901f \
 //x=41.795 //y=0 //x2=41.26 //y2=0.365
cc_780 ( N_GND_c_11_p N_noxref_42_M25_noxref_s ) capacitor c=0.058339f \
 //x=40.7 //y=0 //x2=41.26 //y2=0.365
cc_781 ( N_GND_c_12_p N_noxref_42_M25_noxref_s ) capacitor c=0.00198098f \
 //x=44.03 //y=0 //x2=41.26 //y2=0.365
cc_782 ( N_GND_M25_noxref_d N_noxref_42_M25_noxref_s ) capacitor c=0.0334197f \
 //x=41.69 //y=0.865 //x2=41.26 //y2=0.365
cc_783 ( N_GND_c_24_p N_noxref_43_c_10050_n ) capacitor c=0.00517576f \
 //x=84.73 //y=0 //x2=45.505 //y2=1.59
cc_784 ( N_GND_c_188_p N_noxref_43_c_10050_n ) capacitor c=0.00111448f \
 //x=45.02 //y=0 //x2=45.505 //y2=1.59
cc_785 ( N_GND_c_195_p N_noxref_43_c_10050_n ) capacitor c=0.00180612f \
 //x=48.67 //y=0 //x2=45.505 //y2=1.59
cc_786 ( N_GND_M27_noxref_d N_noxref_43_c_10050_n ) capacitor c=0.00853078f \
 //x=44.915 //y=0.875 //x2=45.505 //y2=1.59
cc_787 ( N_GND_c_24_p N_noxref_43_c_10054_n ) capacitor c=0.00254475f \
 //x=84.73 //y=0 //x2=45.59 //y2=0.625
cc_788 ( N_GND_c_195_p N_noxref_43_c_10054_n ) capacitor c=0.0140928f \
 //x=48.67 //y=0 //x2=45.59 //y2=0.625
cc_789 ( N_GND_M27_noxref_d N_noxref_43_c_10054_n ) capacitor c=0.033954f \
 //x=44.915 //y=0.875 //x2=45.59 //y2=0.625
cc_790 ( N_GND_c_24_p N_noxref_43_c_10057_n ) capacitor c=0.0104386f //x=84.73 \
 //y=0 //x2=46.475 //y2=0.54
cc_791 ( N_GND_c_195_p N_noxref_43_c_10057_n ) capacitor c=0.0360726f \
 //x=48.67 //y=0 //x2=46.475 //y2=0.54
cc_792 ( N_GND_c_24_p N_noxref_43_M27_noxref_s ) capacitor c=0.00507657f \
 //x=84.73 //y=0 //x2=44.485 //y2=0.375
cc_793 ( N_GND_c_188_p N_noxref_43_M27_noxref_s ) capacitor c=0.0140928f \
 //x=45.02 //y=0 //x2=44.485 //y2=0.375
cc_794 ( N_GND_c_195_p N_noxref_43_M27_noxref_s ) capacitor c=0.0131437f \
 //x=48.67 //y=0 //x2=44.485 //y2=0.375
cc_795 ( N_GND_c_12_p N_noxref_43_M27_noxref_s ) capacitor c=0.0696963f \
 //x=44.03 //y=0 //x2=44.485 //y2=0.375
cc_796 ( N_GND_c_13_p N_noxref_43_M27_noxref_s ) capacitor c=3.31601e-19 \
 //x=48.84 //y=0 //x2=44.485 //y2=0.375
cc_797 ( N_GND_M27_noxref_d N_noxref_43_M27_noxref_s ) capacitor c=0.033718f \
 //x=44.915 //y=0.875 //x2=44.485 //y2=0.375
cc_798 ( N_GND_c_24_p N_noxref_44_c_10102_n ) capacitor c=0.00352952f \
 //x=84.73 //y=0 //x2=47.045 //y2=0.995
cc_799 ( N_GND_c_195_p N_noxref_44_c_10102_n ) capacitor c=0.00934524f \
 //x=48.67 //y=0 //x2=47.045 //y2=0.995
cc_800 ( N_GND_c_24_p N_noxref_44_c_10104_n ) capacitor c=0.00254475f \
 //x=84.73 //y=0 //x2=47.13 //y2=0.625
cc_801 ( N_GND_c_195_p N_noxref_44_c_10104_n ) capacitor c=0.0140928f \
 //x=48.67 //y=0 //x2=47.13 //y2=0.625
cc_802 ( N_GND_M27_noxref_d N_noxref_44_c_10104_n ) capacitor c=6.21394e-19 \
 //x=44.915 //y=0.875 //x2=47.13 //y2=0.625
cc_803 ( N_GND_c_24_p N_noxref_44_c_10107_n ) capacitor c=0.0105317f //x=84.73 \
 //y=0 //x2=48.015 //y2=0.54
cc_804 ( N_GND_c_195_p N_noxref_44_c_10107_n ) capacitor c=0.0364215f \
 //x=48.67 //y=0 //x2=48.015 //y2=0.54
cc_805 ( N_GND_c_24_p N_noxref_44_c_10109_n ) capacitor c=0.00254232f \
 //x=84.73 //y=0 //x2=48.1 //y2=0.625
cc_806 ( N_GND_c_195_p N_noxref_44_c_10109_n ) capacitor c=0.0140304f \
 //x=48.67 //y=0 //x2=48.1 //y2=0.625
cc_807 ( N_GND_c_13_p N_noxref_44_c_10109_n ) capacitor c=0.0404137f //x=48.84 \
 //y=0 //x2=48.1 //y2=0.625
cc_808 ( N_GND_M27_noxref_d N_noxref_44_M28_noxref_d ) capacitor c=0.00162435f \
 //x=44.915 //y=0.875 //x2=45.89 //y2=0.91
cc_809 ( N_GND_c_12_p N_noxref_44_M29_noxref_s ) capacitor c=8.16352e-19 \
 //x=44.03 //y=0 //x2=46.995 //y2=0.375
cc_810 ( N_GND_c_13_p N_noxref_44_M29_noxref_s ) capacitor c=0.00183576f \
 //x=48.84 //y=0 //x2=46.995 //y2=0.375
cc_811 ( N_GND_c_24_p N_noxref_45_c_10154_n ) capacitor c=0.00517234f \
 //x=84.73 //y=0 //x2=50.42 //y2=1.58
cc_812 ( N_GND_c_269_p N_noxref_45_c_10154_n ) capacitor c=0.00112872f \
 //x=49.935 //y=0 //x2=50.42 //y2=1.58
cc_813 ( N_GND_c_276_p N_noxref_45_c_10154_n ) capacitor c=0.0018229f //x=52 \
 //y=0 //x2=50.42 //y2=1.58
cc_814 ( N_GND_M30_noxref_d N_noxref_45_c_10154_n ) capacitor c=0.008625f \
 //x=49.83 //y=0.865 //x2=50.42 //y2=1.58
cc_815 ( N_GND_c_24_p N_noxref_45_c_10158_n ) capacitor c=0.00259029f \
 //x=84.73 //y=0 //x2=50.505 //y2=0.615
cc_816 ( N_GND_c_276_p N_noxref_45_c_10158_n ) capacitor c=0.0146901f //x=52 \
 //y=0 //x2=50.505 //y2=0.615
cc_817 ( N_GND_M30_noxref_d N_noxref_45_c_10158_n ) capacitor c=0.033812f \
 //x=49.83 //y=0.865 //x2=50.505 //y2=0.615
cc_818 ( N_GND_c_13_p N_noxref_45_c_10161_n ) capacitor c=2.91423e-19 \
 //x=48.84 //y=0 //x2=50.505 //y2=1.495
cc_819 ( N_GND_c_24_p N_noxref_45_c_10162_n ) capacitor c=0.0106919f //x=84.73 \
 //y=0 //x2=51.39 //y2=0.53
cc_820 ( N_GND_c_276_p N_noxref_45_c_10162_n ) capacitor c=0.0374253f //x=52 \
 //y=0 //x2=51.39 //y2=0.53
cc_821 ( N_GND_c_24_p N_noxref_45_c_10164_n ) capacitor c=0.00258845f \
 //x=84.73 //y=0 //x2=51.475 //y2=0.615
cc_822 ( N_GND_c_276_p N_noxref_45_c_10164_n ) capacitor c=0.0146256f //x=52 \
 //y=0 //x2=51.475 //y2=0.615
cc_823 ( N_GND_c_14_p N_noxref_45_c_10164_n ) capacitor c=0.0431718f //x=52.17 \
 //y=0 //x2=51.475 //y2=0.615
cc_824 ( N_GND_c_24_p N_noxref_45_M30_noxref_s ) capacitor c=0.00259029f \
 //x=84.73 //y=0 //x2=49.4 //y2=0.365
cc_825 ( N_GND_c_269_p N_noxref_45_M30_noxref_s ) capacitor c=0.0146901f \
 //x=49.935 //y=0 //x2=49.4 //y2=0.365
cc_826 ( N_GND_c_13_p N_noxref_45_M30_noxref_s ) capacitor c=0.0583534f \
 //x=48.84 //y=0 //x2=49.4 //y2=0.365
cc_827 ( N_GND_c_14_p N_noxref_45_M30_noxref_s ) capacitor c=0.00198098f \
 //x=52.17 //y=0 //x2=49.4 //y2=0.365
cc_828 ( N_GND_M30_noxref_d N_noxref_45_M30_noxref_s ) capacitor c=0.0334197f \
 //x=49.83 //y=0.865 //x2=49.4 //y2=0.365
cc_829 ( N_GND_c_24_p N_noxref_46_c_10205_n ) capacitor c=0.00517576f \
 //x=84.73 //y=0 //x2=53.645 //y2=1.59
cc_830 ( N_GND_c_288_p N_noxref_46_c_10205_n ) capacitor c=0.00111448f \
 //x=53.16 //y=0 //x2=53.645 //y2=1.59
cc_831 ( N_GND_c_295_p N_noxref_46_c_10205_n ) capacitor c=0.00180612f \
 //x=56.81 //y=0 //x2=53.645 //y2=1.59
cc_832 ( N_GND_M32_noxref_d N_noxref_46_c_10205_n ) capacitor c=0.00853078f \
 //x=53.055 //y=0.875 //x2=53.645 //y2=1.59
cc_833 ( N_GND_c_24_p N_noxref_46_c_10209_n ) capacitor c=0.00254475f \
 //x=84.73 //y=0 //x2=53.73 //y2=0.625
cc_834 ( N_GND_c_295_p N_noxref_46_c_10209_n ) capacitor c=0.0140928f \
 //x=56.81 //y=0 //x2=53.73 //y2=0.625
cc_835 ( N_GND_M32_noxref_d N_noxref_46_c_10209_n ) capacitor c=0.033954f \
 //x=53.055 //y=0.875 //x2=53.73 //y2=0.625
cc_836 ( N_GND_c_24_p N_noxref_46_c_10212_n ) capacitor c=0.0104506f //x=84.73 \
 //y=0 //x2=54.615 //y2=0.54
cc_837 ( N_GND_c_295_p N_noxref_46_c_10212_n ) capacitor c=0.0360726f \
 //x=56.81 //y=0 //x2=54.615 //y2=0.54
cc_838 ( N_GND_c_24_p N_noxref_46_M32_noxref_s ) capacitor c=0.00507657f \
 //x=84.73 //y=0 //x2=52.625 //y2=0.375
cc_839 ( N_GND_c_288_p N_noxref_46_M32_noxref_s ) capacitor c=0.0140928f \
 //x=53.16 //y=0 //x2=52.625 //y2=0.375
cc_840 ( N_GND_c_295_p N_noxref_46_M32_noxref_s ) capacitor c=0.0131437f \
 //x=56.81 //y=0 //x2=52.625 //y2=0.375
cc_841 ( N_GND_c_14_p N_noxref_46_M32_noxref_s ) capacitor c=0.0696963f \
 //x=52.17 //y=0 //x2=52.625 //y2=0.375
cc_842 ( N_GND_c_15_p N_noxref_46_M32_noxref_s ) capacitor c=3.31601e-19 \
 //x=56.98 //y=0 //x2=52.625 //y2=0.375
cc_843 ( N_GND_M32_noxref_d N_noxref_46_M32_noxref_s ) capacitor c=0.033718f \
 //x=53.055 //y=0.875 //x2=52.625 //y2=0.375
cc_844 ( N_GND_c_24_p N_noxref_47_c_10254_n ) capacitor c=0.00352952f \
 //x=84.73 //y=0 //x2=55.185 //y2=0.995
cc_845 ( N_GND_c_295_p N_noxref_47_c_10254_n ) capacitor c=0.00934524f \
 //x=56.81 //y=0 //x2=55.185 //y2=0.995
cc_846 ( N_GND_c_24_p N_noxref_47_c_10256_n ) capacitor c=0.00254475f \
 //x=84.73 //y=0 //x2=55.27 //y2=0.625
cc_847 ( N_GND_c_295_p N_noxref_47_c_10256_n ) capacitor c=0.0140928f \
 //x=56.81 //y=0 //x2=55.27 //y2=0.625
cc_848 ( N_GND_M32_noxref_d N_noxref_47_c_10256_n ) capacitor c=6.21394e-19 \
 //x=53.055 //y=0.875 //x2=55.27 //y2=0.625
cc_849 ( N_GND_c_24_p N_noxref_47_c_10259_n ) capacitor c=0.010529f //x=84.73 \
 //y=0 //x2=56.155 //y2=0.54
cc_850 ( N_GND_c_295_p N_noxref_47_c_10259_n ) capacitor c=0.0364674f \
 //x=56.81 //y=0 //x2=56.155 //y2=0.54
cc_851 ( N_GND_c_24_p N_noxref_47_c_10261_n ) capacitor c=0.00254232f \
 //x=84.73 //y=0 //x2=56.24 //y2=0.625
cc_852 ( N_GND_c_295_p N_noxref_47_c_10261_n ) capacitor c=0.0140304f \
 //x=56.81 //y=0 //x2=56.24 //y2=0.625
cc_853 ( N_GND_c_15_p N_noxref_47_c_10261_n ) capacitor c=0.0404137f //x=56.98 \
 //y=0 //x2=56.24 //y2=0.625
cc_854 ( N_GND_M32_noxref_d N_noxref_47_M33_noxref_d ) capacitor c=0.00162435f \
 //x=53.055 //y=0.875 //x2=54.03 //y2=0.91
cc_855 ( N_GND_c_14_p N_noxref_47_M34_noxref_s ) capacitor c=8.16352e-19 \
 //x=52.17 //y=0 //x2=55.135 //y2=0.375
cc_856 ( N_GND_c_15_p N_noxref_47_M34_noxref_s ) capacitor c=0.00180469f \
 //x=56.98 //y=0 //x2=55.135 //y2=0.375
cc_857 ( N_GND_c_24_p N_noxref_48_c_10306_n ) capacitor c=0.00517576f \
 //x=84.73 //y=0 //x2=58.455 //y2=1.59
cc_858 ( N_GND_c_298_p N_noxref_48_c_10306_n ) capacitor c=0.00111448f \
 //x=57.97 //y=0 //x2=58.455 //y2=1.59
cc_859 ( N_GND_c_305_p N_noxref_48_c_10306_n ) capacitor c=0.00180612f \
 //x=61.62 //y=0 //x2=58.455 //y2=1.59
cc_860 ( N_GND_M35_noxref_d N_noxref_48_c_10306_n ) capacitor c=0.00853078f \
 //x=57.865 //y=0.875 //x2=58.455 //y2=1.59
cc_861 ( N_GND_c_24_p N_noxref_48_c_10310_n ) capacitor c=0.00254475f \
 //x=84.73 //y=0 //x2=58.54 //y2=0.625
cc_862 ( N_GND_c_305_p N_noxref_48_c_10310_n ) capacitor c=0.0140928f \
 //x=61.62 //y=0 //x2=58.54 //y2=0.625
cc_863 ( N_GND_M35_noxref_d N_noxref_48_c_10310_n ) capacitor c=0.033954f \
 //x=57.865 //y=0.875 //x2=58.54 //y2=0.625
cc_864 ( N_GND_c_24_p N_noxref_48_c_10313_n ) capacitor c=0.0104386f //x=84.73 \
 //y=0 //x2=59.425 //y2=0.54
cc_865 ( N_GND_c_305_p N_noxref_48_c_10313_n ) capacitor c=0.0360726f \
 //x=61.62 //y=0 //x2=59.425 //y2=0.54
cc_866 ( N_GND_c_24_p N_noxref_48_M35_noxref_s ) capacitor c=0.00507657f \
 //x=84.73 //y=0 //x2=57.435 //y2=0.375
cc_867 ( N_GND_c_298_p N_noxref_48_M35_noxref_s ) capacitor c=0.0140928f \
 //x=57.97 //y=0 //x2=57.435 //y2=0.375
cc_868 ( N_GND_c_305_p N_noxref_48_M35_noxref_s ) capacitor c=0.0131437f \
 //x=61.62 //y=0 //x2=57.435 //y2=0.375
cc_869 ( N_GND_c_15_p N_noxref_48_M35_noxref_s ) capacitor c=0.0696963f \
 //x=56.98 //y=0 //x2=57.435 //y2=0.375
cc_870 ( N_GND_c_16_p N_noxref_48_M35_noxref_s ) capacitor c=3.31601e-19 \
 //x=61.79 //y=0 //x2=57.435 //y2=0.375
cc_871 ( N_GND_M35_noxref_d N_noxref_48_M35_noxref_s ) capacitor c=0.033718f \
 //x=57.865 //y=0.875 //x2=57.435 //y2=0.375
cc_872 ( N_GND_c_24_p N_noxref_49_c_10358_n ) capacitor c=0.00352952f \
 //x=84.73 //y=0 //x2=59.995 //y2=0.995
cc_873 ( N_GND_c_305_p N_noxref_49_c_10358_n ) capacitor c=0.00934524f \
 //x=61.62 //y=0 //x2=59.995 //y2=0.995
cc_874 ( N_GND_c_24_p N_noxref_49_c_10360_n ) capacitor c=0.00254475f \
 //x=84.73 //y=0 //x2=60.08 //y2=0.625
cc_875 ( N_GND_c_305_p N_noxref_49_c_10360_n ) capacitor c=0.0140928f \
 //x=61.62 //y=0 //x2=60.08 //y2=0.625
cc_876 ( N_GND_M35_noxref_d N_noxref_49_c_10360_n ) capacitor c=6.21394e-19 \
 //x=57.865 //y=0.875 //x2=60.08 //y2=0.625
cc_877 ( N_GND_c_24_p N_noxref_49_c_10363_n ) capacitor c=0.0105317f //x=84.73 \
 //y=0 //x2=60.965 //y2=0.54
cc_878 ( N_GND_c_305_p N_noxref_49_c_10363_n ) capacitor c=0.0364215f \
 //x=61.62 //y=0 //x2=60.965 //y2=0.54
cc_879 ( N_GND_c_24_p N_noxref_49_c_10365_n ) capacitor c=0.00254232f \
 //x=84.73 //y=0 //x2=61.05 //y2=0.625
cc_880 ( N_GND_c_305_p N_noxref_49_c_10365_n ) capacitor c=0.0140304f \
 //x=61.62 //y=0 //x2=61.05 //y2=0.625
cc_881 ( N_GND_c_16_p N_noxref_49_c_10365_n ) capacitor c=0.0404137f //x=61.79 \
 //y=0 //x2=61.05 //y2=0.625
cc_882 ( N_GND_M35_noxref_d N_noxref_49_M36_noxref_d ) capacitor c=0.00162435f \
 //x=57.865 //y=0.875 //x2=58.84 //y2=0.91
cc_883 ( N_GND_c_15_p N_noxref_49_M37_noxref_s ) capacitor c=8.16352e-19 \
 //x=56.98 //y=0 //x2=59.945 //y2=0.375
cc_884 ( N_GND_c_16_p N_noxref_49_M37_noxref_s ) capacitor c=0.00183576f \
 //x=61.79 //y=0 //x2=59.945 //y2=0.375
cc_885 ( N_GND_c_24_p N_noxref_50_c_10410_n ) capacitor c=0.00517234f \
 //x=84.73 //y=0 //x2=63.37 //y2=1.58
cc_886 ( N_GND_c_316_p N_noxref_50_c_10410_n ) capacitor c=0.00112872f \
 //x=62.885 //y=0 //x2=63.37 //y2=1.58
cc_887 ( N_GND_c_323_p N_noxref_50_c_10410_n ) capacitor c=0.0018229f \
 //x=64.95 //y=0 //x2=63.37 //y2=1.58
cc_888 ( N_GND_M38_noxref_d N_noxref_50_c_10410_n ) capacitor c=0.008625f \
 //x=62.78 //y=0.865 //x2=63.37 //y2=1.58
cc_889 ( N_GND_c_24_p N_noxref_50_c_10414_n ) capacitor c=0.00259029f \
 //x=84.73 //y=0 //x2=63.455 //y2=0.615
cc_890 ( N_GND_c_323_p N_noxref_50_c_10414_n ) capacitor c=0.0146901f \
 //x=64.95 //y=0 //x2=63.455 //y2=0.615
cc_891 ( N_GND_M38_noxref_d N_noxref_50_c_10414_n ) capacitor c=0.033812f \
 //x=62.78 //y=0.865 //x2=63.455 //y2=0.615
cc_892 ( N_GND_c_16_p N_noxref_50_c_10417_n ) capacitor c=2.91423e-19 \
 //x=61.79 //y=0 //x2=63.455 //y2=1.495
cc_893 ( N_GND_c_24_p N_noxref_50_c_10418_n ) capacitor c=0.0106919f //x=84.73 \
 //y=0 //x2=64.34 //y2=0.53
cc_894 ( N_GND_c_323_p N_noxref_50_c_10418_n ) capacitor c=0.0374253f \
 //x=64.95 //y=0 //x2=64.34 //y2=0.53
cc_895 ( N_GND_c_24_p N_noxref_50_c_10420_n ) capacitor c=0.00258845f \
 //x=84.73 //y=0 //x2=64.425 //y2=0.615
cc_896 ( N_GND_c_323_p N_noxref_50_c_10420_n ) capacitor c=0.0146256f \
 //x=64.95 //y=0 //x2=64.425 //y2=0.615
cc_897 ( N_GND_c_17_p N_noxref_50_c_10420_n ) capacitor c=0.0431718f //x=65.12 \
 //y=0 //x2=64.425 //y2=0.615
cc_898 ( N_GND_c_24_p N_noxref_50_M38_noxref_s ) capacitor c=0.00259029f \
 //x=84.73 //y=0 //x2=62.35 //y2=0.365
cc_899 ( N_GND_c_316_p N_noxref_50_M38_noxref_s ) capacitor c=0.0146901f \
 //x=62.885 //y=0 //x2=62.35 //y2=0.365
cc_900 ( N_GND_c_16_p N_noxref_50_M38_noxref_s ) capacitor c=0.0583534f \
 //x=61.79 //y=0 //x2=62.35 //y2=0.365
cc_901 ( N_GND_c_17_p N_noxref_50_M38_noxref_s ) capacitor c=0.00198043f \
 //x=65.12 //y=0 //x2=62.35 //y2=0.365
cc_902 ( N_GND_M38_noxref_d N_noxref_50_M38_noxref_s ) capacitor c=0.0334197f \
 //x=62.78 //y=0.865 //x2=62.35 //y2=0.365
cc_903 ( N_GND_c_24_p N_noxref_51_c_10461_n ) capacitor c=0.00517234f \
 //x=84.73 //y=0 //x2=66.7 //y2=1.58
cc_904 ( N_GND_c_340_p N_noxref_51_c_10461_n ) capacitor c=0.00112872f \
 //x=66.215 //y=0 //x2=66.7 //y2=1.58
cc_905 ( N_GND_c_347_p N_noxref_51_c_10461_n ) capacitor c=0.0018229f \
 //x=68.28 //y=0 //x2=66.7 //y2=1.58
cc_906 ( N_GND_M40_noxref_d N_noxref_51_c_10461_n ) capacitor c=0.008625f \
 //x=66.11 //y=0.865 //x2=66.7 //y2=1.58
cc_907 ( N_GND_c_24_p N_noxref_51_c_10465_n ) capacitor c=0.00259029f \
 //x=84.73 //y=0 //x2=66.785 //y2=0.615
cc_908 ( N_GND_c_347_p N_noxref_51_c_10465_n ) capacitor c=0.0146901f \
 //x=68.28 //y=0 //x2=66.785 //y2=0.615
cc_909 ( N_GND_M40_noxref_d N_noxref_51_c_10465_n ) capacitor c=0.033812f \
 //x=66.11 //y=0.865 //x2=66.785 //y2=0.615
cc_910 ( N_GND_c_17_p N_noxref_51_c_10468_n ) capacitor c=2.91423e-19 \
 //x=65.12 //y=0 //x2=66.785 //y2=1.495
cc_911 ( N_GND_c_24_p N_noxref_51_c_10469_n ) capacitor c=0.0106919f //x=84.73 \
 //y=0 //x2=67.67 //y2=0.53
cc_912 ( N_GND_c_347_p N_noxref_51_c_10469_n ) capacitor c=0.0374253f \
 //x=68.28 //y=0 //x2=67.67 //y2=0.53
cc_913 ( N_GND_c_24_p N_noxref_51_c_10471_n ) capacitor c=0.00258845f \
 //x=84.73 //y=0 //x2=67.755 //y2=0.615
cc_914 ( N_GND_c_347_p N_noxref_51_c_10471_n ) capacitor c=0.0146256f \
 //x=68.28 //y=0 //x2=67.755 //y2=0.615
cc_915 ( N_GND_c_18_p N_noxref_51_c_10471_n ) capacitor c=0.0431718f //x=68.45 \
 //y=0 //x2=67.755 //y2=0.615
cc_916 ( N_GND_c_24_p N_noxref_51_M40_noxref_s ) capacitor c=0.00259029f \
 //x=84.73 //y=0 //x2=65.68 //y2=0.365
cc_917 ( N_GND_c_340_p N_noxref_51_M40_noxref_s ) capacitor c=0.0146901f \
 //x=66.215 //y=0 //x2=65.68 //y2=0.365
cc_918 ( N_GND_c_17_p N_noxref_51_M40_noxref_s ) capacitor c=0.058339f \
 //x=65.12 //y=0 //x2=65.68 //y2=0.365
cc_919 ( N_GND_c_18_p N_noxref_51_M40_noxref_s ) capacitor c=0.00198098f \
 //x=68.45 //y=0 //x2=65.68 //y2=0.365
cc_920 ( N_GND_M40_noxref_d N_noxref_51_M40_noxref_s ) capacitor c=0.0334197f \
 //x=66.11 //y=0.865 //x2=65.68 //y2=0.365
cc_921 ( N_GND_c_24_p N_noxref_52_c_10512_n ) capacitor c=0.00517576f \
 //x=84.73 //y=0 //x2=69.925 //y2=1.59
cc_922 ( N_GND_c_354_p N_noxref_52_c_10512_n ) capacitor c=0.00111448f \
 //x=69.44 //y=0 //x2=69.925 //y2=1.59
cc_923 ( N_GND_c_212_p N_noxref_52_c_10512_n ) capacitor c=0.00180612f \
 //x=73.09 //y=0 //x2=69.925 //y2=1.59
cc_924 ( N_GND_M42_noxref_d N_noxref_52_c_10512_n ) capacitor c=0.00853078f \
 //x=69.335 //y=0.875 //x2=69.925 //y2=1.59
cc_925 ( N_GND_c_24_p N_noxref_52_c_10516_n ) capacitor c=0.00254475f \
 //x=84.73 //y=0 //x2=70.01 //y2=0.625
cc_926 ( N_GND_c_212_p N_noxref_52_c_10516_n ) capacitor c=0.0140928f \
 //x=73.09 //y=0 //x2=70.01 //y2=0.625
cc_927 ( N_GND_M42_noxref_d N_noxref_52_c_10516_n ) capacitor c=0.033954f \
 //x=69.335 //y=0.875 //x2=70.01 //y2=0.625
cc_928 ( N_GND_c_24_p N_noxref_52_c_10519_n ) capacitor c=0.0105304f //x=84.73 \
 //y=0 //x2=70.895 //y2=0.54
cc_929 ( N_GND_c_212_p N_noxref_52_c_10519_n ) capacitor c=0.0361183f \
 //x=73.09 //y=0 //x2=70.895 //y2=0.54
cc_930 ( N_GND_c_24_p N_noxref_52_M42_noxref_s ) capacitor c=0.00531539f \
 //x=84.73 //y=0 //x2=68.905 //y2=0.375
cc_931 ( N_GND_c_354_p N_noxref_52_M42_noxref_s ) capacitor c=0.0140928f \
 //x=69.44 //y=0 //x2=68.905 //y2=0.375
cc_932 ( N_GND_c_212_p N_noxref_52_M42_noxref_s ) capacitor c=0.0138368f \
 //x=73.09 //y=0 //x2=68.905 //y2=0.375
cc_933 ( N_GND_c_18_p N_noxref_52_M42_noxref_s ) capacitor c=0.0696963f \
 //x=68.45 //y=0 //x2=68.905 //y2=0.375
cc_934 ( N_GND_c_19_p N_noxref_52_M42_noxref_s ) capacitor c=3.31601e-19 \
 //x=73.26 //y=0 //x2=68.905 //y2=0.375
cc_935 ( N_GND_M42_noxref_d N_noxref_52_M42_noxref_s ) capacitor c=0.033718f \
 //x=69.335 //y=0.875 //x2=68.905 //y2=0.375
cc_936 ( N_GND_c_24_p N_noxref_53_c_10563_n ) capacitor c=0.00375441f \
 //x=84.73 //y=0 //x2=71.465 //y2=0.995
cc_937 ( N_GND_c_212_p N_noxref_53_c_10563_n ) capacitor c=0.00944862f \
 //x=73.09 //y=0 //x2=71.465 //y2=0.995
cc_938 ( N_GND_c_24_p N_noxref_53_c_10565_n ) capacitor c=0.00277579f \
 //x=84.73 //y=0 //x2=71.55 //y2=0.625
cc_939 ( N_GND_c_212_p N_noxref_53_c_10565_n ) capacitor c=0.0142586f \
 //x=73.09 //y=0 //x2=71.55 //y2=0.625
cc_940 ( N_GND_M42_noxref_d N_noxref_53_c_10565_n ) capacitor c=6.21394e-19 \
 //x=69.335 //y=0.875 //x2=71.55 //y2=0.625
cc_941 ( N_GND_c_24_p N_noxref_53_c_10568_n ) capacitor c=0.0114469f //x=84.73 \
 //y=0 //x2=72.435 //y2=0.54
cc_942 ( N_GND_c_212_p N_noxref_53_c_10568_n ) capacitor c=0.0365589f \
 //x=73.09 //y=0 //x2=72.435 //y2=0.54
cc_943 ( N_GND_c_24_p N_noxref_53_c_10570_n ) capacitor c=0.00277442f \
 //x=84.73 //y=0 //x2=72.52 //y2=0.625
cc_944 ( N_GND_c_212_p N_noxref_53_c_10570_n ) capacitor c=0.014197f //x=73.09 \
 //y=0 //x2=72.52 //y2=0.625
cc_945 ( N_GND_c_19_p N_noxref_53_c_10570_n ) capacitor c=0.0400472f //x=73.26 \
 //y=0 //x2=72.52 //y2=0.625
cc_946 ( N_GND_M42_noxref_d N_noxref_53_M43_noxref_d ) capacitor c=0.00162435f \
 //x=69.335 //y=0.875 //x2=70.31 //y2=0.91
cc_947 ( N_GND_c_18_p N_noxref_53_M44_noxref_s ) capacitor c=8.16352e-19 \
 //x=68.45 //y=0 //x2=71.415 //y2=0.375
cc_948 ( N_GND_c_19_p N_noxref_53_M44_noxref_s ) capacitor c=0.00183576f \
 //x=73.26 //y=0 //x2=71.415 //y2=0.375
cc_949 ( N_GND_c_24_p N_noxref_54_c_10615_n ) capacitor c=0.00547799f \
 //x=84.73 //y=0 //x2=74.84 //y2=1.58
cc_950 ( N_GND_c_213_p N_noxref_54_c_10615_n ) capacitor c=0.00112964f \
 //x=74.355 //y=0 //x2=74.84 //y2=1.58
cc_951 ( N_GND_c_451_p N_noxref_54_c_10615_n ) capacitor c=0.00182382f \
 //x=76.42 //y=0 //x2=74.84 //y2=1.58
cc_952 ( N_GND_M45_noxref_d N_noxref_54_c_10615_n ) capacitor c=0.0092166f \
 //x=74.25 //y=0.865 //x2=74.84 //y2=1.58
cc_953 ( N_GND_c_24_p N_noxref_54_c_10619_n ) capacitor c=0.00282859f \
 //x=84.73 //y=0 //x2=74.925 //y2=0.615
cc_954 ( N_GND_c_451_p N_noxref_54_c_10619_n ) capacitor c=0.0148634f \
 //x=76.42 //y=0 //x2=74.925 //y2=0.615
cc_955 ( N_GND_M45_noxref_d N_noxref_54_c_10619_n ) capacitor c=0.0336822f \
 //x=74.25 //y=0.865 //x2=74.925 //y2=0.615
cc_956 ( N_GND_c_19_p N_noxref_54_c_10622_n ) capacitor c=2.91423e-19 \
 //x=73.26 //y=0 //x2=74.925 //y2=1.495
cc_957 ( N_GND_c_24_p N_noxref_54_c_10623_n ) capacitor c=0.00972362f \
 //x=84.73 //y=0 //x2=75.81 //y2=0.53
cc_958 ( N_GND_c_451_p N_noxref_54_c_10623_n ) capacitor c=0.0375226f \
 //x=76.42 //y=0 //x2=75.81 //y2=0.53
cc_959 ( N_GND_c_24_p N_noxref_54_c_10625_n ) capacitor c=0.00212661f \
 //x=84.73 //y=0 //x2=75.895 //y2=0.615
cc_960 ( N_GND_c_451_p N_noxref_54_c_10625_n ) capacitor c=0.0143168f \
 //x=76.42 //y=0 //x2=75.895 //y2=0.615
cc_961 ( N_GND_c_20_p N_noxref_54_c_10625_n ) capacitor c=0.0554337f //x=76.59 \
 //y=0 //x2=75.895 //y2=0.615
cc_962 ( N_GND_c_24_p N_noxref_54_M45_noxref_s ) capacitor c=0.00282937f \
 //x=84.73 //y=0 //x2=73.82 //y2=0.365
cc_963 ( N_GND_c_213_p N_noxref_54_M45_noxref_s ) capacitor c=0.0148639f \
 //x=74.355 //y=0 //x2=73.82 //y2=0.365
cc_964 ( N_GND_c_19_p N_noxref_54_M45_noxref_s ) capacitor c=0.058813f \
 //x=73.26 //y=0 //x2=73.82 //y2=0.365
cc_965 ( N_GND_c_20_p N_noxref_54_M45_noxref_s ) capacitor c=0.00181744f \
 //x=76.59 //y=0 //x2=73.82 //y2=0.365
cc_966 ( N_GND_M45_noxref_d N_noxref_54_M45_noxref_s ) capacitor c=0.0333456f \
 //x=74.25 //y=0.865 //x2=73.82 //y2=0.365
cc_967 ( N_GND_c_454_p N_noxref_55_c_10672_n ) capacitor c=8.01905e-19 \
 //x=77.685 //y=0 //x2=78.17 //y2=1.58
cc_968 ( N_GND_c_460_p N_noxref_55_c_10672_n ) capacitor c=0.00161527f \
 //x=79.75 //y=0 //x2=78.17 //y2=1.58
cc_969 ( N_GND_M47_noxref_d N_noxref_55_c_10672_n ) capacitor c=0.0073276f \
 //x=77.58 //y=0.865 //x2=78.17 //y2=1.58
cc_970 ( N_GND_c_24_p N_noxref_55_c_10675_n ) capacitor c=0.00212661f \
 //x=84.73 //y=0 //x2=78.255 //y2=0.615
cc_971 ( N_GND_c_460_p N_noxref_55_c_10675_n ) capacitor c=0.0143168f \
 //x=79.75 //y=0 //x2=78.255 //y2=0.615
cc_972 ( N_GND_M47_noxref_d N_noxref_55_c_10675_n ) capacitor c=0.0336587f \
 //x=77.58 //y=0.865 //x2=78.255 //y2=0.615
cc_973 ( N_GND_c_20_p N_noxref_55_c_10678_n ) capacitor c=2.91423e-19 \
 //x=76.59 //y=0 //x2=78.255 //y2=1.495
cc_974 ( N_GND_c_24_p N_noxref_55_c_10679_n ) capacitor c=0.00884129f \
 //x=84.73 //y=0 //x2=79.14 //y2=0.53
cc_975 ( N_GND_c_460_p N_noxref_55_c_10679_n ) capacitor c=0.0373651f \
 //x=79.75 //y=0 //x2=79.14 //y2=0.53
cc_976 ( N_GND_c_24_p N_noxref_55_c_10681_n ) capacitor c=0.00212661f \
 //x=84.73 //y=0 //x2=79.225 //y2=0.615
cc_977 ( N_GND_c_460_p N_noxref_55_c_10681_n ) capacitor c=0.0143168f \
 //x=79.75 //y=0 //x2=79.225 //y2=0.615
cc_978 ( N_GND_c_21_p N_noxref_55_c_10681_n ) capacitor c=0.0548042f //x=79.92 \
 //y=0 //x2=79.225 //y2=0.615
cc_979 ( N_GND_c_24_p N_noxref_55_M47_noxref_s ) capacitor c=0.00212661f \
 //x=84.73 //y=0 //x2=77.15 //y2=0.365
cc_980 ( N_GND_c_454_p N_noxref_55_M47_noxref_s ) capacitor c=0.0143168f \
 //x=77.685 //y=0 //x2=77.15 //y2=0.365
cc_981 ( N_GND_c_20_p N_noxref_55_M47_noxref_s ) capacitor c=0.0561194f \
 //x=76.59 //y=0 //x2=77.15 //y2=0.365
cc_982 ( N_GND_c_21_p N_noxref_55_M47_noxref_s ) capacitor c=0.0022128f \
 //x=79.92 //y=0 //x2=77.15 //y2=0.365
cc_983 ( N_GND_M47_noxref_d N_noxref_55_M47_noxref_s ) capacitor c=0.0332904f \
 //x=77.58 //y=0.865 //x2=77.15 //y2=0.365
cc_984 ( N_GND_c_476_p N_noxref_56_c_10727_n ) capacitor c=8.01912e-19 \
 //x=81.015 //y=0 //x2=81.5 //y2=1.58
cc_985 ( N_GND_c_482_p N_noxref_56_c_10727_n ) capacitor c=0.00161527f \
 //x=83.08 //y=0 //x2=81.5 //y2=1.58
cc_986 ( N_GND_M49_noxref_d N_noxref_56_c_10727_n ) capacitor c=0.0073482f \
 //x=80.91 //y=0.865 //x2=81.5 //y2=1.58
cc_987 ( N_GND_c_24_p N_noxref_56_c_10730_n ) capacitor c=0.00212661f \
 //x=84.73 //y=0 //x2=81.585 //y2=0.615
cc_988 ( N_GND_c_482_p N_noxref_56_c_10730_n ) capacitor c=0.0143168f \
 //x=83.08 //y=0 //x2=81.585 //y2=0.615
cc_989 ( N_GND_M49_noxref_d N_noxref_56_c_10730_n ) capacitor c=0.0336587f \
 //x=80.91 //y=0.865 //x2=81.585 //y2=0.615
cc_990 ( N_GND_c_21_p N_noxref_56_c_10733_n ) capacitor c=2.91423e-19 \
 //x=79.92 //y=0 //x2=81.585 //y2=1.495
cc_991 ( N_GND_c_24_p N_noxref_56_c_10734_n ) capacitor c=0.0119802f //x=84.73 \
 //y=0 //x2=82.47 //y2=0.53
cc_992 ( N_GND_c_482_p N_noxref_56_c_10734_n ) capacitor c=0.0371788f \
 //x=83.08 //y=0 //x2=82.47 //y2=0.53
cc_993 ( N_GND_c_24_p N_noxref_56_c_10736_n ) capacitor c=0.00579412f \
 //x=84.73 //y=0 //x2=82.555 //y2=0.615
cc_994 ( N_GND_c_482_p N_noxref_56_c_10736_n ) capacitor c=0.0144285f \
 //x=83.08 //y=0 //x2=82.555 //y2=0.615
cc_995 ( N_GND_c_995_p N_noxref_56_c_10736_n ) capacitor c=0.00114292f \
 //x=83.88 //y=0.45 //x2=82.555 //y2=0.615
cc_996 ( N_GND_c_22_p N_noxref_56_c_10736_n ) capacitor c=0.042944f //x=83.25 \
 //y=0 //x2=82.555 //y2=0.615
cc_997 ( N_GND_c_24_p N_noxref_56_M49_noxref_s ) capacitor c=0.00212661f \
 //x=84.73 //y=0 //x2=80.48 //y2=0.365
cc_998 ( N_GND_c_476_p N_noxref_56_M49_noxref_s ) capacitor c=0.0143168f \
 //x=81.015 //y=0 //x2=80.48 //y2=0.365
cc_999 ( N_GND_c_21_p N_noxref_56_M49_noxref_s ) capacitor c=0.0555228f \
 //x=79.92 //y=0 //x2=80.48 //y2=0.365
cc_1000 ( N_GND_c_22_p N_noxref_56_M49_noxref_s ) capacitor c=0.00201114f \
 //x=83.25 //y=0 //x2=80.48 //y2=0.365
cc_1001 ( N_GND_M49_noxref_d N_noxref_56_M49_noxref_s ) capacitor c=0.0332904f \
 //x=80.91 //y=0.865 //x2=80.48 //y2=0.365
cc_1002 ( N_GND_M51_noxref_s N_noxref_56_M49_noxref_s ) capacitor \
 c=0.00114292f //x=83.745 //y=0.37 //x2=80.48 //y2=0.365
cc_1003 ( N_GND_c_22_p Q ) capacitor c=8.10282e-19 //x=83.25 //y=0 //x2=84.73 \
 //y2=2.22
cc_1004 ( N_GND_c_24_p N_Q_c_10784_n ) capacitor c=0.00180637f //x=84.73 //y=0 \
 //x2=84.645 //y2=2.08
cc_1005 ( N_GND_c_23_p N_Q_c_10784_n ) capacitor c=0.0301661f //x=84.85 //y=0 \
 //x2=84.645 //y2=2.08
cc_1006 ( N_GND_M51_noxref_s N_Q_c_10784_n ) capacitor c=0.00999304f \
 //x=83.745 //y=0.37 //x2=84.645 //y2=2.08
cc_1007 ( N_GND_c_24_p N_Q_M51_noxref_d ) capacitor c=0.00194883f //x=84.73 \
 //y=0 //x2=84.175 //y2=0.91
cc_1008 ( N_GND_c_511_p N_Q_M51_noxref_d ) capacitor c=0.0146043f //x=84.28 \
 //y=0.535 //x2=84.175 //y2=0.91
cc_1009 ( N_GND_c_22_p N_Q_M51_noxref_d ) capacitor c=0.00923478f //x=83.25 \
 //y=0 //x2=84.175 //y2=0.91
cc_1010 ( N_GND_c_23_p N_Q_M51_noxref_d ) capacitor c=0.00950401f //x=84.85 \
 //y=0 //x2=84.175 //y2=0.91
cc_1011 ( N_GND_M51_noxref_s N_Q_M51_noxref_d ) capacitor c=0.0768153f \
 //x=83.745 //y=0.37 //x2=84.175 //y2=0.91
cc_1012 ( N_VDD_c_1035_p N_noxref_3_c_2157_n ) capacitor c=0.00469095f \
 //x=84.73 //y=7.4 //x2=2.025 //y2=5.2
cc_1013 ( N_VDD_c_1036_p N_noxref_3_c_2157_n ) capacitor c=4.3394e-19 \
 //x=1.585 //y=7.4 //x2=2.025 //y2=5.2
cc_1014 ( N_VDD_c_1037_p N_noxref_3_c_2157_n ) capacitor c=4.48693e-19 \
 //x=2.465 //y=7.4 //x2=2.025 //y2=5.2
cc_1015 ( N_VDD_M53_noxref_d N_noxref_3_c_2157_n ) capacitor c=0.0128947f \
 //x=1.525 //y=5.02 //x2=2.025 //y2=5.2
cc_1016 ( N_VDD_c_1012_n N_noxref_3_c_2161_n ) capacitor c=0.00989999f \
 //x=0.74 //y=7.4 //x2=1.315 //y2=5.2
cc_1017 ( N_VDD_M52_noxref_s N_noxref_3_c_2161_n ) capacitor c=0.087833f \
 //x=0.655 //y=5.02 //x2=1.315 //y2=5.2
cc_1018 ( N_VDD_c_1035_p N_noxref_3_c_2163_n ) capacitor c=0.00307195f \
 //x=84.73 //y=7.4 //x2=2.505 //y2=5.2
cc_1019 ( N_VDD_c_1037_p N_noxref_3_c_2163_n ) capacitor c=7.73167e-19 \
 //x=2.465 //y=7.4 //x2=2.505 //y2=5.2
cc_1020 ( N_VDD_M55_noxref_d N_noxref_3_c_2163_n ) capacitor c=0.0161518f \
 //x=2.405 //y=5.02 //x2=2.505 //y2=5.2
cc_1021 ( N_VDD_c_1012_n N_noxref_3_c_2130_n ) capacitor c=0.00159771f \
 //x=0.74 //y=7.4 //x2=2.59 //y2=2.59
cc_1022 ( N_VDD_c_1013_n N_noxref_3_c_2130_n ) capacitor c=0.0452382f //x=3.33 \
 //y=7.4 //x2=2.59 //y2=2.59
cc_1023 ( N_VDD_c_1035_p N_noxref_3_c_2132_n ) capacitor c=9.23542e-19 \
 //x=84.73 //y=7.4 //x2=4.44 //y2=2.08
cc_1024 ( N_VDD_c_1013_n N_noxref_3_c_2132_n ) capacitor c=0.0157357f //x=3.33 \
 //y=7.4 //x2=4.44 //y2=2.08
cc_1025 ( N_VDD_M56_noxref_s N_noxref_3_c_2132_n ) capacitor c=0.0123142f \
 //x=4.285 //y=5.02 //x2=4.44 //y2=2.08
cc_1026 ( N_VDD_c_1035_p N_noxref_3_c_2133_n ) capacitor c=9.10347e-19 \
 //x=84.73 //y=7.4 //x2=9.25 //y2=2.08
cc_1027 ( N_VDD_c_1014_n N_noxref_3_c_2133_n ) capacitor c=0.013427f //x=8.14 \
 //y=7.4 //x2=9.25 //y2=2.08
cc_1028 ( N_VDD_M62_noxref_s N_noxref_3_c_2133_n ) capacitor c=0.0125322f \
 //x=9.095 //y=5.02 //x2=9.25 //y2=2.08
cc_1029 ( N_VDD_c_1052_p N_noxref_3_M56_noxref_g ) capacitor c=0.00749687f \
 //x=5.215 //y=7.4 //x2=4.64 //y2=6.02
cc_1030 ( N_VDD_M56_noxref_s N_noxref_3_M56_noxref_g ) capacitor c=0.0477201f \
 //x=4.285 //y=5.02 //x2=4.64 //y2=6.02
cc_1031 ( N_VDD_c_1052_p N_noxref_3_M57_noxref_g ) capacitor c=0.00675175f \
 //x=5.215 //y=7.4 //x2=5.08 //y2=6.02
cc_1032 ( N_VDD_M57_noxref_d N_noxref_3_M57_noxref_g ) capacitor c=0.015318f \
 //x=5.155 //y=5.02 //x2=5.08 //y2=6.02
cc_1033 ( N_VDD_c_1056_p N_noxref_3_M62_noxref_g ) capacitor c=0.00749687f \
 //x=10.025 //y=7.4 //x2=9.45 //y2=6.02
cc_1034 ( N_VDD_M62_noxref_s N_noxref_3_M62_noxref_g ) capacitor c=0.0477201f \
 //x=9.095 //y=5.02 //x2=9.45 //y2=6.02
cc_1035 ( N_VDD_c_1056_p N_noxref_3_M63_noxref_g ) capacitor c=0.00675175f \
 //x=10.025 //y=7.4 //x2=9.89 //y2=6.02
cc_1036 ( N_VDD_M63_noxref_d N_noxref_3_M63_noxref_g ) capacitor c=0.015318f \
 //x=9.965 //y=5.02 //x2=9.89 //y2=6.02
cc_1037 ( N_VDD_c_1013_n N_noxref_3_c_2182_n ) capacitor c=0.00757682f \
 //x=3.33 //y=7.4 //x2=4.715 //y2=4.79
cc_1038 ( N_VDD_M56_noxref_s N_noxref_3_c_2182_n ) capacitor c=0.00445134f \
 //x=4.285 //y=5.02 //x2=4.715 //y2=4.79
cc_1039 ( N_VDD_c_1014_n N_noxref_3_c_2184_n ) capacitor c=0.00757682f \
 //x=8.14 //y=7.4 //x2=9.525 //y2=4.79
cc_1040 ( N_VDD_M62_noxref_s N_noxref_3_c_2184_n ) capacitor c=0.00444914f \
 //x=9.095 //y=5.02 //x2=9.525 //y2=4.79
cc_1041 ( N_VDD_c_1035_p N_noxref_3_M52_noxref_d ) capacitor c=0.00582349f \
 //x=84.73 //y=7.4 //x2=1.085 //y2=5.02
cc_1042 ( N_VDD_c_1036_p N_noxref_3_M52_noxref_d ) capacitor c=0.0138103f \
 //x=1.585 //y=7.4 //x2=1.085 //y2=5.02
cc_1043 ( N_VDD_c_1013_n N_noxref_3_M52_noxref_d ) capacitor c=6.94454e-19 \
 //x=3.33 //y=7.4 //x2=1.085 //y2=5.02
cc_1044 ( N_VDD_M53_noxref_d N_noxref_3_M52_noxref_d ) capacitor c=0.0664752f \
 //x=1.525 //y=5.02 //x2=1.085 //y2=5.02
cc_1045 ( N_VDD_c_1035_p N_noxref_3_M54_noxref_d ) capacitor c=0.00285083f \
 //x=84.73 //y=7.4 //x2=1.965 //y2=5.02
cc_1046 ( N_VDD_c_1037_p N_noxref_3_M54_noxref_d ) capacitor c=0.0140984f \
 //x=2.465 //y=7.4 //x2=1.965 //y2=5.02
cc_1047 ( N_VDD_c_1013_n N_noxref_3_M54_noxref_d ) capacitor c=0.0120541f \
 //x=3.33 //y=7.4 //x2=1.965 //y2=5.02
cc_1048 ( N_VDD_M52_noxref_s N_noxref_3_M54_noxref_d ) capacitor c=0.00111971f \
 //x=0.655 //y=5.02 //x2=1.965 //y2=5.02
cc_1049 ( N_VDD_M53_noxref_d N_noxref_3_M54_noxref_d ) capacitor c=0.0664752f \
 //x=1.525 //y=5.02 //x2=1.965 //y2=5.02
cc_1050 ( N_VDD_M55_noxref_d N_noxref_3_M54_noxref_d ) capacitor c=0.0664752f \
 //x=2.405 //y=5.02 //x2=1.965 //y2=5.02
cc_1051 ( N_VDD_M56_noxref_s N_noxref_3_M54_noxref_d ) capacitor c=3.73257e-19 \
 //x=4.285 //y=5.02 //x2=1.965 //y2=5.02
cc_1052 ( N_VDD_c_1035_p N_noxref_4_c_2377_n ) capacitor c=0.00444892f \
 //x=84.73 //y=7.4 //x2=10.465 //y2=5.155
cc_1053 ( N_VDD_c_1056_p N_noxref_4_c_2377_n ) capacitor c=4.31931e-19 \
 //x=10.025 //y=7.4 //x2=10.465 //y2=5.155
cc_1054 ( N_VDD_c_1077_p N_noxref_4_c_2377_n ) capacitor c=4.31931e-19 \
 //x=10.905 //y=7.4 //x2=10.465 //y2=5.155
cc_1055 ( N_VDD_M63_noxref_d N_noxref_4_c_2377_n ) capacitor c=0.0112985f \
 //x=9.965 //y=5.02 //x2=10.465 //y2=5.155
cc_1056 ( N_VDD_c_1014_n N_noxref_4_c_2381_n ) capacitor c=0.00863585f \
 //x=8.14 //y=7.4 //x2=9.755 //y2=5.155
cc_1057 ( N_VDD_M62_noxref_s N_noxref_4_c_2381_n ) capacitor c=0.0831083f \
 //x=9.095 //y=5.02 //x2=9.755 //y2=5.155
cc_1058 ( N_VDD_c_1035_p N_noxref_4_c_2383_n ) capacitor c=0.0044221f \
 //x=84.73 //y=7.4 //x2=11.345 //y2=5.155
cc_1059 ( N_VDD_c_1077_p N_noxref_4_c_2383_n ) capacitor c=4.31931e-19 \
 //x=10.905 //y=7.4 //x2=11.345 //y2=5.155
cc_1060 ( N_VDD_c_1083_p N_noxref_4_c_2383_n ) capacitor c=4.31931e-19 \
 //x=11.785 //y=7.4 //x2=11.345 //y2=5.155
cc_1061 ( N_VDD_M65_noxref_d N_noxref_4_c_2383_n ) capacitor c=0.0112985f \
 //x=10.845 //y=5.02 //x2=11.345 //y2=5.155
cc_1062 ( N_VDD_c_1035_p N_noxref_4_c_2387_n ) capacitor c=0.00434174f \
 //x=84.73 //y=7.4 //x2=12.125 //y2=5.155
cc_1063 ( N_VDD_c_1083_p N_noxref_4_c_2387_n ) capacitor c=7.46626e-19 \
 //x=11.785 //y=7.4 //x2=12.125 //y2=5.155
cc_1064 ( N_VDD_c_1087_p N_noxref_4_c_2387_n ) capacitor c=0.00198565f \
 //x=12.78 //y=7.4 //x2=12.125 //y2=5.155
cc_1065 ( N_VDD_M67_noxref_d N_noxref_4_c_2387_n ) capacitor c=0.0112985f \
 //x=11.725 //y=5.02 //x2=12.125 //y2=5.155
cc_1066 ( N_VDD_c_1015_n N_noxref_4_c_2364_n ) capacitor c=0.042636f //x=12.95 \
 //y=7.4 //x2=12.21 //y2=2.59
cc_1067 ( N_VDD_c_1035_p N_noxref_4_c_2365_n ) capacitor c=0.00125279f \
 //x=84.73 //y=7.4 //x2=14.06 //y2=2.08
cc_1068 ( N_VDD_c_1091_p N_noxref_4_c_2365_n ) capacitor c=2.87256e-19 \
 //x=14.535 //y=7.4 //x2=14.06 //y2=2.08
cc_1069 ( N_VDD_c_1015_n N_noxref_4_c_2365_n ) capacitor c=0.0133961f \
 //x=12.95 //y=7.4 //x2=14.06 //y2=2.08
cc_1070 ( N_VDD_c_1091_p N_noxref_4_M68_noxref_g ) capacitor c=0.00726866f \
 //x=14.535 //y=7.4 //x2=13.96 //y2=6.02
cc_1071 ( N_VDD_M68_noxref_s N_noxref_4_M68_noxref_g ) capacitor c=0.054195f \
 //x=13.605 //y=5.02 //x2=13.96 //y2=6.02
cc_1072 ( N_VDD_c_1091_p N_noxref_4_M69_noxref_g ) capacitor c=0.00672952f \
 //x=14.535 //y=7.4 //x2=14.4 //y2=6.02
cc_1073 ( N_VDD_M69_noxref_d N_noxref_4_M69_noxref_g ) capacitor c=0.015318f \
 //x=14.475 //y=5.02 //x2=14.4 //y2=6.02
cc_1074 ( N_VDD_c_1015_n N_noxref_4_c_2399_n ) capacitor c=0.015293f //x=12.95 \
 //y=7.4 //x2=14.06 //y2=4.7
cc_1075 ( N_VDD_c_1035_p N_noxref_4_M62_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=9.525 //y2=5.02
cc_1076 ( N_VDD_c_1056_p N_noxref_4_M62_noxref_d ) capacitor c=0.014035f \
 //x=10.025 //y=7.4 //x2=9.525 //y2=5.02
cc_1077 ( N_VDD_M63_noxref_d N_noxref_4_M62_noxref_d ) capacitor c=0.0664752f \
 //x=9.965 //y=5.02 //x2=9.525 //y2=5.02
cc_1078 ( N_VDD_c_1035_p N_noxref_4_M64_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=10.405 //y2=5.02
cc_1079 ( N_VDD_c_1077_p N_noxref_4_M64_noxref_d ) capacitor c=0.014035f \
 //x=10.905 //y=7.4 //x2=10.405 //y2=5.02
cc_1080 ( N_VDD_c_1015_n N_noxref_4_M64_noxref_d ) capacitor c=4.9285e-19 \
 //x=12.95 //y=7.4 //x2=10.405 //y2=5.02
cc_1081 ( N_VDD_M62_noxref_s N_noxref_4_M64_noxref_d ) capacitor c=0.00130656f \
 //x=9.095 //y=5.02 //x2=10.405 //y2=5.02
cc_1082 ( N_VDD_M63_noxref_d N_noxref_4_M64_noxref_d ) capacitor c=0.0664752f \
 //x=9.965 //y=5.02 //x2=10.405 //y2=5.02
cc_1083 ( N_VDD_M65_noxref_d N_noxref_4_M64_noxref_d ) capacitor c=0.0664752f \
 //x=10.845 //y=5.02 //x2=10.405 //y2=5.02
cc_1084 ( N_VDD_c_1035_p N_noxref_4_M66_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=11.285 //y2=5.02
cc_1085 ( N_VDD_c_1083_p N_noxref_4_M66_noxref_d ) capacitor c=0.014035f \
 //x=11.785 //y=7.4 //x2=11.285 //y2=5.02
cc_1086 ( N_VDD_c_1015_n N_noxref_4_M66_noxref_d ) capacitor c=0.00939849f \
 //x=12.95 //y=7.4 //x2=11.285 //y2=5.02
cc_1087 ( N_VDD_M65_noxref_d N_noxref_4_M66_noxref_d ) capacitor c=0.0664752f \
 //x=10.845 //y=5.02 //x2=11.285 //y2=5.02
cc_1088 ( N_VDD_M67_noxref_d N_noxref_4_M66_noxref_d ) capacitor c=0.0664752f \
 //x=11.725 //y=5.02 //x2=11.285 //y2=5.02
cc_1089 ( N_VDD_M68_noxref_s N_noxref_4_M66_noxref_d ) capacitor c=4.52683e-19 \
 //x=13.605 //y=5.02 //x2=11.285 //y2=5.02
cc_1090 ( N_VDD_c_1035_p N_noxref_5_c_2540_n ) capacitor c=0.0316681f \
 //x=84.73 //y=7.4 //x2=7.28 //y2=4.07
cc_1091 ( N_VDD_c_1114_p N_noxref_5_c_2540_n ) capacitor c=0.00168692f \
 //x=3.16 //y=7.4 //x2=7.28 //y2=4.07
cc_1092 ( N_VDD_c_1115_p N_noxref_5_c_2540_n ) capacitor c=0.0027159f \
 //x=4.335 //y=7.4 //x2=7.28 //y2=4.07
cc_1093 ( N_VDD_c_1052_p N_noxref_5_c_2540_n ) capacitor c=0.00113459f \
 //x=5.215 //y=7.4 //x2=7.28 //y2=4.07
cc_1094 ( N_VDD_c_1013_n N_noxref_5_c_2540_n ) capacitor c=0.0274508f //x=3.33 \
 //y=7.4 //x2=7.28 //y2=4.07
cc_1095 ( N_VDD_M55_noxref_d N_noxref_5_c_2540_n ) capacitor c=5.05307e-19 \
 //x=2.405 //y=5.02 //x2=7.28 //y2=4.07
cc_1096 ( N_VDD_M56_noxref_s N_noxref_5_c_2540_n ) capacitor c=0.00122826f \
 //x=4.285 //y=5.02 //x2=7.28 //y2=4.07
cc_1097 ( N_VDD_c_1035_p N_noxref_5_c_2547_n ) capacitor c=0.00181362f \
 //x=84.73 //y=7.4 //x2=1.965 //y2=4.07
cc_1098 ( N_VDD_c_1014_n N_noxref_5_c_2548_n ) capacitor c=0.0140578f //x=8.14 \
 //y=7.4 //x2=17.275 //y2=4.07
cc_1099 ( N_VDD_c_1015_n N_noxref_5_c_2548_n ) capacitor c=0.0140578f \
 //x=12.95 //y=7.4 //x2=17.275 //y2=4.07
cc_1100 ( N_VDD_c_1016_n N_noxref_5_c_2548_n ) capacitor c=0.014632f //x=16.28 \
 //y=7.4 //x2=17.275 //y2=4.07
cc_1101 ( N_VDD_c_1014_n N_noxref_5_c_2551_n ) capacitor c=0.00104411f \
 //x=8.14 //y=7.4 //x2=7.51 //y2=4.07
cc_1102 ( N_VDD_c_1012_n N_noxref_5_c_2525_n ) capacitor c=6.87732e-19 \
 //x=0.74 //y=7.4 //x2=1.85 //y2=2.08
cc_1103 ( N_VDD_c_1013_n N_noxref_5_c_2525_n ) capacitor c=5.66013e-19 \
 //x=3.33 //y=7.4 //x2=1.85 //y2=2.08
cc_1104 ( N_VDD_c_1035_p N_noxref_5_c_2554_n ) capacitor c=0.00449316f \
 //x=84.73 //y=7.4 //x2=5.655 //y2=5.155
cc_1105 ( N_VDD_c_1052_p N_noxref_5_c_2554_n ) capacitor c=4.32228e-19 \
 //x=5.215 //y=7.4 //x2=5.655 //y2=5.155
cc_1106 ( N_VDD_c_1129_p N_noxref_5_c_2554_n ) capacitor c=4.31906e-19 \
 //x=6.095 //y=7.4 //x2=5.655 //y2=5.155
cc_1107 ( N_VDD_M57_noxref_d N_noxref_5_c_2554_n ) capacitor c=0.0115147f \
 //x=5.155 //y=5.02 //x2=5.655 //y2=5.155
cc_1108 ( N_VDD_c_1013_n N_noxref_5_c_2558_n ) capacitor c=0.00863585f \
 //x=3.33 //y=7.4 //x2=4.945 //y2=5.155
cc_1109 ( N_VDD_M56_noxref_s N_noxref_5_c_2558_n ) capacitor c=0.0831083f \
 //x=4.285 //y=5.02 //x2=4.945 //y2=5.155
cc_1110 ( N_VDD_c_1035_p N_noxref_5_c_2560_n ) capacitor c=0.0044221f \
 //x=84.73 //y=7.4 //x2=6.535 //y2=5.155
cc_1111 ( N_VDD_c_1129_p N_noxref_5_c_2560_n ) capacitor c=4.31931e-19 \
 //x=6.095 //y=7.4 //x2=6.535 //y2=5.155
cc_1112 ( N_VDD_c_1135_p N_noxref_5_c_2560_n ) capacitor c=4.31931e-19 \
 //x=6.975 //y=7.4 //x2=6.535 //y2=5.155
cc_1113 ( N_VDD_M59_noxref_d N_noxref_5_c_2560_n ) capacitor c=0.0112985f \
 //x=6.035 //y=5.02 //x2=6.535 //y2=5.155
cc_1114 ( N_VDD_c_1035_p N_noxref_5_c_2564_n ) capacitor c=0.00433242f \
 //x=84.73 //y=7.4 //x2=7.315 //y2=5.155
cc_1115 ( N_VDD_c_1135_p N_noxref_5_c_2564_n ) capacitor c=7.46626e-19 \
 //x=6.975 //y=7.4 //x2=7.315 //y2=5.155
cc_1116 ( N_VDD_c_1139_p N_noxref_5_c_2564_n ) capacitor c=0.00198565f \
 //x=7.97 //y=7.4 //x2=7.315 //y2=5.155
cc_1117 ( N_VDD_M61_noxref_d N_noxref_5_c_2564_n ) capacitor c=0.0112985f \
 //x=6.915 //y=5.02 //x2=7.315 //y2=5.155
cc_1118 ( N_VDD_c_1035_p N_noxref_5_c_2528_n ) capacitor c=0.00125279f \
 //x=84.73 //y=7.4 //x2=17.39 //y2=2.08
cc_1119 ( N_VDD_c_1142_p N_noxref_5_c_2528_n ) capacitor c=2.87256e-19 \
 //x=17.865 //y=7.4 //x2=17.39 //y2=2.08
cc_1120 ( N_VDD_c_1016_n N_noxref_5_c_2528_n ) capacitor c=0.0132802f \
 //x=16.28 //y=7.4 //x2=17.39 //y2=2.08
cc_1121 ( N_VDD_c_1014_n N_noxref_5_c_2571_n ) capacitor c=0.0427201f //x=8.14 \
 //y=7.4 //x2=7.395 //y2=4.07
cc_1122 ( N_VDD_c_1037_p N_noxref_5_M54_noxref_g ) capacitor c=0.00673971f \
 //x=2.465 //y=7.4 //x2=1.89 //y2=6.02
cc_1123 ( N_VDD_M53_noxref_d N_noxref_5_M54_noxref_g ) capacitor c=0.015318f \
 //x=1.525 //y=5.02 //x2=1.89 //y2=6.02
cc_1124 ( N_VDD_c_1037_p N_noxref_5_M55_noxref_g ) capacitor c=0.00672952f \
 //x=2.465 //y=7.4 //x2=2.33 //y2=6.02
cc_1125 ( N_VDD_c_1013_n N_noxref_5_M55_noxref_g ) capacitor c=0.00928743f \
 //x=3.33 //y=7.4 //x2=2.33 //y2=6.02
cc_1126 ( N_VDD_M55_noxref_d N_noxref_5_M55_noxref_g ) capacitor c=0.0430452f \
 //x=2.405 //y=5.02 //x2=2.33 //y2=6.02
cc_1127 ( N_VDD_c_1142_p N_noxref_5_M72_noxref_g ) capacitor c=0.00726866f \
 //x=17.865 //y=7.4 //x2=17.29 //y2=6.02
cc_1128 ( N_VDD_M72_noxref_s N_noxref_5_M72_noxref_g ) capacitor c=0.054195f \
 //x=16.935 //y=5.02 //x2=17.29 //y2=6.02
cc_1129 ( N_VDD_c_1142_p N_noxref_5_M73_noxref_g ) capacitor c=0.00672952f \
 //x=17.865 //y=7.4 //x2=17.73 //y2=6.02
cc_1130 ( N_VDD_M73_noxref_d N_noxref_5_M73_noxref_g ) capacitor c=0.015318f \
 //x=17.805 //y=5.02 //x2=17.73 //y2=6.02
cc_1131 ( N_VDD_c_1016_n N_noxref_5_c_2581_n ) capacitor c=0.0149273f \
 //x=16.28 //y=7.4 //x2=17.39 //y2=4.7
cc_1132 ( N_VDD_c_1035_p N_noxref_5_M56_noxref_d ) capacitor c=0.00285091f \
 //x=84.73 //y=7.4 //x2=4.715 //y2=5.02
cc_1133 ( N_VDD_c_1052_p N_noxref_5_M56_noxref_d ) capacitor c=0.0141016f \
 //x=5.215 //y=7.4 //x2=4.715 //y2=5.02
cc_1134 ( N_VDD_M57_noxref_d N_noxref_5_M56_noxref_d ) capacitor c=0.0664752f \
 //x=5.155 //y=5.02 //x2=4.715 //y2=5.02
cc_1135 ( N_VDD_c_1035_p N_noxref_5_M58_noxref_d ) capacitor c=0.00275186f \
 //x=84.73 //y=7.4 //x2=5.595 //y2=5.02
cc_1136 ( N_VDD_c_1129_p N_noxref_5_M58_noxref_d ) capacitor c=0.0140346f \
 //x=6.095 //y=7.4 //x2=5.595 //y2=5.02
cc_1137 ( N_VDD_c_1014_n N_noxref_5_M58_noxref_d ) capacitor c=4.9285e-19 \
 //x=8.14 //y=7.4 //x2=5.595 //y2=5.02
cc_1138 ( N_VDD_M56_noxref_s N_noxref_5_M58_noxref_d ) capacitor c=0.00130656f \
 //x=4.285 //y=5.02 //x2=5.595 //y2=5.02
cc_1139 ( N_VDD_M57_noxref_d N_noxref_5_M58_noxref_d ) capacitor c=0.0664752f \
 //x=5.155 //y=5.02 //x2=5.595 //y2=5.02
cc_1140 ( N_VDD_M59_noxref_d N_noxref_5_M58_noxref_d ) capacitor c=0.0664752f \
 //x=6.035 //y=5.02 //x2=5.595 //y2=5.02
cc_1141 ( N_VDD_c_1035_p N_noxref_5_M60_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=6.475 //y2=5.02
cc_1142 ( N_VDD_c_1135_p N_noxref_5_M60_noxref_d ) capacitor c=0.014035f \
 //x=6.975 //y=7.4 //x2=6.475 //y2=5.02
cc_1143 ( N_VDD_c_1014_n N_noxref_5_M60_noxref_d ) capacitor c=0.00939849f \
 //x=8.14 //y=7.4 //x2=6.475 //y2=5.02
cc_1144 ( N_VDD_M59_noxref_d N_noxref_5_M60_noxref_d ) capacitor c=0.0664752f \
 //x=6.035 //y=5.02 //x2=6.475 //y2=5.02
cc_1145 ( N_VDD_M61_noxref_d N_noxref_5_M60_noxref_d ) capacitor c=0.0664752f \
 //x=6.915 //y=5.02 //x2=6.475 //y2=5.02
cc_1146 ( N_VDD_M62_noxref_s N_noxref_5_M60_noxref_d ) capacitor c=3.57641e-19 \
 //x=9.095 //y=5.02 //x2=6.475 //y2=5.02
cc_1147 ( N_VDD_c_1017_n N_noxref_6_c_2819_n ) capacitor c=0.014416f //x=19.61 \
 //y=7.4 //x2=20.605 //y2=4.07
cc_1148 ( N_VDD_c_1017_n N_noxref_6_c_2820_n ) capacitor c=5.12647e-19 \
 //x=19.61 //y=7.4 //x2=18.985 //y2=4.07
cc_1149 ( N_VDD_c_1035_p N_noxref_6_c_2821_n ) capacitor c=0.00453663f \
 //x=84.73 //y=7.4 //x2=18.305 //y2=5.2
cc_1150 ( N_VDD_c_1142_p N_noxref_6_c_2821_n ) capacitor c=4.48391e-19 \
 //x=17.865 //y=7.4 //x2=18.305 //y2=5.2
cc_1151 ( N_VDD_c_1174_p N_noxref_6_c_2821_n ) capacitor c=4.48391e-19 \
 //x=18.745 //y=7.4 //x2=18.305 //y2=5.2
cc_1152 ( N_VDD_M73_noxref_d N_noxref_6_c_2821_n ) capacitor c=0.0124542f \
 //x=17.805 //y=5.02 //x2=18.305 //y2=5.2
cc_1153 ( N_VDD_c_1016_n N_noxref_6_c_2825_n ) capacitor c=0.00985474f \
 //x=16.28 //y=7.4 //x2=17.595 //y2=5.2
cc_1154 ( N_VDD_M72_noxref_s N_noxref_6_c_2825_n ) capacitor c=0.087833f \
 //x=16.935 //y=5.02 //x2=17.595 //y2=5.2
cc_1155 ( N_VDD_c_1035_p N_noxref_6_c_2827_n ) capacitor c=0.00301575f \
 //x=84.73 //y=7.4 //x2=18.785 //y2=5.2
cc_1156 ( N_VDD_c_1174_p N_noxref_6_c_2827_n ) capacitor c=7.72068e-19 \
 //x=18.745 //y=7.4 //x2=18.785 //y2=5.2
cc_1157 ( N_VDD_M75_noxref_d N_noxref_6_c_2827_n ) capacitor c=0.0158515f \
 //x=18.685 //y=5.02 //x2=18.785 //y2=5.2
cc_1158 ( N_VDD_c_1016_n N_noxref_6_c_2804_n ) capacitor c=0.00151618f \
 //x=16.28 //y=7.4 //x2=18.87 //y2=4.07
cc_1159 ( N_VDD_c_1017_n N_noxref_6_c_2804_n ) capacitor c=0.0433528f \
 //x=19.61 //y=7.4 //x2=18.87 //y2=4.07
cc_1160 ( N_VDD_c_1035_p N_noxref_6_c_2805_n ) capacitor c=9.10347e-19 \
 //x=84.73 //y=7.4 //x2=20.72 //y2=2.08
cc_1161 ( N_VDD_c_1017_n N_noxref_6_c_2805_n ) capacitor c=0.0134111f \
 //x=19.61 //y=7.4 //x2=20.72 //y2=2.08
cc_1162 ( N_VDD_M76_noxref_s N_noxref_6_c_2805_n ) capacitor c=0.0120327f \
 //x=20.565 //y=5.02 //x2=20.72 //y2=2.08
cc_1163 ( N_VDD_c_1186_p N_noxref_6_M76_noxref_g ) capacitor c=0.00749687f \
 //x=21.495 //y=7.4 //x2=20.92 //y2=6.02
cc_1164 ( N_VDD_M76_noxref_s N_noxref_6_M76_noxref_g ) capacitor c=0.0477201f \
 //x=20.565 //y=5.02 //x2=20.92 //y2=6.02
cc_1165 ( N_VDD_c_1186_p N_noxref_6_M77_noxref_g ) capacitor c=0.00675175f \
 //x=21.495 //y=7.4 //x2=21.36 //y2=6.02
cc_1166 ( N_VDD_M77_noxref_d N_noxref_6_M77_noxref_g ) capacitor c=0.015318f \
 //x=21.435 //y=5.02 //x2=21.36 //y2=6.02
cc_1167 ( N_VDD_c_1017_n N_noxref_6_c_2839_n ) capacitor c=0.0076931f \
 //x=19.61 //y=7.4 //x2=20.995 //y2=4.79
cc_1168 ( N_VDD_M76_noxref_s N_noxref_6_c_2839_n ) capacitor c=0.00444914f \
 //x=20.565 //y=5.02 //x2=20.995 //y2=4.79
cc_1169 ( N_VDD_c_1035_p N_noxref_6_M72_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=17.365 //y2=5.02
cc_1170 ( N_VDD_c_1142_p N_noxref_6_M72_noxref_d ) capacitor c=0.0140317f \
 //x=17.865 //y=7.4 //x2=17.365 //y2=5.02
cc_1171 ( N_VDD_c_1017_n N_noxref_6_M72_noxref_d ) capacitor c=6.94454e-19 \
 //x=19.61 //y=7.4 //x2=17.365 //y2=5.02
cc_1172 ( N_VDD_M73_noxref_d N_noxref_6_M72_noxref_d ) capacitor c=0.0664752f \
 //x=17.805 //y=5.02 //x2=17.365 //y2=5.02
cc_1173 ( N_VDD_c_1035_p N_noxref_6_M74_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=18.245 //y2=5.02
cc_1174 ( N_VDD_c_1174_p N_noxref_6_M74_noxref_d ) capacitor c=0.0140317f \
 //x=18.745 //y=7.4 //x2=18.245 //y2=5.02
cc_1175 ( N_VDD_c_1017_n N_noxref_6_M74_noxref_d ) capacitor c=0.0120541f \
 //x=19.61 //y=7.4 //x2=18.245 //y2=5.02
cc_1176 ( N_VDD_M72_noxref_s N_noxref_6_M74_noxref_d ) capacitor c=0.00111971f \
 //x=16.935 //y=5.02 //x2=18.245 //y2=5.02
cc_1177 ( N_VDD_M73_noxref_d N_noxref_6_M74_noxref_d ) capacitor c=0.0664752f \
 //x=17.805 //y=5.02 //x2=18.245 //y2=5.02
cc_1178 ( N_VDD_M75_noxref_d N_noxref_6_M74_noxref_d ) capacitor c=0.0664752f \
 //x=18.685 //y=5.02 //x2=18.245 //y2=5.02
cc_1179 ( N_VDD_M76_noxref_s N_noxref_6_M74_noxref_d ) capacitor c=3.73257e-19 \
 //x=20.565 //y=5.02 //x2=18.245 //y2=5.02
cc_1180 ( N_VDD_c_1014_n N_noxref_7_c_2955_n ) capacitor c=7.21808e-19 \
 //x=8.14 //y=7.4 //x2=6.66 //y2=2.08
cc_1181 ( N_VDD_c_1015_n N_noxref_7_c_2956_n ) capacitor c=6.21611e-19 \
 //x=12.95 //y=7.4 //x2=11.47 //y2=2.08
cc_1182 ( N_VDD_c_1035_p N_noxref_7_c_2965_n ) capacitor c=0.00453473f \
 //x=84.73 //y=7.4 //x2=14.975 //y2=5.2
cc_1183 ( N_VDD_c_1091_p N_noxref_7_c_2965_n ) capacitor c=4.48391e-19 \
 //x=14.535 //y=7.4 //x2=14.975 //y2=5.2
cc_1184 ( N_VDD_c_1207_p N_noxref_7_c_2965_n ) capacitor c=4.48377e-19 \
 //x=15.415 //y=7.4 //x2=14.975 //y2=5.2
cc_1185 ( N_VDD_M69_noxref_d N_noxref_7_c_2965_n ) capacitor c=0.0124506f \
 //x=14.475 //y=5.02 //x2=14.975 //y2=5.2
cc_1186 ( N_VDD_c_1015_n N_noxref_7_c_2969_n ) capacitor c=0.00985474f \
 //x=12.95 //y=7.4 //x2=14.265 //y2=5.2
cc_1187 ( N_VDD_M68_noxref_s N_noxref_7_c_2969_n ) capacitor c=0.087833f \
 //x=13.605 //y=5.02 //x2=14.265 //y2=5.2
cc_1188 ( N_VDD_c_1035_p N_noxref_7_c_2971_n ) capacitor c=0.00301575f \
 //x=84.73 //y=7.4 //x2=15.455 //y2=5.2
cc_1189 ( N_VDD_c_1207_p N_noxref_7_c_2971_n ) capacitor c=7.72068e-19 \
 //x=15.415 //y=7.4 //x2=15.455 //y2=5.2
cc_1190 ( N_VDD_M71_noxref_d N_noxref_7_c_2971_n ) capacitor c=0.0158515f \
 //x=15.355 //y=5.02 //x2=15.455 //y2=5.2
cc_1191 ( N_VDD_M72_noxref_s N_noxref_7_c_2971_n ) capacitor c=2.44532e-19 \
 //x=16.935 //y=5.02 //x2=15.455 //y2=5.2
cc_1192 ( N_VDD_c_1015_n N_noxref_7_c_2958_n ) capacitor c=0.00151618f \
 //x=12.95 //y=7.4 //x2=15.54 //y2=3.7
cc_1193 ( N_VDD_c_1016_n N_noxref_7_c_2958_n ) capacitor c=0.0427716f \
 //x=16.28 //y=7.4 //x2=15.54 //y2=3.7
cc_1194 ( N_VDD_c_1018_n N_noxref_7_c_2959_n ) capacitor c=7.28883e-19 \
 //x=24.42 //y=7.4 //x2=22.94 //y2=2.08
cc_1195 ( N_VDD_c_1135_p N_noxref_7_M60_noxref_g ) capacitor c=0.00675175f \
 //x=6.975 //y=7.4 //x2=6.4 //y2=6.02
cc_1196 ( N_VDD_M59_noxref_d N_noxref_7_M60_noxref_g ) capacitor c=0.015318f \
 //x=6.035 //y=5.02 //x2=6.4 //y2=6.02
cc_1197 ( N_VDD_c_1135_p N_noxref_7_M61_noxref_g ) capacitor c=0.00675379f \
 //x=6.975 //y=7.4 //x2=6.84 //y2=6.02
cc_1198 ( N_VDD_M61_noxref_d N_noxref_7_M61_noxref_g ) capacitor c=0.0394719f \
 //x=6.915 //y=5.02 //x2=6.84 //y2=6.02
cc_1199 ( N_VDD_c_1083_p N_noxref_7_M66_noxref_g ) capacitor c=0.00675175f \
 //x=11.785 //y=7.4 //x2=11.21 //y2=6.02
cc_1200 ( N_VDD_M65_noxref_d N_noxref_7_M66_noxref_g ) capacitor c=0.015318f \
 //x=10.845 //y=5.02 //x2=11.21 //y2=6.02
cc_1201 ( N_VDD_c_1083_p N_noxref_7_M67_noxref_g ) capacitor c=0.00675379f \
 //x=11.785 //y=7.4 //x2=11.65 //y2=6.02
cc_1202 ( N_VDD_M67_noxref_d N_noxref_7_M67_noxref_g ) capacitor c=0.0394719f \
 //x=11.725 //y=5.02 //x2=11.65 //y2=6.02
cc_1203 ( N_VDD_c_1226_p N_noxref_7_M80_noxref_g ) capacitor c=0.00675175f \
 //x=23.255 //y=7.4 //x2=22.68 //y2=6.02
cc_1204 ( N_VDD_M79_noxref_d N_noxref_7_M80_noxref_g ) capacitor c=0.015318f \
 //x=22.315 //y=5.02 //x2=22.68 //y2=6.02
cc_1205 ( N_VDD_c_1226_p N_noxref_7_M81_noxref_g ) capacitor c=0.00675379f \
 //x=23.255 //y=7.4 //x2=23.12 //y2=6.02
cc_1206 ( N_VDD_M81_noxref_d N_noxref_7_M81_noxref_g ) capacitor c=0.0394719f \
 //x=23.195 //y=5.02 //x2=23.12 //y2=6.02
cc_1207 ( N_VDD_c_1035_p N_noxref_7_M68_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=14.035 //y2=5.02
cc_1208 ( N_VDD_c_1091_p N_noxref_7_M68_noxref_d ) capacitor c=0.0140317f \
 //x=14.535 //y=7.4 //x2=14.035 //y2=5.02
cc_1209 ( N_VDD_c_1016_n N_noxref_7_M68_noxref_d ) capacitor c=6.94454e-19 \
 //x=16.28 //y=7.4 //x2=14.035 //y2=5.02
cc_1210 ( N_VDD_M69_noxref_d N_noxref_7_M68_noxref_d ) capacitor c=0.0664752f \
 //x=14.475 //y=5.02 //x2=14.035 //y2=5.02
cc_1211 ( N_VDD_c_1035_p N_noxref_7_M70_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=14.915 //y2=5.02
cc_1212 ( N_VDD_c_1207_p N_noxref_7_M70_noxref_d ) capacitor c=0.0140317f \
 //x=15.415 //y=7.4 //x2=14.915 //y2=5.02
cc_1213 ( N_VDD_c_1016_n N_noxref_7_M70_noxref_d ) capacitor c=0.0120541f \
 //x=16.28 //y=7.4 //x2=14.915 //y2=5.02
cc_1214 ( N_VDD_M68_noxref_s N_noxref_7_M70_noxref_d ) capacitor c=0.00111971f \
 //x=13.605 //y=5.02 //x2=14.915 //y2=5.02
cc_1215 ( N_VDD_M69_noxref_d N_noxref_7_M70_noxref_d ) capacitor c=0.0664752f \
 //x=14.475 //y=5.02 //x2=14.915 //y2=5.02
cc_1216 ( N_VDD_M71_noxref_d N_noxref_7_M70_noxref_d ) capacitor c=0.0664752f \
 //x=15.355 //y=5.02 //x2=14.915 //y2=5.02
cc_1217 ( N_VDD_M72_noxref_s N_noxref_7_M70_noxref_d ) capacitor c=4.54516e-19 \
 //x=16.935 //y=5.02 //x2=14.915 //y2=5.02
cc_1218 ( N_VDD_c_1035_p N_noxref_8_c_3309_n ) capacitor c=0.00453663f \
 //x=84.73 //y=7.4 //x2=26.445 //y2=5.2
cc_1219 ( N_VDD_c_1242_p N_noxref_8_c_3309_n ) capacitor c=4.48391e-19 \
 //x=26.005 //y=7.4 //x2=26.445 //y2=5.2
cc_1220 ( N_VDD_c_1243_p N_noxref_8_c_3309_n ) capacitor c=4.48391e-19 \
 //x=26.885 //y=7.4 //x2=26.445 //y2=5.2
cc_1221 ( N_VDD_M83_noxref_d N_noxref_8_c_3309_n ) capacitor c=0.0124542f \
 //x=25.945 //y=5.02 //x2=26.445 //y2=5.2
cc_1222 ( N_VDD_c_1018_n N_noxref_8_c_3313_n ) capacitor c=0.00985474f \
 //x=24.42 //y=7.4 //x2=25.735 //y2=5.2
cc_1223 ( N_VDD_M82_noxref_s N_noxref_8_c_3313_n ) capacitor c=0.087833f \
 //x=25.075 //y=5.02 //x2=25.735 //y2=5.2
cc_1224 ( N_VDD_c_1035_p N_noxref_8_c_3315_n ) capacitor c=0.00301575f \
 //x=84.73 //y=7.4 //x2=26.925 //y2=5.2
cc_1225 ( N_VDD_c_1243_p N_noxref_8_c_3315_n ) capacitor c=7.72068e-19 \
 //x=26.885 //y=7.4 //x2=26.925 //y2=5.2
cc_1226 ( N_VDD_M85_noxref_d N_noxref_8_c_3315_n ) capacitor c=0.0158515f \
 //x=26.825 //y=5.02 //x2=26.925 //y2=5.2
cc_1227 ( N_VDD_c_1018_n N_noxref_8_c_3282_n ) capacitor c=0.00151618f \
 //x=24.42 //y=7.4 //x2=27.01 //y2=2.59
cc_1228 ( N_VDD_c_1019_n N_noxref_8_c_3282_n ) capacitor c=0.0428942f \
 //x=27.75 //y=7.4 //x2=27.01 //y2=2.59
cc_1229 ( N_VDD_c_1035_p N_noxref_8_c_3284_n ) capacitor c=9.10347e-19 \
 //x=84.73 //y=7.4 //x2=28.86 //y2=2.08
cc_1230 ( N_VDD_c_1019_n N_noxref_8_c_3284_n ) capacitor c=0.0133749f \
 //x=27.75 //y=7.4 //x2=28.86 //y2=2.08
cc_1231 ( N_VDD_M86_noxref_s N_noxref_8_c_3284_n ) capacitor c=0.0125322f \
 //x=28.705 //y=5.02 //x2=28.86 //y2=2.08
cc_1232 ( N_VDD_c_1035_p N_noxref_8_c_3285_n ) capacitor c=9.10347e-19 \
 //x=84.73 //y=7.4 //x2=33.67 //y2=2.08
cc_1233 ( N_VDD_c_1020_n N_noxref_8_c_3285_n ) capacitor c=0.013427f //x=32.56 \
 //y=7.4 //x2=33.67 //y2=2.08
cc_1234 ( N_VDD_M92_noxref_s N_noxref_8_c_3285_n ) capacitor c=0.0126798f \
 //x=33.515 //y=5.02 //x2=33.67 //y2=2.08
cc_1235 ( N_VDD_c_1258_p N_noxref_8_M86_noxref_g ) capacitor c=0.00749687f \
 //x=29.635 //y=7.4 //x2=29.06 //y2=6.02
cc_1236 ( N_VDD_M86_noxref_s N_noxref_8_M86_noxref_g ) capacitor c=0.0477201f \
 //x=28.705 //y=5.02 //x2=29.06 //y2=6.02
cc_1237 ( N_VDD_c_1258_p N_noxref_8_M87_noxref_g ) capacitor c=0.00675175f \
 //x=29.635 //y=7.4 //x2=29.5 //y2=6.02
cc_1238 ( N_VDD_M87_noxref_d N_noxref_8_M87_noxref_g ) capacitor c=0.015318f \
 //x=29.575 //y=5.02 //x2=29.5 //y2=6.02
cc_1239 ( N_VDD_c_1262_p N_noxref_8_M92_noxref_g ) capacitor c=0.00749687f \
 //x=34.445 //y=7.4 //x2=33.87 //y2=6.02
cc_1240 ( N_VDD_M92_noxref_s N_noxref_8_M92_noxref_g ) capacitor c=0.0477201f \
 //x=33.515 //y=5.02 //x2=33.87 //y2=6.02
cc_1241 ( N_VDD_c_1262_p N_noxref_8_M93_noxref_g ) capacitor c=0.00675175f \
 //x=34.445 //y=7.4 //x2=34.31 //y2=6.02
cc_1242 ( N_VDD_M93_noxref_d N_noxref_8_M93_noxref_g ) capacitor c=0.015318f \
 //x=34.385 //y=5.02 //x2=34.31 //y2=6.02
cc_1243 ( N_VDD_c_1019_n N_noxref_8_c_3334_n ) capacitor c=0.00757682f \
 //x=27.75 //y=7.4 //x2=29.135 //y2=4.79
cc_1244 ( N_VDD_M86_noxref_s N_noxref_8_c_3334_n ) capacitor c=0.00444914f \
 //x=28.705 //y=5.02 //x2=29.135 //y2=4.79
cc_1245 ( N_VDD_c_1020_n N_noxref_8_c_3336_n ) capacitor c=0.00757682f \
 //x=32.56 //y=7.4 //x2=33.945 //y2=4.79
cc_1246 ( N_VDD_M92_noxref_s N_noxref_8_c_3336_n ) capacitor c=0.00444914f \
 //x=33.515 //y=5.02 //x2=33.945 //y2=4.79
cc_1247 ( N_VDD_c_1035_p N_noxref_8_M82_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=25.505 //y2=5.02
cc_1248 ( N_VDD_c_1242_p N_noxref_8_M82_noxref_d ) capacitor c=0.0140317f \
 //x=26.005 //y=7.4 //x2=25.505 //y2=5.02
cc_1249 ( N_VDD_c_1019_n N_noxref_8_M82_noxref_d ) capacitor c=6.94454e-19 \
 //x=27.75 //y=7.4 //x2=25.505 //y2=5.02
cc_1250 ( N_VDD_M83_noxref_d N_noxref_8_M82_noxref_d ) capacitor c=0.0664752f \
 //x=25.945 //y=5.02 //x2=25.505 //y2=5.02
cc_1251 ( N_VDD_c_1035_p N_noxref_8_M84_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=26.385 //y2=5.02
cc_1252 ( N_VDD_c_1243_p N_noxref_8_M84_noxref_d ) capacitor c=0.0140317f \
 //x=26.885 //y=7.4 //x2=26.385 //y2=5.02
cc_1253 ( N_VDD_c_1019_n N_noxref_8_M84_noxref_d ) capacitor c=0.0120541f \
 //x=27.75 //y=7.4 //x2=26.385 //y2=5.02
cc_1254 ( N_VDD_M82_noxref_s N_noxref_8_M84_noxref_d ) capacitor c=0.00111971f \
 //x=25.075 //y=5.02 //x2=26.385 //y2=5.02
cc_1255 ( N_VDD_M83_noxref_d N_noxref_8_M84_noxref_d ) capacitor c=0.0664752f \
 //x=25.945 //y=5.02 //x2=26.385 //y2=5.02
cc_1256 ( N_VDD_M85_noxref_d N_noxref_8_M84_noxref_d ) capacitor c=0.0664752f \
 //x=26.825 //y=5.02 //x2=26.385 //y2=5.02
cc_1257 ( N_VDD_M86_noxref_s N_noxref_8_M84_noxref_d ) capacitor c=3.73257e-19 \
 //x=28.705 //y=5.02 //x2=26.385 //y2=5.02
cc_1258 ( N_VDD_c_1035_p N_noxref_9_c_3525_n ) capacitor c=0.00444892f \
 //x=84.73 //y=7.4 //x2=34.885 //y2=5.155
cc_1259 ( N_VDD_c_1262_p N_noxref_9_c_3525_n ) capacitor c=4.31931e-19 \
 //x=34.445 //y=7.4 //x2=34.885 //y2=5.155
cc_1260 ( N_VDD_c_1283_p N_noxref_9_c_3525_n ) capacitor c=4.31931e-19 \
 //x=35.325 //y=7.4 //x2=34.885 //y2=5.155
cc_1261 ( N_VDD_M93_noxref_d N_noxref_9_c_3525_n ) capacitor c=0.0112985f \
 //x=34.385 //y=5.02 //x2=34.885 //y2=5.155
cc_1262 ( N_VDD_c_1020_n N_noxref_9_c_3529_n ) capacitor c=0.00863585f \
 //x=32.56 //y=7.4 //x2=34.175 //y2=5.155
cc_1263 ( N_VDD_M92_noxref_s N_noxref_9_c_3529_n ) capacitor c=0.0831083f \
 //x=33.515 //y=5.02 //x2=34.175 //y2=5.155
cc_1264 ( N_VDD_c_1035_p N_noxref_9_c_3531_n ) capacitor c=0.0044221f \
 //x=84.73 //y=7.4 //x2=35.765 //y2=5.155
cc_1265 ( N_VDD_c_1283_p N_noxref_9_c_3531_n ) capacitor c=4.31931e-19 \
 //x=35.325 //y=7.4 //x2=35.765 //y2=5.155
cc_1266 ( N_VDD_c_1289_p N_noxref_9_c_3531_n ) capacitor c=4.31931e-19 \
 //x=36.205 //y=7.4 //x2=35.765 //y2=5.155
cc_1267 ( N_VDD_M95_noxref_d N_noxref_9_c_3531_n ) capacitor c=0.0112985f \
 //x=35.265 //y=5.02 //x2=35.765 //y2=5.155
cc_1268 ( N_VDD_c_1035_p N_noxref_9_c_3535_n ) capacitor c=0.00434174f \
 //x=84.73 //y=7.4 //x2=36.545 //y2=5.155
cc_1269 ( N_VDD_c_1289_p N_noxref_9_c_3535_n ) capacitor c=7.46626e-19 \
 //x=36.205 //y=7.4 //x2=36.545 //y2=5.155
cc_1270 ( N_VDD_c_1293_p N_noxref_9_c_3535_n ) capacitor c=0.00198565f \
 //x=37.2 //y=7.4 //x2=36.545 //y2=5.155
cc_1271 ( N_VDD_M97_noxref_d N_noxref_9_c_3535_n ) capacitor c=0.0112985f \
 //x=36.145 //y=5.02 //x2=36.545 //y2=5.155
cc_1272 ( N_VDD_c_1021_n N_noxref_9_c_3512_n ) capacitor c=0.042636f //x=37.37 \
 //y=7.4 //x2=36.63 //y2=2.59
cc_1273 ( N_VDD_c_1035_p N_noxref_9_c_3513_n ) capacitor c=0.00125279f \
 //x=84.73 //y=7.4 //x2=38.48 //y2=2.08
cc_1274 ( N_VDD_c_1297_p N_noxref_9_c_3513_n ) capacitor c=2.87256e-19 \
 //x=38.955 //y=7.4 //x2=38.48 //y2=2.08
cc_1275 ( N_VDD_c_1021_n N_noxref_9_c_3513_n ) capacitor c=0.0133961f \
 //x=37.37 //y=7.4 //x2=38.48 //y2=2.08
cc_1276 ( N_VDD_c_1297_p N_noxref_9_M98_noxref_g ) capacitor c=0.00726866f \
 //x=38.955 //y=7.4 //x2=38.38 //y2=6.02
cc_1277 ( N_VDD_M98_noxref_s N_noxref_9_M98_noxref_g ) capacitor c=0.054195f \
 //x=38.025 //y=5.02 //x2=38.38 //y2=6.02
cc_1278 ( N_VDD_c_1297_p N_noxref_9_M99_noxref_g ) capacitor c=0.00672952f \
 //x=38.955 //y=7.4 //x2=38.82 //y2=6.02
cc_1279 ( N_VDD_M99_noxref_d N_noxref_9_M99_noxref_g ) capacitor c=0.015318f \
 //x=38.895 //y=5.02 //x2=38.82 //y2=6.02
cc_1280 ( N_VDD_c_1021_n N_noxref_9_c_3547_n ) capacitor c=0.015293f //x=37.37 \
 //y=7.4 //x2=38.48 //y2=4.7
cc_1281 ( N_VDD_c_1035_p N_noxref_9_M92_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=33.945 //y2=5.02
cc_1282 ( N_VDD_c_1262_p N_noxref_9_M92_noxref_d ) capacitor c=0.014035f \
 //x=34.445 //y=7.4 //x2=33.945 //y2=5.02
cc_1283 ( N_VDD_M93_noxref_d N_noxref_9_M92_noxref_d ) capacitor c=0.0664752f \
 //x=34.385 //y=5.02 //x2=33.945 //y2=5.02
cc_1284 ( N_VDD_c_1035_p N_noxref_9_M94_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=34.825 //y2=5.02
cc_1285 ( N_VDD_c_1283_p N_noxref_9_M94_noxref_d ) capacitor c=0.014035f \
 //x=35.325 //y=7.4 //x2=34.825 //y2=5.02
cc_1286 ( N_VDD_c_1021_n N_noxref_9_M94_noxref_d ) capacitor c=4.9285e-19 \
 //x=37.37 //y=7.4 //x2=34.825 //y2=5.02
cc_1287 ( N_VDD_M92_noxref_s N_noxref_9_M94_noxref_d ) capacitor c=0.00130656f \
 //x=33.515 //y=5.02 //x2=34.825 //y2=5.02
cc_1288 ( N_VDD_M93_noxref_d N_noxref_9_M94_noxref_d ) capacitor c=0.0664752f \
 //x=34.385 //y=5.02 //x2=34.825 //y2=5.02
cc_1289 ( N_VDD_M95_noxref_d N_noxref_9_M94_noxref_d ) capacitor c=0.0664752f \
 //x=35.265 //y=5.02 //x2=34.825 //y2=5.02
cc_1290 ( N_VDD_c_1035_p N_noxref_9_M96_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=35.705 //y2=5.02
cc_1291 ( N_VDD_c_1289_p N_noxref_9_M96_noxref_d ) capacitor c=0.014035f \
 //x=36.205 //y=7.4 //x2=35.705 //y2=5.02
cc_1292 ( N_VDD_c_1021_n N_noxref_9_M96_noxref_d ) capacitor c=0.00939849f \
 //x=37.37 //y=7.4 //x2=35.705 //y2=5.02
cc_1293 ( N_VDD_M95_noxref_d N_noxref_9_M96_noxref_d ) capacitor c=0.0664752f \
 //x=35.265 //y=5.02 //x2=35.705 //y2=5.02
cc_1294 ( N_VDD_M97_noxref_d N_noxref_9_M96_noxref_d ) capacitor c=0.0664752f \
 //x=36.145 //y=5.02 //x2=35.705 //y2=5.02
cc_1295 ( N_VDD_M98_noxref_s N_noxref_9_M96_noxref_d ) capacitor c=4.52683e-19 \
 //x=38.025 //y=5.02 //x2=35.705 //y2=5.02
cc_1296 ( N_VDD_c_1019_n N_noxref_10_c_3690_n ) capacitor c=0.0143396f \
 //x=27.75 //y=7.4 //x2=31.7 //y2=4.07
cc_1297 ( N_VDD_c_1020_n N_noxref_10_c_3691_n ) capacitor c=0.0140578f \
 //x=32.56 //y=7.4 //x2=41.695 //y2=4.07
cc_1298 ( N_VDD_c_1021_n N_noxref_10_c_3691_n ) capacitor c=0.0140578f \
 //x=37.37 //y=7.4 //x2=41.695 //y2=4.07
cc_1299 ( N_VDD_c_1022_n N_noxref_10_c_3691_n ) capacitor c=0.014632f //x=40.7 \
 //y=7.4 //x2=41.695 //y2=4.07
cc_1300 ( N_VDD_c_1020_n N_noxref_10_c_3694_n ) capacitor c=0.00104411f \
 //x=32.56 //y=7.4 //x2=31.93 //y2=4.07
cc_1301 ( N_VDD_c_1018_n N_noxref_10_c_3675_n ) capacitor c=5.18578e-19 \
 //x=24.42 //y=7.4 //x2=26.27 //y2=2.08
cc_1302 ( N_VDD_c_1019_n N_noxref_10_c_3675_n ) capacitor c=3.21957e-19 \
 //x=27.75 //y=7.4 //x2=26.27 //y2=2.08
cc_1303 ( N_VDD_c_1035_p N_noxref_10_c_3697_n ) capacitor c=0.00444751f \
 //x=84.73 //y=7.4 //x2=30.075 //y2=5.155
cc_1304 ( N_VDD_c_1258_p N_noxref_10_c_3697_n ) capacitor c=4.31931e-19 \
 //x=29.635 //y=7.4 //x2=30.075 //y2=5.155
cc_1305 ( N_VDD_c_1328_p N_noxref_10_c_3697_n ) capacitor c=4.31906e-19 \
 //x=30.515 //y=7.4 //x2=30.075 //y2=5.155
cc_1306 ( N_VDD_M87_noxref_d N_noxref_10_c_3697_n ) capacitor c=0.0112985f \
 //x=29.575 //y=5.02 //x2=30.075 //y2=5.155
cc_1307 ( N_VDD_c_1019_n N_noxref_10_c_3701_n ) capacitor c=0.00863585f \
 //x=27.75 //y=7.4 //x2=29.365 //y2=5.155
cc_1308 ( N_VDD_M86_noxref_s N_noxref_10_c_3701_n ) capacitor c=0.0831083f \
 //x=28.705 //y=5.02 //x2=29.365 //y2=5.155
cc_1309 ( N_VDD_c_1035_p N_noxref_10_c_3703_n ) capacitor c=0.0044221f \
 //x=84.73 //y=7.4 //x2=30.955 //y2=5.155
cc_1310 ( N_VDD_c_1328_p N_noxref_10_c_3703_n ) capacitor c=4.31931e-19 \
 //x=30.515 //y=7.4 //x2=30.955 //y2=5.155
cc_1311 ( N_VDD_c_1334_p N_noxref_10_c_3703_n ) capacitor c=4.31931e-19 \
 //x=31.395 //y=7.4 //x2=30.955 //y2=5.155
cc_1312 ( N_VDD_M89_noxref_d N_noxref_10_c_3703_n ) capacitor c=0.0112985f \
 //x=30.455 //y=5.02 //x2=30.955 //y2=5.155
cc_1313 ( N_VDD_c_1035_p N_noxref_10_c_3707_n ) capacitor c=0.00433242f \
 //x=84.73 //y=7.4 //x2=31.735 //y2=5.155
cc_1314 ( N_VDD_c_1334_p N_noxref_10_c_3707_n ) capacitor c=7.46626e-19 \
 //x=31.395 //y=7.4 //x2=31.735 //y2=5.155
cc_1315 ( N_VDD_c_1338_p N_noxref_10_c_3707_n ) capacitor c=0.00198565f \
 //x=32.39 //y=7.4 //x2=31.735 //y2=5.155
cc_1316 ( N_VDD_M91_noxref_d N_noxref_10_c_3707_n ) capacitor c=0.0112985f \
 //x=31.335 //y=5.02 //x2=31.735 //y2=5.155
cc_1317 ( N_VDD_c_1035_p N_noxref_10_c_3678_n ) capacitor c=0.00125279f \
 //x=84.73 //y=7.4 //x2=41.81 //y2=2.08
cc_1318 ( N_VDD_c_1341_p N_noxref_10_c_3678_n ) capacitor c=2.87256e-19 \
 //x=42.285 //y=7.4 //x2=41.81 //y2=2.08
cc_1319 ( N_VDD_c_1022_n N_noxref_10_c_3678_n ) capacitor c=0.0132802f \
 //x=40.7 //y=7.4 //x2=41.81 //y2=2.08
cc_1320 ( N_VDD_c_1020_n N_noxref_10_c_3714_n ) capacitor c=0.0427201f \
 //x=32.56 //y=7.4 //x2=31.815 //y2=4.07
cc_1321 ( N_VDD_c_1243_p N_noxref_10_M84_noxref_g ) capacitor c=0.00673971f \
 //x=26.885 //y=7.4 //x2=26.31 //y2=6.02
cc_1322 ( N_VDD_M83_noxref_d N_noxref_10_M84_noxref_g ) capacitor c=0.015318f \
 //x=25.945 //y=5.02 //x2=26.31 //y2=6.02
cc_1323 ( N_VDD_c_1243_p N_noxref_10_M85_noxref_g ) capacitor c=0.00672952f \
 //x=26.885 //y=7.4 //x2=26.75 //y2=6.02
cc_1324 ( N_VDD_c_1019_n N_noxref_10_M85_noxref_g ) capacitor c=0.00928743f \
 //x=27.75 //y=7.4 //x2=26.75 //y2=6.02
cc_1325 ( N_VDD_M85_noxref_d N_noxref_10_M85_noxref_g ) capacitor c=0.0430452f \
 //x=26.825 //y=5.02 //x2=26.75 //y2=6.02
cc_1326 ( N_VDD_c_1341_p N_noxref_10_M102_noxref_g ) capacitor c=0.00726866f \
 //x=42.285 //y=7.4 //x2=41.71 //y2=6.02
cc_1327 ( N_VDD_M102_noxref_s N_noxref_10_M102_noxref_g ) capacitor \
 c=0.054195f //x=41.355 //y=5.02 //x2=41.71 //y2=6.02
cc_1328 ( N_VDD_c_1341_p N_noxref_10_M103_noxref_g ) capacitor c=0.00672952f \
 //x=42.285 //y=7.4 //x2=42.15 //y2=6.02
cc_1329 ( N_VDD_M103_noxref_d N_noxref_10_M103_noxref_g ) capacitor \
 c=0.015318f //x=42.225 //y=5.02 //x2=42.15 //y2=6.02
cc_1330 ( N_VDD_c_1022_n N_noxref_10_c_3724_n ) capacitor c=0.0149273f \
 //x=40.7 //y=7.4 //x2=41.81 //y2=4.7
cc_1331 ( N_VDD_c_1035_p N_noxref_10_M86_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=29.135 //y2=5.02
cc_1332 ( N_VDD_c_1258_p N_noxref_10_M86_noxref_d ) capacitor c=0.014035f \
 //x=29.635 //y=7.4 //x2=29.135 //y2=5.02
cc_1333 ( N_VDD_M87_noxref_d N_noxref_10_M86_noxref_d ) capacitor c=0.0664752f \
 //x=29.575 //y=5.02 //x2=29.135 //y2=5.02
cc_1334 ( N_VDD_c_1035_p N_noxref_10_M88_noxref_d ) capacitor c=0.00275186f \
 //x=84.73 //y=7.4 //x2=30.015 //y2=5.02
cc_1335 ( N_VDD_c_1328_p N_noxref_10_M88_noxref_d ) capacitor c=0.0140346f \
 //x=30.515 //y=7.4 //x2=30.015 //y2=5.02
cc_1336 ( N_VDD_c_1020_n N_noxref_10_M88_noxref_d ) capacitor c=4.9285e-19 \
 //x=32.56 //y=7.4 //x2=30.015 //y2=5.02
cc_1337 ( N_VDD_M86_noxref_s N_noxref_10_M88_noxref_d ) capacitor \
 c=0.00130656f //x=28.705 //y=5.02 //x2=30.015 //y2=5.02
cc_1338 ( N_VDD_M87_noxref_d N_noxref_10_M88_noxref_d ) capacitor c=0.0664752f \
 //x=29.575 //y=5.02 //x2=30.015 //y2=5.02
cc_1339 ( N_VDD_M89_noxref_d N_noxref_10_M88_noxref_d ) capacitor c=0.0664752f \
 //x=30.455 //y=5.02 //x2=30.015 //y2=5.02
cc_1340 ( N_VDD_c_1035_p N_noxref_10_M90_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=30.895 //y2=5.02
cc_1341 ( N_VDD_c_1334_p N_noxref_10_M90_noxref_d ) capacitor c=0.014035f \
 //x=31.395 //y=7.4 //x2=30.895 //y2=5.02
cc_1342 ( N_VDD_c_1020_n N_noxref_10_M90_noxref_d ) capacitor c=0.00939849f \
 //x=32.56 //y=7.4 //x2=30.895 //y2=5.02
cc_1343 ( N_VDD_M89_noxref_d N_noxref_10_M90_noxref_d ) capacitor c=0.0664752f \
 //x=30.455 //y=5.02 //x2=30.895 //y2=5.02
cc_1344 ( N_VDD_M91_noxref_d N_noxref_10_M90_noxref_d ) capacitor c=0.0664752f \
 //x=31.335 //y=5.02 //x2=30.895 //y2=5.02
cc_1345 ( N_VDD_M92_noxref_s N_noxref_10_M90_noxref_d ) capacitor \
 c=3.57641e-19 //x=33.515 //y=5.02 //x2=30.895 //y2=5.02
cc_1346 ( N_VDD_c_1035_p N_noxref_11_c_3975_n ) capacitor c=0.00453663f \
 //x=84.73 //y=7.4 //x2=42.725 //y2=5.2
cc_1347 ( N_VDD_c_1341_p N_noxref_11_c_3975_n ) capacitor c=4.48391e-19 \
 //x=42.285 //y=7.4 //x2=42.725 //y2=5.2
cc_1348 ( N_VDD_c_1371_p N_noxref_11_c_3975_n ) capacitor c=4.48391e-19 \
 //x=43.165 //y=7.4 //x2=42.725 //y2=5.2
cc_1349 ( N_VDD_M103_noxref_d N_noxref_11_c_3975_n ) capacitor c=0.0124542f \
 //x=42.225 //y=5.02 //x2=42.725 //y2=5.2
cc_1350 ( N_VDD_c_1022_n N_noxref_11_c_3979_n ) capacitor c=0.00985474f \
 //x=40.7 //y=7.4 //x2=42.015 //y2=5.2
cc_1351 ( N_VDD_M102_noxref_s N_noxref_11_c_3979_n ) capacitor c=0.087833f \
 //x=41.355 //y=5.02 //x2=42.015 //y2=5.2
cc_1352 ( N_VDD_c_1035_p N_noxref_11_c_3981_n ) capacitor c=0.00301575f \
 //x=84.73 //y=7.4 //x2=43.205 //y2=5.2
cc_1353 ( N_VDD_c_1371_p N_noxref_11_c_3981_n ) capacitor c=7.72068e-19 \
 //x=43.165 //y=7.4 //x2=43.205 //y2=5.2
cc_1354 ( N_VDD_M105_noxref_d N_noxref_11_c_3981_n ) capacitor c=0.0158515f \
 //x=43.105 //y=5.02 //x2=43.205 //y2=5.2
cc_1355 ( N_VDD_c_1022_n N_noxref_11_c_3959_n ) capacitor c=0.00151618f \
 //x=40.7 //y=7.4 //x2=43.29 //y2=2.59
cc_1356 ( N_VDD_c_1023_n N_noxref_11_c_3959_n ) capacitor c=0.0429885f \
 //x=44.03 //y=7.4 //x2=43.29 //y2=2.59
cc_1357 ( N_VDD_c_1035_p N_noxref_11_c_3961_n ) capacitor c=9.10347e-19 \
 //x=84.73 //y=7.4 //x2=45.14 //y2=2.08
cc_1358 ( N_VDD_c_1023_n N_noxref_11_c_3961_n ) capacitor c=0.0134348f \
 //x=44.03 //y=7.4 //x2=45.14 //y2=2.08
cc_1359 ( N_VDD_M106_noxref_s N_noxref_11_c_3961_n ) capacitor c=0.0126798f \
 //x=44.985 //y=5.02 //x2=45.14 //y2=2.08
cc_1360 ( N_VDD_c_1383_p N_noxref_11_M106_noxref_g ) capacitor c=0.00749687f \
 //x=45.915 //y=7.4 //x2=45.34 //y2=6.02
cc_1361 ( N_VDD_M106_noxref_s N_noxref_11_M106_noxref_g ) capacitor \
 c=0.0477201f //x=44.985 //y=5.02 //x2=45.34 //y2=6.02
cc_1362 ( N_VDD_c_1383_p N_noxref_11_M107_noxref_g ) capacitor c=0.00675175f \
 //x=45.915 //y=7.4 //x2=45.78 //y2=6.02
cc_1363 ( N_VDD_M107_noxref_d N_noxref_11_M107_noxref_g ) capacitor \
 c=0.015318f //x=45.855 //y=5.02 //x2=45.78 //y2=6.02
cc_1364 ( N_VDD_c_1023_n N_noxref_11_c_3993_n ) capacitor c=0.0076931f \
 //x=44.03 //y=7.4 //x2=45.415 //y2=4.79
cc_1365 ( N_VDD_M106_noxref_s N_noxref_11_c_3993_n ) capacitor c=0.00444914f \
 //x=44.985 //y=5.02 //x2=45.415 //y2=4.79
cc_1366 ( N_VDD_c_1035_p N_noxref_11_M102_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=41.785 //y2=5.02
cc_1367 ( N_VDD_c_1341_p N_noxref_11_M102_noxref_d ) capacitor c=0.0140317f \
 //x=42.285 //y=7.4 //x2=41.785 //y2=5.02
cc_1368 ( N_VDD_c_1023_n N_noxref_11_M102_noxref_d ) capacitor c=6.94454e-19 \
 //x=44.03 //y=7.4 //x2=41.785 //y2=5.02
cc_1369 ( N_VDD_M103_noxref_d N_noxref_11_M102_noxref_d ) capacitor \
 c=0.0664752f //x=42.225 //y=5.02 //x2=41.785 //y2=5.02
cc_1370 ( N_VDD_c_1035_p N_noxref_11_M104_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=42.665 //y2=5.02
cc_1371 ( N_VDD_c_1371_p N_noxref_11_M104_noxref_d ) capacitor c=0.0140317f \
 //x=43.165 //y=7.4 //x2=42.665 //y2=5.02
cc_1372 ( N_VDD_c_1023_n N_noxref_11_M104_noxref_d ) capacitor c=0.0120541f \
 //x=44.03 //y=7.4 //x2=42.665 //y2=5.02
cc_1373 ( N_VDD_M102_noxref_s N_noxref_11_M104_noxref_d ) capacitor \
 c=0.00111971f //x=41.355 //y=5.02 //x2=42.665 //y2=5.02
cc_1374 ( N_VDD_M103_noxref_d N_noxref_11_M104_noxref_d ) capacitor \
 c=0.0664752f //x=42.225 //y=5.02 //x2=42.665 //y2=5.02
cc_1375 ( N_VDD_M105_noxref_d N_noxref_11_M104_noxref_d ) capacitor \
 c=0.0664752f //x=43.105 //y=5.02 //x2=42.665 //y2=5.02
cc_1376 ( N_VDD_M106_noxref_s N_noxref_11_M104_noxref_d ) capacitor \
 c=3.73257e-19 //x=44.985 //y=5.02 //x2=42.665 //y2=5.02
cc_1377 ( N_VDD_c_1020_n N_noxref_12_c_4111_n ) capacitor c=7.21808e-19 \
 //x=32.56 //y=7.4 //x2=31.08 //y2=2.08
cc_1378 ( N_VDD_c_1021_n N_noxref_12_c_4112_n ) capacitor c=6.21611e-19 \
 //x=37.37 //y=7.4 //x2=35.89 //y2=2.08
cc_1379 ( N_VDD_c_1035_p N_noxref_12_c_4121_n ) capacitor c=0.00453473f \
 //x=84.73 //y=7.4 //x2=39.395 //y2=5.2
cc_1380 ( N_VDD_c_1297_p N_noxref_12_c_4121_n ) capacitor c=4.48391e-19 \
 //x=38.955 //y=7.4 //x2=39.395 //y2=5.2
cc_1381 ( N_VDD_c_1404_p N_noxref_12_c_4121_n ) capacitor c=4.48377e-19 \
 //x=39.835 //y=7.4 //x2=39.395 //y2=5.2
cc_1382 ( N_VDD_M99_noxref_d N_noxref_12_c_4121_n ) capacitor c=0.0124506f \
 //x=38.895 //y=5.02 //x2=39.395 //y2=5.2
cc_1383 ( N_VDD_c_1021_n N_noxref_12_c_4125_n ) capacitor c=0.00985474f \
 //x=37.37 //y=7.4 //x2=38.685 //y2=5.2
cc_1384 ( N_VDD_M98_noxref_s N_noxref_12_c_4125_n ) capacitor c=0.087833f \
 //x=38.025 //y=5.02 //x2=38.685 //y2=5.2
cc_1385 ( N_VDD_c_1035_p N_noxref_12_c_4127_n ) capacitor c=0.00301575f \
 //x=84.73 //y=7.4 //x2=39.875 //y2=5.2
cc_1386 ( N_VDD_c_1404_p N_noxref_12_c_4127_n ) capacitor c=7.72068e-19 \
 //x=39.835 //y=7.4 //x2=39.875 //y2=5.2
cc_1387 ( N_VDD_M101_noxref_d N_noxref_12_c_4127_n ) capacitor c=0.0158515f \
 //x=39.775 //y=5.02 //x2=39.875 //y2=5.2
cc_1388 ( N_VDD_M102_noxref_s N_noxref_12_c_4127_n ) capacitor c=2.44532e-19 \
 //x=41.355 //y=5.02 //x2=39.875 //y2=5.2
cc_1389 ( N_VDD_c_1021_n N_noxref_12_c_4114_n ) capacitor c=0.00151618f \
 //x=37.37 //y=7.4 //x2=39.96 //y2=3.7
cc_1390 ( N_VDD_c_1022_n N_noxref_12_c_4114_n ) capacitor c=0.0427716f \
 //x=40.7 //y=7.4 //x2=39.96 //y2=3.7
cc_1391 ( N_VDD_c_1024_n N_noxref_12_c_4115_n ) capacitor c=7.21739e-19 \
 //x=48.84 //y=7.4 //x2=47.36 //y2=2.08
cc_1392 ( N_VDD_c_1334_p N_noxref_12_M90_noxref_g ) capacitor c=0.00675175f \
 //x=31.395 //y=7.4 //x2=30.82 //y2=6.02
cc_1393 ( N_VDD_M89_noxref_d N_noxref_12_M90_noxref_g ) capacitor c=0.015318f \
 //x=30.455 //y=5.02 //x2=30.82 //y2=6.02
cc_1394 ( N_VDD_c_1334_p N_noxref_12_M91_noxref_g ) capacitor c=0.00675379f \
 //x=31.395 //y=7.4 //x2=31.26 //y2=6.02
cc_1395 ( N_VDD_M91_noxref_d N_noxref_12_M91_noxref_g ) capacitor c=0.0394719f \
 //x=31.335 //y=5.02 //x2=31.26 //y2=6.02
cc_1396 ( N_VDD_c_1289_p N_noxref_12_M96_noxref_g ) capacitor c=0.00675175f \
 //x=36.205 //y=7.4 //x2=35.63 //y2=6.02
cc_1397 ( N_VDD_M95_noxref_d N_noxref_12_M96_noxref_g ) capacitor c=0.015318f \
 //x=35.265 //y=5.02 //x2=35.63 //y2=6.02
cc_1398 ( N_VDD_c_1289_p N_noxref_12_M97_noxref_g ) capacitor c=0.00675379f \
 //x=36.205 //y=7.4 //x2=36.07 //y2=6.02
cc_1399 ( N_VDD_M97_noxref_d N_noxref_12_M97_noxref_g ) capacitor c=0.0394719f \
 //x=36.145 //y=5.02 //x2=36.07 //y2=6.02
cc_1400 ( N_VDD_c_1423_p N_noxref_12_M110_noxref_g ) capacitor c=0.00675175f \
 //x=47.675 //y=7.4 //x2=47.1 //y2=6.02
cc_1401 ( N_VDD_M109_noxref_d N_noxref_12_M110_noxref_g ) capacitor \
 c=0.015318f //x=46.735 //y=5.02 //x2=47.1 //y2=6.02
cc_1402 ( N_VDD_c_1423_p N_noxref_12_M111_noxref_g ) capacitor c=0.00675379f \
 //x=47.675 //y=7.4 //x2=47.54 //y2=6.02
cc_1403 ( N_VDD_M111_noxref_d N_noxref_12_M111_noxref_g ) capacitor \
 c=0.0394719f //x=47.615 //y=5.02 //x2=47.54 //y2=6.02
cc_1404 ( N_VDD_c_1035_p N_noxref_12_M98_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=38.455 //y2=5.02
cc_1405 ( N_VDD_c_1297_p N_noxref_12_M98_noxref_d ) capacitor c=0.0140317f \
 //x=38.955 //y=7.4 //x2=38.455 //y2=5.02
cc_1406 ( N_VDD_c_1022_n N_noxref_12_M98_noxref_d ) capacitor c=6.94454e-19 \
 //x=40.7 //y=7.4 //x2=38.455 //y2=5.02
cc_1407 ( N_VDD_M99_noxref_d N_noxref_12_M98_noxref_d ) capacitor c=0.0664752f \
 //x=38.895 //y=5.02 //x2=38.455 //y2=5.02
cc_1408 ( N_VDD_c_1035_p N_noxref_12_M100_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=39.335 //y2=5.02
cc_1409 ( N_VDD_c_1404_p N_noxref_12_M100_noxref_d ) capacitor c=0.0140317f \
 //x=39.835 //y=7.4 //x2=39.335 //y2=5.02
cc_1410 ( N_VDD_c_1022_n N_noxref_12_M100_noxref_d ) capacitor c=0.0120541f \
 //x=40.7 //y=7.4 //x2=39.335 //y2=5.02
cc_1411 ( N_VDD_M98_noxref_s N_noxref_12_M100_noxref_d ) capacitor \
 c=0.00111971f //x=38.025 //y=5.02 //x2=39.335 //y2=5.02
cc_1412 ( N_VDD_M99_noxref_d N_noxref_12_M100_noxref_d ) capacitor \
 c=0.0664752f //x=38.895 //y=5.02 //x2=39.335 //y2=5.02
cc_1413 ( N_VDD_M101_noxref_d N_noxref_12_M100_noxref_d ) capacitor \
 c=0.0664752f //x=39.775 //y=5.02 //x2=39.335 //y2=5.02
cc_1414 ( N_VDD_M102_noxref_s N_noxref_12_M100_noxref_d ) capacitor \
 c=4.54516e-19 //x=41.355 //y=5.02 //x2=39.335 //y2=5.02
cc_1415 ( N_VDD_c_1023_n N_noxref_13_c_4455_n ) capacitor c=0.0140578f \
 //x=44.03 //y=7.4 //x2=47.985 //y2=4.07
cc_1416 ( N_VDD_c_1024_n N_noxref_13_c_4455_n ) capacitor c=0.00168281f \
 //x=48.84 //y=7.4 //x2=47.985 //y2=4.07
cc_1417 ( N_VDD_c_1035_p N_noxref_13_c_4444_n ) capacitor c=0.0151699f \
 //x=84.73 //y=7.4 //x2=81.655 //y2=4.07
cc_1418 ( N_VDD_c_1441_p N_noxref_13_c_4444_n ) capacitor c=4.075e-19 \
 //x=83.08 //y=7.4 //x2=81.655 //y2=4.07
cc_1419 ( N_VDD_c_1031_n N_noxref_13_c_4444_n ) capacitor c=0.014826f \
 //x=76.59 //y=7.4 //x2=81.655 //y2=4.07
cc_1420 ( N_VDD_c_1032_n N_noxref_13_c_4444_n ) capacitor c=0.0225025f \
 //x=79.92 //y=7.4 //x2=81.655 //y2=4.07
cc_1421 ( N_VDD_c_1031_n N_noxref_13_c_4461_n ) capacitor c=5.4458e-19 \
 //x=76.59 //y=7.4 //x2=75.225 //y2=4.07
cc_1422 ( N_VDD_c_1022_n N_noxref_13_c_4445_n ) capacitor c=5.02639e-19 \
 //x=40.7 //y=7.4 //x2=42.55 //y2=2.08
cc_1423 ( N_VDD_c_1023_n N_noxref_13_c_4445_n ) capacitor c=3.21957e-19 \
 //x=44.03 //y=7.4 //x2=42.55 //y2=2.08
cc_1424 ( N_VDD_c_1035_p N_noxref_13_c_4464_n ) capacitor c=0.00444892f \
 //x=84.73 //y=7.4 //x2=46.355 //y2=5.155
cc_1425 ( N_VDD_c_1383_p N_noxref_13_c_4464_n ) capacitor c=4.31931e-19 \
 //x=45.915 //y=7.4 //x2=46.355 //y2=5.155
cc_1426 ( N_VDD_c_1449_p N_noxref_13_c_4464_n ) capacitor c=4.31931e-19 \
 //x=46.795 //y=7.4 //x2=46.355 //y2=5.155
cc_1427 ( N_VDD_M107_noxref_d N_noxref_13_c_4464_n ) capacitor c=0.0112985f \
 //x=45.855 //y=5.02 //x2=46.355 //y2=5.155
cc_1428 ( N_VDD_c_1023_n N_noxref_13_c_4468_n ) capacitor c=0.00863585f \
 //x=44.03 //y=7.4 //x2=45.645 //y2=5.155
cc_1429 ( N_VDD_M106_noxref_s N_noxref_13_c_4468_n ) capacitor c=0.0831083f \
 //x=44.985 //y=5.02 //x2=45.645 //y2=5.155
cc_1430 ( N_VDD_c_1035_p N_noxref_13_c_4470_n ) capacitor c=0.0044221f \
 //x=84.73 //y=7.4 //x2=47.235 //y2=5.155
cc_1431 ( N_VDD_c_1449_p N_noxref_13_c_4470_n ) capacitor c=4.31931e-19 \
 //x=46.795 //y=7.4 //x2=47.235 //y2=5.155
cc_1432 ( N_VDD_c_1423_p N_noxref_13_c_4470_n ) capacitor c=4.31931e-19 \
 //x=47.675 //y=7.4 //x2=47.235 //y2=5.155
cc_1433 ( N_VDD_M109_noxref_d N_noxref_13_c_4470_n ) capacitor c=0.0112985f \
 //x=46.735 //y=5.02 //x2=47.235 //y2=5.155
cc_1434 ( N_VDD_c_1035_p N_noxref_13_c_4474_n ) capacitor c=0.00434174f \
 //x=84.73 //y=7.4 //x2=48.015 //y2=5.155
cc_1435 ( N_VDD_c_1423_p N_noxref_13_c_4474_n ) capacitor c=7.46626e-19 \
 //x=47.675 //y=7.4 //x2=48.015 //y2=5.155
cc_1436 ( N_VDD_c_1459_p N_noxref_13_c_4474_n ) capacitor c=0.00198565f \
 //x=48.67 //y=7.4 //x2=48.015 //y2=5.155
cc_1437 ( N_VDD_M111_noxref_d N_noxref_13_c_4474_n ) capacitor c=0.0112985f \
 //x=47.615 //y=5.02 //x2=48.015 //y2=5.155
cc_1438 ( N_VDD_c_1024_n N_noxref_13_c_4448_n ) capacitor c=0.0433404f \
 //x=48.84 //y=7.4 //x2=48.1 //y2=2.59
cc_1439 ( N_VDD_c_1031_n N_noxref_13_c_4479_n ) capacitor c=0.00491684f \
 //x=76.59 //y=7.4 //x2=75.11 //y2=4.54
cc_1440 ( N_VDD_c_1030_n N_noxref_13_c_4449_n ) capacitor c=8.10235e-19 \
 //x=73.26 //y=7.4 //x2=75.11 //y2=2.08
cc_1441 ( N_VDD_c_1031_n N_noxref_13_c_4449_n ) capacitor c=0.0042566f \
 //x=76.59 //y=7.4 //x2=75.11 //y2=2.08
cc_1442 ( N_VDD_c_1032_n N_noxref_13_c_4451_n ) capacitor c=0.00116377f \
 //x=79.92 //y=7.4 //x2=81.77 //y2=2.08
cc_1443 ( N_VDD_c_1033_n N_noxref_13_c_4451_n ) capacitor c=5.67082e-19 \
 //x=83.25 //y=7.4 //x2=81.77 //y2=2.08
cc_1444 ( N_VDD_c_1371_p N_noxref_13_M104_noxref_g ) capacitor c=0.00673971f \
 //x=43.165 //y=7.4 //x2=42.59 //y2=6.02
cc_1445 ( N_VDD_M103_noxref_d N_noxref_13_M104_noxref_g ) capacitor \
 c=0.015318f //x=42.225 //y=5.02 //x2=42.59 //y2=6.02
cc_1446 ( N_VDD_c_1371_p N_noxref_13_M105_noxref_g ) capacitor c=0.00672952f \
 //x=43.165 //y=7.4 //x2=43.03 //y2=6.02
cc_1447 ( N_VDD_c_1023_n N_noxref_13_M105_noxref_g ) capacitor c=0.00928743f \
 //x=44.03 //y=7.4 //x2=43.03 //y2=6.02
cc_1448 ( N_VDD_M105_noxref_d N_noxref_13_M105_noxref_g ) capacitor \
 c=0.0430452f //x=43.105 //y=5.02 //x2=43.03 //y2=6.02
cc_1449 ( N_VDD_c_1472_p N_noxref_13_M144_noxref_g ) capacitor c=0.0067918f \
 //x=75.725 //y=7.4 //x2=75.15 //y2=6.025
cc_1450 ( N_VDD_M143_noxref_d N_noxref_13_M144_noxref_g ) capacitor \
 c=0.015526f //x=74.785 //y=5.025 //x2=75.15 //y2=6.025
cc_1451 ( N_VDD_c_1472_p N_noxref_13_M145_noxref_g ) capacitor c=0.00754867f \
 //x=75.725 //y=7.4 //x2=75.59 //y2=6.025
cc_1452 ( N_VDD_M145_noxref_d N_noxref_13_M145_noxref_g ) capacitor \
 c=0.0537676f //x=75.665 //y=5.025 //x2=75.59 //y2=6.025
cc_1453 ( N_VDD_c_1441_p N_noxref_13_M152_noxref_g ) capacitor c=0.00513565f \
 //x=83.08 //y=7.4 //x2=81.81 //y2=6.025
cc_1454 ( N_VDD_c_1441_p N_noxref_13_M153_noxref_g ) capacitor c=0.00512552f \
 //x=83.08 //y=7.4 //x2=82.25 //y2=6.025
cc_1455 ( N_VDD_c_1033_n N_noxref_13_M153_noxref_g ) capacitor c=0.0113524f \
 //x=83.25 //y=7.4 //x2=82.25 //y2=6.025
cc_1456 ( N_VDD_c_1031_n N_noxref_13_c_4496_n ) capacitor c=0.00985898f \
 //x=76.59 //y=7.4 //x2=75.515 //y2=4.795
cc_1457 ( N_VDD_c_1031_n N_noxref_13_c_4497_n ) capacitor c=2.76772e-19 \
 //x=76.59 //y=7.4 //x2=75.15 //y2=4.705
cc_1458 ( N_VDD_c_1035_p N_noxref_13_M106_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=45.415 //y2=5.02
cc_1459 ( N_VDD_c_1383_p N_noxref_13_M106_noxref_d ) capacitor c=0.014035f \
 //x=45.915 //y=7.4 //x2=45.415 //y2=5.02
cc_1460 ( N_VDD_M107_noxref_d N_noxref_13_M106_noxref_d ) capacitor \
 c=0.0664752f //x=45.855 //y=5.02 //x2=45.415 //y2=5.02
cc_1461 ( N_VDD_c_1035_p N_noxref_13_M108_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=46.295 //y2=5.02
cc_1462 ( N_VDD_c_1449_p N_noxref_13_M108_noxref_d ) capacitor c=0.014035f \
 //x=46.795 //y=7.4 //x2=46.295 //y2=5.02
cc_1463 ( N_VDD_c_1024_n N_noxref_13_M108_noxref_d ) capacitor c=4.9285e-19 \
 //x=48.84 //y=7.4 //x2=46.295 //y2=5.02
cc_1464 ( N_VDD_M106_noxref_s N_noxref_13_M108_noxref_d ) capacitor \
 c=0.00130656f //x=44.985 //y=5.02 //x2=46.295 //y2=5.02
cc_1465 ( N_VDD_M107_noxref_d N_noxref_13_M108_noxref_d ) capacitor \
 c=0.0664752f //x=45.855 //y=5.02 //x2=46.295 //y2=5.02
cc_1466 ( N_VDD_M109_noxref_d N_noxref_13_M108_noxref_d ) capacitor \
 c=0.0664752f //x=46.735 //y=5.02 //x2=46.295 //y2=5.02
cc_1467 ( N_VDD_c_1035_p N_noxref_13_M110_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=47.175 //y2=5.02
cc_1468 ( N_VDD_c_1423_p N_noxref_13_M110_noxref_d ) capacitor c=0.014035f \
 //x=47.675 //y=7.4 //x2=47.175 //y2=5.02
cc_1469 ( N_VDD_c_1024_n N_noxref_13_M110_noxref_d ) capacitor c=0.00939849f \
 //x=48.84 //y=7.4 //x2=47.175 //y2=5.02
cc_1470 ( N_VDD_M109_noxref_d N_noxref_13_M110_noxref_d ) capacitor \
 c=0.0664752f //x=46.735 //y=5.02 //x2=47.175 //y2=5.02
cc_1471 ( N_VDD_M111_noxref_d N_noxref_13_M110_noxref_d ) capacitor \
 c=0.0664752f //x=47.615 //y=5.02 //x2=47.175 //y2=5.02
cc_1472 ( N_VDD_M112_noxref_s N_noxref_13_M110_noxref_d ) capacitor \
 c=4.52683e-19 //x=49.495 //y=5.02 //x2=47.175 //y2=5.02
cc_1473 ( N_VDD_c_1035_p N_D_c_4900_n ) capacitor c=0.00593968f //x=84.73 \
 //y=7.4 //x2=25.415 //y2=2.96
cc_1474 ( N_VDD_c_1035_p N_D_c_4908_n ) capacitor c=0.00134996f //x=84.73 \
 //y=7.4 //x2=1.225 //y2=2.96
cc_1475 ( N_VDD_c_1035_p N_D_c_4915_n ) capacitor c=0.00128597f //x=84.73 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_1476 ( N_VDD_c_1036_p N_D_c_4915_n ) capacitor c=2.63811e-19 //x=1.585 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_1477 ( N_VDD_c_1012_n N_D_c_4915_n ) capacitor c=0.01673f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_1478 ( N_VDD_c_1035_p N_D_c_4916_n ) capacitor c=0.00125279f //x=84.73 \
 //y=7.4 //x2=25.53 //y2=2.08
cc_1479 ( N_VDD_c_1242_p N_D_c_4916_n ) capacitor c=2.87256e-19 //x=26.005 \
 //y=7.4 //x2=25.53 //y2=2.08
cc_1480 ( N_VDD_c_1018_n N_D_c_4916_n ) capacitor c=0.0140375f //x=24.42 \
 //y=7.4 //x2=25.53 //y2=2.08
cc_1481 ( N_VDD_c_1035_p N_D_c_4917_n ) capacitor c=0.00125279f //x=84.73 \
 //y=7.4 //x2=49.95 //y2=2.08
cc_1482 ( N_VDD_c_1505_p N_D_c_4917_n ) capacitor c=2.87256e-19 //x=50.425 \
 //y=7.4 //x2=49.95 //y2=2.08
cc_1483 ( N_VDD_c_1024_n N_D_c_4917_n ) capacitor c=0.0139262f //x=48.84 \
 //y=7.4 //x2=49.95 //y2=2.08
cc_1484 ( N_VDD_c_1036_p N_D_M52_noxref_g ) capacitor c=0.00726866f //x=1.585 \
 //y=7.4 //x2=1.01 //y2=6.02
cc_1485 ( N_VDD_M52_noxref_s N_D_M52_noxref_g ) capacitor c=0.054195f \
 //x=0.655 //y=5.02 //x2=1.01 //y2=6.02
cc_1486 ( N_VDD_c_1036_p N_D_M53_noxref_g ) capacitor c=0.00672952f //x=1.585 \
 //y=7.4 //x2=1.45 //y2=6.02
cc_1487 ( N_VDD_M53_noxref_d N_D_M53_noxref_g ) capacitor c=0.015318f \
 //x=1.525 //y=5.02 //x2=1.45 //y2=6.02
cc_1488 ( N_VDD_c_1242_p N_D_M82_noxref_g ) capacitor c=0.00726866f //x=26.005 \
 //y=7.4 //x2=25.43 //y2=6.02
cc_1489 ( N_VDD_M82_noxref_s N_D_M82_noxref_g ) capacitor c=0.054195f \
 //x=25.075 //y=5.02 //x2=25.43 //y2=6.02
cc_1490 ( N_VDD_c_1242_p N_D_M83_noxref_g ) capacitor c=0.00672952f //x=26.005 \
 //y=7.4 //x2=25.87 //y2=6.02
cc_1491 ( N_VDD_M83_noxref_d N_D_M83_noxref_g ) capacitor c=0.015318f \
 //x=25.945 //y=5.02 //x2=25.87 //y2=6.02
cc_1492 ( N_VDD_c_1505_p N_D_M112_noxref_g ) capacitor c=0.00726866f \
 //x=50.425 //y=7.4 //x2=49.85 //y2=6.02
cc_1493 ( N_VDD_M112_noxref_s N_D_M112_noxref_g ) capacitor c=0.054195f \
 //x=49.495 //y=5.02 //x2=49.85 //y2=6.02
cc_1494 ( N_VDD_c_1505_p N_D_M113_noxref_g ) capacitor c=0.00672952f \
 //x=50.425 //y=7.4 //x2=50.29 //y2=6.02
cc_1495 ( N_VDD_M113_noxref_d N_D_M113_noxref_g ) capacitor c=0.015318f \
 //x=50.365 //y=5.02 //x2=50.29 //y2=6.02
cc_1496 ( N_VDD_c_1012_n N_D_c_4971_n ) capacitor c=0.0292267f //x=0.74 \
 //y=7.4 //x2=1.11 //y2=4.7
cc_1497 ( N_VDD_c_1018_n N_D_c_4972_n ) capacitor c=0.0154093f //x=24.42 \
 //y=7.4 //x2=25.53 //y2=4.7
cc_1498 ( N_VDD_c_1024_n N_D_c_4973_n ) capacitor c=0.0154093f //x=48.84 \
 //y=7.4 //x2=49.95 //y2=4.7
cc_1499 ( N_VDD_c_1035_p N_noxref_15_c_5253_n ) capacitor c=0.00453663f \
 //x=84.73 //y=7.4 //x2=50.865 //y2=5.2
cc_1500 ( N_VDD_c_1505_p N_noxref_15_c_5253_n ) capacitor c=4.48391e-19 \
 //x=50.425 //y=7.4 //x2=50.865 //y2=5.2
cc_1501 ( N_VDD_c_1524_p N_noxref_15_c_5253_n ) capacitor c=4.48391e-19 \
 //x=51.305 //y=7.4 //x2=50.865 //y2=5.2
cc_1502 ( N_VDD_M113_noxref_d N_noxref_15_c_5253_n ) capacitor c=0.0124542f \
 //x=50.365 //y=5.02 //x2=50.865 //y2=5.2
cc_1503 ( N_VDD_c_1024_n N_noxref_15_c_5257_n ) capacitor c=0.00985474f \
 //x=48.84 //y=7.4 //x2=50.155 //y2=5.2
cc_1504 ( N_VDD_M112_noxref_s N_noxref_15_c_5257_n ) capacitor c=0.087833f \
 //x=49.495 //y=5.02 //x2=50.155 //y2=5.2
cc_1505 ( N_VDD_c_1035_p N_noxref_15_c_5259_n ) capacitor c=0.00301575f \
 //x=84.73 //y=7.4 //x2=51.345 //y2=5.2
cc_1506 ( N_VDD_c_1524_p N_noxref_15_c_5259_n ) capacitor c=7.72068e-19 \
 //x=51.305 //y=7.4 //x2=51.345 //y2=5.2
cc_1507 ( N_VDD_M115_noxref_d N_noxref_15_c_5259_n ) capacitor c=0.0158515f \
 //x=51.245 //y=5.02 //x2=51.345 //y2=5.2
cc_1508 ( N_VDD_c_1024_n N_noxref_15_c_5226_n ) capacitor c=0.00151618f \
 //x=48.84 //y=7.4 //x2=51.43 //y2=2.59
cc_1509 ( N_VDD_c_1025_n N_noxref_15_c_5226_n ) capacitor c=0.0428942f \
 //x=52.17 //y=7.4 //x2=51.43 //y2=2.59
cc_1510 ( N_VDD_c_1035_p N_noxref_15_c_5228_n ) capacitor c=9.10347e-19 \
 //x=84.73 //y=7.4 //x2=53.28 //y2=2.08
cc_1511 ( N_VDD_c_1025_n N_noxref_15_c_5228_n ) capacitor c=0.0133749f \
 //x=52.17 //y=7.4 //x2=53.28 //y2=2.08
cc_1512 ( N_VDD_M116_noxref_s N_noxref_15_c_5228_n ) capacitor c=0.0125322f \
 //x=53.125 //y=5.02 //x2=53.28 //y2=2.08
cc_1513 ( N_VDD_c_1035_p N_noxref_15_c_5229_n ) capacitor c=9.10347e-19 \
 //x=84.73 //y=7.4 //x2=58.09 //y2=2.08
cc_1514 ( N_VDD_c_1026_n N_noxref_15_c_5229_n ) capacitor c=0.013427f \
 //x=56.98 //y=7.4 //x2=58.09 //y2=2.08
cc_1515 ( N_VDD_M122_noxref_s N_noxref_15_c_5229_n ) capacitor c=0.0126798f \
 //x=57.935 //y=5.02 //x2=58.09 //y2=2.08
cc_1516 ( N_VDD_c_1539_p N_noxref_15_M116_noxref_g ) capacitor c=0.00749687f \
 //x=54.055 //y=7.4 //x2=53.48 //y2=6.02
cc_1517 ( N_VDD_M116_noxref_s N_noxref_15_M116_noxref_g ) capacitor \
 c=0.0477201f //x=53.125 //y=5.02 //x2=53.48 //y2=6.02
cc_1518 ( N_VDD_c_1539_p N_noxref_15_M117_noxref_g ) capacitor c=0.00675175f \
 //x=54.055 //y=7.4 //x2=53.92 //y2=6.02
cc_1519 ( N_VDD_M117_noxref_d N_noxref_15_M117_noxref_g ) capacitor \
 c=0.015318f //x=53.995 //y=5.02 //x2=53.92 //y2=6.02
cc_1520 ( N_VDD_c_1543_p N_noxref_15_M122_noxref_g ) capacitor c=0.00749687f \
 //x=58.865 //y=7.4 //x2=58.29 //y2=6.02
cc_1521 ( N_VDD_M122_noxref_s N_noxref_15_M122_noxref_g ) capacitor \
 c=0.0477201f //x=57.935 //y=5.02 //x2=58.29 //y2=6.02
cc_1522 ( N_VDD_c_1543_p N_noxref_15_M123_noxref_g ) capacitor c=0.00675175f \
 //x=58.865 //y=7.4 //x2=58.73 //y2=6.02
cc_1523 ( N_VDD_M123_noxref_d N_noxref_15_M123_noxref_g ) capacitor \
 c=0.015318f //x=58.805 //y=5.02 //x2=58.73 //y2=6.02
cc_1524 ( N_VDD_c_1025_n N_noxref_15_c_5278_n ) capacitor c=0.00757682f \
 //x=52.17 //y=7.4 //x2=53.555 //y2=4.79
cc_1525 ( N_VDD_M116_noxref_s N_noxref_15_c_5278_n ) capacitor c=0.00444914f \
 //x=53.125 //y=5.02 //x2=53.555 //y2=4.79
cc_1526 ( N_VDD_c_1026_n N_noxref_15_c_5280_n ) capacitor c=0.00757682f \
 //x=56.98 //y=7.4 //x2=58.365 //y2=4.79
cc_1527 ( N_VDD_M122_noxref_s N_noxref_15_c_5280_n ) capacitor c=0.00444914f \
 //x=57.935 //y=5.02 //x2=58.365 //y2=4.79
cc_1528 ( N_VDD_c_1035_p N_noxref_15_M112_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=49.925 //y2=5.02
cc_1529 ( N_VDD_c_1505_p N_noxref_15_M112_noxref_d ) capacitor c=0.0140317f \
 //x=50.425 //y=7.4 //x2=49.925 //y2=5.02
cc_1530 ( N_VDD_c_1025_n N_noxref_15_M112_noxref_d ) capacitor c=6.94454e-19 \
 //x=52.17 //y=7.4 //x2=49.925 //y2=5.02
cc_1531 ( N_VDD_M113_noxref_d N_noxref_15_M112_noxref_d ) capacitor \
 c=0.0664752f //x=50.365 //y=5.02 //x2=49.925 //y2=5.02
cc_1532 ( N_VDD_c_1035_p N_noxref_15_M114_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=50.805 //y2=5.02
cc_1533 ( N_VDD_c_1524_p N_noxref_15_M114_noxref_d ) capacitor c=0.0140317f \
 //x=51.305 //y=7.4 //x2=50.805 //y2=5.02
cc_1534 ( N_VDD_c_1025_n N_noxref_15_M114_noxref_d ) capacitor c=0.0120541f \
 //x=52.17 //y=7.4 //x2=50.805 //y2=5.02
cc_1535 ( N_VDD_M112_noxref_s N_noxref_15_M114_noxref_d ) capacitor \
 c=0.00111971f //x=49.495 //y=5.02 //x2=50.805 //y2=5.02
cc_1536 ( N_VDD_M113_noxref_d N_noxref_15_M114_noxref_d ) capacitor \
 c=0.0664752f //x=50.365 //y=5.02 //x2=50.805 //y2=5.02
cc_1537 ( N_VDD_M115_noxref_d N_noxref_15_M114_noxref_d ) capacitor \
 c=0.0664752f //x=51.245 //y=5.02 //x2=50.805 //y2=5.02
cc_1538 ( N_VDD_M116_noxref_s N_noxref_15_M114_noxref_d ) capacitor \
 c=3.73257e-19 //x=53.125 //y=5.02 //x2=50.805 //y2=5.02
cc_1539 ( N_VDD_c_1035_p N_noxref_16_c_5474_n ) capacitor c=0.00444892f \
 //x=84.73 //y=7.4 //x2=59.305 //y2=5.155
cc_1540 ( N_VDD_c_1543_p N_noxref_16_c_5474_n ) capacitor c=4.31931e-19 \
 //x=58.865 //y=7.4 //x2=59.305 //y2=5.155
cc_1541 ( N_VDD_c_1564_p N_noxref_16_c_5474_n ) capacitor c=4.31931e-19 \
 //x=59.745 //y=7.4 //x2=59.305 //y2=5.155
cc_1542 ( N_VDD_M123_noxref_d N_noxref_16_c_5474_n ) capacitor c=0.0112985f \
 //x=58.805 //y=5.02 //x2=59.305 //y2=5.155
cc_1543 ( N_VDD_c_1026_n N_noxref_16_c_5478_n ) capacitor c=0.00863585f \
 //x=56.98 //y=7.4 //x2=58.595 //y2=5.155
cc_1544 ( N_VDD_M122_noxref_s N_noxref_16_c_5478_n ) capacitor c=0.0831083f \
 //x=57.935 //y=5.02 //x2=58.595 //y2=5.155
cc_1545 ( N_VDD_c_1035_p N_noxref_16_c_5480_n ) capacitor c=0.0044221f \
 //x=84.73 //y=7.4 //x2=60.185 //y2=5.155
cc_1546 ( N_VDD_c_1564_p N_noxref_16_c_5480_n ) capacitor c=4.31931e-19 \
 //x=59.745 //y=7.4 //x2=60.185 //y2=5.155
cc_1547 ( N_VDD_c_1570_p N_noxref_16_c_5480_n ) capacitor c=4.31931e-19 \
 //x=60.625 //y=7.4 //x2=60.185 //y2=5.155
cc_1548 ( N_VDD_M125_noxref_d N_noxref_16_c_5480_n ) capacitor c=0.0112985f \
 //x=59.685 //y=5.02 //x2=60.185 //y2=5.155
cc_1549 ( N_VDD_c_1035_p N_noxref_16_c_5484_n ) capacitor c=0.00434174f \
 //x=84.73 //y=7.4 //x2=60.965 //y2=5.155
cc_1550 ( N_VDD_c_1570_p N_noxref_16_c_5484_n ) capacitor c=7.46626e-19 \
 //x=60.625 //y=7.4 //x2=60.965 //y2=5.155
cc_1551 ( N_VDD_c_1574_p N_noxref_16_c_5484_n ) capacitor c=0.00198565f \
 //x=61.62 //y=7.4 //x2=60.965 //y2=5.155
cc_1552 ( N_VDD_M127_noxref_d N_noxref_16_c_5484_n ) capacitor c=0.0112985f \
 //x=60.565 //y=5.02 //x2=60.965 //y2=5.155
cc_1553 ( N_VDD_c_1027_n N_noxref_16_c_5461_n ) capacitor c=0.042636f \
 //x=61.79 //y=7.4 //x2=61.05 //y2=2.59
cc_1554 ( N_VDD_c_1035_p N_noxref_16_c_5462_n ) capacitor c=0.00125279f \
 //x=84.73 //y=7.4 //x2=62.9 //y2=2.08
cc_1555 ( N_VDD_c_1578_p N_noxref_16_c_5462_n ) capacitor c=2.87256e-19 \
 //x=63.375 //y=7.4 //x2=62.9 //y2=2.08
cc_1556 ( N_VDD_c_1027_n N_noxref_16_c_5462_n ) capacitor c=0.0133961f \
 //x=61.79 //y=7.4 //x2=62.9 //y2=2.08
cc_1557 ( N_VDD_c_1578_p N_noxref_16_M128_noxref_g ) capacitor c=0.00726866f \
 //x=63.375 //y=7.4 //x2=62.8 //y2=6.02
cc_1558 ( N_VDD_M128_noxref_s N_noxref_16_M128_noxref_g ) capacitor \
 c=0.054195f //x=62.445 //y=5.02 //x2=62.8 //y2=6.02
cc_1559 ( N_VDD_c_1578_p N_noxref_16_M129_noxref_g ) capacitor c=0.00672952f \
 //x=63.375 //y=7.4 //x2=63.24 //y2=6.02
cc_1560 ( N_VDD_M129_noxref_d N_noxref_16_M129_noxref_g ) capacitor \
 c=0.015318f //x=63.315 //y=5.02 //x2=63.24 //y2=6.02
cc_1561 ( N_VDD_c_1027_n N_noxref_16_c_5496_n ) capacitor c=0.015293f \
 //x=61.79 //y=7.4 //x2=62.9 //y2=4.7
cc_1562 ( N_VDD_c_1035_p N_noxref_16_M122_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=58.365 //y2=5.02
cc_1563 ( N_VDD_c_1543_p N_noxref_16_M122_noxref_d ) capacitor c=0.014035f \
 //x=58.865 //y=7.4 //x2=58.365 //y2=5.02
cc_1564 ( N_VDD_M123_noxref_d N_noxref_16_M122_noxref_d ) capacitor \
 c=0.0664752f //x=58.805 //y=5.02 //x2=58.365 //y2=5.02
cc_1565 ( N_VDD_c_1035_p N_noxref_16_M124_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=59.245 //y2=5.02
cc_1566 ( N_VDD_c_1564_p N_noxref_16_M124_noxref_d ) capacitor c=0.014035f \
 //x=59.745 //y=7.4 //x2=59.245 //y2=5.02
cc_1567 ( N_VDD_c_1027_n N_noxref_16_M124_noxref_d ) capacitor c=4.9285e-19 \
 //x=61.79 //y=7.4 //x2=59.245 //y2=5.02
cc_1568 ( N_VDD_M122_noxref_s N_noxref_16_M124_noxref_d ) capacitor \
 c=0.00130656f //x=57.935 //y=5.02 //x2=59.245 //y2=5.02
cc_1569 ( N_VDD_M123_noxref_d N_noxref_16_M124_noxref_d ) capacitor \
 c=0.0664752f //x=58.805 //y=5.02 //x2=59.245 //y2=5.02
cc_1570 ( N_VDD_M125_noxref_d N_noxref_16_M124_noxref_d ) capacitor \
 c=0.0664752f //x=59.685 //y=5.02 //x2=59.245 //y2=5.02
cc_1571 ( N_VDD_c_1035_p N_noxref_16_M126_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=60.125 //y2=5.02
cc_1572 ( N_VDD_c_1570_p N_noxref_16_M126_noxref_d ) capacitor c=0.014035f \
 //x=60.625 //y=7.4 //x2=60.125 //y2=5.02
cc_1573 ( N_VDD_c_1027_n N_noxref_16_M126_noxref_d ) capacitor c=0.00939849f \
 //x=61.79 //y=7.4 //x2=60.125 //y2=5.02
cc_1574 ( N_VDD_M125_noxref_d N_noxref_16_M126_noxref_d ) capacitor \
 c=0.0664752f //x=59.685 //y=5.02 //x2=60.125 //y2=5.02
cc_1575 ( N_VDD_M127_noxref_d N_noxref_16_M126_noxref_d ) capacitor \
 c=0.0664752f //x=60.565 //y=5.02 //x2=60.125 //y2=5.02
cc_1576 ( N_VDD_M128_noxref_s N_noxref_16_M126_noxref_d ) capacitor \
 c=4.52683e-19 //x=62.445 //y=5.02 //x2=60.125 //y2=5.02
cc_1577 ( N_VDD_c_1035_p N_CLK_c_5631_n ) capacitor c=0.0679008f //x=84.73 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_1578 ( N_VDD_c_1139_p N_CLK_c_5631_n ) capacitor c=0.00258496f //x=7.97 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_1579 ( N_VDD_c_1602_p N_CLK_c_5631_n ) capacitor c=0.00328994f //x=9.145 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_1580 ( N_VDD_c_1056_p N_CLK_c_5631_n ) capacitor c=0.00135925f //x=10.025 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_1581 ( N_VDD_c_1087_p N_CLK_c_5631_n ) capacitor c=0.00258496f //x=12.78 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_1582 ( N_VDD_c_1605_p N_CLK_c_5631_n ) capacitor c=0.00209689f //x=13.655 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_1583 ( N_VDD_c_1091_p N_CLK_c_5631_n ) capacitor c=7.81728e-19 //x=14.535 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_1584 ( N_VDD_c_1014_n N_CLK_c_5631_n ) capacitor c=0.0389825f //x=8.14 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_1585 ( N_VDD_c_1015_n N_CLK_c_5631_n ) capacitor c=0.0389825f //x=12.95 \
 //y=7.4 //x2=14.685 //y2=4.44
cc_1586 ( N_VDD_M62_noxref_s N_CLK_c_5631_n ) capacitor c=0.00179496f \
 //x=9.095 //y=5.02 //x2=14.685 //y2=4.44
cc_1587 ( N_VDD_M68_noxref_s N_CLK_c_5631_n ) capacitor c=0.00541054f \
 //x=13.605 //y=5.02 //x2=14.685 //y2=4.44
cc_1588 ( N_VDD_c_1035_p N_CLK_c_5642_n ) capacitor c=0.00146064f //x=84.73 \
 //y=7.4 //x2=5.665 //y2=4.44
cc_1589 ( N_VDD_c_1035_p N_CLK_c_5643_n ) capacitor c=0.111938f //x=84.73 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1590 ( N_VDD_c_1613_p N_CLK_c_5643_n ) capacitor c=0.00205475f //x=16.11 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1591 ( N_VDD_c_1614_p N_CLK_c_5643_n ) capacitor c=0.00209689f //x=16.985 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1592 ( N_VDD_c_1142_p N_CLK_c_5643_n ) capacitor c=7.81728e-19 //x=17.865 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1593 ( N_VDD_c_1616_p N_CLK_c_5643_n ) capacitor c=0.00205475f //x=19.44 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1594 ( N_VDD_c_1617_p N_CLK_c_5643_n ) capacitor c=0.00328994f //x=20.615 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1595 ( N_VDD_c_1186_p N_CLK_c_5643_n ) capacitor c=0.00135925f //x=21.495 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1596 ( N_VDD_c_1619_p N_CLK_c_5643_n ) capacitor c=0.00258496f //x=24.25 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1597 ( N_VDD_c_1620_p N_CLK_c_5643_n ) capacitor c=0.00209689f //x=25.125 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1598 ( N_VDD_c_1242_p N_CLK_c_5643_n ) capacitor c=7.81728e-19 //x=26.005 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1599 ( N_VDD_c_1622_p N_CLK_c_5643_n ) capacitor c=0.00205475f //x=27.58 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1600 ( N_VDD_c_1623_p N_CLK_c_5643_n ) capacitor c=0.00328994f //x=28.755 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1601 ( N_VDD_c_1258_p N_CLK_c_5643_n ) capacitor c=0.00135925f //x=29.635 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1602 ( N_VDD_c_1016_n N_CLK_c_5643_n ) capacitor c=0.0389825f //x=16.28 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1603 ( N_VDD_c_1017_n N_CLK_c_5643_n ) capacitor c=0.0389825f //x=19.61 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1604 ( N_VDD_c_1018_n N_CLK_c_5643_n ) capacitor c=0.0392569f //x=24.42 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1605 ( N_VDD_c_1019_n N_CLK_c_5643_n ) capacitor c=0.0389825f //x=27.75 \
 //y=7.4 //x2=29.855 //y2=4.44
cc_1606 ( N_VDD_M71_noxref_d N_CLK_c_5643_n ) capacitor c=6.7165e-19 \
 //x=15.355 //y=5.02 //x2=29.855 //y2=4.44
cc_1607 ( N_VDD_M72_noxref_s N_CLK_c_5643_n ) capacitor c=0.00541054f \
 //x=16.935 //y=5.02 //x2=29.855 //y2=4.44
cc_1608 ( N_VDD_M75_noxref_d N_CLK_c_5643_n ) capacitor c=6.7165e-19 \
 //x=18.685 //y=5.02 //x2=29.855 //y2=4.44
cc_1609 ( N_VDD_M76_noxref_s N_CLK_c_5643_n ) capacitor c=0.00179496f \
 //x=20.565 //y=5.02 //x2=29.855 //y2=4.44
cc_1610 ( N_VDD_M82_noxref_s N_CLK_c_5643_n ) capacitor c=0.00541054f \
 //x=25.075 //y=5.02 //x2=29.855 //y2=4.44
cc_1611 ( N_VDD_M85_noxref_d N_CLK_c_5643_n ) capacitor c=6.7165e-19 \
 //x=26.825 //y=5.02 //x2=29.855 //y2=4.44
cc_1612 ( N_VDD_M86_noxref_s N_CLK_c_5643_n ) capacitor c=0.00179496f \
 //x=28.705 //y=5.02 //x2=29.855 //y2=4.44
cc_1613 ( N_VDD_c_1035_p N_CLK_c_5667_n ) capacitor c=0.00123805f //x=84.73 \
 //y=7.4 //x2=14.915 //y2=4.44
cc_1614 ( N_VDD_c_1035_p N_CLK_c_5668_n ) capacitor c=0.0679008f //x=84.73 \
 //y=7.4 //x2=39.105 //y2=4.44
cc_1615 ( N_VDD_c_1338_p N_CLK_c_5668_n ) capacitor c=0.00258496f //x=32.39 \
 //y=7.4 //x2=39.105 //y2=4.44
cc_1616 ( N_VDD_c_1639_p N_CLK_c_5668_n ) capacitor c=0.00328994f //x=33.565 \
 //y=7.4 //x2=39.105 //y2=4.44
cc_1617 ( N_VDD_c_1262_p N_CLK_c_5668_n ) capacitor c=0.00135925f //x=34.445 \
 //y=7.4 //x2=39.105 //y2=4.44
cc_1618 ( N_VDD_c_1293_p N_CLK_c_5668_n ) capacitor c=0.00258496f //x=37.2 \
 //y=7.4 //x2=39.105 //y2=4.44
cc_1619 ( N_VDD_c_1642_p N_CLK_c_5668_n ) capacitor c=0.00209689f //x=38.075 \
 //y=7.4 //x2=39.105 //y2=4.44
cc_1620 ( N_VDD_c_1297_p N_CLK_c_5668_n ) capacitor c=7.81728e-19 //x=38.955 \
 //y=7.4 //x2=39.105 //y2=4.44
cc_1621 ( N_VDD_c_1020_n N_CLK_c_5668_n ) capacitor c=0.0389825f //x=32.56 \
 //y=7.4 //x2=39.105 //y2=4.44
cc_1622 ( N_VDD_c_1021_n N_CLK_c_5668_n ) capacitor c=0.0389825f //x=37.37 \
 //y=7.4 //x2=39.105 //y2=4.44
cc_1623 ( N_VDD_M92_noxref_s N_CLK_c_5668_n ) capacitor c=0.00179496f \
 //x=33.515 //y=5.02 //x2=39.105 //y2=4.44
cc_1624 ( N_VDD_M98_noxref_s N_CLK_c_5668_n ) capacitor c=0.00541054f \
 //x=38.025 //y=5.02 //x2=39.105 //y2=4.44
cc_1625 ( N_VDD_c_1035_p N_CLK_c_5679_n ) capacitor c=0.00120845f //x=84.73 \
 //y=7.4 //x2=30.085 //y2=4.44
cc_1626 ( N_VDD_c_1035_p N_CLK_c_5680_n ) capacitor c=0.111938f //x=84.73 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1627 ( N_VDD_c_1650_p N_CLK_c_5680_n ) capacitor c=0.00205475f //x=40.53 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1628 ( N_VDD_c_1651_p N_CLK_c_5680_n ) capacitor c=0.00209689f //x=41.405 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1629 ( N_VDD_c_1341_p N_CLK_c_5680_n ) capacitor c=7.81728e-19 //x=42.285 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1630 ( N_VDD_c_1653_p N_CLK_c_5680_n ) capacitor c=0.00205475f //x=43.86 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1631 ( N_VDD_c_1654_p N_CLK_c_5680_n ) capacitor c=0.00328994f //x=45.035 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1632 ( N_VDD_c_1383_p N_CLK_c_5680_n ) capacitor c=0.00135925f //x=45.915 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1633 ( N_VDD_c_1459_p N_CLK_c_5680_n ) capacitor c=0.00258496f //x=48.67 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1634 ( N_VDD_c_1657_p N_CLK_c_5680_n ) capacitor c=0.00209689f //x=49.545 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1635 ( N_VDD_c_1505_p N_CLK_c_5680_n ) capacitor c=7.81728e-19 //x=50.425 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1636 ( N_VDD_c_1659_p N_CLK_c_5680_n ) capacitor c=0.00205475f //x=52 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1637 ( N_VDD_c_1660_p N_CLK_c_5680_n ) capacitor c=0.00328994f //x=53.175 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1638 ( N_VDD_c_1539_p N_CLK_c_5680_n ) capacitor c=0.00135925f //x=54.055 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1639 ( N_VDD_c_1022_n N_CLK_c_5680_n ) capacitor c=0.0389825f //x=40.7 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1640 ( N_VDD_c_1023_n N_CLK_c_5680_n ) capacitor c=0.0389825f //x=44.03 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1641 ( N_VDD_c_1024_n N_CLK_c_5680_n ) capacitor c=0.0392569f //x=48.84 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1642 ( N_VDD_c_1025_n N_CLK_c_5680_n ) capacitor c=0.0389825f //x=52.17 \
 //y=7.4 //x2=54.275 //y2=4.44
cc_1643 ( N_VDD_M101_noxref_d N_CLK_c_5680_n ) capacitor c=6.7165e-19 \
 //x=39.775 //y=5.02 //x2=54.275 //y2=4.44
cc_1644 ( N_VDD_M102_noxref_s N_CLK_c_5680_n ) capacitor c=0.00541054f \
 //x=41.355 //y=5.02 //x2=54.275 //y2=4.44
cc_1645 ( N_VDD_M105_noxref_d N_CLK_c_5680_n ) capacitor c=6.7165e-19 \
 //x=43.105 //y=5.02 //x2=54.275 //y2=4.44
cc_1646 ( N_VDD_M106_noxref_s N_CLK_c_5680_n ) capacitor c=0.00179496f \
 //x=44.985 //y=5.02 //x2=54.275 //y2=4.44
cc_1647 ( N_VDD_M112_noxref_s N_CLK_c_5680_n ) capacitor c=0.00541054f \
 //x=49.495 //y=5.02 //x2=54.275 //y2=4.44
cc_1648 ( N_VDD_M115_noxref_d N_CLK_c_5680_n ) capacitor c=6.7165e-19 \
 //x=51.245 //y=5.02 //x2=54.275 //y2=4.44
cc_1649 ( N_VDD_M116_noxref_s N_CLK_c_5680_n ) capacitor c=0.00179496f \
 //x=53.125 //y=5.02 //x2=54.275 //y2=4.44
cc_1650 ( N_VDD_c_1035_p N_CLK_c_5704_n ) capacitor c=0.00123805f //x=84.73 \
 //y=7.4 //x2=39.335 //y2=4.44
cc_1651 ( N_VDD_c_1035_p N_CLK_c_5705_n ) capacitor c=0.0693925f //x=84.73 \
 //y=7.4 //x2=63.525 //y2=4.44
cc_1652 ( N_VDD_c_1675_p N_CLK_c_5705_n ) capacitor c=0.00258496f //x=56.81 \
 //y=7.4 //x2=63.525 //y2=4.44
cc_1653 ( N_VDD_c_1676_p N_CLK_c_5705_n ) capacitor c=0.00328994f //x=57.985 \
 //y=7.4 //x2=63.525 //y2=4.44
cc_1654 ( N_VDD_c_1543_p N_CLK_c_5705_n ) capacitor c=0.00135925f //x=58.865 \
 //y=7.4 //x2=63.525 //y2=4.44
cc_1655 ( N_VDD_c_1574_p N_CLK_c_5705_n ) capacitor c=0.00258496f //x=61.62 \
 //y=7.4 //x2=63.525 //y2=4.44
cc_1656 ( N_VDD_c_1679_p N_CLK_c_5705_n ) capacitor c=0.00209689f //x=62.495 \
 //y=7.4 //x2=63.525 //y2=4.44
cc_1657 ( N_VDD_c_1578_p N_CLK_c_5705_n ) capacitor c=7.81728e-19 //x=63.375 \
 //y=7.4 //x2=63.525 //y2=4.44
cc_1658 ( N_VDD_c_1026_n N_CLK_c_5705_n ) capacitor c=0.0389825f //x=56.98 \
 //y=7.4 //x2=63.525 //y2=4.44
cc_1659 ( N_VDD_c_1027_n N_CLK_c_5705_n ) capacitor c=0.0389825f //x=61.79 \
 //y=7.4 //x2=63.525 //y2=4.44
cc_1660 ( N_VDD_M122_noxref_s N_CLK_c_5705_n ) capacitor c=0.00179496f \
 //x=57.935 //y=5.02 //x2=63.525 //y2=4.44
cc_1661 ( N_VDD_M128_noxref_s N_CLK_c_5705_n ) capacitor c=0.00541054f \
 //x=62.445 //y=5.02 //x2=63.525 //y2=4.44
cc_1662 ( N_VDD_c_1035_p N_CLK_c_5716_n ) capacitor c=0.00120845f //x=84.73 \
 //y=7.4 //x2=54.505 //y2=4.44
cc_1663 ( N_VDD_c_1035_p N_CLK_c_5622_n ) capacitor c=2.03287e-19 //x=84.73 \
 //y=7.4 //x2=5.55 //y2=2.08
cc_1664 ( N_VDD_c_1013_n N_CLK_c_5622_n ) capacitor c=8.47879e-19 //x=3.33 \
 //y=7.4 //x2=5.55 //y2=2.08
cc_1665 ( N_VDD_c_1015_n N_CLK_c_5623_n ) capacitor c=4.60777e-19 //x=12.95 \
 //y=7.4 //x2=14.8 //y2=2.08
cc_1666 ( N_VDD_c_1016_n N_CLK_c_5623_n ) capacitor c=3.65649e-19 //x=16.28 \
 //y=7.4 //x2=14.8 //y2=2.08
cc_1667 ( N_VDD_c_1035_p N_CLK_c_5625_n ) capacitor c=2.03287e-19 //x=84.73 \
 //y=7.4 //x2=29.97 //y2=2.08
cc_1668 ( N_VDD_c_1019_n N_CLK_c_5625_n ) capacitor c=6.15921e-19 //x=27.75 \
 //y=7.4 //x2=29.97 //y2=2.08
cc_1669 ( N_VDD_c_1021_n N_CLK_c_5626_n ) capacitor c=4.60777e-19 //x=37.37 \
 //y=7.4 //x2=39.22 //y2=2.08
cc_1670 ( N_VDD_c_1022_n N_CLK_c_5626_n ) capacitor c=3.65649e-19 //x=40.7 \
 //y=7.4 //x2=39.22 //y2=2.08
cc_1671 ( N_VDD_c_1035_p N_CLK_c_5628_n ) capacitor c=2.03287e-19 //x=84.73 \
 //y=7.4 //x2=54.39 //y2=2.08
cc_1672 ( N_VDD_c_1025_n N_CLK_c_5628_n ) capacitor c=6.15921e-19 //x=52.17 \
 //y=7.4 //x2=54.39 //y2=2.08
cc_1673 ( N_VDD_c_1027_n N_CLK_c_5629_n ) capacitor c=4.60777e-19 //x=61.79 \
 //y=7.4 //x2=63.64 //y2=2.08
cc_1674 ( N_VDD_c_1028_n N_CLK_c_5629_n ) capacitor c=7.28243e-19 //x=65.12 \
 //y=7.4 //x2=63.64 //y2=2.08
cc_1675 ( N_VDD_c_1129_p N_CLK_M58_noxref_g ) capacitor c=0.00676195f \
 //x=6.095 //y=7.4 //x2=5.52 //y2=6.02
cc_1676 ( N_VDD_M57_noxref_d N_CLK_M58_noxref_g ) capacitor c=0.015318f \
 //x=5.155 //y=5.02 //x2=5.52 //y2=6.02
cc_1677 ( N_VDD_c_1129_p N_CLK_M59_noxref_g ) capacitor c=0.00675175f \
 //x=6.095 //y=7.4 //x2=5.96 //y2=6.02
cc_1678 ( N_VDD_M59_noxref_d N_CLK_M59_noxref_g ) capacitor c=0.015318f \
 //x=6.035 //y=5.02 //x2=5.96 //y2=6.02
cc_1679 ( N_VDD_c_1207_p N_CLK_M70_noxref_g ) capacitor c=0.00673971f \
 //x=15.415 //y=7.4 //x2=14.84 //y2=6.02
cc_1680 ( N_VDD_M69_noxref_d N_CLK_M70_noxref_g ) capacitor c=0.015318f \
 //x=14.475 //y=5.02 //x2=14.84 //y2=6.02
cc_1681 ( N_VDD_c_1207_p N_CLK_M71_noxref_g ) capacitor c=0.00672952f \
 //x=15.415 //y=7.4 //x2=15.28 //y2=6.02
cc_1682 ( N_VDD_c_1016_n N_CLK_M71_noxref_g ) capacitor c=0.00864163f \
 //x=16.28 //y=7.4 //x2=15.28 //y2=6.02
cc_1683 ( N_VDD_M71_noxref_d N_CLK_M71_noxref_g ) capacitor c=0.0430452f \
 //x=15.355 //y=5.02 //x2=15.28 //y2=6.02
cc_1684 ( N_VDD_c_1328_p N_CLK_M88_noxref_g ) capacitor c=0.00676195f \
 //x=30.515 //y=7.4 //x2=29.94 //y2=6.02
cc_1685 ( N_VDD_M87_noxref_d N_CLK_M88_noxref_g ) capacitor c=0.015318f \
 //x=29.575 //y=5.02 //x2=29.94 //y2=6.02
cc_1686 ( N_VDD_c_1328_p N_CLK_M89_noxref_g ) capacitor c=0.00675175f \
 //x=30.515 //y=7.4 //x2=30.38 //y2=6.02
cc_1687 ( N_VDD_M89_noxref_d N_CLK_M89_noxref_g ) capacitor c=0.015318f \
 //x=30.455 //y=5.02 //x2=30.38 //y2=6.02
cc_1688 ( N_VDD_c_1404_p N_CLK_M100_noxref_g ) capacitor c=0.00673971f \
 //x=39.835 //y=7.4 //x2=39.26 //y2=6.02
cc_1689 ( N_VDD_M99_noxref_d N_CLK_M100_noxref_g ) capacitor c=0.015318f \
 //x=38.895 //y=5.02 //x2=39.26 //y2=6.02
cc_1690 ( N_VDD_c_1404_p N_CLK_M101_noxref_g ) capacitor c=0.00672952f \
 //x=39.835 //y=7.4 //x2=39.7 //y2=6.02
cc_1691 ( N_VDD_c_1022_n N_CLK_M101_noxref_g ) capacitor c=0.00864163f \
 //x=40.7 //y=7.4 //x2=39.7 //y2=6.02
cc_1692 ( N_VDD_M101_noxref_d N_CLK_M101_noxref_g ) capacitor c=0.0430452f \
 //x=39.775 //y=5.02 //x2=39.7 //y2=6.02
cc_1693 ( N_VDD_c_1716_p N_CLK_M118_noxref_g ) capacitor c=0.00676195f \
 //x=54.935 //y=7.4 //x2=54.36 //y2=6.02
cc_1694 ( N_VDD_M117_noxref_d N_CLK_M118_noxref_g ) capacitor c=0.015318f \
 //x=53.995 //y=5.02 //x2=54.36 //y2=6.02
cc_1695 ( N_VDD_c_1716_p N_CLK_M119_noxref_g ) capacitor c=0.00675175f \
 //x=54.935 //y=7.4 //x2=54.8 //y2=6.02
cc_1696 ( N_VDD_M119_noxref_d N_CLK_M119_noxref_g ) capacitor c=0.015318f \
 //x=54.875 //y=5.02 //x2=54.8 //y2=6.02
cc_1697 ( N_VDD_c_1720_p N_CLK_M130_noxref_g ) capacitor c=0.00673971f \
 //x=64.255 //y=7.4 //x2=63.68 //y2=6.02
cc_1698 ( N_VDD_M129_noxref_d N_CLK_M130_noxref_g ) capacitor c=0.015318f \
 //x=63.315 //y=5.02 //x2=63.68 //y2=6.02
cc_1699 ( N_VDD_c_1720_p N_CLK_M131_noxref_g ) capacitor c=0.00672952f \
 //x=64.255 //y=7.4 //x2=64.12 //y2=6.02
cc_1700 ( N_VDD_c_1028_n N_CLK_M131_noxref_g ) capacitor c=0.00829014f \
 //x=65.12 //y=7.4 //x2=64.12 //y2=6.02
cc_1701 ( N_VDD_M131_noxref_d N_CLK_M131_noxref_g ) capacitor c=0.0430452f \
 //x=64.195 //y=5.02 //x2=64.12 //y2=6.02
cc_1702 ( N_VDD_c_1025_n N_noxref_18_c_6392_n ) capacitor c=0.0143396f \
 //x=52.17 //y=7.4 //x2=56.12 //y2=4.07
cc_1703 ( N_VDD_c_1035_p N_noxref_18_c_6393_n ) capacitor c=0.046539f \
 //x=84.73 //y=7.4 //x2=66.115 //y2=4.07
cc_1704 ( N_VDD_c_1727_p N_noxref_18_c_6393_n ) capacitor c=0.00168692f \
 //x=64.95 //y=7.4 //x2=66.115 //y2=4.07
cc_1705 ( N_VDD_c_1728_p N_noxref_18_c_6393_n ) capacitor c=0.00172186f \
 //x=65.825 //y=7.4 //x2=66.115 //y2=4.07
cc_1706 ( N_VDD_c_1729_p N_noxref_18_c_6393_n ) capacitor c=6.62004e-19 \
 //x=66.705 //y=7.4 //x2=66.115 //y2=4.07
cc_1707 ( N_VDD_c_1026_n N_noxref_18_c_6393_n ) capacitor c=0.0140578f \
 //x=56.98 //y=7.4 //x2=66.115 //y2=4.07
cc_1708 ( N_VDD_c_1027_n N_noxref_18_c_6393_n ) capacitor c=0.0140578f \
 //x=61.79 //y=7.4 //x2=66.115 //y2=4.07
cc_1709 ( N_VDD_c_1028_n N_noxref_18_c_6393_n ) capacitor c=0.0277022f \
 //x=65.12 //y=7.4 //x2=66.115 //y2=4.07
cc_1710 ( N_VDD_M131_noxref_d N_noxref_18_c_6393_n ) capacitor c=5.05307e-19 \
 //x=64.195 //y=5.02 //x2=66.115 //y2=4.07
cc_1711 ( N_VDD_M132_noxref_s N_noxref_18_c_6393_n ) capacitor c=0.00363031f \
 //x=65.775 //y=5.02 //x2=66.115 //y2=4.07
cc_1712 ( N_VDD_c_1026_n N_noxref_18_c_6402_n ) capacitor c=0.00104411f \
 //x=56.98 //y=7.4 //x2=56.35 //y2=4.07
cc_1713 ( N_VDD_c_1024_n N_noxref_18_c_6377_n ) capacitor c=5.18578e-19 \
 //x=48.84 //y=7.4 //x2=50.69 //y2=2.08
cc_1714 ( N_VDD_c_1025_n N_noxref_18_c_6377_n ) capacitor c=3.21957e-19 \
 //x=52.17 //y=7.4 //x2=50.69 //y2=2.08
cc_1715 ( N_VDD_c_1035_p N_noxref_18_c_6405_n ) capacitor c=0.00444751f \
 //x=84.73 //y=7.4 //x2=54.495 //y2=5.155
cc_1716 ( N_VDD_c_1539_p N_noxref_18_c_6405_n ) capacitor c=4.31931e-19 \
 //x=54.055 //y=7.4 //x2=54.495 //y2=5.155
cc_1717 ( N_VDD_c_1716_p N_noxref_18_c_6405_n ) capacitor c=4.31906e-19 \
 //x=54.935 //y=7.4 //x2=54.495 //y2=5.155
cc_1718 ( N_VDD_M117_noxref_d N_noxref_18_c_6405_n ) capacitor c=0.0112985f \
 //x=53.995 //y=5.02 //x2=54.495 //y2=5.155
cc_1719 ( N_VDD_c_1025_n N_noxref_18_c_6409_n ) capacitor c=0.00863585f \
 //x=52.17 //y=7.4 //x2=53.785 //y2=5.155
cc_1720 ( N_VDD_M116_noxref_s N_noxref_18_c_6409_n ) capacitor c=0.0831083f \
 //x=53.125 //y=5.02 //x2=53.785 //y2=5.155
cc_1721 ( N_VDD_c_1035_p N_noxref_18_c_6411_n ) capacitor c=0.0044221f \
 //x=84.73 //y=7.4 //x2=55.375 //y2=5.155
cc_1722 ( N_VDD_c_1716_p N_noxref_18_c_6411_n ) capacitor c=4.31931e-19 \
 //x=54.935 //y=7.4 //x2=55.375 //y2=5.155
cc_1723 ( N_VDD_c_1746_p N_noxref_18_c_6411_n ) capacitor c=4.31931e-19 \
 //x=55.815 //y=7.4 //x2=55.375 //y2=5.155
cc_1724 ( N_VDD_M119_noxref_d N_noxref_18_c_6411_n ) capacitor c=0.0112985f \
 //x=54.875 //y=5.02 //x2=55.375 //y2=5.155
cc_1725 ( N_VDD_c_1035_p N_noxref_18_c_6415_n ) capacitor c=0.00433242f \
 //x=84.73 //y=7.4 //x2=56.155 //y2=5.155
cc_1726 ( N_VDD_c_1746_p N_noxref_18_c_6415_n ) capacitor c=7.46626e-19 \
 //x=55.815 //y=7.4 //x2=56.155 //y2=5.155
cc_1727 ( N_VDD_c_1675_p N_noxref_18_c_6415_n ) capacitor c=0.00198565f \
 //x=56.81 //y=7.4 //x2=56.155 //y2=5.155
cc_1728 ( N_VDD_M121_noxref_d N_noxref_18_c_6415_n ) capacitor c=0.0112985f \
 //x=55.755 //y=5.02 //x2=56.155 //y2=5.155
cc_1729 ( N_VDD_c_1035_p N_noxref_18_c_6380_n ) capacitor c=0.00126142f \
 //x=84.73 //y=7.4 //x2=66.23 //y2=2.08
cc_1730 ( N_VDD_c_1729_p N_noxref_18_c_6380_n ) capacitor c=2.8777e-19 \
 //x=66.705 //y=7.4 //x2=66.23 //y2=2.08
cc_1731 ( N_VDD_c_1028_n N_noxref_18_c_6380_n ) capacitor c=0.0152982f \
 //x=65.12 //y=7.4 //x2=66.23 //y2=2.08
cc_1732 ( N_VDD_c_1026_n N_noxref_18_c_6422_n ) capacitor c=0.0427201f \
 //x=56.98 //y=7.4 //x2=56.235 //y2=4.07
cc_1733 ( N_VDD_c_1524_p N_noxref_18_M114_noxref_g ) capacitor c=0.00673971f \
 //x=51.305 //y=7.4 //x2=50.73 //y2=6.02
cc_1734 ( N_VDD_M113_noxref_d N_noxref_18_M114_noxref_g ) capacitor \
 c=0.015318f //x=50.365 //y=5.02 //x2=50.73 //y2=6.02
cc_1735 ( N_VDD_c_1524_p N_noxref_18_M115_noxref_g ) capacitor c=0.00672952f \
 //x=51.305 //y=7.4 //x2=51.17 //y2=6.02
cc_1736 ( N_VDD_c_1025_n N_noxref_18_M115_noxref_g ) capacitor c=0.00928743f \
 //x=52.17 //y=7.4 //x2=51.17 //y2=6.02
cc_1737 ( N_VDD_M115_noxref_d N_noxref_18_M115_noxref_g ) capacitor \
 c=0.0430452f //x=51.245 //y=5.02 //x2=51.17 //y2=6.02
cc_1738 ( N_VDD_c_1729_p N_noxref_18_M132_noxref_g ) capacitor c=0.00726866f \
 //x=66.705 //y=7.4 //x2=66.13 //y2=6.02
cc_1739 ( N_VDD_M132_noxref_s N_noxref_18_M132_noxref_g ) capacitor \
 c=0.054195f //x=65.775 //y=5.02 //x2=66.13 //y2=6.02
cc_1740 ( N_VDD_c_1729_p N_noxref_18_M133_noxref_g ) capacitor c=0.00672952f \
 //x=66.705 //y=7.4 //x2=66.57 //y2=6.02
cc_1741 ( N_VDD_M133_noxref_d N_noxref_18_M133_noxref_g ) capacitor \
 c=0.015318f //x=66.645 //y=5.02 //x2=66.57 //y2=6.02
cc_1742 ( N_VDD_c_1028_n N_noxref_18_c_6432_n ) capacitor c=0.0137692f \
 //x=65.12 //y=7.4 //x2=66.23 //y2=4.7
cc_1743 ( N_VDD_c_1035_p N_noxref_18_M116_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=53.555 //y2=5.02
cc_1744 ( N_VDD_c_1539_p N_noxref_18_M116_noxref_d ) capacitor c=0.014035f \
 //x=54.055 //y=7.4 //x2=53.555 //y2=5.02
cc_1745 ( N_VDD_M117_noxref_d N_noxref_18_M116_noxref_d ) capacitor \
 c=0.0664752f //x=53.995 //y=5.02 //x2=53.555 //y2=5.02
cc_1746 ( N_VDD_c_1035_p N_noxref_18_M118_noxref_d ) capacitor c=0.00275186f \
 //x=84.73 //y=7.4 //x2=54.435 //y2=5.02
cc_1747 ( N_VDD_c_1716_p N_noxref_18_M118_noxref_d ) capacitor c=0.0140346f \
 //x=54.935 //y=7.4 //x2=54.435 //y2=5.02
cc_1748 ( N_VDD_c_1026_n N_noxref_18_M118_noxref_d ) capacitor c=4.9285e-19 \
 //x=56.98 //y=7.4 //x2=54.435 //y2=5.02
cc_1749 ( N_VDD_M116_noxref_s N_noxref_18_M118_noxref_d ) capacitor \
 c=0.00130656f //x=53.125 //y=5.02 //x2=54.435 //y2=5.02
cc_1750 ( N_VDD_M117_noxref_d N_noxref_18_M118_noxref_d ) capacitor \
 c=0.0664752f //x=53.995 //y=5.02 //x2=54.435 //y2=5.02
cc_1751 ( N_VDD_M119_noxref_d N_noxref_18_M118_noxref_d ) capacitor \
 c=0.0664752f //x=54.875 //y=5.02 //x2=54.435 //y2=5.02
cc_1752 ( N_VDD_c_1035_p N_noxref_18_M120_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=55.315 //y2=5.02
cc_1753 ( N_VDD_c_1746_p N_noxref_18_M120_noxref_d ) capacitor c=0.014035f \
 //x=55.815 //y=7.4 //x2=55.315 //y2=5.02
cc_1754 ( N_VDD_c_1026_n N_noxref_18_M120_noxref_d ) capacitor c=0.00939849f \
 //x=56.98 //y=7.4 //x2=55.315 //y2=5.02
cc_1755 ( N_VDD_M119_noxref_d N_noxref_18_M120_noxref_d ) capacitor \
 c=0.0664752f //x=54.875 //y=5.02 //x2=55.315 //y2=5.02
cc_1756 ( N_VDD_M121_noxref_d N_noxref_18_M120_noxref_d ) capacitor \
 c=0.0664752f //x=55.755 //y=5.02 //x2=55.315 //y2=5.02
cc_1757 ( N_VDD_M122_noxref_s N_noxref_18_M120_noxref_d ) capacitor \
 c=3.57641e-19 //x=57.935 //y=5.02 //x2=55.315 //y2=5.02
cc_1758 ( N_VDD_c_1035_p N_noxref_19_c_6684_n ) capacitor c=0.017007f \
 //x=84.73 //y=7.4 //x2=69.445 //y2=4.81
cc_1759 ( N_VDD_c_1782_p N_noxref_19_c_6684_n ) capacitor c=0.00238461f \
 //x=68.28 //y=7.4 //x2=69.445 //y2=4.81
cc_1760 ( N_VDD_c_1783_p N_noxref_19_c_6684_n ) capacitor c=0.00393349f \
 //x=69.455 //y=7.4 //x2=69.445 //y2=4.81
cc_1761 ( N_VDD_c_1784_p N_noxref_19_c_6684_n ) capacitor c=2.77727e-19 \
 //x=70.335 //y=7.4 //x2=69.445 //y2=4.81
cc_1762 ( N_VDD_c_1029_n N_noxref_19_c_6684_n ) capacitor c=0.0394216f \
 //x=68.45 //y=7.4 //x2=69.445 //y2=4.81
cc_1763 ( N_VDD_M136_noxref_s N_noxref_19_c_6684_n ) capacitor c=0.00294577f \
 //x=69.405 //y=5.02 //x2=69.445 //y2=4.81
cc_1764 ( N_VDD_c_1035_p N_noxref_19_c_6690_n ) capacitor c=0.00240887f \
 //x=84.73 //y=7.4 //x2=67.825 //y2=4.81
cc_1765 ( N_VDD_c_1028_n N_noxref_19_c_6690_n ) capacitor c=4.80672e-19 \
 //x=65.12 //y=7.4 //x2=67.825 //y2=4.81
cc_1766 ( N_VDD_c_1029_n N_noxref_19_c_6690_n ) capacitor c=0.00102529f \
 //x=68.45 //y=7.4 //x2=67.825 //y2=4.81
cc_1767 ( N_VDD_M135_noxref_d N_noxref_19_c_6690_n ) capacitor c=0.00101443f \
 //x=67.525 //y=5.02 //x2=67.825 //y2=4.81
cc_1768 ( N_VDD_c_1035_p N_noxref_19_c_6694_n ) capacitor c=0.00460596f \
 //x=84.73 //y=7.4 //x2=67.145 //y2=5.2
cc_1769 ( N_VDD_c_1729_p N_noxref_19_c_6694_n ) capacitor c=4.3394e-19 \
 //x=66.705 //y=7.4 //x2=67.145 //y2=5.2
cc_1770 ( N_VDD_c_1793_p N_noxref_19_c_6694_n ) capacitor c=4.48377e-19 \
 //x=67.585 //y=7.4 //x2=67.145 //y2=5.2
cc_1771 ( N_VDD_M133_noxref_d N_noxref_19_c_6694_n ) capacitor c=0.0127013f \
 //x=66.645 //y=5.02 //x2=67.145 //y2=5.2
cc_1772 ( N_VDD_c_1028_n N_noxref_19_c_6698_n ) capacitor c=0.00985474f \
 //x=65.12 //y=7.4 //x2=66.435 //y2=5.2
cc_1773 ( N_VDD_M132_noxref_s N_noxref_19_c_6698_n ) capacitor c=0.087833f \
 //x=65.775 //y=5.02 //x2=66.435 //y2=5.2
cc_1774 ( N_VDD_c_1035_p N_noxref_19_c_6700_n ) capacitor c=0.00297776f \
 //x=84.73 //y=7.4 //x2=67.625 //y2=5.2
cc_1775 ( N_VDD_c_1793_p N_noxref_19_c_6700_n ) capacitor c=7.72068e-19 \
 //x=67.585 //y=7.4 //x2=67.625 //y2=5.2
cc_1776 ( N_VDD_M135_noxref_d N_noxref_19_c_6700_n ) capacitor c=0.0153695f \
 //x=67.525 //y=5.02 //x2=67.625 //y2=5.2
cc_1777 ( N_VDD_c_1028_n N_noxref_19_c_6669_n ) capacitor c=0.0013137f \
 //x=65.12 //y=7.4 //x2=67.71 //y2=4.81
cc_1778 ( N_VDD_c_1029_n N_noxref_19_c_6669_n ) capacitor c=0.0412116f \
 //x=68.45 //y=7.4 //x2=67.71 //y2=4.81
cc_1779 ( N_VDD_M135_noxref_d N_noxref_19_c_6669_n ) capacitor c=3.11243e-19 \
 //x=67.525 //y=5.02 //x2=67.71 //y2=4.81
cc_1780 ( N_VDD_c_1035_p N_noxref_19_c_6670_n ) capacitor c=4.53525e-19 \
 //x=84.73 //y=7.4 //x2=69.56 //y2=2.08
cc_1781 ( N_VDD_c_1029_n N_noxref_19_c_6670_n ) capacitor c=0.0144919f \
 //x=68.45 //y=7.4 //x2=69.56 //y2=2.08
cc_1782 ( N_VDD_M136_noxref_s N_noxref_19_c_6670_n ) capacitor c=0.0192205f \
 //x=69.405 //y=5.02 //x2=69.56 //y2=2.08
cc_1783 ( N_VDD_c_1784_p N_noxref_19_M136_noxref_g ) capacitor c=0.00749687f \
 //x=70.335 //y=7.4 //x2=69.76 //y2=6.02
cc_1784 ( N_VDD_M136_noxref_s N_noxref_19_M136_noxref_g ) capacitor \
 c=0.0477201f //x=69.405 //y=5.02 //x2=69.76 //y2=6.02
cc_1785 ( N_VDD_c_1784_p N_noxref_19_M137_noxref_g ) capacitor c=0.00675175f \
 //x=70.335 //y=7.4 //x2=70.2 //y2=6.02
cc_1786 ( N_VDD_M137_noxref_d N_noxref_19_M137_noxref_g ) capacitor \
 c=0.015318f //x=70.275 //y=5.02 //x2=70.2 //y2=6.02
cc_1787 ( N_VDD_c_1029_n N_noxref_19_c_6713_n ) capacitor c=0.00511046f \
 //x=68.45 //y=7.4 //x2=69.835 //y2=4.79
cc_1788 ( N_VDD_M136_noxref_s N_noxref_19_c_6713_n ) capacitor c=0.00293141f \
 //x=69.405 //y=5.02 //x2=69.835 //y2=4.79
cc_1789 ( N_VDD_c_1035_p N_noxref_19_M132_noxref_d ) capacitor c=0.00287944f \
 //x=84.73 //y=7.4 //x2=66.205 //y2=5.02
cc_1790 ( N_VDD_c_1729_p N_noxref_19_M132_noxref_d ) capacitor c=0.014004f \
 //x=66.705 //y=7.4 //x2=66.205 //y2=5.02
cc_1791 ( N_VDD_c_1029_n N_noxref_19_M132_noxref_d ) capacitor c=6.94454e-19 \
 //x=68.45 //y=7.4 //x2=66.205 //y2=5.02
cc_1792 ( N_VDD_M133_noxref_d N_noxref_19_M132_noxref_d ) capacitor \
 c=0.0664752f //x=66.645 //y=5.02 //x2=66.205 //y2=5.02
cc_1793 ( N_VDD_c_1035_p N_noxref_19_M134_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=67.085 //y2=5.02
cc_1794 ( N_VDD_c_1793_p N_noxref_19_M134_noxref_d ) capacitor c=0.0140317f \
 //x=67.585 //y=7.4 //x2=67.085 //y2=5.02
cc_1795 ( N_VDD_c_1029_n N_noxref_19_M134_noxref_d ) capacitor c=0.0120541f \
 //x=68.45 //y=7.4 //x2=67.085 //y2=5.02
cc_1796 ( N_VDD_M132_noxref_s N_noxref_19_M134_noxref_d ) capacitor \
 c=0.00111971f //x=65.775 //y=5.02 //x2=67.085 //y2=5.02
cc_1797 ( N_VDD_M133_noxref_d N_noxref_19_M134_noxref_d ) capacitor \
 c=0.0664752f //x=66.645 //y=5.02 //x2=67.085 //y2=5.02
cc_1798 ( N_VDD_M135_noxref_d N_noxref_19_M134_noxref_d ) capacitor \
 c=0.0664752f //x=67.525 //y=5.02 //x2=67.085 //y2=5.02
cc_1799 ( N_VDD_M136_noxref_s N_noxref_19_M134_noxref_d ) capacitor \
 c=3.73257e-19 //x=69.405 //y=5.02 //x2=67.085 //y2=5.02
cc_1800 ( N_VDD_c_1035_p N_SN_c_6888_n ) capacitor c=2.03486e-19 //x=84.73 \
 //y=7.4 //x2=10.36 //y2=2.08
cc_1801 ( N_VDD_c_1014_n N_SN_c_6888_n ) capacitor c=6.15069e-19 //x=8.14 \
 //y=7.4 //x2=10.36 //y2=2.08
cc_1802 ( N_VDD_c_1035_p N_SN_c_6889_n ) capacitor c=2.03486e-19 //x=84.73 \
 //y=7.4 //x2=21.83 //y2=2.08
cc_1803 ( N_VDD_c_1017_n N_SN_c_6889_n ) capacitor c=6.85864e-19 //x=19.61 \
 //y=7.4 //x2=21.83 //y2=2.08
cc_1804 ( N_VDD_c_1035_p N_SN_c_6890_n ) capacitor c=2.03486e-19 //x=84.73 \
 //y=7.4 //x2=34.78 //y2=2.08
cc_1805 ( N_VDD_c_1020_n N_SN_c_6890_n ) capacitor c=6.15069e-19 //x=32.56 \
 //y=7.4 //x2=34.78 //y2=2.08
cc_1806 ( N_VDD_c_1035_p N_SN_c_6891_n ) capacitor c=2.03486e-19 //x=84.73 \
 //y=7.4 //x2=46.25 //y2=2.08
cc_1807 ( N_VDD_c_1023_n N_SN_c_6891_n ) capacitor c=5.89117e-19 //x=44.03 \
 //y=7.4 //x2=46.25 //y2=2.08
cc_1808 ( N_VDD_c_1035_p N_SN_c_6892_n ) capacitor c=2.03486e-19 //x=84.73 \
 //y=7.4 //x2=59.2 //y2=2.08
cc_1809 ( N_VDD_c_1026_n N_SN_c_6892_n ) capacitor c=6.15069e-19 //x=56.98 \
 //y=7.4 //x2=59.2 //y2=2.08
cc_1810 ( N_VDD_c_1035_p N_SN_c_6893_n ) capacitor c=2.03486e-19 //x=84.73 \
 //y=7.4 //x2=70.67 //y2=2.08
cc_1811 ( N_VDD_c_1029_n N_SN_c_6893_n ) capacitor c=4.25577e-19 //x=68.45 \
 //y=7.4 //x2=70.67 //y2=2.08
cc_1812 ( N_VDD_c_1077_p N_SN_M64_noxref_g ) capacitor c=0.00676195f \
 //x=10.905 //y=7.4 //x2=10.33 //y2=6.02
cc_1813 ( N_VDD_M63_noxref_d N_SN_M64_noxref_g ) capacitor c=0.015318f \
 //x=9.965 //y=5.02 //x2=10.33 //y2=6.02
cc_1814 ( N_VDD_c_1077_p N_SN_M65_noxref_g ) capacitor c=0.00675175f \
 //x=10.905 //y=7.4 //x2=10.77 //y2=6.02
cc_1815 ( N_VDD_M65_noxref_d N_SN_M65_noxref_g ) capacitor c=0.015318f \
 //x=10.845 //y=5.02 //x2=10.77 //y2=6.02
cc_1816 ( N_VDD_c_1839_p N_SN_M78_noxref_g ) capacitor c=0.00676195f \
 //x=22.375 //y=7.4 //x2=21.8 //y2=6.02
cc_1817 ( N_VDD_M77_noxref_d N_SN_M78_noxref_g ) capacitor c=0.015318f \
 //x=21.435 //y=5.02 //x2=21.8 //y2=6.02
cc_1818 ( N_VDD_c_1839_p N_SN_M79_noxref_g ) capacitor c=0.00675175f \
 //x=22.375 //y=7.4 //x2=22.24 //y2=6.02
cc_1819 ( N_VDD_M79_noxref_d N_SN_M79_noxref_g ) capacitor c=0.015318f \
 //x=22.315 //y=5.02 //x2=22.24 //y2=6.02
cc_1820 ( N_VDD_c_1283_p N_SN_M94_noxref_g ) capacitor c=0.00676195f \
 //x=35.325 //y=7.4 //x2=34.75 //y2=6.02
cc_1821 ( N_VDD_M93_noxref_d N_SN_M94_noxref_g ) capacitor c=0.015318f \
 //x=34.385 //y=5.02 //x2=34.75 //y2=6.02
cc_1822 ( N_VDD_c_1283_p N_SN_M95_noxref_g ) capacitor c=0.00675175f \
 //x=35.325 //y=7.4 //x2=35.19 //y2=6.02
cc_1823 ( N_VDD_M95_noxref_d N_SN_M95_noxref_g ) capacitor c=0.015318f \
 //x=35.265 //y=5.02 //x2=35.19 //y2=6.02
cc_1824 ( N_VDD_c_1449_p N_SN_M108_noxref_g ) capacitor c=0.00676195f \
 //x=46.795 //y=7.4 //x2=46.22 //y2=6.02
cc_1825 ( N_VDD_M107_noxref_d N_SN_M108_noxref_g ) capacitor c=0.015318f \
 //x=45.855 //y=5.02 //x2=46.22 //y2=6.02
cc_1826 ( N_VDD_c_1449_p N_SN_M109_noxref_g ) capacitor c=0.00675175f \
 //x=46.795 //y=7.4 //x2=46.66 //y2=6.02
cc_1827 ( N_VDD_M109_noxref_d N_SN_M109_noxref_g ) capacitor c=0.015318f \
 //x=46.735 //y=5.02 //x2=46.66 //y2=6.02
cc_1828 ( N_VDD_c_1564_p N_SN_M124_noxref_g ) capacitor c=0.00676195f \
 //x=59.745 //y=7.4 //x2=59.17 //y2=6.02
cc_1829 ( N_VDD_M123_noxref_d N_SN_M124_noxref_g ) capacitor c=0.015318f \
 //x=58.805 //y=5.02 //x2=59.17 //y2=6.02
cc_1830 ( N_VDD_c_1564_p N_SN_M125_noxref_g ) capacitor c=0.00675175f \
 //x=59.745 //y=7.4 //x2=59.61 //y2=6.02
cc_1831 ( N_VDD_M125_noxref_d N_SN_M125_noxref_g ) capacitor c=0.015318f \
 //x=59.685 //y=5.02 //x2=59.61 //y2=6.02
cc_1832 ( N_VDD_c_1855_p N_SN_M138_noxref_g ) capacitor c=0.00676195f \
 //x=71.215 //y=7.4 //x2=70.64 //y2=6.02
cc_1833 ( N_VDD_M137_noxref_d N_SN_M138_noxref_g ) capacitor c=0.015318f \
 //x=70.275 //y=5.02 //x2=70.64 //y2=6.02
cc_1834 ( N_VDD_c_1855_p N_SN_M139_noxref_g ) capacitor c=0.00675175f \
 //x=71.215 //y=7.4 //x2=71.08 //y2=6.02
cc_1835 ( N_VDD_M139_noxref_d N_SN_M139_noxref_g ) capacitor c=0.015318f \
 //x=71.155 //y=5.02 //x2=71.08 //y2=6.02
cc_1836 ( N_VDD_c_1035_p N_noxref_21_c_7656_n ) capacitor c=0.0145792f \
 //x=84.73 //y=7.4 //x2=71.665 //y2=3.7
cc_1837 ( N_VDD_c_1029_n N_noxref_21_c_7656_n ) capacitor c=0.00686843f \
 //x=68.45 //y=7.4 //x2=71.665 //y2=3.7
cc_1838 ( N_VDD_c_1026_n N_noxref_21_c_7648_n ) capacitor c=7.21808e-19 \
 //x=56.98 //y=7.4 //x2=55.5 //y2=2.08
cc_1839 ( N_VDD_c_1027_n N_noxref_21_c_7649_n ) capacitor c=6.21611e-19 \
 //x=61.79 //y=7.4 //x2=60.31 //y2=2.08
cc_1840 ( N_VDD_c_1035_p N_noxref_21_c_7660_n ) capacitor c=0.00453473f \
 //x=84.73 //y=7.4 //x2=63.815 //y2=5.2
cc_1841 ( N_VDD_c_1578_p N_noxref_21_c_7660_n ) capacitor c=4.48391e-19 \
 //x=63.375 //y=7.4 //x2=63.815 //y2=5.2
cc_1842 ( N_VDD_c_1720_p N_noxref_21_c_7660_n ) capacitor c=4.48377e-19 \
 //x=64.255 //y=7.4 //x2=63.815 //y2=5.2
cc_1843 ( N_VDD_M129_noxref_d N_noxref_21_c_7660_n ) capacitor c=0.0124506f \
 //x=63.315 //y=5.02 //x2=63.815 //y2=5.2
cc_1844 ( N_VDD_c_1027_n N_noxref_21_c_7664_n ) capacitor c=0.00985474f \
 //x=61.79 //y=7.4 //x2=63.105 //y2=5.2
cc_1845 ( N_VDD_M128_noxref_s N_noxref_21_c_7664_n ) capacitor c=0.087833f \
 //x=62.445 //y=5.02 //x2=63.105 //y2=5.2
cc_1846 ( N_VDD_c_1035_p N_noxref_21_c_7666_n ) capacitor c=0.00307195f \
 //x=84.73 //y=7.4 //x2=64.295 //y2=5.2
cc_1847 ( N_VDD_c_1720_p N_noxref_21_c_7666_n ) capacitor c=7.73167e-19 \
 //x=64.255 //y=7.4 //x2=64.295 //y2=5.2
cc_1848 ( N_VDD_M131_noxref_d N_noxref_21_c_7666_n ) capacitor c=0.0161518f \
 //x=64.195 //y=5.02 //x2=64.295 //y2=5.2
cc_1849 ( N_VDD_M132_noxref_s N_noxref_21_c_7666_n ) capacitor c=2.44532e-19 \
 //x=65.775 //y=5.02 //x2=64.295 //y2=5.2
cc_1850 ( N_VDD_c_1027_n N_noxref_21_c_7651_n ) capacitor c=0.00151618f \
 //x=61.79 //y=7.4 //x2=64.38 //y2=3.7
cc_1851 ( N_VDD_c_1028_n N_noxref_21_c_7651_n ) capacitor c=0.0441967f \
 //x=65.12 //y=7.4 //x2=64.38 //y2=3.7
cc_1852 ( N_VDD_c_1030_n N_noxref_21_c_7652_n ) capacitor c=8.34234e-19 \
 //x=73.26 //y=7.4 //x2=71.78 //y2=2.08
cc_1853 ( N_VDD_c_1746_p N_noxref_21_M120_noxref_g ) capacitor c=0.00675175f \
 //x=55.815 //y=7.4 //x2=55.24 //y2=6.02
cc_1854 ( N_VDD_M119_noxref_d N_noxref_21_M120_noxref_g ) capacitor \
 c=0.015318f //x=54.875 //y=5.02 //x2=55.24 //y2=6.02
cc_1855 ( N_VDD_c_1746_p N_noxref_21_M121_noxref_g ) capacitor c=0.00675379f \
 //x=55.815 //y=7.4 //x2=55.68 //y2=6.02
cc_1856 ( N_VDD_M121_noxref_d N_noxref_21_M121_noxref_g ) capacitor \
 c=0.0394719f //x=55.755 //y=5.02 //x2=55.68 //y2=6.02
cc_1857 ( N_VDD_c_1570_p N_noxref_21_M126_noxref_g ) capacitor c=0.00675175f \
 //x=60.625 //y=7.4 //x2=60.05 //y2=6.02
cc_1858 ( N_VDD_M125_noxref_d N_noxref_21_M126_noxref_g ) capacitor \
 c=0.015318f //x=59.685 //y=5.02 //x2=60.05 //y2=6.02
cc_1859 ( N_VDD_c_1570_p N_noxref_21_M127_noxref_g ) capacitor c=0.00675379f \
 //x=60.625 //y=7.4 //x2=60.49 //y2=6.02
cc_1860 ( N_VDD_M127_noxref_d N_noxref_21_M127_noxref_g ) capacitor \
 c=0.0394719f //x=60.565 //y=5.02 //x2=60.49 //y2=6.02
cc_1861 ( N_VDD_c_1884_p N_noxref_21_M140_noxref_g ) capacitor c=0.00675175f \
 //x=72.095 //y=7.4 //x2=71.52 //y2=6.02
cc_1862 ( N_VDD_M139_noxref_d N_noxref_21_M140_noxref_g ) capacitor \
 c=0.015318f //x=71.155 //y=5.02 //x2=71.52 //y2=6.02
cc_1863 ( N_VDD_c_1884_p N_noxref_21_M141_noxref_g ) capacitor c=0.00675379f \
 //x=72.095 //y=7.4 //x2=71.96 //y2=6.02
cc_1864 ( N_VDD_M141_noxref_d N_noxref_21_M141_noxref_g ) capacitor \
 c=0.0394719f //x=72.035 //y=5.02 //x2=71.96 //y2=6.02
cc_1865 ( N_VDD_c_1035_p N_noxref_21_M128_noxref_d ) capacitor c=0.00275225f \
 //x=84.73 //y=7.4 //x2=62.875 //y2=5.02
cc_1866 ( N_VDD_c_1578_p N_noxref_21_M128_noxref_d ) capacitor c=0.0140317f \
 //x=63.375 //y=7.4 //x2=62.875 //y2=5.02
cc_1867 ( N_VDD_c_1028_n N_noxref_21_M128_noxref_d ) capacitor c=6.94454e-19 \
 //x=65.12 //y=7.4 //x2=62.875 //y2=5.02
cc_1868 ( N_VDD_M129_noxref_d N_noxref_21_M128_noxref_d ) capacitor \
 c=0.0664752f //x=63.315 //y=5.02 //x2=62.875 //y2=5.02
cc_1869 ( N_VDD_c_1035_p N_noxref_21_M130_noxref_d ) capacitor c=0.00285083f \
 //x=84.73 //y=7.4 //x2=63.755 //y2=5.02
cc_1870 ( N_VDD_c_1720_p N_noxref_21_M130_noxref_d ) capacitor c=0.0140984f \
 //x=64.255 //y=7.4 //x2=63.755 //y2=5.02
cc_1871 ( N_VDD_c_1028_n N_noxref_21_M130_noxref_d ) capacitor c=0.0120541f \
 //x=65.12 //y=7.4 //x2=63.755 //y2=5.02
cc_1872 ( N_VDD_M128_noxref_s N_noxref_21_M130_noxref_d ) capacitor \
 c=0.00111971f //x=62.445 //y=5.02 //x2=63.755 //y2=5.02
cc_1873 ( N_VDD_M129_noxref_d N_noxref_21_M130_noxref_d ) capacitor \
 c=0.0664752f //x=63.315 //y=5.02 //x2=63.755 //y2=5.02
cc_1874 ( N_VDD_M131_noxref_d N_noxref_21_M130_noxref_d ) capacitor \
 c=0.0664752f //x=64.195 //y=5.02 //x2=63.755 //y2=5.02
cc_1875 ( N_VDD_M132_noxref_s N_noxref_21_M130_noxref_d ) capacitor \
 c=4.54516e-19 //x=65.775 //y=5.02 //x2=63.755 //y2=5.02
cc_1876 ( N_VDD_c_1035_p N_noxref_22_c_7969_n ) capacitor c=0.0206457f \
 //x=84.73 //y=7.4 //x2=77.255 //y2=5.21
cc_1877 ( N_VDD_c_1472_p N_noxref_22_c_7969_n ) capacitor c=0.00213763f \
 //x=75.725 //y=7.4 //x2=77.255 //y2=5.21
cc_1878 ( N_VDD_c_1901_p N_noxref_22_c_7969_n ) capacitor c=0.003172f \
 //x=76.42 //y=7.4 //x2=77.255 //y2=5.21
cc_1879 ( N_VDD_c_1902_p N_noxref_22_c_7969_n ) capacitor c=0.00424633f \
 //x=79.75 //y=7.4 //x2=77.255 //y2=5.21
cc_1880 ( N_VDD_c_1031_n N_noxref_22_c_7969_n ) capacitor c=0.0430305f \
 //x=76.59 //y=7.4 //x2=77.255 //y2=5.21
cc_1881 ( N_VDD_M145_noxref_d N_noxref_22_c_7969_n ) capacitor c=0.0197937f \
 //x=75.665 //y=5.025 //x2=77.255 //y2=5.21
cc_1882 ( N_VDD_c_1035_p N_noxref_22_c_7975_n ) capacitor c=0.00274812f \
 //x=84.73 //y=7.4 //x2=75.485 //y2=5.21
cc_1883 ( N_VDD_c_1472_p N_noxref_22_c_7975_n ) capacitor c=0.00107267f \
 //x=75.725 //y=7.4 //x2=75.485 //y2=5.21
cc_1884 ( N_VDD_c_1030_n N_noxref_22_c_7975_n ) capacitor c=2.89592e-19 \
 //x=73.26 //y=7.4 //x2=75.485 //y2=5.21
cc_1885 ( N_VDD_c_1031_n N_noxref_22_c_7975_n ) capacitor c=3.35418e-19 \
 //x=76.59 //y=7.4 //x2=75.485 //y2=5.21
cc_1886 ( N_VDD_M145_noxref_d N_noxref_22_c_7975_n ) capacitor c=6.02701e-19 \
 //x=75.665 //y=5.025 //x2=75.485 //y2=5.21
cc_1887 ( N_VDD_c_1035_p N_noxref_22_c_7980_n ) capacitor c=0.00453889f \
 //x=84.73 //y=7.4 //x2=75.285 //y2=5.21
cc_1888 ( N_VDD_c_1911_p N_noxref_22_c_7980_n ) capacitor c=4.52207e-19 \
 //x=74.845 //y=7.4 //x2=75.285 //y2=5.21
cc_1889 ( N_VDD_c_1472_p N_noxref_22_c_7980_n ) capacitor c=4.11408e-19 \
 //x=75.725 //y=7.4 //x2=75.285 //y2=5.21
cc_1890 ( N_VDD_M143_noxref_d N_noxref_22_c_7980_n ) capacitor c=0.0127968f \
 //x=74.785 //y=5.025 //x2=75.285 //y2=5.21
cc_1891 ( N_VDD_c_1030_n N_noxref_22_c_7984_n ) capacitor c=0.00914165f \
 //x=73.26 //y=7.4 //x2=74.575 //y2=5.21
cc_1892 ( N_VDD_M142_noxref_s N_noxref_22_c_7984_n ) capacitor c=0.0872987f \
 //x=73.915 //y=5.025 //x2=74.575 //y2=5.21
cc_1893 ( N_VDD_c_1030_n N_noxref_22_c_7986_n ) capacitor c=6.3991e-19 \
 //x=73.26 //y=7.4 //x2=75.37 //y2=5.295
cc_1894 ( N_VDD_c_1031_n N_noxref_22_c_7986_n ) capacitor c=0.00985441f \
 //x=76.59 //y=7.4 //x2=75.37 //y2=5.295
cc_1895 ( N_VDD_M145_noxref_d N_noxref_22_c_7986_n ) capacitor c=0.0873334f \
 //x=75.665 //y=5.025 //x2=75.37 //y2=5.295
cc_1896 ( N_VDD_c_1031_n N_noxref_22_c_7989_n ) capacitor c=0.0674112f \
 //x=76.59 //y=7.4 //x2=77.37 //y2=5.21
cc_1897 ( N_VDD_M145_noxref_d N_noxref_22_c_7989_n ) capacitor c=0.00235009f \
 //x=75.665 //y=5.025 //x2=77.37 //y2=5.21
cc_1898 ( N_VDD_c_1035_p N_noxref_22_c_7991_n ) capacitor c=0.0296174f \
 //x=84.73 //y=7.4 //x2=77.455 //y2=6.91
cc_1899 ( N_VDD_c_1902_p N_noxref_22_c_7991_n ) capacitor c=0.109938f \
 //x=79.75 //y=7.4 //x2=77.455 //y2=6.91
cc_1900 ( N_VDD_c_1035_p N_noxref_22_M142_noxref_d ) capacitor c=0.00291898f \
 //x=84.73 //y=7.4 //x2=74.345 //y2=5.025
cc_1901 ( N_VDD_c_1911_p N_noxref_22_M142_noxref_d ) capacitor c=0.0137097f \
 //x=74.845 //y=7.4 //x2=74.345 //y2=5.025
cc_1902 ( N_VDD_M143_noxref_d N_noxref_22_M142_noxref_d ) capacitor \
 c=0.067695f //x=74.785 //y=5.025 //x2=74.345 //y2=5.025
cc_1903 ( N_VDD_M145_noxref_d N_noxref_22_M142_noxref_d ) capacitor \
 c=0.00105738f //x=75.665 //y=5.025 //x2=74.345 //y2=5.025
cc_1904 ( N_VDD_c_1035_p N_noxref_22_M144_noxref_d ) capacitor c=0.00241371f \
 //x=84.73 //y=7.4 //x2=75.225 //y2=5.025
cc_1905 ( N_VDD_c_1472_p N_noxref_22_M144_noxref_d ) capacitor c=0.01268f \
 //x=75.725 //y=7.4 //x2=75.225 //y2=5.025
cc_1906 ( N_VDD_M142_noxref_s N_noxref_22_M144_noxref_d ) capacitor \
 c=0.00103189f //x=73.915 //y=5.025 //x2=75.225 //y2=5.025
cc_1907 ( N_VDD_M143_noxref_d N_noxref_22_M144_noxref_d ) capacitor \
 c=0.0653408f //x=74.785 //y=5.025 //x2=75.225 //y2=5.025
cc_1908 ( N_VDD_c_1031_n N_noxref_22_M147_noxref_d ) capacitor c=8.96067e-19 \
 //x=76.59 //y=7.4 //x2=78.105 //y2=5.025
cc_1909 ( N_VDD_c_1032_n N_noxref_22_M147_noxref_d ) capacitor c=8.88629e-19 \
 //x=79.92 //y=7.4 //x2=78.105 //y2=5.025
cc_1910 ( N_VDD_c_1032_n N_noxref_22_M149_noxref_d ) capacitor c=0.0575594f \
 //x=79.92 //y=7.4 //x2=78.985 //y2=5.025
cc_1911 ( N_VDD_c_1035_p N_noxref_23_c_8089_n ) capacitor c=0.031581f \
 //x=84.73 //y=7.4 //x2=72.405 //y2=4.44
cc_1912 ( N_VDD_c_1784_p N_noxref_23_c_8089_n ) capacitor c=0.00123284f \
 //x=70.335 //y=7.4 //x2=72.405 //y2=4.44
cc_1913 ( N_VDD_c_1029_n N_noxref_23_c_8089_n ) capacitor c=0.0249242f \
 //x=68.45 //y=7.4 //x2=72.405 //y2=4.44
cc_1914 ( N_VDD_c_1035_p N_noxref_23_c_8092_n ) capacitor c=0.00149097f \
 //x=84.73 //y=7.4 //x2=67.085 //y2=4.44
cc_1915 ( N_VDD_c_1035_p N_noxref_23_c_8093_n ) capacitor c=0.00963266f \
 //x=84.73 //y=7.4 //x2=73.885 //y2=4.44
cc_1916 ( N_VDD_c_1939_p N_noxref_23_c_8093_n ) capacitor c=0.00197825f \
 //x=73.09 //y=7.4 //x2=73.885 //y2=4.44
cc_1917 ( N_VDD_c_1940_p N_noxref_23_c_8093_n ) capacitor c=0.00196539f \
 //x=73.965 //y=7.4 //x2=73.885 //y2=4.44
cc_1918 ( N_VDD_c_1030_n N_noxref_23_c_8093_n ) capacitor c=0.0380101f \
 //x=73.26 //y=7.4 //x2=73.885 //y2=4.44
cc_1919 ( N_VDD_c_1035_p N_noxref_23_c_8097_n ) capacitor c=0.00193828f \
 //x=84.73 //y=7.4 //x2=72.635 //y2=4.44
cc_1920 ( N_VDD_c_1939_p N_noxref_23_c_8097_n ) capacitor c=6.06662e-19 \
 //x=73.09 //y=7.4 //x2=72.635 //y2=4.44
cc_1921 ( N_VDD_c_1030_n N_noxref_23_c_8097_n ) capacitor c=9.11674e-19 \
 //x=73.26 //y=7.4 //x2=72.635 //y2=4.44
cc_1922 ( N_VDD_c_1035_p N_noxref_23_c_8100_n ) capacitor c=0.014626f \
 //x=84.73 //y=7.4 //x2=77.585 //y2=4.44
cc_1923 ( N_VDD_c_1911_p N_noxref_23_c_8100_n ) capacitor c=0.00134165f \
 //x=74.845 //y=7.4 //x2=77.585 //y2=4.44
cc_1924 ( N_VDD_c_1031_n N_noxref_23_c_8100_n ) capacitor c=0.03415f //x=76.59 \
 //y=7.4 //x2=77.585 //y2=4.44
cc_1925 ( N_VDD_M142_noxref_s N_noxref_23_c_8100_n ) capacitor c=6.29527e-19 \
 //x=73.915 //y=5.025 //x2=77.585 //y2=4.44
cc_1926 ( N_VDD_M145_noxref_d N_noxref_23_c_8100_n ) capacitor c=0.0033086f \
 //x=75.665 //y=5.025 //x2=77.585 //y2=4.44
cc_1927 ( N_VDD_c_1035_p N_noxref_23_c_8105_n ) capacitor c=0.00140297f \
 //x=84.73 //y=7.4 //x2=74.115 //y2=4.44
cc_1928 ( N_VDD_c_1940_p N_noxref_23_c_8105_n ) capacitor c=3.1987e-19 \
 //x=73.965 //y=7.4 //x2=74.115 //y2=4.44
cc_1929 ( N_VDD_c_1030_n N_noxref_23_c_8105_n ) capacitor c=0.00100472f \
 //x=73.26 //y=7.4 //x2=74.115 //y2=4.44
cc_1930 ( N_VDD_M142_noxref_s N_noxref_23_c_8105_n ) capacitor c=0.00225389f \
 //x=73.915 //y=5.025 //x2=74.115 //y2=4.44
cc_1931 ( N_VDD_c_1028_n N_noxref_23_c_8060_n ) capacitor c=8.15787e-19 \
 //x=65.12 //y=7.4 //x2=66.97 //y2=2.08
cc_1932 ( N_VDD_c_1029_n N_noxref_23_c_8060_n ) capacitor c=4.99817e-19 \
 //x=68.45 //y=7.4 //x2=66.97 //y2=2.08
cc_1933 ( N_VDD_c_1035_p N_noxref_23_c_8111_n ) capacitor c=0.00444892f \
 //x=84.73 //y=7.4 //x2=70.775 //y2=5.155
cc_1934 ( N_VDD_c_1784_p N_noxref_23_c_8111_n ) capacitor c=4.31931e-19 \
 //x=70.335 //y=7.4 //x2=70.775 //y2=5.155
cc_1935 ( N_VDD_c_1855_p N_noxref_23_c_8111_n ) capacitor c=4.31931e-19 \
 //x=71.215 //y=7.4 //x2=70.775 //y2=5.155
cc_1936 ( N_VDD_M137_noxref_d N_noxref_23_c_8111_n ) capacitor c=0.0112985f \
 //x=70.275 //y=5.02 //x2=70.775 //y2=5.155
cc_1937 ( N_VDD_c_1029_n N_noxref_23_c_8115_n ) capacitor c=0.00863585f \
 //x=68.45 //y=7.4 //x2=70.065 //y2=5.155
cc_1938 ( N_VDD_M136_noxref_s N_noxref_23_c_8115_n ) capacitor c=0.0831083f \
 //x=69.405 //y=5.02 //x2=70.065 //y2=5.155
cc_1939 ( N_VDD_c_1035_p N_noxref_23_c_8117_n ) capacitor c=0.0044221f \
 //x=84.73 //y=7.4 //x2=71.655 //y2=5.155
cc_1940 ( N_VDD_c_1855_p N_noxref_23_c_8117_n ) capacitor c=4.31931e-19 \
 //x=71.215 //y=7.4 //x2=71.655 //y2=5.155
cc_1941 ( N_VDD_c_1884_p N_noxref_23_c_8117_n ) capacitor c=4.31931e-19 \
 //x=72.095 //y=7.4 //x2=71.655 //y2=5.155
cc_1942 ( N_VDD_M139_noxref_d N_noxref_23_c_8117_n ) capacitor c=0.0112985f \
 //x=71.155 //y=5.02 //x2=71.655 //y2=5.155
cc_1943 ( N_VDD_c_1035_p N_noxref_23_c_8121_n ) capacitor c=0.00434009f \
 //x=84.73 //y=7.4 //x2=72.435 //y2=5.155
cc_1944 ( N_VDD_c_1884_p N_noxref_23_c_8121_n ) capacitor c=7.46626e-19 \
 //x=72.095 //y=7.4 //x2=72.435 //y2=5.155
cc_1945 ( N_VDD_c_1939_p N_noxref_23_c_8121_n ) capacitor c=0.00198541f \
 //x=73.09 //y=7.4 //x2=72.435 //y2=5.155
cc_1946 ( N_VDD_M141_noxref_d N_noxref_23_c_8121_n ) capacitor c=0.0112985f \
 //x=72.035 //y=5.02 //x2=72.435 //y2=5.155
cc_1947 ( N_VDD_M142_noxref_s N_noxref_23_c_8121_n ) capacitor c=4.06494e-19 \
 //x=73.915 //y=5.025 //x2=72.435 //y2=5.155
cc_1948 ( N_VDD_c_1030_n N_noxref_23_c_8126_n ) capacitor c=0.0430788f \
 //x=73.26 //y=7.4 //x2=72.52 //y2=4.44
cc_1949 ( N_VDD_c_1035_p N_noxref_23_c_8063_n ) capacitor c=0.00142825f \
 //x=84.73 //y=7.4 //x2=74 //y2=2.08
cc_1950 ( N_VDD_c_1030_n N_noxref_23_c_8063_n ) capacitor c=0.0247009f \
 //x=73.26 //y=7.4 //x2=74 //y2=2.08
cc_1951 ( N_VDD_c_1031_n N_noxref_23_c_8063_n ) capacitor c=4.17679e-19 \
 //x=76.59 //y=7.4 //x2=74 //y2=2.08
cc_1952 ( N_VDD_M142_noxref_s N_noxref_23_c_8063_n ) capacitor c=0.0119799f \
 //x=73.915 //y=5.025 //x2=74 //y2=2.08
cc_1953 ( N_VDD_c_1031_n N_noxref_23_c_8066_n ) capacitor c=0.0131686f \
 //x=76.59 //y=7.4 //x2=77.7 //y2=2.08
cc_1954 ( N_VDD_c_1032_n N_noxref_23_c_8066_n ) capacitor c=0.00133861f \
 //x=79.92 //y=7.4 //x2=77.7 //y2=2.08
cc_1955 ( N_VDD_c_1793_p N_noxref_23_M134_noxref_g ) capacitor c=0.00673971f \
 //x=67.585 //y=7.4 //x2=67.01 //y2=6.02
cc_1956 ( N_VDD_M133_noxref_d N_noxref_23_M134_noxref_g ) capacitor \
 c=0.015318f //x=66.645 //y=5.02 //x2=67.01 //y2=6.02
cc_1957 ( N_VDD_c_1793_p N_noxref_23_M135_noxref_g ) capacitor c=0.00672952f \
 //x=67.585 //y=7.4 //x2=67.45 //y2=6.02
cc_1958 ( N_VDD_c_1029_n N_noxref_23_M135_noxref_g ) capacitor c=0.00839945f \
 //x=68.45 //y=7.4 //x2=67.45 //y2=6.02
cc_1959 ( N_VDD_M135_noxref_d N_noxref_23_M135_noxref_g ) capacitor \
 c=0.0430452f //x=67.525 //y=5.02 //x2=67.45 //y2=6.02
cc_1960 ( N_VDD_c_1911_p N_noxref_23_M142_noxref_g ) capacitor c=0.00754867f \
 //x=74.845 //y=7.4 //x2=74.27 //y2=6.025
cc_1961 ( N_VDD_c_1030_n N_noxref_23_M142_noxref_g ) capacitor c=0.00694765f \
 //x=73.26 //y=7.4 //x2=74.27 //y2=6.025
cc_1962 ( N_VDD_M142_noxref_s N_noxref_23_M142_noxref_g ) capacitor \
 c=0.0547553f //x=73.915 //y=5.025 //x2=74.27 //y2=6.025
cc_1963 ( N_VDD_c_1911_p N_noxref_23_M143_noxref_g ) capacitor c=0.00678153f \
 //x=74.845 //y=7.4 //x2=74.71 //y2=6.025
cc_1964 ( N_VDD_M143_noxref_d N_noxref_23_M143_noxref_g ) capacitor \
 c=0.015501f //x=74.785 //y=5.025 //x2=74.71 //y2=6.025
cc_1965 ( N_VDD_c_1902_p N_noxref_23_M146_noxref_g ) capacitor c=0.00513227f \
 //x=79.75 //y=7.4 //x2=77.59 //y2=6.025
cc_1966 ( N_VDD_c_1031_n N_noxref_23_M146_noxref_g ) capacitor c=0.00316281f \
 //x=76.59 //y=7.4 //x2=77.59 //y2=6.025
cc_1967 ( N_VDD_c_1902_p N_noxref_23_M147_noxref_g ) capacitor c=0.00512552f \
 //x=79.75 //y=7.4 //x2=78.03 //y2=6.025
cc_1968 ( N_VDD_c_1030_n N_noxref_23_c_8146_n ) capacitor c=0.0110236f \
 //x=73.26 //y=7.4 //x2=74.345 //y2=4.795
cc_1969 ( N_VDD_M142_noxref_s N_noxref_23_c_8146_n ) capacitor c=0.00628155f \
 //x=73.915 //y=5.025 //x2=74.345 //y2=4.795
cc_1970 ( N_VDD_c_1031_n N_noxref_23_c_8148_n ) capacitor c=0.0115029f \
 //x=76.59 //y=7.4 //x2=77.7 //y2=4.705
cc_1971 ( N_VDD_c_1035_p N_noxref_23_M136_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=69.835 //y2=5.02
cc_1972 ( N_VDD_c_1784_p N_noxref_23_M136_noxref_d ) capacitor c=0.014035f \
 //x=70.335 //y=7.4 //x2=69.835 //y2=5.02
cc_1973 ( N_VDD_M137_noxref_d N_noxref_23_M136_noxref_d ) capacitor \
 c=0.0664752f //x=70.275 //y=5.02 //x2=69.835 //y2=5.02
cc_1974 ( N_VDD_c_1035_p N_noxref_23_M138_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=70.715 //y2=5.02
cc_1975 ( N_VDD_c_1855_p N_noxref_23_M138_noxref_d ) capacitor c=0.014035f \
 //x=71.215 //y=7.4 //x2=70.715 //y2=5.02
cc_1976 ( N_VDD_c_1030_n N_noxref_23_M138_noxref_d ) capacitor c=4.9285e-19 \
 //x=73.26 //y=7.4 //x2=70.715 //y2=5.02
cc_1977 ( N_VDD_M136_noxref_s N_noxref_23_M138_noxref_d ) capacitor \
 c=0.00130656f //x=69.405 //y=5.02 //x2=70.715 //y2=5.02
cc_1978 ( N_VDD_M137_noxref_d N_noxref_23_M138_noxref_d ) capacitor \
 c=0.0664752f //x=70.275 //y=5.02 //x2=70.715 //y2=5.02
cc_1979 ( N_VDD_M139_noxref_d N_noxref_23_M138_noxref_d ) capacitor \
 c=0.0664752f //x=71.155 //y=5.02 //x2=70.715 //y2=5.02
cc_1980 ( N_VDD_c_1035_p N_noxref_23_M140_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=71.595 //y2=5.02
cc_1981 ( N_VDD_c_1884_p N_noxref_23_M140_noxref_d ) capacitor c=0.0137384f \
 //x=72.095 //y=7.4 //x2=71.595 //y2=5.02
cc_1982 ( N_VDD_c_1030_n N_noxref_23_M140_noxref_d ) capacitor c=0.00939849f \
 //x=73.26 //y=7.4 //x2=71.595 //y2=5.02
cc_1983 ( N_VDD_M139_noxref_d N_noxref_23_M140_noxref_d ) capacitor \
 c=0.0664752f //x=71.155 //y=5.02 //x2=71.595 //y2=5.02
cc_1984 ( N_VDD_M141_noxref_d N_noxref_23_M140_noxref_d ) capacitor \
 c=0.0664752f //x=72.035 //y=5.02 //x2=71.595 //y2=5.02
cc_1985 ( N_VDD_M142_noxref_s N_noxref_23_M140_noxref_d ) capacitor \
 c=4.52683e-19 //x=73.915 //y=5.025 //x2=71.595 //y2=5.02
cc_1986 ( N_VDD_c_1018_n N_noxref_24_c_8424_n ) capacitor c=0.0045786f \
 //x=24.42 //y=7.4 //x2=79.065 //y2=3.33
cc_1987 ( N_VDD_c_1024_n N_noxref_24_c_8424_n ) capacitor c=0.0045786f \
 //x=48.84 //y=7.4 //x2=79.065 //y2=3.33
cc_1988 ( N_VDD_c_1030_n N_noxref_24_c_8424_n ) capacitor c=0.0045786f \
 //x=73.26 //y=7.4 //x2=79.065 //y2=3.33
cc_1989 ( N_VDD_c_1016_n N_noxref_24_c_8428_n ) capacitor c=6.20324e-19 \
 //x=16.28 //y=7.4 //x2=18.13 //y2=2.08
cc_1990 ( N_VDD_c_1017_n N_noxref_24_c_8428_n ) capacitor c=4.33828e-19 \
 //x=19.61 //y=7.4 //x2=18.13 //y2=2.08
cc_1991 ( N_VDD_c_1035_p N_noxref_24_c_8451_n ) capacitor c=0.00444892f \
 //x=84.73 //y=7.4 //x2=21.935 //y2=5.155
cc_1992 ( N_VDD_c_1186_p N_noxref_24_c_8451_n ) capacitor c=4.31931e-19 \
 //x=21.495 //y=7.4 //x2=21.935 //y2=5.155
cc_1993 ( N_VDD_c_1839_p N_noxref_24_c_8451_n ) capacitor c=4.31931e-19 \
 //x=22.375 //y=7.4 //x2=21.935 //y2=5.155
cc_1994 ( N_VDD_M77_noxref_d N_noxref_24_c_8451_n ) capacitor c=0.0112985f \
 //x=21.435 //y=5.02 //x2=21.935 //y2=5.155
cc_1995 ( N_VDD_c_1017_n N_noxref_24_c_8455_n ) capacitor c=0.00863585f \
 //x=19.61 //y=7.4 //x2=21.225 //y2=5.155
cc_1996 ( N_VDD_M76_noxref_s N_noxref_24_c_8455_n ) capacitor c=0.0831083f \
 //x=20.565 //y=5.02 //x2=21.225 //y2=5.155
cc_1997 ( N_VDD_c_1035_p N_noxref_24_c_8457_n ) capacitor c=0.0044221f \
 //x=84.73 //y=7.4 //x2=22.815 //y2=5.155
cc_1998 ( N_VDD_c_1839_p N_noxref_24_c_8457_n ) capacitor c=4.31931e-19 \
 //x=22.375 //y=7.4 //x2=22.815 //y2=5.155
cc_1999 ( N_VDD_c_1226_p N_noxref_24_c_8457_n ) capacitor c=4.31931e-19 \
 //x=23.255 //y=7.4 //x2=22.815 //y2=5.155
cc_2000 ( N_VDD_M79_noxref_d N_noxref_24_c_8457_n ) capacitor c=0.0112985f \
 //x=22.315 //y=5.02 //x2=22.815 //y2=5.155
cc_2001 ( N_VDD_c_1035_p N_noxref_24_c_8461_n ) capacitor c=0.00434174f \
 //x=84.73 //y=7.4 //x2=23.595 //y2=5.155
cc_2002 ( N_VDD_c_1226_p N_noxref_24_c_8461_n ) capacitor c=7.46626e-19 \
 //x=23.255 //y=7.4 //x2=23.595 //y2=5.155
cc_2003 ( N_VDD_c_1619_p N_noxref_24_c_8461_n ) capacitor c=0.00198565f \
 //x=24.25 //y=7.4 //x2=23.595 //y2=5.155
cc_2004 ( N_VDD_M81_noxref_d N_noxref_24_c_8461_n ) capacitor c=0.0112985f \
 //x=23.195 //y=5.02 //x2=23.595 //y2=5.155
cc_2005 ( N_VDD_c_1018_n N_noxref_24_c_8465_n ) capacitor c=0.0433018f \
 //x=24.42 //y=7.4 //x2=23.68 //y2=3.33
cc_2006 ( N_VDD_c_1031_n N_noxref_24_c_8431_n ) capacitor c=7.57423e-19 \
 //x=76.59 //y=7.4 //x2=79.18 //y2=2.08
cc_2007 ( N_VDD_c_1032_n N_noxref_24_c_8431_n ) capacitor c=0.0263215f \
 //x=79.92 //y=7.4 //x2=79.18 //y2=2.08
cc_2008 ( N_VDD_c_1032_n N_noxref_24_c_8433_n ) capacitor c=0.0263871f \
 //x=79.92 //y=7.4 //x2=80.66 //y2=2.08
cc_2009 ( N_VDD_c_1174_p N_noxref_24_M74_noxref_g ) capacitor c=0.00673971f \
 //x=18.745 //y=7.4 //x2=18.17 //y2=6.02
cc_2010 ( N_VDD_M73_noxref_d N_noxref_24_M74_noxref_g ) capacitor c=0.015318f \
 //x=17.805 //y=5.02 //x2=18.17 //y2=6.02
cc_2011 ( N_VDD_c_1174_p N_noxref_24_M75_noxref_g ) capacitor c=0.00672952f \
 //x=18.745 //y=7.4 //x2=18.61 //y2=6.02
cc_2012 ( N_VDD_c_1017_n N_noxref_24_M75_noxref_g ) capacitor c=0.00928743f \
 //x=19.61 //y=7.4 //x2=18.61 //y2=6.02
cc_2013 ( N_VDD_M75_noxref_d N_noxref_24_M75_noxref_g ) capacitor c=0.0430452f \
 //x=18.685 //y=5.02 //x2=18.61 //y2=6.02
cc_2014 ( N_VDD_c_1902_p N_noxref_24_M148_noxref_g ) capacitor c=0.00512552f \
 //x=79.75 //y=7.4 //x2=78.47 //y2=6.025
cc_2015 ( N_VDD_c_1902_p N_noxref_24_M149_noxref_g ) capacitor c=0.00512552f \
 //x=79.75 //y=7.4 //x2=78.91 //y2=6.025
cc_2016 ( N_VDD_c_1032_n N_noxref_24_M149_noxref_g ) capacitor c=0.010355f \
 //x=79.92 //y=7.4 //x2=78.91 //y2=6.025
cc_2017 ( N_VDD_c_1441_p N_noxref_24_M150_noxref_g ) capacitor c=0.00512552f \
 //x=83.08 //y=7.4 //x2=80.93 //y2=6.025
cc_2018 ( N_VDD_c_1032_n N_noxref_24_M150_noxref_g ) capacitor c=0.00767856f \
 //x=79.92 //y=7.4 //x2=80.93 //y2=6.025
cc_2019 ( N_VDD_c_1441_p N_noxref_24_M151_noxref_g ) capacitor c=0.00512552f \
 //x=83.08 //y=7.4 //x2=81.37 //y2=6.025
cc_2020 ( N_VDD_c_1032_n N_noxref_24_c_8480_n ) capacitor c=0.00803198f \
 //x=79.92 //y=7.4 //x2=78.91 //y2=4.87
cc_2021 ( N_VDD_c_1032_n N_noxref_24_c_8481_n ) capacitor c=0.00803198f \
 //x=79.92 //y=7.4 //x2=81.005 //y2=4.795
cc_2022 ( N_VDD_c_1035_p N_noxref_24_M76_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=20.995 //y2=5.02
cc_2023 ( N_VDD_c_1186_p N_noxref_24_M76_noxref_d ) capacitor c=0.014035f \
 //x=21.495 //y=7.4 //x2=20.995 //y2=5.02
cc_2024 ( N_VDD_M77_noxref_d N_noxref_24_M76_noxref_d ) capacitor c=0.0664752f \
 //x=21.435 //y=5.02 //x2=20.995 //y2=5.02
cc_2025 ( N_VDD_c_1035_p N_noxref_24_M78_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=21.875 //y2=5.02
cc_2026 ( N_VDD_c_1839_p N_noxref_24_M78_noxref_d ) capacitor c=0.014035f \
 //x=22.375 //y=7.4 //x2=21.875 //y2=5.02
cc_2027 ( N_VDD_c_1018_n N_noxref_24_M78_noxref_d ) capacitor c=4.9285e-19 \
 //x=24.42 //y=7.4 //x2=21.875 //y2=5.02
cc_2028 ( N_VDD_M76_noxref_s N_noxref_24_M78_noxref_d ) capacitor \
 c=0.00130656f //x=20.565 //y=5.02 //x2=21.875 //y2=5.02
cc_2029 ( N_VDD_M77_noxref_d N_noxref_24_M78_noxref_d ) capacitor c=0.0664752f \
 //x=21.435 //y=5.02 //x2=21.875 //y2=5.02
cc_2030 ( N_VDD_M79_noxref_d N_noxref_24_M78_noxref_d ) capacitor c=0.0664752f \
 //x=22.315 //y=5.02 //x2=21.875 //y2=5.02
cc_2031 ( N_VDD_c_1035_p N_noxref_24_M80_noxref_d ) capacitor c=0.00275235f \
 //x=84.73 //y=7.4 //x2=22.755 //y2=5.02
cc_2032 ( N_VDD_c_1226_p N_noxref_24_M80_noxref_d ) capacitor c=0.0137384f \
 //x=23.255 //y=7.4 //x2=22.755 //y2=5.02
cc_2033 ( N_VDD_c_1018_n N_noxref_24_M80_noxref_d ) capacitor c=0.00939849f \
 //x=24.42 //y=7.4 //x2=22.755 //y2=5.02
cc_2034 ( N_VDD_M79_noxref_d N_noxref_24_M80_noxref_d ) capacitor c=0.0664752f \
 //x=22.315 //y=5.02 //x2=22.755 //y2=5.02
cc_2035 ( N_VDD_M81_noxref_d N_noxref_24_M80_noxref_d ) capacitor c=0.0664752f \
 //x=23.195 //y=5.02 //x2=22.755 //y2=5.02
cc_2036 ( N_VDD_M82_noxref_s N_noxref_24_M80_noxref_d ) capacitor \
 c=4.52683e-19 //x=25.075 //y=5.02 //x2=22.755 //y2=5.02
cc_2037 ( N_VDD_c_1035_p N_noxref_25_c_8898_n ) capacitor c=0.0212729f \
 //x=84.73 //y=7.4 //x2=80.595 //y2=5.21
cc_2038 ( N_VDD_c_1902_p N_noxref_25_c_8898_n ) capacitor c=0.00386143f \
 //x=79.75 //y=7.4 //x2=80.595 //y2=5.21
cc_2039 ( N_VDD_c_1441_p N_noxref_25_c_8898_n ) capacitor c=0.00403412f \
 //x=83.08 //y=7.4 //x2=80.595 //y2=5.21
cc_2040 ( N_VDD_c_1032_n N_noxref_25_c_8898_n ) capacitor c=0.0473381f \
 //x=79.92 //y=7.4 //x2=80.595 //y2=5.21
cc_2041 ( N_VDD_c_1035_p N_noxref_25_c_8902_n ) capacitor c=0.00264311f \
 //x=84.73 //y=7.4 //x2=78.805 //y2=5.21
cc_2042 ( N_VDD_c_1032_n N_noxref_25_c_8902_n ) capacitor c=6.67754e-19 \
 //x=79.92 //y=7.4 //x2=78.805 //y2=5.21
cc_2043 ( N_VDD_c_1031_n N_noxref_25_c_8904_n ) capacitor c=0.00662411f \
 //x=76.59 //y=7.4 //x2=77.895 //y2=5.21
cc_2044 ( N_VDD_c_1032_n N_noxref_25_c_8905_n ) capacitor c=0.00999961f \
 //x=79.92 //y=7.4 //x2=78.69 //y2=5.295
cc_2045 ( N_VDD_c_1032_n N_noxref_25_c_8906_n ) capacitor c=0.0664301f \
 //x=79.92 //y=7.4 //x2=80.71 //y2=5.21
cc_2046 ( N_VDD_c_1033_n N_noxref_25_c_8906_n ) capacitor c=6.48751e-19 \
 //x=83.25 //y=7.4 //x2=80.71 //y2=5.21
cc_2047 ( N_VDD_c_1035_p N_noxref_25_c_8908_n ) capacitor c=0.0387208f \
 //x=84.73 //y=7.4 //x2=80.795 //y2=6.91
cc_2048 ( N_VDD_c_1441_p N_noxref_25_c_8908_n ) capacitor c=0.108798f \
 //x=83.08 //y=7.4 //x2=80.795 //y2=6.91
cc_2049 ( N_VDD_c_1032_n N_noxref_25_M151_noxref_d ) capacitor c=8.88629e-19 \
 //x=79.92 //y=7.4 //x2=81.445 //y2=5.025
cc_2050 ( N_VDD_c_1033_n N_noxref_25_M151_noxref_d ) capacitor c=8.96067e-19 \
 //x=83.25 //y=7.4 //x2=81.445 //y2=5.025
cc_2051 ( N_VDD_c_1033_n N_noxref_25_M153_noxref_d ) capacitor c=0.0521707f \
 //x=83.25 //y=7.4 //x2=82.325 //y2=5.025
cc_2052 ( N_VDD_M154_noxref_s N_noxref_25_M153_noxref_d ) capacitor \
 c=0.00227726f //x=83.79 //y=5.02 //x2=82.325 //y2=5.025
cc_2053 ( N_VDD_c_1035_p N_noxref_26_c_9004_n ) capacitor c=0.010492f \
 //x=84.73 //y=7.4 //x2=83.875 //y2=4.07
cc_2054 ( N_VDD_c_1441_p N_noxref_26_c_9004_n ) capacitor c=0.00161566f \
 //x=83.08 //y=7.4 //x2=83.875 //y2=4.07
cc_2055 ( N_VDD_c_2078_p N_noxref_26_c_9004_n ) capacitor c=0.00128378f \
 //x=83.84 //y=7.4 //x2=83.875 //y2=4.07
cc_2056 ( N_VDD_c_2079_p N_noxref_26_c_9004_n ) capacitor c=2.49117e-19 \
 //x=84.72 //y=7.4 //x2=83.875 //y2=4.07
cc_2057 ( N_VDD_c_1033_n N_noxref_26_c_9004_n ) capacitor c=0.0302435f \
 //x=83.25 //y=7.4 //x2=83.875 //y2=4.07
cc_2058 ( N_VDD_M154_noxref_s N_noxref_26_c_9004_n ) capacitor c=0.00194099f \
 //x=83.79 //y=5.02 //x2=83.875 //y2=4.07
cc_2059 ( N_VDD_c_1035_p N_noxref_26_c_9007_n ) capacitor c=0.00178785f \
 //x=84.73 //y=7.4 //x2=82.625 //y2=4.07
cc_2060 ( N_VDD_c_1441_p N_noxref_26_c_9007_n ) capacitor c=2.6378e-19 \
 //x=83.08 //y=7.4 //x2=82.625 //y2=4.07
cc_2061 ( N_VDD_c_1033_n N_noxref_26_c_9007_n ) capacitor c=4.55837e-19 \
 //x=83.25 //y=7.4 //x2=82.625 //y2=4.07
cc_2062 ( N_VDD_c_1032_n N_noxref_26_c_9045_n ) capacitor c=0.00660621f \
 //x=79.92 //y=7.4 //x2=81.235 //y2=5.21
cc_2063 ( N_VDD_c_1035_p N_noxref_26_c_9046_n ) capacitor c=0.0017748f \
 //x=84.73 //y=7.4 //x2=82.425 //y2=5.21
cc_2064 ( N_VDD_c_1441_p N_noxref_26_c_9046_n ) capacitor c=0.00139502f \
 //x=83.08 //y=7.4 //x2=82.425 //y2=5.21
cc_2065 ( N_VDD_M154_noxref_s N_noxref_26_c_9046_n ) capacitor c=3.59303e-19 \
 //x=83.79 //y=5.02 //x2=82.425 //y2=5.21
cc_2066 ( N_VDD_c_1032_n N_noxref_26_c_9010_n ) capacitor c=0.00147633f \
 //x=79.92 //y=7.4 //x2=82.51 //y2=4.07
cc_2067 ( N_VDD_c_1033_n N_noxref_26_c_9010_n ) capacitor c=0.0460801f \
 //x=83.25 //y=7.4 //x2=82.51 //y2=4.07
cc_2068 ( N_VDD_c_1035_p N_noxref_26_c_9011_n ) capacitor c=0.00157744f \
 //x=84.73 //y=7.4 //x2=83.99 //y2=2.085
cc_2069 ( N_VDD_c_1033_n N_noxref_26_c_9011_n ) capacitor c=0.0268729f \
 //x=83.25 //y=7.4 //x2=83.99 //y2=2.085
cc_2070 ( N_VDD_c_1034_n N_noxref_26_c_9011_n ) capacitor c=0.00150056f \
 //x=84.73 //y=7.4 //x2=83.99 //y2=2.085
cc_2071 ( N_VDD_M154_noxref_s N_noxref_26_c_9011_n ) capacitor c=0.00896093f \
 //x=83.79 //y=5.02 //x2=83.99 //y2=2.085
cc_2072 ( N_VDD_c_2079_p N_noxref_26_M154_noxref_g ) capacitor c=0.00748034f \
 //x=84.72 //y=7.4 //x2=84.145 //y2=6.02
cc_2073 ( N_VDD_c_1033_n N_noxref_26_M154_noxref_g ) capacitor c=0.00952235f \
 //x=83.25 //y=7.4 //x2=84.145 //y2=6.02
cc_2074 ( N_VDD_M154_noxref_s N_noxref_26_M154_noxref_g ) capacitor \
 c=0.0528676f //x=83.79 //y=5.02 //x2=84.145 //y2=6.02
cc_2075 ( N_VDD_c_2079_p N_noxref_26_M155_noxref_g ) capacitor c=0.00697478f \
 //x=84.72 //y=7.4 //x2=84.585 //y2=6.02
cc_2076 ( N_VDD_M155_noxref_d N_noxref_26_M155_noxref_g ) capacitor \
 c=0.0528676f //x=84.66 //y=5.02 //x2=84.585 //y2=6.02
cc_2077 ( N_VDD_c_1034_n N_noxref_26_c_9060_n ) capacitor c=0.0287802f \
 //x=84.73 //y=7.4 //x2=84.51 //y2=4.79
cc_2078 ( N_VDD_c_1033_n N_noxref_26_c_9061_n ) capacitor c=0.011132f \
 //x=83.25 //y=7.4 //x2=84.22 //y2=4.79
cc_2079 ( N_VDD_M154_noxref_s N_noxref_26_c_9061_n ) capacitor c=0.00524527f \
 //x=83.79 //y=5.02 //x2=84.22 //y2=4.79
cc_2080 ( N_VDD_c_1033_n N_noxref_26_M150_noxref_d ) capacitor c=6.67979e-19 \
 //x=83.25 //y=7.4 //x2=81.005 //y2=5.025
cc_2081 ( N_VDD_c_1033_n N_noxref_26_M152_noxref_d ) capacitor c=0.00965467f \
 //x=83.25 //y=7.4 //x2=81.885 //y2=5.025
cc_2082 ( N_VDD_M154_noxref_s N_noxref_26_M152_noxref_d ) capacitor \
 c=5.3724e-19 //x=83.79 //y=5.02 //x2=81.885 //y2=5.025
cc_2083 ( N_VDD_c_1033_n Q ) capacitor c=5.49291e-19 //x=83.25 //y=7.4 \
 //x2=84.73 //y2=2.22
cc_2084 ( N_VDD_c_1034_n Q ) capacitor c=0.0230793f //x=84.73 //y=7.4 \
 //x2=84.73 //y2=2.22
cc_2085 ( N_VDD_c_1035_p N_Q_c_10794_n ) capacitor c=0.00190861f //x=84.73 \
 //y=7.4 //x2=84.645 //y2=4.58
cc_2086 ( N_VDD_c_2079_p N_Q_c_10794_n ) capacitor c=8.8179e-19 //x=84.72 \
 //y=7.4 //x2=84.645 //y2=4.58
cc_2087 ( N_VDD_M155_noxref_d N_Q_c_10794_n ) capacitor c=0.00641434f \
 //x=84.66 //y=5.02 //x2=84.645 //y2=4.58
cc_2088 ( N_VDD_c_1033_n N_Q_c_10797_n ) capacitor c=0.017572f //x=83.25 \
 //y=7.4 //x2=84.45 //y2=4.58
cc_2089 ( N_VDD_c_1035_p N_Q_M154_noxref_d ) capacitor c=0.00708604f //x=84.73 \
 //y=7.4 //x2=84.22 //y2=5.02
cc_2090 ( N_VDD_c_2079_p N_Q_M154_noxref_d ) capacitor c=0.0139004f //x=84.72 \
 //y=7.4 //x2=84.22 //y2=5.02
cc_2091 ( N_VDD_c_1034_n N_Q_M154_noxref_d ) capacitor c=0.0205533f //x=84.73 \
 //y=7.4 //x2=84.22 //y2=5.02
cc_2092 ( N_VDD_M154_noxref_s N_Q_M154_noxref_d ) capacitor c=0.0843065f \
 //x=83.79 //y=5.02 //x2=84.22 //y2=5.02
cc_2093 ( N_VDD_M155_noxref_d N_Q_M154_noxref_d ) capacitor c=0.0832641f \
 //x=84.66 //y=5.02 //x2=84.22 //y2=5.02
cc_2094 ( N_noxref_3_c_2123_n N_noxref_4_c_2362_n ) capacitor c=0.00564994f \
 //x=9.135 //y=2.59 //x2=12.325 //y2=2.59
cc_2095 ( N_noxref_3_M63_noxref_g N_noxref_4_c_2377_n ) capacitor c=0.0168349f \
 //x=9.89 //y=6.02 //x2=10.465 //y2=5.155
cc_2096 ( N_noxref_3_M62_noxref_g N_noxref_4_c_2381_n ) capacitor c=0.0213876f \
 //x=9.45 //y=6.02 //x2=9.755 //y2=5.155
cc_2097 ( N_noxref_3_c_2200_p N_noxref_4_c_2381_n ) capacitor c=0.00428486f \
 //x=9.815 //y=4.79 //x2=9.755 //y2=5.155
cc_2098 ( N_noxref_3_M63_noxref_g N_noxref_4_M62_noxref_d ) capacitor \
 c=0.0180032f //x=9.89 //y=6.02 //x2=9.525 //y2=5.02
cc_2099 ( N_noxref_3_c_2117_n N_noxref_5_c_2540_n ) capacitor c=0.0043123f \
 //x=4.295 //y=2.59 //x2=7.28 //y2=4.07
cc_2100 ( N_noxref_3_c_2121_n N_noxref_5_c_2540_n ) capacitor c=5.62763e-19 \
 //x=2.705 //y=2.59 //x2=7.28 //y2=4.07
cc_2101 ( N_noxref_3_c_2127_n N_noxref_5_c_2540_n ) capacitor c=0.0121673f \
 //x=4.705 //y=2.59 //x2=7.28 //y2=4.07
cc_2102 ( N_noxref_3_c_2157_n N_noxref_5_c_2540_n ) capacitor c=0.0132304f \
 //x=2.025 //y=5.2 //x2=7.28 //y2=4.07
cc_2103 ( N_noxref_3_c_2130_n N_noxref_5_c_2540_n ) capacitor c=0.0270562f \
 //x=2.59 //y=2.59 //x2=7.28 //y2=4.07
cc_2104 ( N_noxref_3_c_2132_n N_noxref_5_c_2540_n ) capacitor c=0.027299f \
 //x=4.44 //y=2.08 //x2=7.28 //y2=4.07
cc_2105 ( N_noxref_3_c_2182_n N_noxref_5_c_2540_n ) capacitor c=0.0116469f \
 //x=4.715 //y=4.79 //x2=7.28 //y2=4.07
cc_2106 ( N_noxref_3_c_2157_n N_noxref_5_c_2547_n ) capacitor c=0.00204264f \
 //x=2.025 //y=5.2 //x2=1.965 //y2=4.07
cc_2107 ( N_noxref_3_c_2130_n N_noxref_5_c_2547_n ) capacitor c=0.00179385f \
 //x=2.59 //y=2.59 //x2=1.965 //y2=4.07
cc_2108 ( N_noxref_3_c_2133_n N_noxref_5_c_2548_n ) capacitor c=0.0194977f \
 //x=9.25 //y=2.08 //x2=17.275 //y2=4.07
cc_2109 ( N_noxref_3_c_2133_n N_noxref_5_c_2551_n ) capacitor c=3.49381e-19 \
 //x=9.25 //y=2.08 //x2=7.51 //y2=4.07
cc_2110 ( N_noxref_3_c_2157_n N_noxref_5_c_2608_n ) capacitor c=0.0129205f \
 //x=2.025 //y=5.2 //x2=1.85 //y2=4.535
cc_2111 ( N_noxref_3_c_2130_n N_noxref_5_c_2608_n ) capacitor c=0.0101115f \
 //x=2.59 //y=2.59 //x2=1.85 //y2=4.535
cc_2112 ( N_noxref_3_c_2121_n N_noxref_5_c_2525_n ) capacitor c=0.00691549f \
 //x=2.705 //y=2.59 //x2=1.85 //y2=2.08
cc_2113 ( N_noxref_3_c_2130_n N_noxref_5_c_2525_n ) capacitor c=0.0760197f \
 //x=2.59 //y=2.59 //x2=1.85 //y2=2.08
cc_2114 ( N_noxref_3_c_2132_n N_noxref_5_c_2525_n ) capacitor c=8.08904e-19 \
 //x=4.44 //y=2.08 //x2=1.85 //y2=2.08
cc_2115 ( N_noxref_3_M57_noxref_g N_noxref_5_c_2554_n ) capacitor c=0.0178794f \
 //x=5.08 //y=6.02 //x2=5.655 //y2=5.155
cc_2116 ( N_noxref_3_c_2130_n N_noxref_5_c_2558_n ) capacitor c=2.97874e-19 \
 //x=2.59 //y=2.59 //x2=4.945 //y2=5.155
cc_2117 ( N_noxref_3_M56_noxref_g N_noxref_5_c_2558_n ) capacitor c=0.0213876f \
 //x=4.64 //y=6.02 //x2=4.945 //y2=5.155
cc_2118 ( N_noxref_3_c_2221_p N_noxref_5_c_2558_n ) capacitor c=0.00429591f \
 //x=5.005 //y=4.79 //x2=4.945 //y2=5.155
cc_2119 ( N_noxref_3_c_2123_n N_noxref_5_c_2617_n ) capacitor c=0.011558f \
 //x=9.135 //y=2.59 //x2=7 //y2=1.665
cc_2120 ( N_noxref_3_c_2123_n N_noxref_5_c_2618_n ) capacitor c=0.0209737f \
 //x=9.135 //y=2.59 //x2=7.397 //y2=3.905
cc_2121 ( N_noxref_3_c_2133_n N_noxref_5_c_2618_n ) capacitor c=0.0130551f \
 //x=9.25 //y=2.08 //x2=7.397 //y2=3.905
cc_2122 ( N_noxref_3_c_2157_n N_noxref_5_M54_noxref_g ) capacitor c=0.0166421f \
 //x=2.025 //y=5.2 //x2=1.89 //y2=6.02
cc_2123 ( N_noxref_3_M54_noxref_d N_noxref_5_M54_noxref_g ) capacitor \
 c=0.0173476f //x=1.965 //y=5.02 //x2=1.89 //y2=6.02
cc_2124 ( N_noxref_3_c_2163_n N_noxref_5_M55_noxref_g ) capacitor c=0.0199348f \
 //x=2.505 //y=5.2 //x2=2.33 //y2=6.02
cc_2125 ( N_noxref_3_M54_noxref_d N_noxref_5_M55_noxref_g ) capacitor \
 c=0.0179769f //x=1.965 //y=5.02 //x2=2.33 //y2=6.02
cc_2126 ( N_noxref_3_M1_noxref_d N_noxref_5_c_2624_n ) capacitor c=0.00217566f \
 //x=1.96 //y=0.905 //x2=1.885 //y2=0.905
cc_2127 ( N_noxref_3_M1_noxref_d N_noxref_5_c_2625_n ) capacitor c=0.0034598f \
 //x=1.96 //y=0.905 //x2=1.885 //y2=1.25
cc_2128 ( N_noxref_3_M1_noxref_d N_noxref_5_c_2626_n ) capacitor c=0.0065582f \
 //x=1.96 //y=0.905 //x2=1.885 //y2=1.56
cc_2129 ( N_noxref_3_c_2130_n N_noxref_5_c_2627_n ) capacitor c=0.0142673f \
 //x=2.59 //y=2.59 //x2=2.255 //y2=4.79
cc_2130 ( N_noxref_3_c_2233_p N_noxref_5_c_2627_n ) capacitor c=0.00408717f \
 //x=2.11 //y=5.2 //x2=2.255 //y2=4.79
cc_2131 ( N_noxref_3_M1_noxref_d N_noxref_5_c_2629_n ) capacitor c=0.00241102f \
 //x=1.96 //y=0.905 //x2=2.26 //y2=0.75
cc_2132 ( N_noxref_3_c_2129_n N_noxref_5_c_2630_n ) capacitor c=0.00359704f \
 //x=2.505 //y=1.655 //x2=2.26 //y2=1.405
cc_2133 ( N_noxref_3_M1_noxref_d N_noxref_5_c_2630_n ) capacitor c=0.0138845f \
 //x=1.96 //y=0.905 //x2=2.26 //y2=1.405
cc_2134 ( N_noxref_3_M1_noxref_d N_noxref_5_c_2632_n ) capacitor c=0.00132245f \
 //x=1.96 //y=0.905 //x2=2.415 //y2=0.905
cc_2135 ( N_noxref_3_c_2129_n N_noxref_5_c_2633_n ) capacitor c=0.00457401f \
 //x=2.505 //y=1.655 //x2=2.415 //y2=1.25
cc_2136 ( N_noxref_3_M1_noxref_d N_noxref_5_c_2633_n ) capacitor c=0.00566463f \
 //x=1.96 //y=0.905 //x2=2.415 //y2=1.25
cc_2137 ( N_noxref_3_c_2130_n N_noxref_5_c_2635_n ) capacitor c=0.00877984f \
 //x=2.59 //y=2.59 //x2=1.85 //y2=2.08
cc_2138 ( N_noxref_3_c_2130_n N_noxref_5_c_2636_n ) capacitor c=0.00306024f \
 //x=2.59 //y=2.59 //x2=1.85 //y2=1.915
cc_2139 ( N_noxref_3_M1_noxref_d N_noxref_5_c_2636_n ) capacitor c=0.00660593f \
 //x=1.96 //y=0.905 //x2=1.85 //y2=1.915
cc_2140 ( N_noxref_3_c_2157_n N_noxref_5_c_2638_n ) capacitor c=0.00346627f \
 //x=2.025 //y=5.2 //x2=1.88 //y2=4.7
cc_2141 ( N_noxref_3_c_2130_n N_noxref_5_c_2638_n ) capacitor c=0.00517969f \
 //x=2.59 //y=2.59 //x2=1.88 //y2=4.7
cc_2142 ( N_noxref_3_M57_noxref_g N_noxref_5_M56_noxref_d ) capacitor \
 c=0.0180032f //x=5.08 //y=6.02 //x2=4.715 //y2=5.02
cc_2143 ( N_noxref_3_c_2123_n N_noxref_7_c_3001_n ) capacitor c=0.0105654f \
 //x=9.135 //y=2.59 //x2=11.355 //y2=3.7
cc_2144 ( N_noxref_3_c_2133_n N_noxref_7_c_3001_n ) capacitor c=0.0221017f \
 //x=9.25 //y=2.08 //x2=11.355 //y2=3.7
cc_2145 ( N_noxref_3_c_2123_n N_noxref_7_c_3003_n ) capacitor c=6.33807e-19 \
 //x=9.135 //y=2.59 //x2=6.775 //y2=3.7
cc_2146 ( N_noxref_3_c_2123_n N_noxref_7_c_2955_n ) capacitor c=0.021502f \
 //x=9.135 //y=2.59 //x2=6.66 //y2=2.08
cc_2147 ( N_noxref_3_c_2132_n N_noxref_7_c_2955_n ) capacitor c=0.00140336f \
 //x=4.44 //y=2.08 //x2=6.66 //y2=2.08
cc_2148 ( N_noxref_3_c_2133_n N_noxref_7_c_2955_n ) capacitor c=6.98184e-19 \
 //x=9.25 //y=2.08 //x2=6.66 //y2=2.08
cc_2149 ( N_noxref_3_c_2133_n N_noxref_7_c_2956_n ) capacitor c=0.00118478f \
 //x=9.25 //y=2.08 //x2=11.47 //y2=2.08
cc_2150 ( N_noxref_3_c_2123_n N_noxref_7_c_3008_n ) capacitor c=0.0021022f \
 //x=9.135 //y=2.59 //x2=6.66 //y2=2.08
cc_2151 ( N_noxref_3_c_2117_n N_D_c_4900_n ) capacitor c=0.143317f //x=4.295 \
 //y=2.59 //x2=25.415 //y2=2.96
cc_2152 ( N_noxref_3_c_2121_n N_D_c_4900_n ) capacitor c=0.0293646f //x=2.705 \
 //y=2.59 //x2=25.415 //y2=2.96
cc_2153 ( N_noxref_3_c_2123_n N_D_c_4900_n ) capacitor c=0.0294578f //x=9.135 \
 //y=2.59 //x2=25.415 //y2=2.96
cc_2154 ( N_noxref_3_c_2127_n N_D_c_4900_n ) capacitor c=0.426576f //x=4.705 \
 //y=2.59 //x2=25.415 //y2=2.96
cc_2155 ( N_noxref_3_c_2161_n N_D_c_4900_n ) capacitor c=0.00639146f //x=1.315 \
 //y=5.2 //x2=25.415 //y2=2.96
cc_2156 ( N_noxref_3_c_2259_p N_D_c_4900_n ) capacitor c=0.00647243f //x=2.235 \
 //y=1.655 //x2=25.415 //y2=2.96
cc_2157 ( N_noxref_3_c_2130_n N_D_c_4900_n ) capacitor c=0.0244616f //x=2.59 \
 //y=2.59 //x2=25.415 //y2=2.96
cc_2158 ( N_noxref_3_c_2132_n N_D_c_4900_n ) capacitor c=0.0254538f //x=4.44 \
 //y=2.08 //x2=25.415 //y2=2.96
cc_2159 ( N_noxref_3_c_2133_n N_D_c_4900_n ) capacitor c=0.0239333f //x=9.25 \
 //y=2.08 //x2=25.415 //y2=2.96
cc_2160 ( N_noxref_3_c_2161_n N_D_c_4908_n ) capacitor c=2.77803e-19 //x=1.315 \
 //y=5.2 //x2=1.225 //y2=2.96
cc_2161 ( N_noxref_3_c_2161_n N_D_c_4915_n ) capacitor c=0.00563876f //x=1.315 \
 //y=5.2 //x2=1.11 //y2=2.08
cc_2162 ( N_noxref_3_c_2130_n N_D_c_4915_n ) capacitor c=0.00408104f //x=2.59 \
 //y=2.59 //x2=1.11 //y2=2.08
cc_2163 ( N_noxref_3_c_2161_n N_D_M52_noxref_g ) capacitor c=0.0177326f \
 //x=1.315 //y=5.2 //x2=1.01 //y2=6.02
cc_2164 ( N_noxref_3_c_2157_n N_D_M53_noxref_g ) capacitor c=0.0195934f \
 //x=2.025 //y=5.2 //x2=1.45 //y2=6.02
cc_2165 ( N_noxref_3_M52_noxref_d N_D_M53_noxref_g ) capacitor c=0.0173476f \
 //x=1.085 //y=5.02 //x2=1.45 //y2=6.02
cc_2166 ( N_noxref_3_c_2161_n N_D_c_4971_n ) capacitor c=0.00589848f //x=1.315 \
 //y=5.2 //x2=1.11 //y2=4.7
cc_2167 ( N_noxref_3_c_2133_n N_CLK_c_5631_n ) capacitor c=0.0208709f //x=9.25 \
 //y=2.08 //x2=14.685 //y2=4.44
cc_2168 ( N_noxref_3_c_2184_n N_CLK_c_5631_n ) capacitor c=0.0166984f \
 //x=9.525 //y=4.79 //x2=14.685 //y2=4.44
cc_2169 ( N_noxref_3_c_2132_n N_CLK_c_5642_n ) capacitor c=0.00551083f \
 //x=4.44 //y=2.08 //x2=5.665 //y2=4.44
cc_2170 ( N_noxref_3_c_2123_n N_CLK_c_5622_n ) capacitor c=0.0225267f \
 //x=9.135 //y=2.59 //x2=5.55 //y2=2.08
cc_2171 ( N_noxref_3_c_2127_n N_CLK_c_5622_n ) capacitor c=0.00103784f \
 //x=4.705 //y=2.59 //x2=5.55 //y2=2.08
cc_2172 ( N_noxref_3_c_2130_n N_CLK_c_5622_n ) capacitor c=4.30656e-19 \
 //x=2.59 //y=2.59 //x2=5.55 //y2=2.08
cc_2173 ( N_noxref_3_c_2132_n N_CLK_c_5622_n ) capacitor c=0.0487715f //x=4.44 \
 //y=2.08 //x2=5.55 //y2=2.08
cc_2174 ( N_noxref_3_c_2138_n N_CLK_c_5622_n ) capacitor c=0.00238338f \
 //x=4.14 //y=1.915 //x2=5.55 //y2=2.08
cc_2175 ( N_noxref_3_c_2221_p N_CLK_c_5622_n ) capacitor c=0.00147352f \
 //x=5.005 //y=4.79 //x2=5.55 //y2=2.08
cc_2176 ( N_noxref_3_c_2182_n N_CLK_c_5622_n ) capacitor c=0.00141297f \
 //x=4.715 //y=4.79 //x2=5.55 //y2=2.08
cc_2177 ( N_noxref_3_M56_noxref_g N_CLK_M58_noxref_g ) capacitor c=0.0105869f \
 //x=4.64 //y=6.02 //x2=5.52 //y2=6.02
cc_2178 ( N_noxref_3_M57_noxref_g N_CLK_M58_noxref_g ) capacitor c=0.10632f \
 //x=5.08 //y=6.02 //x2=5.52 //y2=6.02
cc_2179 ( N_noxref_3_M57_noxref_g N_CLK_M59_noxref_g ) capacitor c=0.0101598f \
 //x=5.08 //y=6.02 //x2=5.96 //y2=6.02
cc_2180 ( N_noxref_3_c_2134_n N_CLK_c_5769_n ) capacitor c=5.72482e-19 \
 //x=4.14 //y=0.875 //x2=5.115 //y2=0.91
cc_2181 ( N_noxref_3_c_2136_n N_CLK_c_5769_n ) capacitor c=0.00149976f \
 //x=4.14 //y=1.22 //x2=5.115 //y2=0.91
cc_2182 ( N_noxref_3_c_2141_n N_CLK_c_5769_n ) capacitor c=0.0160123f //x=4.67 \
 //y=0.875 //x2=5.115 //y2=0.91
cc_2183 ( N_noxref_3_c_2137_n N_CLK_c_5772_n ) capacitor c=0.00111227f \
 //x=4.14 //y=1.53 //x2=5.115 //y2=1.22
cc_2184 ( N_noxref_3_c_2143_n N_CLK_c_5772_n ) capacitor c=0.0124075f //x=4.67 \
 //y=1.22 //x2=5.115 //y2=1.22
cc_2185 ( N_noxref_3_c_2141_n N_CLK_c_5774_n ) capacitor c=0.00103227f \
 //x=4.67 //y=0.875 //x2=5.64 //y2=0.91
cc_2186 ( N_noxref_3_c_2143_n N_CLK_c_5775_n ) capacitor c=0.0010154f //x=4.67 \
 //y=1.22 //x2=5.64 //y2=1.22
cc_2187 ( N_noxref_3_c_2143_n N_CLK_c_5776_n ) capacitor c=9.23422e-19 \
 //x=4.67 //y=1.22 //x2=5.64 //y2=1.45
cc_2188 ( N_noxref_3_c_2123_n N_CLK_c_5777_n ) capacitor c=0.0030046f \
 //x=9.135 //y=2.59 //x2=5.64 //y2=1.915
cc_2189 ( N_noxref_3_c_2132_n N_CLK_c_5777_n ) capacitor c=0.00231304f \
 //x=4.44 //y=2.08 //x2=5.64 //y2=1.915
cc_2190 ( N_noxref_3_c_2138_n N_CLK_c_5777_n ) capacitor c=0.00964411f \
 //x=4.14 //y=1.915 //x2=5.64 //y2=1.915
cc_2191 ( N_noxref_3_c_2132_n N_CLK_c_5780_n ) capacitor c=0.00183762f \
 //x=4.44 //y=2.08 //x2=5.55 //y2=4.7
cc_2192 ( N_noxref_3_c_2221_p N_CLK_c_5780_n ) capacitor c=0.0168581f \
 //x=5.005 //y=4.79 //x2=5.55 //y2=4.7
cc_2193 ( N_noxref_3_c_2182_n N_CLK_c_5780_n ) capacitor c=0.00484466f \
 //x=4.715 //y=4.79 //x2=5.55 //y2=4.7
cc_2194 ( N_noxref_3_c_2133_n N_SN_c_6843_n ) capacitor c=0.00558344f //x=9.25 \
 //y=2.08 //x2=10.475 //y2=2.22
cc_2195 ( N_noxref_3_c_2148_n N_SN_c_6843_n ) capacitor c=0.00341397f //x=8.95 \
 //y=1.915 //x2=10.475 //y2=2.22
cc_2196 ( N_noxref_3_c_2123_n N_SN_c_6888_n ) capacitor c=0.00311593f \
 //x=9.135 //y=2.59 //x2=10.36 //y2=2.08
cc_2197 ( N_noxref_3_c_2133_n N_SN_c_6888_n ) capacitor c=0.0458067f //x=9.25 \
 //y=2.08 //x2=10.36 //y2=2.08
cc_2198 ( N_noxref_3_c_2148_n N_SN_c_6888_n ) capacitor c=0.00228225f //x=8.95 \
 //y=1.915 //x2=10.36 //y2=2.08
cc_2199 ( N_noxref_3_c_2200_p N_SN_c_6888_n ) capacitor c=0.00147352f \
 //x=9.815 //y=4.79 //x2=10.36 //y2=2.08
cc_2200 ( N_noxref_3_c_2184_n N_SN_c_6888_n ) capacitor c=0.00142741f \
 //x=9.525 //y=4.79 //x2=10.36 //y2=2.08
cc_2201 ( N_noxref_3_M62_noxref_g N_SN_M64_noxref_g ) capacitor c=0.0105869f \
 //x=9.45 //y=6.02 //x2=10.33 //y2=6.02
cc_2202 ( N_noxref_3_M63_noxref_g N_SN_M64_noxref_g ) capacitor c=0.10632f \
 //x=9.89 //y=6.02 //x2=10.33 //y2=6.02
cc_2203 ( N_noxref_3_M63_noxref_g N_SN_M65_noxref_g ) capacitor c=0.0101598f \
 //x=9.89 //y=6.02 //x2=10.77 //y2=6.02
cc_2204 ( N_noxref_3_c_2144_n N_SN_c_6940_n ) capacitor c=5.72482e-19 //x=8.95 \
 //y=0.875 //x2=9.925 //y2=0.91
cc_2205 ( N_noxref_3_c_2146_n N_SN_c_6940_n ) capacitor c=0.00149976f //x=8.95 \
 //y=1.22 //x2=9.925 //y2=0.91
cc_2206 ( N_noxref_3_c_2151_n N_SN_c_6940_n ) capacitor c=0.0160123f //x=9.48 \
 //y=0.875 //x2=9.925 //y2=0.91
cc_2207 ( N_noxref_3_c_2147_n N_SN_c_6943_n ) capacitor c=0.00111227f //x=8.95 \
 //y=1.53 //x2=9.925 //y2=1.22
cc_2208 ( N_noxref_3_c_2153_n N_SN_c_6943_n ) capacitor c=0.0124075f //x=9.48 \
 //y=1.22 //x2=9.925 //y2=1.22
cc_2209 ( N_noxref_3_c_2151_n N_SN_c_6945_n ) capacitor c=0.00103227f //x=9.48 \
 //y=0.875 //x2=10.45 //y2=0.91
cc_2210 ( N_noxref_3_c_2153_n N_SN_c_6946_n ) capacitor c=0.0010154f //x=9.48 \
 //y=1.22 //x2=10.45 //y2=1.22
cc_2211 ( N_noxref_3_c_2153_n N_SN_c_6947_n ) capacitor c=9.23422e-19 //x=9.48 \
 //y=1.22 //x2=10.45 //y2=1.45
cc_2212 ( N_noxref_3_c_2133_n N_SN_c_6948_n ) capacitor c=0.00211714f //x=9.25 \
 //y=2.08 //x2=10.45 //y2=1.915
cc_2213 ( N_noxref_3_c_2148_n N_SN_c_6948_n ) capacitor c=0.00909574f //x=8.95 \
 //y=1.915 //x2=10.45 //y2=1.915
cc_2214 ( N_noxref_3_c_2133_n N_SN_c_6950_n ) capacitor c=0.00183762f //x=9.25 \
 //y=2.08 //x2=10.36 //y2=4.7
cc_2215 ( N_noxref_3_c_2200_p N_SN_c_6950_n ) capacitor c=0.0168581f //x=9.815 \
 //y=4.79 //x2=10.36 //y2=4.7
cc_2216 ( N_noxref_3_c_2184_n N_SN_c_6950_n ) capacitor c=0.00484466f \
 //x=9.525 //y=4.79 //x2=10.36 //y2=4.7
cc_2217 ( N_noxref_3_c_2259_p N_noxref_27_c_9246_n ) capacitor c=3.15806e-19 \
 //x=2.235 //y=1.655 //x2=0.695 //y2=1.495
cc_2218 ( N_noxref_3_c_2259_p N_noxref_27_c_9235_n ) capacitor c=0.0201674f \
 //x=2.235 //y=1.655 //x2=1.665 //y2=1.495
cc_2219 ( N_noxref_3_c_2129_n N_noxref_27_c_9236_n ) capacitor c=0.00463594f \
 //x=2.505 //y=1.655 //x2=2.55 //y2=0.53
cc_2220 ( N_noxref_3_M1_noxref_d N_noxref_27_c_9236_n ) capacitor c=0.0117318f \
 //x=1.96 //y=0.905 //x2=2.55 //y2=0.53
cc_2221 ( N_noxref_3_c_2117_n N_noxref_27_M0_noxref_s ) capacitor \
 c=2.68031e-19 //x=4.295 //y=2.59 //x2=0.56 //y2=0.365
cc_2222 ( N_noxref_3_c_2121_n N_noxref_27_M0_noxref_s ) capacitor \
 c=5.97427e-19 //x=2.705 //y=2.59 //x2=0.56 //y2=0.365
cc_2223 ( N_noxref_3_c_2129_n N_noxref_27_M0_noxref_s ) capacitor c=0.0129465f \
 //x=2.505 //y=1.655 //x2=0.56 //y2=0.365
cc_2224 ( N_noxref_3_M1_noxref_d N_noxref_27_M0_noxref_s ) capacitor \
 c=0.0437911f //x=1.96 //y=0.905 //x2=0.56 //y2=0.365
cc_2225 ( N_noxref_3_c_2117_n N_noxref_28_c_9293_n ) capacitor c=0.00448771f \
 //x=4.295 //y=2.59 //x2=3.92 //y2=1.505
cc_2226 ( N_noxref_3_c_2129_n N_noxref_28_c_9293_n ) capacitor c=4.08644e-19 \
 //x=2.505 //y=1.655 //x2=3.92 //y2=1.505
cc_2227 ( N_noxref_3_c_2138_n N_noxref_28_c_9293_n ) capacitor c=0.0034165f \
 //x=4.14 //y=1.915 //x2=3.92 //y2=1.505
cc_2228 ( N_noxref_3_c_2117_n N_noxref_28_c_9278_n ) capacitor c=0.00818794f \
 //x=4.295 //y=2.59 //x2=4.805 //y2=1.59
cc_2229 ( N_noxref_3_c_2123_n N_noxref_28_c_9278_n ) capacitor c=0.00225113f \
 //x=9.135 //y=2.59 //x2=4.805 //y2=1.59
cc_2230 ( N_noxref_3_c_2127_n N_noxref_28_c_9278_n ) capacitor c=0.00603529f \
 //x=4.705 //y=2.59 //x2=4.805 //y2=1.59
cc_2231 ( N_noxref_3_c_2132_n N_noxref_28_c_9278_n ) capacitor c=0.0122403f \
 //x=4.44 //y=2.08 //x2=4.805 //y2=1.59
cc_2232 ( N_noxref_3_c_2137_n N_noxref_28_c_9278_n ) capacitor c=0.00703864f \
 //x=4.14 //y=1.53 //x2=4.805 //y2=1.59
cc_2233 ( N_noxref_3_c_2138_n N_noxref_28_c_9278_n ) capacitor c=0.0215834f \
 //x=4.14 //y=1.915 //x2=4.805 //y2=1.59
cc_2234 ( N_noxref_3_c_2140_n N_noxref_28_c_9278_n ) capacitor c=0.00708583f \
 //x=4.515 //y=1.375 //x2=4.805 //y2=1.59
cc_2235 ( N_noxref_3_c_2143_n N_noxref_28_c_9278_n ) capacitor c=0.00698822f \
 //x=4.67 //y=1.22 //x2=4.805 //y2=1.59
cc_2236 ( N_noxref_3_c_2123_n N_noxref_28_c_9304_n ) capacitor c=0.0144126f \
 //x=9.135 //y=2.59 //x2=5.775 //y2=1.59
cc_2237 ( N_noxref_3_c_2123_n N_noxref_28_M2_noxref_s ) capacitor \
 c=0.00867201f //x=9.135 //y=2.59 //x2=3.785 //y2=0.375
cc_2238 ( N_noxref_3_c_2134_n N_noxref_28_M2_noxref_s ) capacitor c=0.0327271f \
 //x=4.14 //y=0.875 //x2=3.785 //y2=0.375
cc_2239 ( N_noxref_3_c_2137_n N_noxref_28_M2_noxref_s ) capacitor \
 c=7.99997e-19 //x=4.14 //y=1.53 //x2=3.785 //y2=0.375
cc_2240 ( N_noxref_3_c_2138_n N_noxref_28_M2_noxref_s ) capacitor \
 c=0.00122123f //x=4.14 //y=1.915 //x2=3.785 //y2=0.375
cc_2241 ( N_noxref_3_c_2141_n N_noxref_28_M2_noxref_s ) capacitor c=0.0121427f \
 //x=4.67 //y=0.875 //x2=3.785 //y2=0.375
cc_2242 ( N_noxref_3_M1_noxref_d N_noxref_28_M2_noxref_s ) capacitor \
 c=2.53688e-19 //x=1.96 //y=0.905 //x2=3.785 //y2=0.375
cc_2243 ( N_noxref_3_c_2123_n N_noxref_29_c_9329_n ) capacitor c=0.00494691f \
 //x=9.135 //y=2.59 //x2=6.345 //y2=0.995
cc_2244 ( N_noxref_3_c_2123_n N_noxref_29_c_9334_n ) capacitor c=8.29806e-19 \
 //x=9.135 //y=2.59 //x2=7.315 //y2=0.54
cc_2245 ( N_noxref_3_c_2123_n N_noxref_29_M4_noxref_s ) capacitor \
 c=0.00448771f //x=9.135 //y=2.59 //x2=6.295 //y2=0.375
cc_2246 ( N_noxref_3_c_2123_n N_noxref_30_c_9396_n ) capacitor c=0.00448771f \
 //x=9.135 //y=2.59 //x2=8.73 //y2=1.505
cc_2247 ( N_noxref_3_c_2148_n N_noxref_30_c_9396_n ) capacitor c=0.0034165f \
 //x=8.95 //y=1.915 //x2=8.73 //y2=1.505
cc_2248 ( N_noxref_3_c_2123_n N_noxref_30_c_9381_n ) capacitor c=0.0116291f \
 //x=9.135 //y=2.59 //x2=9.615 //y2=1.59
cc_2249 ( N_noxref_3_c_2133_n N_noxref_30_c_9381_n ) capacitor c=0.0117813f \
 //x=9.25 //y=2.08 //x2=9.615 //y2=1.59
cc_2250 ( N_noxref_3_c_2147_n N_noxref_30_c_9381_n ) capacitor c=0.00703864f \
 //x=8.95 //y=1.53 //x2=9.615 //y2=1.59
cc_2251 ( N_noxref_3_c_2148_n N_noxref_30_c_9381_n ) capacitor c=0.0215834f \
 //x=8.95 //y=1.915 //x2=9.615 //y2=1.59
cc_2252 ( N_noxref_3_c_2150_n N_noxref_30_c_9381_n ) capacitor c=0.00708583f \
 //x=9.325 //y=1.375 //x2=9.615 //y2=1.59
cc_2253 ( N_noxref_3_c_2153_n N_noxref_30_c_9381_n ) capacitor c=0.00698822f \
 //x=9.48 //y=1.22 //x2=9.615 //y2=1.59
cc_2254 ( N_noxref_3_c_2144_n N_noxref_30_M5_noxref_s ) capacitor c=0.0327271f \
 //x=8.95 //y=0.875 //x2=8.595 //y2=0.375
cc_2255 ( N_noxref_3_c_2147_n N_noxref_30_M5_noxref_s ) capacitor \
 c=7.99997e-19 //x=8.95 //y=1.53 //x2=8.595 //y2=0.375
cc_2256 ( N_noxref_3_c_2148_n N_noxref_30_M5_noxref_s ) capacitor \
 c=0.00122123f //x=8.95 //y=1.915 //x2=8.595 //y2=0.375
cc_2257 ( N_noxref_3_c_2151_n N_noxref_30_M5_noxref_s ) capacitor c=0.0121427f \
 //x=9.48 //y=0.875 //x2=8.595 //y2=0.375
cc_2258 ( N_noxref_4_c_2364_n N_noxref_5_c_2548_n ) capacitor c=0.0181982f \
 //x=12.21 //y=2.59 //x2=17.275 //y2=4.07
cc_2259 ( N_noxref_4_c_2365_n N_noxref_5_c_2548_n ) capacitor c=0.0184765f \
 //x=14.06 //y=2.08 //x2=17.275 //y2=4.07
cc_2260 ( N_noxref_4_c_2381_n N_noxref_5_c_2564_n ) capacitor c=3.10026e-19 \
 //x=9.755 //y=5.155 //x2=7.315 //y2=5.155
cc_2261 ( N_noxref_4_c_2361_n N_noxref_7_c_3009_n ) capacitor c=0.00668132f \
 //x=13.945 //y=2.59 //x2=15.425 //y2=3.7
cc_2262 ( N_noxref_4_c_2362_n N_noxref_7_c_3009_n ) capacitor c=5.89982e-19 \
 //x=12.325 //y=2.59 //x2=15.425 //y2=3.7
cc_2263 ( N_noxref_4_c_2364_n N_noxref_7_c_3009_n ) capacitor c=0.0211098f \
 //x=12.21 //y=2.59 //x2=15.425 //y2=3.7
cc_2264 ( N_noxref_4_c_2365_n N_noxref_7_c_3009_n ) capacitor c=0.0210875f \
 //x=14.06 //y=2.08 //x2=15.425 //y2=3.7
cc_2265 ( N_noxref_4_c_2364_n N_noxref_7_c_3013_n ) capacitor c=0.00117715f \
 //x=12.21 //y=2.59 //x2=11.585 //y2=3.7
cc_2266 ( N_noxref_4_c_2362_n N_noxref_7_c_2956_n ) capacitor c=0.00456439f \
 //x=12.325 //y=2.59 //x2=11.47 //y2=2.08
cc_2267 ( N_noxref_4_c_2364_n N_noxref_7_c_2956_n ) capacitor c=0.079434f \
 //x=12.21 //y=2.59 //x2=11.47 //y2=2.08
cc_2268 ( N_noxref_4_c_2365_n N_noxref_7_c_2956_n ) capacitor c=6.53477e-19 \
 //x=14.06 //y=2.08 //x2=11.47 //y2=2.08
cc_2269 ( N_noxref_4_c_2431_p N_noxref_7_c_2956_n ) capacitor c=0.016476f \
 //x=11.43 //y=5.155 //x2=11.47 //y2=2.08
cc_2270 ( N_noxref_4_M69_noxref_g N_noxref_7_c_2965_n ) capacitor c=0.0169521f \
 //x=14.4 //y=6.02 //x2=14.975 //y2=5.2
cc_2271 ( N_noxref_4_c_2365_n N_noxref_7_c_2969_n ) capacitor c=0.00539951f \
 //x=14.06 //y=2.08 //x2=14.265 //y2=5.2
cc_2272 ( N_noxref_4_M68_noxref_g N_noxref_7_c_2969_n ) capacitor c=0.0177326f \
 //x=13.96 //y=6.02 //x2=14.265 //y2=5.2
cc_2273 ( N_noxref_4_c_2399_n N_noxref_7_c_2969_n ) capacitor c=0.00581252f \
 //x=14.06 //y=4.7 //x2=14.265 //y2=5.2
cc_2274 ( N_noxref_4_c_2364_n N_noxref_7_c_2958_n ) capacitor c=3.52729e-19 \
 //x=12.21 //y=2.59 //x2=15.54 //y2=3.7
cc_2275 ( N_noxref_4_c_2365_n N_noxref_7_c_2958_n ) capacitor c=0.00315608f \
 //x=14.06 //y=2.08 //x2=15.54 //y2=3.7
cc_2276 ( N_noxref_4_c_2383_n N_noxref_7_M66_noxref_g ) capacitor c=0.01736f \
 //x=11.345 //y=5.155 //x2=11.21 //y2=6.02
cc_2277 ( N_noxref_4_M66_noxref_d N_noxref_7_M66_noxref_g ) capacitor \
 c=0.0180032f //x=11.285 //y=5.02 //x2=11.21 //y2=6.02
cc_2278 ( N_noxref_4_c_2387_n N_noxref_7_M67_noxref_g ) capacitor c=0.0194981f \
 //x=12.125 //y=5.155 //x2=11.65 //y2=6.02
cc_2279 ( N_noxref_4_M66_noxref_d N_noxref_7_M67_noxref_g ) capacitor \
 c=0.0194246f //x=11.285 //y=5.02 //x2=11.65 //y2=6.02
cc_2280 ( N_noxref_4_M7_noxref_d N_noxref_7_c_3028_n ) capacitor c=0.00217566f \
 //x=11.535 //y=0.915 //x2=11.46 //y2=0.915
cc_2281 ( N_noxref_4_M7_noxref_d N_noxref_7_c_3029_n ) capacitor c=0.0034598f \
 //x=11.535 //y=0.915 //x2=11.46 //y2=1.26
cc_2282 ( N_noxref_4_M7_noxref_d N_noxref_7_c_3030_n ) capacitor c=0.00546784f \
 //x=11.535 //y=0.915 //x2=11.46 //y2=1.57
cc_2283 ( N_noxref_4_M7_noxref_d N_noxref_7_c_3031_n ) capacitor c=0.00241102f \
 //x=11.535 //y=0.915 //x2=11.835 //y2=0.76
cc_2284 ( N_noxref_4_c_2363_n N_noxref_7_c_3032_n ) capacitor c=0.00371277f \
 //x=12.125 //y=1.665 //x2=11.835 //y2=1.415
cc_2285 ( N_noxref_4_M7_noxref_d N_noxref_7_c_3032_n ) capacitor c=0.0138621f \
 //x=11.535 //y=0.915 //x2=11.835 //y2=1.415
cc_2286 ( N_noxref_4_M7_noxref_d N_noxref_7_c_3034_n ) capacitor c=0.00219619f \
 //x=11.535 //y=0.915 //x2=11.99 //y2=0.915
cc_2287 ( N_noxref_4_c_2363_n N_noxref_7_c_3035_n ) capacitor c=0.00457401f \
 //x=12.125 //y=1.665 //x2=11.99 //y2=1.26
cc_2288 ( N_noxref_4_M7_noxref_d N_noxref_7_c_3035_n ) capacitor c=0.00603828f \
 //x=11.535 //y=0.915 //x2=11.99 //y2=1.26
cc_2289 ( N_noxref_4_c_2364_n N_noxref_7_c_3037_n ) capacitor c=0.00709342f \
 //x=12.21 //y=2.59 //x2=11.47 //y2=2.08
cc_2290 ( N_noxref_4_c_2364_n N_noxref_7_c_3038_n ) capacitor c=0.00283672f \
 //x=12.21 //y=2.59 //x2=11.47 //y2=1.915
cc_2291 ( N_noxref_4_M7_noxref_d N_noxref_7_c_3038_n ) capacitor c=0.00661782f \
 //x=11.535 //y=0.915 //x2=11.47 //y2=1.915
cc_2292 ( N_noxref_4_c_2387_n N_noxref_7_c_3040_n ) capacitor c=0.00201851f \
 //x=12.125 //y=5.155 //x2=11.47 //y2=4.7
cc_2293 ( N_noxref_4_c_2364_n N_noxref_7_c_3040_n ) capacitor c=0.013693f \
 //x=12.21 //y=2.59 //x2=11.47 //y2=4.7
cc_2294 ( N_noxref_4_c_2431_p N_noxref_7_c_3040_n ) capacitor c=0.00475601f \
 //x=11.43 //y=5.155 //x2=11.47 //y2=4.7
cc_2295 ( N_noxref_4_M69_noxref_g N_noxref_7_M68_noxref_d ) capacitor \
 c=0.0173476f //x=14.4 //y=6.02 //x2=14.035 //y2=5.02
cc_2296 ( N_noxref_4_c_2361_n N_D_c_4900_n ) capacitor c=0.172364f //x=13.945 \
 //y=2.59 //x2=25.415 //y2=2.96
cc_2297 ( N_noxref_4_c_2362_n N_D_c_4900_n ) capacitor c=0.0293832f //x=12.325 \
 //y=2.59 //x2=25.415 //y2=2.96
cc_2298 ( N_noxref_4_c_2364_n N_D_c_4900_n ) capacitor c=0.0229414f //x=12.21 \
 //y=2.59 //x2=25.415 //y2=2.96
cc_2299 ( N_noxref_4_c_2365_n N_D_c_4900_n ) capacitor c=0.0229194f //x=14.06 \
 //y=2.08 //x2=25.415 //y2=2.96
cc_2300 ( N_noxref_4_c_2377_n N_CLK_c_5631_n ) capacitor c=0.032141f \
 //x=10.465 //y=5.155 //x2=14.685 //y2=4.44
cc_2301 ( N_noxref_4_c_2381_n N_CLK_c_5631_n ) capacitor c=0.0230136f \
 //x=9.755 //y=5.155 //x2=14.685 //y2=4.44
cc_2302 ( N_noxref_4_c_2387_n N_CLK_c_5631_n ) capacitor c=0.0183122f \
 //x=12.125 //y=5.155 //x2=14.685 //y2=4.44
cc_2303 ( N_noxref_4_c_2364_n N_CLK_c_5631_n ) capacitor c=0.0210274f \
 //x=12.21 //y=2.59 //x2=14.685 //y2=4.44
cc_2304 ( N_noxref_4_c_2365_n N_CLK_c_5631_n ) capacitor c=0.0198304f \
 //x=14.06 //y=2.08 //x2=14.685 //y2=4.44
cc_2305 ( N_noxref_4_c_2399_n N_CLK_c_5631_n ) capacitor c=0.0107057f \
 //x=14.06 //y=4.7 //x2=14.685 //y2=4.44
cc_2306 ( N_noxref_4_c_2365_n N_CLK_c_5667_n ) capacitor c=0.00168329f \
 //x=14.06 //y=2.08 //x2=14.915 //y2=4.44
cc_2307 ( N_noxref_4_c_2399_n N_CLK_c_5667_n ) capacitor c=2.91071e-19 \
 //x=14.06 //y=4.7 //x2=14.915 //y2=4.44
cc_2308 ( N_noxref_4_c_2365_n N_CLK_c_5791_n ) capacitor c=0.00400249f \
 //x=14.06 //y=2.08 //x2=14.8 //y2=4.535
cc_2309 ( N_noxref_4_c_2399_n N_CLK_c_5791_n ) capacitor c=0.00415951f \
 //x=14.06 //y=4.7 //x2=14.8 //y2=4.535
cc_2310 ( N_noxref_4_c_2361_n N_CLK_c_5623_n ) capacitor c=0.00720056f \
 //x=13.945 //y=2.59 //x2=14.8 //y2=2.08
cc_2311 ( N_noxref_4_c_2364_n N_CLK_c_5623_n ) capacitor c=7.62201e-19 \
 //x=12.21 //y=2.59 //x2=14.8 //y2=2.08
cc_2312 ( N_noxref_4_c_2365_n N_CLK_c_5623_n ) capacitor c=0.0737918f \
 //x=14.06 //y=2.08 //x2=14.8 //y2=2.08
cc_2313 ( N_noxref_4_c_2370_n N_CLK_c_5623_n ) capacitor c=0.00284029f \
 //x=13.865 //y=1.915 //x2=14.8 //y2=2.08
cc_2314 ( N_noxref_4_M68_noxref_g N_CLK_M70_noxref_g ) capacitor c=0.0104611f \
 //x=13.96 //y=6.02 //x2=14.84 //y2=6.02
cc_2315 ( N_noxref_4_M69_noxref_g N_CLK_M70_noxref_g ) capacitor c=0.106811f \
 //x=14.4 //y=6.02 //x2=14.84 //y2=6.02
cc_2316 ( N_noxref_4_M69_noxref_g N_CLK_M71_noxref_g ) capacitor c=0.0100341f \
 //x=14.4 //y=6.02 //x2=15.28 //y2=6.02
cc_2317 ( N_noxref_4_c_2366_n N_CLK_c_5800_n ) capacitor c=4.86506e-19 \
 //x=13.865 //y=0.865 //x2=14.835 //y2=0.905
cc_2318 ( N_noxref_4_c_2368_n N_CLK_c_5800_n ) capacitor c=0.00152104f \
 //x=13.865 //y=1.21 //x2=14.835 //y2=0.905
cc_2319 ( N_noxref_4_c_2373_n N_CLK_c_5800_n ) capacitor c=0.0151475f \
 //x=14.395 //y=0.865 //x2=14.835 //y2=0.905
cc_2320 ( N_noxref_4_c_2369_n N_CLK_c_5803_n ) capacitor c=0.00109982f \
 //x=13.865 //y=1.52 //x2=14.835 //y2=1.25
cc_2321 ( N_noxref_4_c_2375_n N_CLK_c_5803_n ) capacitor c=0.0111064f \
 //x=14.395 //y=1.21 //x2=14.835 //y2=1.25
cc_2322 ( N_noxref_4_c_2369_n N_CLK_c_5805_n ) capacitor c=9.57794e-19 \
 //x=13.865 //y=1.52 //x2=14.835 //y2=1.56
cc_2323 ( N_noxref_4_c_2370_n N_CLK_c_5805_n ) capacitor c=0.00662747f \
 //x=13.865 //y=1.915 //x2=14.835 //y2=1.56
cc_2324 ( N_noxref_4_c_2375_n N_CLK_c_5805_n ) capacitor c=0.00862358f \
 //x=14.395 //y=1.21 //x2=14.835 //y2=1.56
cc_2325 ( N_noxref_4_c_2373_n N_CLK_c_5808_n ) capacitor c=0.00124821f \
 //x=14.395 //y=0.865 //x2=15.365 //y2=0.905
cc_2326 ( N_noxref_4_c_2375_n N_CLK_c_5809_n ) capacitor c=0.00200715f \
 //x=14.395 //y=1.21 //x2=15.365 //y2=1.25
cc_2327 ( N_noxref_4_c_2365_n N_CLK_c_5810_n ) capacitor c=0.00282278f \
 //x=14.06 //y=2.08 //x2=14.8 //y2=2.08
cc_2328 ( N_noxref_4_c_2370_n N_CLK_c_5810_n ) capacitor c=0.0172771f \
 //x=13.865 //y=1.915 //x2=14.8 //y2=2.08
cc_2329 ( N_noxref_4_c_2365_n N_CLK_c_5812_n ) capacitor c=0.00342116f \
 //x=14.06 //y=2.08 //x2=14.83 //y2=4.7
cc_2330 ( N_noxref_4_c_2399_n N_CLK_c_5812_n ) capacitor c=0.0292158f \
 //x=14.06 //y=4.7 //x2=14.83 //y2=4.7
cc_2331 ( N_noxref_4_c_2361_n N_SN_c_6833_n ) capacitor c=0.172308f //x=13.945 \
 //y=2.59 //x2=21.715 //y2=2.22
cc_2332 ( N_noxref_4_c_2362_n N_SN_c_6833_n ) capacitor c=0.0291301f \
 //x=12.325 //y=2.59 //x2=21.715 //y2=2.22
cc_2333 ( N_noxref_4_c_2495_p N_SN_c_6833_n ) capacitor c=0.016327f //x=11.81 \
 //y=1.665 //x2=21.715 //y2=2.22
cc_2334 ( N_noxref_4_c_2364_n N_SN_c_6833_n ) capacitor c=0.0215653f //x=12.21 \
 //y=2.59 //x2=21.715 //y2=2.22
cc_2335 ( N_noxref_4_c_2365_n N_SN_c_6833_n ) capacitor c=0.0203358f //x=14.06 \
 //y=2.08 //x2=21.715 //y2=2.22
cc_2336 ( N_noxref_4_c_2370_n N_SN_c_6833_n ) capacitor c=0.00894156f \
 //x=13.865 //y=1.915 //x2=21.715 //y2=2.22
cc_2337 ( N_noxref_4_c_2377_n N_SN_c_6888_n ) capacitor c=0.0144268f \
 //x=10.465 //y=5.155 //x2=10.36 //y2=2.08
cc_2338 ( N_noxref_4_c_2364_n N_SN_c_6888_n ) capacitor c=0.00253274f \
 //x=12.21 //y=2.59 //x2=10.36 //y2=2.08
cc_2339 ( N_noxref_4_c_2377_n N_SN_M64_noxref_g ) capacitor c=0.0165266f \
 //x=10.465 //y=5.155 //x2=10.33 //y2=6.02
cc_2340 ( N_noxref_4_M64_noxref_d N_SN_M64_noxref_g ) capacitor c=0.0180032f \
 //x=10.405 //y=5.02 //x2=10.33 //y2=6.02
cc_2341 ( N_noxref_4_c_2383_n N_SN_M65_noxref_g ) capacitor c=0.01736f \
 //x=11.345 //y=5.155 //x2=10.77 //y2=6.02
cc_2342 ( N_noxref_4_M64_noxref_d N_SN_M65_noxref_g ) capacitor c=0.0180032f \
 //x=10.405 //y=5.02 //x2=10.77 //y2=6.02
cc_2343 ( N_noxref_4_c_2505_p N_SN_c_6965_n ) capacitor c=0.00426767f \
 //x=10.55 //y=5.155 //x2=10.695 //y2=4.79
cc_2344 ( N_noxref_4_c_2377_n N_SN_c_6950_n ) capacitor c=0.00322054f \
 //x=10.465 //y=5.155 //x2=10.36 //y2=4.7
cc_2345 ( N_noxref_4_M7_noxref_d N_noxref_30_M5_noxref_s ) capacitor \
 c=0.00309936f //x=11.535 //y=0.915 //x2=8.595 //y2=0.375
cc_2346 ( N_noxref_4_c_2363_n N_noxref_31_c_9439_n ) capacitor c=0.00457167f \
 //x=12.125 //y=1.665 //x2=12.125 //y2=0.54
cc_2347 ( N_noxref_4_M7_noxref_d N_noxref_31_c_9439_n ) capacitor c=0.0115903f \
 //x=11.535 //y=0.915 //x2=12.125 //y2=0.54
cc_2348 ( N_noxref_4_c_2495_p N_noxref_31_c_9449_n ) capacitor c=0.020048f \
 //x=11.81 //y=1.665 //x2=11.24 //y2=0.995
cc_2349 ( N_noxref_4_M7_noxref_d N_noxref_31_M6_noxref_d ) capacitor \
 c=5.27807e-19 //x=11.535 //y=0.915 //x2=10 //y2=0.91
cc_2350 ( N_noxref_4_c_2363_n N_noxref_31_M7_noxref_s ) capacitor c=0.0184051f \
 //x=12.125 //y=1.665 //x2=11.105 //y2=0.375
cc_2351 ( N_noxref_4_M7_noxref_d N_noxref_31_M7_noxref_s ) capacitor \
 c=0.0426444f //x=11.535 //y=0.915 //x2=11.105 //y2=0.375
cc_2352 ( N_noxref_4_c_2363_n N_noxref_32_c_9504_n ) capacitor c=3.04182e-19 \
 //x=12.125 //y=1.665 //x2=13.645 //y2=1.495
cc_2353 ( N_noxref_4_c_2370_n N_noxref_32_c_9504_n ) capacitor c=0.0034165f \
 //x=13.865 //y=1.915 //x2=13.645 //y2=1.495
cc_2354 ( N_noxref_4_c_2365_n N_noxref_32_c_9486_n ) capacitor c=0.011618f \
 //x=14.06 //y=2.08 //x2=14.53 //y2=1.58
cc_2355 ( N_noxref_4_c_2369_n N_noxref_32_c_9486_n ) capacitor c=0.00696403f \
 //x=13.865 //y=1.52 //x2=14.53 //y2=1.58
cc_2356 ( N_noxref_4_c_2370_n N_noxref_32_c_9486_n ) capacitor c=0.0174694f \
 //x=13.865 //y=1.915 //x2=14.53 //y2=1.58
cc_2357 ( N_noxref_4_c_2372_n N_noxref_32_c_9486_n ) capacitor c=0.00776811f \
 //x=14.24 //y=1.365 //x2=14.53 //y2=1.58
cc_2358 ( N_noxref_4_c_2375_n N_noxref_32_c_9486_n ) capacitor c=0.00339872f \
 //x=14.395 //y=1.21 //x2=14.53 //y2=1.58
cc_2359 ( N_noxref_4_c_2370_n N_noxref_32_c_9493_n ) capacitor c=6.71402e-19 \
 //x=13.865 //y=1.915 //x2=14.615 //y2=1.495
cc_2360 ( N_noxref_4_c_2366_n N_noxref_32_M8_noxref_s ) capacitor c=0.0327502f \
 //x=13.865 //y=0.865 //x2=13.51 //y2=0.365
cc_2361 ( N_noxref_4_c_2369_n N_noxref_32_M8_noxref_s ) capacitor \
 c=3.48408e-19 //x=13.865 //y=1.52 //x2=13.51 //y2=0.365
cc_2362 ( N_noxref_4_c_2373_n N_noxref_32_M8_noxref_s ) capacitor c=0.0120759f \
 //x=14.395 //y=0.865 //x2=13.51 //y2=0.365
cc_2363 ( N_noxref_5_c_2548_n N_noxref_6_c_2820_n ) capacitor c=0.0114735f \
 //x=17.275 //y=4.07 //x2=18.985 //y2=4.07
cc_2364 ( N_noxref_5_M73_noxref_g N_noxref_6_c_2821_n ) capacitor c=0.0169521f \
 //x=17.73 //y=6.02 //x2=18.305 //y2=5.2
cc_2365 ( N_noxref_5_c_2528_n N_noxref_6_c_2825_n ) capacitor c=0.00521572f \
 //x=17.39 //y=2.08 //x2=17.595 //y2=5.2
cc_2366 ( N_noxref_5_M72_noxref_g N_noxref_6_c_2825_n ) capacitor c=0.0177326f \
 //x=17.29 //y=6.02 //x2=17.595 //y2=5.2
cc_2367 ( N_noxref_5_c_2581_n N_noxref_6_c_2825_n ) capacitor c=0.00581252f \
 //x=17.39 //y=4.7 //x2=17.595 //y2=5.2
cc_2368 ( N_noxref_5_c_2528_n N_noxref_6_c_2804_n ) capacitor c=0.00305506f \
 //x=17.39 //y=2.08 //x2=18.87 //y2=4.07
cc_2369 ( N_noxref_5_M73_noxref_g N_noxref_6_M72_noxref_d ) capacitor \
 c=0.0173476f //x=17.73 //y=6.02 //x2=17.365 //y2=5.02
cc_2370 ( N_noxref_5_c_2540_n N_noxref_7_c_3001_n ) capacitor c=0.044143f \
 //x=7.28 //y=4.07 //x2=11.355 //y2=3.7
cc_2371 ( N_noxref_5_c_2548_n N_noxref_7_c_3001_n ) capacitor c=0.340271f \
 //x=17.275 //y=4.07 //x2=11.355 //y2=3.7
cc_2372 ( N_noxref_5_c_2551_n N_noxref_7_c_3001_n ) capacitor c=0.0267581f \
 //x=7.51 //y=4.07 //x2=11.355 //y2=3.7
cc_2373 ( N_noxref_5_c_2571_n N_noxref_7_c_3001_n ) capacitor c=0.00219785f \
 //x=7.395 //y=4.07 //x2=11.355 //y2=3.7
cc_2374 ( N_noxref_5_c_2618_n N_noxref_7_c_3001_n ) capacitor c=0.0208458f \
 //x=7.397 //y=3.905 //x2=11.355 //y2=3.7
cc_2375 ( N_noxref_5_c_2540_n N_noxref_7_c_3003_n ) capacitor c=0.0292842f \
 //x=7.28 //y=4.07 //x2=6.775 //y2=3.7
cc_2376 ( N_noxref_5_c_2618_n N_noxref_7_c_3003_n ) capacitor c=0.00179385f \
 //x=7.397 //y=3.905 //x2=6.775 //y2=3.7
cc_2377 ( N_noxref_5_c_2548_n N_noxref_7_c_3009_n ) capacitor c=0.339174f \
 //x=17.275 //y=4.07 //x2=15.425 //y2=3.7
cc_2378 ( N_noxref_5_c_2548_n N_noxref_7_c_3013_n ) capacitor c=0.026596f \
 //x=17.275 //y=4.07 //x2=11.585 //y2=3.7
cc_2379 ( N_noxref_5_c_2548_n N_noxref_7_c_3053_n ) capacitor c=0.17615f \
 //x=17.275 //y=4.07 //x2=22.825 //y2=3.7
cc_2380 ( N_noxref_5_c_2528_n N_noxref_7_c_3053_n ) capacitor c=0.0228984f \
 //x=17.39 //y=2.08 //x2=22.825 //y2=3.7
cc_2381 ( N_noxref_5_c_2548_n N_noxref_7_c_3055_n ) capacitor c=0.026743f \
 //x=17.275 //y=4.07 //x2=15.655 //y2=3.7
cc_2382 ( N_noxref_5_c_2528_n N_noxref_7_c_3055_n ) capacitor c=7.01366e-19 \
 //x=17.39 //y=2.08 //x2=15.655 //y2=3.7
cc_2383 ( N_noxref_5_c_2540_n N_noxref_7_c_2955_n ) capacitor c=0.0197867f \
 //x=7.28 //y=4.07 //x2=6.66 //y2=2.08
cc_2384 ( N_noxref_5_c_2551_n N_noxref_7_c_2955_n ) capacitor c=0.00180189f \
 //x=7.51 //y=4.07 //x2=6.66 //y2=2.08
cc_2385 ( N_noxref_5_c_2666_p N_noxref_7_c_2955_n ) capacitor c=0.0163236f \
 //x=7.4 //y=5.07 //x2=6.66 //y2=2.08
cc_2386 ( N_noxref_5_c_2667_p N_noxref_7_c_2955_n ) capacitor c=0.016476f \
 //x=6.62 //y=5.155 //x2=6.66 //y2=2.08
cc_2387 ( N_noxref_5_c_2571_n N_noxref_7_c_2955_n ) capacitor c=0.00966503f \
 //x=7.395 //y=4.07 //x2=6.66 //y2=2.08
cc_2388 ( N_noxref_5_c_2618_n N_noxref_7_c_2955_n ) capacitor c=0.0555125f \
 //x=7.397 //y=3.905 //x2=6.66 //y2=2.08
cc_2389 ( N_noxref_5_c_2548_n N_noxref_7_c_2956_n ) capacitor c=0.0198068f \
 //x=17.275 //y=4.07 //x2=11.47 //y2=2.08
cc_2390 ( N_noxref_5_c_2548_n N_noxref_7_c_2958_n ) capacitor c=0.020307f \
 //x=17.275 //y=4.07 //x2=15.54 //y2=3.7
cc_2391 ( N_noxref_5_c_2528_n N_noxref_7_c_2958_n ) capacitor c=0.0125457f \
 //x=17.39 //y=2.08 //x2=15.54 //y2=3.7
cc_2392 ( N_noxref_5_c_2560_n N_noxref_7_M60_noxref_g ) capacitor c=0.01736f \
 //x=6.535 //y=5.155 //x2=6.4 //y2=6.02
cc_2393 ( N_noxref_5_M60_noxref_d N_noxref_7_M60_noxref_g ) capacitor \
 c=0.0180032f //x=6.475 //y=5.02 //x2=6.4 //y2=6.02
cc_2394 ( N_noxref_5_c_2564_n N_noxref_7_M61_noxref_g ) capacitor c=0.0194981f \
 //x=7.315 //y=5.155 //x2=6.84 //y2=6.02
cc_2395 ( N_noxref_5_M60_noxref_d N_noxref_7_M61_noxref_g ) capacitor \
 c=0.0194246f //x=6.475 //y=5.02 //x2=6.84 //y2=6.02
cc_2396 ( N_noxref_5_M4_noxref_d N_noxref_7_c_3070_n ) capacitor c=0.00217566f \
 //x=6.725 //y=0.915 //x2=6.65 //y2=0.915
cc_2397 ( N_noxref_5_M4_noxref_d N_noxref_7_c_3071_n ) capacitor c=0.0034598f \
 //x=6.725 //y=0.915 //x2=6.65 //y2=1.26
cc_2398 ( N_noxref_5_M4_noxref_d N_noxref_7_c_3072_n ) capacitor c=0.00544291f \
 //x=6.725 //y=0.915 //x2=6.65 //y2=1.57
cc_2399 ( N_noxref_5_M4_noxref_d N_noxref_7_c_3073_n ) capacitor c=0.00241102f \
 //x=6.725 //y=0.915 //x2=7.025 //y2=0.76
cc_2400 ( N_noxref_5_c_2527_n N_noxref_7_c_3074_n ) capacitor c=0.00359704f \
 //x=7.315 //y=1.665 //x2=7.025 //y2=1.415
cc_2401 ( N_noxref_5_M4_noxref_d N_noxref_7_c_3074_n ) capacitor c=0.0140297f \
 //x=6.725 //y=0.915 //x2=7.025 //y2=1.415
cc_2402 ( N_noxref_5_M4_noxref_d N_noxref_7_c_3076_n ) capacitor c=0.00219619f \
 //x=6.725 //y=0.915 //x2=7.18 //y2=0.915
cc_2403 ( N_noxref_5_c_2527_n N_noxref_7_c_3077_n ) capacitor c=0.00457401f \
 //x=7.315 //y=1.665 //x2=7.18 //y2=1.26
cc_2404 ( N_noxref_5_M4_noxref_d N_noxref_7_c_3077_n ) capacitor c=0.00603828f \
 //x=6.725 //y=0.915 //x2=7.18 //y2=1.26
cc_2405 ( N_noxref_5_c_2618_n N_noxref_7_c_3008_n ) capacitor c=0.00772308f \
 //x=7.397 //y=3.905 //x2=6.66 //y2=2.08
cc_2406 ( N_noxref_5_c_2618_n N_noxref_7_c_3080_n ) capacitor c=0.00404774f \
 //x=7.397 //y=3.905 //x2=6.66 //y2=1.915
cc_2407 ( N_noxref_5_M4_noxref_d N_noxref_7_c_3080_n ) capacitor c=0.00661782f \
 //x=6.725 //y=0.915 //x2=6.66 //y2=1.915
cc_2408 ( N_noxref_5_c_2564_n N_noxref_7_c_3082_n ) capacitor c=0.00201851f \
 //x=7.315 //y=5.155 //x2=6.66 //y2=4.7
cc_2409 ( N_noxref_5_c_2666_p N_noxref_7_c_3082_n ) capacitor c=0.0151148f \
 //x=7.4 //y=5.07 //x2=6.66 //y2=4.7
cc_2410 ( N_noxref_5_c_2667_p N_noxref_7_c_3082_n ) capacitor c=0.00475601f \
 //x=6.62 //y=5.155 //x2=6.66 //y2=4.7
cc_2411 ( N_noxref_5_c_2540_n N_D_c_4900_n ) capacitor c=0.13371f //x=7.28 \
 //y=4.07 //x2=25.415 //y2=2.96
cc_2412 ( N_noxref_5_c_2547_n N_D_c_4900_n ) capacitor c=0.0078476f //x=1.965 \
 //y=4.07 //x2=25.415 //y2=2.96
cc_2413 ( N_noxref_5_c_2548_n N_D_c_4900_n ) capacitor c=0.0497735f //x=17.275 \
 //y=4.07 //x2=25.415 //y2=2.96
cc_2414 ( N_noxref_5_c_2551_n N_D_c_4900_n ) capacitor c=3.49201e-19 //x=7.51 \
 //y=4.07 //x2=25.415 //y2=2.96
cc_2415 ( N_noxref_5_c_2525_n N_D_c_4900_n ) capacitor c=0.0253568f //x=1.85 \
 //y=2.08 //x2=25.415 //y2=2.96
cc_2416 ( N_noxref_5_c_2528_n N_D_c_4900_n ) capacitor c=0.0233491f //x=17.39 \
 //y=2.08 //x2=25.415 //y2=2.96
cc_2417 ( N_noxref_5_c_2618_n N_D_c_4900_n ) capacitor c=0.0210801f //x=7.397 \
 //y=3.905 //x2=25.415 //y2=2.96
cc_2418 ( N_noxref_5_c_2635_n N_D_c_4900_n ) capacitor c=0.00172252f //x=1.85 \
 //y=2.08 //x2=25.415 //y2=2.96
cc_2419 ( N_noxref_5_c_2525_n N_D_c_4908_n ) capacitor c=0.00179385f //x=1.85 \
 //y=2.08 //x2=1.225 //y2=2.96
cc_2420 ( N_noxref_5_c_2547_n N_D_c_4915_n ) capacitor c=0.00642908f //x=1.965 \
 //y=4.07 //x2=1.11 //y2=2.08
cc_2421 ( N_noxref_5_c_2608_n N_D_c_4915_n ) capacitor c=0.00400249f //x=1.85 \
 //y=4.535 //x2=1.11 //y2=2.08
cc_2422 ( N_noxref_5_c_2525_n N_D_c_4915_n ) capacitor c=0.0838182f //x=1.85 \
 //y=2.08 //x2=1.11 //y2=2.08
cc_2423 ( N_noxref_5_c_2635_n N_D_c_4915_n ) capacitor c=0.00307062f //x=1.85 \
 //y=2.08 //x2=1.11 //y2=2.08
cc_2424 ( N_noxref_5_c_2638_n N_D_c_4915_n ) capacitor c=0.00344981f //x=1.88 \
 //y=4.7 //x2=1.11 //y2=2.08
cc_2425 ( N_noxref_5_M54_noxref_g N_D_M52_noxref_g ) capacitor c=0.0104611f \
 //x=1.89 //y=6.02 //x2=1.01 //y2=6.02
cc_2426 ( N_noxref_5_M54_noxref_g N_D_M53_noxref_g ) capacitor c=0.106811f \
 //x=1.89 //y=6.02 //x2=1.45 //y2=6.02
cc_2427 ( N_noxref_5_M55_noxref_g N_D_M53_noxref_g ) capacitor c=0.0100341f \
 //x=2.33 //y=6.02 //x2=1.45 //y2=6.02
cc_2428 ( N_noxref_5_c_2624_n N_D_c_4918_n ) capacitor c=4.86506e-19 //x=1.885 \
 //y=0.905 //x2=0.915 //y2=0.865
cc_2429 ( N_noxref_5_c_2624_n N_D_c_4920_n ) capacitor c=0.00152104f //x=1.885 \
 //y=0.905 //x2=0.915 //y2=1.21
cc_2430 ( N_noxref_5_c_2625_n N_D_c_4921_n ) capacitor c=0.00109982f //x=1.885 \
 //y=1.25 //x2=0.915 //y2=1.52
cc_2431 ( N_noxref_5_c_2626_n N_D_c_4921_n ) capacitor c=9.57794e-19 //x=1.885 \
 //y=1.56 //x2=0.915 //y2=1.52
cc_2432 ( N_noxref_5_c_2525_n N_D_c_4922_n ) capacitor c=0.00308814f //x=1.85 \
 //y=2.08 //x2=0.915 //y2=1.915
cc_2433 ( N_noxref_5_c_2626_n N_D_c_4922_n ) capacitor c=0.00662747f //x=1.885 \
 //y=1.56 //x2=0.915 //y2=1.915
cc_2434 ( N_noxref_5_c_2635_n N_D_c_4922_n ) capacitor c=0.0179092f //x=1.85 \
 //y=2.08 //x2=0.915 //y2=1.915
cc_2435 ( N_noxref_5_c_2624_n N_D_c_4925_n ) capacitor c=0.0151475f //x=1.885 \
 //y=0.905 //x2=1.445 //y2=0.865
cc_2436 ( N_noxref_5_c_2632_n N_D_c_4925_n ) capacitor c=0.00124821f //x=2.415 \
 //y=0.905 //x2=1.445 //y2=0.865
cc_2437 ( N_noxref_5_c_2625_n N_D_c_4927_n ) capacitor c=0.0111064f //x=1.885 \
 //y=1.25 //x2=1.445 //y2=1.21
cc_2438 ( N_noxref_5_c_2626_n N_D_c_4927_n ) capacitor c=0.00862358f //x=1.885 \
 //y=1.56 //x2=1.445 //y2=1.21
cc_2439 ( N_noxref_5_c_2633_n N_D_c_4927_n ) capacitor c=0.00200715f //x=2.415 \
 //y=1.25 //x2=1.445 //y2=1.21
cc_2440 ( N_noxref_5_c_2608_n N_D_c_4971_n ) capacitor c=0.00417994f //x=1.85 \
 //y=4.535 //x2=1.11 //y2=4.7
cc_2441 ( N_noxref_5_c_2638_n N_D_c_4971_n ) capacitor c=0.0293367f //x=1.88 \
 //y=4.7 //x2=1.11 //y2=4.7
cc_2442 ( N_noxref_5_c_2540_n N_CLK_c_5631_n ) capacitor c=0.139602f //x=7.28 \
 //y=4.07 //x2=14.685 //y2=4.44
cc_2443 ( N_noxref_5_c_2548_n N_CLK_c_5631_n ) capacitor c=0.625476f \
 //x=17.275 //y=4.07 //x2=14.685 //y2=4.44
cc_2444 ( N_noxref_5_c_2551_n N_CLK_c_5631_n ) capacitor c=0.0265302f //x=7.51 \
 //y=4.07 //x2=14.685 //y2=4.44
cc_2445 ( N_noxref_5_c_2564_n N_CLK_c_5631_n ) capacitor c=0.0182691f \
 //x=7.315 //y=5.155 //x2=14.685 //y2=4.44
cc_2446 ( N_noxref_5_c_2666_p N_CLK_c_5631_n ) capacitor c=0.0207896f //x=7.4 \
 //y=5.07 //x2=14.685 //y2=4.44
cc_2447 ( N_noxref_5_c_2728_p N_CLK_c_5631_n ) capacitor c=0.0311227f //x=5.74 \
 //y=5.155 //x2=14.685 //y2=4.44
cc_2448 ( N_noxref_5_c_2571_n N_CLK_c_5631_n ) capacitor c=0.00215288f \
 //x=7.395 //y=4.07 //x2=14.685 //y2=4.44
cc_2449 ( N_noxref_5_c_2540_n N_CLK_c_5642_n ) capacitor c=0.0291328f //x=7.28 \
 //y=4.07 //x2=5.665 //y2=4.44
cc_2450 ( N_noxref_5_c_2554_n N_CLK_c_5642_n ) capacitor c=0.00330099f \
 //x=5.655 //y=5.155 //x2=5.665 //y2=4.44
cc_2451 ( N_noxref_5_c_2548_n N_CLK_c_5643_n ) capacitor c=0.236351f \
 //x=17.275 //y=4.07 //x2=29.855 //y2=4.44
cc_2452 ( N_noxref_5_c_2528_n N_CLK_c_5643_n ) capacitor c=0.021665f //x=17.39 \
 //y=2.08 //x2=29.855 //y2=4.44
cc_2453 ( N_noxref_5_c_2581_n N_CLK_c_5643_n ) capacitor c=0.0107036f \
 //x=17.39 //y=4.7 //x2=29.855 //y2=4.44
cc_2454 ( N_noxref_5_c_2548_n N_CLK_c_5667_n ) capacitor c=0.0267161f \
 //x=17.275 //y=4.07 //x2=14.915 //y2=4.44
cc_2455 ( N_noxref_5_c_2540_n N_CLK_c_5622_n ) capacitor c=0.0247116f //x=7.28 \
 //y=4.07 //x2=5.55 //y2=2.08
cc_2456 ( N_noxref_5_c_2554_n N_CLK_c_5622_n ) capacitor c=0.0143918f \
 //x=5.655 //y=5.155 //x2=5.55 //y2=2.08
cc_2457 ( N_noxref_5_c_2666_p N_CLK_c_5622_n ) capacitor c=7.17254e-19 //x=7.4 \
 //y=5.07 //x2=5.55 //y2=2.08
cc_2458 ( N_noxref_5_c_2618_n N_CLK_c_5622_n ) capacitor c=0.00197044f \
 //x=7.397 //y=3.905 //x2=5.55 //y2=2.08
cc_2459 ( N_noxref_5_c_2548_n N_CLK_c_5623_n ) capacitor c=0.0187718f \
 //x=17.275 //y=4.07 //x2=14.8 //y2=2.08
cc_2460 ( N_noxref_5_c_2528_n N_CLK_c_5623_n ) capacitor c=0.00105438f \
 //x=17.39 //y=2.08 //x2=14.8 //y2=2.08
cc_2461 ( N_noxref_5_c_2554_n N_CLK_M58_noxref_g ) capacitor c=0.016514f \
 //x=5.655 //y=5.155 //x2=5.52 //y2=6.02
cc_2462 ( N_noxref_5_M58_noxref_d N_CLK_M58_noxref_g ) capacitor c=0.0180032f \
 //x=5.595 //y=5.02 //x2=5.52 //y2=6.02
cc_2463 ( N_noxref_5_c_2560_n N_CLK_M59_noxref_g ) capacitor c=0.01736f \
 //x=6.535 //y=5.155 //x2=5.96 //y2=6.02
cc_2464 ( N_noxref_5_M58_noxref_d N_CLK_M59_noxref_g ) capacitor c=0.0180032f \
 //x=5.595 //y=5.02 //x2=5.96 //y2=6.02
cc_2465 ( N_noxref_5_c_2728_p N_CLK_c_5837_n ) capacitor c=0.00426767f \
 //x=5.74 //y=5.155 //x2=5.885 //y2=4.79
cc_2466 ( N_noxref_5_c_2554_n N_CLK_c_5780_n ) capacitor c=0.00322046f \
 //x=5.655 //y=5.155 //x2=5.55 //y2=4.7
cc_2467 ( N_noxref_5_c_2528_n N_SN_c_6833_n ) capacitor c=0.0208418f //x=17.39 \
 //y=2.08 //x2=21.715 //y2=2.22
cc_2468 ( N_noxref_5_c_2533_n N_SN_c_6833_n ) capacitor c=0.00894156f \
 //x=17.195 //y=1.915 //x2=21.715 //y2=2.22
cc_2469 ( N_noxref_5_c_2548_n N_SN_c_6888_n ) capacitor c=0.0190126f \
 //x=17.275 //y=4.07 //x2=10.36 //y2=2.08
cc_2470 ( N_noxref_5_c_2618_n N_SN_c_6888_n ) capacitor c=3.85853e-19 \
 //x=7.397 //y=3.905 //x2=10.36 //y2=2.08
cc_2471 ( N_noxref_5_c_2528_n N_noxref_24_c_8497_n ) capacitor c=0.00735597f \
 //x=17.39 //y=2.08 //x2=18.245 //y2=3.33
cc_2472 ( N_noxref_5_c_2528_n N_noxref_24_c_8498_n ) capacitor c=0.00400249f \
 //x=17.39 //y=2.08 //x2=18.13 //y2=4.535
cc_2473 ( N_noxref_5_c_2581_n N_noxref_24_c_8498_n ) capacitor c=0.00417994f \
 //x=17.39 //y=4.7 //x2=18.13 //y2=4.535
cc_2474 ( N_noxref_5_c_2548_n N_noxref_24_c_8428_n ) capacitor c=0.00318578f \
 //x=17.275 //y=4.07 //x2=18.13 //y2=2.08
cc_2475 ( N_noxref_5_c_2528_n N_noxref_24_c_8428_n ) capacitor c=0.0752164f \
 //x=17.39 //y=2.08 //x2=18.13 //y2=2.08
cc_2476 ( N_noxref_5_c_2533_n N_noxref_24_c_8428_n ) capacitor c=0.00284029f \
 //x=17.195 //y=1.915 //x2=18.13 //y2=2.08
cc_2477 ( N_noxref_5_M72_noxref_g N_noxref_24_M74_noxref_g ) capacitor \
 c=0.0104611f //x=17.29 //y=6.02 //x2=18.17 //y2=6.02
cc_2478 ( N_noxref_5_M73_noxref_g N_noxref_24_M74_noxref_g ) capacitor \
 c=0.106811f //x=17.73 //y=6.02 //x2=18.17 //y2=6.02
cc_2479 ( N_noxref_5_M73_noxref_g N_noxref_24_M75_noxref_g ) capacitor \
 c=0.0100341f //x=17.73 //y=6.02 //x2=18.61 //y2=6.02
cc_2480 ( N_noxref_5_c_2529_n N_noxref_24_c_8506_n ) capacitor c=4.86506e-19 \
 //x=17.195 //y=0.865 //x2=18.165 //y2=0.905
cc_2481 ( N_noxref_5_c_2531_n N_noxref_24_c_8506_n ) capacitor c=0.00152104f \
 //x=17.195 //y=1.21 //x2=18.165 //y2=0.905
cc_2482 ( N_noxref_5_c_2536_n N_noxref_24_c_8506_n ) capacitor c=0.0151475f \
 //x=17.725 //y=0.865 //x2=18.165 //y2=0.905
cc_2483 ( N_noxref_5_c_2532_n N_noxref_24_c_8509_n ) capacitor c=0.00109982f \
 //x=17.195 //y=1.52 //x2=18.165 //y2=1.25
cc_2484 ( N_noxref_5_c_2538_n N_noxref_24_c_8509_n ) capacitor c=0.0111064f \
 //x=17.725 //y=1.21 //x2=18.165 //y2=1.25
cc_2485 ( N_noxref_5_c_2532_n N_noxref_24_c_8511_n ) capacitor c=9.57794e-19 \
 //x=17.195 //y=1.52 //x2=18.165 //y2=1.56
cc_2486 ( N_noxref_5_c_2533_n N_noxref_24_c_8511_n ) capacitor c=0.00662747f \
 //x=17.195 //y=1.915 //x2=18.165 //y2=1.56
cc_2487 ( N_noxref_5_c_2538_n N_noxref_24_c_8511_n ) capacitor c=0.00862358f \
 //x=17.725 //y=1.21 //x2=18.165 //y2=1.56
cc_2488 ( N_noxref_5_c_2536_n N_noxref_24_c_8514_n ) capacitor c=0.00124821f \
 //x=17.725 //y=0.865 //x2=18.695 //y2=0.905
cc_2489 ( N_noxref_5_c_2538_n N_noxref_24_c_8515_n ) capacitor c=0.00200715f \
 //x=17.725 //y=1.21 //x2=18.695 //y2=1.25
cc_2490 ( N_noxref_5_c_2528_n N_noxref_24_c_8516_n ) capacitor c=0.00282278f \
 //x=17.39 //y=2.08 //x2=18.13 //y2=2.08
cc_2491 ( N_noxref_5_c_2533_n N_noxref_24_c_8516_n ) capacitor c=0.0172771f \
 //x=17.195 //y=1.915 //x2=18.13 //y2=2.08
cc_2492 ( N_noxref_5_c_2528_n N_noxref_24_c_8518_n ) capacitor c=0.00344981f \
 //x=17.39 //y=2.08 //x2=18.16 //y2=4.7
cc_2493 ( N_noxref_5_c_2581_n N_noxref_24_c_8518_n ) capacitor c=0.0293367f \
 //x=17.39 //y=4.7 //x2=18.16 //y2=4.7
cc_2494 ( N_noxref_5_c_2626_n N_noxref_27_c_9235_n ) capacitor c=0.00623646f \
 //x=1.885 //y=1.56 //x2=1.665 //y2=1.495
cc_2495 ( N_noxref_5_c_2635_n N_noxref_27_c_9235_n ) capacitor c=0.00174428f \
 //x=1.85 //y=2.08 //x2=1.665 //y2=1.495
cc_2496 ( N_noxref_5_c_2525_n N_noxref_27_c_9236_n ) capacitor c=0.00159235f \
 //x=1.85 //y=2.08 //x2=2.55 //y2=0.53
cc_2497 ( N_noxref_5_c_2624_n N_noxref_27_c_9236_n ) capacitor c=0.0188655f \
 //x=1.885 //y=0.905 //x2=2.55 //y2=0.53
cc_2498 ( N_noxref_5_c_2632_n N_noxref_27_c_9236_n ) capacitor c=0.00656458f \
 //x=2.415 //y=0.905 //x2=2.55 //y2=0.53
cc_2499 ( N_noxref_5_c_2635_n N_noxref_27_c_9236_n ) capacitor c=2.1838e-19 \
 //x=1.85 //y=2.08 //x2=2.55 //y2=0.53
cc_2500 ( N_noxref_5_c_2624_n N_noxref_27_M0_noxref_s ) capacitor \
 c=0.00623646f //x=1.885 //y=0.905 //x2=0.56 //y2=0.365
cc_2501 ( N_noxref_5_c_2632_n N_noxref_27_M0_noxref_s ) capacitor c=0.0143002f \
 //x=2.415 //y=0.905 //x2=0.56 //y2=0.365
cc_2502 ( N_noxref_5_c_2633_n N_noxref_27_M0_noxref_s ) capacitor \
 c=0.00290153f //x=2.415 //y=1.25 //x2=0.56 //y2=0.365
cc_2503 ( N_noxref_5_M4_noxref_d N_noxref_28_M2_noxref_s ) capacitor \
 c=0.00309936f //x=6.725 //y=0.915 //x2=3.785 //y2=0.375
cc_2504 ( N_noxref_5_c_2527_n N_noxref_29_c_9334_n ) capacitor c=0.00461497f \
 //x=7.315 //y=1.665 //x2=7.315 //y2=0.54
cc_2505 ( N_noxref_5_M4_noxref_d N_noxref_29_c_9334_n ) capacitor c=0.0116817f \
 //x=6.725 //y=0.915 //x2=7.315 //y2=0.54
cc_2506 ( N_noxref_5_c_2617_n N_noxref_29_c_9347_n ) capacitor c=0.0200405f \
 //x=7 //y=1.665 //x2=6.43 //y2=0.995
cc_2507 ( N_noxref_5_M4_noxref_d N_noxref_29_M3_noxref_d ) capacitor \
 c=5.27807e-19 //x=6.725 //y=0.915 //x2=5.19 //y2=0.91
cc_2508 ( N_noxref_5_c_2527_n N_noxref_29_M4_noxref_s ) capacitor c=0.0201579f \
 //x=7.315 //y=1.665 //x2=6.295 //y2=0.375
cc_2509 ( N_noxref_5_M4_noxref_d N_noxref_29_M4_noxref_s ) capacitor \
 c=0.0426368f //x=6.725 //y=0.915 //x2=6.295 //y2=0.375
cc_2510 ( N_noxref_5_c_2527_n N_noxref_30_c_9396_n ) capacitor c=3.83325e-19 \
 //x=7.315 //y=1.665 //x2=8.73 //y2=1.505
cc_2511 ( N_noxref_5_M4_noxref_d N_noxref_30_M5_noxref_s ) capacitor \
 c=2.55333e-19 //x=6.725 //y=0.915 //x2=8.595 //y2=0.375
cc_2512 ( N_noxref_5_c_2533_n N_noxref_33_c_9555_n ) capacitor c=0.0034165f \
 //x=17.195 //y=1.915 //x2=16.975 //y2=1.495
cc_2513 ( N_noxref_5_c_2528_n N_noxref_33_c_9537_n ) capacitor c=0.011618f \
 //x=17.39 //y=2.08 //x2=17.86 //y2=1.58
cc_2514 ( N_noxref_5_c_2532_n N_noxref_33_c_9537_n ) capacitor c=0.00696403f \
 //x=17.195 //y=1.52 //x2=17.86 //y2=1.58
cc_2515 ( N_noxref_5_c_2533_n N_noxref_33_c_9537_n ) capacitor c=0.0174694f \
 //x=17.195 //y=1.915 //x2=17.86 //y2=1.58
cc_2516 ( N_noxref_5_c_2535_n N_noxref_33_c_9537_n ) capacitor c=0.00776811f \
 //x=17.57 //y=1.365 //x2=17.86 //y2=1.58
cc_2517 ( N_noxref_5_c_2538_n N_noxref_33_c_9537_n ) capacitor c=0.00339872f \
 //x=17.725 //y=1.21 //x2=17.86 //y2=1.58
cc_2518 ( N_noxref_5_c_2533_n N_noxref_33_c_9544_n ) capacitor c=6.71402e-19 \
 //x=17.195 //y=1.915 //x2=17.945 //y2=1.495
cc_2519 ( N_noxref_5_c_2529_n N_noxref_33_M10_noxref_s ) capacitor \
 c=0.0326577f //x=17.195 //y=0.865 //x2=16.84 //y2=0.365
cc_2520 ( N_noxref_5_c_2532_n N_noxref_33_M10_noxref_s ) capacitor \
 c=3.48408e-19 //x=17.195 //y=1.52 //x2=16.84 //y2=0.365
cc_2521 ( N_noxref_5_c_2536_n N_noxref_33_M10_noxref_s ) capacitor \
 c=0.0120759f //x=17.725 //y=0.865 //x2=16.84 //y2=0.365
cc_2522 ( N_noxref_6_c_2819_n N_noxref_7_c_3053_n ) capacitor c=0.176578f \
 //x=20.605 //y=4.07 //x2=22.825 //y2=3.7
cc_2523 ( N_noxref_6_c_2820_n N_noxref_7_c_3053_n ) capacitor c=0.0293059f \
 //x=18.985 //y=4.07 //x2=22.825 //y2=3.7
cc_2524 ( N_noxref_6_c_2804_n N_noxref_7_c_3053_n ) capacitor c=0.0206035f \
 //x=18.87 //y=4.07 //x2=22.825 //y2=3.7
cc_2525 ( N_noxref_6_c_2805_n N_noxref_7_c_3053_n ) capacitor c=0.021626f \
 //x=20.72 //y=2.08 //x2=22.825 //y2=3.7
cc_2526 ( N_noxref_6_c_2804_n N_noxref_7_c_2958_n ) capacitor c=3.49822e-19 \
 //x=18.87 //y=4.07 //x2=15.54 //y2=3.7
cc_2527 ( N_noxref_6_c_2805_n N_noxref_7_c_2959_n ) capacitor c=0.00117332f \
 //x=20.72 //y=2.08 //x2=22.94 //y2=2.08
cc_2528 ( N_noxref_6_c_2804_n N_D_c_4900_n ) capacitor c=0.0211011f //x=18.87 \
 //y=4.07 //x2=25.415 //y2=2.96
cc_2529 ( N_noxref_6_c_2805_n N_D_c_4900_n ) capacitor c=0.0220754f //x=20.72 \
 //y=2.08 //x2=25.415 //y2=2.96
cc_2530 ( N_noxref_6_c_2819_n N_CLK_c_5643_n ) capacitor c=0.172396f \
 //x=20.605 //y=4.07 //x2=29.855 //y2=4.44
cc_2531 ( N_noxref_6_c_2820_n N_CLK_c_5643_n ) capacitor c=0.029188f \
 //x=18.985 //y=4.07 //x2=29.855 //y2=4.44
cc_2532 ( N_noxref_6_c_2821_n N_CLK_c_5643_n ) capacitor c=0.0185297f \
 //x=18.305 //y=5.2 //x2=29.855 //y2=4.44
cc_2533 ( N_noxref_6_c_2825_n N_CLK_c_5643_n ) capacitor c=0.018142f \
 //x=17.595 //y=5.2 //x2=29.855 //y2=4.44
cc_2534 ( N_noxref_6_c_2804_n N_CLK_c_5643_n ) capacitor c=0.0226667f \
 //x=18.87 //y=4.07 //x2=29.855 //y2=4.44
cc_2535 ( N_noxref_6_c_2805_n N_CLK_c_5643_n ) capacitor c=0.0227055f \
 //x=20.72 //y=2.08 //x2=29.855 //y2=4.44
cc_2536 ( N_noxref_6_c_2839_n N_CLK_c_5643_n ) capacitor c=0.016871f \
 //x=20.995 //y=4.79 //x2=29.855 //y2=4.44
cc_2537 ( N_noxref_6_c_2874_p N_SN_c_6833_n ) capacitor c=0.0146822f \
 //x=18.515 //y=1.655 //x2=21.715 //y2=2.22
cc_2538 ( N_noxref_6_c_2804_n N_SN_c_6833_n ) capacitor c=0.0222456f //x=18.87 \
 //y=4.07 //x2=21.715 //y2=2.22
cc_2539 ( N_noxref_6_c_2805_n N_SN_c_6833_n ) capacitor c=0.0216101f //x=20.72 \
 //y=2.08 //x2=21.715 //y2=2.22
cc_2540 ( N_noxref_6_c_2810_n N_SN_c_6833_n ) capacitor c=0.011987f //x=20.42 \
 //y=1.915 //x2=21.715 //y2=2.22
cc_2541 ( N_noxref_6_c_2805_n N_SN_c_6854_n ) capacitor c=0.00165648f \
 //x=20.72 //y=2.08 //x2=21.945 //y2=2.22
cc_2542 ( N_noxref_6_c_2810_n N_SN_c_6854_n ) capacitor c=2.3323e-19 //x=20.42 \
 //y=1.915 //x2=21.945 //y2=2.22
cc_2543 ( N_noxref_6_c_2819_n N_SN_c_6889_n ) capacitor c=0.00520283f \
 //x=20.605 //y=4.07 //x2=21.83 //y2=2.08
cc_2544 ( N_noxref_6_c_2804_n N_SN_c_6889_n ) capacitor c=4.44801e-19 \
 //x=18.87 //y=4.07 //x2=21.83 //y2=2.08
cc_2545 ( N_noxref_6_c_2805_n N_SN_c_6889_n ) capacitor c=0.0446072f //x=20.72 \
 //y=2.08 //x2=21.83 //y2=2.08
cc_2546 ( N_noxref_6_c_2810_n N_SN_c_6889_n ) capacitor c=0.00208635f \
 //x=20.42 //y=1.915 //x2=21.83 //y2=2.08
cc_2547 ( N_noxref_6_c_2884_p N_SN_c_6889_n ) capacitor c=0.00147352f \
 //x=21.285 //y=4.79 //x2=21.83 //y2=2.08
cc_2548 ( N_noxref_6_c_2839_n N_SN_c_6889_n ) capacitor c=0.00142741f \
 //x=20.995 //y=4.79 //x2=21.83 //y2=2.08
cc_2549 ( N_noxref_6_M76_noxref_g N_SN_M78_noxref_g ) capacitor c=0.0105869f \
 //x=20.92 //y=6.02 //x2=21.8 //y2=6.02
cc_2550 ( N_noxref_6_M77_noxref_g N_SN_M78_noxref_g ) capacitor c=0.10632f \
 //x=21.36 //y=6.02 //x2=21.8 //y2=6.02
cc_2551 ( N_noxref_6_M77_noxref_g N_SN_M79_noxref_g ) capacitor c=0.0101598f \
 //x=21.36 //y=6.02 //x2=22.24 //y2=6.02
cc_2552 ( N_noxref_6_c_2806_n N_SN_c_6986_n ) capacitor c=5.72482e-19 \
 //x=20.42 //y=0.875 //x2=21.395 //y2=0.91
cc_2553 ( N_noxref_6_c_2808_n N_SN_c_6986_n ) capacitor c=0.00149976f \
 //x=20.42 //y=1.22 //x2=21.395 //y2=0.91
cc_2554 ( N_noxref_6_c_2813_n N_SN_c_6986_n ) capacitor c=0.0160123f //x=20.95 \
 //y=0.875 //x2=21.395 //y2=0.91
cc_2555 ( N_noxref_6_c_2809_n N_SN_c_6989_n ) capacitor c=0.00111227f \
 //x=20.42 //y=1.53 //x2=21.395 //y2=1.22
cc_2556 ( N_noxref_6_c_2815_n N_SN_c_6989_n ) capacitor c=0.0124075f //x=20.95 \
 //y=1.22 //x2=21.395 //y2=1.22
cc_2557 ( N_noxref_6_c_2813_n N_SN_c_6991_n ) capacitor c=0.00103227f \
 //x=20.95 //y=0.875 //x2=21.92 //y2=0.91
cc_2558 ( N_noxref_6_c_2815_n N_SN_c_6992_n ) capacitor c=0.0010154f //x=20.95 \
 //y=1.22 //x2=21.92 //y2=1.22
cc_2559 ( N_noxref_6_c_2815_n N_SN_c_6993_n ) capacitor c=9.23422e-19 \
 //x=20.95 //y=1.22 //x2=21.92 //y2=1.45
cc_2560 ( N_noxref_6_c_2805_n N_SN_c_6994_n ) capacitor c=0.00203769f \
 //x=20.72 //y=2.08 //x2=21.92 //y2=1.915
cc_2561 ( N_noxref_6_c_2810_n N_SN_c_6994_n ) capacitor c=0.00834532f \
 //x=20.42 //y=1.915 //x2=21.92 //y2=1.915
cc_2562 ( N_noxref_6_c_2805_n N_SN_c_6996_n ) capacitor c=0.00183762f \
 //x=20.72 //y=2.08 //x2=21.83 //y2=4.7
cc_2563 ( N_noxref_6_c_2884_p N_SN_c_6996_n ) capacitor c=0.0168581f \
 //x=21.285 //y=4.79 //x2=21.83 //y2=4.7
cc_2564 ( N_noxref_6_c_2839_n N_SN_c_6996_n ) capacitor c=0.00484466f \
 //x=20.995 //y=4.79 //x2=21.83 //y2=4.7
cc_2565 ( N_noxref_6_c_2819_n N_noxref_24_c_8520_n ) capacitor c=0.0107182f \
 //x=20.605 //y=4.07 //x2=23.565 //y2=3.33
cc_2566 ( N_noxref_6_c_2820_n N_noxref_24_c_8520_n ) capacitor c=8.94954e-19 \
 //x=18.985 //y=4.07 //x2=23.565 //y2=3.33
cc_2567 ( N_noxref_6_c_2804_n N_noxref_24_c_8520_n ) capacitor c=0.0187691f \
 //x=18.87 //y=4.07 //x2=23.565 //y2=3.33
cc_2568 ( N_noxref_6_c_2805_n N_noxref_24_c_8520_n ) capacitor c=0.0197803f \
 //x=20.72 //y=2.08 //x2=23.565 //y2=3.33
cc_2569 ( N_noxref_6_c_2804_n N_noxref_24_c_8497_n ) capacitor c=0.00179385f \
 //x=18.87 //y=4.07 //x2=18.245 //y2=3.33
cc_2570 ( N_noxref_6_c_2821_n N_noxref_24_c_8498_n ) capacitor c=0.0127164f \
 //x=18.305 //y=5.2 //x2=18.13 //y2=4.535
cc_2571 ( N_noxref_6_c_2804_n N_noxref_24_c_8498_n ) capacitor c=0.0101115f \
 //x=18.87 //y=4.07 //x2=18.13 //y2=4.535
cc_2572 ( N_noxref_6_c_2820_n N_noxref_24_c_8428_n ) capacitor c=0.00329059f \
 //x=18.985 //y=4.07 //x2=18.13 //y2=2.08
cc_2573 ( N_noxref_6_c_2804_n N_noxref_24_c_8428_n ) capacitor c=0.0696067f \
 //x=18.87 //y=4.07 //x2=18.13 //y2=2.08
cc_2574 ( N_noxref_6_c_2805_n N_noxref_24_c_8428_n ) capacitor c=7.5121e-19 \
 //x=20.72 //y=2.08 //x2=18.13 //y2=2.08
cc_2575 ( N_noxref_6_M77_noxref_g N_noxref_24_c_8451_n ) capacitor \
 c=0.0168349f //x=21.36 //y=6.02 //x2=21.935 //y2=5.155
cc_2576 ( N_noxref_6_c_2804_n N_noxref_24_c_8455_n ) capacitor c=2.97874e-19 \
 //x=18.87 //y=4.07 //x2=21.225 //y2=5.155
cc_2577 ( N_noxref_6_M76_noxref_g N_noxref_24_c_8455_n ) capacitor \
 c=0.0213876f //x=20.92 //y=6.02 //x2=21.225 //y2=5.155
cc_2578 ( N_noxref_6_c_2884_p N_noxref_24_c_8455_n ) capacitor c=0.00428486f \
 //x=21.285 //y=4.79 //x2=21.225 //y2=5.155
cc_2579 ( N_noxref_6_c_2821_n N_noxref_24_M74_noxref_g ) capacitor \
 c=0.0166421f //x=18.305 //y=5.2 //x2=18.17 //y2=6.02
cc_2580 ( N_noxref_6_M74_noxref_d N_noxref_24_M74_noxref_g ) capacitor \
 c=0.0173476f //x=18.245 //y=5.02 //x2=18.17 //y2=6.02
cc_2581 ( N_noxref_6_c_2827_n N_noxref_24_M75_noxref_g ) capacitor c=0.018922f \
 //x=18.785 //y=5.2 //x2=18.61 //y2=6.02
cc_2582 ( N_noxref_6_M74_noxref_d N_noxref_24_M75_noxref_g ) capacitor \
 c=0.0179769f //x=18.245 //y=5.02 //x2=18.61 //y2=6.02
cc_2583 ( N_noxref_6_M11_noxref_d N_noxref_24_c_8506_n ) capacitor \
 c=0.00217566f //x=18.24 //y=0.905 //x2=18.165 //y2=0.905
cc_2584 ( N_noxref_6_M11_noxref_d N_noxref_24_c_8509_n ) capacitor \
 c=0.0034598f //x=18.24 //y=0.905 //x2=18.165 //y2=1.25
cc_2585 ( N_noxref_6_M11_noxref_d N_noxref_24_c_8511_n ) capacitor \
 c=0.00669531f //x=18.24 //y=0.905 //x2=18.165 //y2=1.56
cc_2586 ( N_noxref_6_c_2804_n N_noxref_24_c_8541_n ) capacitor c=0.0142673f \
 //x=18.87 //y=4.07 //x2=18.535 //y2=4.79
cc_2587 ( N_noxref_6_c_2924_p N_noxref_24_c_8541_n ) capacitor c=0.00407665f \
 //x=18.39 //y=5.2 //x2=18.535 //y2=4.79
cc_2588 ( N_noxref_6_M11_noxref_d N_noxref_24_c_8543_n ) capacitor \
 c=0.00241102f //x=18.24 //y=0.905 //x2=18.54 //y2=0.75
cc_2589 ( N_noxref_6_c_2803_n N_noxref_24_c_8544_n ) capacitor c=0.00371277f \
 //x=18.785 //y=1.655 //x2=18.54 //y2=1.405
cc_2590 ( N_noxref_6_M11_noxref_d N_noxref_24_c_8544_n ) capacitor \
 c=0.0137169f //x=18.24 //y=0.905 //x2=18.54 //y2=1.405
cc_2591 ( N_noxref_6_M11_noxref_d N_noxref_24_c_8514_n ) capacitor \
 c=0.00132245f //x=18.24 //y=0.905 //x2=18.695 //y2=0.905
cc_2592 ( N_noxref_6_c_2803_n N_noxref_24_c_8515_n ) capacitor c=0.00457401f \
 //x=18.785 //y=1.655 //x2=18.695 //y2=1.25
cc_2593 ( N_noxref_6_M11_noxref_d N_noxref_24_c_8515_n ) capacitor \
 c=0.00566463f //x=18.24 //y=0.905 //x2=18.695 //y2=1.25
cc_2594 ( N_noxref_6_c_2804_n N_noxref_24_c_8516_n ) capacitor c=0.00709342f \
 //x=18.87 //y=4.07 //x2=18.13 //y2=2.08
cc_2595 ( N_noxref_6_c_2804_n N_noxref_24_c_8550_n ) capacitor c=0.00306024f \
 //x=18.87 //y=4.07 //x2=18.13 //y2=1.915
cc_2596 ( N_noxref_6_M11_noxref_d N_noxref_24_c_8550_n ) capacitor \
 c=0.00660593f //x=18.24 //y=0.905 //x2=18.13 //y2=1.915
cc_2597 ( N_noxref_6_c_2821_n N_noxref_24_c_8518_n ) capacitor c=0.00346527f \
 //x=18.305 //y=5.2 //x2=18.16 //y2=4.7
cc_2598 ( N_noxref_6_c_2804_n N_noxref_24_c_8518_n ) capacitor c=0.00533692f \
 //x=18.87 //y=4.07 //x2=18.16 //y2=4.7
cc_2599 ( N_noxref_6_M77_noxref_g N_noxref_24_M76_noxref_d ) capacitor \
 c=0.0180032f //x=21.36 //y=6.02 //x2=20.995 //y2=5.02
cc_2600 ( N_noxref_6_c_2874_p N_noxref_33_c_9555_n ) capacitor c=3.15806e-19 \
 //x=18.515 //y=1.655 //x2=16.975 //y2=1.495
cc_2601 ( N_noxref_6_c_2874_p N_noxref_33_c_9544_n ) capacitor c=0.0203424f \
 //x=18.515 //y=1.655 //x2=17.945 //y2=1.495
cc_2602 ( N_noxref_6_c_2803_n N_noxref_33_c_9545_n ) capacitor c=0.00457164f \
 //x=18.785 //y=1.655 //x2=18.83 //y2=0.53
cc_2603 ( N_noxref_6_M11_noxref_d N_noxref_33_c_9545_n ) capacitor \
 c=0.0115831f //x=18.24 //y=0.905 //x2=18.83 //y2=0.53
cc_2604 ( N_noxref_6_c_2803_n N_noxref_33_M10_noxref_s ) capacitor c=0.013435f \
 //x=18.785 //y=1.655 //x2=16.84 //y2=0.365
cc_2605 ( N_noxref_6_M11_noxref_d N_noxref_33_M10_noxref_s ) capacitor \
 c=0.043966f //x=18.24 //y=0.905 //x2=16.84 //y2=0.365
cc_2606 ( N_noxref_6_c_2803_n N_noxref_34_c_9603_n ) capacitor c=4.08644e-19 \
 //x=18.785 //y=1.655 //x2=20.2 //y2=1.505
cc_2607 ( N_noxref_6_c_2810_n N_noxref_34_c_9603_n ) capacitor c=0.0034165f \
 //x=20.42 //y=1.915 //x2=20.2 //y2=1.505
cc_2608 ( N_noxref_6_c_2805_n N_noxref_34_c_9588_n ) capacitor c=0.0115578f \
 //x=20.72 //y=2.08 //x2=21.085 //y2=1.59
cc_2609 ( N_noxref_6_c_2809_n N_noxref_34_c_9588_n ) capacitor c=0.00697148f \
 //x=20.42 //y=1.53 //x2=21.085 //y2=1.59
cc_2610 ( N_noxref_6_c_2810_n N_noxref_34_c_9588_n ) capacitor c=0.0204849f \
 //x=20.42 //y=1.915 //x2=21.085 //y2=1.59
cc_2611 ( N_noxref_6_c_2812_n N_noxref_34_c_9588_n ) capacitor c=0.00610316f \
 //x=20.795 //y=1.375 //x2=21.085 //y2=1.59
cc_2612 ( N_noxref_6_c_2815_n N_noxref_34_c_9588_n ) capacitor c=0.00698822f \
 //x=20.95 //y=1.22 //x2=21.085 //y2=1.59
cc_2613 ( N_noxref_6_c_2806_n N_noxref_34_M12_noxref_s ) capacitor \
 c=0.0327271f //x=20.42 //y=0.875 //x2=20.065 //y2=0.375
cc_2614 ( N_noxref_6_c_2809_n N_noxref_34_M12_noxref_s ) capacitor \
 c=7.99997e-19 //x=20.42 //y=1.53 //x2=20.065 //y2=0.375
cc_2615 ( N_noxref_6_c_2810_n N_noxref_34_M12_noxref_s ) capacitor \
 c=0.00122123f //x=20.42 //y=1.915 //x2=20.065 //y2=0.375
cc_2616 ( N_noxref_6_c_2813_n N_noxref_34_M12_noxref_s ) capacitor \
 c=0.0121427f //x=20.95 //y=0.875 //x2=20.065 //y2=0.375
cc_2617 ( N_noxref_6_M11_noxref_d N_noxref_34_M12_noxref_s ) capacitor \
 c=2.53688e-19 //x=18.24 //y=0.905 //x2=20.065 //y2=0.375
cc_2618 ( N_noxref_7_c_3001_n N_D_c_4900_n ) capacitor c=0.197056f //x=11.355 \
 //y=3.7 //x2=25.415 //y2=2.96
cc_2619 ( N_noxref_7_c_3003_n N_D_c_4900_n ) capacitor c=0.0135066f //x=6.775 \
 //y=3.7 //x2=25.415 //y2=2.96
cc_2620 ( N_noxref_7_c_3009_n N_D_c_4900_n ) capacitor c=0.164935f //x=15.425 \
 //y=3.7 //x2=25.415 //y2=2.96
cc_2621 ( N_noxref_7_c_3013_n N_D_c_4900_n ) capacitor c=0.0121555f //x=11.585 \
 //y=3.7 //x2=25.415 //y2=2.96
cc_2622 ( N_noxref_7_c_3053_n N_D_c_4900_n ) capacitor c=0.140524f //x=22.825 \
 //y=3.7 //x2=25.415 //y2=2.96
cc_2623 ( N_noxref_7_c_3055_n N_D_c_4900_n ) capacitor c=0.0120929f //x=15.655 \
 //y=3.7 //x2=25.415 //y2=2.96
cc_2624 ( N_noxref_7_c_2955_n N_D_c_4900_n ) capacitor c=0.0206487f //x=6.66 \
 //y=2.08 //x2=25.415 //y2=2.96
cc_2625 ( N_noxref_7_c_2956_n N_D_c_4900_n ) capacitor c=0.0229425f //x=11.47 \
 //y=2.08 //x2=25.415 //y2=2.96
cc_2626 ( N_noxref_7_c_2958_n N_D_c_4900_n ) capacitor c=0.0237328f //x=15.54 \
 //y=3.7 //x2=25.415 //y2=2.96
cc_2627 ( N_noxref_7_c_2959_n N_D_c_4900_n ) capacitor c=0.0202855f //x=22.94 \
 //y=2.08 //x2=25.415 //y2=2.96
cc_2628 ( N_noxref_7_c_2959_n N_D_c_4916_n ) capacitor c=0.00106956f //x=22.94 \
 //y=2.08 //x2=25.53 //y2=2.08
cc_2629 ( N_noxref_7_c_3001_n N_CLK_c_5631_n ) capacitor c=0.0345106f \
 //x=11.355 //y=3.7 //x2=14.685 //y2=4.44
cc_2630 ( N_noxref_7_c_3003_n N_CLK_c_5631_n ) capacitor c=7.0371e-19 \
 //x=6.775 //y=3.7 //x2=14.685 //y2=4.44
cc_2631 ( N_noxref_7_c_3009_n N_CLK_c_5631_n ) capacitor c=0.02107f //x=15.425 \
 //y=3.7 //x2=14.685 //y2=4.44
cc_2632 ( N_noxref_7_c_3013_n N_CLK_c_5631_n ) capacitor c=4.78625e-19 \
 //x=11.585 //y=3.7 //x2=14.685 //y2=4.44
cc_2633 ( N_noxref_7_c_2955_n N_CLK_c_5631_n ) capacitor c=0.0200057f //x=6.66 \
 //y=2.08 //x2=14.685 //y2=4.44
cc_2634 ( N_noxref_7_c_2956_n N_CLK_c_5631_n ) capacitor c=0.0200057f \
 //x=11.47 //y=2.08 //x2=14.685 //y2=4.44
cc_2635 ( N_noxref_7_c_2969_n N_CLK_c_5631_n ) capacitor c=0.0172877f \
 //x=14.265 //y=5.2 //x2=14.685 //y2=4.44
cc_2636 ( N_noxref_7_c_3082_n N_CLK_c_5631_n ) capacitor c=0.0111881f //x=6.66 \
 //y=4.7 //x2=14.685 //y2=4.44
cc_2637 ( N_noxref_7_c_3040_n N_CLK_c_5631_n ) capacitor c=0.0111881f \
 //x=11.47 //y=4.7 //x2=14.685 //y2=4.44
cc_2638 ( N_noxref_7_c_2955_n N_CLK_c_5642_n ) capacitor c=0.00153281f \
 //x=6.66 //y=2.08 //x2=5.665 //y2=4.44
cc_2639 ( N_noxref_7_c_3009_n N_CLK_c_5643_n ) capacitor c=0.0050622f \
 //x=15.425 //y=3.7 //x2=29.855 //y2=4.44
cc_2640 ( N_noxref_7_c_3053_n N_CLK_c_5643_n ) capacitor c=0.166022f \
 //x=22.825 //y=3.7 //x2=29.855 //y2=4.44
cc_2641 ( N_noxref_7_c_3055_n N_CLK_c_5643_n ) capacitor c=5.69483e-19 \
 //x=15.655 //y=3.7 //x2=29.855 //y2=4.44
cc_2642 ( N_noxref_7_c_2965_n N_CLK_c_5643_n ) capacitor c=0.0173598f \
 //x=14.975 //y=5.2 //x2=29.855 //y2=4.44
cc_2643 ( N_noxref_7_c_2958_n N_CLK_c_5643_n ) capacitor c=0.0208321f \
 //x=15.54 //y=3.7 //x2=29.855 //y2=4.44
cc_2644 ( N_noxref_7_c_2959_n N_CLK_c_5643_n ) capacitor c=0.0226638f \
 //x=22.94 //y=2.08 //x2=29.855 //y2=4.44
cc_2645 ( N_noxref_7_c_3118_p N_CLK_c_5643_n ) capacitor c=0.0104371f \
 //x=22.94 //y=4.7 //x2=29.855 //y2=4.44
cc_2646 ( N_noxref_7_c_3009_n N_CLK_c_5667_n ) capacitor c=5.12294e-19 \
 //x=15.425 //y=3.7 //x2=14.915 //y2=4.44
cc_2647 ( N_noxref_7_c_2965_n N_CLK_c_5667_n ) capacitor c=0.0023575f \
 //x=14.975 //y=5.2 //x2=14.915 //y2=4.44
cc_2648 ( N_noxref_7_c_2958_n N_CLK_c_5667_n ) capacitor c=0.00151334f \
 //x=15.54 //y=3.7 //x2=14.915 //y2=4.44
cc_2649 ( N_noxref_7_c_3003_n N_CLK_c_5622_n ) capacitor c=0.00526349f \
 //x=6.775 //y=3.7 //x2=5.55 //y2=2.08
cc_2650 ( N_noxref_7_c_2955_n N_CLK_c_5622_n ) capacitor c=0.0466131f //x=6.66 \
 //y=2.08 //x2=5.55 //y2=2.08
cc_2651 ( N_noxref_7_c_3008_n N_CLK_c_5622_n ) capacitor c=0.00228632f \
 //x=6.66 //y=2.08 //x2=5.55 //y2=2.08
cc_2652 ( N_noxref_7_c_3082_n N_CLK_c_5622_n ) capacitor c=0.00218014f \
 //x=6.66 //y=4.7 //x2=5.55 //y2=2.08
cc_2653 ( N_noxref_7_c_2965_n N_CLK_c_5791_n ) capacitor c=0.0126416f \
 //x=14.975 //y=5.2 //x2=14.8 //y2=4.535
cc_2654 ( N_noxref_7_c_2958_n N_CLK_c_5791_n ) capacitor c=0.00923416f \
 //x=15.54 //y=3.7 //x2=14.8 //y2=4.535
cc_2655 ( N_noxref_7_c_3009_n N_CLK_c_5623_n ) capacitor c=0.0193001f \
 //x=15.425 //y=3.7 //x2=14.8 //y2=2.08
cc_2656 ( N_noxref_7_c_3055_n N_CLK_c_5623_n ) capacitor c=0.00117715f \
 //x=15.655 //y=3.7 //x2=14.8 //y2=2.08
cc_2657 ( N_noxref_7_c_2965_n N_CLK_c_5623_n ) capacitor c=3.74769e-19 \
 //x=14.975 //y=5.2 //x2=14.8 //y2=2.08
cc_2658 ( N_noxref_7_c_2958_n N_CLK_c_5623_n ) capacitor c=0.0701851f \
 //x=15.54 //y=3.7 //x2=14.8 //y2=2.08
cc_2659 ( N_noxref_7_M60_noxref_g N_CLK_M58_noxref_g ) capacitor c=0.0101598f \
 //x=6.4 //y=6.02 //x2=5.52 //y2=6.02
cc_2660 ( N_noxref_7_M60_noxref_g N_CLK_M59_noxref_g ) capacitor c=0.0602553f \
 //x=6.4 //y=6.02 //x2=5.96 //y2=6.02
cc_2661 ( N_noxref_7_M61_noxref_g N_CLK_M59_noxref_g ) capacitor c=0.0101598f \
 //x=6.84 //y=6.02 //x2=5.96 //y2=6.02
cc_2662 ( N_noxref_7_c_2965_n N_CLK_M70_noxref_g ) capacitor c=0.0166421f \
 //x=14.975 //y=5.2 //x2=14.84 //y2=6.02
cc_2663 ( N_noxref_7_M70_noxref_d N_CLK_M70_noxref_g ) capacitor c=0.0173476f \
 //x=14.915 //y=5.02 //x2=14.84 //y2=6.02
cc_2664 ( N_noxref_7_c_2971_n N_CLK_M71_noxref_g ) capacitor c=0.018922f \
 //x=15.455 //y=5.2 //x2=15.28 //y2=6.02
cc_2665 ( N_noxref_7_M70_noxref_d N_CLK_M71_noxref_g ) capacitor c=0.0179769f \
 //x=14.915 //y=5.02 //x2=15.28 //y2=6.02
cc_2666 ( N_noxref_7_c_3070_n N_CLK_c_5774_n ) capacitor c=0.00456962f \
 //x=6.65 //y=0.915 //x2=5.64 //y2=0.91
cc_2667 ( N_noxref_7_c_3071_n N_CLK_c_5775_n ) capacitor c=0.00438372f \
 //x=6.65 //y=1.26 //x2=5.64 //y2=1.22
cc_2668 ( N_noxref_7_c_3072_n N_CLK_c_5776_n ) capacitor c=0.00438372f \
 //x=6.65 //y=1.57 //x2=5.64 //y2=1.45
cc_2669 ( N_noxref_7_c_2955_n N_CLK_c_5777_n ) capacitor c=0.0023343f //x=6.66 \
 //y=2.08 //x2=5.64 //y2=1.915
cc_2670 ( N_noxref_7_c_3008_n N_CLK_c_5777_n ) capacitor c=0.00933826f \
 //x=6.66 //y=2.08 //x2=5.64 //y2=1.915
cc_2671 ( N_noxref_7_c_3080_n N_CLK_c_5777_n ) capacitor c=0.00438372f \
 //x=6.66 //y=1.915 //x2=5.64 //y2=1.915
cc_2672 ( N_noxref_7_c_3082_n N_CLK_c_5837_n ) capacitor c=0.0611812f //x=6.66 \
 //y=4.7 //x2=5.885 //y2=4.79
cc_2673 ( N_noxref_7_M9_noxref_d N_CLK_c_5800_n ) capacitor c=0.00217566f \
 //x=14.91 //y=0.905 //x2=14.835 //y2=0.905
cc_2674 ( N_noxref_7_M9_noxref_d N_CLK_c_5803_n ) capacitor c=0.0034598f \
 //x=14.91 //y=0.905 //x2=14.835 //y2=1.25
cc_2675 ( N_noxref_7_M9_noxref_d N_CLK_c_5805_n ) capacitor c=0.00669531f \
 //x=14.91 //y=0.905 //x2=14.835 //y2=1.56
cc_2676 ( N_noxref_7_c_2958_n N_CLK_c_5893_n ) capacitor c=0.0142673f \
 //x=15.54 //y=3.7 //x2=15.205 //y2=4.79
cc_2677 ( N_noxref_7_c_3150_p N_CLK_c_5893_n ) capacitor c=0.00407665f \
 //x=15.06 //y=5.2 //x2=15.205 //y2=4.79
cc_2678 ( N_noxref_7_M9_noxref_d N_CLK_c_5895_n ) capacitor c=0.00241102f \
 //x=14.91 //y=0.905 //x2=15.21 //y2=0.75
cc_2679 ( N_noxref_7_c_2957_n N_CLK_c_5896_n ) capacitor c=0.00371277f \
 //x=15.455 //y=1.655 //x2=15.21 //y2=1.405
cc_2680 ( N_noxref_7_M9_noxref_d N_CLK_c_5896_n ) capacitor c=0.0137169f \
 //x=14.91 //y=0.905 //x2=15.21 //y2=1.405
cc_2681 ( N_noxref_7_M9_noxref_d N_CLK_c_5808_n ) capacitor c=0.00132245f \
 //x=14.91 //y=0.905 //x2=15.365 //y2=0.905
cc_2682 ( N_noxref_7_c_2957_n N_CLK_c_5809_n ) capacitor c=0.00457401f \
 //x=15.455 //y=1.655 //x2=15.365 //y2=1.25
cc_2683 ( N_noxref_7_M9_noxref_d N_CLK_c_5809_n ) capacitor c=0.00566463f \
 //x=14.91 //y=0.905 //x2=15.365 //y2=1.25
cc_2684 ( N_noxref_7_c_2955_n N_CLK_c_5780_n ) capacitor c=0.00142741f \
 //x=6.66 //y=2.08 //x2=5.55 //y2=4.7
cc_2685 ( N_noxref_7_c_3082_n N_CLK_c_5780_n ) capacitor c=0.00487508f \
 //x=6.66 //y=4.7 //x2=5.55 //y2=4.7
cc_2686 ( N_noxref_7_c_2958_n N_CLK_c_5810_n ) capacitor c=0.00731987f \
 //x=15.54 //y=3.7 //x2=14.8 //y2=2.08
cc_2687 ( N_noxref_7_c_2958_n N_CLK_c_5904_n ) capacitor c=0.00306024f \
 //x=15.54 //y=3.7 //x2=14.8 //y2=1.915
cc_2688 ( N_noxref_7_M9_noxref_d N_CLK_c_5904_n ) capacitor c=0.00660593f \
 //x=14.91 //y=0.905 //x2=14.8 //y2=1.915
cc_2689 ( N_noxref_7_c_2965_n N_CLK_c_5812_n ) capacitor c=0.00346519f \
 //x=14.975 //y=5.2 //x2=14.83 //y2=4.7
cc_2690 ( N_noxref_7_c_2958_n N_CLK_c_5812_n ) capacitor c=0.00518077f \
 //x=15.54 //y=3.7 //x2=14.83 //y2=4.7
cc_2691 ( N_noxref_7_c_3001_n N_SN_c_6833_n ) capacitor c=0.00443649f \
 //x=11.355 //y=3.7 //x2=21.715 //y2=2.22
cc_2692 ( N_noxref_7_c_3009_n N_SN_c_6833_n ) capacitor c=0.00777081f \
 //x=15.425 //y=3.7 //x2=21.715 //y2=2.22
cc_2693 ( N_noxref_7_c_3013_n N_SN_c_6833_n ) capacitor c=2.8328e-19 \
 //x=11.585 //y=3.7 //x2=21.715 //y2=2.22
cc_2694 ( N_noxref_7_c_3053_n N_SN_c_6833_n ) capacitor c=0.00665925f \
 //x=22.825 //y=3.7 //x2=21.715 //y2=2.22
cc_2695 ( N_noxref_7_c_3055_n N_SN_c_6833_n ) capacitor c=2.67441e-19 \
 //x=15.655 //y=3.7 //x2=21.715 //y2=2.22
cc_2696 ( N_noxref_7_c_2956_n N_SN_c_6833_n ) capacitor c=0.0209607f //x=11.47 \
 //y=2.08 //x2=21.715 //y2=2.22
cc_2697 ( N_noxref_7_c_3170_p N_SN_c_6833_n ) capacitor c=0.0146822f \
 //x=15.185 //y=1.655 //x2=21.715 //y2=2.22
cc_2698 ( N_noxref_7_c_2958_n N_SN_c_6833_n ) capacitor c=0.0222456f //x=15.54 \
 //y=3.7 //x2=21.715 //y2=2.22
cc_2699 ( N_noxref_7_c_3032_n N_SN_c_6833_n ) capacitor c=3.13485e-19 \
 //x=11.835 //y=1.415 //x2=21.715 //y2=2.22
cc_2700 ( N_noxref_7_c_3037_n N_SN_c_6833_n ) capacitor c=0.00584491f \
 //x=11.47 //y=2.08 //x2=21.715 //y2=2.22
cc_2701 ( N_noxref_7_c_3001_n N_SN_c_6843_n ) capacitor c=4.71779e-19 \
 //x=11.355 //y=3.7 //x2=10.475 //y2=2.22
cc_2702 ( N_noxref_7_c_2956_n N_SN_c_6843_n ) capacitor c=0.00165648f \
 //x=11.47 //y=2.08 //x2=10.475 //y2=2.22
cc_2703 ( N_noxref_7_c_3037_n N_SN_c_6843_n ) capacitor c=2.3323e-19 //x=11.47 \
 //y=2.08 //x2=10.475 //y2=2.22
cc_2704 ( N_noxref_7_c_2959_n N_SN_c_6844_n ) capacitor c=0.0209607f //x=22.94 \
 //y=2.08 //x2=34.665 //y2=2.22
cc_2705 ( N_noxref_7_c_3178_p N_SN_c_6844_n ) capacitor c=3.13485e-19 \
 //x=23.305 //y=1.415 //x2=34.665 //y2=2.22
cc_2706 ( N_noxref_7_c_3179_p N_SN_c_6844_n ) capacitor c=0.00584491f \
 //x=22.94 //y=2.08 //x2=34.665 //y2=2.22
cc_2707 ( N_noxref_7_c_2959_n N_SN_c_6854_n ) capacitor c=0.00165648f \
 //x=22.94 //y=2.08 //x2=21.945 //y2=2.22
cc_2708 ( N_noxref_7_c_3179_p N_SN_c_6854_n ) capacitor c=2.3323e-19 //x=22.94 \
 //y=2.08 //x2=21.945 //y2=2.22
cc_2709 ( N_noxref_7_c_3001_n N_SN_c_6888_n ) capacitor c=0.0213788f \
 //x=11.355 //y=3.7 //x2=10.36 //y2=2.08
cc_2710 ( N_noxref_7_c_3013_n N_SN_c_6888_n ) capacitor c=0.00128547f \
 //x=11.585 //y=3.7 //x2=10.36 //y2=2.08
cc_2711 ( N_noxref_7_c_2956_n N_SN_c_6888_n ) capacitor c=0.0457045f //x=11.47 \
 //y=2.08 //x2=10.36 //y2=2.08
cc_2712 ( N_noxref_7_c_3037_n N_SN_c_6888_n ) capacitor c=0.0019893f //x=11.47 \
 //y=2.08 //x2=10.36 //y2=2.08
cc_2713 ( N_noxref_7_c_3040_n N_SN_c_6888_n ) capacitor c=0.00219458f \
 //x=11.47 //y=4.7 //x2=10.36 //y2=2.08
cc_2714 ( N_noxref_7_c_3053_n N_SN_c_6889_n ) capacitor c=0.0226304f \
 //x=22.825 //y=3.7 //x2=21.83 //y2=2.08
cc_2715 ( N_noxref_7_c_2959_n N_SN_c_6889_n ) capacitor c=0.0459308f //x=22.94 \
 //y=2.08 //x2=21.83 //y2=2.08
cc_2716 ( N_noxref_7_c_3179_p N_SN_c_6889_n ) capacitor c=0.0019893f //x=22.94 \
 //y=2.08 //x2=21.83 //y2=2.08
cc_2717 ( N_noxref_7_c_3118_p N_SN_c_6889_n ) capacitor c=0.00219458f \
 //x=22.94 //y=4.7 //x2=21.83 //y2=2.08
cc_2718 ( N_noxref_7_M66_noxref_g N_SN_M64_noxref_g ) capacitor c=0.0101598f \
 //x=11.21 //y=6.02 //x2=10.33 //y2=6.02
cc_2719 ( N_noxref_7_M66_noxref_g N_SN_M65_noxref_g ) capacitor c=0.0602553f \
 //x=11.21 //y=6.02 //x2=10.77 //y2=6.02
cc_2720 ( N_noxref_7_M67_noxref_g N_SN_M65_noxref_g ) capacitor c=0.0101598f \
 //x=11.65 //y=6.02 //x2=10.77 //y2=6.02
cc_2721 ( N_noxref_7_M80_noxref_g N_SN_M78_noxref_g ) capacitor c=0.0101598f \
 //x=22.68 //y=6.02 //x2=21.8 //y2=6.02
cc_2722 ( N_noxref_7_M80_noxref_g N_SN_M79_noxref_g ) capacitor c=0.0602553f \
 //x=22.68 //y=6.02 //x2=22.24 //y2=6.02
cc_2723 ( N_noxref_7_M81_noxref_g N_SN_M79_noxref_g ) capacitor c=0.0101598f \
 //x=23.12 //y=6.02 //x2=22.24 //y2=6.02
cc_2724 ( N_noxref_7_c_3028_n N_SN_c_6945_n ) capacitor c=0.00456962f \
 //x=11.46 //y=0.915 //x2=10.45 //y2=0.91
cc_2725 ( N_noxref_7_c_3029_n N_SN_c_6946_n ) capacitor c=0.00438372f \
 //x=11.46 //y=1.26 //x2=10.45 //y2=1.22
cc_2726 ( N_noxref_7_c_3030_n N_SN_c_6947_n ) capacitor c=0.00438372f \
 //x=11.46 //y=1.57 //x2=10.45 //y2=1.45
cc_2727 ( N_noxref_7_c_2956_n N_SN_c_6948_n ) capacitor c=0.00205895f \
 //x=11.47 //y=2.08 //x2=10.45 //y2=1.915
cc_2728 ( N_noxref_7_c_3037_n N_SN_c_6948_n ) capacitor c=0.00828003f \
 //x=11.47 //y=2.08 //x2=10.45 //y2=1.915
cc_2729 ( N_noxref_7_c_3038_n N_SN_c_6948_n ) capacitor c=0.00438372f \
 //x=11.47 //y=1.915 //x2=10.45 //y2=1.915
cc_2730 ( N_noxref_7_c_3040_n N_SN_c_6965_n ) capacitor c=0.0611812f //x=11.47 \
 //y=4.7 //x2=10.695 //y2=4.79
cc_2731 ( N_noxref_7_c_3204_p N_SN_c_6991_n ) capacitor c=0.00456962f \
 //x=22.93 //y=0.915 //x2=21.92 //y2=0.91
cc_2732 ( N_noxref_7_c_3205_p N_SN_c_6992_n ) capacitor c=0.00438372f \
 //x=22.93 //y=1.26 //x2=21.92 //y2=1.22
cc_2733 ( N_noxref_7_c_3206_p N_SN_c_6993_n ) capacitor c=0.00438372f \
 //x=22.93 //y=1.57 //x2=21.92 //y2=1.45
cc_2734 ( N_noxref_7_c_2959_n N_SN_c_6994_n ) capacitor c=0.00205895f \
 //x=22.94 //y=2.08 //x2=21.92 //y2=1.915
cc_2735 ( N_noxref_7_c_3179_p N_SN_c_6994_n ) capacitor c=0.00828003f \
 //x=22.94 //y=2.08 //x2=21.92 //y2=1.915
cc_2736 ( N_noxref_7_c_3209_p N_SN_c_6994_n ) capacitor c=0.00438372f \
 //x=22.94 //y=1.915 //x2=21.92 //y2=1.915
cc_2737 ( N_noxref_7_c_3118_p N_SN_c_7045_n ) capacitor c=0.0611812f //x=22.94 \
 //y=4.7 //x2=22.165 //y2=4.79
cc_2738 ( N_noxref_7_c_2956_n N_SN_c_6950_n ) capacitor c=0.00142741f \
 //x=11.47 //y=2.08 //x2=10.36 //y2=4.7
cc_2739 ( N_noxref_7_c_3040_n N_SN_c_6950_n ) capacitor c=0.00487508f \
 //x=11.47 //y=4.7 //x2=10.36 //y2=4.7
cc_2740 ( N_noxref_7_c_2959_n N_SN_c_6996_n ) capacitor c=0.00142741f \
 //x=22.94 //y=2.08 //x2=21.83 //y2=4.7
cc_2741 ( N_noxref_7_c_3118_p N_SN_c_6996_n ) capacitor c=0.00487508f \
 //x=22.94 //y=4.7 //x2=21.83 //y2=4.7
cc_2742 ( N_noxref_7_c_3053_n N_noxref_24_c_8520_n ) capacitor c=0.433921f \
 //x=22.825 //y=3.7 //x2=23.565 //y2=3.33
cc_2743 ( N_noxref_7_c_2959_n N_noxref_24_c_8520_n ) capacitor c=0.0198536f \
 //x=22.94 //y=2.08 //x2=23.565 //y2=3.33
cc_2744 ( N_noxref_7_c_3053_n N_noxref_24_c_8497_n ) capacitor c=0.0291821f \
 //x=22.825 //y=3.7 //x2=18.245 //y2=3.33
cc_2745 ( N_noxref_7_c_2959_n N_noxref_24_c_8558_n ) capacitor c=0.00179385f \
 //x=22.94 //y=2.08 //x2=23.795 //y2=3.33
cc_2746 ( N_noxref_7_c_3053_n N_noxref_24_c_8428_n ) capacitor c=0.0210992f \
 //x=22.825 //y=3.7 //x2=18.13 //y2=2.08
cc_2747 ( N_noxref_7_c_2958_n N_noxref_24_c_8428_n ) capacitor c=9.43705e-19 \
 //x=15.54 //y=3.7 //x2=18.13 //y2=2.08
cc_2748 ( N_noxref_7_M80_noxref_g N_noxref_24_c_8457_n ) capacitor c=0.01736f \
 //x=22.68 //y=6.02 //x2=22.815 //y2=5.155
cc_2749 ( N_noxref_7_M81_noxref_g N_noxref_24_c_8461_n ) capacitor \
 c=0.0194981f //x=23.12 //y=6.02 //x2=23.595 //y2=5.155
cc_2750 ( N_noxref_7_c_3118_p N_noxref_24_c_8461_n ) capacitor c=0.00201851f \
 //x=22.94 //y=4.7 //x2=23.595 //y2=5.155
cc_2751 ( N_noxref_7_c_3178_p N_noxref_24_c_8430_n ) capacitor c=0.00371277f \
 //x=23.305 //y=1.415 //x2=23.595 //y2=1.665
cc_2752 ( N_noxref_7_c_3225_p N_noxref_24_c_8430_n ) capacitor c=0.00457401f \
 //x=23.46 //y=1.26 //x2=23.595 //y2=1.665
cc_2753 ( N_noxref_7_c_3053_n N_noxref_24_c_8465_n ) capacitor c=0.00735597f \
 //x=22.825 //y=3.7 //x2=23.68 //y2=3.33
cc_2754 ( N_noxref_7_c_2959_n N_noxref_24_c_8465_n ) capacitor c=0.0803969f \
 //x=22.94 //y=2.08 //x2=23.68 //y2=3.33
cc_2755 ( N_noxref_7_c_3179_p N_noxref_24_c_8465_n ) capacitor c=0.00709342f \
 //x=22.94 //y=2.08 //x2=23.68 //y2=3.33
cc_2756 ( N_noxref_7_c_3209_p N_noxref_24_c_8465_n ) capacitor c=0.00283672f \
 //x=22.94 //y=1.915 //x2=23.68 //y2=3.33
cc_2757 ( N_noxref_7_c_3118_p N_noxref_24_c_8465_n ) capacitor c=0.013844f \
 //x=22.94 //y=4.7 //x2=23.68 //y2=3.33
cc_2758 ( N_noxref_7_c_2959_n N_noxref_24_c_8571_n ) capacitor c=0.016476f \
 //x=22.94 //y=2.08 //x2=22.9 //y2=5.155
cc_2759 ( N_noxref_7_c_3118_p N_noxref_24_c_8571_n ) capacitor c=0.00475601f \
 //x=22.94 //y=4.7 //x2=22.9 //y2=5.155
cc_2760 ( N_noxref_7_c_3204_p N_noxref_24_M14_noxref_d ) capacitor \
 c=0.00217566f //x=22.93 //y=0.915 //x2=23.005 //y2=0.915
cc_2761 ( N_noxref_7_c_3205_p N_noxref_24_M14_noxref_d ) capacitor \
 c=0.0034598f //x=22.93 //y=1.26 //x2=23.005 //y2=0.915
cc_2762 ( N_noxref_7_c_3206_p N_noxref_24_M14_noxref_d ) capacitor \
 c=0.00546784f //x=22.93 //y=1.57 //x2=23.005 //y2=0.915
cc_2763 ( N_noxref_7_c_3236_p N_noxref_24_M14_noxref_d ) capacitor \
 c=0.00241102f //x=23.305 //y=0.76 //x2=23.005 //y2=0.915
cc_2764 ( N_noxref_7_c_3178_p N_noxref_24_M14_noxref_d ) capacitor \
 c=0.0138621f //x=23.305 //y=1.415 //x2=23.005 //y2=0.915
cc_2765 ( N_noxref_7_c_3238_p N_noxref_24_M14_noxref_d ) capacitor \
 c=0.00219619f //x=23.46 //y=0.915 //x2=23.005 //y2=0.915
cc_2766 ( N_noxref_7_c_3225_p N_noxref_24_M14_noxref_d ) capacitor \
 c=0.00603828f //x=23.46 //y=1.26 //x2=23.005 //y2=0.915
cc_2767 ( N_noxref_7_c_3209_p N_noxref_24_M14_noxref_d ) capacitor \
 c=0.00661782f //x=22.94 //y=1.915 //x2=23.005 //y2=0.915
cc_2768 ( N_noxref_7_M80_noxref_g N_noxref_24_M80_noxref_d ) capacitor \
 c=0.0180032f //x=22.68 //y=6.02 //x2=22.755 //y2=5.02
cc_2769 ( N_noxref_7_M81_noxref_g N_noxref_24_M80_noxref_d ) capacitor \
 c=0.0194246f //x=23.12 //y=6.02 //x2=22.755 //y2=5.02
cc_2770 ( N_noxref_7_c_2955_n N_noxref_29_c_9334_n ) capacitor c=0.0020642f \
 //x=6.66 //y=2.08 //x2=7.315 //y2=0.54
cc_2771 ( N_noxref_7_c_3070_n N_noxref_29_c_9334_n ) capacitor c=0.0194423f \
 //x=6.65 //y=0.915 //x2=7.315 //y2=0.54
cc_2772 ( N_noxref_7_c_3076_n N_noxref_29_c_9334_n ) capacitor c=0.00656458f \
 //x=7.18 //y=0.915 //x2=7.315 //y2=0.54
cc_2773 ( N_noxref_7_c_3008_n N_noxref_29_c_9334_n ) capacitor c=2.20712e-19 \
 //x=6.66 //y=2.08 //x2=7.315 //y2=0.54
cc_2774 ( N_noxref_7_c_3071_n N_noxref_29_c_9347_n ) capacitor c=0.00538033f \
 //x=6.65 //y=1.26 //x2=6.43 //y2=0.995
cc_2775 ( N_noxref_7_c_3070_n N_noxref_29_M4_noxref_s ) capacitor \
 c=0.00538033f //x=6.65 //y=0.915 //x2=6.295 //y2=0.375
cc_2776 ( N_noxref_7_c_3072_n N_noxref_29_M4_noxref_s ) capacitor \
 c=0.00538033f //x=6.65 //y=1.57 //x2=6.295 //y2=0.375
cc_2777 ( N_noxref_7_c_3076_n N_noxref_29_M4_noxref_s ) capacitor c=0.0143002f \
 //x=7.18 //y=0.915 //x2=6.295 //y2=0.375
cc_2778 ( N_noxref_7_c_3077_n N_noxref_29_M4_noxref_s ) capacitor \
 c=0.00290153f //x=7.18 //y=1.26 //x2=6.295 //y2=0.375
cc_2779 ( N_noxref_7_c_2956_n N_noxref_31_c_9439_n ) capacitor c=0.00204385f \
 //x=11.47 //y=2.08 //x2=12.125 //y2=0.54
cc_2780 ( N_noxref_7_c_3028_n N_noxref_31_c_9439_n ) capacitor c=0.0194423f \
 //x=11.46 //y=0.915 //x2=12.125 //y2=0.54
cc_2781 ( N_noxref_7_c_3034_n N_noxref_31_c_9439_n ) capacitor c=0.00656458f \
 //x=11.99 //y=0.915 //x2=12.125 //y2=0.54
cc_2782 ( N_noxref_7_c_3037_n N_noxref_31_c_9439_n ) capacitor c=2.20712e-19 \
 //x=11.47 //y=2.08 //x2=12.125 //y2=0.54
cc_2783 ( N_noxref_7_c_3029_n N_noxref_31_c_9449_n ) capacitor c=0.00538829f \
 //x=11.46 //y=1.26 //x2=11.24 //y2=0.995
cc_2784 ( N_noxref_7_c_3028_n N_noxref_31_M7_noxref_s ) capacitor \
 c=0.00538829f //x=11.46 //y=0.915 //x2=11.105 //y2=0.375
cc_2785 ( N_noxref_7_c_3030_n N_noxref_31_M7_noxref_s ) capacitor \
 c=0.00538829f //x=11.46 //y=1.57 //x2=11.105 //y2=0.375
cc_2786 ( N_noxref_7_c_3034_n N_noxref_31_M7_noxref_s ) capacitor c=0.0143002f \
 //x=11.99 //y=0.915 //x2=11.105 //y2=0.375
cc_2787 ( N_noxref_7_c_3035_n N_noxref_31_M7_noxref_s ) capacitor \
 c=0.00290153f //x=11.99 //y=1.26 //x2=11.105 //y2=0.375
cc_2788 ( N_noxref_7_c_3170_p N_noxref_32_c_9504_n ) capacitor c=3.15806e-19 \
 //x=15.185 //y=1.655 //x2=13.645 //y2=1.495
cc_2789 ( N_noxref_7_c_3170_p N_noxref_32_c_9493_n ) capacitor c=0.020324f \
 //x=15.185 //y=1.655 //x2=14.615 //y2=1.495
cc_2790 ( N_noxref_7_c_2957_n N_noxref_32_c_9494_n ) capacitor c=0.00457164f \
 //x=15.455 //y=1.655 //x2=15.5 //y2=0.53
cc_2791 ( N_noxref_7_M9_noxref_d N_noxref_32_c_9494_n ) capacitor c=0.0115831f \
 //x=14.91 //y=0.905 //x2=15.5 //y2=0.53
cc_2792 ( N_noxref_7_c_2957_n N_noxref_32_M8_noxref_s ) capacitor c=0.013435f \
 //x=15.455 //y=1.655 //x2=13.51 //y2=0.365
cc_2793 ( N_noxref_7_M9_noxref_d N_noxref_32_M8_noxref_s ) capacitor \
 c=0.0439476f //x=14.91 //y=0.905 //x2=13.51 //y2=0.365
cc_2794 ( N_noxref_7_c_2957_n N_noxref_33_c_9555_n ) capacitor c=3.22188e-19 \
 //x=15.455 //y=1.655 //x2=16.975 //y2=1.495
cc_2795 ( N_noxref_7_c_2959_n N_noxref_35_c_9645_n ) capacitor c=0.00204385f \
 //x=22.94 //y=2.08 //x2=23.595 //y2=0.54
cc_2796 ( N_noxref_7_c_3204_p N_noxref_35_c_9645_n ) capacitor c=0.0194423f \
 //x=22.93 //y=0.915 //x2=23.595 //y2=0.54
cc_2797 ( N_noxref_7_c_3238_p N_noxref_35_c_9645_n ) capacitor c=0.00656458f \
 //x=23.46 //y=0.915 //x2=23.595 //y2=0.54
cc_2798 ( N_noxref_7_c_3179_p N_noxref_35_c_9645_n ) capacitor c=2.20712e-19 \
 //x=22.94 //y=2.08 //x2=23.595 //y2=0.54
cc_2799 ( N_noxref_7_c_3205_p N_noxref_35_c_9657_n ) capacitor c=0.00538829f \
 //x=22.93 //y=1.26 //x2=22.71 //y2=0.995
cc_2800 ( N_noxref_7_c_3204_p N_noxref_35_M14_noxref_s ) capacitor \
 c=0.00538829f //x=22.93 //y=0.915 //x2=22.575 //y2=0.375
cc_2801 ( N_noxref_7_c_3206_p N_noxref_35_M14_noxref_s ) capacitor \
 c=0.00538829f //x=22.93 //y=1.57 //x2=22.575 //y2=0.375
cc_2802 ( N_noxref_7_c_3238_p N_noxref_35_M14_noxref_s ) capacitor \
 c=0.0143002f //x=23.46 //y=0.915 //x2=22.575 //y2=0.375
cc_2803 ( N_noxref_7_c_3225_p N_noxref_35_M14_noxref_s ) capacitor \
 c=0.00290153f //x=23.46 //y=1.26 //x2=22.575 //y2=0.375
cc_2804 ( N_noxref_8_c_3279_n N_noxref_9_c_3510_n ) capacitor c=0.00564994f \
 //x=33.555 //y=2.59 //x2=36.745 //y2=2.59
cc_2805 ( N_noxref_8_M93_noxref_g N_noxref_9_c_3525_n ) capacitor c=0.0168349f \
 //x=34.31 //y=6.02 //x2=34.885 //y2=5.155
cc_2806 ( N_noxref_8_M92_noxref_g N_noxref_9_c_3529_n ) capacitor c=0.0213876f \
 //x=33.87 //y=6.02 //x2=34.175 //y2=5.155
cc_2807 ( N_noxref_8_c_3352_p N_noxref_9_c_3529_n ) capacitor c=0.00428486f \
 //x=34.235 //y=4.79 //x2=34.175 //y2=5.155
cc_2808 ( N_noxref_8_M93_noxref_g N_noxref_9_M92_noxref_d ) capacitor \
 c=0.0180032f //x=34.31 //y=6.02 //x2=33.945 //y2=5.02
cc_2809 ( N_noxref_8_c_3282_n N_noxref_10_c_3690_n ) capacitor c=0.0205341f \
 //x=27.01 //y=2.59 //x2=31.7 //y2=4.07
cc_2810 ( N_noxref_8_c_3284_n N_noxref_10_c_3690_n ) capacitor c=0.021838f \
 //x=28.86 //y=2.08 //x2=31.7 //y2=4.07
cc_2811 ( N_noxref_8_c_3282_n N_noxref_10_c_3742_n ) capacitor c=0.00179385f \
 //x=27.01 //y=2.59 //x2=26.385 //y2=4.07
cc_2812 ( N_noxref_8_c_3285_n N_noxref_10_c_3691_n ) capacitor c=0.0194977f \
 //x=33.67 //y=2.08 //x2=41.695 //y2=4.07
cc_2813 ( N_noxref_8_c_3285_n N_noxref_10_c_3694_n ) capacitor c=3.49381e-19 \
 //x=33.67 //y=2.08 //x2=31.93 //y2=4.07
cc_2814 ( N_noxref_8_c_3309_n N_noxref_10_c_3745_n ) capacitor c=0.0126603f \
 //x=26.445 //y=5.2 //x2=26.27 //y2=4.535
cc_2815 ( N_noxref_8_c_3282_n N_noxref_10_c_3745_n ) capacitor c=0.0101115f \
 //x=27.01 //y=2.59 //x2=26.27 //y2=4.535
cc_2816 ( N_noxref_8_c_3278_n N_noxref_10_c_3675_n ) capacitor c=0.00691549f \
 //x=27.125 //y=2.59 //x2=26.27 //y2=2.08
cc_2817 ( N_noxref_8_c_3282_n N_noxref_10_c_3675_n ) capacitor c=0.0688093f \
 //x=27.01 //y=2.59 //x2=26.27 //y2=2.08
cc_2818 ( N_noxref_8_c_3284_n N_noxref_10_c_3675_n ) capacitor c=6.88047e-19 \
 //x=28.86 //y=2.08 //x2=26.27 //y2=2.08
cc_2819 ( N_noxref_8_M87_noxref_g N_noxref_10_c_3697_n ) capacitor \
 c=0.0168349f //x=29.5 //y=6.02 //x2=30.075 //y2=5.155
cc_2820 ( N_noxref_8_c_3282_n N_noxref_10_c_3701_n ) capacitor c=2.97874e-19 \
 //x=27.01 //y=2.59 //x2=29.365 //y2=5.155
cc_2821 ( N_noxref_8_M86_noxref_g N_noxref_10_c_3701_n ) capacitor \
 c=0.0213876f //x=29.06 //y=6.02 //x2=29.365 //y2=5.155
cc_2822 ( N_noxref_8_c_3367_p N_noxref_10_c_3701_n ) capacitor c=0.00428486f \
 //x=29.425 //y=4.79 //x2=29.365 //y2=5.155
cc_2823 ( N_noxref_8_c_3279_n N_noxref_10_c_3754_n ) capacitor c=0.0165903f \
 //x=33.555 //y=2.59 //x2=31.817 //y2=3.905
cc_2824 ( N_noxref_8_c_3285_n N_noxref_10_c_3754_n ) capacitor c=0.0109272f \
 //x=33.67 //y=2.08 //x2=31.817 //y2=3.905
cc_2825 ( N_noxref_8_c_3309_n N_noxref_10_M84_noxref_g ) capacitor \
 c=0.0166421f //x=26.445 //y=5.2 //x2=26.31 //y2=6.02
cc_2826 ( N_noxref_8_M84_noxref_d N_noxref_10_M84_noxref_g ) capacitor \
 c=0.0173476f //x=26.385 //y=5.02 //x2=26.31 //y2=6.02
cc_2827 ( N_noxref_8_c_3315_n N_noxref_10_M85_noxref_g ) capacitor c=0.018922f \
 //x=26.925 //y=5.2 //x2=26.75 //y2=6.02
cc_2828 ( N_noxref_8_M84_noxref_d N_noxref_10_M85_noxref_g ) capacitor \
 c=0.0179769f //x=26.385 //y=5.02 //x2=26.75 //y2=6.02
cc_2829 ( N_noxref_8_M16_noxref_d N_noxref_10_c_3760_n ) capacitor \
 c=0.00217566f //x=26.38 //y=0.905 //x2=26.305 //y2=0.905
cc_2830 ( N_noxref_8_M16_noxref_d N_noxref_10_c_3761_n ) capacitor \
 c=0.0034598f //x=26.38 //y=0.905 //x2=26.305 //y2=1.25
cc_2831 ( N_noxref_8_M16_noxref_d N_noxref_10_c_3762_n ) capacitor \
 c=0.00669531f //x=26.38 //y=0.905 //x2=26.305 //y2=1.56
cc_2832 ( N_noxref_8_c_3282_n N_noxref_10_c_3763_n ) capacitor c=0.0142673f \
 //x=27.01 //y=2.59 //x2=26.675 //y2=4.79
cc_2833 ( N_noxref_8_c_3378_p N_noxref_10_c_3763_n ) capacitor c=0.00407665f \
 //x=26.53 //y=5.2 //x2=26.675 //y2=4.79
cc_2834 ( N_noxref_8_M16_noxref_d N_noxref_10_c_3765_n ) capacitor \
 c=0.00241102f //x=26.38 //y=0.905 //x2=26.68 //y2=0.75
cc_2835 ( N_noxref_8_c_3281_n N_noxref_10_c_3766_n ) capacitor c=0.00371277f \
 //x=26.925 //y=1.655 //x2=26.68 //y2=1.405
cc_2836 ( N_noxref_8_M16_noxref_d N_noxref_10_c_3766_n ) capacitor \
 c=0.0137169f //x=26.38 //y=0.905 //x2=26.68 //y2=1.405
cc_2837 ( N_noxref_8_M16_noxref_d N_noxref_10_c_3768_n ) capacitor \
 c=0.00132245f //x=26.38 //y=0.905 //x2=26.835 //y2=0.905
cc_2838 ( N_noxref_8_c_3281_n N_noxref_10_c_3769_n ) capacitor c=0.00457401f \
 //x=26.925 //y=1.655 //x2=26.835 //y2=1.25
cc_2839 ( N_noxref_8_M16_noxref_d N_noxref_10_c_3769_n ) capacitor \
 c=0.00566463f //x=26.38 //y=0.905 //x2=26.835 //y2=1.25
cc_2840 ( N_noxref_8_c_3282_n N_noxref_10_c_3771_n ) capacitor c=0.00731987f \
 //x=27.01 //y=2.59 //x2=26.27 //y2=2.08
cc_2841 ( N_noxref_8_c_3282_n N_noxref_10_c_3772_n ) capacitor c=0.00306024f \
 //x=27.01 //y=2.59 //x2=26.27 //y2=1.915
cc_2842 ( N_noxref_8_M16_noxref_d N_noxref_10_c_3772_n ) capacitor \
 c=0.00660593f //x=26.38 //y=0.905 //x2=26.27 //y2=1.915
cc_2843 ( N_noxref_8_c_3309_n N_noxref_10_c_3774_n ) capacitor c=0.00346527f \
 //x=26.445 //y=5.2 //x2=26.3 //y2=4.7
cc_2844 ( N_noxref_8_c_3282_n N_noxref_10_c_3774_n ) capacitor c=0.00517969f \
 //x=27.01 //y=2.59 //x2=26.3 //y2=4.7
cc_2845 ( N_noxref_8_M87_noxref_g N_noxref_10_M86_noxref_d ) capacitor \
 c=0.0180032f //x=29.5 //y=6.02 //x2=29.135 //y2=5.02
cc_2846 ( N_noxref_8_c_3285_n N_noxref_12_c_4157_n ) capacitor c=0.0197627f \
 //x=33.67 //y=2.08 //x2=35.775 //y2=3.7
cc_2847 ( N_noxref_8_c_3279_n N_noxref_12_c_4111_n ) capacitor c=0.0179628f \
 //x=33.555 //y=2.59 //x2=31.08 //y2=2.08
cc_2848 ( N_noxref_8_c_3284_n N_noxref_12_c_4111_n ) capacitor c=0.00108806f \
 //x=28.86 //y=2.08 //x2=31.08 //y2=2.08
cc_2849 ( N_noxref_8_c_3285_n N_noxref_12_c_4111_n ) capacitor c=5.77326e-19 \
 //x=33.67 //y=2.08 //x2=31.08 //y2=2.08
cc_2850 ( N_noxref_8_c_3285_n N_noxref_12_c_4112_n ) capacitor c=0.00102099f \
 //x=33.67 //y=2.08 //x2=35.89 //y2=2.08
cc_2851 ( N_noxref_8_c_3277_n N_D_c_4909_n ) capacitor c=0.143317f //x=28.715 \
 //y=2.59 //x2=49.835 //y2=2.96
cc_2852 ( N_noxref_8_c_3278_n N_D_c_4909_n ) capacitor c=0.0293646f //x=27.125 \
 //y=2.59 //x2=49.835 //y2=2.96
cc_2853 ( N_noxref_8_c_3279_n N_D_c_4909_n ) capacitor c=0.0294578f //x=33.555 \
 //y=2.59 //x2=49.835 //y2=2.96
cc_2854 ( N_noxref_8_c_3280_n N_D_c_4909_n ) capacitor c=0.426576f //x=29.125 \
 //y=2.59 //x2=49.835 //y2=2.96
cc_2855 ( N_noxref_8_c_3282_n N_D_c_4909_n ) capacitor c=0.0206018f //x=27.01 \
 //y=2.59 //x2=49.835 //y2=2.96
cc_2856 ( N_noxref_8_c_3284_n N_D_c_4909_n ) capacitor c=0.0215953f //x=28.86 \
 //y=2.08 //x2=49.835 //y2=2.96
cc_2857 ( N_noxref_8_c_3285_n N_D_c_4909_n ) capacitor c=0.0215933f //x=33.67 \
 //y=2.08 //x2=49.835 //y2=2.96
cc_2858 ( N_noxref_8_c_3313_n N_D_c_4916_n ) capacitor c=0.00539951f \
 //x=25.735 //y=5.2 //x2=25.53 //y2=2.08
cc_2859 ( N_noxref_8_c_3282_n N_D_c_4916_n ) capacitor c=0.00347311f //x=27.01 \
 //y=2.59 //x2=25.53 //y2=2.08
cc_2860 ( N_noxref_8_c_3313_n N_D_M82_noxref_g ) capacitor c=0.0177326f \
 //x=25.735 //y=5.2 //x2=25.43 //y2=6.02
cc_2861 ( N_noxref_8_c_3309_n N_D_M83_noxref_g ) capacitor c=0.0169521f \
 //x=26.445 //y=5.2 //x2=25.87 //y2=6.02
cc_2862 ( N_noxref_8_M82_noxref_d N_D_M83_noxref_g ) capacitor c=0.0173476f \
 //x=25.505 //y=5.02 //x2=25.87 //y2=6.02
cc_2863 ( N_noxref_8_c_3313_n N_D_c_4972_n ) capacitor c=0.00581252f \
 //x=25.735 //y=5.2 //x2=25.53 //y2=4.7
cc_2864 ( N_noxref_8_c_3309_n N_CLK_c_5643_n ) capacitor c=0.0185297f \
 //x=26.445 //y=5.2 //x2=29.855 //y2=4.44
cc_2865 ( N_noxref_8_c_3313_n N_CLK_c_5643_n ) capacitor c=0.0181237f \
 //x=25.735 //y=5.2 //x2=29.855 //y2=4.44
cc_2866 ( N_noxref_8_c_3282_n N_CLK_c_5643_n ) capacitor c=0.0208321f \
 //x=27.01 //y=2.59 //x2=29.855 //y2=4.44
cc_2867 ( N_noxref_8_c_3284_n N_CLK_c_5643_n ) capacitor c=0.0208709f \
 //x=28.86 //y=2.08 //x2=29.855 //y2=4.44
cc_2868 ( N_noxref_8_c_3334_n N_CLK_c_5643_n ) capacitor c=0.0166984f \
 //x=29.135 //y=4.79 //x2=29.855 //y2=4.44
cc_2869 ( N_noxref_8_c_3285_n N_CLK_c_5668_n ) capacitor c=0.0208709f \
 //x=33.67 //y=2.08 //x2=39.105 //y2=4.44
cc_2870 ( N_noxref_8_c_3336_n N_CLK_c_5668_n ) capacitor c=0.0166984f \
 //x=33.945 //y=4.79 //x2=39.105 //y2=4.44
cc_2871 ( N_noxref_8_c_3284_n N_CLK_c_5679_n ) capacitor c=0.00153281f \
 //x=28.86 //y=2.08 //x2=30.085 //y2=4.44
cc_2872 ( N_noxref_8_c_3279_n N_CLK_c_5625_n ) capacitor c=0.0190006f \
 //x=33.555 //y=2.59 //x2=29.97 //y2=2.08
cc_2873 ( N_noxref_8_c_3280_n N_CLK_c_5625_n ) capacitor c=0.00103784f \
 //x=29.125 //y=2.59 //x2=29.97 //y2=2.08
cc_2874 ( N_noxref_8_c_3282_n N_CLK_c_5625_n ) capacitor c=3.63796e-19 \
 //x=27.01 //y=2.59 //x2=29.97 //y2=2.08
cc_2875 ( N_noxref_8_c_3284_n N_CLK_c_5625_n ) capacitor c=0.0435204f \
 //x=28.86 //y=2.08 //x2=29.97 //y2=2.08
cc_2876 ( N_noxref_8_c_3290_n N_CLK_c_5625_n ) capacitor c=0.00210802f \
 //x=28.56 //y=1.915 //x2=29.97 //y2=2.08
cc_2877 ( N_noxref_8_c_3367_p N_CLK_c_5625_n ) capacitor c=0.00147352f \
 //x=29.425 //y=4.79 //x2=29.97 //y2=2.08
cc_2878 ( N_noxref_8_c_3334_n N_CLK_c_5625_n ) capacitor c=0.00141297f \
 //x=29.135 //y=4.79 //x2=29.97 //y2=2.08
cc_2879 ( N_noxref_8_M86_noxref_g N_CLK_M88_noxref_g ) capacitor c=0.0105869f \
 //x=29.06 //y=6.02 //x2=29.94 //y2=6.02
cc_2880 ( N_noxref_8_M87_noxref_g N_CLK_M88_noxref_g ) capacitor c=0.10632f \
 //x=29.5 //y=6.02 //x2=29.94 //y2=6.02
cc_2881 ( N_noxref_8_M87_noxref_g N_CLK_M89_noxref_g ) capacitor c=0.0101598f \
 //x=29.5 //y=6.02 //x2=30.38 //y2=6.02
cc_2882 ( N_noxref_8_c_3286_n N_CLK_c_5926_n ) capacitor c=5.72482e-19 \
 //x=28.56 //y=0.875 //x2=29.535 //y2=0.91
cc_2883 ( N_noxref_8_c_3288_n N_CLK_c_5926_n ) capacitor c=0.00149976f \
 //x=28.56 //y=1.22 //x2=29.535 //y2=0.91
cc_2884 ( N_noxref_8_c_3293_n N_CLK_c_5926_n ) capacitor c=0.0160123f \
 //x=29.09 //y=0.875 //x2=29.535 //y2=0.91
cc_2885 ( N_noxref_8_c_3289_n N_CLK_c_5929_n ) capacitor c=0.00111227f \
 //x=28.56 //y=1.53 //x2=29.535 //y2=1.22
cc_2886 ( N_noxref_8_c_3295_n N_CLK_c_5929_n ) capacitor c=0.0124075f \
 //x=29.09 //y=1.22 //x2=29.535 //y2=1.22
cc_2887 ( N_noxref_8_c_3293_n N_CLK_c_5931_n ) capacitor c=0.00103227f \
 //x=29.09 //y=0.875 //x2=30.06 //y2=0.91
cc_2888 ( N_noxref_8_c_3295_n N_CLK_c_5932_n ) capacitor c=0.0010154f \
 //x=29.09 //y=1.22 //x2=30.06 //y2=1.22
cc_2889 ( N_noxref_8_c_3295_n N_CLK_c_5933_n ) capacitor c=9.23422e-19 \
 //x=29.09 //y=1.22 //x2=30.06 //y2=1.45
cc_2890 ( N_noxref_8_c_3284_n N_CLK_c_5934_n ) capacitor c=0.00203769f \
 //x=28.86 //y=2.08 //x2=30.06 //y2=1.915
cc_2891 ( N_noxref_8_c_3290_n N_CLK_c_5934_n ) capacitor c=0.00834532f \
 //x=28.56 //y=1.915 //x2=30.06 //y2=1.915
cc_2892 ( N_noxref_8_c_3284_n N_CLK_c_5936_n ) capacitor c=0.00183762f \
 //x=28.86 //y=2.08 //x2=29.97 //y2=4.7
cc_2893 ( N_noxref_8_c_3367_p N_CLK_c_5936_n ) capacitor c=0.0168581f \
 //x=29.425 //y=4.79 //x2=29.97 //y2=4.7
cc_2894 ( N_noxref_8_c_3334_n N_CLK_c_5936_n ) capacitor c=0.00484466f \
 //x=29.135 //y=4.79 //x2=29.97 //y2=4.7
cc_2895 ( N_noxref_8_c_3277_n N_SN_c_6844_n ) capacitor c=0.140806f //x=28.715 \
 //y=2.59 //x2=34.665 //y2=2.22
cc_2896 ( N_noxref_8_c_3278_n N_SN_c_6844_n ) capacitor c=0.0290445f \
 //x=27.125 //y=2.59 //x2=34.665 //y2=2.22
cc_2897 ( N_noxref_8_c_3279_n N_SN_c_6844_n ) capacitor c=0.414292f //x=33.555 \
 //y=2.59 //x2=34.665 //y2=2.22
cc_2898 ( N_noxref_8_c_3280_n N_SN_c_6844_n ) capacitor c=0.0429267f \
 //x=29.125 //y=2.59 //x2=34.665 //y2=2.22
cc_2899 ( N_noxref_8_c_3444_p N_SN_c_6844_n ) capacitor c=0.0146822f \
 //x=26.655 //y=1.655 //x2=34.665 //y2=2.22
cc_2900 ( N_noxref_8_c_3282_n N_SN_c_6844_n ) capacitor c=0.0217395f //x=27.01 \
 //y=2.59 //x2=34.665 //y2=2.22
cc_2901 ( N_noxref_8_c_3284_n N_SN_c_6844_n ) capacitor c=0.0211309f //x=28.86 \
 //y=2.08 //x2=34.665 //y2=2.22
cc_2902 ( N_noxref_8_c_3285_n N_SN_c_6844_n ) capacitor c=0.021104f //x=33.67 \
 //y=2.08 //x2=34.665 //y2=2.22
cc_2903 ( N_noxref_8_c_3290_n N_SN_c_6844_n ) capacitor c=0.011987f //x=28.56 \
 //y=1.915 //x2=34.665 //y2=2.22
cc_2904 ( N_noxref_8_c_3300_n N_SN_c_6844_n ) capacitor c=0.011987f //x=33.37 \
 //y=1.915 //x2=34.665 //y2=2.22
cc_2905 ( N_noxref_8_c_3285_n N_SN_c_6865_n ) capacitor c=0.00165648f \
 //x=33.67 //y=2.08 //x2=34.895 //y2=2.22
cc_2906 ( N_noxref_8_c_3300_n N_SN_c_6865_n ) capacitor c=2.3323e-19 //x=33.37 \
 //y=1.915 //x2=34.895 //y2=2.22
cc_2907 ( N_noxref_8_c_3279_n N_SN_c_6890_n ) capacitor c=0.00311593f \
 //x=33.555 //y=2.59 //x2=34.78 //y2=2.08
cc_2908 ( N_noxref_8_c_3285_n N_SN_c_6890_n ) capacitor c=0.0428203f //x=33.67 \
 //y=2.08 //x2=34.78 //y2=2.08
cc_2909 ( N_noxref_8_c_3300_n N_SN_c_6890_n ) capacitor c=0.00208635f \
 //x=33.37 //y=1.915 //x2=34.78 //y2=2.08
cc_2910 ( N_noxref_8_c_3352_p N_SN_c_6890_n ) capacitor c=0.00147352f \
 //x=34.235 //y=4.79 //x2=34.78 //y2=2.08
cc_2911 ( N_noxref_8_c_3336_n N_SN_c_6890_n ) capacitor c=0.00142741f \
 //x=33.945 //y=4.79 //x2=34.78 //y2=2.08
cc_2912 ( N_noxref_8_M92_noxref_g N_SN_M94_noxref_g ) capacitor c=0.0105869f \
 //x=33.87 //y=6.02 //x2=34.75 //y2=6.02
cc_2913 ( N_noxref_8_M93_noxref_g N_SN_M94_noxref_g ) capacitor c=0.10632f \
 //x=34.31 //y=6.02 //x2=34.75 //y2=6.02
cc_2914 ( N_noxref_8_M93_noxref_g N_SN_M95_noxref_g ) capacitor c=0.0101598f \
 //x=34.31 //y=6.02 //x2=35.19 //y2=6.02
cc_2915 ( N_noxref_8_c_3296_n N_SN_c_7070_n ) capacitor c=5.72482e-19 \
 //x=33.37 //y=0.875 //x2=34.345 //y2=0.91
cc_2916 ( N_noxref_8_c_3298_n N_SN_c_7070_n ) capacitor c=0.00149976f \
 //x=33.37 //y=1.22 //x2=34.345 //y2=0.91
cc_2917 ( N_noxref_8_c_3303_n N_SN_c_7070_n ) capacitor c=0.0160123f //x=33.9 \
 //y=0.875 //x2=34.345 //y2=0.91
cc_2918 ( N_noxref_8_c_3299_n N_SN_c_7073_n ) capacitor c=0.00111227f \
 //x=33.37 //y=1.53 //x2=34.345 //y2=1.22
cc_2919 ( N_noxref_8_c_3305_n N_SN_c_7073_n ) capacitor c=0.0124075f //x=33.9 \
 //y=1.22 //x2=34.345 //y2=1.22
cc_2920 ( N_noxref_8_c_3303_n N_SN_c_7075_n ) capacitor c=0.00103227f //x=33.9 \
 //y=0.875 //x2=34.87 //y2=0.91
cc_2921 ( N_noxref_8_c_3305_n N_SN_c_7076_n ) capacitor c=0.0010154f //x=33.9 \
 //y=1.22 //x2=34.87 //y2=1.22
cc_2922 ( N_noxref_8_c_3305_n N_SN_c_7077_n ) capacitor c=9.23422e-19 //x=33.9 \
 //y=1.22 //x2=34.87 //y2=1.45
cc_2923 ( N_noxref_8_c_3285_n N_SN_c_7078_n ) capacitor c=0.00203769f \
 //x=33.67 //y=2.08 //x2=34.87 //y2=1.915
cc_2924 ( N_noxref_8_c_3300_n N_SN_c_7078_n ) capacitor c=0.00834532f \
 //x=33.37 //y=1.915 //x2=34.87 //y2=1.915
cc_2925 ( N_noxref_8_c_3285_n N_SN_c_7080_n ) capacitor c=0.00183762f \
 //x=33.67 //y=2.08 //x2=34.78 //y2=4.7
cc_2926 ( N_noxref_8_c_3352_p N_SN_c_7080_n ) capacitor c=0.0168581f \
 //x=34.235 //y=4.79 //x2=34.78 //y2=4.7
cc_2927 ( N_noxref_8_c_3336_n N_SN_c_7080_n ) capacitor c=0.00484466f \
 //x=33.945 //y=4.79 //x2=34.78 //y2=4.7
cc_2928 ( N_noxref_8_c_3277_n N_noxref_24_c_8424_n ) capacitor c=0.0111379f \
 //x=28.715 //y=2.59 //x2=79.065 //y2=3.33
cc_2929 ( N_noxref_8_c_3278_n N_noxref_24_c_8424_n ) capacitor c=8.86511e-19 \
 //x=27.125 //y=2.59 //x2=79.065 //y2=3.33
cc_2930 ( N_noxref_8_c_3279_n N_noxref_24_c_8424_n ) capacitor c=7.63975e-19 \
 //x=33.555 //y=2.59 //x2=79.065 //y2=3.33
cc_2931 ( N_noxref_8_c_3280_n N_noxref_24_c_8424_n ) capacitor c=0.036868f \
 //x=29.125 //y=2.59 //x2=79.065 //y2=3.33
cc_2932 ( N_noxref_8_c_3282_n N_noxref_24_c_8424_n ) capacitor c=0.0211091f \
 //x=27.01 //y=2.59 //x2=79.065 //y2=3.33
cc_2933 ( N_noxref_8_c_3284_n N_noxref_24_c_8424_n ) capacitor c=0.0221447f \
 //x=28.86 //y=2.08 //x2=79.065 //y2=3.33
cc_2934 ( N_noxref_8_c_3285_n N_noxref_24_c_8424_n ) capacitor c=0.0197803f \
 //x=33.67 //y=2.08 //x2=79.065 //y2=3.33
cc_2935 ( N_noxref_8_c_3282_n N_noxref_24_c_8465_n ) capacitor c=3.52729e-19 \
 //x=27.01 //y=2.59 //x2=23.68 //y2=3.33
cc_2936 ( N_noxref_8_c_3444_p N_noxref_36_c_9710_n ) capacitor c=3.15806e-19 \
 //x=26.655 //y=1.655 //x2=25.115 //y2=1.495
cc_2937 ( N_noxref_8_c_3444_p N_noxref_36_c_9699_n ) capacitor c=0.020324f \
 //x=26.655 //y=1.655 //x2=26.085 //y2=1.495
cc_2938 ( N_noxref_8_c_3281_n N_noxref_36_c_9700_n ) capacitor c=0.00457164f \
 //x=26.925 //y=1.655 //x2=26.97 //y2=0.53
cc_2939 ( N_noxref_8_M16_noxref_d N_noxref_36_c_9700_n ) capacitor \
 c=0.0115831f //x=26.38 //y=0.905 //x2=26.97 //y2=0.53
cc_2940 ( N_noxref_8_c_3281_n N_noxref_36_M15_noxref_s ) capacitor \
 c=0.0126484f //x=26.925 //y=1.655 //x2=24.98 //y2=0.365
cc_2941 ( N_noxref_8_M16_noxref_d N_noxref_36_M15_noxref_s ) capacitor \
 c=0.0439476f //x=26.38 //y=0.905 //x2=24.98 //y2=0.365
cc_2942 ( N_noxref_8_c_3281_n N_noxref_37_c_9758_n ) capacitor c=4.08644e-19 \
 //x=26.925 //y=1.655 //x2=28.34 //y2=1.505
cc_2943 ( N_noxref_8_c_3290_n N_noxref_37_c_9758_n ) capacitor c=0.0034165f \
 //x=28.56 //y=1.915 //x2=28.34 //y2=1.505
cc_2944 ( N_noxref_8_c_3284_n N_noxref_37_c_9743_n ) capacitor c=0.0115578f \
 //x=28.86 //y=2.08 //x2=29.225 //y2=1.59
cc_2945 ( N_noxref_8_c_3289_n N_noxref_37_c_9743_n ) capacitor c=0.00697148f \
 //x=28.56 //y=1.53 //x2=29.225 //y2=1.59
cc_2946 ( N_noxref_8_c_3290_n N_noxref_37_c_9743_n ) capacitor c=0.0204849f \
 //x=28.56 //y=1.915 //x2=29.225 //y2=1.59
cc_2947 ( N_noxref_8_c_3292_n N_noxref_37_c_9743_n ) capacitor c=0.00610316f \
 //x=28.935 //y=1.375 //x2=29.225 //y2=1.59
cc_2948 ( N_noxref_8_c_3295_n N_noxref_37_c_9743_n ) capacitor c=0.00698822f \
 //x=29.09 //y=1.22 //x2=29.225 //y2=1.59
cc_2949 ( N_noxref_8_c_3286_n N_noxref_37_M17_noxref_s ) capacitor \
 c=0.0327271f //x=28.56 //y=0.875 //x2=28.205 //y2=0.375
cc_2950 ( N_noxref_8_c_3289_n N_noxref_37_M17_noxref_s ) capacitor \
 c=7.99997e-19 //x=28.56 //y=1.53 //x2=28.205 //y2=0.375
cc_2951 ( N_noxref_8_c_3290_n N_noxref_37_M17_noxref_s ) capacitor \
 c=0.00122123f //x=28.56 //y=1.915 //x2=28.205 //y2=0.375
cc_2952 ( N_noxref_8_c_3293_n N_noxref_37_M17_noxref_s ) capacitor \
 c=0.0121427f //x=29.09 //y=0.875 //x2=28.205 //y2=0.375
cc_2953 ( N_noxref_8_M16_noxref_d N_noxref_37_M17_noxref_s ) capacitor \
 c=2.53688e-19 //x=26.38 //y=0.905 //x2=28.205 //y2=0.375
cc_2954 ( N_noxref_8_c_3300_n N_noxref_39_c_9859_n ) capacitor c=0.0034165f \
 //x=33.37 //y=1.915 //x2=33.15 //y2=1.505
cc_2955 ( N_noxref_8_c_3285_n N_noxref_39_c_9844_n ) capacitor c=0.0115578f \
 //x=33.67 //y=2.08 //x2=34.035 //y2=1.59
cc_2956 ( N_noxref_8_c_3299_n N_noxref_39_c_9844_n ) capacitor c=0.00697148f \
 //x=33.37 //y=1.53 //x2=34.035 //y2=1.59
cc_2957 ( N_noxref_8_c_3300_n N_noxref_39_c_9844_n ) capacitor c=0.0204849f \
 //x=33.37 //y=1.915 //x2=34.035 //y2=1.59
cc_2958 ( N_noxref_8_c_3302_n N_noxref_39_c_9844_n ) capacitor c=0.00610316f \
 //x=33.745 //y=1.375 //x2=34.035 //y2=1.59
cc_2959 ( N_noxref_8_c_3305_n N_noxref_39_c_9844_n ) capacitor c=0.00698822f \
 //x=33.9 //y=1.22 //x2=34.035 //y2=1.59
cc_2960 ( N_noxref_8_c_3296_n N_noxref_39_M20_noxref_s ) capacitor \
 c=0.0327271f //x=33.37 //y=0.875 //x2=33.015 //y2=0.375
cc_2961 ( N_noxref_8_c_3299_n N_noxref_39_M20_noxref_s ) capacitor \
 c=7.99997e-19 //x=33.37 //y=1.53 //x2=33.015 //y2=0.375
cc_2962 ( N_noxref_8_c_3300_n N_noxref_39_M20_noxref_s ) capacitor \
 c=0.00122123f //x=33.37 //y=1.915 //x2=33.015 //y2=0.375
cc_2963 ( N_noxref_8_c_3303_n N_noxref_39_M20_noxref_s ) capacitor \
 c=0.0121427f //x=33.9 //y=0.875 //x2=33.015 //y2=0.375
cc_2964 ( N_noxref_9_c_3512_n N_noxref_10_c_3691_n ) capacitor c=0.0181982f \
 //x=36.63 //y=2.59 //x2=41.695 //y2=4.07
cc_2965 ( N_noxref_9_c_3513_n N_noxref_10_c_3691_n ) capacitor c=0.0184765f \
 //x=38.48 //y=2.08 //x2=41.695 //y2=4.07
cc_2966 ( N_noxref_9_c_3529_n N_noxref_10_c_3707_n ) capacitor c=3.10026e-19 \
 //x=34.175 //y=5.155 //x2=31.735 //y2=5.155
cc_2967 ( N_noxref_9_c_3512_n N_noxref_12_c_4162_n ) capacitor c=0.0187698f \
 //x=36.63 //y=2.59 //x2=39.845 //y2=3.7
cc_2968 ( N_noxref_9_c_3513_n N_noxref_12_c_4162_n ) capacitor c=0.0187484f \
 //x=38.48 //y=2.08 //x2=39.845 //y2=3.7
cc_2969 ( N_noxref_9_c_3512_n N_noxref_12_c_4164_n ) capacitor c=0.00117715f \
 //x=36.63 //y=2.59 //x2=36.005 //y2=3.7
cc_2970 ( N_noxref_9_c_3510_n N_noxref_12_c_4112_n ) capacitor c=0.00456439f \
 //x=36.745 //y=2.59 //x2=35.89 //y2=2.08
cc_2971 ( N_noxref_9_c_3512_n N_noxref_12_c_4112_n ) capacitor c=0.076937f \
 //x=36.63 //y=2.59 //x2=35.89 //y2=2.08
cc_2972 ( N_noxref_9_c_3513_n N_noxref_12_c_4112_n ) capacitor c=5.32619e-19 \
 //x=38.48 //y=2.08 //x2=35.89 //y2=2.08
cc_2973 ( N_noxref_9_c_3577_p N_noxref_12_c_4112_n ) capacitor c=0.016476f \
 //x=35.85 //y=5.155 //x2=35.89 //y2=2.08
cc_2974 ( N_noxref_9_M99_noxref_g N_noxref_12_c_4121_n ) capacitor \
 c=0.0169521f //x=38.82 //y=6.02 //x2=39.395 //y2=5.2
cc_2975 ( N_noxref_9_c_3513_n N_noxref_12_c_4125_n ) capacitor c=0.00539951f \
 //x=38.48 //y=2.08 //x2=38.685 //y2=5.2
cc_2976 ( N_noxref_9_M98_noxref_g N_noxref_12_c_4125_n ) capacitor \
 c=0.0177326f //x=38.38 //y=6.02 //x2=38.685 //y2=5.2
cc_2977 ( N_noxref_9_c_3547_n N_noxref_12_c_4125_n ) capacitor c=0.00581252f \
 //x=38.48 //y=4.7 //x2=38.685 //y2=5.2
cc_2978 ( N_noxref_9_c_3512_n N_noxref_12_c_4114_n ) capacitor c=3.52729e-19 \
 //x=36.63 //y=2.59 //x2=39.96 //y2=3.7
cc_2979 ( N_noxref_9_c_3513_n N_noxref_12_c_4114_n ) capacitor c=0.00294763f \
 //x=38.48 //y=2.08 //x2=39.96 //y2=3.7
cc_2980 ( N_noxref_9_c_3531_n N_noxref_12_M96_noxref_g ) capacitor c=0.01736f \
 //x=35.765 //y=5.155 //x2=35.63 //y2=6.02
cc_2981 ( N_noxref_9_M96_noxref_d N_noxref_12_M96_noxref_g ) capacitor \
 c=0.0180032f //x=35.705 //y=5.02 //x2=35.63 //y2=6.02
cc_2982 ( N_noxref_9_c_3535_n N_noxref_12_M97_noxref_g ) capacitor \
 c=0.0194981f //x=36.545 //y=5.155 //x2=36.07 //y2=6.02
cc_2983 ( N_noxref_9_M96_noxref_d N_noxref_12_M97_noxref_g ) capacitor \
 c=0.0194246f //x=35.705 //y=5.02 //x2=36.07 //y2=6.02
cc_2984 ( N_noxref_9_M22_noxref_d N_noxref_12_c_4179_n ) capacitor \
 c=0.00217566f //x=35.955 //y=0.915 //x2=35.88 //y2=0.915
cc_2985 ( N_noxref_9_M22_noxref_d N_noxref_12_c_4180_n ) capacitor \
 c=0.0034598f //x=35.955 //y=0.915 //x2=35.88 //y2=1.26
cc_2986 ( N_noxref_9_M22_noxref_d N_noxref_12_c_4181_n ) capacitor \
 c=0.00546784f //x=35.955 //y=0.915 //x2=35.88 //y2=1.57
cc_2987 ( N_noxref_9_M22_noxref_d N_noxref_12_c_4182_n ) capacitor \
 c=0.00241102f //x=35.955 //y=0.915 //x2=36.255 //y2=0.76
cc_2988 ( N_noxref_9_c_3511_n N_noxref_12_c_4183_n ) capacitor c=0.00371277f \
 //x=36.545 //y=1.665 //x2=36.255 //y2=1.415
cc_2989 ( N_noxref_9_M22_noxref_d N_noxref_12_c_4183_n ) capacitor \
 c=0.0138621f //x=35.955 //y=0.915 //x2=36.255 //y2=1.415
cc_2990 ( N_noxref_9_M22_noxref_d N_noxref_12_c_4185_n ) capacitor \
 c=0.00219619f //x=35.955 //y=0.915 //x2=36.41 //y2=0.915
cc_2991 ( N_noxref_9_c_3511_n N_noxref_12_c_4186_n ) capacitor c=0.00457401f \
 //x=36.545 //y=1.665 //x2=36.41 //y2=1.26
cc_2992 ( N_noxref_9_M22_noxref_d N_noxref_12_c_4186_n ) capacitor \
 c=0.00603828f //x=35.955 //y=0.915 //x2=36.41 //y2=1.26
cc_2993 ( N_noxref_9_c_3512_n N_noxref_12_c_4188_n ) capacitor c=0.00709342f \
 //x=36.63 //y=2.59 //x2=35.89 //y2=2.08
cc_2994 ( N_noxref_9_c_3512_n N_noxref_12_c_4189_n ) capacitor c=0.00283672f \
 //x=36.63 //y=2.59 //x2=35.89 //y2=1.915
cc_2995 ( N_noxref_9_M22_noxref_d N_noxref_12_c_4189_n ) capacitor \
 c=0.00661782f //x=35.955 //y=0.915 //x2=35.89 //y2=1.915
cc_2996 ( N_noxref_9_c_3535_n N_noxref_12_c_4191_n ) capacitor c=0.00201851f \
 //x=36.545 //y=5.155 //x2=35.89 //y2=4.7
cc_2997 ( N_noxref_9_c_3512_n N_noxref_12_c_4191_n ) capacitor c=0.013693f \
 //x=36.63 //y=2.59 //x2=35.89 //y2=4.7
cc_2998 ( N_noxref_9_c_3577_p N_noxref_12_c_4191_n ) capacitor c=0.00475601f \
 //x=35.85 //y=5.155 //x2=35.89 //y2=4.7
cc_2999 ( N_noxref_9_M99_noxref_g N_noxref_12_M98_noxref_d ) capacitor \
 c=0.0173476f //x=38.82 //y=6.02 //x2=38.455 //y2=5.02
cc_3000 ( N_noxref_9_c_3509_n N_D_c_4909_n ) capacitor c=0.172364f //x=38.365 \
 //y=2.59 //x2=49.835 //y2=2.96
cc_3001 ( N_noxref_9_c_3510_n N_D_c_4909_n ) capacitor c=0.0293832f //x=36.745 \
 //y=2.59 //x2=49.835 //y2=2.96
cc_3002 ( N_noxref_9_c_3512_n N_D_c_4909_n ) capacitor c=0.0206007f //x=36.63 \
 //y=2.59 //x2=49.835 //y2=2.96
cc_3003 ( N_noxref_9_c_3513_n N_D_c_4909_n ) capacitor c=0.0205791f //x=38.48 \
 //y=2.08 //x2=49.835 //y2=2.96
cc_3004 ( N_noxref_9_c_3525_n N_CLK_c_5668_n ) capacitor c=0.032141f \
 //x=34.885 //y=5.155 //x2=39.105 //y2=4.44
cc_3005 ( N_noxref_9_c_3529_n N_CLK_c_5668_n ) capacitor c=0.0230136f \
 //x=34.175 //y=5.155 //x2=39.105 //y2=4.44
cc_3006 ( N_noxref_9_c_3535_n N_CLK_c_5668_n ) capacitor c=0.0183122f \
 //x=36.545 //y=5.155 //x2=39.105 //y2=4.44
cc_3007 ( N_noxref_9_c_3512_n N_CLK_c_5668_n ) capacitor c=0.0210274f \
 //x=36.63 //y=2.59 //x2=39.105 //y2=4.44
cc_3008 ( N_noxref_9_c_3513_n N_CLK_c_5668_n ) capacitor c=0.0198304f \
 //x=38.48 //y=2.08 //x2=39.105 //y2=4.44
cc_3009 ( N_noxref_9_c_3547_n N_CLK_c_5668_n ) capacitor c=0.0107057f \
 //x=38.48 //y=4.7 //x2=39.105 //y2=4.44
cc_3010 ( N_noxref_9_c_3513_n N_CLK_c_5704_n ) capacitor c=0.00168329f \
 //x=38.48 //y=2.08 //x2=39.335 //y2=4.44
cc_3011 ( N_noxref_9_c_3547_n N_CLK_c_5704_n ) capacitor c=2.91071e-19 \
 //x=38.48 //y=4.7 //x2=39.335 //y2=4.44
cc_3012 ( N_noxref_9_c_3513_n N_CLK_c_5947_n ) capacitor c=0.00400249f \
 //x=38.48 //y=2.08 //x2=39.22 //y2=4.535
cc_3013 ( N_noxref_9_c_3547_n N_CLK_c_5947_n ) capacitor c=0.00415951f \
 //x=38.48 //y=4.7 //x2=39.22 //y2=4.535
cc_3014 ( N_noxref_9_c_3509_n N_CLK_c_5626_n ) capacitor c=0.00720056f \
 //x=38.365 //y=2.59 //x2=39.22 //y2=2.08
cc_3015 ( N_noxref_9_c_3512_n N_CLK_c_5626_n ) capacitor c=6.41343e-19 \
 //x=36.63 //y=2.59 //x2=39.22 //y2=2.08
cc_3016 ( N_noxref_9_c_3513_n N_CLK_c_5626_n ) capacitor c=0.0712948f \
 //x=38.48 //y=2.08 //x2=39.22 //y2=2.08
cc_3017 ( N_noxref_9_c_3518_n N_CLK_c_5626_n ) capacitor c=0.00284029f \
 //x=38.285 //y=1.915 //x2=39.22 //y2=2.08
cc_3018 ( N_noxref_9_M98_noxref_g N_CLK_M100_noxref_g ) capacitor c=0.0104611f \
 //x=38.38 //y=6.02 //x2=39.26 //y2=6.02
cc_3019 ( N_noxref_9_M99_noxref_g N_CLK_M100_noxref_g ) capacitor c=0.106811f \
 //x=38.82 //y=6.02 //x2=39.26 //y2=6.02
cc_3020 ( N_noxref_9_M99_noxref_g N_CLK_M101_noxref_g ) capacitor c=0.0100341f \
 //x=38.82 //y=6.02 //x2=39.7 //y2=6.02
cc_3021 ( N_noxref_9_c_3514_n N_CLK_c_5956_n ) capacitor c=4.86506e-19 \
 //x=38.285 //y=0.865 //x2=39.255 //y2=0.905
cc_3022 ( N_noxref_9_c_3516_n N_CLK_c_5956_n ) capacitor c=0.00152104f \
 //x=38.285 //y=1.21 //x2=39.255 //y2=0.905
cc_3023 ( N_noxref_9_c_3521_n N_CLK_c_5956_n ) capacitor c=0.0151475f \
 //x=38.815 //y=0.865 //x2=39.255 //y2=0.905
cc_3024 ( N_noxref_9_c_3517_n N_CLK_c_5959_n ) capacitor c=0.00109982f \
 //x=38.285 //y=1.52 //x2=39.255 //y2=1.25
cc_3025 ( N_noxref_9_c_3523_n N_CLK_c_5959_n ) capacitor c=0.0111064f \
 //x=38.815 //y=1.21 //x2=39.255 //y2=1.25
cc_3026 ( N_noxref_9_c_3517_n N_CLK_c_5961_n ) capacitor c=9.57794e-19 \
 //x=38.285 //y=1.52 //x2=39.255 //y2=1.56
cc_3027 ( N_noxref_9_c_3518_n N_CLK_c_5961_n ) capacitor c=0.00662747f \
 //x=38.285 //y=1.915 //x2=39.255 //y2=1.56
cc_3028 ( N_noxref_9_c_3523_n N_CLK_c_5961_n ) capacitor c=0.00862358f \
 //x=38.815 //y=1.21 //x2=39.255 //y2=1.56
cc_3029 ( N_noxref_9_c_3521_n N_CLK_c_5964_n ) capacitor c=0.00124821f \
 //x=38.815 //y=0.865 //x2=39.785 //y2=0.905
cc_3030 ( N_noxref_9_c_3523_n N_CLK_c_5965_n ) capacitor c=0.00200715f \
 //x=38.815 //y=1.21 //x2=39.785 //y2=1.25
cc_3031 ( N_noxref_9_c_3513_n N_CLK_c_5966_n ) capacitor c=0.00282278f \
 //x=38.48 //y=2.08 //x2=39.22 //y2=2.08
cc_3032 ( N_noxref_9_c_3518_n N_CLK_c_5966_n ) capacitor c=0.0172771f \
 //x=38.285 //y=1.915 //x2=39.22 //y2=2.08
cc_3033 ( N_noxref_9_c_3513_n N_CLK_c_5968_n ) capacitor c=0.00342116f \
 //x=38.48 //y=2.08 //x2=39.25 //y2=4.7
cc_3034 ( N_noxref_9_c_3547_n N_CLK_c_5968_n ) capacitor c=0.0292158f \
 //x=38.48 //y=4.7 //x2=39.25 //y2=4.7
cc_3035 ( N_noxref_9_c_3509_n N_SN_c_6855_n ) capacitor c=0.172308f //x=38.365 \
 //y=2.59 //x2=46.135 //y2=2.22
cc_3036 ( N_noxref_9_c_3510_n N_SN_c_6855_n ) capacitor c=0.0291301f \
 //x=36.745 //y=2.59 //x2=46.135 //y2=2.22
cc_3037 ( N_noxref_9_c_3641_p N_SN_c_6855_n ) capacitor c=0.016327f //x=36.23 \
 //y=1.665 //x2=46.135 //y2=2.22
cc_3038 ( N_noxref_9_c_3512_n N_SN_c_6855_n ) capacitor c=0.0215653f //x=36.63 \
 //y=2.59 //x2=46.135 //y2=2.22
cc_3039 ( N_noxref_9_c_3513_n N_SN_c_6855_n ) capacitor c=0.0203358f //x=38.48 \
 //y=2.08 //x2=46.135 //y2=2.22
cc_3040 ( N_noxref_9_c_3518_n N_SN_c_6855_n ) capacitor c=0.00894156f \
 //x=38.285 //y=1.915 //x2=46.135 //y2=2.22
cc_3041 ( N_noxref_9_c_3525_n N_SN_c_6890_n ) capacitor c=0.0146f //x=34.885 \
 //y=5.155 //x2=34.78 //y2=2.08
cc_3042 ( N_noxref_9_c_3512_n N_SN_c_6890_n ) capacitor c=0.00237834f \
 //x=36.63 //y=2.59 //x2=34.78 //y2=2.08
cc_3043 ( N_noxref_9_c_3525_n N_SN_M94_noxref_g ) capacitor c=0.0165266f \
 //x=34.885 //y=5.155 //x2=34.75 //y2=6.02
cc_3044 ( N_noxref_9_M94_noxref_d N_SN_M94_noxref_g ) capacitor c=0.0180032f \
 //x=34.825 //y=5.02 //x2=34.75 //y2=6.02
cc_3045 ( N_noxref_9_c_3531_n N_SN_M95_noxref_g ) capacitor c=0.01736f \
 //x=35.765 //y=5.155 //x2=35.19 //y2=6.02
cc_3046 ( N_noxref_9_M94_noxref_d N_SN_M95_noxref_g ) capacitor c=0.0180032f \
 //x=34.825 //y=5.02 //x2=35.19 //y2=6.02
cc_3047 ( N_noxref_9_c_3651_p N_SN_c_7095_n ) capacitor c=0.00426767f \
 //x=34.97 //y=5.155 //x2=35.115 //y2=4.79
cc_3048 ( N_noxref_9_c_3525_n N_SN_c_7080_n ) capacitor c=0.00322054f \
 //x=34.885 //y=5.155 //x2=34.78 //y2=4.7
cc_3049 ( N_noxref_9_c_3509_n N_noxref_24_c_8424_n ) capacitor c=0.0125435f \
 //x=38.365 //y=2.59 //x2=79.065 //y2=3.33
cc_3050 ( N_noxref_9_c_3510_n N_noxref_24_c_8424_n ) capacitor c=8.87672e-19 \
 //x=36.745 //y=2.59 //x2=79.065 //y2=3.33
cc_3051 ( N_noxref_9_c_3512_n N_noxref_24_c_8424_n ) capacitor c=0.018769f \
 //x=36.63 //y=2.59 //x2=79.065 //y2=3.33
cc_3052 ( N_noxref_9_c_3513_n N_noxref_24_c_8424_n ) capacitor c=0.0187666f \
 //x=38.48 //y=2.08 //x2=79.065 //y2=3.33
cc_3053 ( N_noxref_9_M22_noxref_d N_noxref_39_M20_noxref_s ) capacitor \
 c=0.00309936f //x=35.955 //y=0.915 //x2=33.015 //y2=0.375
cc_3054 ( N_noxref_9_c_3511_n N_noxref_40_c_9901_n ) capacitor c=0.00457167f \
 //x=36.545 //y=1.665 //x2=36.545 //y2=0.54
cc_3055 ( N_noxref_9_M22_noxref_d N_noxref_40_c_9901_n ) capacitor \
 c=0.0115903f //x=35.955 //y=0.915 //x2=36.545 //y2=0.54
cc_3056 ( N_noxref_9_c_3641_p N_noxref_40_c_9911_n ) capacitor c=0.020048f \
 //x=36.23 //y=1.665 //x2=35.66 //y2=0.995
cc_3057 ( N_noxref_9_M22_noxref_d N_noxref_40_M21_noxref_d ) capacitor \
 c=5.27807e-19 //x=35.955 //y=0.915 //x2=34.42 //y2=0.91
cc_3058 ( N_noxref_9_c_3511_n N_noxref_40_M22_noxref_s ) capacitor \
 c=0.0184051f //x=36.545 //y=1.665 //x2=35.525 //y2=0.375
cc_3059 ( N_noxref_9_M22_noxref_d N_noxref_40_M22_noxref_s ) capacitor \
 c=0.0426444f //x=35.955 //y=0.915 //x2=35.525 //y2=0.375
cc_3060 ( N_noxref_9_c_3511_n N_noxref_41_c_9966_n ) capacitor c=3.04182e-19 \
 //x=36.545 //y=1.665 //x2=38.065 //y2=1.495
cc_3061 ( N_noxref_9_c_3518_n N_noxref_41_c_9966_n ) capacitor c=0.0034165f \
 //x=38.285 //y=1.915 //x2=38.065 //y2=1.495
cc_3062 ( N_noxref_9_c_3513_n N_noxref_41_c_9948_n ) capacitor c=0.0111916f \
 //x=38.48 //y=2.08 //x2=38.95 //y2=1.58
cc_3063 ( N_noxref_9_c_3517_n N_noxref_41_c_9948_n ) capacitor c=0.00696403f \
 //x=38.285 //y=1.52 //x2=38.95 //y2=1.58
cc_3064 ( N_noxref_9_c_3518_n N_noxref_41_c_9948_n ) capacitor c=0.0174694f \
 //x=38.285 //y=1.915 //x2=38.95 //y2=1.58
cc_3065 ( N_noxref_9_c_3520_n N_noxref_41_c_9948_n ) capacitor c=0.00776811f \
 //x=38.66 //y=1.365 //x2=38.95 //y2=1.58
cc_3066 ( N_noxref_9_c_3523_n N_noxref_41_c_9948_n ) capacitor c=0.00339872f \
 //x=38.815 //y=1.21 //x2=38.95 //y2=1.58
cc_3067 ( N_noxref_9_c_3518_n N_noxref_41_c_9955_n ) capacitor c=6.71402e-19 \
 //x=38.285 //y=1.915 //x2=39.035 //y2=1.495
cc_3068 ( N_noxref_9_c_3514_n N_noxref_41_M23_noxref_s ) capacitor \
 c=0.0327502f //x=38.285 //y=0.865 //x2=37.93 //y2=0.365
cc_3069 ( N_noxref_9_c_3517_n N_noxref_41_M23_noxref_s ) capacitor \
 c=3.48408e-19 //x=38.285 //y=1.52 //x2=37.93 //y2=0.365
cc_3070 ( N_noxref_9_c_3521_n N_noxref_41_M23_noxref_s ) capacitor \
 c=0.0120759f //x=38.815 //y=0.865 //x2=37.93 //y2=0.365
cc_3071 ( N_noxref_10_M103_noxref_g N_noxref_11_c_3975_n ) capacitor \
 c=0.0169521f //x=42.15 //y=6.02 //x2=42.725 //y2=5.2
cc_3072 ( N_noxref_10_c_3678_n N_noxref_11_c_3979_n ) capacitor c=0.00521572f \
 //x=41.81 //y=2.08 //x2=42.015 //y2=5.2
cc_3073 ( N_noxref_10_M102_noxref_g N_noxref_11_c_3979_n ) capacitor \
 c=0.0177326f //x=41.71 //y=6.02 //x2=42.015 //y2=5.2
cc_3074 ( N_noxref_10_c_3724_n N_noxref_11_c_3979_n ) capacitor c=0.00581252f \
 //x=41.81 //y=4.7 //x2=42.015 //y2=5.2
cc_3075 ( N_noxref_10_c_3678_n N_noxref_11_c_3959_n ) capacitor c=0.00286703f \
 //x=41.81 //y=2.08 //x2=43.29 //y2=2.59
cc_3076 ( N_noxref_10_M103_noxref_g N_noxref_11_M102_noxref_d ) capacitor \
 c=0.0173476f //x=42.15 //y=6.02 //x2=41.785 //y2=5.02
cc_3077 ( N_noxref_10_c_3690_n N_noxref_12_c_4157_n ) capacitor c=0.044143f \
 //x=31.7 //y=4.07 //x2=35.775 //y2=3.7
cc_3078 ( N_noxref_10_c_3691_n N_noxref_12_c_4157_n ) capacitor c=0.340271f \
 //x=41.695 //y=4.07 //x2=35.775 //y2=3.7
cc_3079 ( N_noxref_10_c_3694_n N_noxref_12_c_4157_n ) capacitor c=0.0267581f \
 //x=31.93 //y=4.07 //x2=35.775 //y2=3.7
cc_3080 ( N_noxref_10_c_3714_n N_noxref_12_c_4157_n ) capacitor c=0.00219785f \
 //x=31.815 //y=4.07 //x2=35.775 //y2=3.7
cc_3081 ( N_noxref_10_c_3754_n N_noxref_12_c_4157_n ) capacitor c=0.0185057f \
 //x=31.817 //y=3.905 //x2=35.775 //y2=3.7
cc_3082 ( N_noxref_10_c_3690_n N_noxref_12_c_4200_n ) capacitor c=0.0292842f \
 //x=31.7 //y=4.07 //x2=31.195 //y2=3.7
cc_3083 ( N_noxref_10_c_3754_n N_noxref_12_c_4200_n ) capacitor c=0.00179385f \
 //x=31.817 //y=3.905 //x2=31.195 //y2=3.7
cc_3084 ( N_noxref_10_c_3691_n N_noxref_12_c_4162_n ) capacitor c=0.339174f \
 //x=41.695 //y=4.07 //x2=39.845 //y2=3.7
cc_3085 ( N_noxref_10_c_3691_n N_noxref_12_c_4164_n ) capacitor c=0.026596f \
 //x=41.695 //y=4.07 //x2=36.005 //y2=3.7
cc_3086 ( N_noxref_10_c_3691_n N_noxref_12_c_4204_n ) capacitor c=0.17615f \
 //x=41.695 //y=4.07 //x2=47.245 //y2=3.7
cc_3087 ( N_noxref_10_c_3678_n N_noxref_12_c_4204_n ) capacitor c=0.0205593f \
 //x=41.81 //y=2.08 //x2=47.245 //y2=3.7
cc_3088 ( N_noxref_10_c_3691_n N_noxref_12_c_4206_n ) capacitor c=0.026743f \
 //x=41.695 //y=4.07 //x2=40.075 //y2=3.7
cc_3089 ( N_noxref_10_c_3678_n N_noxref_12_c_4206_n ) capacitor c=7.01366e-19 \
 //x=41.81 //y=2.08 //x2=40.075 //y2=3.7
cc_3090 ( N_noxref_10_c_3690_n N_noxref_12_c_4111_n ) capacitor c=0.0197867f \
 //x=31.7 //y=4.07 //x2=31.08 //y2=2.08
cc_3091 ( N_noxref_10_c_3694_n N_noxref_12_c_4111_n ) capacitor c=0.00180189f \
 //x=31.93 //y=4.07 //x2=31.08 //y2=2.08
cc_3092 ( N_noxref_10_c_3801_p N_noxref_12_c_4111_n ) capacitor c=0.0163236f \
 //x=31.82 //y=5.07 //x2=31.08 //y2=2.08
cc_3093 ( N_noxref_10_c_3802_p N_noxref_12_c_4111_n ) capacitor c=0.016476f \
 //x=31.04 //y=5.155 //x2=31.08 //y2=2.08
cc_3094 ( N_noxref_10_c_3714_n N_noxref_12_c_4111_n ) capacitor c=0.00966503f \
 //x=31.815 //y=4.07 //x2=31.08 //y2=2.08
cc_3095 ( N_noxref_10_c_3754_n N_noxref_12_c_4111_n ) capacitor c=0.0508802f \
 //x=31.817 //y=3.905 //x2=31.08 //y2=2.08
cc_3096 ( N_noxref_10_c_3691_n N_noxref_12_c_4112_n ) capacitor c=0.0198068f \
 //x=41.695 //y=4.07 //x2=35.89 //y2=2.08
cc_3097 ( N_noxref_10_c_3691_n N_noxref_12_c_4114_n ) capacitor c=0.020307f \
 //x=41.695 //y=4.07 //x2=39.96 //y2=3.7
cc_3098 ( N_noxref_10_c_3678_n N_noxref_12_c_4114_n ) capacitor c=0.0112452f \
 //x=41.81 //y=2.08 //x2=39.96 //y2=3.7
cc_3099 ( N_noxref_10_c_3703_n N_noxref_12_M90_noxref_g ) capacitor c=0.01736f \
 //x=30.955 //y=5.155 //x2=30.82 //y2=6.02
cc_3100 ( N_noxref_10_M90_noxref_d N_noxref_12_M90_noxref_g ) capacitor \
 c=0.0180032f //x=30.895 //y=5.02 //x2=30.82 //y2=6.02
cc_3101 ( N_noxref_10_c_3707_n N_noxref_12_M91_noxref_g ) capacitor \
 c=0.0194981f //x=31.735 //y=5.155 //x2=31.26 //y2=6.02
cc_3102 ( N_noxref_10_M90_noxref_d N_noxref_12_M91_noxref_g ) capacitor \
 c=0.0194246f //x=30.895 //y=5.02 //x2=31.26 //y2=6.02
cc_3103 ( N_noxref_10_M19_noxref_d N_noxref_12_c_4221_n ) capacitor \
 c=0.00217566f //x=31.145 //y=0.915 //x2=31.07 //y2=0.915
cc_3104 ( N_noxref_10_M19_noxref_d N_noxref_12_c_4222_n ) capacitor \
 c=0.0034598f //x=31.145 //y=0.915 //x2=31.07 //y2=1.26
cc_3105 ( N_noxref_10_M19_noxref_d N_noxref_12_c_4223_n ) capacitor \
 c=0.00546784f //x=31.145 //y=0.915 //x2=31.07 //y2=1.57
cc_3106 ( N_noxref_10_M19_noxref_d N_noxref_12_c_4224_n ) capacitor \
 c=0.00241102f //x=31.145 //y=0.915 //x2=31.445 //y2=0.76
cc_3107 ( N_noxref_10_c_3677_n N_noxref_12_c_4225_n ) capacitor c=0.00371277f \
 //x=31.735 //y=1.665 //x2=31.445 //y2=1.415
cc_3108 ( N_noxref_10_M19_noxref_d N_noxref_12_c_4225_n ) capacitor \
 c=0.0138621f //x=31.145 //y=0.915 //x2=31.445 //y2=1.415
cc_3109 ( N_noxref_10_M19_noxref_d N_noxref_12_c_4227_n ) capacitor \
 c=0.00219619f //x=31.145 //y=0.915 //x2=31.6 //y2=0.915
cc_3110 ( N_noxref_10_c_3677_n N_noxref_12_c_4228_n ) capacitor c=0.00457401f \
 //x=31.735 //y=1.665 //x2=31.6 //y2=1.26
cc_3111 ( N_noxref_10_M19_noxref_d N_noxref_12_c_4228_n ) capacitor \
 c=0.00603828f //x=31.145 //y=0.915 //x2=31.6 //y2=1.26
cc_3112 ( N_noxref_10_c_3754_n N_noxref_12_c_4230_n ) capacitor c=0.00709342f \
 //x=31.817 //y=3.905 //x2=31.08 //y2=2.08
cc_3113 ( N_noxref_10_c_3754_n N_noxref_12_c_4231_n ) capacitor c=0.00404774f \
 //x=31.817 //y=3.905 //x2=31.08 //y2=1.915
cc_3114 ( N_noxref_10_M19_noxref_d N_noxref_12_c_4231_n ) capacitor \
 c=0.00661782f //x=31.145 //y=0.915 //x2=31.08 //y2=1.915
cc_3115 ( N_noxref_10_c_3707_n N_noxref_12_c_4233_n ) capacitor c=0.00201851f \
 //x=31.735 //y=5.155 //x2=31.08 //y2=4.7
cc_3116 ( N_noxref_10_c_3801_p N_noxref_12_c_4233_n ) capacitor c=0.0151148f \
 //x=31.82 //y=5.07 //x2=31.08 //y2=4.7
cc_3117 ( N_noxref_10_c_3802_p N_noxref_12_c_4233_n ) capacitor c=0.00475601f \
 //x=31.04 //y=5.155 //x2=31.08 //y2=4.7
cc_3118 ( N_noxref_10_c_3691_n N_noxref_13_c_4513_n ) capacitor c=0.0244534f \
 //x=41.695 //y=4.07 //x2=42.665 //y2=4.07
cc_3119 ( N_noxref_10_c_3678_n N_noxref_13_c_4513_n ) capacitor c=0.00246068f \
 //x=41.81 //y=2.08 //x2=42.665 //y2=4.07
cc_3120 ( N_noxref_10_c_3678_n N_noxref_13_c_4515_n ) capacitor c=0.00400249f \
 //x=41.81 //y=2.08 //x2=42.55 //y2=4.535
cc_3121 ( N_noxref_10_c_3724_n N_noxref_13_c_4515_n ) capacitor c=0.00417994f \
 //x=41.81 //y=4.7 //x2=42.55 //y2=4.535
cc_3122 ( N_noxref_10_c_3691_n N_noxref_13_c_4445_n ) capacitor c=0.00246068f \
 //x=41.695 //y=4.07 //x2=42.55 //y2=2.08
cc_3123 ( N_noxref_10_c_3678_n N_noxref_13_c_4445_n ) capacitor c=0.0742507f \
 //x=41.81 //y=2.08 //x2=42.55 //y2=2.08
cc_3124 ( N_noxref_10_c_3683_n N_noxref_13_c_4445_n ) capacitor c=0.00284029f \
 //x=41.615 //y=1.915 //x2=42.55 //y2=2.08
cc_3125 ( N_noxref_10_M102_noxref_g N_noxref_13_M104_noxref_g ) capacitor \
 c=0.0104611f //x=41.71 //y=6.02 //x2=42.59 //y2=6.02
cc_3126 ( N_noxref_10_M103_noxref_g N_noxref_13_M104_noxref_g ) capacitor \
 c=0.106811f //x=42.15 //y=6.02 //x2=42.59 //y2=6.02
cc_3127 ( N_noxref_10_M103_noxref_g N_noxref_13_M105_noxref_g ) capacitor \
 c=0.0100341f //x=42.15 //y=6.02 //x2=43.03 //y2=6.02
cc_3128 ( N_noxref_10_c_3679_n N_noxref_13_c_4523_n ) capacitor c=4.86506e-19 \
 //x=41.615 //y=0.865 //x2=42.585 //y2=0.905
cc_3129 ( N_noxref_10_c_3681_n N_noxref_13_c_4523_n ) capacitor c=0.00152104f \
 //x=41.615 //y=1.21 //x2=42.585 //y2=0.905
cc_3130 ( N_noxref_10_c_3686_n N_noxref_13_c_4523_n ) capacitor c=0.0151475f \
 //x=42.145 //y=0.865 //x2=42.585 //y2=0.905
cc_3131 ( N_noxref_10_c_3682_n N_noxref_13_c_4526_n ) capacitor c=0.00109982f \
 //x=41.615 //y=1.52 //x2=42.585 //y2=1.25
cc_3132 ( N_noxref_10_c_3688_n N_noxref_13_c_4526_n ) capacitor c=0.0111064f \
 //x=42.145 //y=1.21 //x2=42.585 //y2=1.25
cc_3133 ( N_noxref_10_c_3682_n N_noxref_13_c_4528_n ) capacitor c=9.57794e-19 \
 //x=41.615 //y=1.52 //x2=42.585 //y2=1.56
cc_3134 ( N_noxref_10_c_3683_n N_noxref_13_c_4528_n ) capacitor c=0.00662747f \
 //x=41.615 //y=1.915 //x2=42.585 //y2=1.56
cc_3135 ( N_noxref_10_c_3688_n N_noxref_13_c_4528_n ) capacitor c=0.00862358f \
 //x=42.145 //y=1.21 //x2=42.585 //y2=1.56
cc_3136 ( N_noxref_10_c_3686_n N_noxref_13_c_4531_n ) capacitor c=0.00124821f \
 //x=42.145 //y=0.865 //x2=43.115 //y2=0.905
cc_3137 ( N_noxref_10_c_3688_n N_noxref_13_c_4532_n ) capacitor c=0.00200715f \
 //x=42.145 //y=1.21 //x2=43.115 //y2=1.25
cc_3138 ( N_noxref_10_c_3678_n N_noxref_13_c_4533_n ) capacitor c=0.00282278f \
 //x=41.81 //y=2.08 //x2=42.55 //y2=2.08
cc_3139 ( N_noxref_10_c_3683_n N_noxref_13_c_4533_n ) capacitor c=0.0172771f \
 //x=41.615 //y=1.915 //x2=42.55 //y2=2.08
cc_3140 ( N_noxref_10_c_3678_n N_noxref_13_c_4535_n ) capacitor c=0.00344981f \
 //x=41.81 //y=2.08 //x2=42.58 //y2=4.7
cc_3141 ( N_noxref_10_c_3724_n N_noxref_13_c_4535_n ) capacitor c=0.0293367f \
 //x=41.81 //y=4.7 //x2=42.58 //y2=4.7
cc_3142 ( N_noxref_10_c_3690_n N_D_c_4909_n ) capacitor c=0.0249192f //x=31.7 \
 //y=4.07 //x2=49.835 //y2=2.96
cc_3143 ( N_noxref_10_c_3742_n N_D_c_4909_n ) capacitor c=6.36028e-19 \
 //x=26.385 //y=4.07 //x2=49.835 //y2=2.96
cc_3144 ( N_noxref_10_c_3675_n N_D_c_4909_n ) capacitor c=0.0192451f //x=26.27 \
 //y=2.08 //x2=49.835 //y2=2.96
cc_3145 ( N_noxref_10_c_3678_n N_D_c_4909_n ) capacitor c=0.0210088f //x=41.81 \
 //y=2.08 //x2=49.835 //y2=2.96
cc_3146 ( N_noxref_10_c_3754_n N_D_c_4909_n ) capacitor c=0.0187394f \
 //x=31.817 //y=3.905 //x2=49.835 //y2=2.96
cc_3147 ( N_noxref_10_c_3675_n N_D_c_5060_n ) capacitor c=0.00179385f \
 //x=26.27 //y=2.08 //x2=25.645 //y2=2.96
cc_3148 ( N_noxref_10_c_3742_n N_D_c_4916_n ) capacitor c=0.00735597f \
 //x=26.385 //y=4.07 //x2=25.53 //y2=2.08
cc_3149 ( N_noxref_10_c_3745_n N_D_c_4916_n ) capacitor c=0.00400249f \
 //x=26.27 //y=4.535 //x2=25.53 //y2=2.08
cc_3150 ( N_noxref_10_c_3675_n N_D_c_4916_n ) capacitor c=0.0756279f //x=26.27 \
 //y=2.08 //x2=25.53 //y2=2.08
cc_3151 ( N_noxref_10_c_3771_n N_D_c_4916_n ) capacitor c=0.00282278f \
 //x=26.27 //y=2.08 //x2=25.53 //y2=2.08
cc_3152 ( N_noxref_10_c_3774_n N_D_c_4916_n ) capacitor c=0.00344981f //x=26.3 \
 //y=4.7 //x2=25.53 //y2=2.08
cc_3153 ( N_noxref_10_M84_noxref_g N_D_M82_noxref_g ) capacitor c=0.0104611f \
 //x=26.31 //y=6.02 //x2=25.43 //y2=6.02
cc_3154 ( N_noxref_10_M84_noxref_g N_D_M83_noxref_g ) capacitor c=0.106811f \
 //x=26.31 //y=6.02 //x2=25.87 //y2=6.02
cc_3155 ( N_noxref_10_M85_noxref_g N_D_M83_noxref_g ) capacitor c=0.0100341f \
 //x=26.75 //y=6.02 //x2=25.87 //y2=6.02
cc_3156 ( N_noxref_10_c_3760_n N_D_c_4928_n ) capacitor c=4.86506e-19 \
 //x=26.305 //y=0.905 //x2=25.335 //y2=0.865
cc_3157 ( N_noxref_10_c_3760_n N_D_c_4930_n ) capacitor c=0.00152104f \
 //x=26.305 //y=0.905 //x2=25.335 //y2=1.21
cc_3158 ( N_noxref_10_c_3761_n N_D_c_4931_n ) capacitor c=0.00109982f \
 //x=26.305 //y=1.25 //x2=25.335 //y2=1.52
cc_3159 ( N_noxref_10_c_3762_n N_D_c_4931_n ) capacitor c=9.57794e-19 \
 //x=26.305 //y=1.56 //x2=25.335 //y2=1.52
cc_3160 ( N_noxref_10_c_3675_n N_D_c_4932_n ) capacitor c=0.00284029f \
 //x=26.27 //y=2.08 //x2=25.335 //y2=1.915
cc_3161 ( N_noxref_10_c_3762_n N_D_c_4932_n ) capacitor c=0.00662747f \
 //x=26.305 //y=1.56 //x2=25.335 //y2=1.915
cc_3162 ( N_noxref_10_c_3771_n N_D_c_4932_n ) capacitor c=0.0172771f //x=26.27 \
 //y=2.08 //x2=25.335 //y2=1.915
cc_3163 ( N_noxref_10_c_3760_n N_D_c_4935_n ) capacitor c=0.0151475f \
 //x=26.305 //y=0.905 //x2=25.865 //y2=0.865
cc_3164 ( N_noxref_10_c_3768_n N_D_c_4935_n ) capacitor c=0.00124821f \
 //x=26.835 //y=0.905 //x2=25.865 //y2=0.865
cc_3165 ( N_noxref_10_c_3761_n N_D_c_4937_n ) capacitor c=0.0111064f \
 //x=26.305 //y=1.25 //x2=25.865 //y2=1.21
cc_3166 ( N_noxref_10_c_3762_n N_D_c_4937_n ) capacitor c=0.00862358f \
 //x=26.305 //y=1.56 //x2=25.865 //y2=1.21
cc_3167 ( N_noxref_10_c_3769_n N_D_c_4937_n ) capacitor c=0.00200715f \
 //x=26.835 //y=1.25 //x2=25.865 //y2=1.21
cc_3168 ( N_noxref_10_c_3745_n N_D_c_4972_n ) capacitor c=0.00417994f \
 //x=26.27 //y=4.535 //x2=25.53 //y2=4.7
cc_3169 ( N_noxref_10_c_3774_n N_D_c_4972_n ) capacitor c=0.0293367f //x=26.3 \
 //y=4.7 //x2=25.53 //y2=4.7
cc_3170 ( N_noxref_10_c_3690_n N_CLK_c_5643_n ) capacitor c=0.302855f //x=31.7 \
 //y=4.07 //x2=29.855 //y2=4.44
cc_3171 ( N_noxref_10_c_3742_n N_CLK_c_5643_n ) capacitor c=0.028941f \
 //x=26.385 //y=4.07 //x2=29.855 //y2=4.44
cc_3172 ( N_noxref_10_c_3745_n N_CLK_c_5643_n ) capacitor c=0.0016972f \
 //x=26.27 //y=4.535 //x2=29.855 //y2=4.44
cc_3173 ( N_noxref_10_c_3675_n N_CLK_c_5643_n ) capacitor c=0.0207534f \
 //x=26.27 //y=2.08 //x2=29.855 //y2=4.44
cc_3174 ( N_noxref_10_c_3701_n N_CLK_c_5643_n ) capacitor c=0.0219114f \
 //x=29.365 //y=5.155 //x2=29.855 //y2=4.44
cc_3175 ( N_noxref_10_c_3763_n N_CLK_c_5643_n ) capacitor c=0.00960248f \
 //x=26.675 //y=4.79 //x2=29.855 //y2=4.44
cc_3176 ( N_noxref_10_c_3774_n N_CLK_c_5643_n ) capacitor c=0.00203982f \
 //x=26.3 //y=4.7 //x2=29.855 //y2=4.44
cc_3177 ( N_noxref_10_c_3690_n N_CLK_c_5668_n ) capacitor c=0.139602f //x=31.7 \
 //y=4.07 //x2=39.105 //y2=4.44
cc_3178 ( N_noxref_10_c_3691_n N_CLK_c_5668_n ) capacitor c=0.625476f \
 //x=41.695 //y=4.07 //x2=39.105 //y2=4.44
cc_3179 ( N_noxref_10_c_3694_n N_CLK_c_5668_n ) capacitor c=0.0265302f \
 //x=31.93 //y=4.07 //x2=39.105 //y2=4.44
cc_3180 ( N_noxref_10_c_3707_n N_CLK_c_5668_n ) capacitor c=0.0182691f \
 //x=31.735 //y=5.155 //x2=39.105 //y2=4.44
cc_3181 ( N_noxref_10_c_3801_p N_CLK_c_5668_n ) capacitor c=0.0207896f \
 //x=31.82 //y=5.07 //x2=39.105 //y2=4.44
cc_3182 ( N_noxref_10_c_3891_p N_CLK_c_5668_n ) capacitor c=0.0311227f \
 //x=30.16 //y=5.155 //x2=39.105 //y2=4.44
cc_3183 ( N_noxref_10_c_3714_n N_CLK_c_5668_n ) capacitor c=0.00215288f \
 //x=31.815 //y=4.07 //x2=39.105 //y2=4.44
cc_3184 ( N_noxref_10_c_3690_n N_CLK_c_5679_n ) capacitor c=0.026534f //x=31.7 \
 //y=4.07 //x2=30.085 //y2=4.44
cc_3185 ( N_noxref_10_c_3697_n N_CLK_c_5679_n ) capacitor c=0.00241768f \
 //x=30.075 //y=5.155 //x2=30.085 //y2=4.44
cc_3186 ( N_noxref_10_c_3691_n N_CLK_c_5680_n ) capacitor c=0.236351f \
 //x=41.695 //y=4.07 //x2=54.275 //y2=4.44
cc_3187 ( N_noxref_10_c_3678_n N_CLK_c_5680_n ) capacitor c=0.021665f \
 //x=41.81 //y=2.08 //x2=54.275 //y2=4.44
cc_3188 ( N_noxref_10_c_3724_n N_CLK_c_5680_n ) capacitor c=0.0107036f \
 //x=41.81 //y=4.7 //x2=54.275 //y2=4.44
cc_3189 ( N_noxref_10_c_3691_n N_CLK_c_5704_n ) capacitor c=0.0267161f \
 //x=41.695 //y=4.07 //x2=39.335 //y2=4.44
cc_3190 ( N_noxref_10_c_3690_n N_CLK_c_5625_n ) capacitor c=0.0231929f \
 //x=31.7 //y=4.07 //x2=29.97 //y2=2.08
cc_3191 ( N_noxref_10_c_3697_n N_CLK_c_5625_n ) capacitor c=0.014564f \
 //x=30.075 //y=5.155 //x2=29.97 //y2=2.08
cc_3192 ( N_noxref_10_c_3801_p N_CLK_c_5625_n ) capacitor c=7.17254e-19 \
 //x=31.82 //y=5.07 //x2=29.97 //y2=2.08
cc_3193 ( N_noxref_10_c_3754_n N_CLK_c_5625_n ) capacitor c=0.00157145f \
 //x=31.817 //y=3.905 //x2=29.97 //y2=2.08
cc_3194 ( N_noxref_10_c_3691_n N_CLK_c_5626_n ) capacitor c=0.0187718f \
 //x=41.695 //y=4.07 //x2=39.22 //y2=2.08
cc_3195 ( N_noxref_10_c_3678_n N_CLK_c_5626_n ) capacitor c=6.57265e-19 \
 //x=41.81 //y=2.08 //x2=39.22 //y2=2.08
cc_3196 ( N_noxref_10_c_3697_n N_CLK_M88_noxref_g ) capacitor c=0.016514f \
 //x=30.075 //y=5.155 //x2=29.94 //y2=6.02
cc_3197 ( N_noxref_10_M88_noxref_d N_CLK_M88_noxref_g ) capacitor c=0.0180032f \
 //x=30.015 //y=5.02 //x2=29.94 //y2=6.02
cc_3198 ( N_noxref_10_c_3703_n N_CLK_M89_noxref_g ) capacitor c=0.01736f \
 //x=30.955 //y=5.155 //x2=30.38 //y2=6.02
cc_3199 ( N_noxref_10_M88_noxref_d N_CLK_M89_noxref_g ) capacitor c=0.0180032f \
 //x=30.015 //y=5.02 //x2=30.38 //y2=6.02
cc_3200 ( N_noxref_10_c_3891_p N_CLK_c_6000_n ) capacitor c=0.00426767f \
 //x=30.16 //y=5.155 //x2=30.305 //y2=4.79
cc_3201 ( N_noxref_10_c_3697_n N_CLK_c_5936_n ) capacitor c=0.00322046f \
 //x=30.075 //y=5.155 //x2=29.97 //y2=4.7
cc_3202 ( N_noxref_10_c_3675_n N_SN_c_6844_n ) capacitor c=0.0201924f \
 //x=26.27 //y=2.08 //x2=34.665 //y2=2.22
cc_3203 ( N_noxref_10_c_3912_p N_SN_c_6844_n ) capacitor c=0.0163057f \
 //x=31.42 //y=1.665 //x2=34.665 //y2=2.22
cc_3204 ( N_noxref_10_c_3754_n N_SN_c_6844_n ) capacitor c=0.0197307f \
 //x=31.817 //y=3.905 //x2=34.665 //y2=2.22
cc_3205 ( N_noxref_10_c_3766_n N_SN_c_6844_n ) capacitor c=3.11115e-19 \
 //x=26.68 //y=1.405 //x2=34.665 //y2=2.22
cc_3206 ( N_noxref_10_c_3771_n N_SN_c_6844_n ) capacitor c=0.00570799f \
 //x=26.27 //y=2.08 //x2=34.665 //y2=2.22
cc_3207 ( N_noxref_10_c_3678_n N_SN_c_6855_n ) capacitor c=0.0208418f \
 //x=41.81 //y=2.08 //x2=46.135 //y2=2.22
cc_3208 ( N_noxref_10_c_3683_n N_SN_c_6855_n ) capacitor c=0.00894156f \
 //x=41.615 //y=1.915 //x2=46.135 //y2=2.22
cc_3209 ( N_noxref_10_c_3691_n N_SN_c_6890_n ) capacitor c=0.0190126f \
 //x=41.695 //y=4.07 //x2=34.78 //y2=2.08
cc_3210 ( N_noxref_10_c_3754_n N_SN_c_6890_n ) capacitor c=3.18993e-19 \
 //x=31.817 //y=3.905 //x2=34.78 //y2=2.08
cc_3211 ( N_noxref_10_c_3690_n N_noxref_24_c_8424_n ) capacitor c=0.202797f \
 //x=31.7 //y=4.07 //x2=79.065 //y2=3.33
cc_3212 ( N_noxref_10_c_3742_n N_noxref_24_c_8424_n ) capacitor c=0.0136135f \
 //x=26.385 //y=4.07 //x2=79.065 //y2=3.33
cc_3213 ( N_noxref_10_c_3691_n N_noxref_24_c_8424_n ) capacitor c=0.0684106f \
 //x=41.695 //y=4.07 //x2=79.065 //y2=3.33
cc_3214 ( N_noxref_10_c_3694_n N_noxref_24_c_8424_n ) capacitor c=4.80497e-19 \
 //x=31.93 //y=4.07 //x2=79.065 //y2=3.33
cc_3215 ( N_noxref_10_c_3675_n N_noxref_24_c_8424_n ) capacitor c=0.019633f \
 //x=26.27 //y=2.08 //x2=79.065 //y2=3.33
cc_3216 ( N_noxref_10_c_3678_n N_noxref_24_c_8424_n ) capacitor c=0.0187404f \
 //x=41.81 //y=2.08 //x2=79.065 //y2=3.33
cc_3217 ( N_noxref_10_c_3754_n N_noxref_24_c_8424_n ) capacitor c=0.0187428f \
 //x=31.817 //y=3.905 //x2=79.065 //y2=3.33
cc_3218 ( N_noxref_10_c_3675_n N_noxref_24_c_8465_n ) capacitor c=0.00116483f \
 //x=26.27 //y=2.08 //x2=23.68 //y2=3.33
cc_3219 ( N_noxref_10_c_3762_n N_noxref_36_c_9699_n ) capacitor c=0.00623646f \
 //x=26.305 //y=1.56 //x2=26.085 //y2=1.495
cc_3220 ( N_noxref_10_c_3771_n N_noxref_36_c_9699_n ) capacitor c=0.00173579f \
 //x=26.27 //y=2.08 //x2=26.085 //y2=1.495
cc_3221 ( N_noxref_10_c_3675_n N_noxref_36_c_9700_n ) capacitor c=0.00156605f \
 //x=26.27 //y=2.08 //x2=26.97 //y2=0.53
cc_3222 ( N_noxref_10_c_3760_n N_noxref_36_c_9700_n ) capacitor c=0.0188655f \
 //x=26.305 //y=0.905 //x2=26.97 //y2=0.53
cc_3223 ( N_noxref_10_c_3768_n N_noxref_36_c_9700_n ) capacitor c=0.00656458f \
 //x=26.835 //y=0.905 //x2=26.97 //y2=0.53
cc_3224 ( N_noxref_10_c_3771_n N_noxref_36_c_9700_n ) capacitor c=2.1838e-19 \
 //x=26.27 //y=2.08 //x2=26.97 //y2=0.53
cc_3225 ( N_noxref_10_c_3760_n N_noxref_36_M15_noxref_s ) capacitor \
 c=0.00623646f //x=26.305 //y=0.905 //x2=24.98 //y2=0.365
cc_3226 ( N_noxref_10_c_3768_n N_noxref_36_M15_noxref_s ) capacitor \
 c=0.0143002f //x=26.835 //y=0.905 //x2=24.98 //y2=0.365
cc_3227 ( N_noxref_10_c_3769_n N_noxref_36_M15_noxref_s ) capacitor \
 c=0.00290153f //x=26.835 //y=1.25 //x2=24.98 //y2=0.365
cc_3228 ( N_noxref_10_M19_noxref_d N_noxref_37_M17_noxref_s ) capacitor \
 c=0.00309936f //x=31.145 //y=0.915 //x2=28.205 //y2=0.375
cc_3229 ( N_noxref_10_c_3677_n N_noxref_38_c_9797_n ) capacitor c=0.00457167f \
 //x=31.735 //y=1.665 //x2=31.735 //y2=0.54
cc_3230 ( N_noxref_10_M19_noxref_d N_noxref_38_c_9797_n ) capacitor \
 c=0.0115903f //x=31.145 //y=0.915 //x2=31.735 //y2=0.54
cc_3231 ( N_noxref_10_c_3912_p N_noxref_38_c_9807_n ) capacitor c=0.0200405f \
 //x=31.42 //y=1.665 //x2=30.85 //y2=0.995
cc_3232 ( N_noxref_10_M19_noxref_d N_noxref_38_M18_noxref_d ) capacitor \
 c=5.27807e-19 //x=31.145 //y=0.915 //x2=29.61 //y2=0.91
cc_3233 ( N_noxref_10_c_3677_n N_noxref_38_M19_noxref_s ) capacitor \
 c=0.0196084f //x=31.735 //y=1.665 //x2=30.715 //y2=0.375
cc_3234 ( N_noxref_10_M19_noxref_d N_noxref_38_M19_noxref_s ) capacitor \
 c=0.0426368f //x=31.145 //y=0.915 //x2=30.715 //y2=0.375
cc_3235 ( N_noxref_10_c_3677_n N_noxref_39_c_9859_n ) capacitor c=3.83325e-19 \
 //x=31.735 //y=1.665 //x2=33.15 //y2=1.505
cc_3236 ( N_noxref_10_M19_noxref_d N_noxref_39_M20_noxref_s ) capacitor \
 c=2.55333e-19 //x=31.145 //y=0.915 //x2=33.015 //y2=0.375
cc_3237 ( N_noxref_10_c_3683_n N_noxref_42_c_10017_n ) capacitor c=0.0034165f \
 //x=41.615 //y=1.915 //x2=41.395 //y2=1.495
cc_3238 ( N_noxref_10_c_3678_n N_noxref_42_c_9999_n ) capacitor c=0.011618f \
 //x=41.81 //y=2.08 //x2=42.28 //y2=1.58
cc_3239 ( N_noxref_10_c_3682_n N_noxref_42_c_9999_n ) capacitor c=0.00696403f \
 //x=41.615 //y=1.52 //x2=42.28 //y2=1.58
cc_3240 ( N_noxref_10_c_3683_n N_noxref_42_c_9999_n ) capacitor c=0.0174694f \
 //x=41.615 //y=1.915 //x2=42.28 //y2=1.58
cc_3241 ( N_noxref_10_c_3685_n N_noxref_42_c_9999_n ) capacitor c=0.00776811f \
 //x=41.99 //y=1.365 //x2=42.28 //y2=1.58
cc_3242 ( N_noxref_10_c_3688_n N_noxref_42_c_9999_n ) capacitor c=0.00339872f \
 //x=42.145 //y=1.21 //x2=42.28 //y2=1.58
cc_3243 ( N_noxref_10_c_3683_n N_noxref_42_c_10006_n ) capacitor c=6.71402e-19 \
 //x=41.615 //y=1.915 //x2=42.365 //y2=1.495
cc_3244 ( N_noxref_10_c_3679_n N_noxref_42_M25_noxref_s ) capacitor \
 c=0.0326577f //x=41.615 //y=0.865 //x2=41.26 //y2=0.365
cc_3245 ( N_noxref_10_c_3682_n N_noxref_42_M25_noxref_s ) capacitor \
 c=3.48408e-19 //x=41.615 //y=1.52 //x2=41.26 //y2=0.365
cc_3246 ( N_noxref_10_c_3686_n N_noxref_42_M25_noxref_s ) capacitor \
 c=0.0120759f //x=42.145 //y=0.865 //x2=41.26 //y2=0.365
cc_3247 ( N_noxref_11_c_3959_n N_noxref_12_c_4204_n ) capacitor c=0.0187688f \
 //x=43.29 //y=2.59 //x2=47.245 //y2=3.7
cc_3248 ( N_noxref_11_c_3961_n N_noxref_12_c_4204_n ) capacitor c=0.0197889f \
 //x=45.14 //y=2.08 //x2=47.245 //y2=3.7
cc_3249 ( N_noxref_11_c_3959_n N_noxref_12_c_4114_n ) capacitor c=3.49822e-19 \
 //x=43.29 //y=2.59 //x2=39.96 //y2=3.7
cc_3250 ( N_noxref_11_c_3961_n N_noxref_12_c_4115_n ) capacitor c=0.00107283f \
 //x=45.14 //y=2.08 //x2=47.36 //y2=2.08
cc_3251 ( N_noxref_11_c_3959_n N_noxref_13_c_4455_n ) capacitor c=0.0181936f \
 //x=43.29 //y=2.59 //x2=47.985 //y2=4.07
cc_3252 ( N_noxref_11_c_3961_n N_noxref_13_c_4455_n ) capacitor c=0.0194977f \
 //x=45.14 //y=2.08 //x2=47.985 //y2=4.07
cc_3253 ( N_noxref_11_c_3959_n N_noxref_13_c_4513_n ) capacitor c=0.00131333f \
 //x=43.29 //y=2.59 //x2=42.665 //y2=4.07
cc_3254 ( N_noxref_11_c_3956_n N_noxref_13_c_4434_n ) capacitor c=0.00564994f \
 //x=45.025 //y=2.59 //x2=48.215 //y2=2.59
cc_3255 ( N_noxref_11_c_3975_n N_noxref_13_c_4515_n ) capacitor c=0.0127164f \
 //x=42.725 //y=5.2 //x2=42.55 //y2=4.535
cc_3256 ( N_noxref_11_c_3959_n N_noxref_13_c_4515_n ) capacitor c=0.0101115f \
 //x=43.29 //y=2.59 //x2=42.55 //y2=4.535
cc_3257 ( N_noxref_11_c_3957_n N_noxref_13_c_4445_n ) capacitor c=0.00720056f \
 //x=43.405 //y=2.59 //x2=42.55 //y2=2.08
cc_3258 ( N_noxref_11_c_3959_n N_noxref_13_c_4445_n ) capacitor c=0.0664516f \
 //x=43.29 //y=2.59 //x2=42.55 //y2=2.08
cc_3259 ( N_noxref_11_c_3961_n N_noxref_13_c_4445_n ) capacitor c=5.34685e-19 \
 //x=45.14 //y=2.08 //x2=42.55 //y2=2.08
cc_3260 ( N_noxref_11_M107_noxref_g N_noxref_13_c_4464_n ) capacitor \
 c=0.0168349f //x=45.78 //y=6.02 //x2=46.355 //y2=5.155
cc_3261 ( N_noxref_11_c_3959_n N_noxref_13_c_4468_n ) capacitor c=2.97874e-19 \
 //x=43.29 //y=2.59 //x2=45.645 //y2=5.155
cc_3262 ( N_noxref_11_M106_noxref_g N_noxref_13_c_4468_n ) capacitor \
 c=0.0213876f //x=45.34 //y=6.02 //x2=45.645 //y2=5.155
cc_3263 ( N_noxref_11_c_4028_p N_noxref_13_c_4468_n ) capacitor c=0.00428486f \
 //x=45.705 //y=4.79 //x2=45.645 //y2=5.155
cc_3264 ( N_noxref_11_c_3975_n N_noxref_13_M104_noxref_g ) capacitor \
 c=0.0166421f //x=42.725 //y=5.2 //x2=42.59 //y2=6.02
cc_3265 ( N_noxref_11_M104_noxref_d N_noxref_13_M104_noxref_g ) capacitor \
 c=0.0173476f //x=42.665 //y=5.02 //x2=42.59 //y2=6.02
cc_3266 ( N_noxref_11_c_3981_n N_noxref_13_M105_noxref_g ) capacitor \
 c=0.018922f //x=43.205 //y=5.2 //x2=43.03 //y2=6.02
cc_3267 ( N_noxref_11_M104_noxref_d N_noxref_13_M105_noxref_g ) capacitor \
 c=0.0179769f //x=42.665 //y=5.02 //x2=43.03 //y2=6.02
cc_3268 ( N_noxref_11_M26_noxref_d N_noxref_13_c_4523_n ) capacitor \
 c=0.00217566f //x=42.66 //y=0.905 //x2=42.585 //y2=0.905
cc_3269 ( N_noxref_11_M26_noxref_d N_noxref_13_c_4526_n ) capacitor \
 c=0.0034598f //x=42.66 //y=0.905 //x2=42.585 //y2=1.25
cc_3270 ( N_noxref_11_M26_noxref_d N_noxref_13_c_4528_n ) capacitor \
 c=0.00669531f //x=42.66 //y=0.905 //x2=42.585 //y2=1.56
cc_3271 ( N_noxref_11_c_3959_n N_noxref_13_c_4557_n ) capacitor c=0.0142673f \
 //x=43.29 //y=2.59 //x2=42.955 //y2=4.79
cc_3272 ( N_noxref_11_c_4037_p N_noxref_13_c_4557_n ) capacitor c=0.00407665f \
 //x=42.81 //y=5.2 //x2=42.955 //y2=4.79
cc_3273 ( N_noxref_11_M26_noxref_d N_noxref_13_c_4559_n ) capacitor \
 c=0.00241102f //x=42.66 //y=0.905 //x2=42.96 //y2=0.75
cc_3274 ( N_noxref_11_c_3958_n N_noxref_13_c_4560_n ) capacitor c=0.00371277f \
 //x=43.205 //y=1.655 //x2=42.96 //y2=1.405
cc_3275 ( N_noxref_11_M26_noxref_d N_noxref_13_c_4560_n ) capacitor \
 c=0.0137169f //x=42.66 //y=0.905 //x2=42.96 //y2=1.405
cc_3276 ( N_noxref_11_M26_noxref_d N_noxref_13_c_4531_n ) capacitor \
 c=0.00132245f //x=42.66 //y=0.905 //x2=43.115 //y2=0.905
cc_3277 ( N_noxref_11_c_3958_n N_noxref_13_c_4532_n ) capacitor c=0.00457401f \
 //x=43.205 //y=1.655 //x2=43.115 //y2=1.25
cc_3278 ( N_noxref_11_M26_noxref_d N_noxref_13_c_4532_n ) capacitor \
 c=0.00566463f //x=42.66 //y=0.905 //x2=43.115 //y2=1.25
cc_3279 ( N_noxref_11_c_3959_n N_noxref_13_c_4533_n ) capacitor c=0.00709342f \
 //x=43.29 //y=2.59 //x2=42.55 //y2=2.08
cc_3280 ( N_noxref_11_c_3959_n N_noxref_13_c_4566_n ) capacitor c=0.00306024f \
 //x=43.29 //y=2.59 //x2=42.55 //y2=1.915
cc_3281 ( N_noxref_11_M26_noxref_d N_noxref_13_c_4566_n ) capacitor \
 c=0.00660593f //x=42.66 //y=0.905 //x2=42.55 //y2=1.915
cc_3282 ( N_noxref_11_c_3975_n N_noxref_13_c_4535_n ) capacitor c=0.00346527f \
 //x=42.725 //y=5.2 //x2=42.58 //y2=4.7
cc_3283 ( N_noxref_11_c_3959_n N_noxref_13_c_4535_n ) capacitor c=0.00533692f \
 //x=43.29 //y=2.59 //x2=42.58 //y2=4.7
cc_3284 ( N_noxref_11_M107_noxref_g N_noxref_13_M106_noxref_d ) capacitor \
 c=0.0180032f //x=45.78 //y=6.02 //x2=45.415 //y2=5.02
cc_3285 ( N_noxref_11_c_3956_n N_D_c_4909_n ) capacitor c=0.172771f //x=45.025 \
 //y=2.59 //x2=49.835 //y2=2.96
cc_3286 ( N_noxref_11_c_3957_n N_D_c_4909_n ) capacitor c=0.0293646f \
 //x=43.405 //y=2.59 //x2=49.835 //y2=2.96
cc_3287 ( N_noxref_11_c_3959_n N_D_c_4909_n ) capacitor c=0.0206018f //x=43.29 \
 //y=2.59 //x2=49.835 //y2=2.96
cc_3288 ( N_noxref_11_c_3961_n N_D_c_4909_n ) capacitor c=0.0216195f //x=45.14 \
 //y=2.08 //x2=49.835 //y2=2.96
cc_3289 ( N_noxref_11_c_3975_n N_CLK_c_5680_n ) capacitor c=0.0185297f \
 //x=42.725 //y=5.2 //x2=54.275 //y2=4.44
cc_3290 ( N_noxref_11_c_3979_n N_CLK_c_5680_n ) capacitor c=0.018142f \
 //x=42.015 //y=5.2 //x2=54.275 //y2=4.44
cc_3291 ( N_noxref_11_c_3959_n N_CLK_c_5680_n ) capacitor c=0.0208321f \
 //x=43.29 //y=2.59 //x2=54.275 //y2=4.44
cc_3292 ( N_noxref_11_c_3961_n N_CLK_c_5680_n ) capacitor c=0.0208709f \
 //x=45.14 //y=2.08 //x2=54.275 //y2=4.44
cc_3293 ( N_noxref_11_c_3993_n N_CLK_c_5680_n ) capacitor c=0.0166984f \
 //x=45.415 //y=4.79 //x2=54.275 //y2=4.44
cc_3294 ( N_noxref_11_c_3956_n N_SN_c_6855_n ) capacitor c=0.172576f \
 //x=45.025 //y=2.59 //x2=46.135 //y2=2.22
cc_3295 ( N_noxref_11_c_3957_n N_SN_c_6855_n ) capacitor c=0.0290445f \
 //x=43.405 //y=2.59 //x2=46.135 //y2=2.22
cc_3296 ( N_noxref_11_c_4061_p N_SN_c_6855_n ) capacitor c=0.0146822f \
 //x=42.935 //y=1.655 //x2=46.135 //y2=2.22
cc_3297 ( N_noxref_11_c_3959_n N_SN_c_6855_n ) capacitor c=0.0217395f \
 //x=43.29 //y=2.59 //x2=46.135 //y2=2.22
cc_3298 ( N_noxref_11_c_3961_n N_SN_c_6855_n ) capacitor c=0.021104f //x=45.14 \
 //y=2.08 //x2=46.135 //y2=2.22
cc_3299 ( N_noxref_11_c_3966_n N_SN_c_6855_n ) capacitor c=0.011987f //x=44.84 \
 //y=1.915 //x2=46.135 //y2=2.22
cc_3300 ( N_noxref_11_c_3961_n N_SN_c_6876_n ) capacitor c=0.00165648f \
 //x=45.14 //y=2.08 //x2=46.365 //y2=2.22
cc_3301 ( N_noxref_11_c_3966_n N_SN_c_6876_n ) capacitor c=2.3323e-19 \
 //x=44.84 //y=1.915 //x2=46.365 //y2=2.22
cc_3302 ( N_noxref_11_c_3956_n N_SN_c_6891_n ) capacitor c=0.00320677f \
 //x=45.025 //y=2.59 //x2=46.25 //y2=2.08
cc_3303 ( N_noxref_11_c_3959_n N_SN_c_6891_n ) capacitor c=2.96936e-19 \
 //x=43.29 //y=2.59 //x2=46.25 //y2=2.08
cc_3304 ( N_noxref_11_c_3961_n N_SN_c_6891_n ) capacitor c=0.0428203f \
 //x=45.14 //y=2.08 //x2=46.25 //y2=2.08
cc_3305 ( N_noxref_11_c_3966_n N_SN_c_6891_n ) capacitor c=0.00208635f \
 //x=44.84 //y=1.915 //x2=46.25 //y2=2.08
cc_3306 ( N_noxref_11_c_4028_p N_SN_c_6891_n ) capacitor c=0.00147352f \
 //x=45.705 //y=4.79 //x2=46.25 //y2=2.08
cc_3307 ( N_noxref_11_c_3993_n N_SN_c_6891_n ) capacitor c=0.00142741f \
 //x=45.415 //y=4.79 //x2=46.25 //y2=2.08
cc_3308 ( N_noxref_11_M106_noxref_g N_SN_M108_noxref_g ) capacitor \
 c=0.0105869f //x=45.34 //y=6.02 //x2=46.22 //y2=6.02
cc_3309 ( N_noxref_11_M107_noxref_g N_SN_M108_noxref_g ) capacitor c=0.10632f \
 //x=45.78 //y=6.02 //x2=46.22 //y2=6.02
cc_3310 ( N_noxref_11_M107_noxref_g N_SN_M109_noxref_g ) capacitor \
 c=0.0101598f //x=45.78 //y=6.02 //x2=46.66 //y2=6.02
cc_3311 ( N_noxref_11_c_3962_n N_SN_c_7123_n ) capacitor c=5.72482e-19 \
 //x=44.84 //y=0.875 //x2=45.815 //y2=0.91
cc_3312 ( N_noxref_11_c_3964_n N_SN_c_7123_n ) capacitor c=0.00149976f \
 //x=44.84 //y=1.22 //x2=45.815 //y2=0.91
cc_3313 ( N_noxref_11_c_3969_n N_SN_c_7123_n ) capacitor c=0.0160123f \
 //x=45.37 //y=0.875 //x2=45.815 //y2=0.91
cc_3314 ( N_noxref_11_c_3965_n N_SN_c_7126_n ) capacitor c=0.00111227f \
 //x=44.84 //y=1.53 //x2=45.815 //y2=1.22
cc_3315 ( N_noxref_11_c_3971_n N_SN_c_7126_n ) capacitor c=0.0124075f \
 //x=45.37 //y=1.22 //x2=45.815 //y2=1.22
cc_3316 ( N_noxref_11_c_3969_n N_SN_c_7128_n ) capacitor c=0.00103227f \
 //x=45.37 //y=0.875 //x2=46.34 //y2=0.91
cc_3317 ( N_noxref_11_c_3971_n N_SN_c_7129_n ) capacitor c=0.0010154f \
 //x=45.37 //y=1.22 //x2=46.34 //y2=1.22
cc_3318 ( N_noxref_11_c_3971_n N_SN_c_7130_n ) capacitor c=9.23422e-19 \
 //x=45.37 //y=1.22 //x2=46.34 //y2=1.45
cc_3319 ( N_noxref_11_c_3961_n N_SN_c_7131_n ) capacitor c=0.00203769f \
 //x=45.14 //y=2.08 //x2=46.34 //y2=1.915
cc_3320 ( N_noxref_11_c_3966_n N_SN_c_7131_n ) capacitor c=0.00834532f \
 //x=44.84 //y=1.915 //x2=46.34 //y2=1.915
cc_3321 ( N_noxref_11_c_3961_n N_SN_c_7133_n ) capacitor c=0.00183762f \
 //x=45.14 //y=2.08 //x2=46.25 //y2=4.7
cc_3322 ( N_noxref_11_c_4028_p N_SN_c_7133_n ) capacitor c=0.0168581f \
 //x=45.705 //y=4.79 //x2=46.25 //y2=4.7
cc_3323 ( N_noxref_11_c_3993_n N_SN_c_7133_n ) capacitor c=0.00484466f \
 //x=45.415 //y=4.79 //x2=46.25 //y2=4.7
cc_3324 ( N_noxref_11_c_3956_n N_noxref_24_c_8424_n ) capacitor c=0.0119017f \
 //x=45.025 //y=2.59 //x2=79.065 //y2=3.33
cc_3325 ( N_noxref_11_c_3957_n N_noxref_24_c_8424_n ) capacitor c=8.86511e-19 \
 //x=43.405 //y=2.59 //x2=79.065 //y2=3.33
cc_3326 ( N_noxref_11_c_3959_n N_noxref_24_c_8424_n ) capacitor c=0.0187691f \
 //x=43.29 //y=2.59 //x2=79.065 //y2=3.33
cc_3327 ( N_noxref_11_c_3961_n N_noxref_24_c_8424_n ) capacitor c=0.0198064f \
 //x=45.14 //y=2.08 //x2=79.065 //y2=3.33
cc_3328 ( N_noxref_11_c_4061_p N_noxref_42_c_10017_n ) capacitor c=3.15806e-19 \
 //x=42.935 //y=1.655 //x2=41.395 //y2=1.495
cc_3329 ( N_noxref_11_c_4061_p N_noxref_42_c_10006_n ) capacitor c=0.0203424f \
 //x=42.935 //y=1.655 //x2=42.365 //y2=1.495
cc_3330 ( N_noxref_11_c_3958_n N_noxref_42_c_10007_n ) capacitor c=0.00457164f \
 //x=43.205 //y=1.655 //x2=43.25 //y2=0.53
cc_3331 ( N_noxref_11_M26_noxref_d N_noxref_42_c_10007_n ) capacitor \
 c=0.0115831f //x=42.66 //y=0.905 //x2=43.25 //y2=0.53
cc_3332 ( N_noxref_11_c_3958_n N_noxref_42_M25_noxref_s ) capacitor \
 c=0.0126484f //x=43.205 //y=1.655 //x2=41.26 //y2=0.365
cc_3333 ( N_noxref_11_M26_noxref_d N_noxref_42_M25_noxref_s ) capacitor \
 c=0.043966f //x=42.66 //y=0.905 //x2=41.26 //y2=0.365
cc_3334 ( N_noxref_11_c_3958_n N_noxref_43_c_10065_n ) capacitor c=4.08644e-19 \
 //x=43.205 //y=1.655 //x2=44.62 //y2=1.505
cc_3335 ( N_noxref_11_c_3966_n N_noxref_43_c_10065_n ) capacitor c=0.0034165f \
 //x=44.84 //y=1.915 //x2=44.62 //y2=1.505
cc_3336 ( N_noxref_11_c_3961_n N_noxref_43_c_10050_n ) capacitor c=0.0115578f \
 //x=45.14 //y=2.08 //x2=45.505 //y2=1.59
cc_3337 ( N_noxref_11_c_3965_n N_noxref_43_c_10050_n ) capacitor c=0.00697148f \
 //x=44.84 //y=1.53 //x2=45.505 //y2=1.59
cc_3338 ( N_noxref_11_c_3966_n N_noxref_43_c_10050_n ) capacitor c=0.0204849f \
 //x=44.84 //y=1.915 //x2=45.505 //y2=1.59
cc_3339 ( N_noxref_11_c_3968_n N_noxref_43_c_10050_n ) capacitor c=0.00610316f \
 //x=45.215 //y=1.375 //x2=45.505 //y2=1.59
cc_3340 ( N_noxref_11_c_3971_n N_noxref_43_c_10050_n ) capacitor c=0.00698822f \
 //x=45.37 //y=1.22 //x2=45.505 //y2=1.59
cc_3341 ( N_noxref_11_c_3962_n N_noxref_43_M27_noxref_s ) capacitor \
 c=0.0327271f //x=44.84 //y=0.875 //x2=44.485 //y2=0.375
cc_3342 ( N_noxref_11_c_3965_n N_noxref_43_M27_noxref_s ) capacitor \
 c=7.99997e-19 //x=44.84 //y=1.53 //x2=44.485 //y2=0.375
cc_3343 ( N_noxref_11_c_3966_n N_noxref_43_M27_noxref_s ) capacitor \
 c=0.00122123f //x=44.84 //y=1.915 //x2=44.485 //y2=0.375
cc_3344 ( N_noxref_11_c_3969_n N_noxref_43_M27_noxref_s ) capacitor \
 c=0.0121427f //x=45.37 //y=0.875 //x2=44.485 //y2=0.375
cc_3345 ( N_noxref_11_M26_noxref_d N_noxref_43_M27_noxref_s ) capacitor \
 c=2.53688e-19 //x=42.66 //y=0.905 //x2=44.485 //y2=0.375
cc_3346 ( N_noxref_12_c_4204_n N_noxref_13_c_4455_n ) capacitor c=0.433231f \
 //x=47.245 //y=3.7 //x2=47.985 //y2=4.07
cc_3347 ( N_noxref_12_c_4115_n N_noxref_13_c_4455_n ) capacitor c=0.0211201f \
 //x=47.36 //y=2.08 //x2=47.985 //y2=4.07
cc_3348 ( N_noxref_12_c_4204_n N_noxref_13_c_4513_n ) capacitor c=0.0294057f \
 //x=47.245 //y=3.7 //x2=42.665 //y2=4.07
cc_3349 ( N_noxref_12_c_4115_n N_noxref_13_c_4434_n ) capacitor c=0.00445416f \
 //x=47.36 //y=2.08 //x2=48.215 //y2=2.59
cc_3350 ( N_noxref_12_c_4204_n N_noxref_13_c_4445_n ) capacitor c=0.0187965f \
 //x=47.245 //y=3.7 //x2=42.55 //y2=2.08
cc_3351 ( N_noxref_12_c_4114_n N_noxref_13_c_4445_n ) capacitor c=5.98835e-19 \
 //x=39.96 //y=3.7 //x2=42.55 //y2=2.08
cc_3352 ( N_noxref_12_M110_noxref_g N_noxref_13_c_4470_n ) capacitor \
 c=0.01736f //x=47.1 //y=6.02 //x2=47.235 //y2=5.155
cc_3353 ( N_noxref_12_M111_noxref_g N_noxref_13_c_4474_n ) capacitor \
 c=0.0194981f //x=47.54 //y=6.02 //x2=48.015 //y2=5.155
cc_3354 ( N_noxref_12_c_4248_p N_noxref_13_c_4474_n ) capacitor c=0.00201851f \
 //x=47.36 //y=4.7 //x2=48.015 //y2=5.155
cc_3355 ( N_noxref_12_c_4249_p N_noxref_13_c_4447_n ) capacitor c=0.00371277f \
 //x=47.725 //y=1.415 //x2=48.015 //y2=1.665
cc_3356 ( N_noxref_12_c_4250_p N_noxref_13_c_4447_n ) capacitor c=0.00457401f \
 //x=47.88 //y=1.26 //x2=48.015 //y2=1.665
cc_3357 ( N_noxref_12_c_4204_n N_noxref_13_c_4448_n ) capacitor c=0.00735597f \
 //x=47.245 //y=3.7 //x2=48.1 //y2=2.59
cc_3358 ( N_noxref_12_c_4115_n N_noxref_13_c_4448_n ) capacitor c=0.0771184f \
 //x=47.36 //y=2.08 //x2=48.1 //y2=2.59
cc_3359 ( N_noxref_12_c_4253_p N_noxref_13_c_4448_n ) capacitor c=0.00709342f \
 //x=47.36 //y=2.08 //x2=48.1 //y2=2.59
cc_3360 ( N_noxref_12_c_4254_p N_noxref_13_c_4448_n ) capacitor c=0.00283672f \
 //x=47.36 //y=1.915 //x2=48.1 //y2=2.59
cc_3361 ( N_noxref_12_c_4248_p N_noxref_13_c_4448_n ) capacitor c=0.013844f \
 //x=47.36 //y=4.7 //x2=48.1 //y2=2.59
cc_3362 ( N_noxref_12_c_4115_n N_noxref_13_c_4587_n ) capacitor c=0.016476f \
 //x=47.36 //y=2.08 //x2=47.32 //y2=5.155
cc_3363 ( N_noxref_12_c_4248_p N_noxref_13_c_4587_n ) capacitor c=0.00475601f \
 //x=47.36 //y=4.7 //x2=47.32 //y2=5.155
cc_3364 ( N_noxref_12_c_4258_p N_noxref_13_M29_noxref_d ) capacitor \
 c=0.00217566f //x=47.35 //y=0.915 //x2=47.425 //y2=0.915
cc_3365 ( N_noxref_12_c_4259_p N_noxref_13_M29_noxref_d ) capacitor \
 c=0.0034598f //x=47.35 //y=1.26 //x2=47.425 //y2=0.915
cc_3366 ( N_noxref_12_c_4260_p N_noxref_13_M29_noxref_d ) capacitor \
 c=0.00546784f //x=47.35 //y=1.57 //x2=47.425 //y2=0.915
cc_3367 ( N_noxref_12_c_4261_p N_noxref_13_M29_noxref_d ) capacitor \
 c=0.00241102f //x=47.725 //y=0.76 //x2=47.425 //y2=0.915
cc_3368 ( N_noxref_12_c_4249_p N_noxref_13_M29_noxref_d ) capacitor \
 c=0.0138621f //x=47.725 //y=1.415 //x2=47.425 //y2=0.915
cc_3369 ( N_noxref_12_c_4263_p N_noxref_13_M29_noxref_d ) capacitor \
 c=0.00219619f //x=47.88 //y=0.915 //x2=47.425 //y2=0.915
cc_3370 ( N_noxref_12_c_4250_p N_noxref_13_M29_noxref_d ) capacitor \
 c=0.00603828f //x=47.88 //y=1.26 //x2=47.425 //y2=0.915
cc_3371 ( N_noxref_12_c_4254_p N_noxref_13_M29_noxref_d ) capacitor \
 c=0.00661782f //x=47.36 //y=1.915 //x2=47.425 //y2=0.915
cc_3372 ( N_noxref_12_M110_noxref_g N_noxref_13_M110_noxref_d ) capacitor \
 c=0.0180032f //x=47.1 //y=6.02 //x2=47.175 //y2=5.02
cc_3373 ( N_noxref_12_M111_noxref_g N_noxref_13_M110_noxref_d ) capacitor \
 c=0.0194246f //x=47.54 //y=6.02 //x2=47.175 //y2=5.02
cc_3374 ( N_noxref_12_c_4157_n N_D_c_4909_n ) capacitor c=0.0358131f \
 //x=35.775 //y=3.7 //x2=49.835 //y2=2.96
cc_3375 ( N_noxref_12_c_4200_n N_D_c_4909_n ) capacitor c=8.32553e-19 \
 //x=31.195 //y=3.7 //x2=49.835 //y2=2.96
cc_3376 ( N_noxref_12_c_4162_n N_D_c_4909_n ) capacitor c=0.0288894f \
 //x=39.845 //y=3.7 //x2=49.835 //y2=2.96
cc_3377 ( N_noxref_12_c_4164_n N_D_c_4909_n ) capacitor c=6.03896e-19 \
 //x=36.005 //y=3.7 //x2=49.835 //y2=2.96
cc_3378 ( N_noxref_12_c_4204_n N_D_c_4909_n ) capacitor c=0.05455f //x=47.245 \
 //y=3.7 //x2=49.835 //y2=2.96
cc_3379 ( N_noxref_12_c_4206_n N_D_c_4909_n ) capacitor c=5.76918e-19 \
 //x=40.075 //y=3.7 //x2=49.835 //y2=2.96
cc_3380 ( N_noxref_12_c_4111_n N_D_c_4909_n ) capacitor c=0.0179917f //x=31.08 \
 //y=2.08 //x2=49.835 //y2=2.96
cc_3381 ( N_noxref_12_c_4112_n N_D_c_4909_n ) capacitor c=0.0202855f //x=35.89 \
 //y=2.08 //x2=49.835 //y2=2.96
cc_3382 ( N_noxref_12_c_4114_n N_D_c_4909_n ) capacitor c=0.021075f //x=39.96 \
 //y=3.7 //x2=49.835 //y2=2.96
cc_3383 ( N_noxref_12_c_4115_n N_D_c_4909_n ) capacitor c=0.0202855f //x=47.36 \
 //y=2.08 //x2=49.835 //y2=2.96
cc_3384 ( N_noxref_12_c_4115_n N_D_c_4917_n ) capacitor c=9.78855e-19 \
 //x=47.36 //y=2.08 //x2=49.95 //y2=2.08
cc_3385 ( N_noxref_12_c_4157_n N_CLK_c_5668_n ) capacitor c=0.0345106f \
 //x=35.775 //y=3.7 //x2=39.105 //y2=4.44
cc_3386 ( N_noxref_12_c_4200_n N_CLK_c_5668_n ) capacitor c=7.0371e-19 \
 //x=31.195 //y=3.7 //x2=39.105 //y2=4.44
cc_3387 ( N_noxref_12_c_4162_n N_CLK_c_5668_n ) capacitor c=0.02107f \
 //x=39.845 //y=3.7 //x2=39.105 //y2=4.44
cc_3388 ( N_noxref_12_c_4164_n N_CLK_c_5668_n ) capacitor c=4.78625e-19 \
 //x=36.005 //y=3.7 //x2=39.105 //y2=4.44
cc_3389 ( N_noxref_12_c_4111_n N_CLK_c_5668_n ) capacitor c=0.0200057f \
 //x=31.08 //y=2.08 //x2=39.105 //y2=4.44
cc_3390 ( N_noxref_12_c_4112_n N_CLK_c_5668_n ) capacitor c=0.0200057f \
 //x=35.89 //y=2.08 //x2=39.105 //y2=4.44
cc_3391 ( N_noxref_12_c_4125_n N_CLK_c_5668_n ) capacitor c=0.0172877f \
 //x=38.685 //y=5.2 //x2=39.105 //y2=4.44
cc_3392 ( N_noxref_12_c_4233_n N_CLK_c_5668_n ) capacitor c=0.0111881f \
 //x=31.08 //y=4.7 //x2=39.105 //y2=4.44
cc_3393 ( N_noxref_12_c_4191_n N_CLK_c_5668_n ) capacitor c=0.0111881f \
 //x=35.89 //y=4.7 //x2=39.105 //y2=4.44
cc_3394 ( N_noxref_12_c_4111_n N_CLK_c_5679_n ) capacitor c=0.00153281f \
 //x=31.08 //y=2.08 //x2=30.085 //y2=4.44
cc_3395 ( N_noxref_12_c_4162_n N_CLK_c_5680_n ) capacitor c=0.0050622f \
 //x=39.845 //y=3.7 //x2=54.275 //y2=4.44
cc_3396 ( N_noxref_12_c_4204_n N_CLK_c_5680_n ) capacitor c=0.0653647f \
 //x=47.245 //y=3.7 //x2=54.275 //y2=4.44
cc_3397 ( N_noxref_12_c_4206_n N_CLK_c_5680_n ) capacitor c=5.69483e-19 \
 //x=40.075 //y=3.7 //x2=54.275 //y2=4.44
cc_3398 ( N_noxref_12_c_4121_n N_CLK_c_5680_n ) capacitor c=0.0173598f \
 //x=39.395 //y=5.2 //x2=54.275 //y2=4.44
cc_3399 ( N_noxref_12_c_4114_n N_CLK_c_5680_n ) capacitor c=0.0208321f \
 //x=39.96 //y=3.7 //x2=54.275 //y2=4.44
cc_3400 ( N_noxref_12_c_4115_n N_CLK_c_5680_n ) capacitor c=0.0200057f \
 //x=47.36 //y=2.08 //x2=54.275 //y2=4.44
cc_3401 ( N_noxref_12_c_4248_p N_CLK_c_5680_n ) capacitor c=0.0111881f \
 //x=47.36 //y=4.7 //x2=54.275 //y2=4.44
cc_3402 ( N_noxref_12_c_4162_n N_CLK_c_5704_n ) capacitor c=5.12294e-19 \
 //x=39.845 //y=3.7 //x2=39.335 //y2=4.44
cc_3403 ( N_noxref_12_c_4121_n N_CLK_c_5704_n ) capacitor c=0.0023575f \
 //x=39.395 //y=5.2 //x2=39.335 //y2=4.44
cc_3404 ( N_noxref_12_c_4114_n N_CLK_c_5704_n ) capacitor c=0.00151334f \
 //x=39.96 //y=3.7 //x2=39.335 //y2=4.44
cc_3405 ( N_noxref_12_c_4200_n N_CLK_c_5625_n ) capacitor c=0.00526349f \
 //x=31.195 //y=3.7 //x2=29.97 //y2=2.08
cc_3406 ( N_noxref_12_c_4111_n N_CLK_c_5625_n ) capacitor c=0.0422302f \
 //x=31.08 //y=2.08 //x2=29.97 //y2=2.08
cc_3407 ( N_noxref_12_c_4230_n N_CLK_c_5625_n ) capacitor c=0.00201097f \
 //x=31.08 //y=2.08 //x2=29.97 //y2=2.08
cc_3408 ( N_noxref_12_c_4233_n N_CLK_c_5625_n ) capacitor c=0.00218014f \
 //x=31.08 //y=4.7 //x2=29.97 //y2=2.08
cc_3409 ( N_noxref_12_c_4121_n N_CLK_c_5947_n ) capacitor c=0.0126974f \
 //x=39.395 //y=5.2 //x2=39.22 //y2=4.535
cc_3410 ( N_noxref_12_c_4114_n N_CLK_c_5947_n ) capacitor c=0.00923416f \
 //x=39.96 //y=3.7 //x2=39.22 //y2=4.535
cc_3411 ( N_noxref_12_c_4162_n N_CLK_c_5626_n ) capacitor c=0.0169594f \
 //x=39.845 //y=3.7 //x2=39.22 //y2=2.08
cc_3412 ( N_noxref_12_c_4206_n N_CLK_c_5626_n ) capacitor c=0.00117715f \
 //x=40.075 //y=3.7 //x2=39.22 //y2=2.08
cc_3413 ( N_noxref_12_c_4121_n N_CLK_c_5626_n ) capacitor c=3.74769e-19 \
 //x=39.395 //y=5.2 //x2=39.22 //y2=2.08
cc_3414 ( N_noxref_12_c_4114_n N_CLK_c_5626_n ) capacitor c=0.0679995f \
 //x=39.96 //y=3.7 //x2=39.22 //y2=2.08
cc_3415 ( N_noxref_12_M90_noxref_g N_CLK_M88_noxref_g ) capacitor c=0.0101598f \
 //x=30.82 //y=6.02 //x2=29.94 //y2=6.02
cc_3416 ( N_noxref_12_M90_noxref_g N_CLK_M89_noxref_g ) capacitor c=0.0602553f \
 //x=30.82 //y=6.02 //x2=30.38 //y2=6.02
cc_3417 ( N_noxref_12_M91_noxref_g N_CLK_M89_noxref_g ) capacitor c=0.0101598f \
 //x=31.26 //y=6.02 //x2=30.38 //y2=6.02
cc_3418 ( N_noxref_12_c_4121_n N_CLK_M100_noxref_g ) capacitor c=0.0166421f \
 //x=39.395 //y=5.2 //x2=39.26 //y2=6.02
cc_3419 ( N_noxref_12_M100_noxref_d N_CLK_M100_noxref_g ) capacitor \
 c=0.0173476f //x=39.335 //y=5.02 //x2=39.26 //y2=6.02
cc_3420 ( N_noxref_12_c_4127_n N_CLK_M101_noxref_g ) capacitor c=0.018922f \
 //x=39.875 //y=5.2 //x2=39.7 //y2=6.02
cc_3421 ( N_noxref_12_M100_noxref_d N_CLK_M101_noxref_g ) capacitor \
 c=0.0179769f //x=39.335 //y=5.02 //x2=39.7 //y2=6.02
cc_3422 ( N_noxref_12_c_4221_n N_CLK_c_5931_n ) capacitor c=0.00456962f \
 //x=31.07 //y=0.915 //x2=30.06 //y2=0.91
cc_3423 ( N_noxref_12_c_4222_n N_CLK_c_5932_n ) capacitor c=0.00438372f \
 //x=31.07 //y=1.26 //x2=30.06 //y2=1.22
cc_3424 ( N_noxref_12_c_4223_n N_CLK_c_5933_n ) capacitor c=0.00438372f \
 //x=31.07 //y=1.57 //x2=30.06 //y2=1.45
cc_3425 ( N_noxref_12_c_4111_n N_CLK_c_5934_n ) capacitor c=0.00205895f \
 //x=31.08 //y=2.08 //x2=30.06 //y2=1.915
cc_3426 ( N_noxref_12_c_4230_n N_CLK_c_5934_n ) capacitor c=0.00828003f \
 //x=31.08 //y=2.08 //x2=30.06 //y2=1.915
cc_3427 ( N_noxref_12_c_4231_n N_CLK_c_5934_n ) capacitor c=0.00438372f \
 //x=31.08 //y=1.915 //x2=30.06 //y2=1.915
cc_3428 ( N_noxref_12_c_4233_n N_CLK_c_6000_n ) capacitor c=0.0611812f \
 //x=31.08 //y=4.7 //x2=30.305 //y2=4.79
cc_3429 ( N_noxref_12_M24_noxref_d N_CLK_c_5956_n ) capacitor c=0.00217566f \
 //x=39.33 //y=0.905 //x2=39.255 //y2=0.905
cc_3430 ( N_noxref_12_M24_noxref_d N_CLK_c_5959_n ) capacitor c=0.0034598f \
 //x=39.33 //y=0.905 //x2=39.255 //y2=1.25
cc_3431 ( N_noxref_12_M24_noxref_d N_CLK_c_5961_n ) capacitor c=0.00669531f \
 //x=39.33 //y=0.905 //x2=39.255 //y2=1.56
cc_3432 ( N_noxref_12_c_4114_n N_CLK_c_6054_n ) capacitor c=0.0142673f \
 //x=39.96 //y=3.7 //x2=39.625 //y2=4.79
cc_3433 ( N_noxref_12_c_4327_p N_CLK_c_6054_n ) capacitor c=0.00407665f \
 //x=39.48 //y=5.2 //x2=39.625 //y2=4.79
cc_3434 ( N_noxref_12_M24_noxref_d N_CLK_c_6056_n ) capacitor c=0.00241102f \
 //x=39.33 //y=0.905 //x2=39.63 //y2=0.75
cc_3435 ( N_noxref_12_c_4113_n N_CLK_c_6057_n ) capacitor c=0.00371277f \
 //x=39.875 //y=1.655 //x2=39.63 //y2=1.405
cc_3436 ( N_noxref_12_M24_noxref_d N_CLK_c_6057_n ) capacitor c=0.0137169f \
 //x=39.33 //y=0.905 //x2=39.63 //y2=1.405
cc_3437 ( N_noxref_12_M24_noxref_d N_CLK_c_5964_n ) capacitor c=0.00132245f \
 //x=39.33 //y=0.905 //x2=39.785 //y2=0.905
cc_3438 ( N_noxref_12_c_4113_n N_CLK_c_5965_n ) capacitor c=0.00457401f \
 //x=39.875 //y=1.655 //x2=39.785 //y2=1.25
cc_3439 ( N_noxref_12_M24_noxref_d N_CLK_c_5965_n ) capacitor c=0.00566463f \
 //x=39.33 //y=0.905 //x2=39.785 //y2=1.25
cc_3440 ( N_noxref_12_c_4111_n N_CLK_c_5936_n ) capacitor c=0.00142741f \
 //x=31.08 //y=2.08 //x2=29.97 //y2=4.7
cc_3441 ( N_noxref_12_c_4233_n N_CLK_c_5936_n ) capacitor c=0.00487508f \
 //x=31.08 //y=4.7 //x2=29.97 //y2=4.7
cc_3442 ( N_noxref_12_c_4114_n N_CLK_c_5966_n ) capacitor c=0.00731987f \
 //x=39.96 //y=3.7 //x2=39.22 //y2=2.08
cc_3443 ( N_noxref_12_c_4114_n N_CLK_c_6065_n ) capacitor c=0.00306024f \
 //x=39.96 //y=3.7 //x2=39.22 //y2=1.915
cc_3444 ( N_noxref_12_M24_noxref_d N_CLK_c_6065_n ) capacitor c=0.00660593f \
 //x=39.33 //y=0.905 //x2=39.22 //y2=1.915
cc_3445 ( N_noxref_12_c_4121_n N_CLK_c_5968_n ) capacitor c=0.00346519f \
 //x=39.395 //y=5.2 //x2=39.25 //y2=4.7
cc_3446 ( N_noxref_12_c_4114_n N_CLK_c_5968_n ) capacitor c=0.00518077f \
 //x=39.96 //y=3.7 //x2=39.25 //y2=4.7
cc_3447 ( N_noxref_12_c_4111_n N_SN_c_6844_n ) capacitor c=0.0186201f \
 //x=31.08 //y=2.08 //x2=34.665 //y2=2.22
cc_3448 ( N_noxref_12_c_4225_n N_SN_c_6844_n ) capacitor c=3.13485e-19 \
 //x=31.445 //y=1.415 //x2=34.665 //y2=2.22
cc_3449 ( N_noxref_12_c_4230_n N_SN_c_6844_n ) capacitor c=0.00584491f \
 //x=31.08 //y=2.08 //x2=34.665 //y2=2.22
cc_3450 ( N_noxref_12_c_4112_n N_SN_c_6855_n ) capacitor c=0.0209607f \
 //x=35.89 //y=2.08 //x2=46.135 //y2=2.22
cc_3451 ( N_noxref_12_c_4345_p N_SN_c_6855_n ) capacitor c=0.0146822f \
 //x=39.605 //y=1.655 //x2=46.135 //y2=2.22
cc_3452 ( N_noxref_12_c_4114_n N_SN_c_6855_n ) capacitor c=0.0222456f \
 //x=39.96 //y=3.7 //x2=46.135 //y2=2.22
cc_3453 ( N_noxref_12_c_4183_n N_SN_c_6855_n ) capacitor c=3.13485e-19 \
 //x=36.255 //y=1.415 //x2=46.135 //y2=2.22
cc_3454 ( N_noxref_12_c_4188_n N_SN_c_6855_n ) capacitor c=0.00584491f \
 //x=35.89 //y=2.08 //x2=46.135 //y2=2.22
cc_3455 ( N_noxref_12_c_4112_n N_SN_c_6865_n ) capacitor c=0.00165648f \
 //x=35.89 //y=2.08 //x2=34.895 //y2=2.22
cc_3456 ( N_noxref_12_c_4188_n N_SN_c_6865_n ) capacitor c=2.3323e-19 \
 //x=35.89 //y=2.08 //x2=34.895 //y2=2.22
cc_3457 ( N_noxref_12_c_4115_n N_SN_c_6866_n ) capacitor c=0.0209607f \
 //x=47.36 //y=2.08 //x2=59.085 //y2=2.22
cc_3458 ( N_noxref_12_c_4249_p N_SN_c_6866_n ) capacitor c=3.13485e-19 \
 //x=47.725 //y=1.415 //x2=59.085 //y2=2.22
cc_3459 ( N_noxref_12_c_4253_p N_SN_c_6866_n ) capacitor c=0.00584491f \
 //x=47.36 //y=2.08 //x2=59.085 //y2=2.22
cc_3460 ( N_noxref_12_c_4115_n N_SN_c_6876_n ) capacitor c=0.00165648f \
 //x=47.36 //y=2.08 //x2=46.365 //y2=2.22
cc_3461 ( N_noxref_12_c_4253_p N_SN_c_6876_n ) capacitor c=2.3323e-19 \
 //x=47.36 //y=2.08 //x2=46.365 //y2=2.22
cc_3462 ( N_noxref_12_c_4157_n N_SN_c_6890_n ) capacitor c=0.0190398f \
 //x=35.775 //y=3.7 //x2=34.78 //y2=2.08
cc_3463 ( N_noxref_12_c_4164_n N_SN_c_6890_n ) capacitor c=0.00128547f \
 //x=36.005 //y=3.7 //x2=34.78 //y2=2.08
cc_3464 ( N_noxref_12_c_4112_n N_SN_c_6890_n ) capacitor c=0.0433248f \
 //x=35.89 //y=2.08 //x2=34.78 //y2=2.08
cc_3465 ( N_noxref_12_c_4188_n N_SN_c_6890_n ) capacitor c=0.0019893f \
 //x=35.89 //y=2.08 //x2=34.78 //y2=2.08
cc_3466 ( N_noxref_12_c_4191_n N_SN_c_6890_n ) capacitor c=0.00219458f \
 //x=35.89 //y=4.7 //x2=34.78 //y2=2.08
cc_3467 ( N_noxref_12_c_4204_n N_SN_c_6891_n ) capacitor c=0.0203253f \
 //x=47.245 //y=3.7 //x2=46.25 //y2=2.08
cc_3468 ( N_noxref_12_c_4115_n N_SN_c_6891_n ) capacitor c=0.0432458f \
 //x=47.36 //y=2.08 //x2=46.25 //y2=2.08
cc_3469 ( N_noxref_12_c_4253_p N_SN_c_6891_n ) capacitor c=0.0019893f \
 //x=47.36 //y=2.08 //x2=46.25 //y2=2.08
cc_3470 ( N_noxref_12_c_4248_p N_SN_c_6891_n ) capacitor c=0.00219458f \
 //x=47.36 //y=4.7 //x2=46.25 //y2=2.08
cc_3471 ( N_noxref_12_M96_noxref_g N_SN_M94_noxref_g ) capacitor c=0.0101598f \
 //x=35.63 //y=6.02 //x2=34.75 //y2=6.02
cc_3472 ( N_noxref_12_M96_noxref_g N_SN_M95_noxref_g ) capacitor c=0.0602553f \
 //x=35.63 //y=6.02 //x2=35.19 //y2=6.02
cc_3473 ( N_noxref_12_M97_noxref_g N_SN_M95_noxref_g ) capacitor c=0.0101598f \
 //x=36.07 //y=6.02 //x2=35.19 //y2=6.02
cc_3474 ( N_noxref_12_M110_noxref_g N_SN_M108_noxref_g ) capacitor \
 c=0.0101598f //x=47.1 //y=6.02 //x2=46.22 //y2=6.02
cc_3475 ( N_noxref_12_M110_noxref_g N_SN_M109_noxref_g ) capacitor \
 c=0.0602553f //x=47.1 //y=6.02 //x2=46.66 //y2=6.02
cc_3476 ( N_noxref_12_M111_noxref_g N_SN_M109_noxref_g ) capacitor \
 c=0.0101598f //x=47.54 //y=6.02 //x2=46.66 //y2=6.02
cc_3477 ( N_noxref_12_c_4179_n N_SN_c_7075_n ) capacitor c=0.00456962f \
 //x=35.88 //y=0.915 //x2=34.87 //y2=0.91
cc_3478 ( N_noxref_12_c_4180_n N_SN_c_7076_n ) capacitor c=0.00438372f \
 //x=35.88 //y=1.26 //x2=34.87 //y2=1.22
cc_3479 ( N_noxref_12_c_4181_n N_SN_c_7077_n ) capacitor c=0.00438372f \
 //x=35.88 //y=1.57 //x2=34.87 //y2=1.45
cc_3480 ( N_noxref_12_c_4112_n N_SN_c_7078_n ) capacitor c=0.00205895f \
 //x=35.89 //y=2.08 //x2=34.87 //y2=1.915
cc_3481 ( N_noxref_12_c_4188_n N_SN_c_7078_n ) capacitor c=0.00828003f \
 //x=35.89 //y=2.08 //x2=34.87 //y2=1.915
cc_3482 ( N_noxref_12_c_4189_n N_SN_c_7078_n ) capacitor c=0.00438372f \
 //x=35.89 //y=1.915 //x2=34.87 //y2=1.915
cc_3483 ( N_noxref_12_c_4191_n N_SN_c_7095_n ) capacitor c=0.0611812f \
 //x=35.89 //y=4.7 //x2=35.115 //y2=4.79
cc_3484 ( N_noxref_12_c_4258_p N_SN_c_7128_n ) capacitor c=0.00456962f \
 //x=47.35 //y=0.915 //x2=46.34 //y2=0.91
cc_3485 ( N_noxref_12_c_4259_p N_SN_c_7129_n ) capacitor c=0.00438372f \
 //x=47.35 //y=1.26 //x2=46.34 //y2=1.22
cc_3486 ( N_noxref_12_c_4260_p N_SN_c_7130_n ) capacitor c=0.00438372f \
 //x=47.35 //y=1.57 //x2=46.34 //y2=1.45
cc_3487 ( N_noxref_12_c_4115_n N_SN_c_7131_n ) capacitor c=0.00205895f \
 //x=47.36 //y=2.08 //x2=46.34 //y2=1.915
cc_3488 ( N_noxref_12_c_4253_p N_SN_c_7131_n ) capacitor c=0.00828003f \
 //x=47.36 //y=2.08 //x2=46.34 //y2=1.915
cc_3489 ( N_noxref_12_c_4254_p N_SN_c_7131_n ) capacitor c=0.00438372f \
 //x=47.36 //y=1.915 //x2=46.34 //y2=1.915
cc_3490 ( N_noxref_12_c_4248_p N_SN_c_7179_n ) capacitor c=0.0611812f \
 //x=47.36 //y=4.7 //x2=46.585 //y2=4.79
cc_3491 ( N_noxref_12_c_4112_n N_SN_c_7080_n ) capacitor c=0.00142741f \
 //x=35.89 //y=2.08 //x2=34.78 //y2=4.7
cc_3492 ( N_noxref_12_c_4191_n N_SN_c_7080_n ) capacitor c=0.00487508f \
 //x=35.89 //y=4.7 //x2=34.78 //y2=4.7
cc_3493 ( N_noxref_12_c_4115_n N_SN_c_7133_n ) capacitor c=0.00142741f \
 //x=47.36 //y=2.08 //x2=46.25 //y2=4.7
cc_3494 ( N_noxref_12_c_4248_p N_SN_c_7133_n ) capacitor c=0.00487508f \
 //x=47.36 //y=4.7 //x2=46.25 //y2=4.7
cc_3495 ( N_noxref_12_c_4157_n N_noxref_24_c_8424_n ) capacitor c=0.404606f \
 //x=35.775 //y=3.7 //x2=79.065 //y2=3.33
cc_3496 ( N_noxref_12_c_4200_n N_noxref_24_c_8424_n ) capacitor c=0.029444f \
 //x=31.195 //y=3.7 //x2=79.065 //y2=3.33
cc_3497 ( N_noxref_12_c_4162_n N_noxref_24_c_8424_n ) capacitor c=0.338821f \
 //x=39.845 //y=3.7 //x2=79.065 //y2=3.33
cc_3498 ( N_noxref_12_c_4164_n N_noxref_24_c_8424_n ) capacitor c=0.026734f \
 //x=36.005 //y=3.7 //x2=79.065 //y2=3.33
cc_3499 ( N_noxref_12_c_4204_n N_noxref_24_c_8424_n ) capacitor c=0.663837f \
 //x=47.245 //y=3.7 //x2=79.065 //y2=3.33
cc_3500 ( N_noxref_12_c_4206_n N_noxref_24_c_8424_n ) capacitor c=0.0266742f \
 //x=40.075 //y=3.7 //x2=79.065 //y2=3.33
cc_3501 ( N_noxref_12_c_4111_n N_noxref_24_c_8424_n ) capacitor c=0.0198536f \
 //x=31.08 //y=2.08 //x2=79.065 //y2=3.33
cc_3502 ( N_noxref_12_c_4112_n N_noxref_24_c_8424_n ) capacitor c=0.0198536f \
 //x=35.89 //y=2.08 //x2=79.065 //y2=3.33
cc_3503 ( N_noxref_12_c_4114_n N_noxref_24_c_8424_n ) capacitor c=0.0205775f \
 //x=39.96 //y=3.7 //x2=79.065 //y2=3.33
cc_3504 ( N_noxref_12_c_4115_n N_noxref_24_c_8424_n ) capacitor c=0.0198536f \
 //x=47.36 //y=2.08 //x2=79.065 //y2=3.33
cc_3505 ( N_noxref_12_c_4111_n N_noxref_38_c_9797_n ) capacitor c=0.00204385f \
 //x=31.08 //y=2.08 //x2=31.735 //y2=0.54
cc_3506 ( N_noxref_12_c_4221_n N_noxref_38_c_9797_n ) capacitor c=0.0194423f \
 //x=31.07 //y=0.915 //x2=31.735 //y2=0.54
cc_3507 ( N_noxref_12_c_4227_n N_noxref_38_c_9797_n ) capacitor c=0.00656458f \
 //x=31.6 //y=0.915 //x2=31.735 //y2=0.54
cc_3508 ( N_noxref_12_c_4230_n N_noxref_38_c_9797_n ) capacitor c=2.20712e-19 \
 //x=31.08 //y=2.08 //x2=31.735 //y2=0.54
cc_3509 ( N_noxref_12_c_4222_n N_noxref_38_c_9807_n ) capacitor c=0.00538033f \
 //x=31.07 //y=1.26 //x2=30.85 //y2=0.995
cc_3510 ( N_noxref_12_c_4221_n N_noxref_38_M19_noxref_s ) capacitor \
 c=0.00538033f //x=31.07 //y=0.915 //x2=30.715 //y2=0.375
cc_3511 ( N_noxref_12_c_4223_n N_noxref_38_M19_noxref_s ) capacitor \
 c=0.00538033f //x=31.07 //y=1.57 //x2=30.715 //y2=0.375
cc_3512 ( N_noxref_12_c_4227_n N_noxref_38_M19_noxref_s ) capacitor \
 c=0.0143002f //x=31.6 //y=0.915 //x2=30.715 //y2=0.375
cc_3513 ( N_noxref_12_c_4228_n N_noxref_38_M19_noxref_s ) capacitor \
 c=0.00290153f //x=31.6 //y=1.26 //x2=30.715 //y2=0.375
cc_3514 ( N_noxref_12_c_4112_n N_noxref_40_c_9901_n ) capacitor c=0.00204385f \
 //x=35.89 //y=2.08 //x2=36.545 //y2=0.54
cc_3515 ( N_noxref_12_c_4179_n N_noxref_40_c_9901_n ) capacitor c=0.0194423f \
 //x=35.88 //y=0.915 //x2=36.545 //y2=0.54
cc_3516 ( N_noxref_12_c_4185_n N_noxref_40_c_9901_n ) capacitor c=0.00656458f \
 //x=36.41 //y=0.915 //x2=36.545 //y2=0.54
cc_3517 ( N_noxref_12_c_4188_n N_noxref_40_c_9901_n ) capacitor c=2.20712e-19 \
 //x=35.89 //y=2.08 //x2=36.545 //y2=0.54
cc_3518 ( N_noxref_12_c_4180_n N_noxref_40_c_9911_n ) capacitor c=0.00538829f \
 //x=35.88 //y=1.26 //x2=35.66 //y2=0.995
cc_3519 ( N_noxref_12_c_4179_n N_noxref_40_M22_noxref_s ) capacitor \
 c=0.00538829f //x=35.88 //y=0.915 //x2=35.525 //y2=0.375
cc_3520 ( N_noxref_12_c_4181_n N_noxref_40_M22_noxref_s ) capacitor \
 c=0.00538829f //x=35.88 //y=1.57 //x2=35.525 //y2=0.375
cc_3521 ( N_noxref_12_c_4185_n N_noxref_40_M22_noxref_s ) capacitor \
 c=0.0143002f //x=36.41 //y=0.915 //x2=35.525 //y2=0.375
cc_3522 ( N_noxref_12_c_4186_n N_noxref_40_M22_noxref_s ) capacitor \
 c=0.00290153f //x=36.41 //y=1.26 //x2=35.525 //y2=0.375
cc_3523 ( N_noxref_12_c_4345_p N_noxref_41_c_9966_n ) capacitor c=3.15806e-19 \
 //x=39.605 //y=1.655 //x2=38.065 //y2=1.495
cc_3524 ( N_noxref_12_c_4345_p N_noxref_41_c_9955_n ) capacitor c=0.020324f \
 //x=39.605 //y=1.655 //x2=39.035 //y2=1.495
cc_3525 ( N_noxref_12_c_4113_n N_noxref_41_c_9956_n ) capacitor c=0.00457164f \
 //x=39.875 //y=1.655 //x2=39.92 //y2=0.53
cc_3526 ( N_noxref_12_M24_noxref_d N_noxref_41_c_9956_n ) capacitor \
 c=0.0115831f //x=39.33 //y=0.905 //x2=39.92 //y2=0.53
cc_3527 ( N_noxref_12_c_4113_n N_noxref_41_M23_noxref_s ) capacitor \
 c=0.013435f //x=39.875 //y=1.655 //x2=37.93 //y2=0.365
cc_3528 ( N_noxref_12_M24_noxref_d N_noxref_41_M23_noxref_s ) capacitor \
 c=0.0439476f //x=39.33 //y=0.905 //x2=37.93 //y2=0.365
cc_3529 ( N_noxref_12_c_4113_n N_noxref_42_c_10017_n ) capacitor c=3.22188e-19 \
 //x=39.875 //y=1.655 //x2=41.395 //y2=1.495
cc_3530 ( N_noxref_12_c_4115_n N_noxref_44_c_10107_n ) capacitor c=0.00204385f \
 //x=47.36 //y=2.08 //x2=48.015 //y2=0.54
cc_3531 ( N_noxref_12_c_4258_p N_noxref_44_c_10107_n ) capacitor c=0.0194423f \
 //x=47.35 //y=0.915 //x2=48.015 //y2=0.54
cc_3532 ( N_noxref_12_c_4263_p N_noxref_44_c_10107_n ) capacitor c=0.00656458f \
 //x=47.88 //y=0.915 //x2=48.015 //y2=0.54
cc_3533 ( N_noxref_12_c_4253_p N_noxref_44_c_10107_n ) capacitor c=2.20712e-19 \
 //x=47.36 //y=2.08 //x2=48.015 //y2=0.54
cc_3534 ( N_noxref_12_c_4259_p N_noxref_44_c_10119_n ) capacitor c=0.00538829f \
 //x=47.35 //y=1.26 //x2=47.13 //y2=0.995
cc_3535 ( N_noxref_12_c_4258_p N_noxref_44_M29_noxref_s ) capacitor \
 c=0.00538829f //x=47.35 //y=0.915 //x2=46.995 //y2=0.375
cc_3536 ( N_noxref_12_c_4260_p N_noxref_44_M29_noxref_s ) capacitor \
 c=0.00538829f //x=47.35 //y=1.57 //x2=46.995 //y2=0.375
cc_3537 ( N_noxref_12_c_4263_p N_noxref_44_M29_noxref_s ) capacitor \
 c=0.0143002f //x=47.88 //y=0.915 //x2=46.995 //y2=0.375
cc_3538 ( N_noxref_12_c_4250_p N_noxref_44_M29_noxref_s ) capacitor \
 c=0.00290153f //x=47.88 //y=1.26 //x2=46.995 //y2=0.375
cc_3539 ( N_noxref_13_c_4455_n N_D_c_4909_n ) capacitor c=0.00415759f \
 //x=47.985 //y=4.07 //x2=49.835 //y2=2.96
cc_3540 ( N_noxref_13_c_4433_n N_D_c_4909_n ) capacitor c=0.172149f //x=50.605 \
 //y=2.59 //x2=49.835 //y2=2.96
cc_3541 ( N_noxref_13_c_4434_n N_D_c_4909_n ) capacitor c=0.0293832f \
 //x=48.215 //y=2.59 //x2=49.835 //y2=2.96
cc_3542 ( N_noxref_13_c_4602_p N_D_c_4909_n ) capacitor c=0.00137661f \
 //x=50.69 //y=2.875 //x2=49.835 //y2=2.96
cc_3543 ( N_noxref_13_c_4603_p N_D_c_4909_n ) capacitor c=0.0145308f \
 //x=50.775 //y=2.96 //x2=49.835 //y2=2.96
cc_3544 ( N_noxref_13_c_4445_n N_D_c_4909_n ) capacitor c=0.0192451f //x=42.55 \
 //y=2.08 //x2=49.835 //y2=2.96
cc_3545 ( N_noxref_13_c_4448_n N_D_c_4909_n ) capacitor c=0.0212233f //x=48.1 \
 //y=2.59 //x2=49.835 //y2=2.96
cc_3546 ( N_noxref_13_c_4455_n N_D_c_4917_n ) capacitor c=0.00103915f \
 //x=47.985 //y=4.07 //x2=49.95 //y2=2.08
cc_3547 ( N_noxref_13_c_4433_n N_D_c_4917_n ) capacitor c=0.0196218f \
 //x=50.605 //y=2.59 //x2=49.95 //y2=2.08
cc_3548 ( N_noxref_13_c_4602_p N_D_c_4917_n ) capacitor c=0.00488481f \
 //x=50.69 //y=2.875 //x2=49.95 //y2=2.08
cc_3549 ( N_noxref_13_c_4603_p N_D_c_4917_n ) capacitor c=4.93246e-19 \
 //x=50.775 //y=2.96 //x2=49.95 //y2=2.08
cc_3550 ( N_noxref_13_c_4448_n N_D_c_4917_n ) capacitor c=0.0127927f //x=48.1 \
 //y=2.59 //x2=49.95 //y2=2.08
cc_3551 ( N_noxref_13_c_4435_n N_noxref_15_c_5221_n ) capacitor c=0.143317f \
 //x=74.995 //y=2.96 //x2=53.135 //y2=2.59
cc_3552 ( N_noxref_13_c_4433_n N_noxref_15_c_5222_n ) capacitor c=0.0143981f \
 //x=50.605 //y=2.59 //x2=51.545 //y2=2.59
cc_3553 ( N_noxref_13_c_4434_n N_noxref_15_c_5222_n ) capacitor c=3.63347e-19 \
 //x=48.215 //y=2.59 //x2=51.545 //y2=2.59
cc_3554 ( N_noxref_13_c_4602_p N_noxref_15_c_5222_n ) capacitor c=0.00135108f \
 //x=50.69 //y=2.875 //x2=51.545 //y2=2.59
cc_3555 ( N_noxref_13_c_4435_n N_noxref_15_c_5222_n ) capacitor c=0.0293646f \
 //x=74.995 //y=2.96 //x2=51.545 //y2=2.59
cc_3556 ( N_noxref_13_c_4435_n N_noxref_15_c_5223_n ) capacitor c=0.0294578f \
 //x=74.995 //y=2.96 //x2=57.975 //y2=2.59
cc_3557 ( N_noxref_13_c_4435_n N_noxref_15_c_5224_n ) capacitor c=0.426576f \
 //x=74.995 //y=2.96 //x2=53.545 //y2=2.59
cc_3558 ( N_noxref_13_c_4433_n N_noxref_15_c_5226_n ) capacitor c=0.00186213f \
 //x=50.605 //y=2.59 //x2=51.43 //y2=2.59
cc_3559 ( N_noxref_13_c_4602_p N_noxref_15_c_5226_n ) capacitor c=0.00366495f \
 //x=50.69 //y=2.875 //x2=51.43 //y2=2.59
cc_3560 ( N_noxref_13_c_4435_n N_noxref_15_c_5226_n ) capacitor c=0.0206018f \
 //x=74.995 //y=2.96 //x2=51.43 //y2=2.59
cc_3561 ( N_noxref_13_c_4448_n N_noxref_15_c_5226_n ) capacitor c=3.52729e-19 \
 //x=48.1 //y=2.59 //x2=51.43 //y2=2.59
cc_3562 ( N_noxref_13_c_4435_n N_noxref_15_c_5228_n ) capacitor c=0.0215953f \
 //x=74.995 //y=2.96 //x2=53.28 //y2=2.08
cc_3563 ( N_noxref_13_c_4435_n N_noxref_15_c_5229_n ) capacitor c=0.0215933f \
 //x=74.995 //y=2.96 //x2=58.09 //y2=2.08
cc_3564 ( N_noxref_13_c_4435_n N_noxref_16_c_5458_n ) capacitor c=0.172364f \
 //x=74.995 //y=2.96 //x2=62.785 //y2=2.59
cc_3565 ( N_noxref_13_c_4435_n N_noxref_16_c_5459_n ) capacitor c=0.0293832f \
 //x=74.995 //y=2.96 //x2=61.165 //y2=2.59
cc_3566 ( N_noxref_13_c_4435_n N_noxref_16_c_5461_n ) capacitor c=0.0206007f \
 //x=74.995 //y=2.96 //x2=61.05 //y2=2.59
cc_3567 ( N_noxref_13_c_4435_n N_noxref_16_c_5462_n ) capacitor c=0.0205791f \
 //x=74.995 //y=2.96 //x2=62.9 //y2=2.08
cc_3568 ( N_noxref_13_c_4455_n N_CLK_c_5680_n ) capacitor c=0.491575f \
 //x=47.985 //y=4.07 //x2=54.275 //y2=4.44
cc_3569 ( N_noxref_13_c_4513_n N_CLK_c_5680_n ) capacitor c=0.028941f \
 //x=42.665 //y=4.07 //x2=54.275 //y2=4.44
cc_3570 ( N_noxref_13_c_4433_n N_CLK_c_5680_n ) capacitor c=0.00190208f \
 //x=50.605 //y=2.59 //x2=54.275 //y2=4.44
cc_3571 ( N_noxref_13_c_4515_n N_CLK_c_5680_n ) capacitor c=0.0016972f \
 //x=42.55 //y=4.535 //x2=54.275 //y2=4.44
cc_3572 ( N_noxref_13_c_4445_n N_CLK_c_5680_n ) capacitor c=0.0207534f \
 //x=42.55 //y=2.08 //x2=54.275 //y2=4.44
cc_3573 ( N_noxref_13_c_4464_n N_CLK_c_5680_n ) capacitor c=0.032141f \
 //x=46.355 //y=5.155 //x2=54.275 //y2=4.44
cc_3574 ( N_noxref_13_c_4468_n N_CLK_c_5680_n ) capacitor c=0.0230136f \
 //x=45.645 //y=5.155 //x2=54.275 //y2=4.44
cc_3575 ( N_noxref_13_c_4474_n N_CLK_c_5680_n ) capacitor c=0.0183122f \
 //x=48.015 //y=5.155 //x2=54.275 //y2=4.44
cc_3576 ( N_noxref_13_c_4448_n N_CLK_c_5680_n ) capacitor c=0.022862f //x=48.1 \
 //y=2.59 //x2=54.275 //y2=4.44
cc_3577 ( N_noxref_13_c_4557_n N_CLK_c_5680_n ) capacitor c=0.00960248f \
 //x=42.955 //y=4.79 //x2=54.275 //y2=4.44
cc_3578 ( N_noxref_13_c_4535_n N_CLK_c_5680_n ) capacitor c=0.00203982f \
 //x=42.58 //y=4.7 //x2=54.275 //y2=4.44
cc_3579 ( N_noxref_13_c_4435_n N_CLK_c_5628_n ) capacitor c=0.0190322f \
 //x=74.995 //y=2.96 //x2=54.39 //y2=2.08
cc_3580 ( N_noxref_13_c_4435_n N_CLK_c_5629_n ) capacitor c=0.0192451f \
 //x=74.995 //y=2.96 //x2=63.64 //y2=2.08
cc_3581 ( N_noxref_13_c_4435_n N_noxref_18_c_6392_n ) capacitor c=0.0249192f \
 //x=74.995 //y=2.96 //x2=56.12 //y2=4.07
cc_3582 ( N_noxref_13_c_4455_n N_noxref_18_c_6449_n ) capacitor c=0.00649178f \
 //x=47.985 //y=4.07 //x2=50.805 //y2=4.07
cc_3583 ( N_noxref_13_c_4433_n N_noxref_18_c_6449_n ) capacitor c=2.82712e-19 \
 //x=50.605 //y=2.59 //x2=50.805 //y2=4.07
cc_3584 ( N_noxref_13_c_4433_n N_noxref_18_c_6377_n ) capacitor c=0.0114835f \
 //x=50.605 //y=2.59 //x2=50.69 //y2=2.08
cc_3585 ( N_noxref_13_c_4602_p N_noxref_18_c_6377_n ) capacitor c=0.00862629f \
 //x=50.69 //y=2.875 //x2=50.69 //y2=2.08
cc_3586 ( N_noxref_13_c_4603_p N_noxref_18_c_6377_n ) capacitor c=0.0115443f \
 //x=50.775 //y=2.96 //x2=50.69 //y2=2.08
cc_3587 ( N_noxref_13_c_4448_n N_noxref_18_c_6377_n ) capacitor c=9.45552e-19 \
 //x=48.1 //y=2.59 //x2=50.69 //y2=2.08
cc_3588 ( N_noxref_13_c_4435_n N_noxref_18_c_6380_n ) capacitor c=0.0210088f \
 //x=74.995 //y=2.96 //x2=66.23 //y2=2.08
cc_3589 ( N_noxref_13_c_4435_n N_noxref_18_c_6456_n ) capacitor c=0.0187394f \
 //x=74.995 //y=2.96 //x2=56.237 //y2=3.905
cc_3590 ( N_noxref_13_c_4435_n N_noxref_19_c_6669_n ) capacitor c=0.0211011f \
 //x=74.995 //y=2.96 //x2=67.71 //y2=4.81
cc_3591 ( N_noxref_13_c_4435_n N_noxref_19_c_6670_n ) capacitor c=0.0220754f \
 //x=74.995 //y=2.96 //x2=69.56 //y2=2.08
cc_3592 ( N_noxref_13_c_4445_n N_SN_c_6855_n ) capacitor c=0.0201924f \
 //x=42.55 //y=2.08 //x2=46.135 //y2=2.22
cc_3593 ( N_noxref_13_c_4560_n N_SN_c_6855_n ) capacitor c=3.11115e-19 \
 //x=42.96 //y=1.405 //x2=46.135 //y2=2.22
cc_3594 ( N_noxref_13_c_4533_n N_SN_c_6855_n ) capacitor c=0.00570799f \
 //x=42.55 //y=2.08 //x2=46.135 //y2=2.22
cc_3595 ( N_noxref_13_c_4433_n N_SN_c_6866_n ) capacitor c=0.223946f \
 //x=50.605 //y=2.59 //x2=59.085 //y2=2.22
cc_3596 ( N_noxref_13_c_4434_n N_SN_c_6866_n ) capacitor c=0.0291301f \
 //x=48.215 //y=2.59 //x2=59.085 //y2=2.22
cc_3597 ( N_noxref_13_c_4435_n N_SN_c_6866_n ) capacitor c=0.106844f \
 //x=74.995 //y=2.96 //x2=59.085 //y2=2.22
cc_3598 ( N_noxref_13_c_4658_p N_SN_c_6866_n ) capacitor c=0.016327f //x=47.7 \
 //y=1.665 //x2=59.085 //y2=2.22
cc_3599 ( N_noxref_13_c_4448_n N_SN_c_6866_n ) capacitor c=0.0215653f //x=48.1 \
 //y=2.59 //x2=59.085 //y2=2.22
cc_3600 ( N_noxref_13_c_4435_n N_SN_c_6877_n ) capacitor c=0.408366f \
 //x=74.995 //y=2.96 //x2=70.555 //y2=2.22
cc_3601 ( N_noxref_13_c_4435_n N_SN_c_6887_n ) capacitor c=0.0120222f \
 //x=74.995 //y=2.96 //x2=59.315 //y2=2.22
cc_3602 ( N_noxref_13_c_4455_n N_SN_c_6891_n ) capacitor c=0.0190126f \
 //x=47.985 //y=4.07 //x2=46.25 //y2=2.08
cc_3603 ( N_noxref_13_c_4464_n N_SN_c_6891_n ) capacitor c=0.0146f //x=46.355 \
 //y=5.155 //x2=46.25 //y2=2.08
cc_3604 ( N_noxref_13_c_4448_n N_SN_c_6891_n ) capacitor c=0.00265761f \
 //x=48.1 //y=2.59 //x2=46.25 //y2=2.08
cc_3605 ( N_noxref_13_c_4435_n N_SN_c_6892_n ) capacitor c=0.0216476f \
 //x=74.995 //y=2.96 //x2=59.2 //y2=2.08
cc_3606 ( N_noxref_13_c_4435_n N_SN_c_6893_n ) capacitor c=0.0216476f \
 //x=74.995 //y=2.96 //x2=70.67 //y2=2.08
cc_3607 ( N_noxref_13_c_4464_n N_SN_M108_noxref_g ) capacitor c=0.0165266f \
 //x=46.355 //y=5.155 //x2=46.22 //y2=6.02
cc_3608 ( N_noxref_13_M108_noxref_d N_SN_M108_noxref_g ) capacitor \
 c=0.0180032f //x=46.295 //y=5.02 //x2=46.22 //y2=6.02
cc_3609 ( N_noxref_13_c_4470_n N_SN_M109_noxref_g ) capacitor c=0.01736f \
 //x=47.235 //y=5.155 //x2=46.66 //y2=6.02
cc_3610 ( N_noxref_13_M108_noxref_d N_SN_M109_noxref_g ) capacitor \
 c=0.0180032f //x=46.295 //y=5.02 //x2=46.66 //y2=6.02
cc_3611 ( N_noxref_13_c_4671_p N_SN_c_7179_n ) capacitor c=0.00426767f \
 //x=46.44 //y=5.155 //x2=46.585 //y2=4.79
cc_3612 ( N_noxref_13_c_4435_n N_SN_c_7204_n ) capacitor c=4.10467e-19 \
 //x=74.995 //y=2.96 //x2=70.76 //y2=1.915
cc_3613 ( N_noxref_13_c_4464_n N_SN_c_7133_n ) capacitor c=0.00322054f \
 //x=46.355 //y=5.155 //x2=46.25 //y2=4.7
cc_3614 ( N_noxref_13_c_4435_n N_noxref_21_c_7696_n ) capacitor c=0.0358131f \
 //x=74.995 //y=2.96 //x2=60.195 //y2=3.7
cc_3615 ( N_noxref_13_c_4435_n N_noxref_21_c_7697_n ) capacitor c=8.32553e-19 \
 //x=74.995 //y=2.96 //x2=55.615 //y2=3.7
cc_3616 ( N_noxref_13_c_4435_n N_noxref_21_c_7698_n ) capacitor c=0.0288894f \
 //x=74.995 //y=2.96 //x2=64.265 //y2=3.7
cc_3617 ( N_noxref_13_c_4435_n N_noxref_21_c_7699_n ) capacitor c=6.03896e-19 \
 //x=74.995 //y=2.96 //x2=60.425 //y2=3.7
cc_3618 ( N_noxref_13_c_4435_n N_noxref_21_c_7656_n ) capacitor c=0.0545501f \
 //x=74.995 //y=2.96 //x2=71.665 //y2=3.7
cc_3619 ( N_noxref_13_c_4435_n N_noxref_21_c_7701_n ) capacitor c=5.76918e-19 \
 //x=74.995 //y=2.96 //x2=64.495 //y2=3.7
cc_3620 ( N_noxref_13_c_4435_n N_noxref_21_c_7648_n ) capacitor c=0.0179917f \
 //x=74.995 //y=2.96 //x2=55.5 //y2=2.08
cc_3621 ( N_noxref_13_c_4435_n N_noxref_21_c_7649_n ) capacitor c=0.0202855f \
 //x=74.995 //y=2.96 //x2=60.31 //y2=2.08
cc_3622 ( N_noxref_13_c_4435_n N_noxref_21_c_7651_n ) capacitor c=0.021075f \
 //x=74.995 //y=2.96 //x2=64.38 //y2=3.7
cc_3623 ( N_noxref_13_c_4435_n N_noxref_21_c_7652_n ) capacitor c=0.022447f \
 //x=74.995 //y=2.96 //x2=71.78 //y2=2.08
cc_3624 ( N_noxref_13_c_4435_n N_noxref_21_c_7706_n ) capacitor c=0.0018311f \
 //x=74.995 //y=2.96 //x2=71.78 //y2=2.08
cc_3625 ( N_noxref_13_c_4444_n N_noxref_22_c_7969_n ) capacitor c=0.00923886f \
 //x=81.655 //y=4.07 //x2=77.255 //y2=5.21
cc_3626 ( N_noxref_13_M145_noxref_g N_noxref_22_c_7969_n ) capacitor \
 c=0.0104371f //x=75.59 //y=6.025 //x2=77.255 //y2=5.21
cc_3627 ( N_noxref_13_c_4444_n N_noxref_22_c_7975_n ) capacitor c=0.00122833f \
 //x=81.655 //y=4.07 //x2=75.485 //y2=5.21
cc_3628 ( N_noxref_13_M144_noxref_g N_noxref_22_c_7975_n ) capacitor \
 c=0.0010118f //x=75.15 //y=6.025 //x2=75.485 //y2=5.21
cc_3629 ( N_noxref_13_M145_noxref_g N_noxref_22_c_7975_n ) capacitor \
 c=8.30848e-19 //x=75.59 //y=6.025 //x2=75.485 //y2=5.21
cc_3630 ( N_noxref_13_c_4479_n N_noxref_22_c_7980_n ) capacitor c=0.012748f \
 //x=75.11 //y=4.54 //x2=75.285 //y2=5.21
cc_3631 ( N_noxref_13_M144_noxref_g N_noxref_22_c_7980_n ) capacitor \
 c=0.0161605f //x=75.15 //y=6.025 //x2=75.285 //y2=5.21
cc_3632 ( N_noxref_13_c_4497_n N_noxref_22_c_7980_n ) capacitor c=0.00307538f \
 //x=75.15 //y=4.705 //x2=75.285 //y2=5.21
cc_3633 ( N_noxref_13_M144_noxref_g N_noxref_22_c_7986_n ) capacitor \
 c=0.00226657f //x=75.15 //y=6.025 //x2=75.37 //y2=5.295
cc_3634 ( N_noxref_13_M145_noxref_g N_noxref_22_c_7986_n ) capacitor \
 c=0.0197448f //x=75.59 //y=6.025 //x2=75.37 //y2=5.295
cc_3635 ( N_noxref_13_c_4496_n N_noxref_22_c_7986_n ) capacitor c=0.00458101f \
 //x=75.515 //y=4.795 //x2=75.37 //y2=5.295
cc_3636 ( N_noxref_13_M144_noxref_g N_noxref_22_M144_noxref_d ) capacitor \
 c=0.016914f //x=75.15 //y=6.025 //x2=75.225 //y2=5.025
cc_3637 ( N_noxref_13_c_4435_n N_noxref_23_c_8089_n ) capacitor c=0.00331464f \
 //x=74.995 //y=2.96 //x2=72.405 //y2=4.44
cc_3638 ( N_noxref_13_c_4435_n N_noxref_23_c_8093_n ) capacitor c=0.00429139f \
 //x=74.995 //y=2.96 //x2=73.885 //y2=4.44
cc_3639 ( N_noxref_13_c_4435_n N_noxref_23_c_8097_n ) capacitor c=2.96875e-19 \
 //x=74.995 //y=2.96 //x2=72.635 //y2=4.44
cc_3640 ( N_noxref_13_c_4435_n N_noxref_23_c_8100_n ) capacitor c=0.00512306f \
 //x=74.995 //y=2.96 //x2=77.585 //y2=4.44
cc_3641 ( N_noxref_13_c_4444_n N_noxref_23_c_8100_n ) capacitor c=0.23799f \
 //x=81.655 //y=4.07 //x2=77.585 //y2=4.44
cc_3642 ( N_noxref_13_c_4461_n N_noxref_23_c_8100_n ) capacitor c=0.0289488f \
 //x=75.225 //y=4.07 //x2=77.585 //y2=4.44
cc_3643 ( N_noxref_13_c_4479_n N_noxref_23_c_8100_n ) capacitor c=0.00210648f \
 //x=75.11 //y=4.54 //x2=77.585 //y2=4.44
cc_3644 ( N_noxref_13_c_4449_n N_noxref_23_c_8100_n ) capacitor c=0.0232321f \
 //x=75.11 //y=2.08 //x2=77.585 //y2=4.44
cc_3645 ( N_noxref_13_c_4496_n N_noxref_23_c_8100_n ) capacitor c=0.0069773f \
 //x=75.515 //y=4.795 //x2=77.585 //y2=4.44
cc_3646 ( N_noxref_13_c_4497_n N_noxref_23_c_8100_n ) capacitor c=0.0014023f \
 //x=75.15 //y=4.705 //x2=77.585 //y2=4.44
cc_3647 ( N_noxref_13_c_4435_n N_noxref_23_c_8105_n ) capacitor c=3.35648e-19 \
 //x=74.995 //y=2.96 //x2=74.115 //y2=4.44
cc_3648 ( N_noxref_13_c_4449_n N_noxref_23_c_8105_n ) capacitor c=9.10428e-19 \
 //x=75.11 //y=2.08 //x2=74.115 //y2=4.44
cc_3649 ( N_noxref_13_c_4435_n N_noxref_23_c_8060_n ) capacitor c=0.0192451f \
 //x=74.995 //y=2.96 //x2=66.97 //y2=2.08
cc_3650 ( N_noxref_13_c_4435_n N_noxref_23_c_8177_n ) capacitor c=0.00838703f \
 //x=74.995 //y=2.96 //x2=72.12 //y2=1.665
cc_3651 ( N_noxref_13_c_4435_n N_noxref_23_c_8126_n ) capacitor c=0.0235599f \
 //x=74.995 //y=2.96 //x2=72.52 //y2=4.44
cc_3652 ( N_noxref_13_c_4449_n N_noxref_23_c_8126_n ) capacitor c=7.65096e-19 \
 //x=75.11 //y=2.08 //x2=72.52 //y2=4.44
cc_3653 ( N_noxref_13_c_4435_n N_noxref_23_c_8063_n ) capacitor c=0.0252848f \
 //x=74.995 //y=2.96 //x2=74 //y2=2.08
cc_3654 ( N_noxref_13_c_4461_n N_noxref_23_c_8063_n ) capacitor c=0.00526349f \
 //x=75.225 //y=4.07 //x2=74 //y2=2.08
cc_3655 ( N_noxref_13_c_4479_n N_noxref_23_c_8063_n ) capacitor c=0.00227044f \
 //x=75.11 //y=4.54 //x2=74 //y2=2.08
cc_3656 ( N_noxref_13_c_4449_n N_noxref_23_c_8063_n ) capacitor c=0.0465433f \
 //x=75.11 //y=2.08 //x2=74 //y2=2.08
cc_3657 ( N_noxref_13_c_4453_n N_noxref_23_c_8063_n ) capacitor c=0.00224607f \
 //x=75.11 //y=2.08 //x2=74 //y2=2.08
cc_3658 ( N_noxref_13_c_4497_n N_noxref_23_c_8063_n ) capacitor c=0.00228787f \
 //x=75.15 //y=4.705 //x2=74 //y2=2.08
cc_3659 ( N_noxref_13_c_4435_n N_noxref_23_c_8066_n ) capacitor c=0.00144897f \
 //x=74.995 //y=2.96 //x2=77.7 //y2=2.08
cc_3660 ( N_noxref_13_c_4444_n N_noxref_23_c_8066_n ) capacitor c=0.0242848f \
 //x=81.655 //y=4.07 //x2=77.7 //y2=2.08
cc_3661 ( N_noxref_13_c_4449_n N_noxref_23_c_8066_n ) capacitor c=0.00873163f \
 //x=75.11 //y=2.08 //x2=77.7 //y2=2.08
cc_3662 ( N_noxref_13_M144_noxref_g N_noxref_23_M142_noxref_g ) capacitor \
 c=0.010584f //x=75.15 //y=6.025 //x2=74.27 //y2=6.025
cc_3663 ( N_noxref_13_M144_noxref_g N_noxref_23_M143_noxref_g ) capacitor \
 c=0.106414f //x=75.15 //y=6.025 //x2=74.71 //y2=6.025
cc_3664 ( N_noxref_13_M145_noxref_g N_noxref_23_M143_noxref_g ) capacitor \
 c=0.0102479f //x=75.59 //y=6.025 //x2=74.71 //y2=6.025
cc_3665 ( N_noxref_13_c_4725_p N_noxref_23_c_8068_n ) capacitor c=4.86506e-19 \
 //x=75.145 //y=0.905 //x2=74.175 //y2=0.865
cc_3666 ( N_noxref_13_c_4725_p N_noxref_23_c_8070_n ) capacitor c=0.00152104f \
 //x=75.145 //y=0.905 //x2=74.175 //y2=1.21
cc_3667 ( N_noxref_13_c_4727_p N_noxref_23_c_8071_n ) capacitor c=0.00109982f \
 //x=75.145 //y=1.25 //x2=74.175 //y2=1.52
cc_3668 ( N_noxref_13_c_4728_p N_noxref_23_c_8071_n ) capacitor c=0.00179029f \
 //x=75.145 //y=1.56 //x2=74.175 //y2=1.52
cc_3669 ( N_noxref_13_c_4728_p N_noxref_23_c_8072_n ) capacitor c=0.00662747f \
 //x=75.145 //y=1.56 //x2=74.175 //y2=1.915
cc_3670 ( N_noxref_13_c_4479_n N_noxref_23_c_8197_n ) capacitor c=0.00155256f \
 //x=75.11 //y=4.54 //x2=74.635 //y2=4.795
cc_3671 ( N_noxref_13_c_4497_n N_noxref_23_c_8197_n ) capacitor c=0.0201611f \
 //x=75.15 //y=4.705 //x2=74.635 //y2=4.795
cc_3672 ( N_noxref_13_c_4479_n N_noxref_23_c_8146_n ) capacitor c=0.00180548f \
 //x=75.11 //y=4.54 //x2=74.345 //y2=4.795
cc_3673 ( N_noxref_13_c_4497_n N_noxref_23_c_8146_n ) capacitor c=0.00447195f \
 //x=75.15 //y=4.705 //x2=74.345 //y2=4.795
cc_3674 ( N_noxref_13_c_4725_p N_noxref_23_c_8075_n ) capacitor c=0.0151475f \
 //x=75.145 //y=0.905 //x2=74.705 //y2=0.865
cc_3675 ( N_noxref_13_c_4735_p N_noxref_23_c_8075_n ) capacitor c=0.00124846f \
 //x=75.675 //y=0.905 //x2=74.705 //y2=0.865
cc_3676 ( N_noxref_13_c_4727_p N_noxref_23_c_8077_n ) capacitor c=0.0111064f \
 //x=75.145 //y=1.25 //x2=74.705 //y2=1.21
cc_3677 ( N_noxref_13_c_4728_p N_noxref_23_c_8077_n ) capacitor c=0.00862358f \
 //x=75.145 //y=1.56 //x2=74.705 //y2=1.21
cc_3678 ( N_noxref_13_c_4738_p N_noxref_23_c_8077_n ) capacitor c=0.00168739f \
 //x=75.675 //y=1.25 //x2=74.705 //y2=1.21
cc_3679 ( N_noxref_13_c_4435_n N_noxref_23_c_8087_n ) capacitor c=0.00384973f \
 //x=74.995 //y=2.96 //x2=74 //y2=2.08
cc_3680 ( N_noxref_13_c_4449_n N_noxref_23_c_8087_n ) capacitor c=0.00236728f \
 //x=75.11 //y=2.08 //x2=74 //y2=2.08
cc_3681 ( N_noxref_13_c_4453_n N_noxref_23_c_8087_n ) capacitor c=0.00942627f \
 //x=75.11 //y=2.08 //x2=74 //y2=2.08
cc_3682 ( N_noxref_13_c_4444_n N_noxref_23_c_8148_n ) capacitor c=0.00381677f \
 //x=81.655 //y=4.07 //x2=77.7 //y2=4.705
cc_3683 ( N_noxref_13_c_4455_n N_noxref_24_c_8424_n ) capacitor c=0.0693978f \
 //x=47.985 //y=4.07 //x2=79.065 //y2=3.33
cc_3684 ( N_noxref_13_c_4513_n N_noxref_24_c_8424_n ) capacitor c=8.35979e-19 \
 //x=42.665 //y=4.07 //x2=79.065 //y2=3.33
cc_3685 ( N_noxref_13_c_4433_n N_noxref_24_c_8424_n ) capacitor c=0.0340399f \
 //x=50.605 //y=2.59 //x2=79.065 //y2=3.33
cc_3686 ( N_noxref_13_c_4434_n N_noxref_24_c_8424_n ) capacitor c=8.87672e-19 \
 //x=48.215 //y=2.59 //x2=79.065 //y2=3.33
cc_3687 ( N_noxref_13_c_4435_n N_noxref_24_c_8424_n ) capacitor c=0.0292175f \
 //x=74.995 //y=2.96 //x2=79.065 //y2=3.33
cc_3688 ( N_noxref_13_c_4603_p N_noxref_24_c_8424_n ) capacitor c=2.14003f \
 //x=50.775 //y=2.96 //x2=79.065 //y2=3.33
cc_3689 ( N_noxref_13_c_4444_n N_noxref_24_c_8424_n ) capacitor c=0.185533f \
 //x=81.655 //y=4.07 //x2=79.065 //y2=3.33
cc_3690 ( N_noxref_13_c_4461_n N_noxref_24_c_8424_n ) capacitor c=0.01357f \
 //x=75.225 //y=4.07 //x2=79.065 //y2=3.33
cc_3691 ( N_noxref_13_c_4445_n N_noxref_24_c_8424_n ) capacitor c=0.0169786f \
 //x=42.55 //y=2.08 //x2=79.065 //y2=3.33
cc_3692 ( N_noxref_13_c_4448_n N_noxref_24_c_8424_n ) capacitor c=0.0214009f \
 //x=48.1 //y=2.59 //x2=79.065 //y2=3.33
cc_3693 ( N_noxref_13_c_4449_n N_noxref_24_c_8424_n ) capacitor c=0.0244276f \
 //x=75.11 //y=2.08 //x2=79.065 //y2=3.33
cc_3694 ( N_noxref_13_c_4444_n N_noxref_24_c_8426_n ) capacitor c=0.0234271f \
 //x=81.655 //y=4.07 //x2=80.545 //y2=2.08
cc_3695 ( N_noxref_13_c_4451_n N_noxref_24_c_8426_n ) capacitor c=0.00668632f \
 //x=81.77 //y=2.08 //x2=80.545 //y2=2.08
cc_3696 ( N_noxref_13_c_4756_p N_noxref_24_c_8426_n ) capacitor c=0.00319611f \
 //x=81.77 //y=2.08 //x2=80.545 //y2=2.08
cc_3697 ( N_noxref_13_c_4444_n N_noxref_24_c_8431_n ) capacitor c=0.0248463f \
 //x=81.655 //y=4.07 //x2=79.18 //y2=2.08
cc_3698 ( N_noxref_13_c_4451_n N_noxref_24_c_8431_n ) capacitor c=7.56813e-19 \
 //x=81.77 //y=2.08 //x2=79.18 //y2=2.08
cc_3699 ( N_noxref_13_c_4444_n N_noxref_24_c_8433_n ) capacitor c=0.0282853f \
 //x=81.655 //y=4.07 //x2=80.66 //y2=2.08
cc_3700 ( N_noxref_13_c_4451_n N_noxref_24_c_8433_n ) capacitor c=0.0538261f \
 //x=81.77 //y=2.08 //x2=80.66 //y2=2.08
cc_3701 ( N_noxref_13_c_4756_p N_noxref_24_c_8433_n ) capacitor c=0.00207994f \
 //x=81.77 //y=2.08 //x2=80.66 //y2=2.08
cc_3702 ( N_noxref_13_c_4762_p N_noxref_24_c_8433_n ) capacitor c=0.00196222f \
 //x=81.79 //y=4.705 //x2=80.66 //y2=2.08
cc_3703 ( N_noxref_13_M152_noxref_g N_noxref_24_M150_noxref_g ) capacitor \
 c=0.00932631f //x=81.81 //y=6.025 //x2=80.93 //y2=6.025
cc_3704 ( N_noxref_13_M152_noxref_g N_noxref_24_M151_noxref_g ) capacitor \
 c=0.110179f //x=81.81 //y=6.025 //x2=81.37 //y2=6.025
cc_3705 ( N_noxref_13_M153_noxref_g N_noxref_24_M151_noxref_g ) capacitor \
 c=0.00876656f //x=82.25 //y=6.025 //x2=81.37 //y2=6.025
cc_3706 ( N_noxref_13_c_4444_n N_noxref_24_c_8640_n ) capacitor c=0.00791694f \
 //x=81.655 //y=4.07 //x2=78.545 //y2=4.795
cc_3707 ( N_noxref_13_c_4444_n N_noxref_24_c_8480_n ) capacitor c=0.0014567f \
 //x=81.655 //y=4.07 //x2=78.91 //y2=4.87
cc_3708 ( N_noxref_13_c_4768_p N_noxref_24_c_8435_n ) capacitor c=4.86506e-19 \
 //x=81.805 //y=0.905 //x2=80.835 //y2=0.865
cc_3709 ( N_noxref_13_c_4768_p N_noxref_24_c_8437_n ) capacitor c=0.00101233f \
 //x=81.805 //y=0.905 //x2=80.835 //y2=1.21
cc_3710 ( N_noxref_13_c_4770_p N_noxref_24_c_8644_n ) capacitor c=0.00257836f \
 //x=81.805 //y=1.56 //x2=80.835 //y2=1.52
cc_3711 ( N_noxref_13_c_4770_p N_noxref_24_c_8438_n ) capacitor c=0.00662747f \
 //x=81.805 //y=1.56 //x2=80.835 //y2=1.915
cc_3712 ( N_noxref_13_c_4772_p N_noxref_24_c_8646_n ) capacitor c=0.00168516f \
 //x=81.79 //y=4.705 //x2=81.295 //y2=4.795
cc_3713 ( N_noxref_13_c_4762_p N_noxref_24_c_8646_n ) capacitor c=0.0225854f \
 //x=81.79 //y=4.705 //x2=81.295 //y2=4.795
cc_3714 ( N_noxref_13_c_4444_n N_noxref_24_c_8481_n ) capacitor c=0.0117386f \
 //x=81.655 //y=4.07 //x2=81.005 //y2=4.795
cc_3715 ( N_noxref_13_c_4772_p N_noxref_24_c_8481_n ) capacitor c=0.00143876f \
 //x=81.79 //y=4.705 //x2=81.005 //y2=4.795
cc_3716 ( N_noxref_13_c_4762_p N_noxref_24_c_8481_n ) capacitor c=0.00469886f \
 //x=81.79 //y=4.705 //x2=81.005 //y2=4.795
cc_3717 ( N_noxref_13_c_4768_p N_noxref_24_c_8441_n ) capacitor c=0.0161138f \
 //x=81.805 //y=0.905 //x2=81.365 //y2=0.865
cc_3718 ( N_noxref_13_c_4778_p N_noxref_24_c_8441_n ) capacitor c=0.00130607f \
 //x=82.335 //y=0.905 //x2=81.365 //y2=0.865
cc_3719 ( N_noxref_13_c_4779_p N_noxref_24_c_8443_n ) capacitor c=0.0120728f \
 //x=81.805 //y=1.255 //x2=81.365 //y2=1.21
cc_3720 ( N_noxref_13_c_4770_p N_noxref_24_c_8443_n ) capacitor c=0.00862358f \
 //x=81.805 //y=1.56 //x2=81.365 //y2=1.21
cc_3721 ( N_noxref_13_c_4781_p N_noxref_24_c_8443_n ) capacitor c=4.4593e-19 \
 //x=82.18 //y=1.405 //x2=81.365 //y2=1.21
cc_3722 ( N_noxref_13_c_4782_p N_noxref_24_c_8443_n ) capacitor c=0.00111855f \
 //x=82.335 //y=1.255 //x2=81.365 //y2=1.21
cc_3723 ( N_noxref_13_c_4451_n N_noxref_24_c_8444_n ) capacitor c=0.00218919f \
 //x=81.77 //y=2.08 //x2=80.66 //y2=2.08
cc_3724 ( N_noxref_13_c_4756_p N_noxref_24_c_8444_n ) capacitor c=0.00908973f \
 //x=81.77 //y=2.08 //x2=80.66 //y2=2.08
cc_3725 ( N_noxref_13_c_4444_n N_noxref_25_c_8898_n ) capacitor c=0.0535575f \
 //x=81.655 //y=4.07 //x2=80.595 //y2=5.21
cc_3726 ( N_noxref_13_c_4444_n N_noxref_25_c_8902_n ) capacitor c=0.008149f \
 //x=81.655 //y=4.07 //x2=78.805 //y2=5.21
cc_3727 ( N_noxref_13_c_4444_n N_noxref_25_c_8916_n ) capacitor c=3.2507e-19 \
 //x=81.655 //y=4.07 //x2=78.605 //y2=5.21
cc_3728 ( N_noxref_13_c_4444_n N_noxref_25_c_8904_n ) capacitor c=0.0181202f \
 //x=81.655 //y=4.07 //x2=77.895 //y2=5.21
cc_3729 ( N_noxref_13_c_4444_n N_noxref_25_c_8905_n ) capacitor c=0.00337443f \
 //x=81.655 //y=4.07 //x2=78.69 //y2=5.295
cc_3730 ( N_noxref_13_c_4444_n N_noxref_25_c_8906_n ) capacitor c=0.0011253f \
 //x=81.655 //y=4.07 //x2=80.71 //y2=5.21
cc_3731 ( N_noxref_13_c_4444_n N_noxref_25_c_8920_n ) capacitor c=0.00358031f \
 //x=81.655 //y=4.07 //x2=81.505 //y2=6.91
cc_3732 ( N_noxref_13_M152_noxref_g N_noxref_25_c_8921_n ) capacitor \
 c=0.0150104f //x=81.81 //y=6.025 //x2=82.385 //y2=6.91
cc_3733 ( N_noxref_13_M153_noxref_g N_noxref_25_c_8921_n ) capacitor \
 c=0.0163361f //x=82.25 //y=6.025 //x2=82.385 //y2=6.91
cc_3734 ( N_noxref_13_M152_noxref_g N_noxref_25_M151_noxref_d ) capacitor \
 c=0.0130327f //x=81.81 //y=6.025 //x2=81.445 //y2=5.025
cc_3735 ( N_noxref_13_M153_noxref_g N_noxref_25_M153_noxref_d ) capacitor \
 c=0.0351101f //x=82.25 //y=6.025 //x2=82.325 //y2=5.025
cc_3736 ( N_noxref_13_c_4444_n N_noxref_26_c_8988_n ) capacitor c=0.00477352f \
 //x=81.655 //y=4.07 //x2=78.625 //y2=1.18
cc_3737 ( N_noxref_13_c_4735_p N_noxref_26_c_8988_n ) capacitor c=4.67724e-19 \
 //x=75.675 //y=0.905 //x2=78.625 //y2=1.18
cc_3738 ( N_noxref_13_c_4738_p N_noxref_26_c_8988_n ) capacitor c=0.00747449f \
 //x=75.675 //y=1.25 //x2=78.625 //y2=1.18
cc_3739 ( N_noxref_13_c_4444_n N_noxref_26_c_8995_n ) capacitor c=5.91174e-19 \
 //x=81.655 //y=4.07 //x2=75.525 //y2=1.18
cc_3740 ( N_noxref_13_c_4725_p N_noxref_26_c_8995_n ) capacitor c=3.66947e-19 \
 //x=75.145 //y=0.905 //x2=75.525 //y2=1.18
cc_3741 ( N_noxref_13_c_4727_p N_noxref_26_c_8995_n ) capacitor c=0.00353233f \
 //x=75.145 //y=1.25 //x2=75.525 //y2=1.18
cc_3742 ( N_noxref_13_c_4728_p N_noxref_26_c_8995_n ) capacitor c=0.00292382f \
 //x=75.145 //y=1.56 //x2=75.525 //y2=1.18
cc_3743 ( N_noxref_13_c_4803_p N_noxref_26_c_8995_n ) capacitor c=4.06815e-19 \
 //x=75.52 //y=0.75 //x2=75.525 //y2=1.18
cc_3744 ( N_noxref_13_c_4804_p N_noxref_26_c_8995_n ) capacitor c=7.90416e-19 \
 //x=75.52 //y=1.405 //x2=75.525 //y2=1.18
cc_3745 ( N_noxref_13_c_4738_p N_noxref_26_c_8995_n ) capacitor c=0.0013439f \
 //x=75.675 //y=1.25 //x2=75.525 //y2=1.18
cc_3746 ( N_noxref_13_c_4444_n N_noxref_26_c_8996_n ) capacitor c=0.0114358f \
 //x=81.655 //y=4.07 //x2=81.955 //y2=1.18
cc_3747 ( N_noxref_13_c_4451_n N_noxref_26_c_8996_n ) capacitor c=0.00449159f \
 //x=81.77 //y=2.08 //x2=81.955 //y2=1.18
cc_3748 ( N_noxref_13_c_4768_p N_noxref_26_c_8996_n ) capacitor c=6.33948e-19 \
 //x=81.805 //y=0.905 //x2=81.955 //y2=1.18
cc_3749 ( N_noxref_13_c_4779_p N_noxref_26_c_8996_n ) capacitor c=0.0043333f \
 //x=81.805 //y=1.255 //x2=81.955 //y2=1.18
cc_3750 ( N_noxref_13_c_4770_p N_noxref_26_c_8996_n ) capacitor c=0.0040799f \
 //x=81.805 //y=1.56 //x2=81.955 //y2=1.18
cc_3751 ( N_noxref_13_c_4811_p N_noxref_26_c_8996_n ) capacitor c=4.52813e-19 \
 //x=82.18 //y=0.75 //x2=81.955 //y2=1.18
cc_3752 ( N_noxref_13_c_4781_p N_noxref_26_c_8996_n ) capacitor c=0.00296491f \
 //x=82.18 //y=1.405 //x2=81.955 //y2=1.18
cc_3753 ( N_noxref_13_c_4778_p N_noxref_26_c_8996_n ) capacitor c=2.65983e-19 \
 //x=82.335 //y=0.905 //x2=81.955 //y2=1.18
cc_3754 ( N_noxref_13_c_4782_p N_noxref_26_c_8996_n ) capacitor c=0.00362989f \
 //x=82.335 //y=1.255 //x2=81.955 //y2=1.18
cc_3755 ( N_noxref_13_c_4756_p N_noxref_26_c_8996_n ) capacitor c=5.89141e-19 \
 //x=81.77 //y=2.08 //x2=81.955 //y2=1.18
cc_3756 ( N_noxref_13_c_4444_n N_noxref_26_c_9003_n ) capacitor c=5.35864e-19 \
 //x=81.655 //y=4.07 //x2=78.855 //y2=1.18
cc_3757 ( N_noxref_13_c_4444_n N_noxref_26_c_9007_n ) capacitor c=0.0243956f \
 //x=81.655 //y=4.07 //x2=82.625 //y2=4.07
cc_3758 ( N_noxref_13_c_4451_n N_noxref_26_c_9007_n ) capacitor c=0.00197285f \
 //x=81.77 //y=2.08 //x2=82.625 //y2=4.07
cc_3759 ( N_noxref_13_c_4444_n N_noxref_26_c_9089_n ) capacitor c=0.00154966f \
 //x=81.655 //y=4.07 //x2=81.945 //y2=5.21
cc_3760 ( N_noxref_13_c_4772_p N_noxref_26_c_9089_n ) capacitor c=0.0128151f \
 //x=81.79 //y=4.705 //x2=81.945 //y2=5.21
cc_3761 ( N_noxref_13_M152_noxref_g N_noxref_26_c_9089_n ) capacitor \
 c=0.0167296f //x=81.81 //y=6.025 //x2=81.945 //y2=5.21
cc_3762 ( N_noxref_13_c_4762_p N_noxref_26_c_9089_n ) capacitor c=0.00368327f \
 //x=81.79 //y=4.705 //x2=81.945 //y2=5.21
cc_3763 ( N_noxref_13_c_4444_n N_noxref_26_c_9045_n ) capacitor c=0.0138451f \
 //x=81.655 //y=4.07 //x2=81.235 //y2=5.21
cc_3764 ( N_noxref_13_M153_noxref_g N_noxref_26_c_9046_n ) capacitor \
 c=0.0222938f //x=82.25 //y=6.025 //x2=82.425 //y2=5.21
cc_3765 ( N_noxref_13_c_4781_p N_noxref_26_c_9008_n ) capacitor c=0.00810194f \
 //x=82.18 //y=1.405 //x2=82.425 //y2=1.645
cc_3766 ( N_noxref_13_c_4826_p N_noxref_26_c_9096_n ) capacitor c=0.00671029f \
 //x=81.77 //y=1.915 //x2=82.155 //y2=1.645
cc_3767 ( N_noxref_13_c_4444_n N_noxref_26_c_9010_n ) capacitor c=0.00246068f \
 //x=81.655 //y=4.07 //x2=82.51 //y2=4.07
cc_3768 ( N_noxref_13_c_4451_n N_noxref_26_c_9010_n ) capacitor c=0.0817254f \
 //x=81.77 //y=2.08 //x2=82.51 //y2=4.07
cc_3769 ( N_noxref_13_c_4772_p N_noxref_26_c_9010_n ) capacitor c=0.00998395f \
 //x=81.79 //y=4.705 //x2=82.51 //y2=4.07
cc_3770 ( N_noxref_13_c_4830_p N_noxref_26_c_9010_n ) capacitor c=0.0143966f \
 //x=82.175 //y=4.795 //x2=82.51 //y2=4.07
cc_3771 ( N_noxref_13_c_4756_p N_noxref_26_c_9010_n ) capacitor c=0.00704374f \
 //x=81.77 //y=2.08 //x2=82.51 //y2=4.07
cc_3772 ( N_noxref_13_c_4826_p N_noxref_26_c_9010_n ) capacitor c=0.0033061f \
 //x=81.77 //y=1.915 //x2=82.51 //y2=4.07
cc_3773 ( N_noxref_13_c_4762_p N_noxref_26_c_9010_n ) capacitor c=0.00526987f \
 //x=81.79 //y=4.705 //x2=82.51 //y2=4.07
cc_3774 ( N_noxref_13_c_4451_n N_noxref_26_c_9011_n ) capacitor c=9.6769e-19 \
 //x=81.77 //y=2.08 //x2=83.99 //y2=2.085
cc_3775 ( N_noxref_13_c_4830_p N_noxref_26_c_9105_n ) capacitor c=0.00410596f \
 //x=82.175 //y=4.795 //x2=82.03 //y2=5.21
cc_3776 ( N_noxref_13_c_4725_p N_noxref_26_M46_noxref_d ) capacitor \
 c=0.00218556f //x=75.145 //y=0.905 //x2=75.22 //y2=0.905
cc_3777 ( N_noxref_13_c_4727_p N_noxref_26_M46_noxref_d ) capacitor \
 c=0.00327871f //x=75.145 //y=1.25 //x2=75.22 //y2=0.905
cc_3778 ( N_noxref_13_c_4728_p N_noxref_26_M46_noxref_d ) capacitor \
 c=0.00292542f //x=75.145 //y=1.56 //x2=75.22 //y2=0.905
cc_3779 ( N_noxref_13_c_4803_p N_noxref_26_M46_noxref_d ) capacitor \
 c=0.00235569f //x=75.52 //y=0.75 //x2=75.22 //y2=0.905
cc_3780 ( N_noxref_13_c_4804_p N_noxref_26_M46_noxref_d ) capacitor \
 c=0.00613695f //x=75.52 //y=1.405 //x2=75.22 //y2=0.905
cc_3781 ( N_noxref_13_c_4735_p N_noxref_26_M46_noxref_d ) capacitor \
 c=0.00131413f //x=75.675 //y=0.905 //x2=75.22 //y2=0.905
cc_3782 ( N_noxref_13_c_4738_p N_noxref_26_M46_noxref_d ) capacitor \
 c=0.00676348f //x=75.675 //y=1.25 //x2=75.22 //y2=0.905
cc_3783 ( N_noxref_13_c_4768_p N_noxref_26_M50_noxref_d ) capacitor \
 c=0.00226395f //x=81.805 //y=0.905 //x2=81.88 //y2=0.905
cc_3784 ( N_noxref_13_c_4779_p N_noxref_26_M50_noxref_d ) capacitor \
 c=0.004517f //x=81.805 //y=1.255 //x2=81.88 //y2=0.905
cc_3785 ( N_noxref_13_c_4770_p N_noxref_26_M50_noxref_d ) capacitor \
 c=0.00655125f //x=81.805 //y=1.56 //x2=81.88 //y2=0.905
cc_3786 ( N_noxref_13_c_4811_p N_noxref_26_M50_noxref_d ) capacitor \
 c=0.00241003f //x=82.18 //y=0.75 //x2=81.88 //y2=0.905
cc_3787 ( N_noxref_13_c_4781_p N_noxref_26_M50_noxref_d ) capacitor \
 c=0.0159024f //x=82.18 //y=1.405 //x2=81.88 //y2=0.905
cc_3788 ( N_noxref_13_c_4778_p N_noxref_26_M50_noxref_d ) capacitor \
 c=0.00132831f //x=82.335 //y=0.905 //x2=81.88 //y2=0.905
cc_3789 ( N_noxref_13_c_4782_p N_noxref_26_M50_noxref_d ) capacitor \
 c=0.00330743f //x=82.335 //y=1.255 //x2=81.88 //y2=0.905
cc_3790 ( N_noxref_13_M152_noxref_g N_noxref_26_M152_noxref_d ) capacitor \
 c=0.0130327f //x=81.81 //y=6.025 //x2=81.885 //y2=5.025
cc_3791 ( N_noxref_13_M153_noxref_g N_noxref_26_M152_noxref_d ) capacitor \
 c=0.0136385f //x=82.25 //y=6.025 //x2=81.885 //y2=5.025
cc_3792 ( N_noxref_13_c_4528_n N_noxref_42_c_10006_n ) capacitor c=0.00623646f \
 //x=42.585 //y=1.56 //x2=42.365 //y2=1.495
cc_3793 ( N_noxref_13_c_4533_n N_noxref_42_c_10006_n ) capacitor c=0.00173579f \
 //x=42.55 //y=2.08 //x2=42.365 //y2=1.495
cc_3794 ( N_noxref_13_c_4445_n N_noxref_42_c_10007_n ) capacitor c=0.00156605f \
 //x=42.55 //y=2.08 //x2=43.25 //y2=0.53
cc_3795 ( N_noxref_13_c_4523_n N_noxref_42_c_10007_n ) capacitor c=0.0188655f \
 //x=42.585 //y=0.905 //x2=43.25 //y2=0.53
cc_3796 ( N_noxref_13_c_4531_n N_noxref_42_c_10007_n ) capacitor c=0.00656458f \
 //x=43.115 //y=0.905 //x2=43.25 //y2=0.53
cc_3797 ( N_noxref_13_c_4533_n N_noxref_42_c_10007_n ) capacitor c=2.1838e-19 \
 //x=42.55 //y=2.08 //x2=43.25 //y2=0.53
cc_3798 ( N_noxref_13_c_4523_n N_noxref_42_M25_noxref_s ) capacitor \
 c=0.00623646f //x=42.585 //y=0.905 //x2=41.26 //y2=0.365
cc_3799 ( N_noxref_13_c_4531_n N_noxref_42_M25_noxref_s ) capacitor \
 c=0.0143002f //x=43.115 //y=0.905 //x2=41.26 //y2=0.365
cc_3800 ( N_noxref_13_c_4532_n N_noxref_42_M25_noxref_s ) capacitor \
 c=0.00290153f //x=43.115 //y=1.25 //x2=41.26 //y2=0.365
cc_3801 ( N_noxref_13_M29_noxref_d N_noxref_43_M27_noxref_s ) capacitor \
 c=0.00309936f //x=47.425 //y=0.915 //x2=44.485 //y2=0.375
cc_3802 ( N_noxref_13_c_4447_n N_noxref_44_c_10107_n ) capacitor c=0.00457167f \
 //x=48.015 //y=1.665 //x2=48.015 //y2=0.54
cc_3803 ( N_noxref_13_M29_noxref_d N_noxref_44_c_10107_n ) capacitor \
 c=0.0115903f //x=47.425 //y=0.915 //x2=48.015 //y2=0.54
cc_3804 ( N_noxref_13_c_4658_p N_noxref_44_c_10119_n ) capacitor c=0.020048f \
 //x=47.7 //y=1.665 //x2=47.13 //y2=0.995
cc_3805 ( N_noxref_13_M29_noxref_d N_noxref_44_M28_noxref_d ) capacitor \
 c=5.27807e-19 //x=47.425 //y=0.915 //x2=45.89 //y2=0.91
cc_3806 ( N_noxref_13_c_4447_n N_noxref_44_M29_noxref_s ) capacitor \
 c=0.0184051f //x=48.015 //y=1.665 //x2=46.995 //y2=0.375
cc_3807 ( N_noxref_13_M29_noxref_d N_noxref_44_M29_noxref_s ) capacitor \
 c=0.0426444f //x=47.425 //y=0.915 //x2=46.995 //y2=0.375
cc_3808 ( N_noxref_13_c_4447_n N_noxref_45_c_10172_n ) capacitor c=3.04182e-19 \
 //x=48.015 //y=1.665 //x2=49.535 //y2=1.495
cc_3809 ( N_noxref_13_c_4435_n N_noxref_52_c_10527_n ) capacitor c=0.00152987f \
 //x=74.995 //y=2.96 //x2=70.895 //y2=1.59
cc_3810 ( N_noxref_13_c_4435_n N_noxref_52_M42_noxref_s ) capacitor \
 c=0.00302917f //x=74.995 //y=2.96 //x2=68.905 //y2=0.375
cc_3811 ( N_noxref_13_c_4435_n N_noxref_53_c_10563_n ) capacitor c=0.00383675f \
 //x=74.995 //y=2.96 //x2=71.465 //y2=0.995
cc_3812 ( N_noxref_13_c_4435_n N_noxref_53_c_10568_n ) capacitor c=6.69632e-19 \
 //x=74.995 //y=2.96 //x2=72.435 //y2=0.54
cc_3813 ( N_noxref_13_c_4435_n N_noxref_53_M44_noxref_s ) capacitor \
 c=0.00324882f //x=74.995 //y=2.96 //x2=71.415 //y2=0.375
cc_3814 ( N_noxref_13_c_4435_n N_noxref_54_c_10633_n ) capacitor c=8.52215e-19 \
 //x=74.995 //y=2.96 //x2=73.955 //y2=1.495
cc_3815 ( N_noxref_13_c_4435_n N_noxref_54_c_10615_n ) capacitor c=0.0139765f \
 //x=74.995 //y=2.96 //x2=74.84 //y2=1.58
cc_3816 ( N_noxref_13_c_4435_n N_noxref_54_c_10622_n ) capacitor c=0.00323786f \
 //x=74.995 //y=2.96 //x2=74.925 //y2=1.495
cc_3817 ( N_noxref_13_c_4728_p N_noxref_54_c_10622_n ) capacitor c=0.00746306f \
 //x=75.145 //y=1.56 //x2=74.925 //y2=1.495
cc_3818 ( N_noxref_13_c_4453_n N_noxref_54_c_10622_n ) capacitor c=0.00174417f \
 //x=75.11 //y=2.08 //x2=74.925 //y2=1.495
cc_3819 ( N_noxref_13_c_4435_n N_noxref_54_c_10623_n ) capacitor c=4.30845e-19 \
 //x=74.995 //y=2.96 //x2=75.81 //y2=0.53
cc_3820 ( N_noxref_13_c_4449_n N_noxref_54_c_10623_n ) capacitor c=0.00159166f \
 //x=75.11 //y=2.08 //x2=75.81 //y2=0.53
cc_3821 ( N_noxref_13_c_4725_p N_noxref_54_c_10623_n ) capacitor c=0.0200006f \
 //x=75.145 //y=0.905 //x2=75.81 //y2=0.53
cc_3822 ( N_noxref_13_c_4735_p N_noxref_54_c_10623_n ) capacitor c=0.00825432f \
 //x=75.675 //y=0.905 //x2=75.81 //y2=0.53
cc_3823 ( N_noxref_13_c_4453_n N_noxref_54_c_10623_n ) capacitor c=2.1838e-19 \
 //x=75.11 //y=2.08 //x2=75.81 //y2=0.53
cc_3824 ( N_noxref_13_c_4725_p N_noxref_54_M45_noxref_s ) capacitor \
 c=0.00746306f //x=75.145 //y=0.905 //x2=73.82 //y2=0.365
cc_3825 ( N_noxref_13_c_4728_p N_noxref_54_M45_noxref_s ) capacitor \
 c=0.00211573f //x=75.145 //y=1.56 //x2=73.82 //y2=0.365
cc_3826 ( N_noxref_13_c_4735_p N_noxref_54_M45_noxref_s ) capacitor \
 c=0.0133026f //x=75.675 //y=0.905 //x2=73.82 //y2=0.365
cc_3827 ( N_noxref_13_c_4738_p N_noxref_54_M45_noxref_s ) capacitor \
 c=0.00793126f //x=75.675 //y=1.25 //x2=73.82 //y2=0.365
cc_3828 ( N_noxref_13_c_4888_p N_noxref_54_M45_noxref_s ) capacitor \
 c=0.00392195f //x=75.11 //y=1.915 //x2=73.82 //y2=0.365
cc_3829 ( N_noxref_13_c_4444_n N_noxref_56_c_10727_n ) capacitor c=0.00631223f \
 //x=81.655 //y=4.07 //x2=81.5 //y2=1.58
cc_3830 ( N_noxref_13_c_4444_n N_noxref_56_c_10733_n ) capacitor c=0.00108825f \
 //x=81.655 //y=4.07 //x2=81.585 //y2=1.495
cc_3831 ( N_noxref_13_c_4770_p N_noxref_56_c_10733_n ) capacitor c=0.00698471f \
 //x=81.805 //y=1.56 //x2=81.585 //y2=1.495
cc_3832 ( N_noxref_13_c_4756_p N_noxref_56_c_10733_n ) capacitor c=0.00171785f \
 //x=81.77 //y=2.08 //x2=81.585 //y2=1.495
cc_3833 ( N_noxref_13_c_4451_n N_noxref_56_c_10734_n ) capacitor c=0.00118117f \
 //x=81.77 //y=2.08 //x2=82.47 //y2=0.53
cc_3834 ( N_noxref_13_c_4768_p N_noxref_56_c_10734_n ) capacitor c=0.0191024f \
 //x=81.805 //y=0.905 //x2=82.47 //y2=0.53
cc_3835 ( N_noxref_13_c_4778_p N_noxref_56_c_10734_n ) capacitor c=0.00655165f \
 //x=82.335 //y=0.905 //x2=82.47 //y2=0.53
cc_3836 ( N_noxref_13_c_4756_p N_noxref_56_c_10734_n ) capacitor c=2.1838e-19 \
 //x=81.77 //y=2.08 //x2=82.47 //y2=0.53
cc_3837 ( N_noxref_13_c_4768_p N_noxref_56_M49_noxref_s ) capacitor \
 c=0.00698471f //x=81.805 //y=0.905 //x2=80.48 //y2=0.365
cc_3838 ( N_noxref_13_c_4781_p N_noxref_56_M49_noxref_s ) capacitor \
 c=0.00316186f //x=82.18 //y=1.405 //x2=80.48 //y2=0.365
cc_3839 ( N_noxref_13_c_4778_p N_noxref_56_M49_noxref_s ) capacitor \
 c=0.0142835f //x=82.335 //y=0.905 //x2=80.48 //y2=0.365
cc_3840 ( N_D_M113_noxref_g N_noxref_15_c_5253_n ) capacitor c=0.0169521f \
 //x=50.29 //y=6.02 //x2=50.865 //y2=5.2
cc_3841 ( N_D_c_4917_n N_noxref_15_c_5257_n ) capacitor c=0.00539951f \
 //x=49.95 //y=2.08 //x2=50.155 //y2=5.2
cc_3842 ( N_D_M112_noxref_g N_noxref_15_c_5257_n ) capacitor c=0.0177326f \
 //x=49.85 //y=6.02 //x2=50.155 //y2=5.2
cc_3843 ( N_D_c_4973_n N_noxref_15_c_5257_n ) capacitor c=0.00581252f \
 //x=49.95 //y=4.7 //x2=50.155 //y2=5.2
cc_3844 ( N_D_c_4917_n N_noxref_15_c_5226_n ) capacitor c=0.00337041f \
 //x=49.95 //y=2.08 //x2=51.43 //y2=2.59
cc_3845 ( N_D_M113_noxref_g N_noxref_15_M112_noxref_d ) capacitor c=0.0173476f \
 //x=50.29 //y=6.02 //x2=49.925 //y2=5.02
cc_3846 ( N_D_c_4900_n N_CLK_c_5631_n ) capacitor c=0.00594004f //x=25.415 \
 //y=2.96 //x2=14.685 //y2=4.44
cc_3847 ( N_D_c_4900_n N_CLK_c_5642_n ) capacitor c=6.59274e-19 //x=25.415 \
 //y=2.96 //x2=5.665 //y2=4.44
cc_3848 ( N_D_c_4900_n N_CLK_c_5643_n ) capacitor c=0.0121978f //x=25.415 \
 //y=2.96 //x2=29.855 //y2=4.44
cc_3849 ( N_D_c_4909_n N_CLK_c_5643_n ) capacitor c=0.00334314f //x=49.835 \
 //y=2.96 //x2=29.855 //y2=4.44
cc_3850 ( N_D_c_5060_n N_CLK_c_5643_n ) capacitor c=3.52702e-19 //x=25.645 \
 //y=2.96 //x2=29.855 //y2=4.44
cc_3851 ( N_D_c_4916_n N_CLK_c_5643_n ) capacitor c=0.0236903f //x=25.53 \
 //y=2.08 //x2=29.855 //y2=4.44
cc_3852 ( N_D_c_4972_n N_CLK_c_5643_n ) capacitor c=0.00890426f //x=25.53 \
 //y=4.7 //x2=29.855 //y2=4.44
cc_3853 ( N_D_c_4909_n N_CLK_c_5680_n ) capacitor c=0.00675488f //x=49.835 \
 //y=2.96 //x2=54.275 //y2=4.44
cc_3854 ( N_D_c_4917_n N_CLK_c_5680_n ) capacitor c=0.0236903f //x=49.95 \
 //y=2.08 //x2=54.275 //y2=4.44
cc_3855 ( N_D_c_4973_n N_CLK_c_5680_n ) capacitor c=0.00890426f //x=49.95 \
 //y=4.7 //x2=54.275 //y2=4.44
cc_3856 ( N_D_c_4900_n N_CLK_c_5622_n ) capacitor c=0.0228892f //x=25.415 \
 //y=2.96 //x2=5.55 //y2=2.08
cc_3857 ( N_D_c_4900_n N_CLK_c_5623_n ) capacitor c=0.0215847f //x=25.415 \
 //y=2.96 //x2=14.8 //y2=2.08
cc_3858 ( N_D_c_4909_n N_CLK_c_5625_n ) capacitor c=0.0190322f //x=49.835 \
 //y=2.96 //x2=29.97 //y2=2.08
cc_3859 ( N_D_c_4909_n N_CLK_c_5626_n ) capacitor c=0.0192451f //x=49.835 \
 //y=2.96 //x2=39.22 //y2=2.08
cc_3860 ( N_D_c_4917_n N_noxref_18_c_6449_n ) capacitor c=0.00423741f \
 //x=49.95 //y=2.08 //x2=50.805 //y2=4.07
cc_3861 ( N_D_c_4917_n N_noxref_18_c_6458_n ) capacitor c=0.00400249f \
 //x=49.95 //y=2.08 //x2=50.69 //y2=4.535
cc_3862 ( N_D_c_4973_n N_noxref_18_c_6458_n ) capacitor c=0.00417994f \
 //x=49.95 //y=4.7 //x2=50.69 //y2=4.535
cc_3863 ( N_D_c_4909_n N_noxref_18_c_6377_n ) capacitor c=0.00262125f \
 //x=49.835 //y=2.96 //x2=50.69 //y2=2.08
cc_3864 ( N_D_c_4917_n N_noxref_18_c_6377_n ) capacitor c=0.0734198f //x=49.95 \
 //y=2.08 //x2=50.69 //y2=2.08
cc_3865 ( N_D_c_4942_n N_noxref_18_c_6377_n ) capacitor c=0.00284029f \
 //x=49.755 //y=1.915 //x2=50.69 //y2=2.08
cc_3866 ( N_D_M112_noxref_g N_noxref_18_M114_noxref_g ) capacitor c=0.0104611f \
 //x=49.85 //y=6.02 //x2=50.73 //y2=6.02
cc_3867 ( N_D_M113_noxref_g N_noxref_18_M114_noxref_g ) capacitor c=0.106811f \
 //x=50.29 //y=6.02 //x2=50.73 //y2=6.02
cc_3868 ( N_D_M113_noxref_g N_noxref_18_M115_noxref_g ) capacitor c=0.0100341f \
 //x=50.29 //y=6.02 //x2=51.17 //y2=6.02
cc_3869 ( N_D_c_4938_n N_noxref_18_c_6466_n ) capacitor c=4.86506e-19 \
 //x=49.755 //y=0.865 //x2=50.725 //y2=0.905
cc_3870 ( N_D_c_4940_n N_noxref_18_c_6466_n ) capacitor c=0.00152104f \
 //x=49.755 //y=1.21 //x2=50.725 //y2=0.905
cc_3871 ( N_D_c_4945_n N_noxref_18_c_6466_n ) capacitor c=0.0151475f \
 //x=50.285 //y=0.865 //x2=50.725 //y2=0.905
cc_3872 ( N_D_c_4941_n N_noxref_18_c_6469_n ) capacitor c=0.00109982f \
 //x=49.755 //y=1.52 //x2=50.725 //y2=1.25
cc_3873 ( N_D_c_4947_n N_noxref_18_c_6469_n ) capacitor c=0.0111064f \
 //x=50.285 //y=1.21 //x2=50.725 //y2=1.25
cc_3874 ( N_D_c_4941_n N_noxref_18_c_6471_n ) capacitor c=9.57794e-19 \
 //x=49.755 //y=1.52 //x2=50.725 //y2=1.56
cc_3875 ( N_D_c_4942_n N_noxref_18_c_6471_n ) capacitor c=0.00662747f \
 //x=49.755 //y=1.915 //x2=50.725 //y2=1.56
cc_3876 ( N_D_c_4947_n N_noxref_18_c_6471_n ) capacitor c=0.00862358f \
 //x=50.285 //y=1.21 //x2=50.725 //y2=1.56
cc_3877 ( N_D_c_4945_n N_noxref_18_c_6474_n ) capacitor c=0.00124821f \
 //x=50.285 //y=0.865 //x2=51.255 //y2=0.905
cc_3878 ( N_D_c_4947_n N_noxref_18_c_6475_n ) capacitor c=0.00200715f \
 //x=50.285 //y=1.21 //x2=51.255 //y2=1.25
cc_3879 ( N_D_c_4917_n N_noxref_18_c_6476_n ) capacitor c=0.00282278f \
 //x=49.95 //y=2.08 //x2=50.69 //y2=2.08
cc_3880 ( N_D_c_4942_n N_noxref_18_c_6476_n ) capacitor c=0.0172771f \
 //x=49.755 //y=1.915 //x2=50.69 //y2=2.08
cc_3881 ( N_D_c_4917_n N_noxref_18_c_6478_n ) capacitor c=0.00344981f \
 //x=49.95 //y=2.08 //x2=50.72 //y2=4.7
cc_3882 ( N_D_c_4973_n N_noxref_18_c_6478_n ) capacitor c=0.0293367f //x=49.95 \
 //y=4.7 //x2=50.72 //y2=4.7
cc_3883 ( N_D_c_4900_n N_SN_c_6833_n ) capacitor c=0.395089f //x=25.415 \
 //y=2.96 //x2=21.715 //y2=2.22
cc_3884 ( N_D_c_4900_n N_SN_c_6843_n ) capacitor c=0.0132772f //x=25.415 \
 //y=2.96 //x2=10.475 //y2=2.22
cc_3885 ( N_D_c_4900_n N_SN_c_6844_n ) capacitor c=0.146261f //x=25.415 \
 //y=2.96 //x2=34.665 //y2=2.22
cc_3886 ( N_D_c_4909_n N_SN_c_6844_n ) capacitor c=0.13581f //x=49.835 \
 //y=2.96 //x2=34.665 //y2=2.22
cc_3887 ( N_D_c_5060_n N_SN_c_6844_n ) capacitor c=0.0120598f //x=25.645 \
 //y=2.96 //x2=34.665 //y2=2.22
cc_3888 ( N_D_c_4916_n N_SN_c_6844_n ) capacitor c=0.0211592f //x=25.53 \
 //y=2.08 //x2=34.665 //y2=2.22
cc_3889 ( N_D_c_4932_n N_SN_c_6844_n ) capacitor c=0.00894156f //x=25.335 \
 //y=1.915 //x2=34.665 //y2=2.22
cc_3890 ( N_D_c_4900_n N_SN_c_6854_n ) capacitor c=0.0120222f //x=25.415 \
 //y=2.96 //x2=21.945 //y2=2.22
cc_3891 ( N_D_c_4909_n N_SN_c_6855_n ) capacitor c=0.316819f //x=49.835 \
 //y=2.96 //x2=46.135 //y2=2.22
cc_3892 ( N_D_c_4909_n N_SN_c_6865_n ) capacitor c=0.0120222f //x=49.835 \
 //y=2.96 //x2=34.895 //y2=2.22
cc_3893 ( N_D_c_4909_n N_SN_c_6866_n ) capacitor c=0.0792983f //x=49.835 \
 //y=2.96 //x2=59.085 //y2=2.22
cc_3894 ( N_D_c_4917_n N_SN_c_6866_n ) capacitor c=0.0185012f //x=49.95 \
 //y=2.08 //x2=59.085 //y2=2.22
cc_3895 ( N_D_c_4942_n N_SN_c_6866_n ) capacitor c=0.00894156f //x=49.755 \
 //y=1.915 //x2=59.085 //y2=2.22
cc_3896 ( N_D_c_4909_n N_SN_c_6876_n ) capacitor c=0.0120222f //x=49.835 \
 //y=2.96 //x2=46.365 //y2=2.22
cc_3897 ( N_D_c_4900_n N_SN_c_6888_n ) capacitor c=0.0239871f //x=25.415 \
 //y=2.96 //x2=10.36 //y2=2.08
cc_3898 ( N_D_c_4900_n N_SN_c_6889_n ) capacitor c=0.0216476f //x=25.415 \
 //y=2.96 //x2=21.83 //y2=2.08
cc_3899 ( N_D_c_4909_n N_SN_c_6890_n ) capacitor c=0.0216476f //x=49.835 \
 //y=2.96 //x2=34.78 //y2=2.08
cc_3900 ( N_D_c_4909_n N_SN_c_6891_n ) capacitor c=0.0216476f //x=49.835 \
 //y=2.96 //x2=46.25 //y2=2.08
cc_3901 ( N_D_c_4900_n N_noxref_24_c_8520_n ) capacitor c=0.46661f //x=25.415 \
 //y=2.96 //x2=23.565 //y2=3.33
cc_3902 ( N_D_c_4900_n N_noxref_24_c_8497_n ) capacitor c=0.0291053f \
 //x=25.415 //y=2.96 //x2=18.245 //y2=3.33
cc_3903 ( N_D_c_4900_n N_noxref_24_c_8424_n ) capacitor c=0.144311f //x=25.415 \
 //y=2.96 //x2=79.065 //y2=3.33
cc_3904 ( N_D_c_4909_n N_noxref_24_c_8424_n ) capacitor c=2.15187f //x=49.835 \
 //y=2.96 //x2=79.065 //y2=3.33
cc_3905 ( N_D_c_5060_n N_noxref_24_c_8424_n ) capacitor c=0.026764f //x=25.645 \
 //y=2.96 //x2=79.065 //y2=3.33
cc_3906 ( N_D_c_4916_n N_noxref_24_c_8424_n ) capacitor c=0.0244325f //x=25.53 \
 //y=2.08 //x2=79.065 //y2=3.33
cc_3907 ( N_D_c_4917_n N_noxref_24_c_8424_n ) capacitor c=0.0244325f //x=49.95 \
 //y=2.08 //x2=79.065 //y2=3.33
cc_3908 ( N_D_c_4900_n N_noxref_24_c_8558_n ) capacitor c=0.0266688f \
 //x=25.415 //y=2.96 //x2=23.795 //y2=3.33
cc_3909 ( N_D_c_4916_n N_noxref_24_c_8558_n ) capacitor c=7.01366e-19 \
 //x=25.53 //y=2.08 //x2=23.795 //y2=3.33
cc_3910 ( N_D_c_4900_n N_noxref_24_c_8428_n ) capacitor c=0.0210797f \
 //x=25.415 //y=2.96 //x2=18.13 //y2=2.08
cc_3911 ( N_D_c_4900_n N_noxref_24_c_8465_n ) capacitor c=0.0229057f \
 //x=25.415 //y=2.96 //x2=23.68 //y2=3.33
cc_3912 ( N_D_c_5060_n N_noxref_24_c_8465_n ) capacitor c=7.01366e-19 \
 //x=25.645 //y=2.96 //x2=23.68 //y2=3.33
cc_3913 ( N_D_c_4916_n N_noxref_24_c_8465_n ) capacitor c=0.013729f //x=25.53 \
 //y=2.08 //x2=23.68 //y2=3.33
cc_3914 ( N_D_c_4922_n N_noxref_27_c_9246_n ) capacitor c=0.0034165f //x=0.915 \
 //y=1.915 //x2=0.695 //y2=1.495
cc_3915 ( N_D_c_4900_n N_noxref_27_c_9228_n ) capacitor c=0.00547841f \
 //x=25.415 //y=2.96 //x2=1.58 //y2=1.58
cc_3916 ( N_D_c_4908_n N_noxref_27_c_9228_n ) capacitor c=0.00242864f \
 //x=1.225 //y=2.96 //x2=1.58 //y2=1.58
cc_3917 ( N_D_c_4915_n N_noxref_27_c_9228_n ) capacitor c=0.0115783f //x=1.11 \
 //y=2.08 //x2=1.58 //y2=1.58
cc_3918 ( N_D_c_4921_n N_noxref_27_c_9228_n ) capacitor c=0.00703567f \
 //x=0.915 //y=1.52 //x2=1.58 //y2=1.58
cc_3919 ( N_D_c_4922_n N_noxref_27_c_9228_n ) capacitor c=0.0209643f //x=0.915 \
 //y=1.915 //x2=1.58 //y2=1.58
cc_3920 ( N_D_c_4924_n N_noxref_27_c_9228_n ) capacitor c=0.00780629f //x=1.29 \
 //y=1.365 //x2=1.58 //y2=1.58
cc_3921 ( N_D_c_4927_n N_noxref_27_c_9228_n ) capacitor c=0.00339872f \
 //x=1.445 //y=1.21 //x2=1.58 //y2=1.58
cc_3922 ( N_D_c_4900_n N_noxref_27_c_9235_n ) capacitor c=0.00311515f \
 //x=25.415 //y=2.96 //x2=1.665 //y2=1.495
cc_3923 ( N_D_c_4922_n N_noxref_27_c_9235_n ) capacitor c=6.71402e-19 \
 //x=0.915 //y=1.915 //x2=1.665 //y2=1.495
cc_3924 ( N_D_c_4900_n N_noxref_27_c_9236_n ) capacitor c=7.29507e-19 \
 //x=25.415 //y=2.96 //x2=2.55 //y2=0.53
cc_3925 ( N_D_c_4918_n N_noxref_27_M0_noxref_s ) capacitor c=0.0326577f \
 //x=0.915 //y=0.865 //x2=0.56 //y2=0.365
cc_3926 ( N_D_c_4921_n N_noxref_27_M0_noxref_s ) capacitor c=3.48408e-19 \
 //x=0.915 //y=1.52 //x2=0.56 //y2=0.365
cc_3927 ( N_D_c_4925_n N_noxref_27_M0_noxref_s ) capacitor c=0.0120759f \
 //x=1.445 //y=0.865 //x2=0.56 //y2=0.365
cc_3928 ( N_D_c_4900_n N_noxref_30_c_9381_n ) capacitor c=0.00351507f \
 //x=25.415 //y=2.96 //x2=9.615 //y2=1.59
cc_3929 ( N_D_c_4900_n N_noxref_30_c_9412_n ) capacitor c=0.00667312f \
 //x=25.415 //y=2.96 //x2=10.585 //y2=1.59
cc_3930 ( N_D_c_4900_n N_noxref_30_M5_noxref_s ) capacitor c=0.00324882f \
 //x=25.415 //y=2.96 //x2=8.595 //y2=0.375
cc_3931 ( N_D_c_4932_n N_noxref_36_c_9710_n ) capacitor c=0.0034165f \
 //x=25.335 //y=1.915 //x2=25.115 //y2=1.495
cc_3932 ( N_D_c_4916_n N_noxref_36_c_9692_n ) capacitor c=0.0111916f //x=25.53 \
 //y=2.08 //x2=26 //y2=1.58
cc_3933 ( N_D_c_4931_n N_noxref_36_c_9692_n ) capacitor c=0.00696403f \
 //x=25.335 //y=1.52 //x2=26 //y2=1.58
cc_3934 ( N_D_c_4932_n N_noxref_36_c_9692_n ) capacitor c=0.0174694f \
 //x=25.335 //y=1.915 //x2=26 //y2=1.58
cc_3935 ( N_D_c_4934_n N_noxref_36_c_9692_n ) capacitor c=0.00776811f \
 //x=25.71 //y=1.365 //x2=26 //y2=1.58
cc_3936 ( N_D_c_4937_n N_noxref_36_c_9692_n ) capacitor c=0.00339872f \
 //x=25.865 //y=1.21 //x2=26 //y2=1.58
cc_3937 ( N_D_c_4932_n N_noxref_36_c_9699_n ) capacitor c=6.71402e-19 \
 //x=25.335 //y=1.915 //x2=26.085 //y2=1.495
cc_3938 ( N_D_c_4928_n N_noxref_36_M15_noxref_s ) capacitor c=0.0327502f \
 //x=25.335 //y=0.865 //x2=24.98 //y2=0.365
cc_3939 ( N_D_c_4931_n N_noxref_36_M15_noxref_s ) capacitor c=3.48408e-19 \
 //x=25.335 //y=1.52 //x2=24.98 //y2=0.365
cc_3940 ( N_D_c_4935_n N_noxref_36_M15_noxref_s ) capacitor c=0.0120759f \
 //x=25.865 //y=0.865 //x2=24.98 //y2=0.365
cc_3941 ( N_D_c_4942_n N_noxref_45_c_10172_n ) capacitor c=0.0034165f \
 //x=49.755 //y=1.915 //x2=49.535 //y2=1.495
cc_3942 ( N_D_c_4917_n N_noxref_45_c_10154_n ) capacitor c=0.0111916f \
 //x=49.95 //y=2.08 //x2=50.42 //y2=1.58
cc_3943 ( N_D_c_4941_n N_noxref_45_c_10154_n ) capacitor c=0.00696403f \
 //x=49.755 //y=1.52 //x2=50.42 //y2=1.58
cc_3944 ( N_D_c_4942_n N_noxref_45_c_10154_n ) capacitor c=0.0174694f \
 //x=49.755 //y=1.915 //x2=50.42 //y2=1.58
cc_3945 ( N_D_c_4944_n N_noxref_45_c_10154_n ) capacitor c=0.00776811f \
 //x=50.13 //y=1.365 //x2=50.42 //y2=1.58
cc_3946 ( N_D_c_4947_n N_noxref_45_c_10154_n ) capacitor c=0.00339872f \
 //x=50.285 //y=1.21 //x2=50.42 //y2=1.58
cc_3947 ( N_D_c_4942_n N_noxref_45_c_10161_n ) capacitor c=6.71402e-19 \
 //x=49.755 //y=1.915 //x2=50.505 //y2=1.495
cc_3948 ( N_D_c_4938_n N_noxref_45_M30_noxref_s ) capacitor c=0.0327502f \
 //x=49.755 //y=0.865 //x2=49.4 //y2=0.365
cc_3949 ( N_D_c_4941_n N_noxref_45_M30_noxref_s ) capacitor c=3.48408e-19 \
 //x=49.755 //y=1.52 //x2=49.4 //y2=0.365
cc_3950 ( N_D_c_4945_n N_noxref_45_M30_noxref_s ) capacitor c=0.0120759f \
 //x=50.285 //y=0.865 //x2=49.4 //y2=0.365
cc_3951 ( N_noxref_15_c_5223_n N_noxref_16_c_5459_n ) capacitor c=0.00564994f \
 //x=57.975 //y=2.59 //x2=61.165 //y2=2.59
cc_3952 ( N_noxref_15_M123_noxref_g N_noxref_16_c_5474_n ) capacitor \
 c=0.0168349f //x=58.73 //y=6.02 //x2=59.305 //y2=5.155
cc_3953 ( N_noxref_15_M122_noxref_g N_noxref_16_c_5478_n ) capacitor \
 c=0.0213876f //x=58.29 //y=6.02 //x2=58.595 //y2=5.155
cc_3954 ( N_noxref_15_c_5315_p N_noxref_16_c_5478_n ) capacitor c=0.00428486f \
 //x=58.655 //y=4.79 //x2=58.595 //y2=5.155
cc_3955 ( N_noxref_15_M123_noxref_g N_noxref_16_M122_noxref_d ) capacitor \
 c=0.0180032f //x=58.73 //y=6.02 //x2=58.365 //y2=5.02
cc_3956 ( N_noxref_15_c_5253_n N_CLK_c_5680_n ) capacitor c=0.0185297f \
 //x=50.865 //y=5.2 //x2=54.275 //y2=4.44
cc_3957 ( N_noxref_15_c_5257_n N_CLK_c_5680_n ) capacitor c=0.018142f \
 //x=50.155 //y=5.2 //x2=54.275 //y2=4.44
cc_3958 ( N_noxref_15_c_5226_n N_CLK_c_5680_n ) capacitor c=0.0208321f \
 //x=51.43 //y=2.59 //x2=54.275 //y2=4.44
cc_3959 ( N_noxref_15_c_5228_n N_CLK_c_5680_n ) capacitor c=0.0208709f \
 //x=53.28 //y=2.08 //x2=54.275 //y2=4.44
cc_3960 ( N_noxref_15_c_5278_n N_CLK_c_5680_n ) capacitor c=0.0166984f \
 //x=53.555 //y=4.79 //x2=54.275 //y2=4.44
cc_3961 ( N_noxref_15_c_5229_n N_CLK_c_5705_n ) capacitor c=0.0208709f \
 //x=58.09 //y=2.08 //x2=63.525 //y2=4.44
cc_3962 ( N_noxref_15_c_5280_n N_CLK_c_5705_n ) capacitor c=0.0166984f \
 //x=58.365 //y=4.79 //x2=63.525 //y2=4.44
cc_3963 ( N_noxref_15_c_5228_n N_CLK_c_5716_n ) capacitor c=0.00153281f \
 //x=53.28 //y=2.08 //x2=54.505 //y2=4.44
cc_3964 ( N_noxref_15_c_5223_n N_CLK_c_5628_n ) capacitor c=0.0190006f \
 //x=57.975 //y=2.59 //x2=54.39 //y2=2.08
cc_3965 ( N_noxref_15_c_5224_n N_CLK_c_5628_n ) capacitor c=0.00103784f \
 //x=53.545 //y=2.59 //x2=54.39 //y2=2.08
cc_3966 ( N_noxref_15_c_5226_n N_CLK_c_5628_n ) capacitor c=3.63796e-19 \
 //x=51.43 //y=2.59 //x2=54.39 //y2=2.08
cc_3967 ( N_noxref_15_c_5228_n N_CLK_c_5628_n ) capacitor c=0.0435204f \
 //x=53.28 //y=2.08 //x2=54.39 //y2=2.08
cc_3968 ( N_noxref_15_c_5234_n N_CLK_c_5628_n ) capacitor c=0.00210802f \
 //x=52.98 //y=1.915 //x2=54.39 //y2=2.08
cc_3969 ( N_noxref_15_c_5330_p N_CLK_c_5628_n ) capacitor c=0.00147352f \
 //x=53.845 //y=4.79 //x2=54.39 //y2=2.08
cc_3970 ( N_noxref_15_c_5278_n N_CLK_c_5628_n ) capacitor c=0.00141297f \
 //x=53.555 //y=4.79 //x2=54.39 //y2=2.08
cc_3971 ( N_noxref_15_M116_noxref_g N_CLK_M118_noxref_g ) capacitor \
 c=0.0105869f //x=53.48 //y=6.02 //x2=54.36 //y2=6.02
cc_3972 ( N_noxref_15_M117_noxref_g N_CLK_M118_noxref_g ) capacitor c=0.10632f \
 //x=53.92 //y=6.02 //x2=54.36 //y2=6.02
cc_3973 ( N_noxref_15_M117_noxref_g N_CLK_M119_noxref_g ) capacitor \
 c=0.0101598f //x=53.92 //y=6.02 //x2=54.8 //y2=6.02
cc_3974 ( N_noxref_15_c_5230_n N_CLK_c_6114_n ) capacitor c=5.72482e-19 \
 //x=52.98 //y=0.875 //x2=53.955 //y2=0.91
cc_3975 ( N_noxref_15_c_5232_n N_CLK_c_6114_n ) capacitor c=0.00149976f \
 //x=52.98 //y=1.22 //x2=53.955 //y2=0.91
cc_3976 ( N_noxref_15_c_5237_n N_CLK_c_6114_n ) capacitor c=0.0160123f \
 //x=53.51 //y=0.875 //x2=53.955 //y2=0.91
cc_3977 ( N_noxref_15_c_5233_n N_CLK_c_6117_n ) capacitor c=0.00111227f \
 //x=52.98 //y=1.53 //x2=53.955 //y2=1.22
cc_3978 ( N_noxref_15_c_5239_n N_CLK_c_6117_n ) capacitor c=0.0124075f \
 //x=53.51 //y=1.22 //x2=53.955 //y2=1.22
cc_3979 ( N_noxref_15_c_5237_n N_CLK_c_6119_n ) capacitor c=0.00103227f \
 //x=53.51 //y=0.875 //x2=54.48 //y2=0.91
cc_3980 ( N_noxref_15_c_5239_n N_CLK_c_6120_n ) capacitor c=0.0010154f \
 //x=53.51 //y=1.22 //x2=54.48 //y2=1.22
cc_3981 ( N_noxref_15_c_5239_n N_CLK_c_6121_n ) capacitor c=9.23422e-19 \
 //x=53.51 //y=1.22 //x2=54.48 //y2=1.45
cc_3982 ( N_noxref_15_c_5228_n N_CLK_c_6122_n ) capacitor c=0.00203769f \
 //x=53.28 //y=2.08 //x2=54.48 //y2=1.915
cc_3983 ( N_noxref_15_c_5234_n N_CLK_c_6122_n ) capacitor c=0.00834532f \
 //x=52.98 //y=1.915 //x2=54.48 //y2=1.915
cc_3984 ( N_noxref_15_c_5228_n N_CLK_c_6124_n ) capacitor c=0.00183762f \
 //x=53.28 //y=2.08 //x2=54.39 //y2=4.7
cc_3985 ( N_noxref_15_c_5330_p N_CLK_c_6124_n ) capacitor c=0.0168581f \
 //x=53.845 //y=4.79 //x2=54.39 //y2=4.7
cc_3986 ( N_noxref_15_c_5278_n N_CLK_c_6124_n ) capacitor c=0.00484466f \
 //x=53.555 //y=4.79 //x2=54.39 //y2=4.7
cc_3987 ( N_noxref_15_c_5226_n N_noxref_18_c_6392_n ) capacitor c=0.0205341f \
 //x=51.43 //y=2.59 //x2=56.12 //y2=4.07
cc_3988 ( N_noxref_15_c_5228_n N_noxref_18_c_6392_n ) capacitor c=0.021838f \
 //x=53.28 //y=2.08 //x2=56.12 //y2=4.07
cc_3989 ( N_noxref_15_c_5226_n N_noxref_18_c_6449_n ) capacitor c=0.00131333f \
 //x=51.43 //y=2.59 //x2=50.805 //y2=4.07
cc_3990 ( N_noxref_15_c_5229_n N_noxref_18_c_6393_n ) capacitor c=0.0194977f \
 //x=58.09 //y=2.08 //x2=66.115 //y2=4.07
cc_3991 ( N_noxref_15_c_5229_n N_noxref_18_c_6402_n ) capacitor c=3.49381e-19 \
 //x=58.09 //y=2.08 //x2=56.35 //y2=4.07
cc_3992 ( N_noxref_15_c_5253_n N_noxref_18_c_6458_n ) capacitor c=0.0126603f \
 //x=50.865 //y=5.2 //x2=50.69 //y2=4.535
cc_3993 ( N_noxref_15_c_5226_n N_noxref_18_c_6458_n ) capacitor c=0.0101115f \
 //x=51.43 //y=2.59 //x2=50.69 //y2=4.535
cc_3994 ( N_noxref_15_c_5222_n N_noxref_18_c_6377_n ) capacitor c=0.00228021f \
 //x=51.545 //y=2.59 //x2=50.69 //y2=2.08
cc_3995 ( N_noxref_15_c_5226_n N_noxref_18_c_6377_n ) capacitor c=0.0672954f \
 //x=51.43 //y=2.59 //x2=50.69 //y2=2.08
cc_3996 ( N_noxref_15_c_5228_n N_noxref_18_c_6377_n ) capacitor c=6.6118e-19 \
 //x=53.28 //y=2.08 //x2=50.69 //y2=2.08
cc_3997 ( N_noxref_15_M117_noxref_g N_noxref_18_c_6405_n ) capacitor \
 c=0.0168349f //x=53.92 //y=6.02 //x2=54.495 //y2=5.155
cc_3998 ( N_noxref_15_c_5226_n N_noxref_18_c_6409_n ) capacitor c=2.97874e-19 \
 //x=51.43 //y=2.59 //x2=53.785 //y2=5.155
cc_3999 ( N_noxref_15_M116_noxref_g N_noxref_18_c_6409_n ) capacitor \
 c=0.0213876f //x=53.48 //y=6.02 //x2=53.785 //y2=5.155
cc_4000 ( N_noxref_15_c_5330_p N_noxref_18_c_6409_n ) capacitor c=0.00428486f \
 //x=53.845 //y=4.79 //x2=53.785 //y2=5.155
cc_4001 ( N_noxref_15_c_5223_n N_noxref_18_c_6456_n ) capacitor c=0.0165903f \
 //x=57.975 //y=2.59 //x2=56.237 //y2=3.905
cc_4002 ( N_noxref_15_c_5229_n N_noxref_18_c_6456_n ) capacitor c=0.0109272f \
 //x=58.09 //y=2.08 //x2=56.237 //y2=3.905
cc_4003 ( N_noxref_15_c_5253_n N_noxref_18_M114_noxref_g ) capacitor \
 c=0.0166421f //x=50.865 //y=5.2 //x2=50.73 //y2=6.02
cc_4004 ( N_noxref_15_M114_noxref_d N_noxref_18_M114_noxref_g ) capacitor \
 c=0.0173476f //x=50.805 //y=5.02 //x2=50.73 //y2=6.02
cc_4005 ( N_noxref_15_c_5259_n N_noxref_18_M115_noxref_g ) capacitor \
 c=0.018922f //x=51.345 //y=5.2 //x2=51.17 //y2=6.02
cc_4006 ( N_noxref_15_M114_noxref_d N_noxref_18_M115_noxref_g ) capacitor \
 c=0.0179769f //x=50.805 //y=5.02 //x2=51.17 //y2=6.02
cc_4007 ( N_noxref_15_M31_noxref_d N_noxref_18_c_6466_n ) capacitor \
 c=0.00217566f //x=50.8 //y=0.905 //x2=50.725 //y2=0.905
cc_4008 ( N_noxref_15_M31_noxref_d N_noxref_18_c_6469_n ) capacitor \
 c=0.0034598f //x=50.8 //y=0.905 //x2=50.725 //y2=1.25
cc_4009 ( N_noxref_15_M31_noxref_d N_noxref_18_c_6471_n ) capacitor \
 c=0.00669531f //x=50.8 //y=0.905 //x2=50.725 //y2=1.56
cc_4010 ( N_noxref_15_c_5226_n N_noxref_18_c_6503_n ) capacitor c=0.0142673f \
 //x=51.43 //y=2.59 //x2=51.095 //y2=4.79
cc_4011 ( N_noxref_15_c_5372_p N_noxref_18_c_6503_n ) capacitor c=0.00407665f \
 //x=50.95 //y=5.2 //x2=51.095 //y2=4.79
cc_4012 ( N_noxref_15_M31_noxref_d N_noxref_18_c_6505_n ) capacitor \
 c=0.00241102f //x=50.8 //y=0.905 //x2=51.1 //y2=0.75
cc_4013 ( N_noxref_15_c_5225_n N_noxref_18_c_6506_n ) capacitor c=0.00371277f \
 //x=51.345 //y=1.655 //x2=51.1 //y2=1.405
cc_4014 ( N_noxref_15_M31_noxref_d N_noxref_18_c_6506_n ) capacitor \
 c=0.0137169f //x=50.8 //y=0.905 //x2=51.1 //y2=1.405
cc_4015 ( N_noxref_15_M31_noxref_d N_noxref_18_c_6474_n ) capacitor \
 c=0.00132245f //x=50.8 //y=0.905 //x2=51.255 //y2=0.905
cc_4016 ( N_noxref_15_c_5225_n N_noxref_18_c_6475_n ) capacitor c=0.00457401f \
 //x=51.345 //y=1.655 //x2=51.255 //y2=1.25
cc_4017 ( N_noxref_15_M31_noxref_d N_noxref_18_c_6475_n ) capacitor \
 c=0.00566463f //x=50.8 //y=0.905 //x2=51.255 //y2=1.25
cc_4018 ( N_noxref_15_c_5226_n N_noxref_18_c_6476_n ) capacitor c=0.00731987f \
 //x=51.43 //y=2.59 //x2=50.69 //y2=2.08
cc_4019 ( N_noxref_15_c_5226_n N_noxref_18_c_6512_n ) capacitor c=0.00306024f \
 //x=51.43 //y=2.59 //x2=50.69 //y2=1.915
cc_4020 ( N_noxref_15_M31_noxref_d N_noxref_18_c_6512_n ) capacitor \
 c=0.00660593f //x=50.8 //y=0.905 //x2=50.69 //y2=1.915
cc_4021 ( N_noxref_15_c_5253_n N_noxref_18_c_6478_n ) capacitor c=0.00346527f \
 //x=50.865 //y=5.2 //x2=50.72 //y2=4.7
cc_4022 ( N_noxref_15_c_5226_n N_noxref_18_c_6478_n ) capacitor c=0.00517969f \
 //x=51.43 //y=2.59 //x2=50.72 //y2=4.7
cc_4023 ( N_noxref_15_M117_noxref_g N_noxref_18_M116_noxref_d ) capacitor \
 c=0.0180032f //x=53.92 //y=6.02 //x2=53.555 //y2=5.02
cc_4024 ( N_noxref_15_c_5221_n N_SN_c_6866_n ) capacitor c=0.140806f \
 //x=53.135 //y=2.59 //x2=59.085 //y2=2.22
cc_4025 ( N_noxref_15_c_5222_n N_SN_c_6866_n ) capacitor c=0.0290445f \
 //x=51.545 //y=2.59 //x2=59.085 //y2=2.22
cc_4026 ( N_noxref_15_c_5223_n N_SN_c_6866_n ) capacitor c=0.414292f \
 //x=57.975 //y=2.59 //x2=59.085 //y2=2.22
cc_4027 ( N_noxref_15_c_5224_n N_SN_c_6866_n ) capacitor c=0.0429267f \
 //x=53.545 //y=2.59 //x2=59.085 //y2=2.22
cc_4028 ( N_noxref_15_c_5389_p N_SN_c_6866_n ) capacitor c=0.0146822f \
 //x=51.075 //y=1.655 //x2=59.085 //y2=2.22
cc_4029 ( N_noxref_15_c_5226_n N_SN_c_6866_n ) capacitor c=0.0217395f \
 //x=51.43 //y=2.59 //x2=59.085 //y2=2.22
cc_4030 ( N_noxref_15_c_5228_n N_SN_c_6866_n ) capacitor c=0.0211309f \
 //x=53.28 //y=2.08 //x2=59.085 //y2=2.22
cc_4031 ( N_noxref_15_c_5229_n N_SN_c_6866_n ) capacitor c=0.021104f //x=58.09 \
 //y=2.08 //x2=59.085 //y2=2.22
cc_4032 ( N_noxref_15_c_5234_n N_SN_c_6866_n ) capacitor c=0.011987f //x=52.98 \
 //y=1.915 //x2=59.085 //y2=2.22
cc_4033 ( N_noxref_15_c_5244_n N_SN_c_6866_n ) capacitor c=0.011987f //x=57.79 \
 //y=1.915 //x2=59.085 //y2=2.22
cc_4034 ( N_noxref_15_c_5229_n N_SN_c_6887_n ) capacitor c=0.00165648f \
 //x=58.09 //y=2.08 //x2=59.315 //y2=2.22
cc_4035 ( N_noxref_15_c_5244_n N_SN_c_6887_n ) capacitor c=2.3323e-19 \
 //x=57.79 //y=1.915 //x2=59.315 //y2=2.22
cc_4036 ( N_noxref_15_c_5223_n N_SN_c_6892_n ) capacitor c=0.00311593f \
 //x=57.975 //y=2.59 //x2=59.2 //y2=2.08
cc_4037 ( N_noxref_15_c_5229_n N_SN_c_6892_n ) capacitor c=0.0428203f \
 //x=58.09 //y=2.08 //x2=59.2 //y2=2.08
cc_4038 ( N_noxref_15_c_5244_n N_SN_c_6892_n ) capacitor c=0.00208635f \
 //x=57.79 //y=1.915 //x2=59.2 //y2=2.08
cc_4039 ( N_noxref_15_c_5315_p N_SN_c_6892_n ) capacitor c=0.00147352f \
 //x=58.655 //y=4.79 //x2=59.2 //y2=2.08
cc_4040 ( N_noxref_15_c_5280_n N_SN_c_6892_n ) capacitor c=0.00142741f \
 //x=58.365 //y=4.79 //x2=59.2 //y2=2.08
cc_4041 ( N_noxref_15_M122_noxref_g N_SN_M124_noxref_g ) capacitor \
 c=0.0105869f //x=58.29 //y=6.02 //x2=59.17 //y2=6.02
cc_4042 ( N_noxref_15_M123_noxref_g N_SN_M124_noxref_g ) capacitor c=0.10632f \
 //x=58.73 //y=6.02 //x2=59.17 //y2=6.02
cc_4043 ( N_noxref_15_M123_noxref_g N_SN_M125_noxref_g ) capacitor \
 c=0.0101598f //x=58.73 //y=6.02 //x2=59.61 //y2=6.02
cc_4044 ( N_noxref_15_c_5240_n N_SN_c_7244_n ) capacitor c=5.72482e-19 \
 //x=57.79 //y=0.875 //x2=58.765 //y2=0.91
cc_4045 ( N_noxref_15_c_5242_n N_SN_c_7244_n ) capacitor c=0.00149976f \
 //x=57.79 //y=1.22 //x2=58.765 //y2=0.91
cc_4046 ( N_noxref_15_c_5247_n N_SN_c_7244_n ) capacitor c=0.0160123f \
 //x=58.32 //y=0.875 //x2=58.765 //y2=0.91
cc_4047 ( N_noxref_15_c_5243_n N_SN_c_7247_n ) capacitor c=0.00111227f \
 //x=57.79 //y=1.53 //x2=58.765 //y2=1.22
cc_4048 ( N_noxref_15_c_5249_n N_SN_c_7247_n ) capacitor c=0.0124075f \
 //x=58.32 //y=1.22 //x2=58.765 //y2=1.22
cc_4049 ( N_noxref_15_c_5247_n N_SN_c_7249_n ) capacitor c=0.00103227f \
 //x=58.32 //y=0.875 //x2=59.29 //y2=0.91
cc_4050 ( N_noxref_15_c_5249_n N_SN_c_7250_n ) capacitor c=0.0010154f \
 //x=58.32 //y=1.22 //x2=59.29 //y2=1.22
cc_4051 ( N_noxref_15_c_5249_n N_SN_c_7251_n ) capacitor c=9.23422e-19 \
 //x=58.32 //y=1.22 //x2=59.29 //y2=1.45
cc_4052 ( N_noxref_15_c_5229_n N_SN_c_7252_n ) capacitor c=0.00203769f \
 //x=58.09 //y=2.08 //x2=59.29 //y2=1.915
cc_4053 ( N_noxref_15_c_5244_n N_SN_c_7252_n ) capacitor c=0.00834532f \
 //x=57.79 //y=1.915 //x2=59.29 //y2=1.915
cc_4054 ( N_noxref_15_c_5229_n N_SN_c_7254_n ) capacitor c=0.00183762f \
 //x=58.09 //y=2.08 //x2=59.2 //y2=4.7
cc_4055 ( N_noxref_15_c_5315_p N_SN_c_7254_n ) capacitor c=0.0168581f \
 //x=58.655 //y=4.79 //x2=59.2 //y2=4.7
cc_4056 ( N_noxref_15_c_5280_n N_SN_c_7254_n ) capacitor c=0.00484466f \
 //x=58.365 //y=4.79 //x2=59.2 //y2=4.7
cc_4057 ( N_noxref_15_c_5229_n N_noxref_21_c_7696_n ) capacitor c=0.0197627f \
 //x=58.09 //y=2.08 //x2=60.195 //y2=3.7
cc_4058 ( N_noxref_15_c_5223_n N_noxref_21_c_7648_n ) capacitor c=0.0179628f \
 //x=57.975 //y=2.59 //x2=55.5 //y2=2.08
cc_4059 ( N_noxref_15_c_5228_n N_noxref_21_c_7648_n ) capacitor c=0.00108806f \
 //x=53.28 //y=2.08 //x2=55.5 //y2=2.08
cc_4060 ( N_noxref_15_c_5229_n N_noxref_21_c_7648_n ) capacitor c=5.77326e-19 \
 //x=58.09 //y=2.08 //x2=55.5 //y2=2.08
cc_4061 ( N_noxref_15_c_5229_n N_noxref_21_c_7649_n ) capacitor c=0.00102099f \
 //x=58.09 //y=2.08 //x2=60.31 //y2=2.08
cc_4062 ( N_noxref_15_c_5221_n N_noxref_24_c_8424_n ) capacitor c=0.0111379f \
 //x=53.135 //y=2.59 //x2=79.065 //y2=3.33
cc_4063 ( N_noxref_15_c_5222_n N_noxref_24_c_8424_n ) capacitor c=8.86511e-19 \
 //x=51.545 //y=2.59 //x2=79.065 //y2=3.33
cc_4064 ( N_noxref_15_c_5223_n N_noxref_24_c_8424_n ) capacitor c=7.63975e-19 \
 //x=57.975 //y=2.59 //x2=79.065 //y2=3.33
cc_4065 ( N_noxref_15_c_5224_n N_noxref_24_c_8424_n ) capacitor c=0.036868f \
 //x=53.545 //y=2.59 //x2=79.065 //y2=3.33
cc_4066 ( N_noxref_15_c_5226_n N_noxref_24_c_8424_n ) capacitor c=0.0211091f \
 //x=51.43 //y=2.59 //x2=79.065 //y2=3.33
cc_4067 ( N_noxref_15_c_5228_n N_noxref_24_c_8424_n ) capacitor c=0.0221447f \
 //x=53.28 //y=2.08 //x2=79.065 //y2=3.33
cc_4068 ( N_noxref_15_c_5229_n N_noxref_24_c_8424_n ) capacitor c=0.0197803f \
 //x=58.09 //y=2.08 //x2=79.065 //y2=3.33
cc_4069 ( N_noxref_15_c_5389_p N_noxref_45_c_10172_n ) capacitor c=3.15806e-19 \
 //x=51.075 //y=1.655 //x2=49.535 //y2=1.495
cc_4070 ( N_noxref_15_c_5389_p N_noxref_45_c_10161_n ) capacitor c=0.020324f \
 //x=51.075 //y=1.655 //x2=50.505 //y2=1.495
cc_4071 ( N_noxref_15_c_5225_n N_noxref_45_c_10162_n ) capacitor c=0.00457164f \
 //x=51.345 //y=1.655 //x2=51.39 //y2=0.53
cc_4072 ( N_noxref_15_M31_noxref_d N_noxref_45_c_10162_n ) capacitor \
 c=0.0115831f //x=50.8 //y=0.905 //x2=51.39 //y2=0.53
cc_4073 ( N_noxref_15_c_5225_n N_noxref_45_M30_noxref_s ) capacitor \
 c=0.0126484f //x=51.345 //y=1.655 //x2=49.4 //y2=0.365
cc_4074 ( N_noxref_15_M31_noxref_d N_noxref_45_M30_noxref_s ) capacitor \
 c=0.0439476f //x=50.8 //y=0.905 //x2=49.4 //y2=0.365
cc_4075 ( N_noxref_15_c_5225_n N_noxref_46_c_10220_n ) capacitor c=4.08644e-19 \
 //x=51.345 //y=1.655 //x2=52.76 //y2=1.505
cc_4076 ( N_noxref_15_c_5234_n N_noxref_46_c_10220_n ) capacitor c=0.0034165f \
 //x=52.98 //y=1.915 //x2=52.76 //y2=1.505
cc_4077 ( N_noxref_15_c_5228_n N_noxref_46_c_10205_n ) capacitor c=0.0115578f \
 //x=53.28 //y=2.08 //x2=53.645 //y2=1.59
cc_4078 ( N_noxref_15_c_5233_n N_noxref_46_c_10205_n ) capacitor c=0.00697148f \
 //x=52.98 //y=1.53 //x2=53.645 //y2=1.59
cc_4079 ( N_noxref_15_c_5234_n N_noxref_46_c_10205_n ) capacitor c=0.0204849f \
 //x=52.98 //y=1.915 //x2=53.645 //y2=1.59
cc_4080 ( N_noxref_15_c_5236_n N_noxref_46_c_10205_n ) capacitor c=0.00610316f \
 //x=53.355 //y=1.375 //x2=53.645 //y2=1.59
cc_4081 ( N_noxref_15_c_5239_n N_noxref_46_c_10205_n ) capacitor c=0.00698822f \
 //x=53.51 //y=1.22 //x2=53.645 //y2=1.59
cc_4082 ( N_noxref_15_c_5230_n N_noxref_46_M32_noxref_s ) capacitor \
 c=0.0327271f //x=52.98 //y=0.875 //x2=52.625 //y2=0.375
cc_4083 ( N_noxref_15_c_5233_n N_noxref_46_M32_noxref_s ) capacitor \
 c=7.99997e-19 //x=52.98 //y=1.53 //x2=52.625 //y2=0.375
cc_4084 ( N_noxref_15_c_5234_n N_noxref_46_M32_noxref_s ) capacitor \
 c=0.00122123f //x=52.98 //y=1.915 //x2=52.625 //y2=0.375
cc_4085 ( N_noxref_15_c_5237_n N_noxref_46_M32_noxref_s ) capacitor \
 c=0.0121427f //x=53.51 //y=0.875 //x2=52.625 //y2=0.375
cc_4086 ( N_noxref_15_M31_noxref_d N_noxref_46_M32_noxref_s ) capacitor \
 c=2.53688e-19 //x=50.8 //y=0.905 //x2=52.625 //y2=0.375
cc_4087 ( N_noxref_15_c_5244_n N_noxref_48_c_10321_n ) capacitor c=0.0034165f \
 //x=57.79 //y=1.915 //x2=57.57 //y2=1.505
cc_4088 ( N_noxref_15_c_5229_n N_noxref_48_c_10306_n ) capacitor c=0.0115578f \
 //x=58.09 //y=2.08 //x2=58.455 //y2=1.59
cc_4089 ( N_noxref_15_c_5243_n N_noxref_48_c_10306_n ) capacitor c=0.00697148f \
 //x=57.79 //y=1.53 //x2=58.455 //y2=1.59
cc_4090 ( N_noxref_15_c_5244_n N_noxref_48_c_10306_n ) capacitor c=0.0204849f \
 //x=57.79 //y=1.915 //x2=58.455 //y2=1.59
cc_4091 ( N_noxref_15_c_5246_n N_noxref_48_c_10306_n ) capacitor c=0.00610316f \
 //x=58.165 //y=1.375 //x2=58.455 //y2=1.59
cc_4092 ( N_noxref_15_c_5249_n N_noxref_48_c_10306_n ) capacitor c=0.00698822f \
 //x=58.32 //y=1.22 //x2=58.455 //y2=1.59
cc_4093 ( N_noxref_15_c_5240_n N_noxref_48_M35_noxref_s ) capacitor \
 c=0.0327271f //x=57.79 //y=0.875 //x2=57.435 //y2=0.375
cc_4094 ( N_noxref_15_c_5243_n N_noxref_48_M35_noxref_s ) capacitor \
 c=7.99997e-19 //x=57.79 //y=1.53 //x2=57.435 //y2=0.375
cc_4095 ( N_noxref_15_c_5244_n N_noxref_48_M35_noxref_s ) capacitor \
 c=0.00122123f //x=57.79 //y=1.915 //x2=57.435 //y2=0.375
cc_4096 ( N_noxref_15_c_5247_n N_noxref_48_M35_noxref_s ) capacitor \
 c=0.0121427f //x=58.32 //y=0.875 //x2=57.435 //y2=0.375
cc_4097 ( N_noxref_16_c_5474_n N_CLK_c_5705_n ) capacitor c=0.032141f \
 //x=59.305 //y=5.155 //x2=63.525 //y2=4.44
cc_4098 ( N_noxref_16_c_5478_n N_CLK_c_5705_n ) capacitor c=0.0230136f \
 //x=58.595 //y=5.155 //x2=63.525 //y2=4.44
cc_4099 ( N_noxref_16_c_5484_n N_CLK_c_5705_n ) capacitor c=0.0183122f \
 //x=60.965 //y=5.155 //x2=63.525 //y2=4.44
cc_4100 ( N_noxref_16_c_5461_n N_CLK_c_5705_n ) capacitor c=0.0210274f \
 //x=61.05 //y=2.59 //x2=63.525 //y2=4.44
cc_4101 ( N_noxref_16_c_5462_n N_CLK_c_5705_n ) capacitor c=0.0215137f \
 //x=62.9 //y=2.08 //x2=63.525 //y2=4.44
cc_4102 ( N_noxref_16_c_5496_n N_CLK_c_5705_n ) capacitor c=0.0109968f \
 //x=62.9 //y=4.7 //x2=63.525 //y2=4.44
cc_4103 ( N_noxref_16_c_5462_n N_CLK_c_6133_n ) capacitor c=0.00400249f \
 //x=62.9 //y=2.08 //x2=63.64 //y2=4.535
cc_4104 ( N_noxref_16_c_5496_n N_CLK_c_6133_n ) capacitor c=0.00415951f \
 //x=62.9 //y=4.7 //x2=63.64 //y2=4.535
cc_4105 ( N_noxref_16_c_5458_n N_CLK_c_5629_n ) capacitor c=0.00720056f \
 //x=62.785 //y=2.59 //x2=63.64 //y2=2.08
cc_4106 ( N_noxref_16_c_5461_n N_CLK_c_5629_n ) capacitor c=6.41343e-19 \
 //x=61.05 //y=2.59 //x2=63.64 //y2=2.08
cc_4107 ( N_noxref_16_c_5462_n N_CLK_c_5629_n ) capacitor c=0.0712948f \
 //x=62.9 //y=2.08 //x2=63.64 //y2=2.08
cc_4108 ( N_noxref_16_c_5467_n N_CLK_c_5629_n ) capacitor c=0.00284029f \
 //x=62.705 //y=1.915 //x2=63.64 //y2=2.08
cc_4109 ( N_noxref_16_M128_noxref_g N_CLK_M130_noxref_g ) capacitor \
 c=0.0104611f //x=62.8 //y=6.02 //x2=63.68 //y2=6.02
cc_4110 ( N_noxref_16_M129_noxref_g N_CLK_M130_noxref_g ) capacitor \
 c=0.106811f //x=63.24 //y=6.02 //x2=63.68 //y2=6.02
cc_4111 ( N_noxref_16_M129_noxref_g N_CLK_M131_noxref_g ) capacitor \
 c=0.0100341f //x=63.24 //y=6.02 //x2=64.12 //y2=6.02
cc_4112 ( N_noxref_16_c_5463_n N_CLK_c_6142_n ) capacitor c=4.86506e-19 \
 //x=62.705 //y=0.865 //x2=63.675 //y2=0.905
cc_4113 ( N_noxref_16_c_5465_n N_CLK_c_6142_n ) capacitor c=0.00152104f \
 //x=62.705 //y=1.21 //x2=63.675 //y2=0.905
cc_4114 ( N_noxref_16_c_5470_n N_CLK_c_6142_n ) capacitor c=0.0151475f \
 //x=63.235 //y=0.865 //x2=63.675 //y2=0.905
cc_4115 ( N_noxref_16_c_5466_n N_CLK_c_6145_n ) capacitor c=0.00109982f \
 //x=62.705 //y=1.52 //x2=63.675 //y2=1.25
cc_4116 ( N_noxref_16_c_5472_n N_CLK_c_6145_n ) capacitor c=0.0111064f \
 //x=63.235 //y=1.21 //x2=63.675 //y2=1.25
cc_4117 ( N_noxref_16_c_5466_n N_CLK_c_6147_n ) capacitor c=9.57794e-19 \
 //x=62.705 //y=1.52 //x2=63.675 //y2=1.56
cc_4118 ( N_noxref_16_c_5467_n N_CLK_c_6147_n ) capacitor c=0.00662747f \
 //x=62.705 //y=1.915 //x2=63.675 //y2=1.56
cc_4119 ( N_noxref_16_c_5472_n N_CLK_c_6147_n ) capacitor c=0.00862358f \
 //x=63.235 //y=1.21 //x2=63.675 //y2=1.56
cc_4120 ( N_noxref_16_c_5470_n N_CLK_c_6150_n ) capacitor c=0.00124821f \
 //x=63.235 //y=0.865 //x2=64.205 //y2=0.905
cc_4121 ( N_noxref_16_c_5472_n N_CLK_c_6151_n ) capacitor c=0.00200715f \
 //x=63.235 //y=1.21 //x2=64.205 //y2=1.25
cc_4122 ( N_noxref_16_c_5462_n N_CLK_c_6152_n ) capacitor c=0.00282278f \
 //x=62.9 //y=2.08 //x2=63.64 //y2=2.08
cc_4123 ( N_noxref_16_c_5467_n N_CLK_c_6152_n ) capacitor c=0.0172771f \
 //x=62.705 //y=1.915 //x2=63.64 //y2=2.08
cc_4124 ( N_noxref_16_c_5462_n N_CLK_c_6154_n ) capacitor c=0.00342116f \
 //x=62.9 //y=2.08 //x2=63.67 //y2=4.7
cc_4125 ( N_noxref_16_c_5496_n N_CLK_c_6154_n ) capacitor c=0.0292158f \
 //x=62.9 //y=4.7 //x2=63.67 //y2=4.7
cc_4126 ( N_noxref_16_c_5461_n N_noxref_18_c_6393_n ) capacitor c=0.0181982f \
 //x=61.05 //y=2.59 //x2=66.115 //y2=4.07
cc_4127 ( N_noxref_16_c_5462_n N_noxref_18_c_6393_n ) capacitor c=0.0184765f \
 //x=62.9 //y=2.08 //x2=66.115 //y2=4.07
cc_4128 ( N_noxref_16_c_5478_n N_noxref_18_c_6415_n ) capacitor c=3.10026e-19 \
 //x=58.595 //y=5.155 //x2=56.155 //y2=5.155
cc_4129 ( N_noxref_16_c_5458_n N_SN_c_6877_n ) capacitor c=0.172308f \
 //x=62.785 //y=2.59 //x2=70.555 //y2=2.22
cc_4130 ( N_noxref_16_c_5459_n N_SN_c_6877_n ) capacitor c=0.0291301f \
 //x=61.165 //y=2.59 //x2=70.555 //y2=2.22
cc_4131 ( N_noxref_16_c_5555_p N_SN_c_6877_n ) capacitor c=0.016327f //x=60.65 \
 //y=1.665 //x2=70.555 //y2=2.22
cc_4132 ( N_noxref_16_c_5461_n N_SN_c_6877_n ) capacitor c=0.0215653f \
 //x=61.05 //y=2.59 //x2=70.555 //y2=2.22
cc_4133 ( N_noxref_16_c_5462_n N_SN_c_6877_n ) capacitor c=0.0203358f //x=62.9 \
 //y=2.08 //x2=70.555 //y2=2.22
cc_4134 ( N_noxref_16_c_5467_n N_SN_c_6877_n ) capacitor c=0.00894156f \
 //x=62.705 //y=1.915 //x2=70.555 //y2=2.22
cc_4135 ( N_noxref_16_c_5474_n N_SN_c_6892_n ) capacitor c=0.0146f //x=59.305 \
 //y=5.155 //x2=59.2 //y2=2.08
cc_4136 ( N_noxref_16_c_5461_n N_SN_c_6892_n ) capacitor c=0.00237834f \
 //x=61.05 //y=2.59 //x2=59.2 //y2=2.08
cc_4137 ( N_noxref_16_c_5474_n N_SN_M124_noxref_g ) capacitor c=0.0165266f \
 //x=59.305 //y=5.155 //x2=59.17 //y2=6.02
cc_4138 ( N_noxref_16_M124_noxref_d N_SN_M124_noxref_g ) capacitor \
 c=0.0180032f //x=59.245 //y=5.02 //x2=59.17 //y2=6.02
cc_4139 ( N_noxref_16_c_5480_n N_SN_M125_noxref_g ) capacitor c=0.01736f \
 //x=60.185 //y=5.155 //x2=59.61 //y2=6.02
cc_4140 ( N_noxref_16_M124_noxref_d N_SN_M125_noxref_g ) capacitor \
 c=0.0180032f //x=59.245 //y=5.02 //x2=59.61 //y2=6.02
cc_4141 ( N_noxref_16_c_5565_p N_SN_c_7269_n ) capacitor c=0.00426767f \
 //x=59.39 //y=5.155 //x2=59.535 //y2=4.79
cc_4142 ( N_noxref_16_c_5474_n N_SN_c_7254_n ) capacitor c=0.00322054f \
 //x=59.305 //y=5.155 //x2=59.2 //y2=4.7
cc_4143 ( N_noxref_16_c_5461_n N_noxref_21_c_7698_n ) capacitor c=0.0187698f \
 //x=61.05 //y=2.59 //x2=64.265 //y2=3.7
cc_4144 ( N_noxref_16_c_5462_n N_noxref_21_c_7698_n ) capacitor c=0.0187484f \
 //x=62.9 //y=2.08 //x2=64.265 //y2=3.7
cc_4145 ( N_noxref_16_c_5461_n N_noxref_21_c_7699_n ) capacitor c=0.00117715f \
 //x=61.05 //y=2.59 //x2=60.425 //y2=3.7
cc_4146 ( N_noxref_16_c_5459_n N_noxref_21_c_7649_n ) capacitor c=0.00456439f \
 //x=61.165 //y=2.59 //x2=60.31 //y2=2.08
cc_4147 ( N_noxref_16_c_5461_n N_noxref_21_c_7649_n ) capacitor c=0.076937f \
 //x=61.05 //y=2.59 //x2=60.31 //y2=2.08
cc_4148 ( N_noxref_16_c_5462_n N_noxref_21_c_7649_n ) capacitor c=5.32619e-19 \
 //x=62.9 //y=2.08 //x2=60.31 //y2=2.08
cc_4149 ( N_noxref_16_c_5573_p N_noxref_21_c_7649_n ) capacitor c=0.016476f \
 //x=60.27 //y=5.155 //x2=60.31 //y2=2.08
cc_4150 ( N_noxref_16_M129_noxref_g N_noxref_21_c_7660_n ) capacitor \
 c=0.0169521f //x=63.24 //y=6.02 //x2=63.815 //y2=5.2
cc_4151 ( N_noxref_16_c_5462_n N_noxref_21_c_7664_n ) capacitor c=0.00539951f \
 //x=62.9 //y=2.08 //x2=63.105 //y2=5.2
cc_4152 ( N_noxref_16_M128_noxref_g N_noxref_21_c_7664_n ) capacitor \
 c=0.0177326f //x=62.8 //y=6.02 //x2=63.105 //y2=5.2
cc_4153 ( N_noxref_16_c_5496_n N_noxref_21_c_7664_n ) capacitor c=0.00581252f \
 //x=62.9 //y=4.7 //x2=63.105 //y2=5.2
cc_4154 ( N_noxref_16_c_5461_n N_noxref_21_c_7651_n ) capacitor c=3.52729e-19 \
 //x=61.05 //y=2.59 //x2=64.38 //y2=3.7
cc_4155 ( N_noxref_16_c_5462_n N_noxref_21_c_7651_n ) capacitor c=0.00321436f \
 //x=62.9 //y=2.08 //x2=64.38 //y2=3.7
cc_4156 ( N_noxref_16_c_5480_n N_noxref_21_M126_noxref_g ) capacitor \
 c=0.01736f //x=60.185 //y=5.155 //x2=60.05 //y2=6.02
cc_4157 ( N_noxref_16_M126_noxref_d N_noxref_21_M126_noxref_g ) capacitor \
 c=0.0180032f //x=60.125 //y=5.02 //x2=60.05 //y2=6.02
cc_4158 ( N_noxref_16_c_5484_n N_noxref_21_M127_noxref_g ) capacitor \
 c=0.0194981f //x=60.965 //y=5.155 //x2=60.49 //y2=6.02
cc_4159 ( N_noxref_16_M126_noxref_d N_noxref_21_M127_noxref_g ) capacitor \
 c=0.0194246f //x=60.125 //y=5.02 //x2=60.49 //y2=6.02
cc_4160 ( N_noxref_16_M37_noxref_d N_noxref_21_c_7729_n ) capacitor \
 c=0.00217566f //x=60.375 //y=0.915 //x2=60.3 //y2=0.915
cc_4161 ( N_noxref_16_M37_noxref_d N_noxref_21_c_7730_n ) capacitor \
 c=0.0034598f //x=60.375 //y=0.915 //x2=60.3 //y2=1.26
cc_4162 ( N_noxref_16_M37_noxref_d N_noxref_21_c_7731_n ) capacitor \
 c=0.00546784f //x=60.375 //y=0.915 //x2=60.3 //y2=1.57
cc_4163 ( N_noxref_16_M37_noxref_d N_noxref_21_c_7732_n ) capacitor \
 c=0.00241102f //x=60.375 //y=0.915 //x2=60.675 //y2=0.76
cc_4164 ( N_noxref_16_c_5460_n N_noxref_21_c_7733_n ) capacitor c=0.00371277f \
 //x=60.965 //y=1.665 //x2=60.675 //y2=1.415
cc_4165 ( N_noxref_16_M37_noxref_d N_noxref_21_c_7733_n ) capacitor \
 c=0.0138621f //x=60.375 //y=0.915 //x2=60.675 //y2=1.415
cc_4166 ( N_noxref_16_M37_noxref_d N_noxref_21_c_7735_n ) capacitor \
 c=0.00219619f //x=60.375 //y=0.915 //x2=60.83 //y2=0.915
cc_4167 ( N_noxref_16_c_5460_n N_noxref_21_c_7736_n ) capacitor c=0.00457401f \
 //x=60.965 //y=1.665 //x2=60.83 //y2=1.26
cc_4168 ( N_noxref_16_M37_noxref_d N_noxref_21_c_7736_n ) capacitor \
 c=0.00603828f //x=60.375 //y=0.915 //x2=60.83 //y2=1.26
cc_4169 ( N_noxref_16_c_5461_n N_noxref_21_c_7738_n ) capacitor c=0.00709342f \
 //x=61.05 //y=2.59 //x2=60.31 //y2=2.08
cc_4170 ( N_noxref_16_c_5461_n N_noxref_21_c_7739_n ) capacitor c=0.00283672f \
 //x=61.05 //y=2.59 //x2=60.31 //y2=1.915
cc_4171 ( N_noxref_16_M37_noxref_d N_noxref_21_c_7739_n ) capacitor \
 c=0.00661782f //x=60.375 //y=0.915 //x2=60.31 //y2=1.915
cc_4172 ( N_noxref_16_c_5484_n N_noxref_21_c_7741_n ) capacitor c=0.00201851f \
 //x=60.965 //y=5.155 //x2=60.31 //y2=4.7
cc_4173 ( N_noxref_16_c_5461_n N_noxref_21_c_7741_n ) capacitor c=0.013693f \
 //x=61.05 //y=2.59 //x2=60.31 //y2=4.7
cc_4174 ( N_noxref_16_c_5573_p N_noxref_21_c_7741_n ) capacitor c=0.00475601f \
 //x=60.27 //y=5.155 //x2=60.31 //y2=4.7
cc_4175 ( N_noxref_16_M129_noxref_g N_noxref_21_M128_noxref_d ) capacitor \
 c=0.0173476f //x=63.24 //y=6.02 //x2=62.875 //y2=5.02
cc_4176 ( N_noxref_16_c_5458_n N_noxref_24_c_8424_n ) capacitor c=0.0125435f \
 //x=62.785 //y=2.59 //x2=79.065 //y2=3.33
cc_4177 ( N_noxref_16_c_5459_n N_noxref_24_c_8424_n ) capacitor c=8.87672e-19 \
 //x=61.165 //y=2.59 //x2=79.065 //y2=3.33
cc_4178 ( N_noxref_16_c_5461_n N_noxref_24_c_8424_n ) capacitor c=0.018769f \
 //x=61.05 //y=2.59 //x2=79.065 //y2=3.33
cc_4179 ( N_noxref_16_c_5462_n N_noxref_24_c_8424_n ) capacitor c=0.0187666f \
 //x=62.9 //y=2.08 //x2=79.065 //y2=3.33
cc_4180 ( N_noxref_16_M37_noxref_d N_noxref_48_M35_noxref_s ) capacitor \
 c=0.00309936f //x=60.375 //y=0.915 //x2=57.435 //y2=0.375
cc_4181 ( N_noxref_16_c_5460_n N_noxref_49_c_10363_n ) capacitor c=0.00457167f \
 //x=60.965 //y=1.665 //x2=60.965 //y2=0.54
cc_4182 ( N_noxref_16_M37_noxref_d N_noxref_49_c_10363_n ) capacitor \
 c=0.0115903f //x=60.375 //y=0.915 //x2=60.965 //y2=0.54
cc_4183 ( N_noxref_16_c_5555_p N_noxref_49_c_10373_n ) capacitor c=0.020048f \
 //x=60.65 //y=1.665 //x2=60.08 //y2=0.995
cc_4184 ( N_noxref_16_M37_noxref_d N_noxref_49_M36_noxref_d ) capacitor \
 c=5.27807e-19 //x=60.375 //y=0.915 //x2=58.84 //y2=0.91
cc_4185 ( N_noxref_16_c_5460_n N_noxref_49_M37_noxref_s ) capacitor \
 c=0.0184051f //x=60.965 //y=1.665 //x2=59.945 //y2=0.375
cc_4186 ( N_noxref_16_M37_noxref_d N_noxref_49_M37_noxref_s ) capacitor \
 c=0.0426444f //x=60.375 //y=0.915 //x2=59.945 //y2=0.375
cc_4187 ( N_noxref_16_c_5460_n N_noxref_50_c_10428_n ) capacitor c=3.04182e-19 \
 //x=60.965 //y=1.665 //x2=62.485 //y2=1.495
cc_4188 ( N_noxref_16_c_5467_n N_noxref_50_c_10428_n ) capacitor c=0.0034165f \
 //x=62.705 //y=1.915 //x2=62.485 //y2=1.495
cc_4189 ( N_noxref_16_c_5462_n N_noxref_50_c_10410_n ) capacitor c=0.0111916f \
 //x=62.9 //y=2.08 //x2=63.37 //y2=1.58
cc_4190 ( N_noxref_16_c_5466_n N_noxref_50_c_10410_n ) capacitor c=0.00696403f \
 //x=62.705 //y=1.52 //x2=63.37 //y2=1.58
cc_4191 ( N_noxref_16_c_5467_n N_noxref_50_c_10410_n ) capacitor c=0.0174694f \
 //x=62.705 //y=1.915 //x2=63.37 //y2=1.58
cc_4192 ( N_noxref_16_c_5469_n N_noxref_50_c_10410_n ) capacitor c=0.00776811f \
 //x=63.08 //y=1.365 //x2=63.37 //y2=1.58
cc_4193 ( N_noxref_16_c_5472_n N_noxref_50_c_10410_n ) capacitor c=0.00339872f \
 //x=63.235 //y=1.21 //x2=63.37 //y2=1.58
cc_4194 ( N_noxref_16_c_5467_n N_noxref_50_c_10417_n ) capacitor c=6.71402e-19 \
 //x=62.705 //y=1.915 //x2=63.455 //y2=1.495
cc_4195 ( N_noxref_16_c_5463_n N_noxref_50_M38_noxref_s ) capacitor \
 c=0.0327502f //x=62.705 //y=0.865 //x2=62.35 //y2=0.365
cc_4196 ( N_noxref_16_c_5466_n N_noxref_50_M38_noxref_s ) capacitor \
 c=3.48408e-19 //x=62.705 //y=1.52 //x2=62.35 //y2=0.365
cc_4197 ( N_noxref_16_c_5470_n N_noxref_50_M38_noxref_s ) capacitor \
 c=0.0120759f //x=63.235 //y=0.865 //x2=62.35 //y2=0.365
cc_4198 ( N_CLK_c_5680_n N_noxref_18_c_6392_n ) capacitor c=0.302855f \
 //x=54.275 //y=4.44 //x2=56.12 //y2=4.07
cc_4199 ( N_CLK_c_5705_n N_noxref_18_c_6392_n ) capacitor c=0.139602f \
 //x=63.525 //y=4.44 //x2=56.12 //y2=4.07
cc_4200 ( N_CLK_c_5716_n N_noxref_18_c_6392_n ) capacitor c=0.026534f \
 //x=54.505 //y=4.44 //x2=56.12 //y2=4.07
cc_4201 ( N_CLK_c_5628_n N_noxref_18_c_6392_n ) capacitor c=0.0231929f \
 //x=54.39 //y=2.08 //x2=56.12 //y2=4.07
cc_4202 ( N_CLK_c_5680_n N_noxref_18_c_6449_n ) capacitor c=0.028941f \
 //x=54.275 //y=4.44 //x2=50.805 //y2=4.07
cc_4203 ( N_CLK_c_5705_n N_noxref_18_c_6393_n ) capacitor c=0.654862f \
 //x=63.525 //y=4.44 //x2=66.115 //y2=4.07
cc_4204 ( N_CLK_c_5629_n N_noxref_18_c_6393_n ) capacitor c=0.0187718f \
 //x=63.64 //y=2.08 //x2=66.115 //y2=4.07
cc_4205 ( N_CLK_c_6163_p N_noxref_18_c_6393_n ) capacitor c=0.00756255f \
 //x=64.045 //y=4.79 //x2=66.115 //y2=4.07
cc_4206 ( N_CLK_c_6154_n N_noxref_18_c_6393_n ) capacitor c=4.6185e-19 \
 //x=63.67 //y=4.7 //x2=66.115 //y2=4.07
cc_4207 ( N_CLK_c_5705_n N_noxref_18_c_6402_n ) capacitor c=0.0265302f \
 //x=63.525 //y=4.44 //x2=56.35 //y2=4.07
cc_4208 ( N_CLK_c_5680_n N_noxref_18_c_6458_n ) capacitor c=0.0016972f \
 //x=54.275 //y=4.44 //x2=50.69 //y2=4.535
cc_4209 ( N_CLK_c_5680_n N_noxref_18_c_6377_n ) capacitor c=0.0207534f \
 //x=54.275 //y=4.44 //x2=50.69 //y2=2.08
cc_4210 ( N_CLK_c_5716_n N_noxref_18_c_6405_n ) capacitor c=0.00241768f \
 //x=54.505 //y=4.44 //x2=54.495 //y2=5.155
cc_4211 ( N_CLK_c_5628_n N_noxref_18_c_6405_n ) capacitor c=0.014564f \
 //x=54.39 //y=2.08 //x2=54.495 //y2=5.155
cc_4212 ( N_CLK_M118_noxref_g N_noxref_18_c_6405_n ) capacitor c=0.016514f \
 //x=54.36 //y=6.02 //x2=54.495 //y2=5.155
cc_4213 ( N_CLK_c_6124_n N_noxref_18_c_6405_n ) capacitor c=0.00322046f \
 //x=54.39 //y=4.7 //x2=54.495 //y2=5.155
cc_4214 ( N_CLK_c_5680_n N_noxref_18_c_6409_n ) capacitor c=0.0219114f \
 //x=54.275 //y=4.44 //x2=53.785 //y2=5.155
cc_4215 ( N_CLK_M119_noxref_g N_noxref_18_c_6411_n ) capacitor c=0.01736f \
 //x=54.8 //y=6.02 //x2=55.375 //y2=5.155
cc_4216 ( N_CLK_c_5705_n N_noxref_18_c_6415_n ) capacitor c=0.0182691f \
 //x=63.525 //y=4.44 //x2=56.155 //y2=5.155
cc_4217 ( N_CLK_c_5705_n N_noxref_18_c_6539_n ) capacitor c=0.0207896f \
 //x=63.525 //y=4.44 //x2=56.24 //y2=5.07
cc_4218 ( N_CLK_c_5628_n N_noxref_18_c_6539_n ) capacitor c=7.17254e-19 \
 //x=54.39 //y=2.08 //x2=56.24 //y2=5.07
cc_4219 ( N_CLK_c_5629_n N_noxref_18_c_6380_n ) capacitor c=6.57265e-19 \
 //x=63.64 //y=2.08 //x2=66.23 //y2=2.08
cc_4220 ( N_CLK_c_5705_n N_noxref_18_c_6542_n ) capacitor c=0.0311227f \
 //x=63.525 //y=4.44 //x2=54.58 //y2=5.155
cc_4221 ( N_CLK_c_6179_p N_noxref_18_c_6542_n ) capacitor c=0.00426767f \
 //x=54.725 //y=4.79 //x2=54.58 //y2=5.155
cc_4222 ( N_CLK_c_5705_n N_noxref_18_c_6422_n ) capacitor c=0.00215288f \
 //x=63.525 //y=4.44 //x2=56.235 //y2=4.07
cc_4223 ( N_CLK_c_5628_n N_noxref_18_c_6456_n ) capacitor c=0.00157145f \
 //x=54.39 //y=2.08 //x2=56.237 //y2=3.905
cc_4224 ( N_CLK_c_5680_n N_noxref_18_c_6503_n ) capacitor c=0.00960248f \
 //x=54.275 //y=4.44 //x2=51.095 //y2=4.79
cc_4225 ( N_CLK_c_5680_n N_noxref_18_c_6478_n ) capacitor c=0.00203982f \
 //x=54.275 //y=4.44 //x2=50.72 //y2=4.7
cc_4226 ( N_CLK_M118_noxref_g N_noxref_18_M118_noxref_d ) capacitor \
 c=0.0180032f //x=54.36 //y=6.02 //x2=54.435 //y2=5.02
cc_4227 ( N_CLK_M119_noxref_g N_noxref_18_M118_noxref_d ) capacitor \
 c=0.0180032f //x=54.8 //y=6.02 //x2=54.435 //y2=5.02
cc_4228 ( N_CLK_c_5623_n N_SN_c_6833_n ) capacitor c=0.0201924f //x=14.8 \
 //y=2.08 //x2=21.715 //y2=2.22
cc_4229 ( N_CLK_c_5896_n N_SN_c_6833_n ) capacitor c=3.11115e-19 //x=15.21 \
 //y=1.405 //x2=21.715 //y2=2.22
cc_4230 ( N_CLK_c_5810_n N_SN_c_6833_n ) capacitor c=0.00568402f //x=14.8 \
 //y=2.08 //x2=21.715 //y2=2.22
cc_4231 ( N_CLK_c_5625_n N_SN_c_6844_n ) capacitor c=0.0193884f //x=29.97 \
 //y=2.08 //x2=34.665 //y2=2.22
cc_4232 ( N_CLK_c_5934_n N_SN_c_6844_n ) capacitor c=0.00583058f //x=30.06 \
 //y=1.915 //x2=34.665 //y2=2.22
cc_4233 ( N_CLK_c_5626_n N_SN_c_6855_n ) capacitor c=0.0201924f //x=39.22 \
 //y=2.08 //x2=46.135 //y2=2.22
cc_4234 ( N_CLK_c_6057_n N_SN_c_6855_n ) capacitor c=3.11115e-19 //x=39.63 \
 //y=1.405 //x2=46.135 //y2=2.22
cc_4235 ( N_CLK_c_5966_n N_SN_c_6855_n ) capacitor c=0.00568402f //x=39.22 \
 //y=2.08 //x2=46.135 //y2=2.22
cc_4236 ( N_CLK_c_5628_n N_SN_c_6866_n ) capacitor c=0.0193884f //x=54.39 \
 //y=2.08 //x2=59.085 //y2=2.22
cc_4237 ( N_CLK_c_6122_n N_SN_c_6866_n ) capacitor c=0.00583058f //x=54.48 \
 //y=1.915 //x2=59.085 //y2=2.22
cc_4238 ( N_CLK_c_5629_n N_SN_c_6877_n ) capacitor c=0.0201924f //x=63.64 \
 //y=2.08 //x2=70.555 //y2=2.22
cc_4239 ( N_CLK_c_6197_p N_SN_c_6877_n ) capacitor c=3.11115e-19 //x=64.05 \
 //y=1.405 //x2=70.555 //y2=2.22
cc_4240 ( N_CLK_c_6152_n N_SN_c_6877_n ) capacitor c=0.00568402f //x=63.64 \
 //y=2.08 //x2=70.555 //y2=2.22
cc_4241 ( N_CLK_c_5631_n N_SN_c_6888_n ) capacitor c=0.0210462f //x=14.685 \
 //y=4.44 //x2=10.36 //y2=2.08
cc_4242 ( N_CLK_c_5643_n N_SN_c_6889_n ) capacitor c=0.0233868f //x=29.855 \
 //y=4.44 //x2=21.83 //y2=2.08
cc_4243 ( N_CLK_c_5668_n N_SN_c_6890_n ) capacitor c=0.0210462f //x=39.105 \
 //y=4.44 //x2=34.78 //y2=2.08
cc_4244 ( N_CLK_c_5680_n N_SN_c_6891_n ) capacitor c=0.0210462f //x=54.275 \
 //y=4.44 //x2=46.25 //y2=2.08
cc_4245 ( N_CLK_c_5705_n N_SN_c_6892_n ) capacitor c=0.0210462f //x=63.525 \
 //y=4.44 //x2=59.2 //y2=2.08
cc_4246 ( N_CLK_c_5631_n N_SN_c_6965_n ) capacitor c=0.0085986f //x=14.685 \
 //y=4.44 //x2=10.695 //y2=4.79
cc_4247 ( N_CLK_c_5643_n N_SN_c_7045_n ) capacitor c=0.0085986f //x=29.855 \
 //y=4.44 //x2=22.165 //y2=4.79
cc_4248 ( N_CLK_c_5668_n N_SN_c_7095_n ) capacitor c=0.0085986f //x=39.105 \
 //y=4.44 //x2=35.115 //y2=4.79
cc_4249 ( N_CLK_c_5680_n N_SN_c_7179_n ) capacitor c=0.0085986f //x=54.275 \
 //y=4.44 //x2=46.585 //y2=4.79
cc_4250 ( N_CLK_c_5705_n N_SN_c_7269_n ) capacitor c=0.0085986f //x=63.525 \
 //y=4.44 //x2=59.535 //y2=4.79
cc_4251 ( N_CLK_c_5631_n N_SN_c_6950_n ) capacitor c=0.00293313f //x=14.685 \
 //y=4.44 //x2=10.36 //y2=4.7
cc_4252 ( N_CLK_c_5643_n N_SN_c_6996_n ) capacitor c=0.00293313f //x=29.855 \
 //y=4.44 //x2=21.83 //y2=4.7
cc_4253 ( N_CLK_c_5668_n N_SN_c_7080_n ) capacitor c=0.00293313f //x=39.105 \
 //y=4.44 //x2=34.78 //y2=4.7
cc_4254 ( N_CLK_c_5680_n N_SN_c_7133_n ) capacitor c=0.00293313f //x=54.275 \
 //y=4.44 //x2=46.25 //y2=4.7
cc_4255 ( N_CLK_c_5705_n N_SN_c_7254_n ) capacitor c=0.00293313f //x=63.525 \
 //y=4.44 //x2=59.2 //y2=4.7
cc_4256 ( N_CLK_c_5705_n N_noxref_21_c_7696_n ) capacitor c=0.0345106f \
 //x=63.525 //y=4.44 //x2=60.195 //y2=3.7
cc_4257 ( N_CLK_c_5705_n N_noxref_21_c_7697_n ) capacitor c=7.0371e-19 \
 //x=63.525 //y=4.44 //x2=55.615 //y2=3.7
cc_4258 ( N_CLK_c_5628_n N_noxref_21_c_7697_n ) capacitor c=0.00526349f \
 //x=54.39 //y=2.08 //x2=55.615 //y2=3.7
cc_4259 ( N_CLK_c_5705_n N_noxref_21_c_7698_n ) capacitor c=0.0218071f \
 //x=63.525 //y=4.44 //x2=64.265 //y2=3.7
cc_4260 ( N_CLK_c_5629_n N_noxref_21_c_7698_n ) capacitor c=0.0169594f \
 //x=63.64 //y=2.08 //x2=64.265 //y2=3.7
cc_4261 ( N_CLK_c_5705_n N_noxref_21_c_7699_n ) capacitor c=4.78625e-19 \
 //x=63.525 //y=4.44 //x2=60.425 //y2=3.7
cc_4262 ( N_CLK_c_5629_n N_noxref_21_c_7701_n ) capacitor c=0.00117715f \
 //x=63.64 //y=2.08 //x2=64.495 //y2=3.7
cc_4263 ( N_CLK_c_5705_n N_noxref_21_c_7648_n ) capacitor c=0.0200057f \
 //x=63.525 //y=4.44 //x2=55.5 //y2=2.08
cc_4264 ( N_CLK_c_5716_n N_noxref_21_c_7648_n ) capacitor c=0.00153281f \
 //x=54.505 //y=4.44 //x2=55.5 //y2=2.08
cc_4265 ( N_CLK_c_5628_n N_noxref_21_c_7648_n ) capacitor c=0.0422302f \
 //x=54.39 //y=2.08 //x2=55.5 //y2=2.08
cc_4266 ( N_CLK_c_6122_n N_noxref_21_c_7648_n ) capacitor c=0.00205895f \
 //x=54.48 //y=1.915 //x2=55.5 //y2=2.08
cc_4267 ( N_CLK_c_6124_n N_noxref_21_c_7648_n ) capacitor c=0.00142741f \
 //x=54.39 //y=4.7 //x2=55.5 //y2=2.08
cc_4268 ( N_CLK_c_5705_n N_noxref_21_c_7649_n ) capacitor c=0.0200057f \
 //x=63.525 //y=4.44 //x2=60.31 //y2=2.08
cc_4269 ( N_CLK_c_5705_n N_noxref_21_c_7660_n ) capacitor c=0.00325337f \
 //x=63.525 //y=4.44 //x2=63.815 //y2=5.2
cc_4270 ( N_CLK_c_6133_n N_noxref_21_c_7660_n ) capacitor c=0.0126974f \
 //x=63.64 //y=4.535 //x2=63.815 //y2=5.2
cc_4271 ( N_CLK_c_5629_n N_noxref_21_c_7660_n ) capacitor c=3.74769e-19 \
 //x=63.64 //y=2.08 //x2=63.815 //y2=5.2
cc_4272 ( N_CLK_M130_noxref_g N_noxref_21_c_7660_n ) capacitor c=0.0166421f \
 //x=63.68 //y=6.02 //x2=63.815 //y2=5.2
cc_4273 ( N_CLK_c_6154_n N_noxref_21_c_7660_n ) capacitor c=0.00346519f \
 //x=63.67 //y=4.7 //x2=63.815 //y2=5.2
cc_4274 ( N_CLK_c_5705_n N_noxref_21_c_7664_n ) capacitor c=0.0172877f \
 //x=63.525 //y=4.44 //x2=63.105 //y2=5.2
cc_4275 ( N_CLK_M131_noxref_g N_noxref_21_c_7666_n ) capacitor c=0.0199348f \
 //x=64.12 //y=6.02 //x2=64.295 //y2=5.2
cc_4276 ( N_CLK_c_6197_p N_noxref_21_c_7650_n ) capacitor c=0.00371277f \
 //x=64.05 //y=1.405 //x2=64.295 //y2=1.655
cc_4277 ( N_CLK_c_6151_n N_noxref_21_c_7650_n ) capacitor c=0.00457401f \
 //x=64.205 //y=1.25 //x2=64.295 //y2=1.655
cc_4278 ( N_CLK_c_5705_n N_noxref_21_c_7651_n ) capacitor c=0.00451182f \
 //x=63.525 //y=4.44 //x2=64.38 //y2=3.7
cc_4279 ( N_CLK_c_6133_n N_noxref_21_c_7651_n ) capacitor c=0.00923416f \
 //x=63.64 //y=4.535 //x2=64.38 //y2=3.7
cc_4280 ( N_CLK_c_5629_n N_noxref_21_c_7651_n ) capacitor c=0.0694656f \
 //x=63.64 //y=2.08 //x2=64.38 //y2=3.7
cc_4281 ( N_CLK_c_6163_p N_noxref_21_c_7651_n ) capacitor c=0.0123615f \
 //x=64.045 //y=4.79 //x2=64.38 //y2=3.7
cc_4282 ( N_CLK_c_6152_n N_noxref_21_c_7651_n ) capacitor c=0.00731987f \
 //x=63.64 //y=2.08 //x2=64.38 //y2=3.7
cc_4283 ( N_CLK_c_6241_p N_noxref_21_c_7651_n ) capacitor c=0.00306024f \
 //x=63.64 //y=1.915 //x2=64.38 //y2=3.7
cc_4284 ( N_CLK_c_6154_n N_noxref_21_c_7651_n ) capacitor c=0.00502355f \
 //x=63.67 //y=4.7 //x2=64.38 //y2=3.7
cc_4285 ( N_CLK_c_6163_p N_noxref_21_c_7774_n ) capacitor c=0.00408717f \
 //x=64.045 //y=4.79 //x2=63.9 //y2=5.2
cc_4286 ( N_CLK_M118_noxref_g N_noxref_21_M120_noxref_g ) capacitor \
 c=0.0101598f //x=54.36 //y=6.02 //x2=55.24 //y2=6.02
cc_4287 ( N_CLK_M119_noxref_g N_noxref_21_M120_noxref_g ) capacitor \
 c=0.0602553f //x=54.8 //y=6.02 //x2=55.24 //y2=6.02
cc_4288 ( N_CLK_M119_noxref_g N_noxref_21_M121_noxref_g ) capacitor \
 c=0.0101598f //x=54.8 //y=6.02 //x2=55.68 //y2=6.02
cc_4289 ( N_CLK_c_6119_n N_noxref_21_c_7778_n ) capacitor c=0.00456962f \
 //x=54.48 //y=0.91 //x2=55.49 //y2=0.915
cc_4290 ( N_CLK_c_6120_n N_noxref_21_c_7779_n ) capacitor c=0.00438372f \
 //x=54.48 //y=1.22 //x2=55.49 //y2=1.26
cc_4291 ( N_CLK_c_6121_n N_noxref_21_c_7780_n ) capacitor c=0.00438372f \
 //x=54.48 //y=1.45 //x2=55.49 //y2=1.57
cc_4292 ( N_CLK_c_5628_n N_noxref_21_c_7781_n ) capacitor c=0.00201097f \
 //x=54.39 //y=2.08 //x2=55.5 //y2=2.08
cc_4293 ( N_CLK_c_6122_n N_noxref_21_c_7781_n ) capacitor c=0.00828003f \
 //x=54.48 //y=1.915 //x2=55.5 //y2=2.08
cc_4294 ( N_CLK_c_6122_n N_noxref_21_c_7783_n ) capacitor c=0.00438372f \
 //x=54.48 //y=1.915 //x2=55.5 //y2=1.915
cc_4295 ( N_CLK_c_5705_n N_noxref_21_c_7784_n ) capacitor c=0.0111881f \
 //x=63.525 //y=4.44 //x2=55.5 //y2=4.7
cc_4296 ( N_CLK_c_5628_n N_noxref_21_c_7784_n ) capacitor c=0.00218014f \
 //x=54.39 //y=2.08 //x2=55.5 //y2=4.7
cc_4297 ( N_CLK_c_6179_p N_noxref_21_c_7784_n ) capacitor c=0.0611812f \
 //x=54.725 //y=4.79 //x2=55.5 //y2=4.7
cc_4298 ( N_CLK_c_6124_n N_noxref_21_c_7784_n ) capacitor c=0.00487508f \
 //x=54.39 //y=4.7 //x2=55.5 //y2=4.7
cc_4299 ( N_CLK_c_5705_n N_noxref_21_c_7741_n ) capacitor c=0.0111881f \
 //x=63.525 //y=4.44 //x2=60.31 //y2=4.7
cc_4300 ( N_CLK_c_6142_n N_noxref_21_M39_noxref_d ) capacitor c=0.00217566f \
 //x=63.675 //y=0.905 //x2=63.75 //y2=0.905
cc_4301 ( N_CLK_c_6145_n N_noxref_21_M39_noxref_d ) capacitor c=0.0034598f \
 //x=63.675 //y=1.25 //x2=63.75 //y2=0.905
cc_4302 ( N_CLK_c_6147_n N_noxref_21_M39_noxref_d ) capacitor c=0.00669531f \
 //x=63.675 //y=1.56 //x2=63.75 //y2=0.905
cc_4303 ( N_CLK_c_6261_p N_noxref_21_M39_noxref_d ) capacitor c=0.00241102f \
 //x=64.05 //y=0.75 //x2=63.75 //y2=0.905
cc_4304 ( N_CLK_c_6197_p N_noxref_21_M39_noxref_d ) capacitor c=0.0137169f \
 //x=64.05 //y=1.405 //x2=63.75 //y2=0.905
cc_4305 ( N_CLK_c_6150_n N_noxref_21_M39_noxref_d ) capacitor c=0.00132245f \
 //x=64.205 //y=0.905 //x2=63.75 //y2=0.905
cc_4306 ( N_CLK_c_6151_n N_noxref_21_M39_noxref_d ) capacitor c=0.00566463f \
 //x=64.205 //y=1.25 //x2=63.75 //y2=0.905
cc_4307 ( N_CLK_c_6241_p N_noxref_21_M39_noxref_d ) capacitor c=0.00660593f \
 //x=63.64 //y=1.915 //x2=63.75 //y2=0.905
cc_4308 ( N_CLK_M130_noxref_g N_noxref_21_M130_noxref_d ) capacitor \
 c=0.0173476f //x=63.68 //y=6.02 //x2=63.755 //y2=5.02
cc_4309 ( N_CLK_M131_noxref_g N_noxref_21_M130_noxref_d ) capacitor \
 c=0.0179769f //x=64.12 //y=6.02 //x2=63.755 //y2=5.02
cc_4310 ( N_CLK_c_5705_n N_noxref_23_c_8092_n ) capacitor c=0.00472509f \
 //x=63.525 //y=4.44 //x2=67.085 //y2=4.44
cc_4311 ( N_CLK_c_5643_n N_noxref_24_c_8520_n ) capacitor c=0.0309065f \
 //x=29.855 //y=4.44 //x2=23.565 //y2=3.33
cc_4312 ( N_CLK_c_5643_n N_noxref_24_c_8497_n ) capacitor c=6.53919e-19 \
 //x=29.855 //y=4.44 //x2=18.245 //y2=3.33
cc_4313 ( N_CLK_c_5643_n N_noxref_24_c_8424_n ) capacitor c=0.08511f \
 //x=29.855 //y=4.44 //x2=79.065 //y2=3.33
cc_4314 ( N_CLK_c_5668_n N_noxref_24_c_8424_n ) capacitor c=0.00667512f \
 //x=39.105 //y=4.44 //x2=79.065 //y2=3.33
cc_4315 ( N_CLK_c_5679_n N_noxref_24_c_8424_n ) capacitor c=5.01525e-19 \
 //x=30.085 //y=4.44 //x2=79.065 //y2=3.33
cc_4316 ( N_CLK_c_5680_n N_noxref_24_c_8424_n ) capacitor c=0.0917934f \
 //x=54.275 //y=4.44 //x2=79.065 //y2=3.33
cc_4317 ( N_CLK_c_5705_n N_noxref_24_c_8424_n ) capacitor c=0.00667512f \
 //x=63.525 //y=4.44 //x2=79.065 //y2=3.33
cc_4318 ( N_CLK_c_5716_n N_noxref_24_c_8424_n ) capacitor c=5.01525e-19 \
 //x=54.505 //y=4.44 //x2=79.065 //y2=3.33
cc_4319 ( N_CLK_c_5625_n N_noxref_24_c_8424_n ) capacitor c=0.0213922f \
 //x=29.97 //y=2.08 //x2=79.065 //y2=3.33
cc_4320 ( N_CLK_c_5626_n N_noxref_24_c_8424_n ) capacitor c=0.0169786f \
 //x=39.22 //y=2.08 //x2=79.065 //y2=3.33
cc_4321 ( N_CLK_c_5628_n N_noxref_24_c_8424_n ) capacitor c=0.0213922f \
 //x=54.39 //y=2.08 //x2=79.065 //y2=3.33
cc_4322 ( N_CLK_c_5629_n N_noxref_24_c_8424_n ) capacitor c=0.0169786f \
 //x=63.64 //y=2.08 //x2=79.065 //y2=3.33
cc_4323 ( N_CLK_c_5643_n N_noxref_24_c_8558_n ) capacitor c=0.00698923f \
 //x=29.855 //y=4.44 //x2=23.795 //y2=3.33
cc_4324 ( N_CLK_c_5643_n N_noxref_24_c_8498_n ) capacitor c=0.0016972f \
 //x=29.855 //y=4.44 //x2=18.13 //y2=4.535
cc_4325 ( N_CLK_c_5643_n N_noxref_24_c_8428_n ) capacitor c=0.0212595f \
 //x=29.855 //y=4.44 //x2=18.13 //y2=2.08
cc_4326 ( N_CLK_c_5643_n N_noxref_24_c_8451_n ) capacitor c=0.032141f \
 //x=29.855 //y=4.44 //x2=21.935 //y2=5.155
cc_4327 ( N_CLK_c_5643_n N_noxref_24_c_8455_n ) capacitor c=0.0230136f \
 //x=29.855 //y=4.44 //x2=21.225 //y2=5.155
cc_4328 ( N_CLK_c_5643_n N_noxref_24_c_8461_n ) capacitor c=0.0183122f \
 //x=29.855 //y=4.44 //x2=23.595 //y2=5.155
cc_4329 ( N_CLK_c_5643_n N_noxref_24_c_8465_n ) capacitor c=0.0249802f \
 //x=29.855 //y=4.44 //x2=23.68 //y2=3.33
cc_4330 ( N_CLK_c_5643_n N_noxref_24_c_8541_n ) capacitor c=0.00960248f \
 //x=29.855 //y=4.44 //x2=18.535 //y2=4.79
cc_4331 ( N_CLK_c_5643_n N_noxref_24_c_8518_n ) capacitor c=0.00203982f \
 //x=29.855 //y=4.44 //x2=18.16 //y2=4.7
cc_4332 ( N_CLK_c_5769_n N_noxref_28_c_9285_n ) capacitor c=0.0167228f \
 //x=5.115 //y=0.91 //x2=5.775 //y2=0.54
cc_4333 ( N_CLK_c_5774_n N_noxref_28_c_9285_n ) capacitor c=0.00534519f \
 //x=5.64 //y=0.91 //x2=5.775 //y2=0.54
cc_4334 ( N_CLK_c_5622_n N_noxref_28_c_9304_n ) capacitor c=0.012334f //x=5.55 \
 //y=2.08 //x2=5.775 //y2=1.59
cc_4335 ( N_CLK_c_5772_n N_noxref_28_c_9304_n ) capacitor c=0.0153476f \
 //x=5.115 //y=1.22 //x2=5.775 //y2=1.59
cc_4336 ( N_CLK_c_5777_n N_noxref_28_c_9304_n ) capacitor c=0.0219329f \
 //x=5.64 //y=1.915 //x2=5.775 //y2=1.59
cc_4337 ( N_CLK_c_5769_n N_noxref_28_M2_noxref_s ) capacitor c=0.00798959f \
 //x=5.115 //y=0.91 //x2=3.785 //y2=0.375
cc_4338 ( N_CLK_c_5776_n N_noxref_28_M2_noxref_s ) capacitor c=0.00212176f \
 //x=5.64 //y=1.45 //x2=3.785 //y2=0.375
cc_4339 ( N_CLK_c_5777_n N_noxref_28_M2_noxref_s ) capacitor c=0.00298115f \
 //x=5.64 //y=1.915 //x2=3.785 //y2=0.375
cc_4340 ( N_CLK_c_6298_p N_noxref_29_c_9329_n ) capacitor c=2.14837e-19 \
 //x=5.485 //y=0.755 //x2=6.345 //y2=0.995
cc_4341 ( N_CLK_c_5774_n N_noxref_29_c_9329_n ) capacitor c=0.00123426f \
 //x=5.64 //y=0.91 //x2=6.345 //y2=0.995
cc_4342 ( N_CLK_c_5775_n N_noxref_29_c_9329_n ) capacitor c=0.0129288f \
 //x=5.64 //y=1.22 //x2=6.345 //y2=0.995
cc_4343 ( N_CLK_c_5776_n N_noxref_29_c_9329_n ) capacitor c=0.00142359f \
 //x=5.64 //y=1.45 //x2=6.345 //y2=0.995
cc_4344 ( N_CLK_c_5769_n N_noxref_29_M3_noxref_d ) capacitor c=0.00223875f \
 //x=5.115 //y=0.91 //x2=5.19 //y2=0.91
cc_4345 ( N_CLK_c_5772_n N_noxref_29_M3_noxref_d ) capacitor c=0.00262485f \
 //x=5.115 //y=1.22 //x2=5.19 //y2=0.91
cc_4346 ( N_CLK_c_6298_p N_noxref_29_M3_noxref_d ) capacitor c=0.00220746f \
 //x=5.485 //y=0.755 //x2=5.19 //y2=0.91
cc_4347 ( N_CLK_c_6305_p N_noxref_29_M3_noxref_d ) capacitor c=0.00194798f \
 //x=5.485 //y=1.375 //x2=5.19 //y2=0.91
cc_4348 ( N_CLK_c_5774_n N_noxref_29_M3_noxref_d ) capacitor c=0.00198465f \
 //x=5.64 //y=0.91 //x2=5.19 //y2=0.91
cc_4349 ( N_CLK_c_5775_n N_noxref_29_M3_noxref_d ) capacitor c=0.00128384f \
 //x=5.64 //y=1.22 //x2=5.19 //y2=0.91
cc_4350 ( N_CLK_c_5774_n N_noxref_29_M4_noxref_s ) capacitor c=7.21316e-19 \
 //x=5.64 //y=0.91 //x2=6.295 //y2=0.375
cc_4351 ( N_CLK_c_5775_n N_noxref_29_M4_noxref_s ) capacitor c=0.00348171f \
 //x=5.64 //y=1.22 //x2=6.295 //y2=0.375
cc_4352 ( N_CLK_c_5805_n N_noxref_32_c_9493_n ) capacitor c=0.00623646f \
 //x=14.835 //y=1.56 //x2=14.615 //y2=1.495
cc_4353 ( N_CLK_c_5810_n N_noxref_32_c_9493_n ) capacitor c=0.00173579f \
 //x=14.8 //y=2.08 //x2=14.615 //y2=1.495
cc_4354 ( N_CLK_c_5623_n N_noxref_32_c_9494_n ) capacitor c=0.00156605f \
 //x=14.8 //y=2.08 //x2=15.5 //y2=0.53
cc_4355 ( N_CLK_c_5800_n N_noxref_32_c_9494_n ) capacitor c=0.0188655f \
 //x=14.835 //y=0.905 //x2=15.5 //y2=0.53
cc_4356 ( N_CLK_c_5808_n N_noxref_32_c_9494_n ) capacitor c=0.00656458f \
 //x=15.365 //y=0.905 //x2=15.5 //y2=0.53
cc_4357 ( N_CLK_c_5810_n N_noxref_32_c_9494_n ) capacitor c=2.1838e-19 \
 //x=14.8 //y=2.08 //x2=15.5 //y2=0.53
cc_4358 ( N_CLK_c_5800_n N_noxref_32_M8_noxref_s ) capacitor c=0.00623646f \
 //x=14.835 //y=0.905 //x2=13.51 //y2=0.365
cc_4359 ( N_CLK_c_5808_n N_noxref_32_M8_noxref_s ) capacitor c=0.0143002f \
 //x=15.365 //y=0.905 //x2=13.51 //y2=0.365
cc_4360 ( N_CLK_c_5809_n N_noxref_32_M8_noxref_s ) capacitor c=0.00290153f \
 //x=15.365 //y=1.25 //x2=13.51 //y2=0.365
cc_4361 ( N_CLK_c_5926_n N_noxref_37_c_9750_n ) capacitor c=0.0167228f \
 //x=29.535 //y=0.91 //x2=30.195 //y2=0.54
cc_4362 ( N_CLK_c_5931_n N_noxref_37_c_9750_n ) capacitor c=0.00534519f \
 //x=30.06 //y=0.91 //x2=30.195 //y2=0.54
cc_4363 ( N_CLK_c_5625_n N_noxref_37_c_9773_n ) capacitor c=0.0117694f \
 //x=29.97 //y=2.08 //x2=30.195 //y2=1.59
cc_4364 ( N_CLK_c_5929_n N_noxref_37_c_9773_n ) capacitor c=0.0157358f \
 //x=29.535 //y=1.22 //x2=30.195 //y2=1.59
cc_4365 ( N_CLK_c_5934_n N_noxref_37_c_9773_n ) capacitor c=0.021347f \
 //x=30.06 //y=1.915 //x2=30.195 //y2=1.59
cc_4366 ( N_CLK_c_5926_n N_noxref_37_M17_noxref_s ) capacitor c=0.00798959f \
 //x=29.535 //y=0.91 //x2=28.205 //y2=0.375
cc_4367 ( N_CLK_c_5933_n N_noxref_37_M17_noxref_s ) capacitor c=0.00212176f \
 //x=30.06 //y=1.45 //x2=28.205 //y2=0.375
cc_4368 ( N_CLK_c_5934_n N_noxref_37_M17_noxref_s ) capacitor c=0.00298115f \
 //x=30.06 //y=1.915 //x2=28.205 //y2=0.375
cc_4369 ( N_CLK_c_6327_p N_noxref_38_c_9792_n ) capacitor c=2.14837e-19 \
 //x=29.905 //y=0.755 //x2=30.765 //y2=0.995
cc_4370 ( N_CLK_c_5931_n N_noxref_38_c_9792_n ) capacitor c=0.00123426f \
 //x=30.06 //y=0.91 //x2=30.765 //y2=0.995
cc_4371 ( N_CLK_c_5932_n N_noxref_38_c_9792_n ) capacitor c=0.0129288f \
 //x=30.06 //y=1.22 //x2=30.765 //y2=0.995
cc_4372 ( N_CLK_c_5933_n N_noxref_38_c_9792_n ) capacitor c=0.00142359f \
 //x=30.06 //y=1.45 //x2=30.765 //y2=0.995
cc_4373 ( N_CLK_c_5926_n N_noxref_38_M18_noxref_d ) capacitor c=0.00223875f \
 //x=29.535 //y=0.91 //x2=29.61 //y2=0.91
cc_4374 ( N_CLK_c_5929_n N_noxref_38_M18_noxref_d ) capacitor c=0.00262485f \
 //x=29.535 //y=1.22 //x2=29.61 //y2=0.91
cc_4375 ( N_CLK_c_6327_p N_noxref_38_M18_noxref_d ) capacitor c=0.00220746f \
 //x=29.905 //y=0.755 //x2=29.61 //y2=0.91
cc_4376 ( N_CLK_c_6334_p N_noxref_38_M18_noxref_d ) capacitor c=0.00194798f \
 //x=29.905 //y=1.375 //x2=29.61 //y2=0.91
cc_4377 ( N_CLK_c_5931_n N_noxref_38_M18_noxref_d ) capacitor c=0.00198465f \
 //x=30.06 //y=0.91 //x2=29.61 //y2=0.91
cc_4378 ( N_CLK_c_5932_n N_noxref_38_M18_noxref_d ) capacitor c=0.00128384f \
 //x=30.06 //y=1.22 //x2=29.61 //y2=0.91
cc_4379 ( N_CLK_c_5931_n N_noxref_38_M19_noxref_s ) capacitor c=7.21316e-19 \
 //x=30.06 //y=0.91 //x2=30.715 //y2=0.375
cc_4380 ( N_CLK_c_5932_n N_noxref_38_M19_noxref_s ) capacitor c=0.00348171f \
 //x=30.06 //y=1.22 //x2=30.715 //y2=0.375
cc_4381 ( N_CLK_c_5961_n N_noxref_41_c_9955_n ) capacitor c=0.00623646f \
 //x=39.255 //y=1.56 //x2=39.035 //y2=1.495
cc_4382 ( N_CLK_c_5966_n N_noxref_41_c_9955_n ) capacitor c=0.00173579f \
 //x=39.22 //y=2.08 //x2=39.035 //y2=1.495
cc_4383 ( N_CLK_c_5626_n N_noxref_41_c_9956_n ) capacitor c=0.00156605f \
 //x=39.22 //y=2.08 //x2=39.92 //y2=0.53
cc_4384 ( N_CLK_c_5956_n N_noxref_41_c_9956_n ) capacitor c=0.0188655f \
 //x=39.255 //y=0.905 //x2=39.92 //y2=0.53
cc_4385 ( N_CLK_c_5964_n N_noxref_41_c_9956_n ) capacitor c=0.00656458f \
 //x=39.785 //y=0.905 //x2=39.92 //y2=0.53
cc_4386 ( N_CLK_c_5966_n N_noxref_41_c_9956_n ) capacitor c=2.1838e-19 \
 //x=39.22 //y=2.08 //x2=39.92 //y2=0.53
cc_4387 ( N_CLK_c_5956_n N_noxref_41_M23_noxref_s ) capacitor c=0.00623646f \
 //x=39.255 //y=0.905 //x2=37.93 //y2=0.365
cc_4388 ( N_CLK_c_5964_n N_noxref_41_M23_noxref_s ) capacitor c=0.0143002f \
 //x=39.785 //y=0.905 //x2=37.93 //y2=0.365
cc_4389 ( N_CLK_c_5965_n N_noxref_41_M23_noxref_s ) capacitor c=0.00290153f \
 //x=39.785 //y=1.25 //x2=37.93 //y2=0.365
cc_4390 ( N_CLK_c_6114_n N_noxref_46_c_10212_n ) capacitor c=0.0167228f \
 //x=53.955 //y=0.91 //x2=54.615 //y2=0.54
cc_4391 ( N_CLK_c_6119_n N_noxref_46_c_10212_n ) capacitor c=0.00534519f \
 //x=54.48 //y=0.91 //x2=54.615 //y2=0.54
cc_4392 ( N_CLK_c_5628_n N_noxref_46_c_10234_n ) capacitor c=0.0117694f \
 //x=54.39 //y=2.08 //x2=54.615 //y2=1.59
cc_4393 ( N_CLK_c_6117_n N_noxref_46_c_10234_n ) capacitor c=0.0157358f \
 //x=53.955 //y=1.22 //x2=54.615 //y2=1.59
cc_4394 ( N_CLK_c_6122_n N_noxref_46_c_10234_n ) capacitor c=0.021347f \
 //x=54.48 //y=1.915 //x2=54.615 //y2=1.59
cc_4395 ( N_CLK_c_6114_n N_noxref_46_M32_noxref_s ) capacitor c=0.00798959f \
 //x=53.955 //y=0.91 //x2=52.625 //y2=0.375
cc_4396 ( N_CLK_c_6121_n N_noxref_46_M32_noxref_s ) capacitor c=0.00212176f \
 //x=54.48 //y=1.45 //x2=52.625 //y2=0.375
cc_4397 ( N_CLK_c_6122_n N_noxref_46_M32_noxref_s ) capacitor c=0.00298115f \
 //x=54.48 //y=1.915 //x2=52.625 //y2=0.375
cc_4398 ( N_CLK_c_6356_p N_noxref_47_c_10254_n ) capacitor c=2.14837e-19 \
 //x=54.325 //y=0.755 //x2=55.185 //y2=0.995
cc_4399 ( N_CLK_c_6119_n N_noxref_47_c_10254_n ) capacitor c=0.00123426f \
 //x=54.48 //y=0.91 //x2=55.185 //y2=0.995
cc_4400 ( N_CLK_c_6120_n N_noxref_47_c_10254_n ) capacitor c=0.0129288f \
 //x=54.48 //y=1.22 //x2=55.185 //y2=0.995
cc_4401 ( N_CLK_c_6121_n N_noxref_47_c_10254_n ) capacitor c=0.00142359f \
 //x=54.48 //y=1.45 //x2=55.185 //y2=0.995
cc_4402 ( N_CLK_c_6114_n N_noxref_47_M33_noxref_d ) capacitor c=0.00223875f \
 //x=53.955 //y=0.91 //x2=54.03 //y2=0.91
cc_4403 ( N_CLK_c_6117_n N_noxref_47_M33_noxref_d ) capacitor c=0.00262485f \
 //x=53.955 //y=1.22 //x2=54.03 //y2=0.91
cc_4404 ( N_CLK_c_6356_p N_noxref_47_M33_noxref_d ) capacitor c=0.00220746f \
 //x=54.325 //y=0.755 //x2=54.03 //y2=0.91
cc_4405 ( N_CLK_c_6363_p N_noxref_47_M33_noxref_d ) capacitor c=0.00194798f \
 //x=54.325 //y=1.375 //x2=54.03 //y2=0.91
cc_4406 ( N_CLK_c_6119_n N_noxref_47_M33_noxref_d ) capacitor c=0.00198465f \
 //x=54.48 //y=0.91 //x2=54.03 //y2=0.91
cc_4407 ( N_CLK_c_6120_n N_noxref_47_M33_noxref_d ) capacitor c=0.00128384f \
 //x=54.48 //y=1.22 //x2=54.03 //y2=0.91
cc_4408 ( N_CLK_c_6119_n N_noxref_47_M34_noxref_s ) capacitor c=7.21316e-19 \
 //x=54.48 //y=0.91 //x2=55.135 //y2=0.375
cc_4409 ( N_CLK_c_6120_n N_noxref_47_M34_noxref_s ) capacitor c=0.00348171f \
 //x=54.48 //y=1.22 //x2=55.135 //y2=0.375
cc_4410 ( N_CLK_c_6147_n N_noxref_50_c_10417_n ) capacitor c=0.00623646f \
 //x=63.675 //y=1.56 //x2=63.455 //y2=1.495
cc_4411 ( N_CLK_c_6152_n N_noxref_50_c_10417_n ) capacitor c=0.00173579f \
 //x=63.64 //y=2.08 //x2=63.455 //y2=1.495
cc_4412 ( N_CLK_c_5629_n N_noxref_50_c_10418_n ) capacitor c=0.00156605f \
 //x=63.64 //y=2.08 //x2=64.34 //y2=0.53
cc_4413 ( N_CLK_c_6142_n N_noxref_50_c_10418_n ) capacitor c=0.0188655f \
 //x=63.675 //y=0.905 //x2=64.34 //y2=0.53
cc_4414 ( N_CLK_c_6150_n N_noxref_50_c_10418_n ) capacitor c=0.00656458f \
 //x=64.205 //y=0.905 //x2=64.34 //y2=0.53
cc_4415 ( N_CLK_c_6152_n N_noxref_50_c_10418_n ) capacitor c=2.1838e-19 \
 //x=63.64 //y=2.08 //x2=64.34 //y2=0.53
cc_4416 ( N_CLK_c_6142_n N_noxref_50_M38_noxref_s ) capacitor c=0.00623646f \
 //x=63.675 //y=0.905 //x2=62.35 //y2=0.365
cc_4417 ( N_CLK_c_6150_n N_noxref_50_M38_noxref_s ) capacitor c=0.0143002f \
 //x=64.205 //y=0.905 //x2=62.35 //y2=0.365
cc_4418 ( N_CLK_c_6151_n N_noxref_50_M38_noxref_s ) capacitor c=0.00290153f \
 //x=64.205 //y=1.25 //x2=62.35 //y2=0.365
cc_4419 ( N_noxref_18_M133_noxref_g N_noxref_19_c_6694_n ) capacitor \
 c=0.0187084f //x=66.57 //y=6.02 //x2=67.145 //y2=5.2
cc_4420 ( N_noxref_18_c_6393_n N_noxref_19_c_6698_n ) capacitor c=0.00144307f \
 //x=66.115 //y=4.07 //x2=66.435 //y2=5.2
cc_4421 ( N_noxref_18_c_6380_n N_noxref_19_c_6698_n ) capacitor c=0.00529872f \
 //x=66.23 //y=2.08 //x2=66.435 //y2=5.2
cc_4422 ( N_noxref_18_M132_noxref_g N_noxref_19_c_6698_n ) capacitor \
 c=0.0177326f //x=66.13 //y=6.02 //x2=66.435 //y2=5.2
cc_4423 ( N_noxref_18_c_6432_n N_noxref_19_c_6698_n ) capacitor c=0.00585724f \
 //x=66.23 //y=4.7 //x2=66.435 //y2=5.2
cc_4424 ( N_noxref_18_c_6380_n N_noxref_19_c_6669_n ) capacitor c=0.00309648f \
 //x=66.23 //y=2.08 //x2=67.71 //y2=4.81
cc_4425 ( N_noxref_18_M133_noxref_g N_noxref_19_M132_noxref_d ) capacitor \
 c=0.0173476f //x=66.57 //y=6.02 //x2=66.205 //y2=5.02
cc_4426 ( N_noxref_18_c_6377_n N_SN_c_6866_n ) capacitor c=0.0178519f \
 //x=50.69 //y=2.08 //x2=59.085 //y2=2.22
cc_4427 ( N_noxref_18_c_6558_p N_SN_c_6866_n ) capacitor c=0.0163057f \
 //x=55.84 //y=1.665 //x2=59.085 //y2=2.22
cc_4428 ( N_noxref_18_c_6456_n N_SN_c_6866_n ) capacitor c=0.0197307f \
 //x=56.237 //y=3.905 //x2=59.085 //y2=2.22
cc_4429 ( N_noxref_18_c_6506_n N_SN_c_6866_n ) capacitor c=3.11115e-19 \
 //x=51.1 //y=1.405 //x2=59.085 //y2=2.22
cc_4430 ( N_noxref_18_c_6476_n N_SN_c_6866_n ) capacitor c=0.00570799f \
 //x=50.69 //y=2.08 //x2=59.085 //y2=2.22
cc_4431 ( N_noxref_18_c_6380_n N_SN_c_6877_n ) capacitor c=0.0208418f \
 //x=66.23 //y=2.08 //x2=70.555 //y2=2.22
cc_4432 ( N_noxref_18_c_6385_n N_SN_c_6877_n ) capacitor c=0.00894156f \
 //x=66.035 //y=1.915 //x2=70.555 //y2=2.22
cc_4433 ( N_noxref_18_c_6393_n N_SN_c_6892_n ) capacitor c=0.0190126f \
 //x=66.115 //y=4.07 //x2=59.2 //y2=2.08
cc_4434 ( N_noxref_18_c_6456_n N_SN_c_6892_n ) capacitor c=3.18993e-19 \
 //x=56.237 //y=3.905 //x2=59.2 //y2=2.08
cc_4435 ( N_noxref_18_c_6392_n N_noxref_21_c_7696_n ) capacitor c=0.044143f \
 //x=56.12 //y=4.07 //x2=60.195 //y2=3.7
cc_4436 ( N_noxref_18_c_6393_n N_noxref_21_c_7696_n ) capacitor c=0.340271f \
 //x=66.115 //y=4.07 //x2=60.195 //y2=3.7
cc_4437 ( N_noxref_18_c_6402_n N_noxref_21_c_7696_n ) capacitor c=0.0267581f \
 //x=56.35 //y=4.07 //x2=60.195 //y2=3.7
cc_4438 ( N_noxref_18_c_6422_n N_noxref_21_c_7696_n ) capacitor c=0.00219785f \
 //x=56.235 //y=4.07 //x2=60.195 //y2=3.7
cc_4439 ( N_noxref_18_c_6456_n N_noxref_21_c_7696_n ) capacitor c=0.0185057f \
 //x=56.237 //y=3.905 //x2=60.195 //y2=3.7
cc_4440 ( N_noxref_18_c_6392_n N_noxref_21_c_7697_n ) capacitor c=0.0292842f \
 //x=56.12 //y=4.07 //x2=55.615 //y2=3.7
cc_4441 ( N_noxref_18_c_6456_n N_noxref_21_c_7697_n ) capacitor c=0.00179385f \
 //x=56.237 //y=3.905 //x2=55.615 //y2=3.7
cc_4442 ( N_noxref_18_c_6393_n N_noxref_21_c_7698_n ) capacitor c=0.339174f \
 //x=66.115 //y=4.07 //x2=64.265 //y2=3.7
cc_4443 ( N_noxref_18_c_6393_n N_noxref_21_c_7699_n ) capacitor c=0.026596f \
 //x=66.115 //y=4.07 //x2=60.425 //y2=3.7
cc_4444 ( N_noxref_18_c_6393_n N_noxref_21_c_7656_n ) capacitor c=0.17615f \
 //x=66.115 //y=4.07 //x2=71.665 //y2=3.7
cc_4445 ( N_noxref_18_c_6380_n N_noxref_21_c_7656_n ) capacitor c=0.0205593f \
 //x=66.23 //y=2.08 //x2=71.665 //y2=3.7
cc_4446 ( N_noxref_18_c_6432_n N_noxref_21_c_7656_n ) capacitor c=0.00463981f \
 //x=66.23 //y=4.7 //x2=71.665 //y2=3.7
cc_4447 ( N_noxref_18_c_6393_n N_noxref_21_c_7701_n ) capacitor c=0.026743f \
 //x=66.115 //y=4.07 //x2=64.495 //y2=3.7
cc_4448 ( N_noxref_18_c_6380_n N_noxref_21_c_7701_n ) capacitor c=7.01366e-19 \
 //x=66.23 //y=2.08 //x2=64.495 //y2=3.7
cc_4449 ( N_noxref_18_c_6392_n N_noxref_21_c_7648_n ) capacitor c=0.0197867f \
 //x=56.12 //y=4.07 //x2=55.5 //y2=2.08
cc_4450 ( N_noxref_18_c_6402_n N_noxref_21_c_7648_n ) capacitor c=0.00180189f \
 //x=56.35 //y=4.07 //x2=55.5 //y2=2.08
cc_4451 ( N_noxref_18_c_6539_n N_noxref_21_c_7648_n ) capacitor c=0.0163236f \
 //x=56.24 //y=5.07 //x2=55.5 //y2=2.08
cc_4452 ( N_noxref_18_c_6583_p N_noxref_21_c_7648_n ) capacitor c=0.016476f \
 //x=55.46 //y=5.155 //x2=55.5 //y2=2.08
cc_4453 ( N_noxref_18_c_6422_n N_noxref_21_c_7648_n ) capacitor c=0.00966503f \
 //x=56.235 //y=4.07 //x2=55.5 //y2=2.08
cc_4454 ( N_noxref_18_c_6456_n N_noxref_21_c_7648_n ) capacitor c=0.0508802f \
 //x=56.237 //y=3.905 //x2=55.5 //y2=2.08
cc_4455 ( N_noxref_18_c_6393_n N_noxref_21_c_7649_n ) capacitor c=0.0198068f \
 //x=66.115 //y=4.07 //x2=60.31 //y2=2.08
cc_4456 ( N_noxref_18_c_6393_n N_noxref_21_c_7660_n ) capacitor c=0.0126022f \
 //x=66.115 //y=4.07 //x2=63.815 //y2=5.2
cc_4457 ( N_noxref_18_c_6393_n N_noxref_21_c_7651_n ) capacitor c=0.0253623f \
 //x=66.115 //y=4.07 //x2=64.38 //y2=3.7
cc_4458 ( N_noxref_18_c_6380_n N_noxref_21_c_7651_n ) capacitor c=0.011807f \
 //x=66.23 //y=2.08 //x2=64.38 //y2=3.7
cc_4459 ( N_noxref_18_c_6411_n N_noxref_21_M120_noxref_g ) capacitor \
 c=0.01736f //x=55.375 //y=5.155 //x2=55.24 //y2=6.02
cc_4460 ( N_noxref_18_M120_noxref_d N_noxref_21_M120_noxref_g ) capacitor \
 c=0.0180032f //x=55.315 //y=5.02 //x2=55.24 //y2=6.02
cc_4461 ( N_noxref_18_c_6415_n N_noxref_21_M121_noxref_g ) capacitor \
 c=0.0194981f //x=56.155 //y=5.155 //x2=55.68 //y2=6.02
cc_4462 ( N_noxref_18_M120_noxref_d N_noxref_21_M121_noxref_g ) capacitor \
 c=0.0194246f //x=55.315 //y=5.02 //x2=55.68 //y2=6.02
cc_4463 ( N_noxref_18_M34_noxref_d N_noxref_21_c_7778_n ) capacitor \
 c=0.00217566f //x=55.565 //y=0.915 //x2=55.49 //y2=0.915
cc_4464 ( N_noxref_18_M34_noxref_d N_noxref_21_c_7779_n ) capacitor \
 c=0.0034598f //x=55.565 //y=0.915 //x2=55.49 //y2=1.26
cc_4465 ( N_noxref_18_M34_noxref_d N_noxref_21_c_7780_n ) capacitor \
 c=0.00546784f //x=55.565 //y=0.915 //x2=55.49 //y2=1.57
cc_4466 ( N_noxref_18_M34_noxref_d N_noxref_21_c_7830_n ) capacitor \
 c=0.00241102f //x=55.565 //y=0.915 //x2=55.865 //y2=0.76
cc_4467 ( N_noxref_18_c_6379_n N_noxref_21_c_7831_n ) capacitor c=0.00371277f \
 //x=56.155 //y=1.665 //x2=55.865 //y2=1.415
cc_4468 ( N_noxref_18_M34_noxref_d N_noxref_21_c_7831_n ) capacitor \
 c=0.0138621f //x=55.565 //y=0.915 //x2=55.865 //y2=1.415
cc_4469 ( N_noxref_18_M34_noxref_d N_noxref_21_c_7833_n ) capacitor \
 c=0.00219619f //x=55.565 //y=0.915 //x2=56.02 //y2=0.915
cc_4470 ( N_noxref_18_c_6379_n N_noxref_21_c_7834_n ) capacitor c=0.00457401f \
 //x=56.155 //y=1.665 //x2=56.02 //y2=1.26
cc_4471 ( N_noxref_18_M34_noxref_d N_noxref_21_c_7834_n ) capacitor \
 c=0.00603828f //x=55.565 //y=0.915 //x2=56.02 //y2=1.26
cc_4472 ( N_noxref_18_c_6456_n N_noxref_21_c_7781_n ) capacitor c=0.00709342f \
 //x=56.237 //y=3.905 //x2=55.5 //y2=2.08
cc_4473 ( N_noxref_18_c_6456_n N_noxref_21_c_7783_n ) capacitor c=0.00404774f \
 //x=56.237 //y=3.905 //x2=55.5 //y2=1.915
cc_4474 ( N_noxref_18_M34_noxref_d N_noxref_21_c_7783_n ) capacitor \
 c=0.00661782f //x=55.565 //y=0.915 //x2=55.5 //y2=1.915
cc_4475 ( N_noxref_18_c_6415_n N_noxref_21_c_7784_n ) capacitor c=0.00201851f \
 //x=56.155 //y=5.155 //x2=55.5 //y2=4.7
cc_4476 ( N_noxref_18_c_6539_n N_noxref_21_c_7784_n ) capacitor c=0.0151148f \
 //x=56.24 //y=5.07 //x2=55.5 //y2=4.7
cc_4477 ( N_noxref_18_c_6583_p N_noxref_21_c_7784_n ) capacitor c=0.00475601f \
 //x=55.46 //y=5.155 //x2=55.5 //y2=4.7
cc_4478 ( N_noxref_18_c_6380_n N_noxref_23_c_8092_n ) capacitor c=0.00470962f \
 //x=66.23 //y=2.08 //x2=67.085 //y2=4.44
cc_4479 ( N_noxref_18_c_6432_n N_noxref_23_c_8092_n ) capacitor c=2.48643e-19 \
 //x=66.23 //y=4.7 //x2=67.085 //y2=4.44
cc_4480 ( N_noxref_18_c_6380_n N_noxref_23_c_8213_n ) capacitor c=0.00371837f \
 //x=66.23 //y=2.08 //x2=66.97 //y2=4.535
cc_4481 ( N_noxref_18_c_6432_n N_noxref_23_c_8213_n ) capacitor c=0.00415951f \
 //x=66.23 //y=4.7 //x2=66.97 //y2=4.535
cc_4482 ( N_noxref_18_c_6393_n N_noxref_23_c_8060_n ) capacitor c=0.00735597f \
 //x=66.115 //y=4.07 //x2=66.97 //y2=2.08
cc_4483 ( N_noxref_18_c_6380_n N_noxref_23_c_8060_n ) capacitor c=0.0754429f \
 //x=66.23 //y=2.08 //x2=66.97 //y2=2.08
cc_4484 ( N_noxref_18_c_6385_n N_noxref_23_c_8060_n ) capacitor c=0.00284029f \
 //x=66.035 //y=1.915 //x2=66.97 //y2=2.08
cc_4485 ( N_noxref_18_M132_noxref_g N_noxref_23_M134_noxref_g ) capacitor \
 c=0.0104611f //x=66.13 //y=6.02 //x2=67.01 //y2=6.02
cc_4486 ( N_noxref_18_M133_noxref_g N_noxref_23_M134_noxref_g ) capacitor \
 c=0.106618f //x=66.57 //y=6.02 //x2=67.01 //y2=6.02
cc_4487 ( N_noxref_18_M133_noxref_g N_noxref_23_M135_noxref_g ) capacitor \
 c=0.0101362f //x=66.57 //y=6.02 //x2=67.45 //y2=6.02
cc_4488 ( N_noxref_18_c_6381_n N_noxref_23_c_8221_n ) capacitor c=4.86506e-19 \
 //x=66.035 //y=0.865 //x2=67.005 //y2=0.905
cc_4489 ( N_noxref_18_c_6383_n N_noxref_23_c_8221_n ) capacitor c=0.00152104f \
 //x=66.035 //y=1.21 //x2=67.005 //y2=0.905
cc_4490 ( N_noxref_18_c_6388_n N_noxref_23_c_8221_n ) capacitor c=0.0151475f \
 //x=66.565 //y=0.865 //x2=67.005 //y2=0.905
cc_4491 ( N_noxref_18_c_6384_n N_noxref_23_c_8224_n ) capacitor c=0.00109982f \
 //x=66.035 //y=1.52 //x2=67.005 //y2=1.25
cc_4492 ( N_noxref_18_c_6390_n N_noxref_23_c_8224_n ) capacitor c=0.0111064f \
 //x=66.565 //y=1.21 //x2=67.005 //y2=1.25
cc_4493 ( N_noxref_18_c_6384_n N_noxref_23_c_8226_n ) capacitor c=9.57794e-19 \
 //x=66.035 //y=1.52 //x2=67.005 //y2=1.56
cc_4494 ( N_noxref_18_c_6385_n N_noxref_23_c_8226_n ) capacitor c=0.00662747f \
 //x=66.035 //y=1.915 //x2=67.005 //y2=1.56
cc_4495 ( N_noxref_18_c_6390_n N_noxref_23_c_8226_n ) capacitor c=0.00862358f \
 //x=66.565 //y=1.21 //x2=67.005 //y2=1.56
cc_4496 ( N_noxref_18_c_6388_n N_noxref_23_c_8229_n ) capacitor c=0.00124821f \
 //x=66.565 //y=0.865 //x2=67.535 //y2=0.905
cc_4497 ( N_noxref_18_c_6390_n N_noxref_23_c_8230_n ) capacitor c=0.00200715f \
 //x=66.565 //y=1.21 //x2=67.535 //y2=1.25
cc_4498 ( N_noxref_18_c_6380_n N_noxref_23_c_8231_n ) capacitor c=0.00282278f \
 //x=66.23 //y=2.08 //x2=66.97 //y2=2.08
cc_4499 ( N_noxref_18_c_6385_n N_noxref_23_c_8231_n ) capacitor c=0.0172771f \
 //x=66.035 //y=1.915 //x2=66.97 //y2=2.08
cc_4500 ( N_noxref_18_c_6380_n N_noxref_23_c_8233_n ) capacitor c=0.00342116f \
 //x=66.23 //y=2.08 //x2=67 //y2=4.7
cc_4501 ( N_noxref_18_c_6432_n N_noxref_23_c_8233_n ) capacitor c=0.0292158f \
 //x=66.23 //y=4.7 //x2=67 //y2=4.7
cc_4502 ( N_noxref_18_c_6392_n N_noxref_24_c_8424_n ) capacitor c=0.202797f \
 //x=56.12 //y=4.07 //x2=79.065 //y2=3.33
cc_4503 ( N_noxref_18_c_6449_n N_noxref_24_c_8424_n ) capacitor c=0.0136135f \
 //x=50.805 //y=4.07 //x2=79.065 //y2=3.33
cc_4504 ( N_noxref_18_c_6393_n N_noxref_24_c_8424_n ) capacitor c=0.0684106f \
 //x=66.115 //y=4.07 //x2=79.065 //y2=3.33
cc_4505 ( N_noxref_18_c_6402_n N_noxref_24_c_8424_n ) capacitor c=4.80497e-19 \
 //x=56.35 //y=4.07 //x2=79.065 //y2=3.33
cc_4506 ( N_noxref_18_c_6377_n N_noxref_24_c_8424_n ) capacitor c=0.019633f \
 //x=50.69 //y=2.08 //x2=79.065 //y2=3.33
cc_4507 ( N_noxref_18_c_6380_n N_noxref_24_c_8424_n ) capacitor c=0.0187404f \
 //x=66.23 //y=2.08 //x2=79.065 //y2=3.33
cc_4508 ( N_noxref_18_c_6456_n N_noxref_24_c_8424_n ) capacitor c=0.0187428f \
 //x=56.237 //y=3.905 //x2=79.065 //y2=3.33
cc_4509 ( N_noxref_18_c_6471_n N_noxref_45_c_10161_n ) capacitor c=0.00623646f \
 //x=50.725 //y=1.56 //x2=50.505 //y2=1.495
cc_4510 ( N_noxref_18_c_6476_n N_noxref_45_c_10161_n ) capacitor c=0.00173579f \
 //x=50.69 //y=2.08 //x2=50.505 //y2=1.495
cc_4511 ( N_noxref_18_c_6377_n N_noxref_45_c_10162_n ) capacitor c=0.00156605f \
 //x=50.69 //y=2.08 //x2=51.39 //y2=0.53
cc_4512 ( N_noxref_18_c_6466_n N_noxref_45_c_10162_n ) capacitor c=0.0188655f \
 //x=50.725 //y=0.905 //x2=51.39 //y2=0.53
cc_4513 ( N_noxref_18_c_6474_n N_noxref_45_c_10162_n ) capacitor c=0.00656458f \
 //x=51.255 //y=0.905 //x2=51.39 //y2=0.53
cc_4514 ( N_noxref_18_c_6476_n N_noxref_45_c_10162_n ) capacitor c=2.1838e-19 \
 //x=50.69 //y=2.08 //x2=51.39 //y2=0.53
cc_4515 ( N_noxref_18_c_6466_n N_noxref_45_M30_noxref_s ) capacitor \
 c=0.00623646f //x=50.725 //y=0.905 //x2=49.4 //y2=0.365
cc_4516 ( N_noxref_18_c_6474_n N_noxref_45_M30_noxref_s ) capacitor \
 c=0.0143002f //x=51.255 //y=0.905 //x2=49.4 //y2=0.365
cc_4517 ( N_noxref_18_c_6475_n N_noxref_45_M30_noxref_s ) capacitor \
 c=0.00290153f //x=51.255 //y=1.25 //x2=49.4 //y2=0.365
cc_4518 ( N_noxref_18_M34_noxref_d N_noxref_46_M32_noxref_s ) capacitor \
 c=0.00309936f //x=55.565 //y=0.915 //x2=52.625 //y2=0.375
cc_4519 ( N_noxref_18_c_6379_n N_noxref_47_c_10259_n ) capacitor c=0.00457167f \
 //x=56.155 //y=1.665 //x2=56.155 //y2=0.54
cc_4520 ( N_noxref_18_M34_noxref_d N_noxref_47_c_10259_n ) capacitor \
 c=0.0115903f //x=55.565 //y=0.915 //x2=56.155 //y2=0.54
cc_4521 ( N_noxref_18_c_6558_p N_noxref_47_c_10281_n ) capacitor c=0.0200405f \
 //x=55.84 //y=1.665 //x2=55.27 //y2=0.995
cc_4522 ( N_noxref_18_M34_noxref_d N_noxref_47_M33_noxref_d ) capacitor \
 c=5.27807e-19 //x=55.565 //y=0.915 //x2=54.03 //y2=0.91
cc_4523 ( N_noxref_18_c_6379_n N_noxref_47_M34_noxref_s ) capacitor \
 c=0.0196084f //x=56.155 //y=1.665 //x2=55.135 //y2=0.375
cc_4524 ( N_noxref_18_M34_noxref_d N_noxref_47_M34_noxref_s ) capacitor \
 c=0.0426368f //x=55.565 //y=0.915 //x2=55.135 //y2=0.375
cc_4525 ( N_noxref_18_c_6379_n N_noxref_48_c_10321_n ) capacitor c=3.83325e-19 \
 //x=56.155 //y=1.665 //x2=57.57 //y2=1.505
cc_4526 ( N_noxref_18_M34_noxref_d N_noxref_48_M35_noxref_s ) capacitor \
 c=2.55333e-19 //x=55.565 //y=0.915 //x2=57.435 //y2=0.375
cc_4527 ( N_noxref_18_c_6385_n N_noxref_51_c_10479_n ) capacitor c=0.0034165f \
 //x=66.035 //y=1.915 //x2=65.815 //y2=1.495
cc_4528 ( N_noxref_18_c_6380_n N_noxref_51_c_10461_n ) capacitor c=0.011618f \
 //x=66.23 //y=2.08 //x2=66.7 //y2=1.58
cc_4529 ( N_noxref_18_c_6384_n N_noxref_51_c_10461_n ) capacitor c=0.00696403f \
 //x=66.035 //y=1.52 //x2=66.7 //y2=1.58
cc_4530 ( N_noxref_18_c_6385_n N_noxref_51_c_10461_n ) capacitor c=0.0174694f \
 //x=66.035 //y=1.915 //x2=66.7 //y2=1.58
cc_4531 ( N_noxref_18_c_6387_n N_noxref_51_c_10461_n ) capacitor c=0.00776811f \
 //x=66.41 //y=1.365 //x2=66.7 //y2=1.58
cc_4532 ( N_noxref_18_c_6390_n N_noxref_51_c_10461_n ) capacitor c=0.00339872f \
 //x=66.565 //y=1.21 //x2=66.7 //y2=1.58
cc_4533 ( N_noxref_18_c_6385_n N_noxref_51_c_10468_n ) capacitor c=6.71402e-19 \
 //x=66.035 //y=1.915 //x2=66.785 //y2=1.495
cc_4534 ( N_noxref_18_c_6381_n N_noxref_51_M40_noxref_s ) capacitor \
 c=0.0326577f //x=66.035 //y=0.865 //x2=65.68 //y2=0.365
cc_4535 ( N_noxref_18_c_6384_n N_noxref_51_M40_noxref_s ) capacitor \
 c=3.48408e-19 //x=66.035 //y=1.52 //x2=65.68 //y2=0.365
cc_4536 ( N_noxref_18_c_6388_n N_noxref_51_M40_noxref_s ) capacitor \
 c=0.0120759f //x=66.565 //y=0.865 //x2=65.68 //y2=0.365
cc_4537 ( N_noxref_19_c_6735_p N_SN_c_6877_n ) capacitor c=0.0146822f \
 //x=67.355 //y=1.655 //x2=70.555 //y2=2.22
cc_4538 ( N_noxref_19_c_6669_n N_SN_c_6877_n ) capacitor c=0.0222456f \
 //x=67.71 //y=4.81 //x2=70.555 //y2=2.22
cc_4539 ( N_noxref_19_c_6670_n N_SN_c_6877_n ) capacitor c=0.0232665f \
 //x=69.56 //y=2.08 //x2=70.555 //y2=2.22
cc_4540 ( N_noxref_19_c_6675_n N_SN_c_6877_n ) capacitor c=0.0122202f \
 //x=69.26 //y=1.915 //x2=70.555 //y2=2.22
cc_4541 ( N_noxref_19_c_6684_n N_SN_c_6893_n ) capacitor c=0.00578357f \
 //x=69.445 //y=4.81 //x2=70.67 //y2=2.08
cc_4542 ( N_noxref_19_c_6669_n N_SN_c_6893_n ) capacitor c=3.46098e-19 \
 //x=67.71 //y=4.81 //x2=70.67 //y2=2.08
cc_4543 ( N_noxref_19_c_6670_n N_SN_c_6893_n ) capacitor c=0.0449298f \
 //x=69.56 //y=2.08 //x2=70.67 //y2=2.08
cc_4544 ( N_noxref_19_c_6675_n N_SN_c_6893_n ) capacitor c=0.00208635f \
 //x=69.26 //y=1.915 //x2=70.67 //y2=2.08
cc_4545 ( N_noxref_19_c_6743_p N_SN_c_6893_n ) capacitor c=0.00147352f \
 //x=70.125 //y=4.79 //x2=70.67 //y2=2.08
cc_4546 ( N_noxref_19_c_6713_n N_SN_c_6893_n ) capacitor c=0.00142741f \
 //x=69.835 //y=4.79 //x2=70.67 //y2=2.08
cc_4547 ( N_noxref_19_M136_noxref_g N_SN_M138_noxref_g ) capacitor c=0.010767f \
 //x=69.76 //y=6.02 //x2=70.64 //y2=6.02
cc_4548 ( N_noxref_19_M137_noxref_g N_SN_M138_noxref_g ) capacitor c=0.105888f \
 //x=70.2 //y=6.02 //x2=70.64 //y2=6.02
cc_4549 ( N_noxref_19_M137_noxref_g N_SN_M139_noxref_g ) capacitor \
 c=0.0101598f //x=70.2 //y=6.02 //x2=71.08 //y2=6.02
cc_4550 ( N_noxref_19_c_6671_n N_SN_c_7321_n ) capacitor c=5.72482e-19 \
 //x=69.26 //y=0.875 //x2=70.235 //y2=0.91
cc_4551 ( N_noxref_19_c_6673_n N_SN_c_7321_n ) capacitor c=0.00149976f \
 //x=69.26 //y=1.22 //x2=70.235 //y2=0.91
cc_4552 ( N_noxref_19_c_6678_n N_SN_c_7321_n ) capacitor c=0.0160123f \
 //x=69.79 //y=0.875 //x2=70.235 //y2=0.91
cc_4553 ( N_noxref_19_c_6674_n N_SN_c_7324_n ) capacitor c=0.00111227f \
 //x=69.26 //y=1.53 //x2=70.235 //y2=1.22
cc_4554 ( N_noxref_19_c_6680_n N_SN_c_7324_n ) capacitor c=0.0124075f \
 //x=69.79 //y=1.22 //x2=70.235 //y2=1.22
cc_4555 ( N_noxref_19_c_6678_n N_SN_c_7326_n ) capacitor c=0.00103227f \
 //x=69.79 //y=0.875 //x2=70.76 //y2=0.91
cc_4556 ( N_noxref_19_c_6680_n N_SN_c_7327_n ) capacitor c=0.0010154f \
 //x=69.79 //y=1.22 //x2=70.76 //y2=1.22
cc_4557 ( N_noxref_19_c_6680_n N_SN_c_7328_n ) capacitor c=9.23422e-19 \
 //x=69.79 //y=1.22 //x2=70.76 //y2=1.45
cc_4558 ( N_noxref_19_c_6670_n N_SN_c_7204_n ) capacitor c=0.00203769f \
 //x=69.56 //y=2.08 //x2=70.76 //y2=1.915
cc_4559 ( N_noxref_19_c_6675_n N_SN_c_7204_n ) capacitor c=0.00834532f \
 //x=69.26 //y=1.915 //x2=70.76 //y2=1.915
cc_4560 ( N_noxref_19_c_6684_n N_SN_c_7331_n ) capacitor c=2.03638e-19 \
 //x=69.445 //y=4.81 //x2=70.67 //y2=4.7
cc_4561 ( N_noxref_19_c_6670_n N_SN_c_7331_n ) capacitor c=0.00171483f \
 //x=69.56 //y=2.08 //x2=70.67 //y2=4.7
cc_4562 ( N_noxref_19_c_6743_p N_SN_c_7331_n ) capacitor c=0.0168581f \
 //x=70.125 //y=4.79 //x2=70.67 //y2=4.7
cc_4563 ( N_noxref_19_c_6713_n N_SN_c_7331_n ) capacitor c=0.00484466f \
 //x=69.835 //y=4.79 //x2=70.67 //y2=4.7
cc_4564 ( N_noxref_19_c_6684_n N_noxref_21_c_7656_n ) capacitor c=0.00623742f \
 //x=69.445 //y=4.81 //x2=71.665 //y2=3.7
cc_4565 ( N_noxref_19_c_6690_n N_noxref_21_c_7656_n ) capacitor c=5.88942e-19 \
 //x=67.825 //y=4.81 //x2=71.665 //y2=3.7
cc_4566 ( N_noxref_19_c_6698_n N_noxref_21_c_7656_n ) capacitor c=0.00902928f \
 //x=66.435 //y=5.2 //x2=71.665 //y2=3.7
cc_4567 ( N_noxref_19_c_6669_n N_noxref_21_c_7656_n ) capacitor c=0.0211071f \
 //x=67.71 //y=4.81 //x2=71.665 //y2=3.7
cc_4568 ( N_noxref_19_c_6670_n N_noxref_21_c_7656_n ) capacitor c=0.022094f \
 //x=69.56 //y=2.08 //x2=71.665 //y2=3.7
cc_4569 ( N_noxref_19_c_6669_n N_noxref_21_c_7651_n ) capacitor c=3.98811e-19 \
 //x=67.71 //y=4.81 //x2=64.38 //y2=3.7
cc_4570 ( N_noxref_19_c_6670_n N_noxref_21_c_7652_n ) capacitor c=0.00109291f \
 //x=69.56 //y=2.08 //x2=71.78 //y2=2.08
cc_4571 ( N_noxref_19_c_6684_n N_noxref_23_c_8089_n ) capacitor c=0.172728f \
 //x=69.445 //y=4.81 //x2=72.405 //y2=4.44
cc_4572 ( N_noxref_19_c_6690_n N_noxref_23_c_8089_n ) capacitor c=0.02932f \
 //x=67.825 //y=4.81 //x2=72.405 //y2=4.44
cc_4573 ( N_noxref_19_c_6694_n N_noxref_23_c_8089_n ) capacitor c=0.0156912f \
 //x=67.145 //y=5.2 //x2=72.405 //y2=4.44
cc_4574 ( N_noxref_19_c_6669_n N_noxref_23_c_8089_n ) capacitor c=0.0207668f \
 //x=67.71 //y=4.81 //x2=72.405 //y2=4.44
cc_4575 ( N_noxref_19_c_6670_n N_noxref_23_c_8089_n ) capacitor c=0.0229719f \
 //x=69.56 //y=2.08 //x2=72.405 //y2=4.44
cc_4576 ( N_noxref_19_c_6713_n N_noxref_23_c_8089_n ) capacitor c=0.0159284f \
 //x=69.835 //y=4.79 //x2=72.405 //y2=4.44
cc_4577 ( N_noxref_19_c_6694_n N_noxref_23_c_8092_n ) capacitor c=0.00319981f \
 //x=67.145 //y=5.2 //x2=67.085 //y2=4.44
cc_4578 ( N_noxref_19_c_6669_n N_noxref_23_c_8092_n ) capacitor c=0.00151334f \
 //x=67.71 //y=4.81 //x2=67.085 //y2=4.44
cc_4579 ( N_noxref_19_c_6690_n N_noxref_23_c_8213_n ) capacitor c=0.00460468f \
 //x=67.825 //y=4.81 //x2=66.97 //y2=4.535
cc_4580 ( N_noxref_19_c_6694_n N_noxref_23_c_8213_n ) capacitor c=0.0126416f \
 //x=67.145 //y=5.2 //x2=66.97 //y2=4.535
cc_4581 ( N_noxref_19_c_6669_n N_noxref_23_c_8213_n ) capacitor c=0.00799018f \
 //x=67.71 //y=4.81 //x2=66.97 //y2=4.535
cc_4582 ( N_noxref_19_c_6694_n N_noxref_23_c_8060_n ) capacitor c=3.74769e-19 \
 //x=67.145 //y=5.2 //x2=66.97 //y2=2.08
cc_4583 ( N_noxref_19_c_6669_n N_noxref_23_c_8060_n ) capacitor c=0.0707506f \
 //x=67.71 //y=4.81 //x2=66.97 //y2=2.08
cc_4584 ( N_noxref_19_c_6670_n N_noxref_23_c_8060_n ) capacitor c=7.09566e-19 \
 //x=69.56 //y=2.08 //x2=66.97 //y2=2.08
cc_4585 ( N_noxref_19_M137_noxref_g N_noxref_23_c_8111_n ) capacitor \
 c=0.0168349f //x=70.2 //y=6.02 //x2=70.775 //y2=5.155
cc_4586 ( N_noxref_19_c_6669_n N_noxref_23_c_8115_n ) capacitor c=2.97874e-19 \
 //x=67.71 //y=4.81 //x2=70.065 //y2=5.155
cc_4587 ( N_noxref_19_M136_noxref_g N_noxref_23_c_8115_n ) capacitor \
 c=0.0213876f //x=69.76 //y=6.02 //x2=70.065 //y2=5.155
cc_4588 ( N_noxref_19_c_6743_p N_noxref_23_c_8115_n ) capacitor c=0.00428486f \
 //x=70.125 //y=4.79 //x2=70.065 //y2=5.155
cc_4589 ( N_noxref_19_c_6684_n N_noxref_23_c_8126_n ) capacitor c=7.70294e-19 \
 //x=69.445 //y=4.81 //x2=72.52 //y2=4.44
cc_4590 ( N_noxref_19_c_6670_n N_noxref_23_c_8126_n ) capacitor c=6.93912e-19 \
 //x=69.56 //y=2.08 //x2=72.52 //y2=4.44
cc_4591 ( N_noxref_19_c_6694_n N_noxref_23_M134_noxref_g ) capacitor \
 c=0.0166421f //x=67.145 //y=5.2 //x2=67.01 //y2=6.02
cc_4592 ( N_noxref_19_M134_noxref_d N_noxref_23_M134_noxref_g ) capacitor \
 c=0.0173476f //x=67.085 //y=5.02 //x2=67.01 //y2=6.02
cc_4593 ( N_noxref_19_c_6690_n N_noxref_23_M135_noxref_g ) capacitor \
 c=6.16494e-19 //x=67.825 //y=4.81 //x2=67.45 //y2=6.02
cc_4594 ( N_noxref_19_c_6700_n N_noxref_23_M135_noxref_g ) capacitor \
 c=0.018922f //x=67.625 //y=5.2 //x2=67.45 //y2=6.02
cc_4595 ( N_noxref_19_M134_noxref_d N_noxref_23_M135_noxref_g ) capacitor \
 c=0.0179769f //x=67.085 //y=5.02 //x2=67.45 //y2=6.02
cc_4596 ( N_noxref_19_M41_noxref_d N_noxref_23_c_8221_n ) capacitor \
 c=0.00217566f //x=67.08 //y=0.905 //x2=67.005 //y2=0.905
cc_4597 ( N_noxref_19_M41_noxref_d N_noxref_23_c_8224_n ) capacitor \
 c=0.0034598f //x=67.08 //y=0.905 //x2=67.005 //y2=1.25
cc_4598 ( N_noxref_19_M41_noxref_d N_noxref_23_c_8226_n ) capacitor \
 c=0.00669531f //x=67.08 //y=0.905 //x2=67.005 //y2=1.56
cc_4599 ( N_noxref_19_c_6690_n N_noxref_23_c_8263_n ) capacitor c=0.00729362f \
 //x=67.825 //y=4.81 //x2=67.375 //y2=4.79
cc_4600 ( N_noxref_19_c_6669_n N_noxref_23_c_8263_n ) capacitor c=0.0118091f \
 //x=67.71 //y=4.81 //x2=67.375 //y2=4.79
cc_4601 ( N_noxref_19_c_6799_p N_noxref_23_c_8263_n ) capacitor c=0.00407665f \
 //x=67.23 //y=5.2 //x2=67.375 //y2=4.79
cc_4602 ( N_noxref_19_M41_noxref_d N_noxref_23_c_8266_n ) capacitor \
 c=0.00241102f //x=67.08 //y=0.905 //x2=67.38 //y2=0.75
cc_4603 ( N_noxref_19_c_6668_n N_noxref_23_c_8267_n ) capacitor c=0.00371277f \
 //x=67.625 //y=1.655 //x2=67.38 //y2=1.405
cc_4604 ( N_noxref_19_M41_noxref_d N_noxref_23_c_8267_n ) capacitor \
 c=0.0137169f //x=67.08 //y=0.905 //x2=67.38 //y2=1.405
cc_4605 ( N_noxref_19_M41_noxref_d N_noxref_23_c_8229_n ) capacitor \
 c=0.00132245f //x=67.08 //y=0.905 //x2=67.535 //y2=0.905
cc_4606 ( N_noxref_19_c_6668_n N_noxref_23_c_8230_n ) capacitor c=0.00457401f \
 //x=67.625 //y=1.655 //x2=67.535 //y2=1.25
cc_4607 ( N_noxref_19_M41_noxref_d N_noxref_23_c_8230_n ) capacitor \
 c=0.00566463f //x=67.08 //y=0.905 //x2=67.535 //y2=1.25
cc_4608 ( N_noxref_19_c_6669_n N_noxref_23_c_8231_n ) capacitor c=0.00709342f \
 //x=67.71 //y=4.81 //x2=66.97 //y2=2.08
cc_4609 ( N_noxref_19_c_6669_n N_noxref_23_c_8273_n ) capacitor c=0.00306024f \
 //x=67.71 //y=4.81 //x2=66.97 //y2=1.915
cc_4610 ( N_noxref_19_M41_noxref_d N_noxref_23_c_8273_n ) capacitor \
 c=0.00660593f //x=67.08 //y=0.905 //x2=66.97 //y2=1.915
cc_4611 ( N_noxref_19_c_6690_n N_noxref_23_c_8233_n ) capacitor c=4.79518e-19 \
 //x=67.825 //y=4.81 //x2=67 //y2=4.7
cc_4612 ( N_noxref_19_c_6694_n N_noxref_23_c_8233_n ) capacitor c=0.00346519f \
 //x=67.145 //y=5.2 //x2=67 //y2=4.7
cc_4613 ( N_noxref_19_c_6669_n N_noxref_23_c_8233_n ) capacitor c=0.00501989f \
 //x=67.71 //y=4.81 //x2=67 //y2=4.7
cc_4614 ( N_noxref_19_M137_noxref_g N_noxref_23_M136_noxref_d ) capacitor \
 c=0.0180032f //x=70.2 //y=6.02 //x2=69.835 //y2=5.02
cc_4615 ( N_noxref_19_c_6669_n N_noxref_24_c_8424_n ) capacitor c=0.0187691f \
 //x=67.71 //y=4.81 //x2=79.065 //y2=3.33
cc_4616 ( N_noxref_19_c_6670_n N_noxref_24_c_8424_n ) capacitor c=0.0198064f \
 //x=69.56 //y=2.08 //x2=79.065 //y2=3.33
cc_4617 ( N_noxref_19_c_6735_p N_noxref_51_c_10479_n ) capacitor c=3.15806e-19 \
 //x=67.355 //y=1.655 //x2=65.815 //y2=1.495
cc_4618 ( N_noxref_19_c_6735_p N_noxref_51_c_10468_n ) capacitor c=0.0203424f \
 //x=67.355 //y=1.655 //x2=66.785 //y2=1.495
cc_4619 ( N_noxref_19_c_6668_n N_noxref_51_c_10469_n ) capacitor c=0.00457164f \
 //x=67.625 //y=1.655 //x2=67.67 //y2=0.53
cc_4620 ( N_noxref_19_M41_noxref_d N_noxref_51_c_10469_n ) capacitor \
 c=0.0115831f //x=67.08 //y=0.905 //x2=67.67 //y2=0.53
cc_4621 ( N_noxref_19_c_6668_n N_noxref_51_M40_noxref_s ) capacitor \
 c=0.013435f //x=67.625 //y=1.655 //x2=65.68 //y2=0.365
cc_4622 ( N_noxref_19_M41_noxref_d N_noxref_51_M40_noxref_s ) capacitor \
 c=0.043966f //x=67.08 //y=0.905 //x2=65.68 //y2=0.365
cc_4623 ( N_noxref_19_c_6668_n N_noxref_52_c_10529_n ) capacitor c=4.08644e-19 \
 //x=67.625 //y=1.655 //x2=69.04 //y2=1.505
cc_4624 ( N_noxref_19_c_6675_n N_noxref_52_c_10529_n ) capacitor c=0.0034165f \
 //x=69.26 //y=1.915 //x2=69.04 //y2=1.505
cc_4625 ( N_noxref_19_c_6670_n N_noxref_52_c_10512_n ) capacitor c=0.0115611f \
 //x=69.56 //y=2.08 //x2=69.925 //y2=1.59
cc_4626 ( N_noxref_19_c_6674_n N_noxref_52_c_10512_n ) capacitor c=0.00697148f \
 //x=69.26 //y=1.53 //x2=69.925 //y2=1.59
cc_4627 ( N_noxref_19_c_6675_n N_noxref_52_c_10512_n ) capacitor c=0.0204849f \
 //x=69.26 //y=1.915 //x2=69.925 //y2=1.59
cc_4628 ( N_noxref_19_c_6677_n N_noxref_52_c_10512_n ) capacitor c=0.00610316f \
 //x=69.635 //y=1.375 //x2=69.925 //y2=1.59
cc_4629 ( N_noxref_19_c_6680_n N_noxref_52_c_10512_n ) capacitor c=0.00698822f \
 //x=69.79 //y=1.22 //x2=69.925 //y2=1.59
cc_4630 ( N_noxref_19_c_6671_n N_noxref_52_M42_noxref_s ) capacitor \
 c=0.0327271f //x=69.26 //y=0.875 //x2=68.905 //y2=0.375
cc_4631 ( N_noxref_19_c_6674_n N_noxref_52_M42_noxref_s ) capacitor \
 c=7.99997e-19 //x=69.26 //y=1.53 //x2=68.905 //y2=0.375
cc_4632 ( N_noxref_19_c_6675_n N_noxref_52_M42_noxref_s ) capacitor \
 c=0.00122123f //x=69.26 //y=1.915 //x2=68.905 //y2=0.375
cc_4633 ( N_noxref_19_c_6678_n N_noxref_52_M42_noxref_s ) capacitor \
 c=0.0121427f //x=69.79 //y=0.875 //x2=68.905 //y2=0.375
cc_4634 ( N_noxref_19_M41_noxref_d N_noxref_52_M42_noxref_s ) capacitor \
 c=2.53688e-19 //x=67.08 //y=0.905 //x2=68.905 //y2=0.375
cc_4635 ( N_SN_c_6892_n N_noxref_21_c_7696_n ) capacitor c=0.0190398f //x=59.2 \
 //y=2.08 //x2=60.195 //y2=3.7
cc_4636 ( N_SN_c_6892_n N_noxref_21_c_7699_n ) capacitor c=0.00128547f \
 //x=59.2 //y=2.08 //x2=60.425 //y2=3.7
cc_4637 ( N_SN_c_6893_n N_noxref_21_c_7656_n ) capacitor c=0.0226304f \
 //x=70.67 //y=2.08 //x2=71.665 //y2=3.7
cc_4638 ( N_SN_c_6866_n N_noxref_21_c_7648_n ) capacitor c=0.0186201f \
 //x=59.085 //y=2.22 //x2=55.5 //y2=2.08
cc_4639 ( N_SN_c_6877_n N_noxref_21_c_7649_n ) capacitor c=0.0209607f \
 //x=70.555 //y=2.22 //x2=60.31 //y2=2.08
cc_4640 ( N_SN_c_6887_n N_noxref_21_c_7649_n ) capacitor c=0.00165648f \
 //x=59.315 //y=2.22 //x2=60.31 //y2=2.08
cc_4641 ( N_SN_c_6892_n N_noxref_21_c_7649_n ) capacitor c=0.0433248f //x=59.2 \
 //y=2.08 //x2=60.31 //y2=2.08
cc_4642 ( N_SN_c_7252_n N_noxref_21_c_7649_n ) capacitor c=0.00205895f \
 //x=59.29 //y=1.915 //x2=60.31 //y2=2.08
cc_4643 ( N_SN_c_7254_n N_noxref_21_c_7649_n ) capacitor c=0.00142741f \
 //x=59.2 //y=4.7 //x2=60.31 //y2=2.08
cc_4644 ( N_SN_c_6877_n N_noxref_21_c_7858_n ) capacitor c=0.0146822f \
 //x=70.555 //y=2.22 //x2=64.025 //y2=1.655
cc_4645 ( N_SN_c_6877_n N_noxref_21_c_7651_n ) capacitor c=0.0222456f \
 //x=70.555 //y=2.22 //x2=64.38 //y2=3.7
cc_4646 ( N_SN_c_6877_n N_noxref_21_c_7652_n ) capacitor c=0.00558344f \
 //x=70.555 //y=2.22 //x2=71.78 //y2=2.08
cc_4647 ( N_SN_c_6893_n N_noxref_21_c_7652_n ) capacitor c=0.0466321f \
 //x=70.67 //y=2.08 //x2=71.78 //y2=2.08
cc_4648 ( N_SN_c_7204_n N_noxref_21_c_7652_n ) capacitor c=0.00213841f \
 //x=70.76 //y=1.915 //x2=71.78 //y2=2.08
cc_4649 ( N_SN_c_7331_n N_noxref_21_c_7652_n ) capacitor c=0.00142741f \
 //x=70.67 //y=4.7 //x2=71.78 //y2=2.08
cc_4650 ( N_SN_M124_noxref_g N_noxref_21_M126_noxref_g ) capacitor \
 c=0.0101598f //x=59.17 //y=6.02 //x2=60.05 //y2=6.02
cc_4651 ( N_SN_M125_noxref_g N_noxref_21_M126_noxref_g ) capacitor \
 c=0.0602553f //x=59.61 //y=6.02 //x2=60.05 //y2=6.02
cc_4652 ( N_SN_M125_noxref_g N_noxref_21_M127_noxref_g ) capacitor \
 c=0.0101598f //x=59.61 //y=6.02 //x2=60.49 //y2=6.02
cc_4653 ( N_SN_M138_noxref_g N_noxref_21_M140_noxref_g ) capacitor \
 c=0.0101598f //x=70.64 //y=6.02 //x2=71.52 //y2=6.02
cc_4654 ( N_SN_M139_noxref_g N_noxref_21_M140_noxref_g ) capacitor \
 c=0.0602553f //x=71.08 //y=6.02 //x2=71.52 //y2=6.02
cc_4655 ( N_SN_M139_noxref_g N_noxref_21_M141_noxref_g ) capacitor \
 c=0.0101598f //x=71.08 //y=6.02 //x2=71.96 //y2=6.02
cc_4656 ( N_SN_c_6866_n N_noxref_21_c_7831_n ) capacitor c=3.13485e-19 \
 //x=59.085 //y=2.22 //x2=55.865 //y2=1.415
cc_4657 ( N_SN_c_7249_n N_noxref_21_c_7729_n ) capacitor c=0.00456962f \
 //x=59.29 //y=0.91 //x2=60.3 //y2=0.915
cc_4658 ( N_SN_c_7250_n N_noxref_21_c_7730_n ) capacitor c=0.00438372f \
 //x=59.29 //y=1.22 //x2=60.3 //y2=1.26
cc_4659 ( N_SN_c_7251_n N_noxref_21_c_7731_n ) capacitor c=0.00438372f \
 //x=59.29 //y=1.45 //x2=60.3 //y2=1.57
cc_4660 ( N_SN_c_6877_n N_noxref_21_c_7733_n ) capacitor c=3.13485e-19 \
 //x=70.555 //y=2.22 //x2=60.675 //y2=1.415
cc_4661 ( N_SN_c_7326_n N_noxref_21_c_7875_n ) capacitor c=0.00456962f \
 //x=70.76 //y=0.91 //x2=71.77 //y2=0.915
cc_4662 ( N_SN_c_7327_n N_noxref_21_c_7876_n ) capacitor c=0.00438372f \
 //x=70.76 //y=1.22 //x2=71.77 //y2=1.26
cc_4663 ( N_SN_c_7328_n N_noxref_21_c_7877_n ) capacitor c=0.00438372f \
 //x=70.76 //y=1.45 //x2=71.77 //y2=1.57
cc_4664 ( N_SN_c_6866_n N_noxref_21_c_7781_n ) capacitor c=0.00584491f \
 //x=59.085 //y=2.22 //x2=55.5 //y2=2.08
cc_4665 ( N_SN_c_6877_n N_noxref_21_c_7738_n ) capacitor c=0.00584491f \
 //x=70.555 //y=2.22 //x2=60.31 //y2=2.08
cc_4666 ( N_SN_c_6887_n N_noxref_21_c_7738_n ) capacitor c=2.3323e-19 \
 //x=59.315 //y=2.22 //x2=60.31 //y2=2.08
cc_4667 ( N_SN_c_6892_n N_noxref_21_c_7738_n ) capacitor c=0.0019893f //x=59.2 \
 //y=2.08 //x2=60.31 //y2=2.08
cc_4668 ( N_SN_c_7252_n N_noxref_21_c_7738_n ) capacitor c=0.00828003f \
 //x=59.29 //y=1.915 //x2=60.31 //y2=2.08
cc_4669 ( N_SN_c_7252_n N_noxref_21_c_7739_n ) capacitor c=0.00438372f \
 //x=59.29 //y=1.915 //x2=60.31 //y2=1.915
cc_4670 ( N_SN_c_6892_n N_noxref_21_c_7741_n ) capacitor c=0.00219458f \
 //x=59.2 //y=2.08 //x2=60.31 //y2=4.7
cc_4671 ( N_SN_c_7269_n N_noxref_21_c_7741_n ) capacitor c=0.0611812f \
 //x=59.535 //y=4.79 //x2=60.31 //y2=4.7
cc_4672 ( N_SN_c_7254_n N_noxref_21_c_7741_n ) capacitor c=0.00487508f \
 //x=59.2 //y=4.7 //x2=60.31 //y2=4.7
cc_4673 ( N_SN_c_6877_n N_noxref_21_c_7706_n ) capacitor c=0.00341397f \
 //x=70.555 //y=2.22 //x2=71.78 //y2=2.08
cc_4674 ( N_SN_c_6893_n N_noxref_21_c_7706_n ) capacitor c=0.0021852f \
 //x=70.67 //y=2.08 //x2=71.78 //y2=2.08
cc_4675 ( N_SN_c_7204_n N_noxref_21_c_7706_n ) capacitor c=0.00896806f \
 //x=70.76 //y=1.915 //x2=71.78 //y2=2.08
cc_4676 ( N_SN_c_7204_n N_noxref_21_c_7890_n ) capacitor c=0.00438372f \
 //x=70.76 //y=1.915 //x2=71.78 //y2=1.915
cc_4677 ( N_SN_c_6893_n N_noxref_21_c_7891_n ) capacitor c=0.00219458f \
 //x=70.67 //y=2.08 //x2=71.78 //y2=4.7
cc_4678 ( N_SN_c_7378_p N_noxref_21_c_7891_n ) capacitor c=0.0611812f \
 //x=71.005 //y=4.79 //x2=71.78 //y2=4.7
cc_4679 ( N_SN_c_7331_n N_noxref_21_c_7891_n ) capacitor c=0.00487508f \
 //x=70.67 //y=4.7 //x2=71.78 //y2=4.7
cc_4680 ( N_SN_c_6893_n N_noxref_23_c_8089_n ) capacitor c=0.0233868f \
 //x=70.67 //y=2.08 //x2=72.405 //y2=4.44
cc_4681 ( N_SN_c_7378_p N_noxref_23_c_8089_n ) capacitor c=0.0085986f \
 //x=71.005 //y=4.79 //x2=72.405 //y2=4.44
cc_4682 ( N_SN_c_7331_n N_noxref_23_c_8089_n ) capacitor c=0.00293313f \
 //x=70.67 //y=4.7 //x2=72.405 //y2=4.44
cc_4683 ( N_SN_c_6877_n N_noxref_23_c_8060_n ) capacitor c=0.0201924f \
 //x=70.555 //y=2.22 //x2=66.97 //y2=2.08
cc_4684 ( N_SN_c_6893_n N_noxref_23_c_8111_n ) capacitor c=0.0144268f \
 //x=70.67 //y=2.08 //x2=70.775 //y2=5.155
cc_4685 ( N_SN_M138_noxref_g N_noxref_23_c_8111_n ) capacitor c=0.0165266f \
 //x=70.64 //y=6.02 //x2=70.775 //y2=5.155
cc_4686 ( N_SN_c_7331_n N_noxref_23_c_8111_n ) capacitor c=0.00322054f \
 //x=70.67 //y=4.7 //x2=70.775 //y2=5.155
cc_4687 ( N_SN_M139_noxref_g N_noxref_23_c_8117_n ) capacitor c=0.01736f \
 //x=71.08 //y=6.02 //x2=71.655 //y2=5.155
cc_4688 ( N_SN_c_6893_n N_noxref_23_c_8126_n ) capacitor c=0.00300717f \
 //x=70.67 //y=2.08 //x2=72.52 //y2=4.44
cc_4689 ( N_SN_c_7378_p N_noxref_23_c_8288_n ) capacitor c=0.00426767f \
 //x=71.005 //y=4.79 //x2=70.86 //y2=5.155
cc_4690 ( N_SN_c_6877_n N_noxref_23_c_8267_n ) capacitor c=3.11115e-19 \
 //x=70.555 //y=2.22 //x2=67.38 //y2=1.405
cc_4691 ( N_SN_c_6877_n N_noxref_23_c_8231_n ) capacitor c=0.00568402f \
 //x=70.555 //y=2.22 //x2=66.97 //y2=2.08
cc_4692 ( N_SN_M138_noxref_g N_noxref_23_M138_noxref_d ) capacitor \
 c=0.0180032f //x=70.64 //y=6.02 //x2=70.715 //y2=5.02
cc_4693 ( N_SN_M139_noxref_g N_noxref_23_M138_noxref_d ) capacitor \
 c=0.0180032f //x=71.08 //y=6.02 //x2=70.715 //y2=5.02
cc_4694 ( N_SN_c_6833_n N_noxref_24_c_8520_n ) capacitor c=0.0205469f \
 //x=21.715 //y=2.22 //x2=23.565 //y2=3.33
cc_4695 ( N_SN_c_6844_n N_noxref_24_c_8520_n ) capacitor c=0.011348f \
 //x=34.665 //y=2.22 //x2=23.565 //y2=3.33
cc_4696 ( N_SN_c_6854_n N_noxref_24_c_8520_n ) capacitor c=4.81986e-19 \
 //x=21.945 //y=2.22 //x2=23.565 //y2=3.33
cc_4697 ( N_SN_c_6889_n N_noxref_24_c_8520_n ) capacitor c=0.0190562f \
 //x=21.83 //y=2.08 //x2=23.565 //y2=3.33
cc_4698 ( N_SN_c_6833_n N_noxref_24_c_8497_n ) capacitor c=7.29504e-19 \
 //x=21.715 //y=2.22 //x2=18.245 //y2=3.33
cc_4699 ( N_SN_c_6844_n N_noxref_24_c_8424_n ) capacitor c=0.0245103f \
 //x=34.665 //y=2.22 //x2=79.065 //y2=3.33
cc_4700 ( N_SN_c_6855_n N_noxref_24_c_8424_n ) capacitor c=0.0442417f \
 //x=46.135 //y=2.22 //x2=79.065 //y2=3.33
cc_4701 ( N_SN_c_6865_n N_noxref_24_c_8424_n ) capacitor c=4.81986e-19 \
 //x=34.895 //y=2.22 //x2=79.065 //y2=3.33
cc_4702 ( N_SN_c_6866_n N_noxref_24_c_8424_n ) capacitor c=0.0254299f \
 //x=59.085 //y=2.22 //x2=79.065 //y2=3.33
cc_4703 ( N_SN_c_6876_n N_noxref_24_c_8424_n ) capacitor c=4.81986e-19 \
 //x=46.365 //y=2.22 //x2=79.065 //y2=3.33
cc_4704 ( N_SN_c_6877_n N_noxref_24_c_8424_n ) capacitor c=0.0554412f \
 //x=70.555 //y=2.22 //x2=79.065 //y2=3.33
cc_4705 ( N_SN_c_6887_n N_noxref_24_c_8424_n ) capacitor c=4.81986e-19 \
 //x=59.315 //y=2.22 //x2=79.065 //y2=3.33
cc_4706 ( N_SN_c_6890_n N_noxref_24_c_8424_n ) capacitor c=0.0190562f \
 //x=34.78 //y=2.08 //x2=79.065 //y2=3.33
cc_4707 ( N_SN_c_6891_n N_noxref_24_c_8424_n ) capacitor c=0.0190562f \
 //x=46.25 //y=2.08 //x2=79.065 //y2=3.33
cc_4708 ( N_SN_c_6892_n N_noxref_24_c_8424_n ) capacitor c=0.0190562f //x=59.2 \
 //y=2.08 //x2=79.065 //y2=3.33
cc_4709 ( N_SN_c_6893_n N_noxref_24_c_8424_n ) capacitor c=0.0190562f \
 //x=70.67 //y=2.08 //x2=79.065 //y2=3.33
cc_4710 ( N_SN_c_6844_n N_noxref_24_c_8558_n ) capacitor c=4.49298e-19 \
 //x=34.665 //y=2.22 //x2=23.795 //y2=3.33
cc_4711 ( N_SN_c_6833_n N_noxref_24_c_8428_n ) capacitor c=0.0201924f \
 //x=21.715 //y=2.22 //x2=18.13 //y2=2.08
cc_4712 ( N_SN_c_6889_n N_noxref_24_c_8451_n ) capacitor c=0.0144268f \
 //x=21.83 //y=2.08 //x2=21.935 //y2=5.155
cc_4713 ( N_SN_M78_noxref_g N_noxref_24_c_8451_n ) capacitor c=0.0165266f \
 //x=21.8 //y=6.02 //x2=21.935 //y2=5.155
cc_4714 ( N_SN_c_6996_n N_noxref_24_c_8451_n ) capacitor c=0.00322054f \
 //x=21.83 //y=4.7 //x2=21.935 //y2=5.155
cc_4715 ( N_SN_M79_noxref_g N_noxref_24_c_8457_n ) capacitor c=0.01736f \
 //x=22.24 //y=6.02 //x2=22.815 //y2=5.155
cc_4716 ( N_SN_c_6844_n N_noxref_24_c_8735_n ) capacitor c=0.016327f \
 //x=34.665 //y=2.22 //x2=23.28 //y2=1.665
cc_4717 ( N_SN_c_6844_n N_noxref_24_c_8465_n ) capacitor c=0.0220713f \
 //x=34.665 //y=2.22 //x2=23.68 //y2=3.33
cc_4718 ( N_SN_c_6889_n N_noxref_24_c_8465_n ) capacitor c=0.00303929f \
 //x=21.83 //y=2.08 //x2=23.68 //y2=3.33
cc_4719 ( N_SN_c_7045_n N_noxref_24_c_8738_n ) capacitor c=0.00426767f \
 //x=22.165 //y=4.79 //x2=22.02 //y2=5.155
cc_4720 ( N_SN_c_6833_n N_noxref_24_c_8544_n ) capacitor c=3.11115e-19 \
 //x=21.715 //y=2.22 //x2=18.54 //y2=1.405
cc_4721 ( N_SN_c_6833_n N_noxref_24_c_8516_n ) capacitor c=0.00570799f \
 //x=21.715 //y=2.22 //x2=18.13 //y2=2.08
cc_4722 ( N_SN_M78_noxref_g N_noxref_24_M78_noxref_d ) capacitor c=0.0180032f \
 //x=21.8 //y=6.02 //x2=21.875 //y2=5.02
cc_4723 ( N_SN_M79_noxref_g N_noxref_24_M78_noxref_d ) capacitor c=0.0180032f \
 //x=22.24 //y=6.02 //x2=21.875 //y2=5.02
cc_4724 ( N_SN_c_6940_n N_noxref_30_c_9388_n ) capacitor c=0.0167228f \
 //x=9.925 //y=0.91 //x2=10.585 //y2=0.54
cc_4725 ( N_SN_c_6945_n N_noxref_30_c_9388_n ) capacitor c=0.00534519f \
 //x=10.45 //y=0.91 //x2=10.585 //y2=0.54
cc_4726 ( N_SN_c_6833_n N_noxref_30_c_9412_n ) capacitor c=0.00387656f \
 //x=21.715 //y=2.22 //x2=10.585 //y2=1.59
cc_4727 ( N_SN_c_6843_n N_noxref_30_c_9412_n ) capacitor c=0.00354473f \
 //x=10.475 //y=2.22 //x2=10.585 //y2=1.59
cc_4728 ( N_SN_c_6888_n N_noxref_30_c_9412_n ) capacitor c=0.011736f //x=10.36 \
 //y=2.08 //x2=10.585 //y2=1.59
cc_4729 ( N_SN_c_6943_n N_noxref_30_c_9412_n ) capacitor c=0.0153695f \
 //x=9.925 //y=1.22 //x2=10.585 //y2=1.59
cc_4730 ( N_SN_c_6948_n N_noxref_30_c_9412_n ) capacitor c=0.0213278f \
 //x=10.45 //y=1.915 //x2=10.585 //y2=1.59
cc_4731 ( N_SN_c_6833_n N_noxref_30_M5_noxref_s ) capacitor c=0.00599513f \
 //x=21.715 //y=2.22 //x2=8.595 //y2=0.375
cc_4732 ( N_SN_c_6940_n N_noxref_30_M5_noxref_s ) capacitor c=0.00798959f \
 //x=9.925 //y=0.91 //x2=8.595 //y2=0.375
cc_4733 ( N_SN_c_6947_n N_noxref_30_M5_noxref_s ) capacitor c=0.00212176f \
 //x=10.45 //y=1.45 //x2=8.595 //y2=0.375
cc_4734 ( N_SN_c_6948_n N_noxref_30_M5_noxref_s ) capacitor c=0.00298115f \
 //x=10.45 //y=1.915 //x2=8.595 //y2=0.375
cc_4735 ( N_SN_c_6833_n N_noxref_31_c_9434_n ) capacitor c=0.00657782f \
 //x=21.715 //y=2.22 //x2=11.155 //y2=0.995
cc_4736 ( N_SN_c_7436_p N_noxref_31_c_9434_n ) capacitor c=2.14837e-19 \
 //x=10.295 //y=0.755 //x2=11.155 //y2=0.995
cc_4737 ( N_SN_c_6945_n N_noxref_31_c_9434_n ) capacitor c=0.00123426f \
 //x=10.45 //y=0.91 //x2=11.155 //y2=0.995
cc_4738 ( N_SN_c_6946_n N_noxref_31_c_9434_n ) capacitor c=0.0129288f \
 //x=10.45 //y=1.22 //x2=11.155 //y2=0.995
cc_4739 ( N_SN_c_6947_n N_noxref_31_c_9434_n ) capacitor c=0.00142359f \
 //x=10.45 //y=1.45 //x2=11.155 //y2=0.995
cc_4740 ( N_SN_c_6833_n N_noxref_31_c_9439_n ) capacitor c=0.00147946f \
 //x=21.715 //y=2.22 //x2=12.125 //y2=0.54
cc_4741 ( N_SN_c_6940_n N_noxref_31_M6_noxref_d ) capacitor c=0.00223875f \
 //x=9.925 //y=0.91 //x2=10 //y2=0.91
cc_4742 ( N_SN_c_6943_n N_noxref_31_M6_noxref_d ) capacitor c=0.00262485f \
 //x=9.925 //y=1.22 //x2=10 //y2=0.91
cc_4743 ( N_SN_c_7436_p N_noxref_31_M6_noxref_d ) capacitor c=0.00220746f \
 //x=10.295 //y=0.755 //x2=10 //y2=0.91
cc_4744 ( N_SN_c_7444_p N_noxref_31_M6_noxref_d ) capacitor c=0.00194798f \
 //x=10.295 //y=1.375 //x2=10 //y2=0.91
cc_4745 ( N_SN_c_6945_n N_noxref_31_M6_noxref_d ) capacitor c=0.00198465f \
 //x=10.45 //y=0.91 //x2=10 //y2=0.91
cc_4746 ( N_SN_c_6946_n N_noxref_31_M6_noxref_d ) capacitor c=0.00128384f \
 //x=10.45 //y=1.22 //x2=10 //y2=0.91
cc_4747 ( N_SN_c_6833_n N_noxref_31_M7_noxref_s ) capacitor c=0.00642985f \
 //x=21.715 //y=2.22 //x2=11.105 //y2=0.375
cc_4748 ( N_SN_c_6945_n N_noxref_31_M7_noxref_s ) capacitor c=7.21316e-19 \
 //x=10.45 //y=0.91 //x2=11.105 //y2=0.375
cc_4749 ( N_SN_c_6946_n N_noxref_31_M7_noxref_s ) capacitor c=0.00348171f \
 //x=10.45 //y=1.22 //x2=11.105 //y2=0.375
cc_4750 ( N_SN_c_6833_n N_noxref_32_c_9504_n ) capacitor c=0.00635755f \
 //x=21.715 //y=2.22 //x2=13.645 //y2=1.495
cc_4751 ( N_SN_c_6833_n N_noxref_32_c_9486_n ) capacitor c=0.0223494f \
 //x=21.715 //y=2.22 //x2=14.53 //y2=1.58
cc_4752 ( N_SN_c_6833_n N_noxref_32_c_9493_n ) capacitor c=0.00649228f \
 //x=21.715 //y=2.22 //x2=14.615 //y2=1.495
cc_4753 ( N_SN_c_6833_n N_noxref_32_c_9494_n ) capacitor c=0.00178534f \
 //x=21.715 //y=2.22 //x2=15.5 //y2=0.53
cc_4754 ( N_SN_c_6833_n N_noxref_32_M8_noxref_s ) capacitor c=0.00113237f \
 //x=21.715 //y=2.22 //x2=13.51 //y2=0.365
cc_4755 ( N_SN_c_6833_n N_noxref_33_c_9555_n ) capacitor c=0.00635755f \
 //x=21.715 //y=2.22 //x2=16.975 //y2=1.495
cc_4756 ( N_SN_c_6833_n N_noxref_33_c_9537_n ) capacitor c=0.0223494f \
 //x=21.715 //y=2.22 //x2=17.86 //y2=1.58
cc_4757 ( N_SN_c_6833_n N_noxref_33_c_9544_n ) capacitor c=0.00649228f \
 //x=21.715 //y=2.22 //x2=17.945 //y2=1.495
cc_4758 ( N_SN_c_6833_n N_noxref_33_c_9545_n ) capacitor c=0.00178534f \
 //x=21.715 //y=2.22 //x2=18.83 //y2=0.53
cc_4759 ( N_SN_c_6833_n N_noxref_33_M10_noxref_s ) capacitor c=0.00113237f \
 //x=21.715 //y=2.22 //x2=16.84 //y2=0.365
cc_4760 ( N_SN_c_6833_n N_noxref_34_c_9603_n ) capacitor c=0.00642985f \
 //x=21.715 //y=2.22 //x2=20.2 //y2=1.505
cc_4761 ( N_SN_c_6833_n N_noxref_34_c_9588_n ) capacitor c=0.0225733f \
 //x=21.715 //y=2.22 //x2=21.085 //y2=1.59
cc_4762 ( N_SN_c_6986_n N_noxref_34_c_9595_n ) capacitor c=0.0167228f \
 //x=21.395 //y=0.91 //x2=22.055 //y2=0.54
cc_4763 ( N_SN_c_6991_n N_noxref_34_c_9595_n ) capacitor c=0.00534519f \
 //x=21.92 //y=0.91 //x2=22.055 //y2=0.54
cc_4764 ( N_SN_c_6833_n N_noxref_34_c_9619_n ) capacitor c=0.0139868f \
 //x=21.715 //y=2.22 //x2=22.055 //y2=1.59
cc_4765 ( N_SN_c_6844_n N_noxref_34_c_9619_n ) capacitor c=0.00387656f \
 //x=34.665 //y=2.22 //x2=22.055 //y2=1.59
cc_4766 ( N_SN_c_6854_n N_noxref_34_c_9619_n ) capacitor c=0.00251375f \
 //x=21.945 //y=2.22 //x2=22.055 //y2=1.59
cc_4767 ( N_SN_c_6889_n N_noxref_34_c_9619_n ) capacitor c=0.011736f //x=21.83 \
 //y=2.08 //x2=22.055 //y2=1.59
cc_4768 ( N_SN_c_6989_n N_noxref_34_c_9619_n ) capacitor c=0.0157358f \
 //x=21.395 //y=1.22 //x2=22.055 //y2=1.59
cc_4769 ( N_SN_c_6994_n N_noxref_34_c_9619_n ) capacitor c=0.0213278f \
 //x=21.92 //y=1.915 //x2=22.055 //y2=1.59
cc_4770 ( N_SN_c_6833_n N_noxref_34_M12_noxref_s ) capacitor c=0.00642985f \
 //x=21.715 //y=2.22 //x2=20.065 //y2=0.375
cc_4771 ( N_SN_c_6844_n N_noxref_34_M12_noxref_s ) capacitor c=0.00599513f \
 //x=34.665 //y=2.22 //x2=20.065 //y2=0.375
cc_4772 ( N_SN_c_6986_n N_noxref_34_M12_noxref_s ) capacitor c=0.00798959f \
 //x=21.395 //y=0.91 //x2=20.065 //y2=0.375
cc_4773 ( N_SN_c_6993_n N_noxref_34_M12_noxref_s ) capacitor c=0.00212176f \
 //x=21.92 //y=1.45 //x2=20.065 //y2=0.375
cc_4774 ( N_SN_c_6994_n N_noxref_34_M12_noxref_s ) capacitor c=0.00298115f \
 //x=21.92 //y=1.915 //x2=20.065 //y2=0.375
cc_4775 ( N_SN_c_6844_n N_noxref_35_c_9640_n ) capacitor c=0.00657782f \
 //x=34.665 //y=2.22 //x2=22.625 //y2=0.995
cc_4776 ( N_SN_c_7476_p N_noxref_35_c_9640_n ) capacitor c=2.14837e-19 \
 //x=21.765 //y=0.755 //x2=22.625 //y2=0.995
cc_4777 ( N_SN_c_6991_n N_noxref_35_c_9640_n ) capacitor c=0.00123426f \
 //x=21.92 //y=0.91 //x2=22.625 //y2=0.995
cc_4778 ( N_SN_c_6992_n N_noxref_35_c_9640_n ) capacitor c=0.0129288f \
 //x=21.92 //y=1.22 //x2=22.625 //y2=0.995
cc_4779 ( N_SN_c_6993_n N_noxref_35_c_9640_n ) capacitor c=0.00142359f \
 //x=21.92 //y=1.45 //x2=22.625 //y2=0.995
cc_4780 ( N_SN_c_6844_n N_noxref_35_c_9645_n ) capacitor c=0.00147946f \
 //x=34.665 //y=2.22 //x2=23.595 //y2=0.54
cc_4781 ( N_SN_c_6986_n N_noxref_35_M13_noxref_d ) capacitor c=0.00223875f \
 //x=21.395 //y=0.91 //x2=21.47 //y2=0.91
cc_4782 ( N_SN_c_6989_n N_noxref_35_M13_noxref_d ) capacitor c=0.00262485f \
 //x=21.395 //y=1.22 //x2=21.47 //y2=0.91
cc_4783 ( N_SN_c_7476_p N_noxref_35_M13_noxref_d ) capacitor c=0.00220746f \
 //x=21.765 //y=0.755 //x2=21.47 //y2=0.91
cc_4784 ( N_SN_c_7484_p N_noxref_35_M13_noxref_d ) capacitor c=0.00194798f \
 //x=21.765 //y=1.375 //x2=21.47 //y2=0.91
cc_4785 ( N_SN_c_6991_n N_noxref_35_M13_noxref_d ) capacitor c=0.00198465f \
 //x=21.92 //y=0.91 //x2=21.47 //y2=0.91
cc_4786 ( N_SN_c_6992_n N_noxref_35_M13_noxref_d ) capacitor c=0.00128384f \
 //x=21.92 //y=1.22 //x2=21.47 //y2=0.91
cc_4787 ( N_SN_c_6844_n N_noxref_35_M14_noxref_s ) capacitor c=0.00642985f \
 //x=34.665 //y=2.22 //x2=22.575 //y2=0.375
cc_4788 ( N_SN_c_6991_n N_noxref_35_M14_noxref_s ) capacitor c=7.21316e-19 \
 //x=21.92 //y=0.91 //x2=22.575 //y2=0.375
cc_4789 ( N_SN_c_6992_n N_noxref_35_M14_noxref_s ) capacitor c=0.00348171f \
 //x=21.92 //y=1.22 //x2=22.575 //y2=0.375
cc_4790 ( N_SN_c_6844_n N_noxref_36_c_9710_n ) capacitor c=0.00635755f \
 //x=34.665 //y=2.22 //x2=25.115 //y2=1.495
cc_4791 ( N_SN_c_6844_n N_noxref_36_c_9692_n ) capacitor c=0.0223494f \
 //x=34.665 //y=2.22 //x2=26 //y2=1.58
cc_4792 ( N_SN_c_6844_n N_noxref_36_c_9699_n ) capacitor c=0.00649228f \
 //x=34.665 //y=2.22 //x2=26.085 //y2=1.495
cc_4793 ( N_SN_c_6844_n N_noxref_36_c_9700_n ) capacitor c=0.00178534f \
 //x=34.665 //y=2.22 //x2=26.97 //y2=0.53
cc_4794 ( N_SN_c_6844_n N_noxref_36_M15_noxref_s ) capacitor c=0.00113237f \
 //x=34.665 //y=2.22 //x2=24.98 //y2=0.365
cc_4795 ( N_SN_c_6844_n N_noxref_37_c_9758_n ) capacitor c=0.00642985f \
 //x=34.665 //y=2.22 //x2=28.34 //y2=1.505
cc_4796 ( N_SN_c_6844_n N_noxref_37_c_9743_n ) capacitor c=0.0225733f \
 //x=34.665 //y=2.22 //x2=29.225 //y2=1.59
cc_4797 ( N_SN_c_6844_n N_noxref_37_c_9773_n ) capacitor c=0.0203655f \
 //x=34.665 //y=2.22 //x2=30.195 //y2=1.59
cc_4798 ( N_SN_c_6844_n N_noxref_37_M17_noxref_s ) capacitor c=0.012425f \
 //x=34.665 //y=2.22 //x2=28.205 //y2=0.375
cc_4799 ( N_SN_c_6844_n N_noxref_38_c_9792_n ) capacitor c=0.00657782f \
 //x=34.665 //y=2.22 //x2=30.765 //y2=0.995
cc_4800 ( N_SN_c_6844_n N_noxref_38_c_9797_n ) capacitor c=0.00147946f \
 //x=34.665 //y=2.22 //x2=31.735 //y2=0.54
cc_4801 ( N_SN_c_6844_n N_noxref_38_M19_noxref_s ) capacitor c=0.00642985f \
 //x=34.665 //y=2.22 //x2=30.715 //y2=0.375
cc_4802 ( N_SN_c_6844_n N_noxref_39_c_9859_n ) capacitor c=0.00642985f \
 //x=34.665 //y=2.22 //x2=33.15 //y2=1.505
cc_4803 ( N_SN_c_6844_n N_noxref_39_c_9844_n ) capacitor c=0.0225733f \
 //x=34.665 //y=2.22 //x2=34.035 //y2=1.59
cc_4804 ( N_SN_c_7070_n N_noxref_39_c_9851_n ) capacitor c=0.0167228f \
 //x=34.345 //y=0.91 //x2=35.005 //y2=0.54
cc_4805 ( N_SN_c_7075_n N_noxref_39_c_9851_n ) capacitor c=0.00534519f \
 //x=34.87 //y=0.91 //x2=35.005 //y2=0.54
cc_4806 ( N_SN_c_6844_n N_noxref_39_c_9876_n ) capacitor c=0.0139868f \
 //x=34.665 //y=2.22 //x2=35.005 //y2=1.59
cc_4807 ( N_SN_c_6855_n N_noxref_39_c_9876_n ) capacitor c=0.00387656f \
 //x=46.135 //y=2.22 //x2=35.005 //y2=1.59
cc_4808 ( N_SN_c_6865_n N_noxref_39_c_9876_n ) capacitor c=0.00251375f \
 //x=34.895 //y=2.22 //x2=35.005 //y2=1.59
cc_4809 ( N_SN_c_6890_n N_noxref_39_c_9876_n ) capacitor c=0.011736f //x=34.78 \
 //y=2.08 //x2=35.005 //y2=1.59
cc_4810 ( N_SN_c_7073_n N_noxref_39_c_9876_n ) capacitor c=0.0157358f \
 //x=34.345 //y=1.22 //x2=35.005 //y2=1.59
cc_4811 ( N_SN_c_7078_n N_noxref_39_c_9876_n ) capacitor c=0.0213278f \
 //x=34.87 //y=1.915 //x2=35.005 //y2=1.59
cc_4812 ( N_SN_c_6844_n N_noxref_39_M20_noxref_s ) capacitor c=0.00642985f \
 //x=34.665 //y=2.22 //x2=33.015 //y2=0.375
cc_4813 ( N_SN_c_6855_n N_noxref_39_M20_noxref_s ) capacitor c=0.00599513f \
 //x=46.135 //y=2.22 //x2=33.015 //y2=0.375
cc_4814 ( N_SN_c_7070_n N_noxref_39_M20_noxref_s ) capacitor c=0.00798959f \
 //x=34.345 //y=0.91 //x2=33.015 //y2=0.375
cc_4815 ( N_SN_c_7077_n N_noxref_39_M20_noxref_s ) capacitor c=0.00212176f \
 //x=34.87 //y=1.45 //x2=33.015 //y2=0.375
cc_4816 ( N_SN_c_7078_n N_noxref_39_M20_noxref_s ) capacitor c=0.00298115f \
 //x=34.87 //y=1.915 //x2=33.015 //y2=0.375
cc_4817 ( N_SN_c_6855_n N_noxref_40_c_9896_n ) capacitor c=0.00657782f \
 //x=46.135 //y=2.22 //x2=35.575 //y2=0.995
cc_4818 ( N_SN_c_7518_p N_noxref_40_c_9896_n ) capacitor c=2.14837e-19 \
 //x=34.715 //y=0.755 //x2=35.575 //y2=0.995
cc_4819 ( N_SN_c_7075_n N_noxref_40_c_9896_n ) capacitor c=0.00123426f \
 //x=34.87 //y=0.91 //x2=35.575 //y2=0.995
cc_4820 ( N_SN_c_7076_n N_noxref_40_c_9896_n ) capacitor c=0.0129288f \
 //x=34.87 //y=1.22 //x2=35.575 //y2=0.995
cc_4821 ( N_SN_c_7077_n N_noxref_40_c_9896_n ) capacitor c=0.00142359f \
 //x=34.87 //y=1.45 //x2=35.575 //y2=0.995
cc_4822 ( N_SN_c_6855_n N_noxref_40_c_9901_n ) capacitor c=0.00147946f \
 //x=46.135 //y=2.22 //x2=36.545 //y2=0.54
cc_4823 ( N_SN_c_7070_n N_noxref_40_M21_noxref_d ) capacitor c=0.00223875f \
 //x=34.345 //y=0.91 //x2=34.42 //y2=0.91
cc_4824 ( N_SN_c_7073_n N_noxref_40_M21_noxref_d ) capacitor c=0.00262485f \
 //x=34.345 //y=1.22 //x2=34.42 //y2=0.91
cc_4825 ( N_SN_c_7518_p N_noxref_40_M21_noxref_d ) capacitor c=0.00220746f \
 //x=34.715 //y=0.755 //x2=34.42 //y2=0.91
cc_4826 ( N_SN_c_7526_p N_noxref_40_M21_noxref_d ) capacitor c=0.00194798f \
 //x=34.715 //y=1.375 //x2=34.42 //y2=0.91
cc_4827 ( N_SN_c_7075_n N_noxref_40_M21_noxref_d ) capacitor c=0.00198465f \
 //x=34.87 //y=0.91 //x2=34.42 //y2=0.91
cc_4828 ( N_SN_c_7076_n N_noxref_40_M21_noxref_d ) capacitor c=0.00128384f \
 //x=34.87 //y=1.22 //x2=34.42 //y2=0.91
cc_4829 ( N_SN_c_6855_n N_noxref_40_M22_noxref_s ) capacitor c=0.00642985f \
 //x=46.135 //y=2.22 //x2=35.525 //y2=0.375
cc_4830 ( N_SN_c_7075_n N_noxref_40_M22_noxref_s ) capacitor c=7.21316e-19 \
 //x=34.87 //y=0.91 //x2=35.525 //y2=0.375
cc_4831 ( N_SN_c_7076_n N_noxref_40_M22_noxref_s ) capacitor c=0.00348171f \
 //x=34.87 //y=1.22 //x2=35.525 //y2=0.375
cc_4832 ( N_SN_c_6855_n N_noxref_41_c_9966_n ) capacitor c=0.00635755f \
 //x=46.135 //y=2.22 //x2=38.065 //y2=1.495
cc_4833 ( N_SN_c_6855_n N_noxref_41_c_9948_n ) capacitor c=0.0223494f \
 //x=46.135 //y=2.22 //x2=38.95 //y2=1.58
cc_4834 ( N_SN_c_6855_n N_noxref_41_c_9955_n ) capacitor c=0.00649228f \
 //x=46.135 //y=2.22 //x2=39.035 //y2=1.495
cc_4835 ( N_SN_c_6855_n N_noxref_41_c_9956_n ) capacitor c=0.00178534f \
 //x=46.135 //y=2.22 //x2=39.92 //y2=0.53
cc_4836 ( N_SN_c_6855_n N_noxref_41_M23_noxref_s ) capacitor c=0.00113237f \
 //x=46.135 //y=2.22 //x2=37.93 //y2=0.365
cc_4837 ( N_SN_c_6855_n N_noxref_42_c_10017_n ) capacitor c=0.00635755f \
 //x=46.135 //y=2.22 //x2=41.395 //y2=1.495
cc_4838 ( N_SN_c_6855_n N_noxref_42_c_9999_n ) capacitor c=0.0223494f \
 //x=46.135 //y=2.22 //x2=42.28 //y2=1.58
cc_4839 ( N_SN_c_6855_n N_noxref_42_c_10006_n ) capacitor c=0.00649228f \
 //x=46.135 //y=2.22 //x2=42.365 //y2=1.495
cc_4840 ( N_SN_c_6855_n N_noxref_42_c_10007_n ) capacitor c=0.00178534f \
 //x=46.135 //y=2.22 //x2=43.25 //y2=0.53
cc_4841 ( N_SN_c_6855_n N_noxref_42_M25_noxref_s ) capacitor c=0.00113237f \
 //x=46.135 //y=2.22 //x2=41.26 //y2=0.365
cc_4842 ( N_SN_c_6855_n N_noxref_43_c_10065_n ) capacitor c=0.00642985f \
 //x=46.135 //y=2.22 //x2=44.62 //y2=1.505
cc_4843 ( N_SN_c_6855_n N_noxref_43_c_10050_n ) capacitor c=0.0225733f \
 //x=46.135 //y=2.22 //x2=45.505 //y2=1.59
cc_4844 ( N_SN_c_7123_n N_noxref_43_c_10057_n ) capacitor c=0.0167228f \
 //x=45.815 //y=0.91 //x2=46.475 //y2=0.54
cc_4845 ( N_SN_c_7128_n N_noxref_43_c_10057_n ) capacitor c=0.00534519f \
 //x=46.34 //y=0.91 //x2=46.475 //y2=0.54
cc_4846 ( N_SN_c_6855_n N_noxref_43_c_10082_n ) capacitor c=0.0139868f \
 //x=46.135 //y=2.22 //x2=46.475 //y2=1.59
cc_4847 ( N_SN_c_6866_n N_noxref_43_c_10082_n ) capacitor c=0.00387656f \
 //x=59.085 //y=2.22 //x2=46.475 //y2=1.59
cc_4848 ( N_SN_c_6876_n N_noxref_43_c_10082_n ) capacitor c=0.00251375f \
 //x=46.365 //y=2.22 //x2=46.475 //y2=1.59
cc_4849 ( N_SN_c_6891_n N_noxref_43_c_10082_n ) capacitor c=0.011736f \
 //x=46.25 //y=2.08 //x2=46.475 //y2=1.59
cc_4850 ( N_SN_c_7126_n N_noxref_43_c_10082_n ) capacitor c=0.0157358f \
 //x=45.815 //y=1.22 //x2=46.475 //y2=1.59
cc_4851 ( N_SN_c_7131_n N_noxref_43_c_10082_n ) capacitor c=0.0213278f \
 //x=46.34 //y=1.915 //x2=46.475 //y2=1.59
cc_4852 ( N_SN_c_6855_n N_noxref_43_M27_noxref_s ) capacitor c=0.00642985f \
 //x=46.135 //y=2.22 //x2=44.485 //y2=0.375
cc_4853 ( N_SN_c_6866_n N_noxref_43_M27_noxref_s ) capacitor c=0.00599513f \
 //x=59.085 //y=2.22 //x2=44.485 //y2=0.375
cc_4854 ( N_SN_c_7123_n N_noxref_43_M27_noxref_s ) capacitor c=0.00798959f \
 //x=45.815 //y=0.91 //x2=44.485 //y2=0.375
cc_4855 ( N_SN_c_7130_n N_noxref_43_M27_noxref_s ) capacitor c=0.00212176f \
 //x=46.34 //y=1.45 //x2=44.485 //y2=0.375
cc_4856 ( N_SN_c_7131_n N_noxref_43_M27_noxref_s ) capacitor c=0.00298115f \
 //x=46.34 //y=1.915 //x2=44.485 //y2=0.375
cc_4857 ( N_SN_c_6866_n N_noxref_44_c_10102_n ) capacitor c=0.00657782f \
 //x=59.085 //y=2.22 //x2=47.045 //y2=0.995
cc_4858 ( N_SN_c_7558_p N_noxref_44_c_10102_n ) capacitor c=2.14837e-19 \
 //x=46.185 //y=0.755 //x2=47.045 //y2=0.995
cc_4859 ( N_SN_c_7128_n N_noxref_44_c_10102_n ) capacitor c=0.00123426f \
 //x=46.34 //y=0.91 //x2=47.045 //y2=0.995
cc_4860 ( N_SN_c_7129_n N_noxref_44_c_10102_n ) capacitor c=0.0129288f \
 //x=46.34 //y=1.22 //x2=47.045 //y2=0.995
cc_4861 ( N_SN_c_7130_n N_noxref_44_c_10102_n ) capacitor c=0.00142359f \
 //x=46.34 //y=1.45 //x2=47.045 //y2=0.995
cc_4862 ( N_SN_c_6866_n N_noxref_44_c_10107_n ) capacitor c=0.00147946f \
 //x=59.085 //y=2.22 //x2=48.015 //y2=0.54
cc_4863 ( N_SN_c_7123_n N_noxref_44_M28_noxref_d ) capacitor c=0.00223875f \
 //x=45.815 //y=0.91 //x2=45.89 //y2=0.91
cc_4864 ( N_SN_c_7126_n N_noxref_44_M28_noxref_d ) capacitor c=0.00262485f \
 //x=45.815 //y=1.22 //x2=45.89 //y2=0.91
cc_4865 ( N_SN_c_7558_p N_noxref_44_M28_noxref_d ) capacitor c=0.00220746f \
 //x=46.185 //y=0.755 //x2=45.89 //y2=0.91
cc_4866 ( N_SN_c_7566_p N_noxref_44_M28_noxref_d ) capacitor c=0.00194798f \
 //x=46.185 //y=1.375 //x2=45.89 //y2=0.91
cc_4867 ( N_SN_c_7128_n N_noxref_44_M28_noxref_d ) capacitor c=0.00198465f \
 //x=46.34 //y=0.91 //x2=45.89 //y2=0.91
cc_4868 ( N_SN_c_7129_n N_noxref_44_M28_noxref_d ) capacitor c=0.00128384f \
 //x=46.34 //y=1.22 //x2=45.89 //y2=0.91
cc_4869 ( N_SN_c_6866_n N_noxref_44_M29_noxref_s ) capacitor c=0.00642985f \
 //x=59.085 //y=2.22 //x2=46.995 //y2=0.375
cc_4870 ( N_SN_c_7128_n N_noxref_44_M29_noxref_s ) capacitor c=7.21316e-19 \
 //x=46.34 //y=0.91 //x2=46.995 //y2=0.375
cc_4871 ( N_SN_c_7129_n N_noxref_44_M29_noxref_s ) capacitor c=0.00348171f \
 //x=46.34 //y=1.22 //x2=46.995 //y2=0.375
cc_4872 ( N_SN_c_6866_n N_noxref_45_c_10172_n ) capacitor c=0.00635755f \
 //x=59.085 //y=2.22 //x2=49.535 //y2=1.495
cc_4873 ( N_SN_c_6866_n N_noxref_45_c_10154_n ) capacitor c=0.0223494f \
 //x=59.085 //y=2.22 //x2=50.42 //y2=1.58
cc_4874 ( N_SN_c_6866_n N_noxref_45_c_10161_n ) capacitor c=0.00649228f \
 //x=59.085 //y=2.22 //x2=50.505 //y2=1.495
cc_4875 ( N_SN_c_6866_n N_noxref_45_c_10162_n ) capacitor c=0.00178534f \
 //x=59.085 //y=2.22 //x2=51.39 //y2=0.53
cc_4876 ( N_SN_c_6866_n N_noxref_45_M30_noxref_s ) capacitor c=0.00113237f \
 //x=59.085 //y=2.22 //x2=49.4 //y2=0.365
cc_4877 ( N_SN_c_6866_n N_noxref_46_c_10220_n ) capacitor c=0.00642985f \
 //x=59.085 //y=2.22 //x2=52.76 //y2=1.505
cc_4878 ( N_SN_c_6866_n N_noxref_46_c_10205_n ) capacitor c=0.0225733f \
 //x=59.085 //y=2.22 //x2=53.645 //y2=1.59
cc_4879 ( N_SN_c_6866_n N_noxref_46_c_10234_n ) capacitor c=0.0203655f \
 //x=59.085 //y=2.22 //x2=54.615 //y2=1.59
cc_4880 ( N_SN_c_6866_n N_noxref_46_M32_noxref_s ) capacitor c=0.012425f \
 //x=59.085 //y=2.22 //x2=52.625 //y2=0.375
cc_4881 ( N_SN_c_6866_n N_noxref_47_c_10254_n ) capacitor c=0.00657782f \
 //x=59.085 //y=2.22 //x2=55.185 //y2=0.995
cc_4882 ( N_SN_c_6866_n N_noxref_47_c_10259_n ) capacitor c=0.00147946f \
 //x=59.085 //y=2.22 //x2=56.155 //y2=0.54
cc_4883 ( N_SN_c_6866_n N_noxref_47_M34_noxref_s ) capacitor c=0.00642985f \
 //x=59.085 //y=2.22 //x2=55.135 //y2=0.375
cc_4884 ( N_SN_c_6866_n N_noxref_48_c_10321_n ) capacitor c=0.00642985f \
 //x=59.085 //y=2.22 //x2=57.57 //y2=1.505
cc_4885 ( N_SN_c_6866_n N_noxref_48_c_10306_n ) capacitor c=0.0225733f \
 //x=59.085 //y=2.22 //x2=58.455 //y2=1.59
cc_4886 ( N_SN_c_7244_n N_noxref_48_c_10313_n ) capacitor c=0.0167228f \
 //x=58.765 //y=0.91 //x2=59.425 //y2=0.54
cc_4887 ( N_SN_c_7249_n N_noxref_48_c_10313_n ) capacitor c=0.00534519f \
 //x=59.29 //y=0.91 //x2=59.425 //y2=0.54
cc_4888 ( N_SN_c_6866_n N_noxref_48_c_10338_n ) capacitor c=0.0139868f \
 //x=59.085 //y=2.22 //x2=59.425 //y2=1.59
cc_4889 ( N_SN_c_6877_n N_noxref_48_c_10338_n ) capacitor c=0.00387656f \
 //x=70.555 //y=2.22 //x2=59.425 //y2=1.59
cc_4890 ( N_SN_c_6887_n N_noxref_48_c_10338_n ) capacitor c=0.00251375f \
 //x=59.315 //y=2.22 //x2=59.425 //y2=1.59
cc_4891 ( N_SN_c_6892_n N_noxref_48_c_10338_n ) capacitor c=0.011736f //x=59.2 \
 //y=2.08 //x2=59.425 //y2=1.59
cc_4892 ( N_SN_c_7247_n N_noxref_48_c_10338_n ) capacitor c=0.0157358f \
 //x=58.765 //y=1.22 //x2=59.425 //y2=1.59
cc_4893 ( N_SN_c_7252_n N_noxref_48_c_10338_n ) capacitor c=0.0213278f \
 //x=59.29 //y=1.915 //x2=59.425 //y2=1.59
cc_4894 ( N_SN_c_6866_n N_noxref_48_M35_noxref_s ) capacitor c=0.00642985f \
 //x=59.085 //y=2.22 //x2=57.435 //y2=0.375
cc_4895 ( N_SN_c_6877_n N_noxref_48_M35_noxref_s ) capacitor c=0.00599513f \
 //x=70.555 //y=2.22 //x2=57.435 //y2=0.375
cc_4896 ( N_SN_c_7244_n N_noxref_48_M35_noxref_s ) capacitor c=0.00798959f \
 //x=58.765 //y=0.91 //x2=57.435 //y2=0.375
cc_4897 ( N_SN_c_7251_n N_noxref_48_M35_noxref_s ) capacitor c=0.00212176f \
 //x=59.29 //y=1.45 //x2=57.435 //y2=0.375
cc_4898 ( N_SN_c_7252_n N_noxref_48_M35_noxref_s ) capacitor c=0.00298115f \
 //x=59.29 //y=1.915 //x2=57.435 //y2=0.375
cc_4899 ( N_SN_c_6877_n N_noxref_49_c_10358_n ) capacitor c=0.00657782f \
 //x=70.555 //y=2.22 //x2=59.995 //y2=0.995
cc_4900 ( N_SN_c_7600_p N_noxref_49_c_10358_n ) capacitor c=2.14837e-19 \
 //x=59.135 //y=0.755 //x2=59.995 //y2=0.995
cc_4901 ( N_SN_c_7249_n N_noxref_49_c_10358_n ) capacitor c=0.00123426f \
 //x=59.29 //y=0.91 //x2=59.995 //y2=0.995
cc_4902 ( N_SN_c_7250_n N_noxref_49_c_10358_n ) capacitor c=0.0129288f \
 //x=59.29 //y=1.22 //x2=59.995 //y2=0.995
cc_4903 ( N_SN_c_7251_n N_noxref_49_c_10358_n ) capacitor c=0.00142359f \
 //x=59.29 //y=1.45 //x2=59.995 //y2=0.995
cc_4904 ( N_SN_c_6877_n N_noxref_49_c_10363_n ) capacitor c=0.00147946f \
 //x=70.555 //y=2.22 //x2=60.965 //y2=0.54
cc_4905 ( N_SN_c_7244_n N_noxref_49_M36_noxref_d ) capacitor c=0.00223875f \
 //x=58.765 //y=0.91 //x2=58.84 //y2=0.91
cc_4906 ( N_SN_c_7247_n N_noxref_49_M36_noxref_d ) capacitor c=0.00262485f \
 //x=58.765 //y=1.22 //x2=58.84 //y2=0.91
cc_4907 ( N_SN_c_7600_p N_noxref_49_M36_noxref_d ) capacitor c=0.00220746f \
 //x=59.135 //y=0.755 //x2=58.84 //y2=0.91
cc_4908 ( N_SN_c_7608_p N_noxref_49_M36_noxref_d ) capacitor c=0.00194798f \
 //x=59.135 //y=1.375 //x2=58.84 //y2=0.91
cc_4909 ( N_SN_c_7249_n N_noxref_49_M36_noxref_d ) capacitor c=0.00198465f \
 //x=59.29 //y=0.91 //x2=58.84 //y2=0.91
cc_4910 ( N_SN_c_7250_n N_noxref_49_M36_noxref_d ) capacitor c=0.00128384f \
 //x=59.29 //y=1.22 //x2=58.84 //y2=0.91
cc_4911 ( N_SN_c_6877_n N_noxref_49_M37_noxref_s ) capacitor c=0.00642985f \
 //x=70.555 //y=2.22 //x2=59.945 //y2=0.375
cc_4912 ( N_SN_c_7249_n N_noxref_49_M37_noxref_s ) capacitor c=7.21316e-19 \
 //x=59.29 //y=0.91 //x2=59.945 //y2=0.375
cc_4913 ( N_SN_c_7250_n N_noxref_49_M37_noxref_s ) capacitor c=0.00348171f \
 //x=59.29 //y=1.22 //x2=59.945 //y2=0.375
cc_4914 ( N_SN_c_6877_n N_noxref_50_c_10428_n ) capacitor c=0.00635755f \
 //x=70.555 //y=2.22 //x2=62.485 //y2=1.495
cc_4915 ( N_SN_c_6877_n N_noxref_50_c_10410_n ) capacitor c=0.0223494f \
 //x=70.555 //y=2.22 //x2=63.37 //y2=1.58
cc_4916 ( N_SN_c_6877_n N_noxref_50_c_10417_n ) capacitor c=0.00649228f \
 //x=70.555 //y=2.22 //x2=63.455 //y2=1.495
cc_4917 ( N_SN_c_6877_n N_noxref_50_c_10418_n ) capacitor c=0.00178534f \
 //x=70.555 //y=2.22 //x2=64.34 //y2=0.53
cc_4918 ( N_SN_c_6877_n N_noxref_50_M38_noxref_s ) capacitor c=0.00113237f \
 //x=70.555 //y=2.22 //x2=62.35 //y2=0.365
cc_4919 ( N_SN_c_6877_n N_noxref_51_c_10479_n ) capacitor c=0.00635755f \
 //x=70.555 //y=2.22 //x2=65.815 //y2=1.495
cc_4920 ( N_SN_c_6877_n N_noxref_51_c_10461_n ) capacitor c=0.0223494f \
 //x=70.555 //y=2.22 //x2=66.7 //y2=1.58
cc_4921 ( N_SN_c_6877_n N_noxref_51_c_10468_n ) capacitor c=0.00649228f \
 //x=70.555 //y=2.22 //x2=66.785 //y2=1.495
cc_4922 ( N_SN_c_6877_n N_noxref_51_c_10469_n ) capacitor c=0.00178534f \
 //x=70.555 //y=2.22 //x2=67.67 //y2=0.53
cc_4923 ( N_SN_c_6877_n N_noxref_51_M40_noxref_s ) capacitor c=0.00113237f \
 //x=70.555 //y=2.22 //x2=65.68 //y2=0.365
cc_4924 ( N_SN_c_6877_n N_noxref_52_c_10529_n ) capacitor c=0.00642985f \
 //x=70.555 //y=2.22 //x2=69.04 //y2=1.505
cc_4925 ( N_SN_c_6877_n N_noxref_52_c_10512_n ) capacitor c=0.0225733f \
 //x=70.555 //y=2.22 //x2=69.925 //y2=1.59
cc_4926 ( N_SN_c_7321_n N_noxref_52_c_10519_n ) capacitor c=0.0167228f \
 //x=70.235 //y=0.91 //x2=70.895 //y2=0.54
cc_4927 ( N_SN_c_7326_n N_noxref_52_c_10519_n ) capacitor c=0.00534519f \
 //x=70.76 //y=0.91 //x2=70.895 //y2=0.54
cc_4928 ( N_SN_c_6877_n N_noxref_52_c_10527_n ) capacitor c=0.0178105f \
 //x=70.555 //y=2.22 //x2=70.895 //y2=1.59
cc_4929 ( N_SN_c_6893_n N_noxref_52_c_10527_n ) capacitor c=0.011736f \
 //x=70.67 //y=2.08 //x2=70.895 //y2=1.59
cc_4930 ( N_SN_c_7324_n N_noxref_52_c_10527_n ) capacitor c=0.0157358f \
 //x=70.235 //y=1.22 //x2=70.895 //y2=1.59
cc_4931 ( N_SN_c_7204_n N_noxref_52_c_10527_n ) capacitor c=0.0215856f \
 //x=70.76 //y=1.915 //x2=70.895 //y2=1.59
cc_4932 ( N_SN_c_6877_n N_noxref_52_M42_noxref_s ) capacitor c=0.00642985f \
 //x=70.555 //y=2.22 //x2=68.905 //y2=0.375
cc_4933 ( N_SN_c_7321_n N_noxref_52_M42_noxref_s ) capacitor c=0.00798959f \
 //x=70.235 //y=0.91 //x2=68.905 //y2=0.375
cc_4934 ( N_SN_c_7328_n N_noxref_52_M42_noxref_s ) capacitor c=0.00212176f \
 //x=70.76 //y=1.45 //x2=68.905 //y2=0.375
cc_4935 ( N_SN_c_7204_n N_noxref_52_M42_noxref_s ) capacitor c=0.00298115f \
 //x=70.76 //y=1.915 //x2=68.905 //y2=0.375
cc_4936 ( N_SN_c_7636_p N_noxref_53_c_10563_n ) capacitor c=2.14837e-19 \
 //x=70.605 //y=0.755 //x2=71.465 //y2=0.995
cc_4937 ( N_SN_c_7326_n N_noxref_53_c_10563_n ) capacitor c=0.00123426f \
 //x=70.76 //y=0.91 //x2=71.465 //y2=0.995
cc_4938 ( N_SN_c_7327_n N_noxref_53_c_10563_n ) capacitor c=0.0129288f \
 //x=70.76 //y=1.22 //x2=71.465 //y2=0.995
cc_4939 ( N_SN_c_7328_n N_noxref_53_c_10563_n ) capacitor c=0.00142359f \
 //x=70.76 //y=1.45 //x2=71.465 //y2=0.995
cc_4940 ( N_SN_c_7321_n N_noxref_53_M43_noxref_d ) capacitor c=0.00223875f \
 //x=70.235 //y=0.91 //x2=70.31 //y2=0.91
cc_4941 ( N_SN_c_7324_n N_noxref_53_M43_noxref_d ) capacitor c=0.00262485f \
 //x=70.235 //y=1.22 //x2=70.31 //y2=0.91
cc_4942 ( N_SN_c_7636_p N_noxref_53_M43_noxref_d ) capacitor c=0.00220746f \
 //x=70.605 //y=0.755 //x2=70.31 //y2=0.91
cc_4943 ( N_SN_c_7643_p N_noxref_53_M43_noxref_d ) capacitor c=0.00194798f \
 //x=70.605 //y=1.375 //x2=70.31 //y2=0.91
cc_4944 ( N_SN_c_7326_n N_noxref_53_M43_noxref_d ) capacitor c=0.00198465f \
 //x=70.76 //y=0.91 //x2=70.31 //y2=0.91
cc_4945 ( N_SN_c_7327_n N_noxref_53_M43_noxref_d ) capacitor c=0.00128384f \
 //x=70.76 //y=1.22 //x2=70.31 //y2=0.91
cc_4946 ( N_SN_c_7326_n N_noxref_53_M44_noxref_s ) capacitor c=7.21316e-19 \
 //x=70.76 //y=0.91 //x2=71.415 //y2=0.375
cc_4947 ( N_SN_c_7327_n N_noxref_53_M44_noxref_s ) capacitor c=0.00348171f \
 //x=70.76 //y=1.22 //x2=71.415 //y2=0.375
cc_4948 ( N_noxref_21_c_7656_n N_noxref_23_c_8089_n ) capacitor c=0.208429f \
 //x=71.665 //y=3.7 //x2=72.405 //y2=4.44
cc_4949 ( N_noxref_21_c_7652_n N_noxref_23_c_8089_n ) capacitor c=0.0226638f \
 //x=71.78 //y=2.08 //x2=72.405 //y2=4.44
cc_4950 ( N_noxref_21_c_7891_n N_noxref_23_c_8089_n ) capacitor c=0.0104371f \
 //x=71.78 //y=4.7 //x2=72.405 //y2=4.44
cc_4951 ( N_noxref_21_c_7656_n N_noxref_23_c_8092_n ) capacitor c=0.0135825f \
 //x=71.665 //y=3.7 //x2=67.085 //y2=4.44
cc_4952 ( N_noxref_21_c_7652_n N_noxref_23_c_8097_n ) capacitor c=0.00136386f \
 //x=71.78 //y=2.08 //x2=72.635 //y2=4.44
cc_4953 ( N_noxref_21_c_7891_n N_noxref_23_c_8097_n ) capacitor c=4.71425e-19 \
 //x=71.78 //y=4.7 //x2=72.635 //y2=4.44
cc_4954 ( N_noxref_21_c_7656_n N_noxref_23_c_8060_n ) capacitor c=0.0195852f \
 //x=71.665 //y=3.7 //x2=66.97 //y2=2.08
cc_4955 ( N_noxref_21_c_7651_n N_noxref_23_c_8060_n ) capacitor c=8.38753e-19 \
 //x=64.38 //y=3.7 //x2=66.97 //y2=2.08
cc_4956 ( N_noxref_21_M140_noxref_g N_noxref_23_c_8117_n ) capacitor \
 c=0.01736f //x=71.52 //y=6.02 //x2=71.655 //y2=5.155
cc_4957 ( N_noxref_21_M141_noxref_g N_noxref_23_c_8121_n ) capacitor \
 c=0.0194981f //x=71.96 //y=6.02 //x2=72.435 //y2=5.155
cc_4958 ( N_noxref_21_c_7891_n N_noxref_23_c_8121_n ) capacitor c=0.00201851f \
 //x=71.78 //y=4.7 //x2=72.435 //y2=5.155
cc_4959 ( N_noxref_21_c_7905_p N_noxref_23_c_8062_n ) capacitor c=0.00359704f \
 //x=72.145 //y=1.415 //x2=72.435 //y2=1.665
cc_4960 ( N_noxref_21_c_7906_p N_noxref_23_c_8062_n ) capacitor c=0.00457401f \
 //x=72.3 //y=1.26 //x2=72.435 //y2=1.665
cc_4961 ( N_noxref_21_c_7656_n N_noxref_23_c_8126_n ) capacitor c=0.00735597f \
 //x=71.665 //y=3.7 //x2=72.52 //y2=4.44
cc_4962 ( N_noxref_21_c_7652_n N_noxref_23_c_8126_n ) capacitor c=0.0826949f \
 //x=71.78 //y=2.08 //x2=72.52 //y2=4.44
cc_4963 ( N_noxref_21_c_7706_n N_noxref_23_c_8126_n ) capacitor c=0.00772308f \
 //x=71.78 //y=2.08 //x2=72.52 //y2=4.44
cc_4964 ( N_noxref_21_c_7890_n N_noxref_23_c_8126_n ) capacitor c=0.00283672f \
 //x=71.78 //y=1.915 //x2=72.52 //y2=4.44
cc_4965 ( N_noxref_21_c_7891_n N_noxref_23_c_8126_n ) capacitor c=0.0121861f \
 //x=71.78 //y=4.7 //x2=72.52 //y2=4.44
cc_4966 ( N_noxref_21_c_7652_n N_noxref_23_c_8063_n ) capacitor c=0.00109179f \
 //x=71.78 //y=2.08 //x2=74 //y2=2.08
cc_4967 ( N_noxref_21_c_7652_n N_noxref_23_c_8312_n ) capacitor c=0.016476f \
 //x=71.78 //y=2.08 //x2=71.74 //y2=5.155
cc_4968 ( N_noxref_21_c_7891_n N_noxref_23_c_8312_n ) capacitor c=0.00475601f \
 //x=71.78 //y=4.7 //x2=71.74 //y2=5.155
cc_4969 ( N_noxref_21_c_7875_n N_noxref_23_M44_noxref_d ) capacitor \
 c=0.00217566f //x=71.77 //y=0.915 //x2=71.845 //y2=0.915
cc_4970 ( N_noxref_21_c_7876_n N_noxref_23_M44_noxref_d ) capacitor \
 c=0.0034598f //x=71.77 //y=1.26 //x2=71.845 //y2=0.915
cc_4971 ( N_noxref_21_c_7877_n N_noxref_23_M44_noxref_d ) capacitor \
 c=0.00544291f //x=71.77 //y=1.57 //x2=71.845 //y2=0.915
cc_4972 ( N_noxref_21_c_7918_p N_noxref_23_M44_noxref_d ) capacitor \
 c=0.00241102f //x=72.145 //y=0.76 //x2=71.845 //y2=0.915
cc_4973 ( N_noxref_21_c_7905_p N_noxref_23_M44_noxref_d ) capacitor \
 c=0.0140297f //x=72.145 //y=1.415 //x2=71.845 //y2=0.915
cc_4974 ( N_noxref_21_c_7920_p N_noxref_23_M44_noxref_d ) capacitor \
 c=0.00219619f //x=72.3 //y=0.915 //x2=71.845 //y2=0.915
cc_4975 ( N_noxref_21_c_7906_p N_noxref_23_M44_noxref_d ) capacitor \
 c=0.00603828f //x=72.3 //y=1.26 //x2=71.845 //y2=0.915
cc_4976 ( N_noxref_21_c_7890_n N_noxref_23_M44_noxref_d ) capacitor \
 c=0.00661782f //x=71.78 //y=1.915 //x2=71.845 //y2=0.915
cc_4977 ( N_noxref_21_M140_noxref_g N_noxref_23_M140_noxref_d ) capacitor \
 c=0.0180032f //x=71.52 //y=6.02 //x2=71.595 //y2=5.02
cc_4978 ( N_noxref_21_M141_noxref_g N_noxref_23_M140_noxref_d ) capacitor \
 c=0.0194246f //x=71.96 //y=6.02 //x2=71.595 //y2=5.02
cc_4979 ( N_noxref_21_c_7696_n N_noxref_24_c_8424_n ) capacitor c=0.404606f \
 //x=60.195 //y=3.7 //x2=79.065 //y2=3.33
cc_4980 ( N_noxref_21_c_7697_n N_noxref_24_c_8424_n ) capacitor c=0.029444f \
 //x=55.615 //y=3.7 //x2=79.065 //y2=3.33
cc_4981 ( N_noxref_21_c_7698_n N_noxref_24_c_8424_n ) capacitor c=0.338821f \
 //x=64.265 //y=3.7 //x2=79.065 //y2=3.33
cc_4982 ( N_noxref_21_c_7699_n N_noxref_24_c_8424_n ) capacitor c=0.026734f \
 //x=60.425 //y=3.7 //x2=79.065 //y2=3.33
cc_4983 ( N_noxref_21_c_7656_n N_noxref_24_c_8424_n ) capacitor c=0.663838f \
 //x=71.665 //y=3.7 //x2=79.065 //y2=3.33
cc_4984 ( N_noxref_21_c_7701_n N_noxref_24_c_8424_n ) capacitor c=0.0266742f \
 //x=64.495 //y=3.7 //x2=79.065 //y2=3.33
cc_4985 ( N_noxref_21_c_7648_n N_noxref_24_c_8424_n ) capacitor c=0.0198536f \
 //x=55.5 //y=2.08 //x2=79.065 //y2=3.33
cc_4986 ( N_noxref_21_c_7649_n N_noxref_24_c_8424_n ) capacitor c=0.0198536f \
 //x=60.31 //y=2.08 //x2=79.065 //y2=3.33
cc_4987 ( N_noxref_21_c_7651_n N_noxref_24_c_8424_n ) capacitor c=0.0205775f \
 //x=64.38 //y=3.7 //x2=79.065 //y2=3.33
cc_4988 ( N_noxref_21_c_7652_n N_noxref_24_c_8424_n ) capacitor c=0.0198536f \
 //x=71.78 //y=2.08 //x2=79.065 //y2=3.33
cc_4989 ( N_noxref_21_c_7648_n N_noxref_47_c_10259_n ) capacitor c=0.00204385f \
 //x=55.5 //y=2.08 //x2=56.155 //y2=0.54
cc_4990 ( N_noxref_21_c_7778_n N_noxref_47_c_10259_n ) capacitor c=0.0194423f \
 //x=55.49 //y=0.915 //x2=56.155 //y2=0.54
cc_4991 ( N_noxref_21_c_7833_n N_noxref_47_c_10259_n ) capacitor c=0.00656458f \
 //x=56.02 //y=0.915 //x2=56.155 //y2=0.54
cc_4992 ( N_noxref_21_c_7781_n N_noxref_47_c_10259_n ) capacitor c=2.20712e-19 \
 //x=55.5 //y=2.08 //x2=56.155 //y2=0.54
cc_4993 ( N_noxref_21_c_7779_n N_noxref_47_c_10281_n ) capacitor c=0.00538033f \
 //x=55.49 //y=1.26 //x2=55.27 //y2=0.995
cc_4994 ( N_noxref_21_c_7778_n N_noxref_47_M34_noxref_s ) capacitor \
 c=0.00538033f //x=55.49 //y=0.915 //x2=55.135 //y2=0.375
cc_4995 ( N_noxref_21_c_7780_n N_noxref_47_M34_noxref_s ) capacitor \
 c=0.00538033f //x=55.49 //y=1.57 //x2=55.135 //y2=0.375
cc_4996 ( N_noxref_21_c_7833_n N_noxref_47_M34_noxref_s ) capacitor \
 c=0.0143002f //x=56.02 //y=0.915 //x2=55.135 //y2=0.375
cc_4997 ( N_noxref_21_c_7834_n N_noxref_47_M34_noxref_s ) capacitor \
 c=0.00290153f //x=56.02 //y=1.26 //x2=55.135 //y2=0.375
cc_4998 ( N_noxref_21_c_7649_n N_noxref_49_c_10363_n ) capacitor c=0.00204385f \
 //x=60.31 //y=2.08 //x2=60.965 //y2=0.54
cc_4999 ( N_noxref_21_c_7729_n N_noxref_49_c_10363_n ) capacitor c=0.0194423f \
 //x=60.3 //y=0.915 //x2=60.965 //y2=0.54
cc_5000 ( N_noxref_21_c_7735_n N_noxref_49_c_10363_n ) capacitor c=0.00656458f \
 //x=60.83 //y=0.915 //x2=60.965 //y2=0.54
cc_5001 ( N_noxref_21_c_7738_n N_noxref_49_c_10363_n ) capacitor c=2.20712e-19 \
 //x=60.31 //y=2.08 //x2=60.965 //y2=0.54
cc_5002 ( N_noxref_21_c_7730_n N_noxref_49_c_10373_n ) capacitor c=0.00538829f \
 //x=60.3 //y=1.26 //x2=60.08 //y2=0.995
cc_5003 ( N_noxref_21_c_7729_n N_noxref_49_M37_noxref_s ) capacitor \
 c=0.00538829f //x=60.3 //y=0.915 //x2=59.945 //y2=0.375
cc_5004 ( N_noxref_21_c_7731_n N_noxref_49_M37_noxref_s ) capacitor \
 c=0.00538829f //x=60.3 //y=1.57 //x2=59.945 //y2=0.375
cc_5005 ( N_noxref_21_c_7735_n N_noxref_49_M37_noxref_s ) capacitor \
 c=0.0143002f //x=60.83 //y=0.915 //x2=59.945 //y2=0.375
cc_5006 ( N_noxref_21_c_7736_n N_noxref_49_M37_noxref_s ) capacitor \
 c=0.00290153f //x=60.83 //y=1.26 //x2=59.945 //y2=0.375
cc_5007 ( N_noxref_21_c_7858_n N_noxref_50_c_10428_n ) capacitor c=3.15806e-19 \
 //x=64.025 //y=1.655 //x2=62.485 //y2=1.495
cc_5008 ( N_noxref_21_c_7858_n N_noxref_50_c_10417_n ) capacitor c=0.020324f \
 //x=64.025 //y=1.655 //x2=63.455 //y2=1.495
cc_5009 ( N_noxref_21_c_7650_n N_noxref_50_c_10418_n ) capacitor c=0.00457164f \
 //x=64.295 //y=1.655 //x2=64.34 //y2=0.53
cc_5010 ( N_noxref_21_M39_noxref_d N_noxref_50_c_10418_n ) capacitor \
 c=0.0115831f //x=63.75 //y=0.905 //x2=64.34 //y2=0.53
cc_5011 ( N_noxref_21_c_7650_n N_noxref_50_M38_noxref_s ) capacitor \
 c=0.013435f //x=64.295 //y=1.655 //x2=62.35 //y2=0.365
cc_5012 ( N_noxref_21_M39_noxref_d N_noxref_50_M38_noxref_s ) capacitor \
 c=0.0439476f //x=63.75 //y=0.905 //x2=62.35 //y2=0.365
cc_5013 ( N_noxref_21_c_7650_n N_noxref_51_c_10479_n ) capacitor c=3.22188e-19 \
 //x=64.295 //y=1.655 //x2=65.815 //y2=1.495
cc_5014 ( N_noxref_21_c_7652_n N_noxref_53_c_10568_n ) capacitor c=0.00207733f \
 //x=71.78 //y=2.08 //x2=72.435 //y2=0.54
cc_5015 ( N_noxref_21_c_7875_n N_noxref_53_c_10568_n ) capacitor c=0.0194423f \
 //x=71.77 //y=0.915 //x2=72.435 //y2=0.54
cc_5016 ( N_noxref_21_c_7920_p N_noxref_53_c_10568_n ) capacitor c=0.00656458f \
 //x=72.3 //y=0.915 //x2=72.435 //y2=0.54
cc_5017 ( N_noxref_21_c_7706_n N_noxref_53_c_10568_n ) capacitor c=2.20712e-19 \
 //x=71.78 //y=2.08 //x2=72.435 //y2=0.54
cc_5018 ( N_noxref_21_c_7876_n N_noxref_53_c_10595_n ) capacitor c=0.00538829f \
 //x=71.77 //y=1.26 //x2=71.55 //y2=0.995
cc_5019 ( N_noxref_21_c_7875_n N_noxref_53_M44_noxref_s ) capacitor \
 c=0.00538829f //x=71.77 //y=0.915 //x2=71.415 //y2=0.375
cc_5020 ( N_noxref_21_c_7877_n N_noxref_53_M44_noxref_s ) capacitor \
 c=0.00538829f //x=71.77 //y=1.57 //x2=71.415 //y2=0.375
cc_5021 ( N_noxref_21_c_7920_p N_noxref_53_M44_noxref_s ) capacitor \
 c=0.0143002f //x=72.3 //y=0.915 //x2=71.415 //y2=0.375
cc_5022 ( N_noxref_21_c_7906_p N_noxref_53_M44_noxref_s ) capacitor \
 c=0.00290153f //x=72.3 //y=1.26 //x2=71.415 //y2=0.375
cc_5023 ( N_noxref_22_c_7969_n N_noxref_23_c_8100_n ) capacitor c=0.0856654f \
 //x=77.255 //y=5.21 //x2=77.585 //y2=4.44
cc_5024 ( N_noxref_22_c_7975_n N_noxref_23_c_8100_n ) capacitor c=0.0130311f \
 //x=75.485 //y=5.21 //x2=77.585 //y2=4.44
cc_5025 ( N_noxref_22_c_7980_n N_noxref_23_c_8100_n ) capacitor c=0.00145992f \
 //x=75.285 //y=5.21 //x2=77.585 //y2=4.44
cc_5026 ( N_noxref_22_c_7984_n N_noxref_23_c_8100_n ) capacitor c=0.0197096f \
 //x=74.575 //y=5.21 //x2=77.585 //y2=4.44
cc_5027 ( N_noxref_22_c_7986_n N_noxref_23_c_8100_n ) capacitor c=0.00467548f \
 //x=75.37 //y=5.295 //x2=77.585 //y2=4.44
cc_5028 ( N_noxref_22_c_7989_n N_noxref_23_c_8100_n ) capacitor c=0.00439121f \
 //x=77.37 //y=5.21 //x2=77.585 //y2=4.44
cc_5029 ( N_noxref_22_c_8022_p N_noxref_23_c_8100_n ) capacitor c=0.00249667f \
 //x=78.165 //y=6.91 //x2=77.585 //y2=4.44
cc_5030 ( N_noxref_22_c_8022_p N_noxref_23_c_8066_n ) capacitor c=8.81369e-19 \
 //x=78.165 //y=6.91 //x2=77.7 //y2=2.08
cc_5031 ( N_noxref_22_c_7984_n N_noxref_23_M142_noxref_g ) capacitor \
 c=0.0172236f //x=74.575 //y=5.21 //x2=74.27 //y2=6.025
cc_5032 ( N_noxref_22_c_7980_n N_noxref_23_M143_noxref_g ) capacitor \
 c=0.0169795f //x=75.285 //y=5.21 //x2=74.71 //y2=6.025
cc_5033 ( N_noxref_22_M142_noxref_d N_noxref_23_M143_noxref_g ) capacitor \
 c=0.0169879f //x=74.345 //y=5.025 //x2=74.71 //y2=6.025
cc_5034 ( N_noxref_22_c_7969_n N_noxref_23_M146_noxref_g ) capacitor \
 c=0.00503498f //x=77.255 //y=5.21 //x2=77.59 //y2=6.025
cc_5035 ( N_noxref_22_c_7989_n N_noxref_23_M146_noxref_g ) capacitor \
 c=0.0481665f //x=77.37 //y=5.21 //x2=77.59 //y2=6.025
cc_5036 ( N_noxref_22_c_8022_p N_noxref_23_M146_noxref_g ) capacitor \
 c=0.0163949f //x=78.165 //y=6.91 //x2=77.59 //y2=6.025
cc_5037 ( N_noxref_22_c_8022_p N_noxref_23_M147_noxref_g ) capacitor \
 c=0.0150104f //x=78.165 //y=6.91 //x2=78.03 //y2=6.025
cc_5038 ( N_noxref_22_M147_noxref_d N_noxref_23_M147_noxref_g ) capacitor \
 c=0.0130327f //x=78.105 //y=5.025 //x2=78.03 //y2=6.025
cc_5039 ( N_noxref_22_c_7984_n N_noxref_23_c_8197_n ) capacitor c=0.00405363f \
 //x=74.575 //y=5.21 //x2=74.635 //y2=4.795
cc_5040 ( N_noxref_22_M149_noxref_d N_noxref_24_c_8431_n ) capacitor \
 c=0.00496677f //x=78.985 //y=5.025 //x2=79.18 //y2=2.08
cc_5041 ( N_noxref_22_c_8034_p N_noxref_24_M148_noxref_g ) capacitor \
 c=0.0150104f //x=79.045 //y=6.91 //x2=78.47 //y2=6.025
cc_5042 ( N_noxref_22_M147_noxref_d N_noxref_24_M148_noxref_g ) capacitor \
 c=0.0130327f //x=78.105 //y=5.025 //x2=78.47 //y2=6.025
cc_5043 ( N_noxref_22_c_8034_p N_noxref_24_M149_noxref_g ) capacitor \
 c=0.0155183f //x=79.045 //y=6.91 //x2=78.91 //y2=6.025
cc_5044 ( N_noxref_22_M149_noxref_d N_noxref_24_M149_noxref_g ) capacitor \
 c=0.0398886f //x=78.985 //y=5.025 //x2=78.91 //y2=6.025
cc_5045 ( N_noxref_22_M149_noxref_d N_noxref_24_c_8480_n ) capacitor \
 c=0.00411435f //x=78.985 //y=5.025 //x2=78.91 //y2=4.87
cc_5046 ( N_noxref_22_c_8034_p N_noxref_25_c_8898_n ) capacitor c=0.00546043f \
 //x=79.045 //y=6.91 //x2=80.595 //y2=5.21
cc_5047 ( N_noxref_22_M149_noxref_d N_noxref_25_c_8898_n ) capacitor \
 c=0.00675852f //x=78.985 //y=5.025 //x2=80.595 //y2=5.21
cc_5048 ( N_noxref_22_c_7969_n N_noxref_25_c_8902_n ) capacitor c=0.0086908f \
 //x=77.255 //y=5.21 //x2=78.805 //y2=5.21
cc_5049 ( N_noxref_22_c_8034_p N_noxref_25_c_8902_n ) capacitor c=9.39989e-19 \
 //x=79.045 //y=6.91 //x2=78.805 //y2=5.21
cc_5050 ( N_noxref_22_c_8022_p N_noxref_25_c_8916_n ) capacitor c=0.00102709f \
 //x=78.165 //y=6.91 //x2=78.605 //y2=5.21
cc_5051 ( N_noxref_22_c_8034_p N_noxref_25_c_8916_n ) capacitor c=9.89472e-19 \
 //x=79.045 //y=6.91 //x2=78.605 //y2=5.21
cc_5052 ( N_noxref_22_M147_noxref_d N_noxref_25_c_8916_n ) capacitor \
 c=0.0124612f //x=78.105 //y=5.025 //x2=78.605 //y2=5.21
cc_5053 ( N_noxref_22_c_7969_n N_noxref_25_c_8904_n ) capacitor c=0.00638395f \
 //x=77.255 //y=5.21 //x2=77.895 //y2=5.21
cc_5054 ( N_noxref_22_c_7989_n N_noxref_25_c_8904_n ) capacitor c=0.0682565f \
 //x=77.37 //y=5.21 //x2=77.895 //y2=5.21
cc_5055 ( N_noxref_22_c_7989_n N_noxref_25_c_8905_n ) capacitor c=9.46973e-19 \
 //x=77.37 //y=5.21 //x2=78.69 //y2=5.295
cc_5056 ( N_noxref_22_M149_noxref_d N_noxref_25_c_8906_n ) capacitor \
 c=0.001104f //x=78.985 //y=5.025 //x2=80.71 //y2=5.21
cc_5057 ( N_noxref_22_c_8034_p N_noxref_25_c_8908_n ) capacitor c=0.001104f \
 //x=79.045 //y=6.91 //x2=80.795 //y2=6.91
cc_5058 ( N_noxref_22_c_7969_n N_noxref_25_M146_noxref_d ) capacitor \
 c=4.76678e-19 //x=77.255 //y=5.21 //x2=77.665 //y2=5.025
cc_5059 ( N_noxref_22_c_8022_p N_noxref_25_M146_noxref_d ) capacitor \
 c=0.0115421f //x=78.165 //y=6.91 //x2=77.665 //y2=5.025
cc_5060 ( N_noxref_22_M147_noxref_d N_noxref_25_M146_noxref_d ) capacitor \
 c=0.0458293f //x=78.105 //y=5.025 //x2=77.665 //y2=5.025
cc_5061 ( N_noxref_22_M149_noxref_d N_noxref_25_M146_noxref_d ) capacitor \
 c=7.47391e-19 //x=78.985 //y=5.025 //x2=77.665 //y2=5.025
cc_5062 ( N_noxref_22_c_7989_n N_noxref_25_M148_noxref_d ) capacitor \
 c=9.55e-19 //x=77.37 //y=5.21 //x2=78.545 //y2=5.025
cc_5063 ( N_noxref_22_c_8034_p N_noxref_25_M148_noxref_d ) capacitor \
 c=0.0115693f //x=79.045 //y=6.91 //x2=78.545 //y2=5.025
cc_5064 ( N_noxref_22_M147_noxref_d N_noxref_25_M148_noxref_d ) capacitor \
 c=0.0458293f //x=78.105 //y=5.025 //x2=78.545 //y2=5.025
cc_5065 ( N_noxref_22_M149_noxref_d N_noxref_25_M148_noxref_d ) capacitor \
 c=0.0550393f //x=78.985 //y=5.025 //x2=78.545 //y2=5.025
cc_5066 ( N_noxref_22_c_7989_n N_noxref_55_c_10689_n ) capacitor c=0.00110943f \
 //x=77.37 //y=5.21 //x2=77.285 //y2=1.495
cc_5067 ( N_noxref_23_c_8089_n N_noxref_24_c_8424_n ) capacitor c=0.0386482f \
 //x=72.405 //y=4.44 //x2=79.065 //y2=3.33
cc_5068 ( N_noxref_23_c_8092_n N_noxref_24_c_8424_n ) capacitor c=6.32406e-19 \
 //x=67.085 //y=4.44 //x2=79.065 //y2=3.33
cc_5069 ( N_noxref_23_c_8093_n N_noxref_24_c_8424_n ) capacitor c=0.0379268f \
 //x=73.885 //y=4.44 //x2=79.065 //y2=3.33
cc_5070 ( N_noxref_23_c_8097_n N_noxref_24_c_8424_n ) capacitor c=0.00699571f \
 //x=72.635 //y=4.44 //x2=79.065 //y2=3.33
cc_5071 ( N_noxref_23_c_8100_n N_noxref_24_c_8424_n ) capacitor c=0.0359616f \
 //x=77.585 //y=4.44 //x2=79.065 //y2=3.33
cc_5072 ( N_noxref_23_c_8105_n N_noxref_24_c_8424_n ) capacitor c=0.00681681f \
 //x=74.115 //y=4.44 //x2=79.065 //y2=3.33
cc_5073 ( N_noxref_23_c_8060_n N_noxref_24_c_8424_n ) capacitor c=0.0169786f \
 //x=66.97 //y=2.08 //x2=79.065 //y2=3.33
cc_5074 ( N_noxref_23_c_8126_n N_noxref_24_c_8424_n ) capacitor c=0.0224844f \
 //x=72.52 //y=4.44 //x2=79.065 //y2=3.33
cc_5075 ( N_noxref_23_c_8063_n N_noxref_24_c_8424_n ) capacitor c=0.0235144f \
 //x=74 //y=2.08 //x2=79.065 //y2=3.33
cc_5076 ( N_noxref_23_c_8066_n N_noxref_24_c_8424_n ) capacitor c=0.0282872f \
 //x=77.7 //y=2.08 //x2=79.065 //y2=3.33
cc_5077 ( N_noxref_23_c_8066_n N_noxref_24_c_8427_n ) capacitor c=0.00622935f \
 //x=77.7 //y=2.08 //x2=79.295 //y2=2.08
cc_5078 ( N_noxref_23_c_8100_n N_noxref_24_c_8431_n ) capacitor c=0.00408423f \
 //x=77.585 //y=4.44 //x2=79.18 //y2=2.08
cc_5079 ( N_noxref_23_c_8066_n N_noxref_24_c_8431_n ) capacitor c=0.0343626f \
 //x=77.7 //y=2.08 //x2=79.18 //y2=2.08
cc_5080 ( N_noxref_23_c_8081_n N_noxref_24_c_8431_n ) capacitor c=2.35599e-19 \
 //x=77.505 //y=1.915 //x2=79.18 //y2=2.08
cc_5081 ( N_noxref_23_c_8148_n N_noxref_24_c_8431_n ) capacitor c=2.35599e-19 \
 //x=77.7 //y=4.705 //x2=79.18 //y2=2.08
cc_5082 ( N_noxref_23_c_8066_n N_noxref_24_c_8433_n ) capacitor c=5.76627e-19 \
 //x=77.7 //y=2.08 //x2=80.66 //y2=2.08
cc_5083 ( N_noxref_23_M146_noxref_g N_noxref_24_M148_noxref_g ) capacitor \
 c=0.009459f //x=77.59 //y=6.025 //x2=78.47 //y2=6.025
cc_5084 ( N_noxref_23_M147_noxref_g N_noxref_24_M148_noxref_g ) capacitor \
 c=0.0626756f //x=78.03 //y=6.025 //x2=78.47 //y2=6.025
cc_5085 ( N_noxref_23_M147_noxref_g N_noxref_24_M149_noxref_g ) capacitor \
 c=0.00899012f //x=78.03 //y=6.025 //x2=78.91 //y2=6.025
cc_5086 ( N_noxref_23_c_8078_n N_noxref_24_c_8778_n ) capacitor c=4.86506e-19 \
 //x=77.505 //y=0.865 //x2=78.475 //y2=0.905
cc_5087 ( N_noxref_23_c_8080_n N_noxref_24_c_8778_n ) capacitor c=0.00101233f \
 //x=77.505 //y=1.21 //x2=78.475 //y2=0.905
cc_5088 ( N_noxref_23_c_8084_n N_noxref_24_c_8778_n ) capacitor c=0.0168844f \
 //x=78.035 //y=0.865 //x2=78.475 //y2=0.905
cc_5089 ( N_noxref_23_c_8363_p N_noxref_24_c_8781_n ) capacitor c=7.88071e-19 \
 //x=77.505 //y=1.52 //x2=78.475 //y2=1.25
cc_5090 ( N_noxref_23_c_8086_n N_noxref_24_c_8781_n ) capacitor c=0.0168218f \
 //x=78.035 //y=1.21 //x2=78.475 //y2=1.25
cc_5091 ( N_noxref_23_c_8066_n N_noxref_24_c_8640_n ) capacitor c=9.39431e-19 \
 //x=77.7 //y=2.08 //x2=78.545 //y2=4.795
cc_5092 ( N_noxref_23_c_8148_n N_noxref_24_c_8640_n ) capacitor c=0.0634092f \
 //x=77.7 //y=4.705 //x2=78.545 //y2=4.795
cc_5093 ( N_noxref_23_c_8066_n N_noxref_24_c_8480_n ) capacitor c=2.35599e-19 \
 //x=77.7 //y=2.08 //x2=78.91 //y2=4.87
cc_5094 ( N_noxref_23_c_8148_n N_noxref_24_c_8480_n ) capacitor c=5.35364e-19 \
 //x=77.7 //y=4.705 //x2=78.91 //y2=4.87
cc_5095 ( N_noxref_23_c_8084_n N_noxref_24_c_8787_n ) capacitor c=0.00124821f \
 //x=78.035 //y=0.865 //x2=79.005 //y2=0.905
cc_5096 ( N_noxref_23_c_8086_n N_noxref_24_c_8788_n ) capacitor c=8.19575e-19 \
 //x=78.035 //y=1.21 //x2=79.005 //y2=1.25
cc_5097 ( N_noxref_23_c_8086_n N_noxref_24_c_8789_n ) capacitor c=3.60397e-19 \
 //x=78.035 //y=1.21 //x2=79.005 //y2=1.56
cc_5098 ( N_noxref_23_c_8081_n N_noxref_24_c_8434_n ) capacitor c=4.61972e-19 \
 //x=77.505 //y=1.915 //x2=79.005 //y2=1.915
cc_5099 ( N_noxref_23_M147_noxref_g N_noxref_25_c_8916_n ) capacitor \
 c=0.0179287f //x=78.03 //y=6.025 //x2=78.605 //y2=5.21
cc_5100 ( N_noxref_23_c_8100_n N_noxref_25_c_8904_n ) capacitor c=0.0021588f \
 //x=77.585 //y=4.44 //x2=77.895 //y2=5.21
cc_5101 ( N_noxref_23_c_8066_n N_noxref_25_c_8904_n ) capacitor c=0.0056513f \
 //x=77.7 //y=2.08 //x2=77.895 //y2=5.21
cc_5102 ( N_noxref_23_M146_noxref_g N_noxref_25_c_8904_n ) capacitor \
 c=0.0132827f //x=77.59 //y=6.025 //x2=77.895 //y2=5.21
cc_5103 ( N_noxref_23_c_8148_n N_noxref_25_c_8904_n ) capacitor c=0.00554802f \
 //x=77.7 //y=4.705 //x2=77.895 //y2=5.21
cc_5104 ( N_noxref_23_M147_noxref_g N_noxref_25_M146_noxref_d ) capacitor \
 c=0.0130327f //x=78.03 //y=6.025 //x2=77.665 //y2=5.025
cc_5105 ( N_noxref_23_c_8080_n N_noxref_26_c_8988_n ) capacitor c=0.00500281f \
 //x=77.505 //y=1.21 //x2=78.625 //y2=1.18
cc_5106 ( N_noxref_23_c_8363_p N_noxref_26_c_8988_n ) capacitor c=0.00352558f \
 //x=77.505 //y=1.52 //x2=78.625 //y2=1.18
cc_5107 ( N_noxref_23_c_8082_n N_noxref_26_c_8988_n ) capacitor c=4.02408e-19 \
 //x=77.88 //y=0.71 //x2=78.625 //y2=1.18
cc_5108 ( N_noxref_23_c_8083_n N_noxref_26_c_8988_n ) capacitor c=0.00341863f \
 //x=77.88 //y=1.365 //x2=78.625 //y2=1.18
cc_5109 ( N_noxref_23_c_8086_n N_noxref_26_c_8988_n ) capacitor c=0.00753876f \
 //x=78.035 //y=1.21 //x2=78.625 //y2=1.18
cc_5110 ( N_noxref_23_c_8226_n N_noxref_51_c_10468_n ) capacitor c=0.00623646f \
 //x=67.005 //y=1.56 //x2=66.785 //y2=1.495
cc_5111 ( N_noxref_23_c_8231_n N_noxref_51_c_10468_n ) capacitor c=0.00173579f \
 //x=66.97 //y=2.08 //x2=66.785 //y2=1.495
cc_5112 ( N_noxref_23_c_8060_n N_noxref_51_c_10469_n ) capacitor c=0.00156605f \
 //x=66.97 //y=2.08 //x2=67.67 //y2=0.53
cc_5113 ( N_noxref_23_c_8221_n N_noxref_51_c_10469_n ) capacitor c=0.0188655f \
 //x=67.005 //y=0.905 //x2=67.67 //y2=0.53
cc_5114 ( N_noxref_23_c_8229_n N_noxref_51_c_10469_n ) capacitor c=0.00656458f \
 //x=67.535 //y=0.905 //x2=67.67 //y2=0.53
cc_5115 ( N_noxref_23_c_8231_n N_noxref_51_c_10469_n ) capacitor c=2.1838e-19 \
 //x=66.97 //y=2.08 //x2=67.67 //y2=0.53
cc_5116 ( N_noxref_23_c_8221_n N_noxref_51_M40_noxref_s ) capacitor \
 c=0.00623646f //x=67.005 //y=0.905 //x2=65.68 //y2=0.365
cc_5117 ( N_noxref_23_c_8229_n N_noxref_51_M40_noxref_s ) capacitor \
 c=0.0143002f //x=67.535 //y=0.905 //x2=65.68 //y2=0.365
cc_5118 ( N_noxref_23_c_8230_n N_noxref_51_M40_noxref_s ) capacitor \
 c=0.00290153f //x=67.535 //y=1.25 //x2=65.68 //y2=0.365
cc_5119 ( N_noxref_23_M44_noxref_d N_noxref_52_M42_noxref_s ) capacitor \
 c=0.00309936f //x=71.845 //y=0.915 //x2=68.905 //y2=0.375
cc_5120 ( N_noxref_23_c_8062_n N_noxref_53_c_10568_n ) capacitor c=0.00464291f \
 //x=72.435 //y=1.665 //x2=72.435 //y2=0.54
cc_5121 ( N_noxref_23_M44_noxref_d N_noxref_53_c_10568_n ) capacitor \
 c=0.0117407f //x=71.845 //y=0.915 //x2=72.435 //y2=0.54
cc_5122 ( N_noxref_23_c_8177_n N_noxref_53_c_10595_n ) capacitor c=0.020048f \
 //x=72.12 //y=1.665 //x2=71.55 //y2=0.995
cc_5123 ( N_noxref_23_M44_noxref_d N_noxref_53_M43_noxref_d ) capacitor \
 c=5.27807e-19 //x=71.845 //y=0.915 //x2=70.31 //y2=0.91
cc_5124 ( N_noxref_23_c_8062_n N_noxref_53_M44_noxref_s ) capacitor \
 c=0.0205269f //x=72.435 //y=1.665 //x2=71.415 //y2=0.375
cc_5125 ( N_noxref_23_M44_noxref_d N_noxref_53_M44_noxref_s ) capacitor \
 c=0.0426134f //x=71.845 //y=0.915 //x2=71.415 //y2=0.375
cc_5126 ( N_noxref_23_c_8062_n N_noxref_54_c_10633_n ) capacitor c=3.04182e-19 \
 //x=72.435 //y=1.665 //x2=73.955 //y2=1.495
cc_5127 ( N_noxref_23_c_8063_n N_noxref_54_c_10633_n ) capacitor c=0.0160451f \
 //x=74 //y=2.08 //x2=73.955 //y2=1.495
cc_5128 ( N_noxref_23_c_8072_n N_noxref_54_c_10633_n ) capacitor c=0.0034165f \
 //x=74.175 //y=1.915 //x2=73.955 //y2=1.495
cc_5129 ( N_noxref_23_c_8087_n N_noxref_54_c_10633_n ) capacitor c=0.00781973f \
 //x=74 //y=2.08 //x2=73.955 //y2=1.495
cc_5130 ( N_noxref_23_c_8063_n N_noxref_54_c_10615_n ) capacitor c=0.00513915f \
 //x=74 //y=2.08 //x2=74.84 //y2=1.58
cc_5131 ( N_noxref_23_c_8071_n N_noxref_54_c_10615_n ) capacitor c=0.00720513f \
 //x=74.175 //y=1.52 //x2=74.84 //y2=1.58
cc_5132 ( N_noxref_23_c_8072_n N_noxref_54_c_10615_n ) capacitor c=0.0140339f \
 //x=74.175 //y=1.915 //x2=74.84 //y2=1.58
cc_5133 ( N_noxref_23_c_8074_n N_noxref_54_c_10615_n ) capacitor c=0.0100869f \
 //x=74.55 //y=1.365 //x2=74.84 //y2=1.58
cc_5134 ( N_noxref_23_c_8077_n N_noxref_54_c_10615_n ) capacitor c=0.00339872f \
 //x=74.705 //y=1.21 //x2=74.84 //y2=1.58
cc_5135 ( N_noxref_23_c_8087_n N_noxref_54_c_10615_n ) capacitor c=0.00324565f \
 //x=74 //y=2.08 //x2=74.84 //y2=1.58
cc_5136 ( N_noxref_23_c_8072_n N_noxref_54_c_10622_n ) capacitor c=6.71402e-19 \
 //x=74.175 //y=1.915 //x2=74.925 //y2=1.495
cc_5137 ( N_noxref_23_c_8068_n N_noxref_54_M45_noxref_s ) capacitor \
 c=0.0326926f //x=74.175 //y=0.865 //x2=73.82 //y2=0.365
cc_5138 ( N_noxref_23_c_8071_n N_noxref_54_M45_noxref_s ) capacitor \
 c=0.00110192f //x=74.175 //y=1.52 //x2=73.82 //y2=0.365
cc_5139 ( N_noxref_23_c_8075_n N_noxref_54_M45_noxref_s ) capacitor \
 c=0.0120759f //x=74.705 //y=0.865 //x2=73.82 //y2=0.365
cc_5140 ( N_noxref_23_c_8081_n N_noxref_55_c_10689_n ) capacitor c=0.0034165f \
 //x=77.505 //y=1.915 //x2=77.285 //y2=1.495
cc_5141 ( N_noxref_23_c_8066_n N_noxref_55_c_10672_n ) capacitor c=0.0112688f \
 //x=77.7 //y=2.08 //x2=78.17 //y2=1.58
cc_5142 ( N_noxref_23_c_8363_p N_noxref_55_c_10672_n ) capacitor c=0.00598984f \
 //x=77.505 //y=1.52 //x2=78.17 //y2=1.58
cc_5143 ( N_noxref_23_c_8081_n N_noxref_55_c_10672_n ) capacitor c=0.0203825f \
 //x=77.505 //y=1.915 //x2=78.17 //y2=1.58
cc_5144 ( N_noxref_23_c_8083_n N_noxref_55_c_10672_n ) capacitor c=0.00767729f \
 //x=77.88 //y=1.365 //x2=78.17 //y2=1.58
cc_5145 ( N_noxref_23_c_8086_n N_noxref_55_c_10672_n ) capacitor c=0.0059368f \
 //x=78.035 //y=1.21 //x2=78.17 //y2=1.58
cc_5146 ( N_noxref_23_c_8081_n N_noxref_55_c_10678_n ) capacitor c=0.00122123f \
 //x=77.505 //y=1.915 //x2=78.255 //y2=1.495
cc_5147 ( N_noxref_23_c_8078_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.0312776f //x=77.505 //y=0.865 //x2=77.15 //y2=0.365
cc_5148 ( N_noxref_23_c_8363_p N_noxref_55_M47_noxref_s ) capacitor \
 c=3.48408e-19 //x=77.505 //y=1.52 //x2=77.15 //y2=0.365
cc_5149 ( N_noxref_23_c_8084_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.0132463f //x=78.035 //y=0.865 //x2=77.15 //y2=0.365
cc_5150 ( N_noxref_24_c_8424_n N_noxref_25_c_8898_n ) capacitor c=9.03043e-19 \
 //x=79.065 //y=3.33 //x2=80.595 //y2=5.21
cc_5151 ( N_noxref_24_c_8426_n N_noxref_25_c_8898_n ) capacitor c=5.48246e-19 \
 //x=80.545 //y=2.08 //x2=80.595 //y2=5.21
cc_5152 ( N_noxref_24_c_8431_n N_noxref_25_c_8898_n ) capacitor c=0.00419026f \
 //x=79.18 //y=2.08 //x2=80.595 //y2=5.21
cc_5153 ( N_noxref_24_c_8433_n N_noxref_25_c_8898_n ) capacitor c=0.0031527f \
 //x=80.66 //y=2.08 //x2=80.595 //y2=5.21
cc_5154 ( N_noxref_24_M149_noxref_g N_noxref_25_c_8898_n ) capacitor \
 c=0.0109874f //x=78.91 //y=6.025 //x2=80.595 //y2=5.21
cc_5155 ( N_noxref_24_M150_noxref_g N_noxref_25_c_8898_n ) capacitor \
 c=0.00645933f //x=80.93 //y=6.025 //x2=80.595 //y2=5.21
cc_5156 ( N_noxref_24_c_8480_n N_noxref_25_c_8898_n ) capacitor c=0.00270424f \
 //x=78.91 //y=4.87 //x2=80.595 //y2=5.21
cc_5157 ( N_noxref_24_c_8481_n N_noxref_25_c_8898_n ) capacitor c=0.00176728f \
 //x=81.005 //y=4.795 //x2=80.595 //y2=5.21
cc_5158 ( N_noxref_24_c_8424_n N_noxref_25_c_8902_n ) capacitor c=5.58709e-19 \
 //x=79.065 //y=3.33 //x2=78.805 //y2=5.21
cc_5159 ( N_noxref_24_M148_noxref_g N_noxref_25_c_8902_n ) capacitor \
 c=6.87102e-19 //x=78.47 //y=6.025 //x2=78.805 //y2=5.21
cc_5160 ( N_noxref_24_M149_noxref_g N_noxref_25_c_8902_n ) capacitor \
 c=8.33934e-19 //x=78.91 //y=6.025 //x2=78.805 //y2=5.21
cc_5161 ( N_noxref_24_M148_noxref_g N_noxref_25_c_8916_n ) capacitor \
 c=0.0179287f //x=78.47 //y=6.025 //x2=78.605 //y2=5.21
cc_5162 ( N_noxref_24_M148_noxref_g N_noxref_25_c_8905_n ) capacitor \
 c=0.0019882f //x=78.47 //y=6.025 //x2=78.69 //y2=5.295
cc_5163 ( N_noxref_24_M149_noxref_g N_noxref_25_c_8905_n ) capacitor \
 c=0.0159381f //x=78.91 //y=6.025 //x2=78.69 //y2=5.295
cc_5164 ( N_noxref_24_c_8805_p N_noxref_25_c_8905_n ) capacitor c=0.00456817f \
 //x=78.835 //y=4.795 //x2=78.69 //y2=5.295
cc_5165 ( N_noxref_24_c_8433_n N_noxref_25_c_8906_n ) capacitor c=0.0183146f \
 //x=80.66 //y=2.08 //x2=80.71 //y2=5.21
cc_5166 ( N_noxref_24_M150_noxref_g N_noxref_25_c_8906_n ) capacitor \
 c=0.0484795f //x=80.93 //y=6.025 //x2=80.71 //y2=5.21
cc_5167 ( N_noxref_24_c_8481_n N_noxref_25_c_8906_n ) capacitor c=0.0078825f \
 //x=81.005 //y=4.795 //x2=80.71 //y2=5.21
cc_5168 ( N_noxref_24_M150_noxref_g N_noxref_25_c_8920_n ) capacitor \
 c=0.0164606f //x=80.93 //y=6.025 //x2=81.505 //y2=6.91
cc_5169 ( N_noxref_24_M151_noxref_g N_noxref_25_c_8920_n ) capacitor \
 c=0.0150104f //x=81.37 //y=6.025 //x2=81.505 //y2=6.91
cc_5170 ( N_noxref_24_M148_noxref_g N_noxref_25_M148_noxref_d ) capacitor \
 c=0.0129738f //x=78.47 //y=6.025 //x2=78.545 //y2=5.025
cc_5171 ( N_noxref_24_M151_noxref_g N_noxref_25_M151_noxref_d ) capacitor \
 c=0.0130327f //x=81.37 //y=6.025 //x2=81.445 //y2=5.025
cc_5172 ( N_noxref_24_c_8424_n N_noxref_26_c_8988_n ) capacitor c=0.0396175f \
 //x=79.065 //y=3.33 //x2=78.625 //y2=1.18
cc_5173 ( N_noxref_24_c_8778_n N_noxref_26_c_8988_n ) capacitor c=5.17481e-19 \
 //x=78.475 //y=0.905 //x2=78.625 //y2=1.18
cc_5174 ( N_noxref_24_c_8781_n N_noxref_26_c_8988_n ) capacitor c=0.00624467f \
 //x=78.475 //y=1.25 //x2=78.625 //y2=1.18
cc_5175 ( N_noxref_24_c_8424_n N_noxref_26_c_8995_n ) capacitor c=0.00382246f \
 //x=79.065 //y=3.33 //x2=75.525 //y2=1.18
cc_5176 ( N_noxref_24_c_8424_n N_noxref_26_c_8996_n ) capacitor c=0.00273991f \
 //x=79.065 //y=3.33 //x2=81.955 //y2=1.18
cc_5177 ( N_noxref_24_c_8426_n N_noxref_26_c_8996_n ) capacitor c=0.053129f \
 //x=80.545 //y=2.08 //x2=81.955 //y2=1.18
cc_5178 ( N_noxref_24_c_8427_n N_noxref_26_c_8996_n ) capacitor c=0.0102038f \
 //x=79.295 //y=2.08 //x2=81.955 //y2=1.18
cc_5179 ( N_noxref_24_c_8431_n N_noxref_26_c_8996_n ) capacitor c=0.00189559f \
 //x=79.18 //y=2.08 //x2=81.955 //y2=1.18
cc_5180 ( N_noxref_24_c_8433_n N_noxref_26_c_8996_n ) capacitor c=0.00134607f \
 //x=80.66 //y=2.08 //x2=81.955 //y2=1.18
cc_5181 ( N_noxref_24_c_8787_n N_noxref_26_c_8996_n ) capacitor c=4.67724e-19 \
 //x=79.005 //y=0.905 //x2=81.955 //y2=1.18
cc_5182 ( N_noxref_24_c_8788_n N_noxref_26_c_8996_n ) capacitor c=0.00591245f \
 //x=79.005 //y=1.25 //x2=81.955 //y2=1.18
cc_5183 ( N_noxref_24_c_8789_n N_noxref_26_c_8996_n ) capacitor c=0.00340173f \
 //x=79.005 //y=1.56 //x2=81.955 //y2=1.18
cc_5184 ( N_noxref_24_c_8434_n N_noxref_26_c_8996_n ) capacitor c=2.04565e-19 \
 //x=79.005 //y=1.915 //x2=81.955 //y2=1.18
cc_5185 ( N_noxref_24_c_8437_n N_noxref_26_c_8996_n ) capacitor c=0.00500281f \
 //x=80.835 //y=1.21 //x2=81.955 //y2=1.18
cc_5186 ( N_noxref_24_c_8644_n N_noxref_26_c_8996_n ) capacitor c=0.00361177f \
 //x=80.835 //y=1.52 //x2=81.955 //y2=1.18
cc_5187 ( N_noxref_24_c_8439_n N_noxref_26_c_8996_n ) capacitor c=4.02408e-19 \
 //x=81.21 //y=0.71 //x2=81.955 //y2=1.18
cc_5188 ( N_noxref_24_c_8440_n N_noxref_26_c_8996_n ) capacitor c=0.0036677f \
 //x=81.21 //y=1.365 //x2=81.955 //y2=1.18
cc_5189 ( N_noxref_24_c_8443_n N_noxref_26_c_8996_n ) capacitor c=0.00776505f \
 //x=81.365 //y=1.21 //x2=81.955 //y2=1.18
cc_5190 ( N_noxref_24_c_8424_n N_noxref_26_c_9003_n ) capacitor c=0.00337373f \
 //x=79.065 //y=3.33 //x2=78.855 //y2=1.18
cc_5191 ( N_noxref_24_c_8781_n N_noxref_26_c_9003_n ) capacitor c=0.00154876f \
 //x=78.475 //y=1.25 //x2=78.855 //y2=1.18
cc_5192 ( N_noxref_24_c_8833_p N_noxref_26_c_9003_n ) capacitor c=4.52813e-19 \
 //x=78.85 //y=0.75 //x2=78.855 //y2=1.18
cc_5193 ( N_noxref_24_c_8834_p N_noxref_26_c_9003_n ) capacitor c=7.90416e-19 \
 //x=78.85 //y=1.405 //x2=78.855 //y2=1.18
cc_5194 ( N_noxref_24_c_8788_n N_noxref_26_c_9003_n ) capacitor c=4.79299e-19 \
 //x=79.005 //y=1.25 //x2=78.855 //y2=1.18
cc_5195 ( N_noxref_24_c_8789_n N_noxref_26_c_9003_n ) capacitor c=9.69054e-19 \
 //x=79.005 //y=1.56 //x2=78.855 //y2=1.18
cc_5196 ( N_noxref_24_M151_noxref_g N_noxref_26_c_9089_n ) capacitor \
 c=0.0179287f //x=81.37 //y=6.025 //x2=81.945 //y2=5.21
cc_5197 ( N_noxref_24_M150_noxref_g N_noxref_26_c_9045_n ) capacitor \
 c=0.0132916f //x=80.93 //y=6.025 //x2=81.235 //y2=5.21
cc_5198 ( N_noxref_24_c_8646_n N_noxref_26_c_9045_n ) capacitor c=0.00405122f \
 //x=81.295 //y=4.795 //x2=81.235 //y2=5.21
cc_5199 ( N_noxref_24_c_8433_n N_noxref_26_c_9010_n ) capacitor c=0.00334764f \
 //x=80.66 //y=2.08 //x2=82.51 //y2=4.07
cc_5200 ( N_noxref_24_c_8424_n N_noxref_26_M46_noxref_d ) capacitor \
 c=0.00415098f //x=79.065 //y=3.33 //x2=75.22 //y2=0.905
cc_5201 ( N_noxref_24_c_8424_n N_noxref_26_M48_noxref_d ) capacitor \
 c=0.00415178f //x=79.065 //y=3.33 //x2=78.55 //y2=0.905
cc_5202 ( N_noxref_24_c_8778_n N_noxref_26_M48_noxref_d ) capacitor \
 c=0.00217566f //x=78.475 //y=0.905 //x2=78.55 //y2=0.905
cc_5203 ( N_noxref_24_c_8781_n N_noxref_26_M48_noxref_d ) capacitor \
 c=0.00711747f //x=78.475 //y=1.25 //x2=78.55 //y2=0.905
cc_5204 ( N_noxref_24_c_8833_p N_noxref_26_M48_noxref_d ) capacitor \
 c=0.00234223f //x=78.85 //y=0.75 //x2=78.55 //y2=0.905
cc_5205 ( N_noxref_24_c_8834_p N_noxref_26_M48_noxref_d ) capacitor \
 c=0.00602848f //x=78.85 //y=1.405 //x2=78.55 //y2=0.905
cc_5206 ( N_noxref_24_c_8787_n N_noxref_26_M48_noxref_d ) capacitor \
 c=0.00132245f //x=79.005 //y=0.905 //x2=78.55 //y2=0.905
cc_5207 ( N_noxref_24_c_8788_n N_noxref_26_M48_noxref_d ) capacitor \
 c=0.004434f //x=79.005 //y=1.25 //x2=78.55 //y2=0.905
cc_5208 ( N_noxref_24_c_8789_n N_noxref_26_M48_noxref_d ) capacitor \
 c=0.00270197f //x=79.005 //y=1.56 //x2=78.55 //y2=0.905
cc_5209 ( N_noxref_24_M151_noxref_g N_noxref_26_M150_noxref_d ) capacitor \
 c=0.0130327f //x=81.37 //y=6.025 //x2=81.005 //y2=5.025
cc_5210 ( N_noxref_24_c_8511_n N_noxref_33_c_9544_n ) capacitor c=0.00623646f \
 //x=18.165 //y=1.56 //x2=17.945 //y2=1.495
cc_5211 ( N_noxref_24_c_8516_n N_noxref_33_c_9544_n ) capacitor c=0.00173579f \
 //x=18.13 //y=2.08 //x2=17.945 //y2=1.495
cc_5212 ( N_noxref_24_c_8428_n N_noxref_33_c_9545_n ) capacitor c=0.00156605f \
 //x=18.13 //y=2.08 //x2=18.83 //y2=0.53
cc_5213 ( N_noxref_24_c_8506_n N_noxref_33_c_9545_n ) capacitor c=0.0188655f \
 //x=18.165 //y=0.905 //x2=18.83 //y2=0.53
cc_5214 ( N_noxref_24_c_8514_n N_noxref_33_c_9545_n ) capacitor c=0.00656458f \
 //x=18.695 //y=0.905 //x2=18.83 //y2=0.53
cc_5215 ( N_noxref_24_c_8516_n N_noxref_33_c_9545_n ) capacitor c=2.1838e-19 \
 //x=18.13 //y=2.08 //x2=18.83 //y2=0.53
cc_5216 ( N_noxref_24_c_8506_n N_noxref_33_M10_noxref_s ) capacitor \
 c=0.00623646f //x=18.165 //y=0.905 //x2=16.84 //y2=0.365
cc_5217 ( N_noxref_24_c_8514_n N_noxref_33_M10_noxref_s ) capacitor \
 c=0.0143002f //x=18.695 //y=0.905 //x2=16.84 //y2=0.365
cc_5218 ( N_noxref_24_c_8515_n N_noxref_33_M10_noxref_s ) capacitor \
 c=0.00290153f //x=18.695 //y=1.25 //x2=16.84 //y2=0.365
cc_5219 ( N_noxref_24_M14_noxref_d N_noxref_34_M12_noxref_s ) capacitor \
 c=0.00309936f //x=23.005 //y=0.915 //x2=20.065 //y2=0.375
cc_5220 ( N_noxref_24_c_8430_n N_noxref_35_c_9645_n ) capacitor c=0.00457167f \
 //x=23.595 //y=1.665 //x2=23.595 //y2=0.54
cc_5221 ( N_noxref_24_M14_noxref_d N_noxref_35_c_9645_n ) capacitor \
 c=0.0115903f //x=23.005 //y=0.915 //x2=23.595 //y2=0.54
cc_5222 ( N_noxref_24_c_8735_n N_noxref_35_c_9657_n ) capacitor c=0.020048f \
 //x=23.28 //y=1.665 //x2=22.71 //y2=0.995
cc_5223 ( N_noxref_24_M14_noxref_d N_noxref_35_M13_noxref_d ) capacitor \
 c=5.27807e-19 //x=23.005 //y=0.915 //x2=21.47 //y2=0.91
cc_5224 ( N_noxref_24_c_8430_n N_noxref_35_M14_noxref_s ) capacitor \
 c=0.0196084f //x=23.595 //y=1.665 //x2=22.575 //y2=0.375
cc_5225 ( N_noxref_24_M14_noxref_d N_noxref_35_M14_noxref_s ) capacitor \
 c=0.0426444f //x=23.005 //y=0.915 //x2=22.575 //y2=0.375
cc_5226 ( N_noxref_24_c_8430_n N_noxref_36_c_9710_n ) capacitor c=3.04182e-19 \
 //x=23.595 //y=1.665 //x2=25.115 //y2=1.495
cc_5227 ( N_noxref_24_c_8424_n N_noxref_54_M45_noxref_s ) capacitor \
 c=0.00218253f //x=79.065 //y=3.33 //x2=73.82 //y2=0.365
cc_5228 ( N_noxref_24_c_8424_n N_noxref_55_c_10689_n ) capacitor c=0.00191103f \
 //x=79.065 //y=3.33 //x2=77.285 //y2=1.495
cc_5229 ( N_noxref_24_c_8424_n N_noxref_55_c_10672_n ) capacitor c=0.0095211f \
 //x=79.065 //y=3.33 //x2=78.17 //y2=1.58
cc_5230 ( N_noxref_24_c_8424_n N_noxref_55_c_10678_n ) capacitor c=0.00218253f \
 //x=79.065 //y=3.33 //x2=78.255 //y2=1.495
cc_5231 ( N_noxref_24_c_8434_n N_noxref_55_c_10678_n ) capacitor c=0.0028747f \
 //x=79.005 //y=1.915 //x2=78.255 //y2=1.495
cc_5232 ( N_noxref_24_c_8778_n N_noxref_55_c_10679_n ) capacitor c=0.021566f \
 //x=78.475 //y=0.905 //x2=79.14 //y2=0.53
cc_5233 ( N_noxref_24_c_8787_n N_noxref_55_c_10679_n ) capacitor c=0.00781103f \
 //x=79.005 //y=0.905 //x2=79.14 //y2=0.53
cc_5234 ( N_noxref_24_c_8426_n N_noxref_55_M47_noxref_s ) capacitor \
 c=5.34178e-19 //x=80.545 //y=2.08 //x2=77.15 //y2=0.365
cc_5235 ( N_noxref_24_c_8427_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.00116116f //x=79.295 //y=2.08 //x2=77.15 //y2=0.365
cc_5236 ( N_noxref_24_c_8431_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.0152989f //x=79.18 //y=2.08 //x2=77.15 //y2=0.365
cc_5237 ( N_noxref_24_c_8778_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.0064603f //x=78.475 //y=0.905 //x2=77.15 //y2=0.365
cc_5238 ( N_noxref_24_c_8781_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.00602248f //x=78.475 //y=1.25 //x2=77.15 //y2=0.365
cc_5239 ( N_noxref_24_c_8787_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.0321601f //x=79.005 //y=0.905 //x2=77.15 //y2=0.365
cc_5240 ( N_noxref_24_c_8789_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.00239072f //x=79.005 //y=1.56 //x2=77.15 //y2=0.365
cc_5241 ( N_noxref_24_c_8434_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.00784558f //x=79.005 //y=1.915 //x2=77.15 //y2=0.365
cc_5242 ( N_noxref_24_c_8426_n N_noxref_56_c_10757_n ) capacitor c=0.00169534f \
 //x=80.545 //y=2.08 //x2=80.615 //y2=1.495
cc_5243 ( N_noxref_24_c_8433_n N_noxref_56_c_10757_n ) capacitor c=0.016698f \
 //x=80.66 //y=2.08 //x2=80.615 //y2=1.495
cc_5244 ( N_noxref_24_c_8438_n N_noxref_56_c_10757_n ) capacitor c=0.0034165f \
 //x=80.835 //y=1.915 //x2=80.615 //y2=1.495
cc_5245 ( N_noxref_24_c_8444_n N_noxref_56_c_10757_n ) capacitor c=0.00531095f \
 //x=80.66 //y=2.08 //x2=80.615 //y2=1.495
cc_5246 ( N_noxref_24_c_8426_n N_noxref_56_c_10727_n ) capacitor c=0.00222439f \
 //x=80.545 //y=2.08 //x2=81.5 //y2=1.58
cc_5247 ( N_noxref_24_c_8433_n N_noxref_56_c_10727_n ) capacitor c=0.00587616f \
 //x=80.66 //y=2.08 //x2=81.5 //y2=1.58
cc_5248 ( N_noxref_24_c_8644_n N_noxref_56_c_10727_n ) capacitor c=0.0061593f \
 //x=80.835 //y=1.52 //x2=81.5 //y2=1.58
cc_5249 ( N_noxref_24_c_8438_n N_noxref_56_c_10727_n ) capacitor c=0.0142098f \
 //x=80.835 //y=1.915 //x2=81.5 //y2=1.58
cc_5250 ( N_noxref_24_c_8440_n N_noxref_56_c_10727_n ) capacitor c=0.00991953f \
 //x=81.21 //y=1.365 //x2=81.5 //y2=1.58
cc_5251 ( N_noxref_24_c_8443_n N_noxref_56_c_10727_n ) capacitor c=0.00339872f \
 //x=81.365 //y=1.21 //x2=81.5 //y2=1.58
cc_5252 ( N_noxref_24_c_8444_n N_noxref_56_c_10727_n ) capacitor c=0.00147967f \
 //x=80.66 //y=2.08 //x2=81.5 //y2=1.58
cc_5253 ( N_noxref_24_c_8438_n N_noxref_56_c_10733_n ) capacitor c=6.71402e-19 \
 //x=80.835 //y=1.915 //x2=81.585 //y2=1.495
cc_5254 ( N_noxref_24_c_8435_n N_noxref_56_M49_noxref_s ) capacitor \
 c=0.0314164f //x=80.835 //y=0.865 //x2=80.48 //y2=0.365
cc_5255 ( N_noxref_24_c_8644_n N_noxref_56_M49_noxref_s ) capacitor \
 c=0.00110192f //x=80.835 //y=1.52 //x2=80.48 //y2=0.365
cc_5256 ( N_noxref_24_c_8441_n N_noxref_56_M49_noxref_s ) capacitor \
 c=0.0132463f //x=81.365 //y=0.865 //x2=80.48 //y2=0.365
cc_5257 ( N_noxref_25_c_8920_n N_noxref_26_c_9089_n ) capacitor c=0.00102709f \
 //x=81.505 //y=6.91 //x2=81.945 //y2=5.21
cc_5258 ( N_noxref_25_c_8921_n N_noxref_26_c_9089_n ) capacitor c=0.00101874f \
 //x=82.385 //y=6.91 //x2=81.945 //y2=5.21
cc_5259 ( N_noxref_25_M151_noxref_d N_noxref_26_c_9089_n ) capacitor \
 c=0.012404f //x=81.445 //y=5.025 //x2=81.945 //y2=5.21
cc_5260 ( N_noxref_25_c_8898_n N_noxref_26_c_9045_n ) capacitor c=0.00602307f \
 //x=80.595 //y=5.21 //x2=81.235 //y2=5.21
cc_5261 ( N_noxref_25_c_8906_n N_noxref_26_c_9045_n ) capacitor c=0.0683084f \
 //x=80.71 //y=5.21 //x2=81.235 //y2=5.21
cc_5262 ( N_noxref_25_c_8921_n N_noxref_26_c_9046_n ) capacitor c=0.00173777f \
 //x=82.385 //y=6.91 //x2=82.425 //y2=5.21
cc_5263 ( N_noxref_25_M153_noxref_d N_noxref_26_c_9046_n ) capacitor \
 c=0.0154399f //x=82.325 //y=5.025 //x2=82.425 //y2=5.21
cc_5264 ( N_noxref_25_c_8906_n N_noxref_26_c_9010_n ) capacitor c=3.02032e-19 \
 //x=80.71 //y=5.21 //x2=82.51 //y2=4.07
cc_5265 ( N_noxref_25_c_8898_n N_noxref_26_M150_noxref_d ) capacitor \
 c=8.04912e-19 //x=80.595 //y=5.21 //x2=81.005 //y2=5.025
cc_5266 ( N_noxref_25_c_8920_n N_noxref_26_M150_noxref_d ) capacitor \
 c=0.0117542f //x=81.505 //y=6.91 //x2=81.005 //y2=5.025
cc_5267 ( N_noxref_25_M151_noxref_d N_noxref_26_M150_noxref_d ) capacitor \
 c=0.0458293f //x=81.445 //y=5.025 //x2=81.005 //y2=5.025
cc_5268 ( N_noxref_25_c_8906_n N_noxref_26_M152_noxref_d ) capacitor \
 c=9.91979e-19 //x=80.71 //y=5.21 //x2=81.885 //y2=5.025
cc_5269 ( N_noxref_25_c_8921_n N_noxref_26_M152_noxref_d ) capacitor \
 c=0.0118172f //x=82.385 //y=6.91 //x2=81.885 //y2=5.025
cc_5270 ( N_noxref_25_M151_noxref_d N_noxref_26_M152_noxref_d ) capacitor \
 c=0.0458293f //x=81.445 //y=5.025 //x2=81.885 //y2=5.025
cc_5271 ( N_noxref_25_M153_noxref_d N_noxref_26_M152_noxref_d ) capacitor \
 c=0.0458293f //x=82.325 //y=5.025 //x2=81.885 //y2=5.025
cc_5272 ( N_noxref_26_c_8988_n N_noxref_54_c_10623_n ) capacitor c=0.00641749f \
 //x=78.625 //y=1.18 //x2=75.81 //y2=0.53
cc_5273 ( N_noxref_26_c_8995_n N_noxref_54_c_10623_n ) capacitor c=0.00219859f \
 //x=75.525 //y=1.18 //x2=75.81 //y2=0.53
cc_5274 ( N_noxref_26_M46_noxref_d N_noxref_54_c_10623_n ) capacitor \
 c=0.0136817f //x=75.22 //y=0.905 //x2=75.81 //y2=0.53
cc_5275 ( N_noxref_26_c_8988_n N_noxref_54_M45_noxref_s ) capacitor \
 c=0.0211151f //x=78.625 //y=1.18 //x2=73.82 //y2=0.365
cc_5276 ( N_noxref_26_c_8995_n N_noxref_54_M45_noxref_s ) capacitor \
 c=0.00804471f //x=75.525 //y=1.18 //x2=73.82 //y2=0.365
cc_5277 ( N_noxref_26_M46_noxref_d N_noxref_54_M45_noxref_s ) capacitor \
 c=0.0458734f //x=75.22 //y=0.905 //x2=73.82 //y2=0.365
cc_5278 ( N_noxref_26_c_8988_n N_noxref_55_c_10672_n ) capacitor c=0.0230023f \
 //x=78.625 //y=1.18 //x2=78.17 //y2=1.58
cc_5279 ( N_noxref_26_c_8988_n N_noxref_55_c_10679_n ) capacitor c=0.00641749f \
 //x=78.625 //y=1.18 //x2=79.14 //y2=0.53
cc_5280 ( N_noxref_26_c_8996_n N_noxref_55_c_10679_n ) capacitor c=0.00641749f \
 //x=81.955 //y=1.18 //x2=79.14 //y2=0.53
cc_5281 ( N_noxref_26_c_9003_n N_noxref_55_c_10679_n ) capacitor c=0.0015838f \
 //x=78.855 //y=1.18 //x2=79.14 //y2=0.53
cc_5282 ( N_noxref_26_M48_noxref_d N_noxref_55_c_10679_n ) capacitor \
 c=0.0130616f //x=78.55 //y=0.905 //x2=79.14 //y2=0.53
cc_5283 ( N_noxref_26_c_8988_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.045024f //x=78.625 //y=1.18 //x2=77.15 //y2=0.365
cc_5284 ( N_noxref_26_c_8996_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.019112f //x=81.955 //y=1.18 //x2=77.15 //y2=0.365
cc_5285 ( N_noxref_26_c_9003_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.00279707f //x=78.855 //y=1.18 //x2=77.15 //y2=0.365
cc_5286 ( N_noxref_26_M48_noxref_d N_noxref_55_M47_noxref_s ) capacitor \
 c=0.0444718f //x=78.55 //y=0.905 //x2=77.15 //y2=0.365
cc_5287 ( N_noxref_26_c_9096_n N_noxref_56_c_10757_n ) capacitor c=2.73698e-19 \
 //x=82.155 //y=1.645 //x2=80.615 //y2=1.495
cc_5288 ( N_noxref_26_c_8996_n N_noxref_56_c_10727_n ) capacitor c=0.0234642f \
 //x=81.955 //y=1.18 //x2=81.5 //y2=1.58
cc_5289 ( N_noxref_26_c_9096_n N_noxref_56_c_10733_n ) capacitor c=0.0195484f \
 //x=82.155 //y=1.645 //x2=81.585 //y2=1.495
cc_5290 ( N_noxref_26_c_8996_n N_noxref_56_c_10734_n ) capacitor c=0.0069137f \
 //x=81.955 //y=1.18 //x2=82.47 //y2=0.53
cc_5291 ( N_noxref_26_c_9008_n N_noxref_56_c_10734_n ) capacitor c=0.00458011f \
 //x=82.425 //y=1.645 //x2=82.47 //y2=0.53
cc_5292 ( N_noxref_26_M50_noxref_d N_noxref_56_c_10734_n ) capacitor \
 c=0.0132979f //x=81.88 //y=0.905 //x2=82.47 //y2=0.53
cc_5293 ( N_noxref_26_c_8996_n N_noxref_56_M49_noxref_s ) capacitor \
 c=0.0513705f //x=81.955 //y=1.18 //x2=80.48 //y2=0.365
cc_5294 ( N_noxref_26_c_9008_n N_noxref_56_M49_noxref_s ) capacitor \
 c=0.0154295f //x=82.425 //y=1.645 //x2=80.48 //y2=0.365
cc_5295 ( N_noxref_26_M50_noxref_d N_noxref_56_M49_noxref_s ) capacitor \
 c=0.0438441f //x=81.88 //y=0.905 //x2=80.48 //y2=0.365
cc_5296 ( N_noxref_26_c_9004_n Q ) capacitor c=0.00467401f //x=83.875 //y=4.07 \
 //x2=84.73 //y2=2.22
cc_5297 ( N_noxref_26_c_9010_n Q ) capacitor c=0.00120943f //x=82.51 //y=4.07 \
 //x2=84.73 //y2=2.22
cc_5298 ( N_noxref_26_c_9011_n Q ) capacitor c=0.0711602f //x=83.99 //y=2.085 \
 //x2=84.73 //y2=2.22
cc_5299 ( N_noxref_26_c_9023_n Q ) capacitor c=8.49451e-19 //x=83.99 //y=2.085 \
 //x2=84.73 //y2=2.22
cc_5300 ( N_noxref_26_c_9208_p N_Q_c_10784_n ) capacitor c=0.0023507f \
 //x=84.475 //y=1.41 //x2=84.645 //y2=2.08
cc_5301 ( N_noxref_26_c_9023_n N_Q_c_10808_n ) capacitor c=0.0167852f \
 //x=83.99 //y=2.085 //x2=84.445 //y2=2.08
cc_5302 ( N_noxref_26_c_9060_n N_Q_c_10794_n ) capacitor c=0.0101013f \
 //x=84.51 //y=4.79 //x2=84.645 //y2=4.58
cc_5303 ( N_noxref_26_c_9011_n N_Q_c_10797_n ) capacitor c=0.0250878f \
 //x=83.99 //y=2.085 //x2=84.45 //y2=4.58
cc_5304 ( N_noxref_26_c_9061_n N_Q_c_10797_n ) capacitor c=0.00962086f \
 //x=84.22 //y=4.79 //x2=84.45 //y2=4.58
cc_5305 ( N_noxref_26_c_9010_n N_Q_M51_noxref_d ) capacitor c=3.32382e-19 \
 //x=82.51 //y=4.07 //x2=84.175 //y2=0.91
cc_5306 ( N_noxref_26_c_9011_n N_Q_M51_noxref_d ) capacitor c=0.0177062f \
 //x=83.99 //y=2.085 //x2=84.175 //y2=0.91
cc_5307 ( N_noxref_26_c_9016_n N_Q_M51_noxref_d ) capacitor c=0.00218556f \
 //x=84.1 //y=0.91 //x2=84.175 //y2=0.91
cc_5308 ( N_noxref_26_c_9216_p N_Q_M51_noxref_d ) capacitor c=0.00347355f \
 //x=84.1 //y=1.255 //x2=84.175 //y2=0.91
cc_5309 ( N_noxref_26_c_9217_p N_Q_M51_noxref_d ) capacitor c=0.00742431f \
 //x=84.1 //y=1.565 //x2=84.175 //y2=0.91
cc_5310 ( N_noxref_26_c_9018_n N_Q_M51_noxref_d ) capacitor c=0.00957707f \
 //x=84.1 //y=1.92 //x2=84.175 //y2=0.91
cc_5311 ( N_noxref_26_c_9019_n N_Q_M51_noxref_d ) capacitor c=0.00220879f \
 //x=84.475 //y=0.755 //x2=84.175 //y2=0.91
cc_5312 ( N_noxref_26_c_9208_p N_Q_M51_noxref_d ) capacitor c=0.0138447f \
 //x=84.475 //y=1.41 //x2=84.175 //y2=0.91
cc_5313 ( N_noxref_26_c_9020_n N_Q_M51_noxref_d ) capacitor c=0.00218624f \
 //x=84.63 //y=0.91 //x2=84.175 //y2=0.91
cc_5314 ( N_noxref_26_c_9022_n N_Q_M51_noxref_d ) capacitor c=0.00601286f \
 //x=84.63 //y=1.255 //x2=84.175 //y2=0.91
cc_5315 ( N_noxref_26_c_9010_n N_Q_M154_noxref_d ) capacitor c=6.32888e-19 \
 //x=82.51 //y=4.07 //x2=84.22 //y2=5.02
cc_5316 ( N_noxref_26_M154_noxref_g N_Q_M154_noxref_d ) capacitor c=0.0219309f \
 //x=84.145 //y=6.02 //x2=84.22 //y2=5.02
cc_5317 ( N_noxref_26_M155_noxref_g N_Q_M154_noxref_d ) capacitor c=0.021902f \
 //x=84.585 //y=6.02 //x2=84.22 //y2=5.02
cc_5318 ( N_noxref_26_c_9060_n N_Q_M154_noxref_d ) capacitor c=0.0148755f \
 //x=84.51 //y=4.79 //x2=84.22 //y2=5.02
cc_5319 ( N_noxref_26_c_9061_n N_Q_M154_noxref_d ) capacitor c=0.00307344f \
 //x=84.22 //y=4.79 //x2=84.22 //y2=5.02
cc_5320 ( N_noxref_27_c_9238_n N_noxref_28_M2_noxref_s ) capacitor \
 c=0.00199452f //x=2.635 //y=0.615 //x2=3.785 //y2=0.375
cc_5321 ( N_noxref_28_c_9285_n N_noxref_29_c_9329_n ) capacitor c=0.0133059f \
 //x=5.775 //y=0.54 //x2=6.345 //y2=0.995
cc_5322 ( N_noxref_28_c_9304_n N_noxref_29_c_9329_n ) capacitor c=0.0100097f \
 //x=5.775 //y=1.59 //x2=6.345 //y2=0.995
cc_5323 ( N_noxref_28_M2_noxref_s N_noxref_29_c_9329_n ) capacitor \
 c=0.0224457f //x=3.785 //y=0.375 //x2=6.345 //y2=0.995
cc_5324 ( N_noxref_28_M2_noxref_s N_noxref_29_c_9331_n ) capacitor \
 c=0.0180035f //x=3.785 //y=0.375 //x2=6.43 //y2=0.625
cc_5325 ( N_noxref_28_c_9285_n N_noxref_29_M3_noxref_d ) capacitor \
 c=0.0128027f //x=5.775 //y=0.54 //x2=5.19 //y2=0.91
cc_5326 ( N_noxref_28_c_9304_n N_noxref_29_M3_noxref_d ) capacitor \
 c=0.00879751f //x=5.775 //y=1.59 //x2=5.19 //y2=0.91
cc_5327 ( N_noxref_28_M2_noxref_s N_noxref_29_M3_noxref_d ) capacitor \
 c=0.0159202f //x=3.785 //y=0.375 //x2=5.19 //y2=0.91
cc_5328 ( N_noxref_28_M2_noxref_s N_noxref_29_M4_noxref_s ) capacitor \
 c=0.0213553f //x=3.785 //y=0.375 //x2=6.295 //y2=0.375
cc_5329 ( N_noxref_29_c_9336_n N_noxref_30_M5_noxref_s ) capacitor \
 c=0.00191848f //x=7.4 //y=0.625 //x2=8.595 //y2=0.375
cc_5330 ( N_noxref_30_c_9388_n N_noxref_31_c_9434_n ) capacitor c=0.0131801f \
 //x=10.585 //y=0.54 //x2=11.155 //y2=0.995
cc_5331 ( N_noxref_30_c_9412_n N_noxref_31_c_9434_n ) capacitor c=0.00980353f \
 //x=10.585 //y=1.59 //x2=11.155 //y2=0.995
cc_5332 ( N_noxref_30_M5_noxref_s N_noxref_31_c_9434_n ) capacitor \
 c=0.0221661f //x=8.595 //y=0.375 //x2=11.155 //y2=0.995
cc_5333 ( N_noxref_30_M5_noxref_s N_noxref_31_c_9436_n ) capacitor \
 c=0.0180035f //x=8.595 //y=0.375 //x2=11.24 //y2=0.625
cc_5334 ( N_noxref_30_c_9388_n N_noxref_31_M6_noxref_d ) capacitor \
 c=0.0128066f //x=10.585 //y=0.54 //x2=10 //y2=0.91
cc_5335 ( N_noxref_30_c_9412_n N_noxref_31_M6_noxref_d ) capacitor \
 c=0.00879078f //x=10.585 //y=1.59 //x2=10 //y2=0.91
cc_5336 ( N_noxref_30_M5_noxref_s N_noxref_31_M6_noxref_d ) capacitor \
 c=0.0159202f //x=8.595 //y=0.375 //x2=10 //y2=0.91
cc_5337 ( N_noxref_30_M5_noxref_s N_noxref_31_M7_noxref_s ) capacitor \
 c=0.0213553f //x=8.595 //y=0.375 //x2=11.105 //y2=0.375
cc_5338 ( N_noxref_31_c_9441_n N_noxref_32_M8_noxref_s ) capacitor \
 c=0.00164795f //x=12.21 //y=0.625 //x2=13.51 //y2=0.365
cc_5339 ( N_noxref_32_c_9496_n N_noxref_33_M10_noxref_s ) capacitor \
 c=0.00174327f //x=15.585 //y=0.615 //x2=16.84 //y2=0.365
cc_5340 ( N_noxref_33_c_9547_n N_noxref_34_M12_noxref_s ) capacitor \
 c=0.00199452f //x=18.915 //y=0.615 //x2=20.065 //y2=0.375
cc_5341 ( N_noxref_34_c_9595_n N_noxref_35_c_9640_n ) capacitor c=0.0131801f \
 //x=22.055 //y=0.54 //x2=22.625 //y2=0.995
cc_5342 ( N_noxref_34_c_9619_n N_noxref_35_c_9640_n ) capacitor c=0.00980353f \
 //x=22.055 //y=1.59 //x2=22.625 //y2=0.995
cc_5343 ( N_noxref_34_M12_noxref_s N_noxref_35_c_9640_n ) capacitor \
 c=0.0221661f //x=20.065 //y=0.375 //x2=22.625 //y2=0.995
cc_5344 ( N_noxref_34_M12_noxref_s N_noxref_35_c_9642_n ) capacitor \
 c=0.0180035f //x=20.065 //y=0.375 //x2=22.71 //y2=0.625
cc_5345 ( N_noxref_34_c_9595_n N_noxref_35_M13_noxref_d ) capacitor \
 c=0.0127176f //x=22.055 //y=0.54 //x2=21.47 //y2=0.91
cc_5346 ( N_noxref_34_c_9619_n N_noxref_35_M13_noxref_d ) capacitor \
 c=0.0086073f //x=22.055 //y=1.59 //x2=21.47 //y2=0.91
cc_5347 ( N_noxref_34_M12_noxref_s N_noxref_35_M13_noxref_d ) capacitor \
 c=0.0159202f //x=20.065 //y=0.375 //x2=21.47 //y2=0.91
cc_5348 ( N_noxref_34_M12_noxref_s N_noxref_35_M14_noxref_s ) capacitor \
 c=0.0213553f //x=20.065 //y=0.375 //x2=22.575 //y2=0.375
cc_5349 ( N_noxref_35_c_9647_n N_noxref_36_M15_noxref_s ) capacitor \
 c=0.00164795f //x=23.68 //y=0.625 //x2=24.98 //y2=0.365
cc_5350 ( N_noxref_36_c_9702_n N_noxref_37_M17_noxref_s ) capacitor \
 c=0.00199452f //x=27.055 //y=0.615 //x2=28.205 //y2=0.375
cc_5351 ( N_noxref_37_c_9750_n N_noxref_38_c_9792_n ) capacitor c=0.0131877f \
 //x=30.195 //y=0.54 //x2=30.765 //y2=0.995
cc_5352 ( N_noxref_37_c_9773_n N_noxref_38_c_9792_n ) capacitor c=0.00981707f \
 //x=30.195 //y=1.59 //x2=30.765 //y2=0.995
cc_5353 ( N_noxref_37_M17_noxref_s N_noxref_38_c_9792_n ) capacitor \
 c=0.0221661f //x=28.205 //y=0.375 //x2=30.765 //y2=0.995
cc_5354 ( N_noxref_37_M17_noxref_s N_noxref_38_c_9794_n ) capacitor \
 c=0.0180035f //x=28.205 //y=0.375 //x2=30.85 //y2=0.625
cc_5355 ( N_noxref_37_c_9750_n N_noxref_38_M18_noxref_d ) capacitor \
 c=0.0127191f //x=30.195 //y=0.54 //x2=29.61 //y2=0.91
cc_5356 ( N_noxref_37_c_9773_n N_noxref_38_M18_noxref_d ) capacitor \
 c=0.00861161f //x=30.195 //y=1.59 //x2=29.61 //y2=0.91
cc_5357 ( N_noxref_37_M17_noxref_s N_noxref_38_M18_noxref_d ) capacitor \
 c=0.0159202f //x=28.205 //y=0.375 //x2=29.61 //y2=0.91
cc_5358 ( N_noxref_37_M17_noxref_s N_noxref_38_M19_noxref_s ) capacitor \
 c=0.0213553f //x=28.205 //y=0.375 //x2=30.715 //y2=0.375
cc_5359 ( N_noxref_38_c_9799_n N_noxref_39_M20_noxref_s ) capacitor \
 c=0.00191848f //x=31.82 //y=0.625 //x2=33.015 //y2=0.375
cc_5360 ( N_noxref_39_c_9851_n N_noxref_40_c_9896_n ) capacitor c=0.0131801f \
 //x=35.005 //y=0.54 //x2=35.575 //y2=0.995
cc_5361 ( N_noxref_39_c_9876_n N_noxref_40_c_9896_n ) capacitor c=0.00980353f \
 //x=35.005 //y=1.59 //x2=35.575 //y2=0.995
cc_5362 ( N_noxref_39_M20_noxref_s N_noxref_40_c_9896_n ) capacitor \
 c=0.0221661f //x=33.015 //y=0.375 //x2=35.575 //y2=0.995
cc_5363 ( N_noxref_39_M20_noxref_s N_noxref_40_c_9898_n ) capacitor \
 c=0.0180035f //x=33.015 //y=0.375 //x2=35.66 //y2=0.625
cc_5364 ( N_noxref_39_c_9851_n N_noxref_40_M21_noxref_d ) capacitor \
 c=0.0127176f //x=35.005 //y=0.54 //x2=34.42 //y2=0.91
cc_5365 ( N_noxref_39_c_9876_n N_noxref_40_M21_noxref_d ) capacitor \
 c=0.0086073f //x=35.005 //y=1.59 //x2=34.42 //y2=0.91
cc_5366 ( N_noxref_39_M20_noxref_s N_noxref_40_M21_noxref_d ) capacitor \
 c=0.0159202f //x=33.015 //y=0.375 //x2=34.42 //y2=0.91
cc_5367 ( N_noxref_39_M20_noxref_s N_noxref_40_M22_noxref_s ) capacitor \
 c=0.0213553f //x=33.015 //y=0.375 //x2=35.525 //y2=0.375
cc_5368 ( N_noxref_40_c_9903_n N_noxref_41_M23_noxref_s ) capacitor \
 c=0.00164795f //x=36.63 //y=0.625 //x2=37.93 //y2=0.365
cc_5369 ( N_noxref_41_c_9958_n N_noxref_42_M25_noxref_s ) capacitor \
 c=0.00174327f //x=40.005 //y=0.615 //x2=41.26 //y2=0.365
cc_5370 ( N_noxref_42_c_10009_n N_noxref_43_M27_noxref_s ) capacitor \
 c=0.00199452f //x=43.335 //y=0.615 //x2=44.485 //y2=0.375
cc_5371 ( N_noxref_43_c_10057_n N_noxref_44_c_10102_n ) capacitor c=0.0131801f \
 //x=46.475 //y=0.54 //x2=47.045 //y2=0.995
cc_5372 ( N_noxref_43_c_10082_n N_noxref_44_c_10102_n ) capacitor \
 c=0.00980353f //x=46.475 //y=1.59 //x2=47.045 //y2=0.995
cc_5373 ( N_noxref_43_M27_noxref_s N_noxref_44_c_10102_n ) capacitor \
 c=0.0221661f //x=44.485 //y=0.375 //x2=47.045 //y2=0.995
cc_5374 ( N_noxref_43_M27_noxref_s N_noxref_44_c_10104_n ) capacitor \
 c=0.0180035f //x=44.485 //y=0.375 //x2=47.13 //y2=0.625
cc_5375 ( N_noxref_43_c_10057_n N_noxref_44_M28_noxref_d ) capacitor \
 c=0.0127176f //x=46.475 //y=0.54 //x2=45.89 //y2=0.91
cc_5376 ( N_noxref_43_c_10082_n N_noxref_44_M28_noxref_d ) capacitor \
 c=0.0086073f //x=46.475 //y=1.59 //x2=45.89 //y2=0.91
cc_5377 ( N_noxref_43_M27_noxref_s N_noxref_44_M28_noxref_d ) capacitor \
 c=0.0159202f //x=44.485 //y=0.375 //x2=45.89 //y2=0.91
cc_5378 ( N_noxref_43_M27_noxref_s N_noxref_44_M29_noxref_s ) capacitor \
 c=0.0213553f //x=44.485 //y=0.375 //x2=46.995 //y2=0.375
cc_5379 ( N_noxref_44_c_10109_n N_noxref_45_M30_noxref_s ) capacitor \
 c=0.00164795f //x=48.1 //y=0.625 //x2=49.4 //y2=0.365
cc_5380 ( N_noxref_45_c_10164_n N_noxref_46_M32_noxref_s ) capacitor \
 c=0.00199452f //x=51.475 //y=0.615 //x2=52.625 //y2=0.375
cc_5381 ( N_noxref_46_c_10212_n N_noxref_47_c_10254_n ) capacitor c=0.0131877f \
 //x=54.615 //y=0.54 //x2=55.185 //y2=0.995
cc_5382 ( N_noxref_46_c_10234_n N_noxref_47_c_10254_n ) capacitor \
 c=0.00981707f //x=54.615 //y=1.59 //x2=55.185 //y2=0.995
cc_5383 ( N_noxref_46_M32_noxref_s N_noxref_47_c_10254_n ) capacitor \
 c=0.0221661f //x=52.625 //y=0.375 //x2=55.185 //y2=0.995
cc_5384 ( N_noxref_46_M32_noxref_s N_noxref_47_c_10256_n ) capacitor \
 c=0.0180035f //x=52.625 //y=0.375 //x2=55.27 //y2=0.625
cc_5385 ( N_noxref_46_c_10212_n N_noxref_47_M33_noxref_d ) capacitor \
 c=0.0127191f //x=54.615 //y=0.54 //x2=54.03 //y2=0.91
cc_5386 ( N_noxref_46_c_10234_n N_noxref_47_M33_noxref_d ) capacitor \
 c=0.00861161f //x=54.615 //y=1.59 //x2=54.03 //y2=0.91
cc_5387 ( N_noxref_46_M32_noxref_s N_noxref_47_M33_noxref_d ) capacitor \
 c=0.0159202f //x=52.625 //y=0.375 //x2=54.03 //y2=0.91
cc_5388 ( N_noxref_46_M32_noxref_s N_noxref_47_M34_noxref_s ) capacitor \
 c=0.0213553f //x=52.625 //y=0.375 //x2=55.135 //y2=0.375
cc_5389 ( N_noxref_47_c_10261_n N_noxref_48_M35_noxref_s ) capacitor \
 c=0.00191848f //x=56.24 //y=0.625 //x2=57.435 //y2=0.375
cc_5390 ( N_noxref_48_c_10313_n N_noxref_49_c_10358_n ) capacitor c=0.0131801f \
 //x=59.425 //y=0.54 //x2=59.995 //y2=0.995
cc_5391 ( N_noxref_48_c_10338_n N_noxref_49_c_10358_n ) capacitor \
 c=0.00980353f //x=59.425 //y=1.59 //x2=59.995 //y2=0.995
cc_5392 ( N_noxref_48_M35_noxref_s N_noxref_49_c_10358_n ) capacitor \
 c=0.0221661f //x=57.435 //y=0.375 //x2=59.995 //y2=0.995
cc_5393 ( N_noxref_48_M35_noxref_s N_noxref_49_c_10360_n ) capacitor \
 c=0.0180035f //x=57.435 //y=0.375 //x2=60.08 //y2=0.625
cc_5394 ( N_noxref_48_c_10313_n N_noxref_49_M36_noxref_d ) capacitor \
 c=0.0127176f //x=59.425 //y=0.54 //x2=58.84 //y2=0.91
cc_5395 ( N_noxref_48_c_10338_n N_noxref_49_M36_noxref_d ) capacitor \
 c=0.0086073f //x=59.425 //y=1.59 //x2=58.84 //y2=0.91
cc_5396 ( N_noxref_48_M35_noxref_s N_noxref_49_M36_noxref_d ) capacitor \
 c=0.0159202f //x=57.435 //y=0.375 //x2=58.84 //y2=0.91
cc_5397 ( N_noxref_48_M35_noxref_s N_noxref_49_M37_noxref_s ) capacitor \
 c=0.0213553f //x=57.435 //y=0.375 //x2=59.945 //y2=0.375
cc_5398 ( N_noxref_49_c_10365_n N_noxref_50_M38_noxref_s ) capacitor \
 c=0.00164795f //x=61.05 //y=0.625 //x2=62.35 //y2=0.365
cc_5399 ( N_noxref_50_c_10420_n N_noxref_51_M40_noxref_s ) capacitor \
 c=0.00174327f //x=64.425 //y=0.615 //x2=65.68 //y2=0.365
cc_5400 ( N_noxref_51_c_10471_n N_noxref_52_M42_noxref_s ) capacitor \
 c=0.00199452f //x=67.755 //y=0.615 //x2=68.905 //y2=0.375
cc_5401 ( N_noxref_52_c_10519_n N_noxref_53_c_10563_n ) capacitor c=0.0132328f \
 //x=70.895 //y=0.54 //x2=71.465 //y2=0.995
cc_5402 ( N_noxref_52_c_10527_n N_noxref_53_c_10563_n ) capacitor \
 c=0.00988406f //x=70.895 //y=1.59 //x2=71.465 //y2=0.995
cc_5403 ( N_noxref_52_M42_noxref_s N_noxref_53_c_10563_n ) capacitor \
 c=0.0226274f //x=68.905 //y=0.375 //x2=71.465 //y2=0.995
cc_5404 ( N_noxref_52_M42_noxref_s N_noxref_53_c_10565_n ) capacitor \
 c=0.0180035f //x=68.905 //y=0.375 //x2=71.55 //y2=0.625
cc_5405 ( N_noxref_52_c_10519_n N_noxref_53_M43_noxref_d ) capacitor \
 c=0.0127176f //x=70.895 //y=0.54 //x2=70.31 //y2=0.91
cc_5406 ( N_noxref_52_c_10527_n N_noxref_53_M43_noxref_d ) capacitor \
 c=0.0086073f //x=70.895 //y=1.59 //x2=70.31 //y2=0.91
cc_5407 ( N_noxref_52_M42_noxref_s N_noxref_53_M43_noxref_d ) capacitor \
 c=0.0159202f //x=68.905 //y=0.375 //x2=70.31 //y2=0.91
cc_5408 ( N_noxref_52_M42_noxref_s N_noxref_53_M44_noxref_s ) capacitor \
 c=0.0213553f //x=68.905 //y=0.375 //x2=71.415 //y2=0.375
cc_5409 ( N_noxref_53_c_10570_n N_noxref_54_M45_noxref_s ) capacitor \
 c=0.00195059f //x=72.52 //y=0.625 //x2=73.82 //y2=0.365
cc_5410 ( N_noxref_54_M45_noxref_s N_noxref_55_c_10689_n ) capacitor \
 c=0.0011299f //x=73.82 //y=0.365 //x2=77.285 //y2=1.495
cc_5411 ( N_noxref_54_c_10625_n N_noxref_55_M47_noxref_s ) capacitor \
 c=0.0011299f //x=75.895 //y=0.615 //x2=77.15 //y2=0.365
cc_5412 ( N_noxref_55_M47_noxref_s N_noxref_56_c_10757_n ) capacitor \
 c=0.0011299f //x=77.15 //y=0.365 //x2=80.615 //y2=1.495
cc_5413 ( N_noxref_55_c_10681_n N_noxref_56_M49_noxref_s ) capacitor \
 c=0.0011299f //x=79.225 //y=0.615 //x2=80.48 //y2=0.365
