* SPICE3 file created from DFFRNQNX1.ext - technology: sky130A

.subckt DFFRNQNX1 QN D CLK RN VPB VNB
X0 VPB CLK a_277_1004# VPB sky130_fd_pr__pfet_01v8 ad=1.24e+13p pd=1.004e+08u as=0p ps=0u w=2e+06u l=150000u M=2
X1 VPB a_277_1004# QN VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.74e+12p ps=1.374e+07u w=2e+06u l=150000u M=2
X2 a_599_943# RN VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X3 QN a_4151_943# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X4 VNB a_147_159# a_91_75# VNB sky130_fd_pr__nfet_01v8 ad=1.0746e+12p pd=9.42e+06u as=0p ps=0u w=3e+06u l=150000u
X5 a_147_159# CLK VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X6 a_4151_943# QN VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X7 QN a_4151_943# a_3924_182# VNB sky130_fd_pr__nfet_01v8 ad=1.791e+11p pd=1.57e+06u as=0p ps=0u w=3e+06u l=150000u
X8 VPB a_599_943# a_277_1004# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X9 VPB a_147_159# a_2141_1004# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X10 VPB a_2141_1004# a_147_159# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X11 a_147_159# RN VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X12 a_4151_943# a_147_159# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X13 a_372_182# CLK a_91_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X14 VNB a_277_1004# a_3643_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X15 a_277_1004# a_147_159# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X16 VNB QN a_4626_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X17 VPB a_277_1004# a_599_943# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X18 a_599_943# RN a_1334_182# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X19 VNB a_599_943# a_2036_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X20 VNB a_2141_1004# a_2681_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X21 a_2141_1004# a_599_943# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X22 a_3924_182# RN a_3643_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X23 VPB a_1304_166# a_599_943# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X24 VPB RN QN VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X25 VNB a_277_1004# a_1053_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X26 a_2962_182# CLK a_2681_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X27 a_1334_182# a_1304_166# a_1053_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X28 a_4151_943# a_147_159# a_4626_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X29 a_2141_1004# a_147_159# a_2036_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X30 a_277_1004# a_599_943# a_372_182# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X31 a_147_159# RN a_2962_182# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
C0 VPB a_147_159# 2.82fF
.ends
