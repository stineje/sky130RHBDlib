* SPICE3 file created from DLATCHN.ext - technology: sky130A

.subckt DLATCHN Q D GATE_N VDD GND
X0 VDD a_1739_182 a_3239_1005 VDD pshort w=2 l=0.15 M=2
X1 a_3905_1005 a_2849_182 a_3451_383 VDD pshort w=2 l=0.15 M=2
X2 VDD D a_629_182 VDD pshort w=2 l=0.15 M=2
X3 a_1105_1004 a_185_182 VDD VDD pshort w=2 l=0.15 M=2
X4 Q a_3451_383 GND GND nshort w=3 l=0.15
X5 a_185_182 GATE_N GND GND nshort w=3 l=0.15
X6 Q a_3451_383 a_3239_1005 VDD pshort w=2 l=0.15 M=2
X7 VDD a_2215_1004 a_2849_182 VDD pshort w=2 l=0.15 M=2
X8 VDD Q a_3905_1005 VDD pshort w=2 l=0.15 M=2
X9 a_1739_182 a_1105_1004 VDD VDD pshort w=2 l=0.15 M=2
X10 VDD GATE_N a_185_182 VDD pshort w=2 l=0.15 M=2
X11 a_2215_1004 a_185_182 VDD VDD pshort w=2 l=0.15 M=2
X12 GND a_629_182 a_1000_73 GND nshort w=3 l=0.15
X13 a_1739_182 a_1105_1004 GND GND nshort w=3 l=0.15
X14 a_2215_1004 D VDD VDD pshort w=2 l=0.15 M=2
X15 VDD a_629_182 a_1105_1004 VDD pshort w=2 l=0.15 M=2
X16 GND a_185_182 a_2110_73 GND nshort w=3 l=0.15
X17 a_629_182 D GND GND nshort w=3 l=0.15
X18 a_2849_182 a_2215_1004 GND GND nshort w=3 l=0.15
X19 a_1105_1004 a_185_182 a_1000_73 GND nshort w=3 l=0.15
X20 a_3451_383 Q GND GND nshort w=3 l=0.15
X21 Q a_1739_182 GND GND nshort w=3 l=0.15
X22 a_3451_383 a_2849_182 GND GND nshort w=3 l=0.15
X23 a_2215_1004 D a_2110_73 GND nshort w=3 l=0.15
C0 VDD GND 10.87fF
.ends
