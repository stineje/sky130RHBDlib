** sch_path: /home/rjridle/OpenRadHardSCL/lib/xschem/Tutorial/Timing_Specifications.sch
**.subckt Timing_Specifications
**.ends
.end
