* SPICE3 file created from NAND3X1.ext - technology: sky130A

.subckt NAND3X1 Y A B VDD VSS
X0 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=0.00226 pd=1.826 as=0.00174 ps=1.374 w=2 l=0.15 M=2
X1 VDD a_599_989 Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X2 Y a_599_989 a_372_210 VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0 ps=0 w=3 l=0.15
X3 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X4 VSS A a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0 ps=0 w=3 l=0.15
X5 a_372_210 B a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
C0 VDD Y 2.50f
.ends
