magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -66 377 3618 897
<< pwell >>
rect 4 43 3538 317
rect -26 -43 3578 43
<< locali >>
rect 44 316 926 363
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3552 831
rect 22 729 136 751
rect 22 695 30 729
rect 64 695 102 729
rect 22 435 136 695
rect 170 453 232 751
rect 268 729 446 735
rect 302 695 340 729
rect 374 695 412 729
rect 268 489 446 695
rect 480 453 542 751
rect 576 729 754 735
rect 610 695 648 729
rect 682 695 720 729
rect 576 489 754 695
rect 788 453 858 751
rect 892 729 1070 735
rect 926 695 964 729
rect 998 695 1036 729
rect 892 489 1070 695
rect 1114 498 1180 751
rect 1114 464 1130 498
rect 1164 464 1180 498
rect 170 397 1070 453
rect 960 282 1070 397
rect 22 119 129 282
rect 163 239 1070 282
rect 163 151 234 239
rect 22 85 23 119
rect 57 85 95 119
rect 268 119 446 205
rect 480 146 558 239
rect 302 85 340 119
rect 374 85 412 119
rect 592 119 771 205
rect 805 146 854 239
rect 592 85 664 119
rect 698 85 736 119
rect 770 85 771 119
rect 888 119 1066 205
rect 1114 158 1180 464
rect 1214 729 1392 751
rect 1248 695 1286 729
rect 1320 695 1358 729
rect 1214 435 1392 695
rect 1426 498 1492 751
rect 1426 464 1442 498
rect 1476 464 1492 498
rect 1232 313 1366 379
rect 888 85 960 119
rect 994 85 1032 119
rect 1214 119 1392 279
rect 1426 158 1492 464
rect 1526 729 1704 751
rect 1560 695 1598 729
rect 1632 695 1670 729
rect 1526 435 1704 695
rect 1738 498 1804 751
rect 1738 464 1754 498
rect 1788 464 1804 498
rect 1544 313 1678 379
rect 1214 85 1286 119
rect 1320 85 1358 119
rect 1526 119 1704 279
rect 1738 158 1804 464
rect 1838 729 2016 751
rect 1872 695 1910 729
rect 1944 695 1982 729
rect 1838 435 2016 695
rect 2050 498 2116 751
rect 2050 464 2066 498
rect 2100 464 2116 498
rect 1856 313 1990 379
rect 1526 85 1598 119
rect 1632 85 1670 119
rect 1838 119 2016 279
rect 2050 158 2116 464
rect 2150 729 2328 751
rect 2184 695 2222 729
rect 2256 695 2294 729
rect 2150 435 2328 695
rect 2362 498 2428 751
rect 2362 464 2378 498
rect 2412 464 2428 498
rect 2168 313 2302 379
rect 1838 85 1910 119
rect 1944 85 1982 119
rect 2150 119 2328 279
rect 2362 158 2428 464
rect 2462 729 2640 751
rect 2496 695 2534 729
rect 2568 695 2606 729
rect 2462 435 2640 695
rect 2674 498 2740 751
rect 2674 464 2690 498
rect 2724 464 2740 498
rect 2480 313 2614 379
rect 2150 85 2222 119
rect 2256 85 2294 119
rect 2462 119 2640 279
rect 2674 158 2740 464
rect 2774 729 2952 751
rect 2808 695 2846 729
rect 2880 695 2918 729
rect 2774 435 2952 695
rect 2986 498 3052 751
rect 2986 464 3002 498
rect 3036 464 3052 498
rect 2792 313 2926 379
rect 2462 85 2534 119
rect 2568 85 2606 119
rect 2774 119 2952 279
rect 2986 158 3052 464
rect 3086 729 3264 751
rect 3120 695 3158 729
rect 3192 695 3230 729
rect 3086 435 3264 695
rect 3298 498 3380 751
rect 3298 464 3314 498
rect 3348 464 3380 498
rect 3104 313 3238 379
rect 2774 85 2846 119
rect 2880 85 2918 119
rect 3086 119 3264 279
rect 3298 158 3380 464
rect 3414 729 3520 751
rect 3448 695 3486 729
rect 3414 435 3520 695
rect 3086 85 3158 119
rect 3192 85 3230 119
rect 3414 119 3520 299
rect 3414 85 3486 119
rect 268 83 446 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 30 695 64 729
rect 102 695 136 729
rect 268 695 302 729
rect 340 695 374 729
rect 412 695 446 729
rect 576 695 610 729
rect 648 695 682 729
rect 720 695 754 729
rect 892 695 926 729
rect 964 695 998 729
rect 1036 695 1070 729
rect 1130 464 1164 498
rect 23 85 57 119
rect 95 85 129 119
rect 268 85 302 119
rect 340 85 374 119
rect 412 85 446 119
rect 664 85 698 119
rect 736 85 770 119
rect 1214 695 1248 729
rect 1286 695 1320 729
rect 1358 695 1392 729
rect 1442 464 1476 498
rect 960 85 994 119
rect 1032 85 1066 119
rect 1526 695 1560 729
rect 1598 695 1632 729
rect 1670 695 1704 729
rect 1754 464 1788 498
rect 1286 85 1320 119
rect 1358 85 1392 119
rect 1838 695 1872 729
rect 1910 695 1944 729
rect 1982 695 2016 729
rect 2066 464 2100 498
rect 1598 85 1632 119
rect 1670 85 1704 119
rect 2150 695 2184 729
rect 2222 695 2256 729
rect 2294 695 2328 729
rect 2378 464 2412 498
rect 1910 85 1944 119
rect 1982 85 2016 119
rect 2462 695 2496 729
rect 2534 695 2568 729
rect 2606 695 2640 729
rect 2690 464 2724 498
rect 2222 85 2256 119
rect 2294 85 2328 119
rect 2774 695 2808 729
rect 2846 695 2880 729
rect 2918 695 2952 729
rect 3002 464 3036 498
rect 2534 85 2568 119
rect 2606 85 2640 119
rect 3086 695 3120 729
rect 3158 695 3192 729
rect 3230 695 3264 729
rect 3314 464 3348 498
rect 2846 85 2880 119
rect 2918 85 2952 119
rect 3414 695 3448 729
rect 3486 695 3520 729
rect 3158 85 3192 119
rect 3230 85 3264 119
rect 3486 85 3520 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
<< metal1 >>
rect 0 831 3552 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3552 831
rect 0 791 3552 797
rect 0 729 3552 763
rect 0 695 30 729
rect 64 695 102 729
rect 136 695 268 729
rect 302 695 340 729
rect 374 695 412 729
rect 446 695 576 729
rect 610 695 648 729
rect 682 695 720 729
rect 754 695 892 729
rect 926 695 964 729
rect 998 695 1036 729
rect 1070 695 1214 729
rect 1248 695 1286 729
rect 1320 695 1358 729
rect 1392 695 1526 729
rect 1560 695 1598 729
rect 1632 695 1670 729
rect 1704 695 1838 729
rect 1872 695 1910 729
rect 1944 695 1982 729
rect 2016 695 2150 729
rect 2184 695 2222 729
rect 2256 695 2294 729
rect 2328 695 2462 729
rect 2496 695 2534 729
rect 2568 695 2606 729
rect 2640 695 2774 729
rect 2808 695 2846 729
rect 2880 695 2918 729
rect 2952 695 3086 729
rect 3120 695 3158 729
rect 3192 695 3230 729
rect 3264 695 3414 729
rect 3448 695 3486 729
rect 3520 695 3552 729
rect 0 689 3552 695
rect 1118 498 1176 504
rect 1430 498 1488 504
rect 1742 498 1800 504
rect 2054 498 2112 504
rect 2366 498 2424 504
rect 2678 498 2736 504
rect 2990 498 3048 504
rect 3302 498 3360 504
rect 1118 464 1130 498
rect 1164 464 1442 498
rect 1476 464 1754 498
rect 1788 464 2066 498
rect 2100 464 2378 498
rect 2412 464 2690 498
rect 2724 464 3002 498
rect 3036 464 3314 498
rect 3348 464 3360 498
rect 1118 458 1176 464
rect 1430 458 1488 464
rect 1742 458 1800 464
rect 2054 458 2112 464
rect 2366 458 2424 464
rect 2678 458 2736 464
rect 2990 458 3048 464
rect 3302 458 3360 464
rect 0 119 3552 125
rect 0 85 23 119
rect 57 85 95 119
rect 129 85 268 119
rect 302 85 340 119
rect 374 85 412 119
rect 446 85 664 119
rect 698 85 736 119
rect 770 85 960 119
rect 994 85 1032 119
rect 1066 85 1286 119
rect 1320 85 1358 119
rect 1392 85 1598 119
rect 1632 85 1670 119
rect 1704 85 1910 119
rect 1944 85 1982 119
rect 2016 85 2222 119
rect 2256 85 2294 119
rect 2328 85 2534 119
rect 2568 85 2606 119
rect 2640 85 2846 119
rect 2880 85 2918 119
rect 2952 85 3158 119
rect 3192 85 3230 119
rect 3264 85 3486 119
rect 3520 85 3552 119
rect 0 51 3552 85
rect 0 17 3552 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3552 17
rect 0 -23 3552 -17
<< obsm1 >>
rect 948 350 1072 356
rect 1234 350 1364 356
rect 1546 350 1676 356
rect 1858 350 1988 356
rect 2170 350 2300 356
rect 2482 350 2612 356
rect 2794 350 2924 356
rect 3106 350 3236 356
rect 948 316 3250 350
rect 948 310 1072 316
rect 1234 310 1364 316
rect 1546 310 1676 316
rect 1858 310 1988 316
rect 2170 310 2300 316
rect 2482 310 2612 316
rect 2794 310 2924 316
rect 3106 310 3236 316
<< labels >>
rlabel locali s 44 316 926 363 6 A
port 1 nsew signal input
rlabel metal1 s 0 51 3552 125 6 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 -23 3552 23 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s -26 -43 3578 43 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 4 43 3538 317 6 VNB
port 3 nsew ground bidirectional
rlabel metal1 s 0 791 3552 837 6 VPB
port 4 nsew power bidirectional
rlabel nwell s -66 377 3618 897 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 689 3552 763 6 VPWR
port 5 nsew power bidirectional
rlabel metal1 s 3302 458 3360 464 6 X
port 6 nsew signal output
rlabel metal1 s 2990 458 3048 464 6 X
port 6 nsew signal output
rlabel metal1 s 2678 458 2736 464 6 X
port 6 nsew signal output
rlabel metal1 s 2366 458 2424 464 6 X
port 6 nsew signal output
rlabel metal1 s 2054 458 2112 464 6 X
port 6 nsew signal output
rlabel metal1 s 1742 458 1800 464 6 X
port 6 nsew signal output
rlabel metal1 s 1430 458 1488 464 6 X
port 6 nsew signal output
rlabel metal1 s 1118 458 1176 464 6 X
port 6 nsew signal output
rlabel metal1 s 1118 464 3360 498 6 X
port 6 nsew signal output
rlabel metal1 s 3302 498 3360 504 6 X
port 6 nsew signal output
rlabel metal1 s 2990 498 3048 504 6 X
port 6 nsew signal output
rlabel metal1 s 2678 498 2736 504 6 X
port 6 nsew signal output
rlabel metal1 s 2366 498 2424 504 6 X
port 6 nsew signal output
rlabel metal1 s 2054 498 2112 504 6 X
port 6 nsew signal output
rlabel metal1 s 1742 498 1800 504 6 X
port 6 nsew signal output
rlabel metal1 s 1430 498 1488 504 6 X
port 6 nsew signal output
rlabel metal1 s 1118 498 1176 504 6 X
port 6 nsew signal output
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 3552 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 1130684
string GDS_START 1091408
<< end >>
