* SPICE3 file created from AOAI4X1.ext - technology: sky130A

.subckt AOAI4X1 YN A B C D VDD GND
X0 VDD aoai4x1_pcell_0/m1_537_501# aoai4x1_pcell_0/nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X1 aoai4x1_pcell_0/m1_1203_501# C aoai4x1_pcell_0/nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X2 aoai4x1_pcell_0/m1_1203_501# aoai4x1_pcell_0/m1_537_501# GND GND nshort w=3 l=0.15
X3 aoai4x1_pcell_0/m1_1203_501# C GND GND nshort w=3 l=0.15
X4 GND A aoai4x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X5 aoai4x1_pcell_0/m1_537_501# B aoai4x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X6 VDD A aoai4x1_pcell_0/m1_537_501# VDD pshort w=2 l=0.15
X7 VDD B aoai4x1_pcell_0/m1_537_501# VDD pshort w=2 l=0.15
X8 GND aoai4x1_pcell_0/m1_1203_501# aoai4x1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X9 YN D aoai4x1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X10 VDD aoai4x1_pcell_0/m1_1203_501# YN VDD pshort w=2 l=0.15
X11 VDD D YN VDD pshort w=2 l=0.15
C0 VDD GND 4.00fF
.ends
