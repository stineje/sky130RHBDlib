// File: dffx1_pcell.spi.DFFX1_PCELL.pxi
// Created: Tue Oct 15 15:56:33 2024
// 
simulator lang=spectre
x_PM_DFFX1_PCELL\%noxref_1 ( N_noxref_1_c_8_p N_noxref_1_c_97_p \
 N_noxref_1_c_1_p N_noxref_1_c_9_p N_noxref_1_c_10_p N_noxref_1_c_11_p \
 N_noxref_1_c_16_p N_noxref_1_c_30_p N_noxref_1_c_38_p N_noxref_1_c_51_p \
 N_noxref_1_c_75_p N_noxref_1_c_82_p N_noxref_1_c_226_p N_noxref_1_c_2_p \
 N_noxref_1_c_3_p N_noxref_1_c_4_p N_noxref_1_c_5_p N_noxref_1_c_6_p \
 N_noxref_1_c_7_p N_noxref_1_M0_noxref_d N_noxref_1_M3_noxref_d \
 N_noxref_1_M5_noxref_d N_noxref_1_M7_noxref_d N_noxref_1_M9_noxref_d \
 N_noxref_1_M11_noxref_d )  PM_DFFX1_PCELL\%noxref_1
x_PM_DFFX1_PCELL\%noxref_2 ( N_noxref_2_c_266_p N_noxref_2_c_258_n \
 N_noxref_2_c_366_p N_noxref_2_c_355_p N_noxref_2_c_281_p N_noxref_2_c_333_p \
 N_noxref_2_c_334_p N_noxref_2_c_267_p N_noxref_2_c_268_p N_noxref_2_c_336_p \
 N_noxref_2_c_337_p N_noxref_2_c_279_p N_noxref_2_c_303_p N_noxref_2_c_339_p \
 N_noxref_2_c_340_p N_noxref_2_c_314_p N_noxref_2_c_359_p N_noxref_2_c_421_p \
 N_noxref_2_c_422_p N_noxref_2_c_384_p N_noxref_2_c_490_p N_noxref_2_c_424_p \
 N_noxref_2_c_425_p N_noxref_2_c_426_p N_noxref_2_c_463_p N_noxref_2_c_259_n \
 N_noxref_2_c_260_n N_noxref_2_c_261_n N_noxref_2_c_262_n N_noxref_2_c_263_n \
 N_noxref_2_c_264_n N_noxref_2_M13_noxref_s N_noxref_2_M14_noxref_d \
 N_noxref_2_M16_noxref_d N_noxref_2_M18_noxref_d N_noxref_2_M19_noxref_s \
 N_noxref_2_M20_noxref_d N_noxref_2_M22_noxref_d N_noxref_2_M23_noxref_s \
 N_noxref_2_M24_noxref_d N_noxref_2_M26_noxref_d N_noxref_2_M27_noxref_s \
 N_noxref_2_M28_noxref_d N_noxref_2_M30_noxref_d N_noxref_2_M31_noxref_s \
 N_noxref_2_M32_noxref_d N_noxref_2_M34_noxref_d N_noxref_2_M35_noxref_s \
 N_noxref_2_M36_noxref_d N_noxref_2_M38_noxref_d )  PM_DFFX1_PCELL\%noxref_2
x_PM_DFFX1_PCELL\%noxref_3 ( N_noxref_3_c_547_n N_noxref_3_c_552_n \
 N_noxref_3_c_553_n N_noxref_3_c_557_n N_noxref_3_c_558_n N_noxref_3_c_576_n \
 N_noxref_3_c_580_n N_noxref_3_c_582_n N_noxref_3_c_559_n N_noxref_3_c_756_p \
 N_noxref_3_c_560_n N_noxref_3_c_561_n N_noxref_3_c_743_p \
 N_noxref_3_M2_noxref_g N_noxref_3_M5_noxref_g N_noxref_3_M17_noxref_g \
 N_noxref_3_M18_noxref_g N_noxref_3_M23_noxref_g N_noxref_3_M24_noxref_g \
 N_noxref_3_c_636_p N_noxref_3_c_637_p N_noxref_3_c_638_p N_noxref_3_c_680_p \
 N_noxref_3_c_657_p N_noxref_3_c_682_p N_noxref_3_c_658_p N_noxref_3_c_562_n \
 N_noxref_3_c_564_n N_noxref_3_c_565_n N_noxref_3_c_566_n N_noxref_3_c_567_n \
 N_noxref_3_c_568_n N_noxref_3_c_569_n N_noxref_3_c_571_n N_noxref_3_c_631_p \
 N_noxref_3_c_641_p N_noxref_3_c_626_p N_noxref_3_c_599_n \
 N_noxref_3_M4_noxref_d N_noxref_3_M19_noxref_d N_noxref_3_M21_noxref_d )  \
 PM_DFFX1_PCELL\%noxref_3
x_PM_DFFX1_PCELL\%noxref_4 ( N_noxref_4_c_779_n N_noxref_4_c_783_n \
 N_noxref_4_c_800_n N_noxref_4_c_804_n N_noxref_4_c_806_n N_noxref_4_c_784_n \
 N_noxref_4_c_869_p N_noxref_4_c_785_n N_noxref_4_c_786_n N_noxref_4_c_896_p \
 N_noxref_4_M7_noxref_g N_noxref_4_M27_noxref_g N_noxref_4_M28_noxref_g \
 N_noxref_4_c_787_n N_noxref_4_c_789_n N_noxref_4_c_790_n N_noxref_4_c_791_n \
 N_noxref_4_c_792_n N_noxref_4_c_793_n N_noxref_4_c_794_n N_noxref_4_c_796_n \
 N_noxref_4_c_819_n N_noxref_4_M6_noxref_d N_noxref_4_M23_noxref_d \
 N_noxref_4_M25_noxref_d )  PM_DFFX1_PCELL\%noxref_4
x_PM_DFFX1_PCELL\%noxref_5 ( N_noxref_5_c_932_n N_noxref_5_c_950_n \
 N_noxref_5_c_929_n N_noxref_5_c_995_n N_noxref_5_c_930_n \
 N_noxref_5_M1_noxref_g N_noxref_5_M8_noxref_g N_noxref_5_M15_noxref_g \
 N_noxref_5_M16_noxref_g N_noxref_5_M29_noxref_g N_noxref_5_M30_noxref_g \
 N_noxref_5_c_1075_p N_noxref_5_c_1077_p N_noxref_5_c_1109_p \
 N_noxref_5_c_1116_p N_noxref_5_c_981_n N_noxref_5_c_982_n N_noxref_5_c_983_n \
 N_noxref_5_c_984_n N_noxref_5_c_987_n N_noxref_5_c_1004_n N_noxref_5_c_1007_n \
 N_noxref_5_c_1009_n N_noxref_5_c_1045_p N_noxref_5_c_1094_p \
 N_noxref_5_c_1062_p N_noxref_5_c_1012_n N_noxref_5_c_1013_n \
 N_noxref_5_c_988_n N_noxref_5_c_1014_n N_noxref_5_c_1069_p \
 N_noxref_5_c_1016_n )  PM_DFFX1_PCELL\%noxref_5
x_PM_DFFX1_PCELL\%noxref_6 ( N_noxref_6_c_1207_n N_noxref_6_c_1208_n \
 N_noxref_6_c_1134_n N_noxref_6_c_1215_n N_noxref_6_c_1161_n \
 N_noxref_6_c_1165_n N_noxref_6_c_1167_n N_noxref_6_c_1171_n \
 N_noxref_6_c_1136_n N_noxref_6_c_1221_n N_noxref_6_c_1175_n \
 N_noxref_6_c_1137_n N_noxref_6_c_1138_n N_noxref_6_c_1269_n \
 N_noxref_6_c_1233_n N_noxref_6_M3_noxref_g N_noxref_6_M9_noxref_g \
 N_noxref_6_M19_noxref_g N_noxref_6_M20_noxref_g N_noxref_6_M31_noxref_g \
 N_noxref_6_M32_noxref_g N_noxref_6_c_1139_n N_noxref_6_c_1141_n \
 N_noxref_6_c_1142_n N_noxref_6_c_1143_n N_noxref_6_c_1144_n \
 N_noxref_6_c_1145_n N_noxref_6_c_1146_n N_noxref_6_c_1148_n \
 N_noxref_6_c_1149_n N_noxref_6_c_1151_n N_noxref_6_c_1152_n \
 N_noxref_6_c_1153_n N_noxref_6_c_1154_n N_noxref_6_c_1155_n \
 N_noxref_6_c_1156_n N_noxref_6_c_1158_n N_noxref_6_c_1190_n \
 N_noxref_6_c_1191_n N_noxref_6_M2_noxref_d N_noxref_6_M13_noxref_d \
 N_noxref_6_M15_noxref_d N_noxref_6_M17_noxref_d )  PM_DFFX1_PCELL\%noxref_6
x_PM_DFFX1_PCELL\%noxref_7 ( N_noxref_7_c_1385_n N_noxref_7_c_1386_n \
 N_noxref_7_c_1416_n N_noxref_7_c_1486_n N_noxref_7_c_1387_n \
 N_noxref_7_c_1430_n N_noxref_7_c_1389_n N_noxref_7_c_1488_n \
 N_noxref_7_c_1390_n N_noxref_7_c_1438_n N_noxref_7_c_1442_n \
 N_noxref_7_c_1444_n N_noxref_7_c_1392_n N_noxref_7_c_1626_n \
 N_noxref_7_c_1393_n N_noxref_7_c_1681_p N_noxref_7_c_1394_n \
 N_noxref_7_c_1581_n N_noxref_7_M0_noxref_g N_noxref_7_M6_noxref_g \
 N_noxref_7_M12_noxref_g N_noxref_7_M13_noxref_g N_noxref_7_M14_noxref_g \
 N_noxref_7_M25_noxref_g N_noxref_7_M26_noxref_g N_noxref_7_M37_noxref_g \
 N_noxref_7_M38_noxref_g N_noxref_7_c_1396_n N_noxref_7_c_1398_n \
 N_noxref_7_c_1399_n N_noxref_7_c_1400_n N_noxref_7_c_1401_n \
 N_noxref_7_c_1402_n N_noxref_7_c_1403_n N_noxref_7_c_1405_n \
 N_noxref_7_c_1595_n N_noxref_7_c_1466_n N_noxref_7_c_1497_n \
 N_noxref_7_c_1500_n N_noxref_7_c_1502_n N_noxref_7_c_1534_n \
 N_noxref_7_c_1536_n N_noxref_7_c_1537_n N_noxref_7_c_1505_n \
 N_noxref_7_c_1506_n N_noxref_7_c_1688_p N_noxref_7_c_1690_p \
 N_noxref_7_c_1691_p N_noxref_7_c_1714_p N_noxref_7_c_1722_p \
 N_noxref_7_c_1709_p N_noxref_7_c_1696_p N_noxref_7_c_1699_p \
 N_noxref_7_c_1507_n N_noxref_7_c_1543_n N_noxref_7_c_1509_n \
 N_noxref_7_c_1683_p N_noxref_7_c_1716_p N_noxref_7_c_1684_p \
 N_noxref_7_M8_noxref_d N_noxref_7_M27_noxref_d N_noxref_7_M29_noxref_d )  \
 PM_DFFX1_PCELL\%noxref_7
x_PM_DFFX1_PCELL\%noxref_8 ( N_noxref_8_c_1766_n N_noxref_8_c_1741_n \
 N_noxref_8_c_1745_n N_noxref_8_c_1748_n N_noxref_8_c_1759_n \
 N_noxref_8_M0_noxref_s )  PM_DFFX1_PCELL\%noxref_8
x_PM_DFFX1_PCELL\%noxref_9 ( N_noxref_9_c_1788_n N_noxref_9_c_1790_n \
 N_noxref_9_c_1793_n N_noxref_9_c_1796_n N_noxref_9_c_1807_n \
 N_noxref_9_M1_noxref_d N_noxref_9_M2_noxref_s )  PM_DFFX1_PCELL\%noxref_9
x_PM_DFFX1_PCELL\%noxref_10 ( N_noxref_10_c_1850_n N_noxref_10_c_1841_n \
 N_noxref_10_M4_noxref_g N_noxref_10_M21_noxref_g N_noxref_10_M22_noxref_g \
 N_noxref_10_c_1860_n N_noxref_10_c_1861_n N_noxref_10_c_1862_n \
 N_noxref_10_c_1863_n N_noxref_10_c_1865_n N_noxref_10_c_1866_n \
 N_noxref_10_c_1868_n N_noxref_10_c_1869_n N_noxref_10_c_1871_n \
 N_noxref_10_c_1872_n N_noxref_10_c_1874_n )  PM_DFFX1_PCELL\%noxref_10
x_PM_DFFX1_PCELL\%noxref_11 ( N_noxref_11_c_1933_n N_noxref_11_c_1914_n \
 N_noxref_11_c_1918_n N_noxref_11_c_1921_n N_noxref_11_c_1922_n \
 N_noxref_11_c_1925_n N_noxref_11_M3_noxref_s )  PM_DFFX1_PCELL\%noxref_11
x_PM_DFFX1_PCELL\%noxref_12 ( N_noxref_12_c_1985_n N_noxref_12_c_1966_n \
 N_noxref_12_c_1970_n N_noxref_12_c_1973_n N_noxref_12_c_1974_n \
 N_noxref_12_c_1977_n N_noxref_12_M5_noxref_s )  PM_DFFX1_PCELL\%noxref_12
x_PM_DFFX1_PCELL\%noxref_13 ( N_noxref_13_c_2038_n N_noxref_13_c_2019_n \
 N_noxref_13_c_2023_n N_noxref_13_c_2026_n N_noxref_13_c_2027_n \
 N_noxref_13_c_2030_n N_noxref_13_M7_noxref_s )  PM_DFFX1_PCELL\%noxref_13
x_PM_DFFX1_PCELL\%noxref_14 ( N_noxref_14_c_2081_n N_noxref_14_c_2072_n \
 N_noxref_14_M10_noxref_g N_noxref_14_M33_noxref_g N_noxref_14_M34_noxref_g \
 N_noxref_14_c_2089_n N_noxref_14_c_2092_n N_noxref_14_c_2094_n \
 N_noxref_14_c_2106_n N_noxref_14_c_2124_p N_noxref_14_c_2112_p \
 N_noxref_14_c_2097_n N_noxref_14_c_2098_n N_noxref_14_c_2099_n \
 N_noxref_14_c_2118_p N_noxref_14_c_2101_n )  PM_DFFX1_PCELL\%noxref_14
x_PM_DFFX1_PCELL\%noxref_15 ( N_noxref_15_c_2146_n N_noxref_15_c_2150_n \
 N_noxref_15_c_2152_n N_noxref_15_c_2141_n N_noxref_15_c_2177_n \
 N_noxref_15_c_2142_n N_noxref_15_c_2193_n N_noxref_15_M10_noxref_d \
 N_noxref_15_M31_noxref_d N_noxref_15_M33_noxref_d )  PM_DFFX1_PCELL\%noxref_15
x_PM_DFFX1_PCELL\%noxref_16 ( N_noxref_16_c_2232_n N_noxref_16_c_2213_n \
 N_noxref_16_c_2217_n N_noxref_16_c_2220_n N_noxref_16_c_2221_n \
 N_noxref_16_c_2224_n N_noxref_16_M9_noxref_s )  PM_DFFX1_PCELL\%noxref_16
x_PM_DFFX1_PCELL\%noxref_17 ( N_noxref_17_c_2265_n N_noxref_17_M11_noxref_g \
 N_noxref_17_M35_noxref_g N_noxref_17_M36_noxref_g N_noxref_17_c_2266_n \
 N_noxref_17_c_2268_n N_noxref_17_c_2269_n N_noxref_17_c_2270_n \
 N_noxref_17_c_2271_n N_noxref_17_c_2272_n N_noxref_17_c_2273_n \
 N_noxref_17_c_2275_n N_noxref_17_c_2283_n )  PM_DFFX1_PCELL\%noxref_17
x_PM_DFFX1_PCELL\%noxref_18 ( N_noxref_18_c_2330_n N_noxref_18_c_2334_n \
 N_noxref_18_c_2336_n N_noxref_18_c_2325_n N_noxref_18_c_2384_p \
 N_noxref_18_c_2326_n N_noxref_18_c_2366_n N_noxref_18_M12_noxref_d \
 N_noxref_18_M35_noxref_d N_noxref_18_M37_noxref_d )  PM_DFFX1_PCELL\%noxref_18
x_PM_DFFX1_PCELL\%noxref_19 ( N_noxref_19_c_2407_n N_noxref_19_c_2390_n \
 N_noxref_19_c_2394_n N_noxref_19_c_2397_n N_noxref_19_c_2398_n \
 N_noxref_19_c_2400_n N_noxref_19_M11_noxref_s )  PM_DFFX1_PCELL\%noxref_19
cc_1 ( N_noxref_1_c_1_p N_noxref_2_c_258_n ) capacitor c=0.00989031f //x=0.74 \
 //y=0 //x2=0.74 //y2=7.4
cc_2 ( N_noxref_1_c_2_p N_noxref_2_c_259_n ) capacitor c=0.00989031f //x=21.09 \
 //y=0 //x2=21.09 //y2=7.4
cc_3 ( N_noxref_1_c_3_p N_noxref_2_c_260_n ) capacitor c=0.00500587f //x=4.81 \
 //y=0 //x2=4.81 //y2=7.4
cc_4 ( N_noxref_1_c_4_p N_noxref_2_c_261_n ) capacitor c=0.00500587f //x=8.14 \
 //y=0 //x2=8.14 //y2=7.4
cc_5 ( N_noxref_1_c_5_p N_noxref_2_c_262_n ) capacitor c=0.00500587f //x=11.47 \
 //y=0 //x2=11.47 //y2=7.4
cc_6 ( N_noxref_1_c_6_p N_noxref_2_c_263_n ) capacitor c=0.00524516f //x=14.8 \
 //y=0 //x2=14.8 //y2=7.4
cc_7 ( N_noxref_1_c_7_p N_noxref_2_c_264_n ) capacitor c=0.0052832f //x=18.13 \
 //y=0 //x2=18.13 //y2=7.4
cc_8 ( N_noxref_1_c_8_p N_noxref_3_c_547_n ) capacitor c=0.0264756f //x=21.09 \
 //y=0 //x2=7.285 //y2=3.33
cc_9 ( N_noxref_1_c_9_p N_noxref_3_c_547_n ) capacitor c=0.00174514f //x=4.64 \
 //y=0 //x2=7.285 //y2=3.33
cc_10 ( N_noxref_1_c_10_p N_noxref_3_c_547_n ) capacitor c=0.00192599f \
 //x=5.905 //y=0 //x2=7.285 //y2=3.33
cc_11 ( N_noxref_1_c_11_p N_noxref_3_c_547_n ) capacitor c=5.39691e-19 \
 //x=7.97 //y=0 //x2=7.285 //y2=3.33
cc_12 ( N_noxref_1_c_3_p N_noxref_3_c_547_n ) capacitor c=0.00820844f //x=4.81 \
 //y=0 //x2=7.285 //y2=3.33
cc_13 ( N_noxref_1_c_8_p N_noxref_3_c_552_n ) capacitor c=0.00172266f \
 //x=21.09 //y=0 //x2=3.445 //y2=3.33
cc_14 ( N_noxref_1_c_8_p N_noxref_3_c_553_n ) capacitor c=0.0143714f //x=21.09 \
 //y=0 //x2=9.135 //y2=3.33
cc_15 ( N_noxref_1_c_11_p N_noxref_3_c_553_n ) capacitor c=0.00157139f \
 //x=7.97 //y=0 //x2=9.135 //y2=3.33
cc_16 ( N_noxref_1_c_16_p N_noxref_3_c_553_n ) capacitor c=0.00189853f \
 //x=9.235 //y=0 //x2=9.135 //y2=3.33
cc_17 ( N_noxref_1_c_4_p N_noxref_3_c_553_n ) capacitor c=0.00820844f //x=8.14 \
 //y=0 //x2=9.135 //y2=3.33
cc_18 ( N_noxref_1_c_8_p N_noxref_3_c_557_n ) capacitor c=0.00153258f \
 //x=21.09 //y=0 //x2=7.515 //y2=3.33
cc_19 ( N_noxref_1_c_3_p N_noxref_3_c_558_n ) capacitor c=9.53263e-19 //x=4.81 \
 //y=0 //x2=3.33 //y2=2.08
cc_20 ( N_noxref_1_c_4_p N_noxref_3_c_559_n ) capacitor c=0.0462817f //x=8.14 \
 //y=0 //x2=7.315 //y2=1.655
cc_21 ( N_noxref_1_c_3_p N_noxref_3_c_560_n ) capacitor c=9.64732e-19 //x=4.81 \
 //y=0 //x2=7.4 //y2=3.33
cc_22 ( N_noxref_1_c_4_p N_noxref_3_c_561_n ) capacitor c=0.0179404f //x=8.14 \
 //y=0 //x2=9.25 //y2=2.08
cc_23 ( N_noxref_1_c_16_p N_noxref_3_c_562_n ) capacitor c=0.00135046f \
 //x=9.235 //y=0 //x2=9.055 //y2=0.865
cc_24 ( N_noxref_1_M5_noxref_d N_noxref_3_c_562_n ) capacitor c=0.00220047f \
 //x=9.13 //y=0.865 //x2=9.055 //y2=0.865
cc_25 ( N_noxref_1_M5_noxref_d N_noxref_3_c_564_n ) capacitor c=0.00255985f \
 //x=9.13 //y=0.865 //x2=9.055 //y2=1.21
cc_26 ( N_noxref_1_c_4_p N_noxref_3_c_565_n ) capacitor c=0.0018059f //x=8.14 \
 //y=0 //x2=9.055 //y2=1.52
cc_27 ( N_noxref_1_c_4_p N_noxref_3_c_566_n ) capacitor c=0.0114883f //x=8.14 \
 //y=0 //x2=9.055 //y2=1.915
cc_28 ( N_noxref_1_M5_noxref_d N_noxref_3_c_567_n ) capacitor c=0.0131326f \
 //x=9.13 //y=0.865 //x2=9.43 //y2=0.71
cc_29 ( N_noxref_1_M5_noxref_d N_noxref_3_c_568_n ) capacitor c=0.00193127f \
 //x=9.13 //y=0.865 //x2=9.43 //y2=1.365
cc_30 ( N_noxref_1_c_30_p N_noxref_3_c_569_n ) capacitor c=0.00130622f \
 //x=11.3 //y=0 //x2=9.585 //y2=0.865
cc_31 ( N_noxref_1_M5_noxref_d N_noxref_3_c_569_n ) capacitor c=0.00257848f \
 //x=9.13 //y=0.865 //x2=9.585 //y2=0.865
cc_32 ( N_noxref_1_M5_noxref_d N_noxref_3_c_571_n ) capacitor c=0.00255985f \
 //x=9.13 //y=0.865 //x2=9.585 //y2=1.21
cc_33 ( N_noxref_1_c_3_p N_noxref_3_M4_noxref_d ) capacitor c=8.58106e-19 \
 //x=4.81 //y=0 //x2=6.77 //y2=0.905
cc_34 ( N_noxref_1_c_4_p N_noxref_3_M4_noxref_d ) capacitor c=0.00616547f \
 //x=8.14 //y=0 //x2=6.77 //y2=0.905
cc_35 ( N_noxref_1_M3_noxref_d N_noxref_3_M4_noxref_d ) capacitor \
 c=0.00143464f //x=5.8 //y=0.865 //x2=6.77 //y2=0.905
cc_36 ( N_noxref_1_c_8_p N_noxref_4_c_779_n ) capacitor c=0.0143714f //x=21.09 \
 //y=0 //x2=12.465 //y2=3.33
cc_37 ( N_noxref_1_c_30_p N_noxref_4_c_779_n ) capacitor c=0.00157139f \
 //x=11.3 //y=0 //x2=12.465 //y2=3.33
cc_38 ( N_noxref_1_c_38_p N_noxref_4_c_779_n ) capacitor c=0.00189853f \
 //x=12.565 //y=0 //x2=12.465 //y2=3.33
cc_39 ( N_noxref_1_c_5_p N_noxref_4_c_779_n ) capacitor c=0.00820844f \
 //x=11.47 //y=0 //x2=12.465 //y2=3.33
cc_40 ( N_noxref_1_c_8_p N_noxref_4_c_783_n ) capacitor c=0.00174211f \
 //x=21.09 //y=0 //x2=10.845 //y2=3.33
cc_41 ( N_noxref_1_c_5_p N_noxref_4_c_784_n ) capacitor c=0.0462817f //x=11.47 \
 //y=0 //x2=10.645 //y2=1.655
cc_42 ( N_noxref_1_c_4_p N_noxref_4_c_785_n ) capacitor c=9.64732e-19 //x=8.14 \
 //y=0 //x2=10.73 //y2=3.33
cc_43 ( N_noxref_1_c_5_p N_noxref_4_c_786_n ) capacitor c=0.0179404f //x=11.47 \
 //y=0 //x2=12.58 //y2=2.08
cc_44 ( N_noxref_1_c_38_p N_noxref_4_c_787_n ) capacitor c=0.00135046f \
 //x=12.565 //y=0 //x2=12.385 //y2=0.865
cc_45 ( N_noxref_1_M7_noxref_d N_noxref_4_c_787_n ) capacitor c=0.00220047f \
 //x=12.46 //y=0.865 //x2=12.385 //y2=0.865
cc_46 ( N_noxref_1_M7_noxref_d N_noxref_4_c_789_n ) capacitor c=0.00255985f \
 //x=12.46 //y=0.865 //x2=12.385 //y2=1.21
cc_47 ( N_noxref_1_c_5_p N_noxref_4_c_790_n ) capacitor c=0.0018059f //x=11.47 \
 //y=0 //x2=12.385 //y2=1.52
cc_48 ( N_noxref_1_c_5_p N_noxref_4_c_791_n ) capacitor c=0.0114883f //x=11.47 \
 //y=0 //x2=12.385 //y2=1.915
cc_49 ( N_noxref_1_M7_noxref_d N_noxref_4_c_792_n ) capacitor c=0.0131326f \
 //x=12.46 //y=0.865 //x2=12.76 //y2=0.71
cc_50 ( N_noxref_1_M7_noxref_d N_noxref_4_c_793_n ) capacitor c=0.00193127f \
 //x=12.46 //y=0.865 //x2=12.76 //y2=1.365
cc_51 ( N_noxref_1_c_51_p N_noxref_4_c_794_n ) capacitor c=0.00130622f \
 //x=14.63 //y=0 //x2=12.915 //y2=0.865
cc_52 ( N_noxref_1_M7_noxref_d N_noxref_4_c_794_n ) capacitor c=0.00257848f \
 //x=12.46 //y=0.865 //x2=12.915 //y2=0.865
cc_53 ( N_noxref_1_M7_noxref_d N_noxref_4_c_796_n ) capacitor c=0.00255985f \
 //x=12.46 //y=0.865 //x2=12.915 //y2=1.21
cc_54 ( N_noxref_1_c_4_p N_noxref_4_M6_noxref_d ) capacitor c=8.58106e-19 \
 //x=8.14 //y=0 //x2=10.1 //y2=0.905
cc_55 ( N_noxref_1_c_5_p N_noxref_4_M6_noxref_d ) capacitor c=0.00616547f \
 //x=11.47 //y=0 //x2=10.1 //y2=0.905
cc_56 ( N_noxref_1_M5_noxref_d N_noxref_4_M6_noxref_d ) capacitor \
 c=0.00143464f //x=9.13 //y=0.865 //x2=10.1 //y2=0.905
cc_57 ( N_noxref_1_c_1_p N_noxref_5_c_929_n ) capacitor c=7.64246e-19 //x=0.74 \
 //y=0 //x2=2.22 //y2=2.08
cc_58 ( N_noxref_1_c_5_p N_noxref_5_c_930_n ) capacitor c=9.2064e-19 //x=11.47 \
 //y=0 //x2=13.32 //y2=2.08
cc_59 ( N_noxref_1_c_6_p N_noxref_5_c_930_n ) capacitor c=9.53263e-19 //x=14.8 \
 //y=0 //x2=13.32 //y2=2.08
cc_60 ( N_noxref_1_c_8_p N_noxref_6_c_1134_n ) capacitor c=0.046817f //x=21.09 \
 //y=0 //x2=15.795 //y2=3.7
cc_61 ( N_noxref_1_c_6_p N_noxref_6_c_1134_n ) capacitor c=0.00533016f \
 //x=14.8 //y=0 //x2=15.795 //y2=3.7
cc_62 ( N_noxref_1_c_3_p N_noxref_6_c_1136_n ) capacitor c=0.0459932f //x=4.81 \
 //y=0 //x2=3.985 //y2=1.665
cc_63 ( N_noxref_1_c_3_p N_noxref_6_c_1137_n ) capacitor c=0.0179404f //x=4.81 \
 //y=0 //x2=5.92 //y2=2.08
cc_64 ( N_noxref_1_c_6_p N_noxref_6_c_1138_n ) capacitor c=0.0179404f //x=14.8 \
 //y=0 //x2=15.91 //y2=2.08
cc_65 ( N_noxref_1_c_10_p N_noxref_6_c_1139_n ) capacitor c=0.00135046f \
 //x=5.905 //y=0 //x2=5.725 //y2=0.865
cc_66 ( N_noxref_1_M3_noxref_d N_noxref_6_c_1139_n ) capacitor c=0.00220047f \
 //x=5.8 //y=0.865 //x2=5.725 //y2=0.865
cc_67 ( N_noxref_1_M3_noxref_d N_noxref_6_c_1141_n ) capacitor c=0.00255985f \
 //x=5.8 //y=0.865 //x2=5.725 //y2=1.21
cc_68 ( N_noxref_1_c_3_p N_noxref_6_c_1142_n ) capacitor c=0.00189421f \
 //x=4.81 //y=0 //x2=5.725 //y2=1.52
cc_69 ( N_noxref_1_c_3_p N_noxref_6_c_1143_n ) capacitor c=0.0114883f //x=4.81 \
 //y=0 //x2=5.725 //y2=1.915
cc_70 ( N_noxref_1_M3_noxref_d N_noxref_6_c_1144_n ) capacitor c=0.0131326f \
 //x=5.8 //y=0.865 //x2=6.1 //y2=0.71
cc_71 ( N_noxref_1_M3_noxref_d N_noxref_6_c_1145_n ) capacitor c=0.00193127f \
 //x=5.8 //y=0.865 //x2=6.1 //y2=1.365
cc_72 ( N_noxref_1_c_11_p N_noxref_6_c_1146_n ) capacitor c=0.00130622f \
 //x=7.97 //y=0 //x2=6.255 //y2=0.865
cc_73 ( N_noxref_1_M3_noxref_d N_noxref_6_c_1146_n ) capacitor c=0.00257848f \
 //x=5.8 //y=0.865 //x2=6.255 //y2=0.865
cc_74 ( N_noxref_1_M3_noxref_d N_noxref_6_c_1148_n ) capacitor c=0.00255985f \
 //x=5.8 //y=0.865 //x2=6.255 //y2=1.21
cc_75 ( N_noxref_1_c_75_p N_noxref_6_c_1149_n ) capacitor c=0.00135046f \
 //x=15.895 //y=0 //x2=15.715 //y2=0.865
cc_76 ( N_noxref_1_M9_noxref_d N_noxref_6_c_1149_n ) capacitor c=0.00220047f \
 //x=15.79 //y=0.865 //x2=15.715 //y2=0.865
cc_77 ( N_noxref_1_M9_noxref_d N_noxref_6_c_1151_n ) capacitor c=0.00255985f \
 //x=15.79 //y=0.865 //x2=15.715 //y2=1.21
cc_78 ( N_noxref_1_c_6_p N_noxref_6_c_1152_n ) capacitor c=0.0018059f //x=14.8 \
 //y=0 //x2=15.715 //y2=1.52
cc_79 ( N_noxref_1_c_6_p N_noxref_6_c_1153_n ) capacitor c=0.0114883f //x=14.8 \
 //y=0 //x2=15.715 //y2=1.915
cc_80 ( N_noxref_1_M9_noxref_d N_noxref_6_c_1154_n ) capacitor c=0.0131326f \
 //x=15.79 //y=0.865 //x2=16.09 //y2=0.71
cc_81 ( N_noxref_1_M9_noxref_d N_noxref_6_c_1155_n ) capacitor c=0.00193127f \
 //x=15.79 //y=0.865 //x2=16.09 //y2=1.365
cc_82 ( N_noxref_1_c_82_p N_noxref_6_c_1156_n ) capacitor c=0.00130622f \
 //x=17.96 //y=0 //x2=16.245 //y2=0.865
cc_83 ( N_noxref_1_M9_noxref_d N_noxref_6_c_1156_n ) capacitor c=0.00257848f \
 //x=15.79 //y=0.865 //x2=16.245 //y2=0.865
cc_84 ( N_noxref_1_M9_noxref_d N_noxref_6_c_1158_n ) capacitor c=0.00255985f \
 //x=15.79 //y=0.865 //x2=16.245 //y2=1.21
cc_85 ( N_noxref_1_c_3_p N_noxref_6_M2_noxref_d ) capacitor c=0.00591582f \
 //x=4.81 //y=0 //x2=3.395 //y2=0.915
cc_86 ( N_noxref_1_c_8_p N_noxref_7_c_1385_n ) capacitor c=0.0147496f \
 //x=21.09 //y=0 //x2=9.875 //y2=4.07
cc_87 ( N_noxref_1_c_8_p N_noxref_7_c_1386_n ) capacitor c=0.0015877f \
 //x=21.09 //y=0 //x2=1.225 //y2=4.07
cc_88 ( N_noxref_1_c_8_p N_noxref_7_c_1387_n ) capacitor c=0.0278143f \
 //x=21.09 //y=0 //x2=19.865 //y2=4.07
cc_89 ( N_noxref_1_c_7_p N_noxref_7_c_1387_n ) capacitor c=0.00363802f \
 //x=18.13 //y=0 //x2=19.865 //y2=4.07
cc_90 ( N_noxref_1_c_1_p N_noxref_7_c_1389_n ) capacitor c=0.0180363f //x=0.74 \
 //y=0 //x2=1.11 //y2=2.08
cc_91 ( N_noxref_1_c_4_p N_noxref_7_c_1390_n ) capacitor c=9.2064e-19 //x=8.14 \
 //y=0 //x2=9.99 //y2=2.08
cc_92 ( N_noxref_1_c_5_p N_noxref_7_c_1390_n ) capacitor c=9.53263e-19 \
 //x=11.47 //y=0 //x2=9.99 //y2=2.08
cc_93 ( N_noxref_1_c_6_p N_noxref_7_c_1392_n ) capacitor c=0.0462817f //x=14.8 \
 //y=0 //x2=13.975 //y2=1.655
cc_94 ( N_noxref_1_c_5_p N_noxref_7_c_1393_n ) capacitor c=9.64732e-19 \
 //x=11.47 //y=0 //x2=14.06 //y2=4.07
cc_95 ( N_noxref_1_c_2_p N_noxref_7_c_1394_n ) capacitor c=9.53263e-19 \
 //x=21.09 //y=0 //x2=19.98 //y2=2.08
cc_96 ( N_noxref_1_c_7_p N_noxref_7_c_1394_n ) capacitor c=9.2064e-19 \
 //x=18.13 //y=0 //x2=19.98 //y2=2.08
cc_97 ( N_noxref_1_c_97_p N_noxref_7_c_1396_n ) capacitor c=0.00132755f \
 //x=0.99 //y=0 //x2=0.81 //y2=0.875
cc_98 ( N_noxref_1_M0_noxref_d N_noxref_7_c_1396_n ) capacitor c=0.00211996f \
 //x=0.885 //y=0.875 //x2=0.81 //y2=0.875
cc_99 ( N_noxref_1_M0_noxref_d N_noxref_7_c_1398_n ) capacitor c=0.00255985f \
 //x=0.885 //y=0.875 //x2=0.81 //y2=1.22
cc_100 ( N_noxref_1_c_1_p N_noxref_7_c_1399_n ) capacitor c=0.00295461f \
 //x=0.74 //y=0 //x2=0.81 //y2=1.53
cc_101 ( N_noxref_1_c_1_p N_noxref_7_c_1400_n ) capacitor c=0.0134214f \
 //x=0.74 //y=0 //x2=0.81 //y2=1.915
cc_102 ( N_noxref_1_M0_noxref_d N_noxref_7_c_1401_n ) capacitor c=0.0131341f \
 //x=0.885 //y=0.875 //x2=1.185 //y2=0.72
cc_103 ( N_noxref_1_M0_noxref_d N_noxref_7_c_1402_n ) capacitor c=0.00193146f \
 //x=0.885 //y=0.875 //x2=1.185 //y2=1.375
cc_104 ( N_noxref_1_c_9_p N_noxref_7_c_1403_n ) capacitor c=0.00129018f \
 //x=4.64 //y=0 //x2=1.34 //y2=0.875
cc_105 ( N_noxref_1_M0_noxref_d N_noxref_7_c_1403_n ) capacitor c=0.00257848f \
 //x=0.885 //y=0.875 //x2=1.34 //y2=0.875
cc_106 ( N_noxref_1_M0_noxref_d N_noxref_7_c_1405_n ) capacitor c=0.00255985f \
 //x=0.885 //y=0.875 //x2=1.34 //y2=1.22
cc_107 ( N_noxref_1_c_5_p N_noxref_7_M8_noxref_d ) capacitor c=8.58106e-19 \
 //x=11.47 //y=0 //x2=13.43 //y2=0.905
cc_108 ( N_noxref_1_c_6_p N_noxref_7_M8_noxref_d ) capacitor c=0.00616547f \
 //x=14.8 //y=0 //x2=13.43 //y2=0.905
cc_109 ( N_noxref_1_M7_noxref_d N_noxref_7_M8_noxref_d ) capacitor \
 c=0.00143464f //x=12.46 //y=0.865 //x2=13.43 //y2=0.905
cc_110 ( N_noxref_1_c_8_p N_noxref_8_c_1741_n ) capacitor c=0.00618812f \
 //x=21.09 //y=0 //x2=1.475 //y2=1.59
cc_111 ( N_noxref_1_c_97_p N_noxref_8_c_1741_n ) capacitor c=0.00110021f \
 //x=0.99 //y=0 //x2=1.475 //y2=1.59
cc_112 ( N_noxref_1_c_9_p N_noxref_8_c_1741_n ) capacitor c=0.00179185f \
 //x=4.64 //y=0 //x2=1.475 //y2=1.59
cc_113 ( N_noxref_1_M0_noxref_d N_noxref_8_c_1741_n ) capacitor c=0.00894788f \
 //x=0.885 //y=0.875 //x2=1.475 //y2=1.59
cc_114 ( N_noxref_1_c_8_p N_noxref_8_c_1745_n ) capacitor c=0.00575184f \
 //x=21.09 //y=0 //x2=1.56 //y2=0.625
cc_115 ( N_noxref_1_c_9_p N_noxref_8_c_1745_n ) capacitor c=0.0140218f \
 //x=4.64 //y=0 //x2=1.56 //y2=0.625
cc_116 ( N_noxref_1_M0_noxref_d N_noxref_8_c_1745_n ) capacitor c=0.033954f \
 //x=0.885 //y=0.875 //x2=1.56 //y2=0.625
cc_117 ( N_noxref_1_c_8_p N_noxref_8_c_1748_n ) capacitor c=0.0139021f \
 //x=21.09 //y=0 //x2=2.445 //y2=0.54
cc_118 ( N_noxref_1_c_9_p N_noxref_8_c_1748_n ) capacitor c=0.0356078f \
 //x=4.64 //y=0 //x2=2.445 //y2=0.54
cc_119 ( N_noxref_1_c_2_p N_noxref_8_c_1748_n ) capacitor c=0.00177725f \
 //x=21.09 //y=0 //x2=2.445 //y2=0.54
cc_120 ( N_noxref_1_c_8_p N_noxref_8_M0_noxref_s ) capacitor c=0.0125336f \
 //x=21.09 //y=0 //x2=0.455 //y2=0.375
cc_121 ( N_noxref_1_c_97_p N_noxref_8_M0_noxref_s ) capacitor c=0.0140218f \
 //x=0.99 //y=0 //x2=0.455 //y2=0.375
cc_122 ( N_noxref_1_c_1_p N_noxref_8_M0_noxref_s ) capacitor c=0.0712607f \
 //x=0.74 //y=0 //x2=0.455 //y2=0.375
cc_123 ( N_noxref_1_c_9_p N_noxref_8_M0_noxref_s ) capacitor c=0.0131422f \
 //x=4.64 //y=0 //x2=0.455 //y2=0.375
cc_124 ( N_noxref_1_c_3_p N_noxref_8_M0_noxref_s ) capacitor c=3.31601e-19 \
 //x=4.81 //y=0 //x2=0.455 //y2=0.375
cc_125 ( N_noxref_1_M0_noxref_d N_noxref_8_M0_noxref_s ) capacitor c=0.033718f \
 //x=0.885 //y=0.875 //x2=0.455 //y2=0.375
cc_126 ( N_noxref_1_c_8_p N_noxref_9_c_1788_n ) capacitor c=0.00402784f \
 //x=21.09 //y=0 //x2=3.015 //y2=0.995
cc_127 ( N_noxref_1_c_9_p N_noxref_9_c_1788_n ) capacitor c=0.00829979f \
 //x=4.64 //y=0 //x2=3.015 //y2=0.995
cc_128 ( N_noxref_1_c_8_p N_noxref_9_c_1790_n ) capacitor c=0.00575184f \
 //x=21.09 //y=0 //x2=3.1 //y2=0.625
cc_129 ( N_noxref_1_c_9_p N_noxref_9_c_1790_n ) capacitor c=0.0140218f \
 //x=4.64 //y=0 //x2=3.1 //y2=0.625
cc_130 ( N_noxref_1_M0_noxref_d N_noxref_9_c_1790_n ) capacitor c=6.21394e-19 \
 //x=0.885 //y=0.875 //x2=3.1 //y2=0.625
cc_131 ( N_noxref_1_c_8_p N_noxref_9_c_1793_n ) capacitor c=0.0118365f \
 //x=21.09 //y=0 //x2=3.985 //y2=0.54
cc_132 ( N_noxref_1_c_9_p N_noxref_9_c_1793_n ) capacitor c=0.0365413f \
 //x=4.64 //y=0 //x2=3.985 //y2=0.54
cc_133 ( N_noxref_1_c_2_p N_noxref_9_c_1793_n ) capacitor c=0.00189848f \
 //x=21.09 //y=0 //x2=3.985 //y2=0.54
cc_134 ( N_noxref_1_c_8_p N_noxref_9_c_1796_n ) capacitor c=0.00287549f \
 //x=21.09 //y=0 //x2=4.07 //y2=0.625
cc_135 ( N_noxref_1_c_9_p N_noxref_9_c_1796_n ) capacitor c=0.0142658f \
 //x=4.64 //y=0 //x2=4.07 //y2=0.625
cc_136 ( N_noxref_1_c_3_p N_noxref_9_c_1796_n ) capacitor c=0.0404137f \
 //x=4.81 //y=0 //x2=4.07 //y2=0.625
cc_137 ( N_noxref_1_M0_noxref_d N_noxref_9_M1_noxref_d ) capacitor \
 c=0.00162435f //x=0.885 //y=0.875 //x2=1.86 //y2=0.91
cc_138 ( N_noxref_1_c_1_p N_noxref_9_M2_noxref_s ) capacitor c=8.16352e-19 \
 //x=0.74 //y=0 //x2=2.965 //y2=0.375
cc_139 ( N_noxref_1_c_3_p N_noxref_9_M2_noxref_s ) capacitor c=0.00183576f \
 //x=4.81 //y=0 //x2=2.965 //y2=0.375
cc_140 ( N_noxref_1_c_3_p N_noxref_10_c_1841_n ) capacitor c=9.2064e-19 \
 //x=4.81 //y=0 //x2=6.66 //y2=2.08
cc_141 ( N_noxref_1_c_4_p N_noxref_10_c_1841_n ) capacitor c=9.53263e-19 \
 //x=8.14 //y=0 //x2=6.66 //y2=2.08
cc_142 ( N_noxref_1_c_8_p N_noxref_11_c_1914_n ) capacitor c=0.00552526f \
 //x=21.09 //y=0 //x2=6.39 //y2=1.58
cc_143 ( N_noxref_1_c_10_p N_noxref_11_c_1914_n ) capacitor c=0.00113001f \
 //x=5.905 //y=0 //x2=6.39 //y2=1.58
cc_144 ( N_noxref_1_c_11_p N_noxref_11_c_1914_n ) capacitor c=0.0018242f \
 //x=7.97 //y=0 //x2=6.39 //y2=1.58
cc_145 ( N_noxref_1_M3_noxref_d N_noxref_11_c_1914_n ) capacitor c=0.00897209f \
 //x=5.8 //y=0.865 //x2=6.39 //y2=1.58
cc_146 ( N_noxref_1_c_8_p N_noxref_11_c_1918_n ) capacitor c=0.00293348f \
 //x=21.09 //y=0 //x2=6.475 //y2=0.615
cc_147 ( N_noxref_1_c_11_p N_noxref_11_c_1918_n ) capacitor c=0.0149357f \
 //x=7.97 //y=0 //x2=6.475 //y2=0.615
cc_148 ( N_noxref_1_M3_noxref_d N_noxref_11_c_1918_n ) capacitor c=0.033812f \
 //x=5.8 //y=0.865 //x2=6.475 //y2=0.615
cc_149 ( N_noxref_1_c_3_p N_noxref_11_c_1921_n ) capacitor c=2.91423e-19 \
 //x=4.81 //y=0 //x2=6.475 //y2=1.495
cc_150 ( N_noxref_1_c_8_p N_noxref_11_c_1922_n ) capacitor c=0.0120397f \
 //x=21.09 //y=0 //x2=7.36 //y2=0.53
cc_151 ( N_noxref_1_c_11_p N_noxref_11_c_1922_n ) capacitor c=0.037553f \
 //x=7.97 //y=0 //x2=7.36 //y2=0.53
cc_152 ( N_noxref_1_c_2_p N_noxref_11_c_1922_n ) capacitor c=0.00198885f \
 //x=21.09 //y=0 //x2=7.36 //y2=0.53
cc_153 ( N_noxref_1_c_8_p N_noxref_11_c_1925_n ) capacitor c=0.00292576f \
 //x=21.09 //y=0 //x2=7.445 //y2=0.615
cc_154 ( N_noxref_1_c_11_p N_noxref_11_c_1925_n ) capacitor c=0.0148673f \
 //x=7.97 //y=0 //x2=7.445 //y2=0.615
cc_155 ( N_noxref_1_c_4_p N_noxref_11_c_1925_n ) capacitor c=0.0431718f \
 //x=8.14 //y=0 //x2=7.445 //y2=0.615
cc_156 ( N_noxref_1_c_8_p N_noxref_11_M3_noxref_s ) capacitor c=0.00293348f \
 //x=21.09 //y=0 //x2=5.37 //y2=0.365
cc_157 ( N_noxref_1_c_10_p N_noxref_11_M3_noxref_s ) capacitor c=0.0149357f \
 //x=5.905 //y=0 //x2=5.37 //y2=0.365
cc_158 ( N_noxref_1_c_3_p N_noxref_11_M3_noxref_s ) capacitor c=0.0583534f \
 //x=4.81 //y=0 //x2=5.37 //y2=0.365
cc_159 ( N_noxref_1_c_4_p N_noxref_11_M3_noxref_s ) capacitor c=0.00198043f \
 //x=8.14 //y=0 //x2=5.37 //y2=0.365
cc_160 ( N_noxref_1_M3_noxref_d N_noxref_11_M3_noxref_s ) capacitor \
 c=0.0334197f //x=5.8 //y=0.865 //x2=5.37 //y2=0.365
cc_161 ( N_noxref_1_c_8_p N_noxref_12_c_1966_n ) capacitor c=0.00556119f \
 //x=21.09 //y=0 //x2=9.72 //y2=1.58
cc_162 ( N_noxref_1_c_16_p N_noxref_12_c_1966_n ) capacitor c=0.00113001f \
 //x=9.235 //y=0 //x2=9.72 //y2=1.58
cc_163 ( N_noxref_1_c_30_p N_noxref_12_c_1966_n ) capacitor c=0.00180846f \
 //x=11.3 //y=0 //x2=9.72 //y2=1.58
cc_164 ( N_noxref_1_M5_noxref_d N_noxref_12_c_1966_n ) capacitor c=0.00897268f \
 //x=9.13 //y=0.865 //x2=9.72 //y2=1.58
cc_165 ( N_noxref_1_c_8_p N_noxref_12_c_1970_n ) capacitor c=0.00302994f \
 //x=21.09 //y=0 //x2=9.805 //y2=0.615
cc_166 ( N_noxref_1_c_30_p N_noxref_12_c_1970_n ) capacitor c=0.0146208f \
 //x=11.3 //y=0 //x2=9.805 //y2=0.615
cc_167 ( N_noxref_1_M5_noxref_d N_noxref_12_c_1970_n ) capacitor c=0.033812f \
 //x=9.13 //y=0.865 //x2=9.805 //y2=0.615
cc_168 ( N_noxref_1_c_4_p N_noxref_12_c_1973_n ) capacitor c=2.91423e-19 \
 //x=8.14 //y=0 //x2=9.805 //y2=1.495
cc_169 ( N_noxref_1_c_8_p N_noxref_12_c_1974_n ) capacitor c=0.0123695f \
 //x=21.09 //y=0 //x2=10.69 //y2=0.53
cc_170 ( N_noxref_1_c_30_p N_noxref_12_c_1974_n ) capacitor c=0.0373121f \
 //x=11.3 //y=0 //x2=10.69 //y2=0.53
cc_171 ( N_noxref_1_c_2_p N_noxref_12_c_1974_n ) capacitor c=0.00198885f \
 //x=21.09 //y=0 //x2=10.69 //y2=0.53
cc_172 ( N_noxref_1_c_8_p N_noxref_12_c_1977_n ) capacitor c=0.00292576f \
 //x=21.09 //y=0 //x2=10.775 //y2=0.615
cc_173 ( N_noxref_1_c_30_p N_noxref_12_c_1977_n ) capacitor c=0.0148673f \
 //x=11.3 //y=0 //x2=10.775 //y2=0.615
cc_174 ( N_noxref_1_c_5_p N_noxref_12_c_1977_n ) capacitor c=0.0431718f \
 //x=11.47 //y=0 //x2=10.775 //y2=0.615
cc_175 ( N_noxref_1_c_8_p N_noxref_12_M5_noxref_s ) capacitor c=0.00293348f \
 //x=21.09 //y=0 //x2=8.7 //y2=0.365
cc_176 ( N_noxref_1_c_16_p N_noxref_12_M5_noxref_s ) capacitor c=0.0149357f \
 //x=9.235 //y=0 //x2=8.7 //y2=0.365
cc_177 ( N_noxref_1_c_4_p N_noxref_12_M5_noxref_s ) capacitor c=0.058339f \
 //x=8.14 //y=0 //x2=8.7 //y2=0.365
cc_178 ( N_noxref_1_c_5_p N_noxref_12_M5_noxref_s ) capacitor c=0.00198043f \
 //x=11.47 //y=0 //x2=8.7 //y2=0.365
cc_179 ( N_noxref_1_M5_noxref_d N_noxref_12_M5_noxref_s ) capacitor \
 c=0.0334197f //x=9.13 //y=0.865 //x2=8.7 //y2=0.365
cc_180 ( N_noxref_1_c_8_p N_noxref_13_c_2019_n ) capacitor c=0.00556119f \
 //x=21.09 //y=0 //x2=13.05 //y2=1.58
cc_181 ( N_noxref_1_c_38_p N_noxref_13_c_2019_n ) capacitor c=0.00113001f \
 //x=12.565 //y=0 //x2=13.05 //y2=1.58
cc_182 ( N_noxref_1_c_51_p N_noxref_13_c_2019_n ) capacitor c=0.00180846f \
 //x=14.63 //y=0 //x2=13.05 //y2=1.58
cc_183 ( N_noxref_1_M7_noxref_d N_noxref_13_c_2019_n ) capacitor c=0.00897268f \
 //x=12.46 //y=0.865 //x2=13.05 //y2=1.58
cc_184 ( N_noxref_1_c_8_p N_noxref_13_c_2023_n ) capacitor c=0.00302994f \
 //x=21.09 //y=0 //x2=13.135 //y2=0.615
cc_185 ( N_noxref_1_c_51_p N_noxref_13_c_2023_n ) capacitor c=0.0146208f \
 //x=14.63 //y=0 //x2=13.135 //y2=0.615
cc_186 ( N_noxref_1_M7_noxref_d N_noxref_13_c_2023_n ) capacitor c=0.033812f \
 //x=12.46 //y=0.865 //x2=13.135 //y2=0.615
cc_187 ( N_noxref_1_c_5_p N_noxref_13_c_2026_n ) capacitor c=2.91423e-19 \
 //x=11.47 //y=0 //x2=13.135 //y2=1.495
cc_188 ( N_noxref_1_c_8_p N_noxref_13_c_2027_n ) capacitor c=0.0124224f \
 //x=21.09 //y=0 //x2=14.02 //y2=0.53
cc_189 ( N_noxref_1_c_51_p N_noxref_13_c_2027_n ) capacitor c=0.0371035f \
 //x=14.63 //y=0 //x2=14.02 //y2=0.53
cc_190 ( N_noxref_1_c_2_p N_noxref_13_c_2027_n ) capacitor c=0.00198885f \
 //x=21.09 //y=0 //x2=14.02 //y2=0.53
cc_191 ( N_noxref_1_c_8_p N_noxref_13_c_2030_n ) capacitor c=0.00303012f \
 //x=21.09 //y=0 //x2=14.105 //y2=0.615
cc_192 ( N_noxref_1_c_51_p N_noxref_13_c_2030_n ) capacitor c=0.0144264f \
 //x=14.63 //y=0 //x2=14.105 //y2=0.615
cc_193 ( N_noxref_1_c_6_p N_noxref_13_c_2030_n ) capacitor c=0.0431718f \
 //x=14.8 //y=0 //x2=14.105 //y2=0.615
cc_194 ( N_noxref_1_c_8_p N_noxref_13_M7_noxref_s ) capacitor c=0.00293348f \
 //x=21.09 //y=0 //x2=12.03 //y2=0.365
cc_195 ( N_noxref_1_c_38_p N_noxref_13_M7_noxref_s ) capacitor c=0.0149357f \
 //x=12.565 //y=0 //x2=12.03 //y2=0.365
cc_196 ( N_noxref_1_c_5_p N_noxref_13_M7_noxref_s ) capacitor c=0.058339f \
 //x=11.47 //y=0 //x2=12.03 //y2=0.365
cc_197 ( N_noxref_1_c_6_p N_noxref_13_M7_noxref_s ) capacitor c=0.00198043f \
 //x=14.8 //y=0 //x2=12.03 //y2=0.365
cc_198 ( N_noxref_1_M7_noxref_d N_noxref_13_M7_noxref_s ) capacitor \
 c=0.0334197f //x=12.46 //y=0.865 //x2=12.03 //y2=0.365
cc_199 ( N_noxref_1_c_6_p N_noxref_14_c_2072_n ) capacitor c=9.2064e-19 \
 //x=14.8 //y=0 //x2=16.65 //y2=2.08
cc_200 ( N_noxref_1_c_7_p N_noxref_14_c_2072_n ) capacitor c=9.53263e-19 \
 //x=18.13 //y=0 //x2=16.65 //y2=2.08
cc_201 ( N_noxref_1_c_7_p N_noxref_15_c_2141_n ) capacitor c=0.0462817f \
 //x=18.13 //y=0 //x2=17.305 //y2=1.655
cc_202 ( N_noxref_1_c_6_p N_noxref_15_c_2142_n ) capacitor c=9.64732e-19 \
 //x=14.8 //y=0 //x2=17.39 //y2=5.115
cc_203 ( N_noxref_1_c_6_p N_noxref_15_M10_noxref_d ) capacitor c=8.58106e-19 \
 //x=14.8 //y=0 //x2=16.76 //y2=0.905
cc_204 ( N_noxref_1_c_7_p N_noxref_15_M10_noxref_d ) capacitor c=0.00616547f \
 //x=18.13 //y=0 //x2=16.76 //y2=0.905
cc_205 ( N_noxref_1_M9_noxref_d N_noxref_15_M10_noxref_d ) capacitor \
 c=0.00143464f //x=15.79 //y=0.865 //x2=16.76 //y2=0.905
cc_206 ( N_noxref_1_c_8_p N_noxref_16_c_2213_n ) capacitor c=0.00565424f \
 //x=21.09 //y=0 //x2=16.38 //y2=1.58
cc_207 ( N_noxref_1_c_75_p N_noxref_16_c_2213_n ) capacitor c=0.00111428f \
 //x=15.895 //y=0 //x2=16.38 //y2=1.58
cc_208 ( N_noxref_1_c_82_p N_noxref_16_c_2213_n ) capacitor c=0.00180846f \
 //x=17.96 //y=0 //x2=16.38 //y2=1.58
cc_209 ( N_noxref_1_M9_noxref_d N_noxref_16_c_2213_n ) capacitor c=0.00901798f \
 //x=15.79 //y=0.865 //x2=16.38 //y2=1.58
cc_210 ( N_noxref_1_c_8_p N_noxref_16_c_2217_n ) capacitor c=0.005846f \
 //x=21.09 //y=0 //x2=16.465 //y2=0.615
cc_211 ( N_noxref_1_c_82_p N_noxref_16_c_2217_n ) capacitor c=0.0146208f \
 //x=17.96 //y=0 //x2=16.465 //y2=0.615
cc_212 ( N_noxref_1_M9_noxref_d N_noxref_16_c_2217_n ) capacitor c=0.033812f \
 //x=15.79 //y=0.865 //x2=16.465 //y2=0.615
cc_213 ( N_noxref_1_c_6_p N_noxref_16_c_2220_n ) capacitor c=2.91423e-19 \
 //x=14.8 //y=0 //x2=16.465 //y2=1.495
cc_214 ( N_noxref_1_c_8_p N_noxref_16_c_2221_n ) capacitor c=0.0145018f \
 //x=21.09 //y=0 //x2=17.35 //y2=0.53
cc_215 ( N_noxref_1_c_82_p N_noxref_16_c_2221_n ) capacitor c=0.0371035f \
 //x=17.96 //y=0 //x2=17.35 //y2=0.53
cc_216 ( N_noxref_1_c_2_p N_noxref_16_c_2221_n ) capacitor c=0.00198885f \
 //x=21.09 //y=0 //x2=17.35 //y2=0.53
cc_217 ( N_noxref_1_c_8_p N_noxref_16_c_2224_n ) capacitor c=0.00579979f \
 //x=21.09 //y=0 //x2=17.435 //y2=0.615
cc_218 ( N_noxref_1_c_82_p N_noxref_16_c_2224_n ) capacitor c=0.0144264f \
 //x=17.96 //y=0 //x2=17.435 //y2=0.615
cc_219 ( N_noxref_1_c_7_p N_noxref_16_c_2224_n ) capacitor c=0.0431718f \
 //x=18.13 //y=0 //x2=17.435 //y2=0.615
cc_220 ( N_noxref_1_c_8_p N_noxref_16_M9_noxref_s ) capacitor c=0.00302994f \
 //x=21.09 //y=0 //x2=15.36 //y2=0.365
cc_221 ( N_noxref_1_c_75_p N_noxref_16_M9_noxref_s ) capacitor c=0.0146208f \
 //x=15.895 //y=0 //x2=15.36 //y2=0.365
cc_222 ( N_noxref_1_c_6_p N_noxref_16_M9_noxref_s ) capacitor c=0.058339f \
 //x=14.8 //y=0 //x2=15.36 //y2=0.365
cc_223 ( N_noxref_1_c_7_p N_noxref_16_M9_noxref_s ) capacitor c=0.00198043f \
 //x=18.13 //y=0 //x2=15.36 //y2=0.365
cc_224 ( N_noxref_1_M9_noxref_d N_noxref_16_M9_noxref_s ) capacitor \
 c=0.0334197f //x=15.79 //y=0.865 //x2=15.36 //y2=0.365
cc_225 ( N_noxref_1_c_7_p N_noxref_17_c_2265_n ) capacitor c=0.0179404f \
 //x=18.13 //y=0 //x2=19.24 //y2=2.08
cc_226 ( N_noxref_1_c_226_p N_noxref_17_c_2266_n ) capacitor c=0.00135046f \
 //x=19.225 //y=0 //x2=19.045 //y2=0.865
cc_227 ( N_noxref_1_M11_noxref_d N_noxref_17_c_2266_n ) capacitor \
 c=0.00220047f //x=19.12 //y=0.865 //x2=19.045 //y2=0.865
cc_228 ( N_noxref_1_M11_noxref_d N_noxref_17_c_2268_n ) capacitor \
 c=0.00255985f //x=19.12 //y=0.865 //x2=19.045 //y2=1.21
cc_229 ( N_noxref_1_c_7_p N_noxref_17_c_2269_n ) capacitor c=0.0018059f \
 //x=18.13 //y=0 //x2=19.045 //y2=1.52
cc_230 ( N_noxref_1_c_7_p N_noxref_17_c_2270_n ) capacitor c=0.0114883f \
 //x=18.13 //y=0 //x2=19.045 //y2=1.915
cc_231 ( N_noxref_1_M11_noxref_d N_noxref_17_c_2271_n ) capacitor c=0.0131326f \
 //x=19.12 //y=0.865 //x2=19.42 //y2=0.71
cc_232 ( N_noxref_1_M11_noxref_d N_noxref_17_c_2272_n ) capacitor \
 c=0.00193127f //x=19.12 //y=0.865 //x2=19.42 //y2=1.365
cc_233 ( N_noxref_1_c_2_p N_noxref_17_c_2273_n ) capacitor c=0.00130622f \
 //x=21.09 //y=0 //x2=19.575 //y2=0.865
cc_234 ( N_noxref_1_M11_noxref_d N_noxref_17_c_2273_n ) capacitor \
 c=0.00257848f //x=19.12 //y=0.865 //x2=19.575 //y2=0.865
cc_235 ( N_noxref_1_M11_noxref_d N_noxref_17_c_2275_n ) capacitor \
 c=0.00255985f //x=19.12 //y=0.865 //x2=19.575 //y2=1.21
cc_236 ( N_noxref_1_c_2_p N_noxref_18_c_2325_n ) capacitor c=0.0468439f \
 //x=21.09 //y=0 //x2=20.635 //y2=1.655
cc_237 ( N_noxref_1_c_7_p N_noxref_18_c_2326_n ) capacitor c=9.64732e-19 \
 //x=18.13 //y=0 //x2=20.72 //y2=5.115
cc_238 ( N_noxref_1_c_2_p N_noxref_18_M12_noxref_d ) capacitor c=0.00618259f \
 //x=21.09 //y=0 //x2=20.09 //y2=0.905
cc_239 ( N_noxref_1_c_7_p N_noxref_18_M12_noxref_d ) capacitor c=8.58106e-19 \
 //x=18.13 //y=0 //x2=20.09 //y2=0.905
cc_240 ( N_noxref_1_M11_noxref_d N_noxref_18_M12_noxref_d ) capacitor \
 c=0.00143464f //x=19.12 //y=0.865 //x2=20.09 //y2=0.905
cc_241 ( N_noxref_1_c_8_p N_noxref_19_c_2390_n ) capacitor c=0.00571027f \
 //x=21.09 //y=0 //x2=19.71 //y2=1.58
cc_242 ( N_noxref_1_c_226_p N_noxref_19_c_2390_n ) capacitor c=0.00111428f \
 //x=19.225 //y=0 //x2=19.71 //y2=1.58
cc_243 ( N_noxref_1_c_2_p N_noxref_19_c_2390_n ) capacitor c=0.00180846f \
 //x=21.09 //y=0 //x2=19.71 //y2=1.58
cc_244 ( N_noxref_1_M11_noxref_d N_noxref_19_c_2390_n ) capacitor \
 c=0.00904677f //x=19.12 //y=0.865 //x2=19.71 //y2=1.58
cc_245 ( N_noxref_1_c_8_p N_noxref_19_c_2394_n ) capacitor c=0.00584537f \
 //x=21.09 //y=0 //x2=19.795 //y2=0.615
cc_246 ( N_noxref_1_c_2_p N_noxref_19_c_2394_n ) capacitor c=0.0146208f \
 //x=21.09 //y=0 //x2=19.795 //y2=0.615
cc_247 ( N_noxref_1_M11_noxref_d N_noxref_19_c_2394_n ) capacitor c=0.033812f \
 //x=19.12 //y=0.865 //x2=19.795 //y2=0.615
cc_248 ( N_noxref_1_c_7_p N_noxref_19_c_2397_n ) capacitor c=2.91423e-19 \
 //x=18.13 //y=0 //x2=19.795 //y2=1.495
cc_249 ( N_noxref_1_c_8_p N_noxref_19_c_2398_n ) capacitor c=0.0182917f \
 //x=21.09 //y=0 //x2=20.68 //y2=0.53
cc_250 ( N_noxref_1_c_2_p N_noxref_19_c_2398_n ) capacitor c=0.0390924f \
 //x=21.09 //y=0 //x2=20.68 //y2=0.53
cc_251 ( N_noxref_1_c_8_p N_noxref_19_c_2400_n ) capacitor c=0.00719615f \
 //x=21.09 //y=0 //x2=20.765 //y2=0.615
cc_252 ( N_noxref_1_c_2_p N_noxref_19_c_2400_n ) capacitor c=0.0584079f \
 //x=21.09 //y=0 //x2=20.765 //y2=0.615
cc_253 ( N_noxref_1_c_8_p N_noxref_19_M11_noxref_s ) capacitor c=0.005846f \
 //x=21.09 //y=0 //x2=18.69 //y2=0.365
cc_254 ( N_noxref_1_c_226_p N_noxref_19_M11_noxref_s ) capacitor c=0.0146208f \
 //x=19.225 //y=0 //x2=18.69 //y2=0.365
cc_255 ( N_noxref_1_c_2_p N_noxref_19_M11_noxref_s ) capacitor c=0.00198482f \
 //x=21.09 //y=0 //x2=18.69 //y2=0.365
cc_256 ( N_noxref_1_c_7_p N_noxref_19_M11_noxref_s ) capacitor c=0.058339f \
 //x=18.13 //y=0 //x2=18.69 //y2=0.365
cc_257 ( N_noxref_1_M11_noxref_d N_noxref_19_M11_noxref_s ) capacitor \
 c=0.0334197f //x=19.12 //y=0.865 //x2=18.69 //y2=0.365
cc_258 ( N_noxref_2_c_260_n N_noxref_3_c_558_n ) capacitor c=6.58823e-19 \
 //x=4.81 //y=7.4 //x2=3.33 //y2=2.08
cc_259 ( N_noxref_2_c_266_p N_noxref_3_c_576_n ) capacitor c=0.00453663f \
 //x=21.09 //y=7.4 //x2=6.835 //y2=5.2
cc_260 ( N_noxref_2_c_267_p N_noxref_3_c_576_n ) capacitor c=4.48391e-19 \
 //x=6.395 //y=7.4 //x2=6.835 //y2=5.2
cc_261 ( N_noxref_2_c_268_p N_noxref_3_c_576_n ) capacitor c=4.48391e-19 \
 //x=7.275 //y=7.4 //x2=6.835 //y2=5.2
cc_262 ( N_noxref_2_M20_noxref_d N_noxref_3_c_576_n ) capacitor c=0.0124542f \
 //x=6.335 //y=5.02 //x2=6.835 //y2=5.2
cc_263 ( N_noxref_2_c_260_n N_noxref_3_c_580_n ) capacitor c=0.00985474f \
 //x=4.81 //y=7.4 //x2=6.125 //y2=5.2
cc_264 ( N_noxref_2_M19_noxref_s N_noxref_3_c_580_n ) capacitor c=0.087833f \
 //x=5.465 //y=5.02 //x2=6.125 //y2=5.2
cc_265 ( N_noxref_2_c_266_p N_noxref_3_c_582_n ) capacitor c=0.00301575f \
 //x=21.09 //y=7.4 //x2=7.315 //y2=5.2
cc_266 ( N_noxref_2_c_268_p N_noxref_3_c_582_n ) capacitor c=7.72068e-19 \
 //x=7.275 //y=7.4 //x2=7.315 //y2=5.2
cc_267 ( N_noxref_2_M22_noxref_d N_noxref_3_c_582_n ) capacitor c=0.0158515f \
 //x=7.215 //y=5.02 //x2=7.315 //y2=5.2
cc_268 ( N_noxref_2_M23_noxref_s N_noxref_3_c_582_n ) capacitor c=2.44532e-19 \
 //x=8.795 //y=5.02 //x2=7.315 //y2=5.2
cc_269 ( N_noxref_2_c_260_n N_noxref_3_c_560_n ) capacitor c=0.00151618f \
 //x=4.81 //y=7.4 //x2=7.4 //y2=3.33
cc_270 ( N_noxref_2_c_261_n N_noxref_3_c_560_n ) capacitor c=0.0429414f \
 //x=8.14 //y=7.4 //x2=7.4 //y2=3.33
cc_271 ( N_noxref_2_c_266_p N_noxref_3_c_561_n ) capacitor c=0.00125279f \
 //x=21.09 //y=7.4 //x2=9.25 //y2=2.08
cc_272 ( N_noxref_2_c_279_p N_noxref_3_c_561_n ) capacitor c=2.87256e-19 \
 //x=9.725 //y=7.4 //x2=9.25 //y2=2.08
cc_273 ( N_noxref_2_c_261_n N_noxref_3_c_561_n ) capacitor c=0.0134208f \
 //x=8.14 //y=7.4 //x2=9.25 //y2=2.08
cc_274 ( N_noxref_2_c_281_p N_noxref_3_M17_noxref_g ) capacitor c=0.00675175f \
 //x=3.645 //y=7.4 //x2=3.07 //y2=6.02
cc_275 ( N_noxref_2_M16_noxref_d N_noxref_3_M17_noxref_g ) capacitor \
 c=0.015318f //x=2.705 //y=5.02 //x2=3.07 //y2=6.02
cc_276 ( N_noxref_2_c_281_p N_noxref_3_M18_noxref_g ) capacitor c=0.00675379f \
 //x=3.645 //y=7.4 //x2=3.51 //y2=6.02
cc_277 ( N_noxref_2_M18_noxref_d N_noxref_3_M18_noxref_g ) capacitor \
 c=0.0394719f //x=3.585 //y=5.02 //x2=3.51 //y2=6.02
cc_278 ( N_noxref_2_c_279_p N_noxref_3_M23_noxref_g ) capacitor c=0.00726866f \
 //x=9.725 //y=7.4 //x2=9.15 //y2=6.02
cc_279 ( N_noxref_2_M23_noxref_s N_noxref_3_M23_noxref_g ) capacitor \
 c=0.054195f //x=8.795 //y=5.02 //x2=9.15 //y2=6.02
cc_280 ( N_noxref_2_c_279_p N_noxref_3_M24_noxref_g ) capacitor c=0.00672952f \
 //x=9.725 //y=7.4 //x2=9.59 //y2=6.02
cc_281 ( N_noxref_2_M24_noxref_d N_noxref_3_M24_noxref_g ) capacitor \
 c=0.015318f //x=9.665 //y=5.02 //x2=9.59 //y2=6.02
cc_282 ( N_noxref_2_c_261_n N_noxref_3_c_599_n ) capacitor c=0.0150435f \
 //x=8.14 //y=7.4 //x2=9.25 //y2=4.7
cc_283 ( N_noxref_2_c_266_p N_noxref_3_M19_noxref_d ) capacitor c=0.00275225f \
 //x=21.09 //y=7.4 //x2=5.895 //y2=5.02
cc_284 ( N_noxref_2_c_267_p N_noxref_3_M19_noxref_d ) capacitor c=0.0140317f \
 //x=6.395 //y=7.4 //x2=5.895 //y2=5.02
cc_285 ( N_noxref_2_c_261_n N_noxref_3_M19_noxref_d ) capacitor c=6.94454e-19 \
 //x=8.14 //y=7.4 //x2=5.895 //y2=5.02
cc_286 ( N_noxref_2_M20_noxref_d N_noxref_3_M19_noxref_d ) capacitor \
 c=0.0664752f //x=6.335 //y=5.02 //x2=5.895 //y2=5.02
cc_287 ( N_noxref_2_c_266_p N_noxref_3_M21_noxref_d ) capacitor c=0.00275225f \
 //x=21.09 //y=7.4 //x2=6.775 //y2=5.02
cc_288 ( N_noxref_2_c_268_p N_noxref_3_M21_noxref_d ) capacitor c=0.0140317f \
 //x=7.275 //y=7.4 //x2=6.775 //y2=5.02
cc_289 ( N_noxref_2_c_261_n N_noxref_3_M21_noxref_d ) capacitor c=0.0120541f \
 //x=8.14 //y=7.4 //x2=6.775 //y2=5.02
cc_290 ( N_noxref_2_M19_noxref_s N_noxref_3_M21_noxref_d ) capacitor \
 c=0.00111971f //x=5.465 //y=5.02 //x2=6.775 //y2=5.02
cc_291 ( N_noxref_2_M20_noxref_d N_noxref_3_M21_noxref_d ) capacitor \
 c=0.0664752f //x=6.335 //y=5.02 //x2=6.775 //y2=5.02
cc_292 ( N_noxref_2_M22_noxref_d N_noxref_3_M21_noxref_d ) capacitor \
 c=0.0664752f //x=7.215 //y=5.02 //x2=6.775 //y2=5.02
cc_293 ( N_noxref_2_M23_noxref_s N_noxref_3_M21_noxref_d ) capacitor \
 c=4.54516e-19 //x=8.795 //y=5.02 //x2=6.775 //y2=5.02
cc_294 ( N_noxref_2_c_266_p N_noxref_4_c_800_n ) capacitor c=0.00453663f \
 //x=21.09 //y=7.4 //x2=10.165 //y2=5.2
cc_295 ( N_noxref_2_c_279_p N_noxref_4_c_800_n ) capacitor c=4.48391e-19 \
 //x=9.725 //y=7.4 //x2=10.165 //y2=5.2
cc_296 ( N_noxref_2_c_303_p N_noxref_4_c_800_n ) capacitor c=4.48391e-19 \
 //x=10.605 //y=7.4 //x2=10.165 //y2=5.2
cc_297 ( N_noxref_2_M24_noxref_d N_noxref_4_c_800_n ) capacitor c=0.0124542f \
 //x=9.665 //y=5.02 //x2=10.165 //y2=5.2
cc_298 ( N_noxref_2_c_261_n N_noxref_4_c_804_n ) capacitor c=0.00985474f \
 //x=8.14 //y=7.4 //x2=9.455 //y2=5.2
cc_299 ( N_noxref_2_M23_noxref_s N_noxref_4_c_804_n ) capacitor c=0.087833f \
 //x=8.795 //y=5.02 //x2=9.455 //y2=5.2
cc_300 ( N_noxref_2_c_266_p N_noxref_4_c_806_n ) capacitor c=0.00301575f \
 //x=21.09 //y=7.4 //x2=10.645 //y2=5.2
cc_301 ( N_noxref_2_c_303_p N_noxref_4_c_806_n ) capacitor c=7.72068e-19 \
 //x=10.605 //y=7.4 //x2=10.645 //y2=5.2
cc_302 ( N_noxref_2_M26_noxref_d N_noxref_4_c_806_n ) capacitor c=0.0158515f \
 //x=10.545 //y=5.02 //x2=10.645 //y2=5.2
cc_303 ( N_noxref_2_M27_noxref_s N_noxref_4_c_806_n ) capacitor c=2.44532e-19 \
 //x=12.125 //y=5.02 //x2=10.645 //y2=5.2
cc_304 ( N_noxref_2_c_261_n N_noxref_4_c_785_n ) capacitor c=0.00151618f \
 //x=8.14 //y=7.4 //x2=10.73 //y2=3.33
cc_305 ( N_noxref_2_c_262_n N_noxref_4_c_785_n ) capacitor c=0.0427674f \
 //x=11.47 //y=7.4 //x2=10.73 //y2=3.33
cc_306 ( N_noxref_2_c_266_p N_noxref_4_c_786_n ) capacitor c=0.00125279f \
 //x=21.09 //y=7.4 //x2=12.58 //y2=2.08
cc_307 ( N_noxref_2_c_314_p N_noxref_4_c_786_n ) capacitor c=2.87256e-19 \
 //x=13.055 //y=7.4 //x2=12.58 //y2=2.08
cc_308 ( N_noxref_2_c_262_n N_noxref_4_c_786_n ) capacitor c=0.0133228f \
 //x=11.47 //y=7.4 //x2=12.58 //y2=2.08
cc_309 ( N_noxref_2_c_314_p N_noxref_4_M27_noxref_g ) capacitor c=0.00726866f \
 //x=13.055 //y=7.4 //x2=12.48 //y2=6.02
cc_310 ( N_noxref_2_M27_noxref_s N_noxref_4_M27_noxref_g ) capacitor \
 c=0.054195f //x=12.125 //y=5.02 //x2=12.48 //y2=6.02
cc_311 ( N_noxref_2_c_314_p N_noxref_4_M28_noxref_g ) capacitor c=0.00672952f \
 //x=13.055 //y=7.4 //x2=12.92 //y2=6.02
cc_312 ( N_noxref_2_M28_noxref_d N_noxref_4_M28_noxref_g ) capacitor \
 c=0.015318f //x=12.995 //y=5.02 //x2=12.92 //y2=6.02
cc_313 ( N_noxref_2_c_262_n N_noxref_4_c_819_n ) capacitor c=0.0149273f \
 //x=11.47 //y=7.4 //x2=12.58 //y2=4.7
cc_314 ( N_noxref_2_c_266_p N_noxref_4_M23_noxref_d ) capacitor c=0.00275225f \
 //x=21.09 //y=7.4 //x2=9.225 //y2=5.02
cc_315 ( N_noxref_2_c_279_p N_noxref_4_M23_noxref_d ) capacitor c=0.0140317f \
 //x=9.725 //y=7.4 //x2=9.225 //y2=5.02
cc_316 ( N_noxref_2_c_262_n N_noxref_4_M23_noxref_d ) capacitor c=6.94454e-19 \
 //x=11.47 //y=7.4 //x2=9.225 //y2=5.02
cc_317 ( N_noxref_2_M24_noxref_d N_noxref_4_M23_noxref_d ) capacitor \
 c=0.0664752f //x=9.665 //y=5.02 //x2=9.225 //y2=5.02
cc_318 ( N_noxref_2_c_266_p N_noxref_4_M25_noxref_d ) capacitor c=0.00275225f \
 //x=21.09 //y=7.4 //x2=10.105 //y2=5.02
cc_319 ( N_noxref_2_c_303_p N_noxref_4_M25_noxref_d ) capacitor c=0.0140317f \
 //x=10.605 //y=7.4 //x2=10.105 //y2=5.02
cc_320 ( N_noxref_2_c_262_n N_noxref_4_M25_noxref_d ) capacitor c=0.0120541f \
 //x=11.47 //y=7.4 //x2=10.105 //y2=5.02
cc_321 ( N_noxref_2_M23_noxref_s N_noxref_4_M25_noxref_d ) capacitor \
 c=0.00111971f //x=8.795 //y=5.02 //x2=10.105 //y2=5.02
cc_322 ( N_noxref_2_M24_noxref_d N_noxref_4_M25_noxref_d ) capacitor \
 c=0.0664752f //x=9.665 //y=5.02 //x2=10.105 //y2=5.02
cc_323 ( N_noxref_2_M26_noxref_d N_noxref_4_M25_noxref_d ) capacitor \
 c=0.0664752f //x=10.545 //y=5.02 //x2=10.105 //y2=5.02
cc_324 ( N_noxref_2_M27_noxref_s N_noxref_4_M25_noxref_d ) capacitor \
 c=4.54516e-19 //x=12.125 //y=5.02 //x2=10.105 //y2=5.02
cc_325 ( N_noxref_2_c_266_p N_noxref_5_c_932_n ) capacitor c=0.0824294f \
 //x=21.09 //y=7.4 //x2=13.205 //y2=4.44
cc_326 ( N_noxref_2_c_333_p N_noxref_5_c_932_n ) capacitor c=0.00258496f \
 //x=4.64 //y=7.4 //x2=13.205 //y2=4.44
cc_327 ( N_noxref_2_c_334_p N_noxref_5_c_932_n ) capacitor c=0.00209689f \
 //x=5.515 //y=7.4 //x2=13.205 //y2=4.44
cc_328 ( N_noxref_2_c_267_p N_noxref_5_c_932_n ) capacitor c=7.81728e-19 \
 //x=6.395 //y=7.4 //x2=13.205 //y2=4.44
cc_329 ( N_noxref_2_c_336_p N_noxref_5_c_932_n ) capacitor c=0.00205475f \
 //x=7.97 //y=7.4 //x2=13.205 //y2=4.44
cc_330 ( N_noxref_2_c_337_p N_noxref_5_c_932_n ) capacitor c=0.00209689f \
 //x=8.845 //y=7.4 //x2=13.205 //y2=4.44
cc_331 ( N_noxref_2_c_279_p N_noxref_5_c_932_n ) capacitor c=7.81728e-19 \
 //x=9.725 //y=7.4 //x2=13.205 //y2=4.44
cc_332 ( N_noxref_2_c_339_p N_noxref_5_c_932_n ) capacitor c=0.00205475f \
 //x=11.3 //y=7.4 //x2=13.205 //y2=4.44
cc_333 ( N_noxref_2_c_340_p N_noxref_5_c_932_n ) capacitor c=0.00209689f \
 //x=12.175 //y=7.4 //x2=13.205 //y2=4.44
cc_334 ( N_noxref_2_c_314_p N_noxref_5_c_932_n ) capacitor c=7.81728e-19 \
 //x=13.055 //y=7.4 //x2=13.205 //y2=4.44
cc_335 ( N_noxref_2_c_260_n N_noxref_5_c_932_n ) capacitor c=0.0389825f \
 //x=4.81 //y=7.4 //x2=13.205 //y2=4.44
cc_336 ( N_noxref_2_c_261_n N_noxref_5_c_932_n ) capacitor c=0.0389825f \
 //x=8.14 //y=7.4 //x2=13.205 //y2=4.44
cc_337 ( N_noxref_2_c_262_n N_noxref_5_c_932_n ) capacitor c=0.0389825f \
 //x=11.47 //y=7.4 //x2=13.205 //y2=4.44
cc_338 ( N_noxref_2_M19_noxref_s N_noxref_5_c_932_n ) capacitor c=0.00541054f \
 //x=5.465 //y=5.02 //x2=13.205 //y2=4.44
cc_339 ( N_noxref_2_M22_noxref_d N_noxref_5_c_932_n ) capacitor c=6.7165e-19 \
 //x=7.215 //y=5.02 //x2=13.205 //y2=4.44
cc_340 ( N_noxref_2_M23_noxref_s N_noxref_5_c_932_n ) capacitor c=0.00541054f \
 //x=8.795 //y=5.02 //x2=13.205 //y2=4.44
cc_341 ( N_noxref_2_M26_noxref_d N_noxref_5_c_932_n ) capacitor c=6.7165e-19 \
 //x=10.545 //y=5.02 //x2=13.205 //y2=4.44
cc_342 ( N_noxref_2_M27_noxref_s N_noxref_5_c_932_n ) capacitor c=0.00541054f \
 //x=12.125 //y=5.02 //x2=13.205 //y2=4.44
cc_343 ( N_noxref_2_c_266_p N_noxref_5_c_950_n ) capacitor c=0.00146064f \
 //x=21.09 //y=7.4 //x2=2.335 //y2=4.44
cc_344 ( N_noxref_2_c_266_p N_noxref_5_c_929_n ) capacitor c=2.03287e-19 \
 //x=21.09 //y=7.4 //x2=2.22 //y2=2.08
cc_345 ( N_noxref_2_c_258_n N_noxref_5_c_929_n ) capacitor c=9.53425e-19 \
 //x=0.74 //y=7.4 //x2=2.22 //y2=2.08
cc_346 ( N_noxref_2_c_262_n N_noxref_5_c_930_n ) capacitor c=5.27482e-19 \
 //x=11.47 //y=7.4 //x2=13.32 //y2=2.08
cc_347 ( N_noxref_2_c_263_n N_noxref_5_c_930_n ) capacitor c=7.54518e-19 \
 //x=14.8 //y=7.4 //x2=13.32 //y2=2.08
cc_348 ( N_noxref_2_c_355_p N_noxref_5_M15_noxref_g ) capacitor c=0.00676195f \
 //x=2.765 //y=7.4 //x2=2.19 //y2=6.02
cc_349 ( N_noxref_2_M14_noxref_d N_noxref_5_M15_noxref_g ) capacitor \
 c=0.015318f //x=1.825 //y=5.02 //x2=2.19 //y2=6.02
cc_350 ( N_noxref_2_c_355_p N_noxref_5_M16_noxref_g ) capacitor c=0.00675175f \
 //x=2.765 //y=7.4 //x2=2.63 //y2=6.02
cc_351 ( N_noxref_2_M16_noxref_d N_noxref_5_M16_noxref_g ) capacitor \
 c=0.015318f //x=2.705 //y=5.02 //x2=2.63 //y2=6.02
cc_352 ( N_noxref_2_c_359_p N_noxref_5_M29_noxref_g ) capacitor c=0.00673971f \
 //x=13.935 //y=7.4 //x2=13.36 //y2=6.02
cc_353 ( N_noxref_2_M28_noxref_d N_noxref_5_M29_noxref_g ) capacitor \
 c=0.015318f //x=12.995 //y=5.02 //x2=13.36 //y2=6.02
cc_354 ( N_noxref_2_c_359_p N_noxref_5_M30_noxref_g ) capacitor c=0.00672952f \
 //x=13.935 //y=7.4 //x2=13.8 //y2=6.02
cc_355 ( N_noxref_2_c_263_n N_noxref_5_M30_noxref_g ) capacitor c=0.00864163f \
 //x=14.8 //y=7.4 //x2=13.8 //y2=6.02
cc_356 ( N_noxref_2_M30_noxref_d N_noxref_5_M30_noxref_g ) capacitor \
 c=0.0430452f //x=13.875 //y=5.02 //x2=13.8 //y2=6.02
cc_357 ( N_noxref_2_c_263_n N_noxref_6_c_1134_n ) capacitor c=0.00290959f \
 //x=14.8 //y=7.4 //x2=15.795 //y2=3.7
cc_358 ( N_noxref_2_c_266_p N_noxref_6_c_1161_n ) capacitor c=0.00449316f \
 //x=21.09 //y=7.4 //x2=2.325 //y2=5.155
cc_359 ( N_noxref_2_c_366_p N_noxref_6_c_1161_n ) capacitor c=4.32228e-19 \
 //x=1.885 //y=7.4 //x2=2.325 //y2=5.155
cc_360 ( N_noxref_2_c_355_p N_noxref_6_c_1161_n ) capacitor c=4.31906e-19 \
 //x=2.765 //y=7.4 //x2=2.325 //y2=5.155
cc_361 ( N_noxref_2_M14_noxref_d N_noxref_6_c_1161_n ) capacitor c=0.0115147f \
 //x=1.825 //y=5.02 //x2=2.325 //y2=5.155
cc_362 ( N_noxref_2_c_258_n N_noxref_6_c_1165_n ) capacitor c=0.00880189f \
 //x=0.74 //y=7.4 //x2=1.615 //y2=5.155
cc_363 ( N_noxref_2_M13_noxref_s N_noxref_6_c_1165_n ) capacitor c=0.0831083f \
 //x=0.955 //y=5.02 //x2=1.615 //y2=5.155
cc_364 ( N_noxref_2_c_266_p N_noxref_6_c_1167_n ) capacitor c=0.0044221f \
 //x=21.09 //y=7.4 //x2=3.205 //y2=5.155
cc_365 ( N_noxref_2_c_355_p N_noxref_6_c_1167_n ) capacitor c=4.31931e-19 \
 //x=2.765 //y=7.4 //x2=3.205 //y2=5.155
cc_366 ( N_noxref_2_c_281_p N_noxref_6_c_1167_n ) capacitor c=4.31931e-19 \
 //x=3.645 //y=7.4 //x2=3.205 //y2=5.155
cc_367 ( N_noxref_2_M16_noxref_d N_noxref_6_c_1167_n ) capacitor c=0.0112985f \
 //x=2.705 //y=5.02 //x2=3.205 //y2=5.155
cc_368 ( N_noxref_2_c_266_p N_noxref_6_c_1171_n ) capacitor c=0.00434174f \
 //x=21.09 //y=7.4 //x2=3.985 //y2=5.155
cc_369 ( N_noxref_2_c_281_p N_noxref_6_c_1171_n ) capacitor c=7.46626e-19 \
 //x=3.645 //y=7.4 //x2=3.985 //y2=5.155
cc_370 ( N_noxref_2_c_333_p N_noxref_6_c_1171_n ) capacitor c=0.00198565f \
 //x=4.64 //y=7.4 //x2=3.985 //y2=5.155
cc_371 ( N_noxref_2_M18_noxref_d N_noxref_6_c_1171_n ) capacitor c=0.0112985f \
 //x=3.585 //y=5.02 //x2=3.985 //y2=5.155
cc_372 ( N_noxref_2_c_260_n N_noxref_6_c_1175_n ) capacitor c=0.0426341f \
 //x=4.81 //y=7.4 //x2=4.07 //y2=3.7
cc_373 ( N_noxref_2_c_266_p N_noxref_6_c_1137_n ) capacitor c=0.00125279f \
 //x=21.09 //y=7.4 //x2=5.92 //y2=2.08
cc_374 ( N_noxref_2_c_267_p N_noxref_6_c_1137_n ) capacitor c=2.87256e-19 \
 //x=6.395 //y=7.4 //x2=5.92 //y2=2.08
cc_375 ( N_noxref_2_c_260_n N_noxref_6_c_1137_n ) capacitor c=0.0134665f \
 //x=4.81 //y=7.4 //x2=5.92 //y2=2.08
cc_376 ( N_noxref_2_c_266_p N_noxref_6_c_1138_n ) capacitor c=0.00126216f \
 //x=21.09 //y=7.4 //x2=15.91 //y2=2.08
cc_377 ( N_noxref_2_c_384_p N_noxref_6_c_1138_n ) capacitor c=2.87813e-19 \
 //x=16.385 //y=7.4 //x2=15.91 //y2=2.08
cc_378 ( N_noxref_2_c_263_n N_noxref_6_c_1138_n ) capacitor c=0.0157486f \
 //x=14.8 //y=7.4 //x2=15.91 //y2=2.08
cc_379 ( N_noxref_2_c_267_p N_noxref_6_M19_noxref_g ) capacitor c=0.00726866f \
 //x=6.395 //y=7.4 //x2=5.82 //y2=6.02
cc_380 ( N_noxref_2_M19_noxref_s N_noxref_6_M19_noxref_g ) capacitor \
 c=0.054195f //x=5.465 //y=5.02 //x2=5.82 //y2=6.02
cc_381 ( N_noxref_2_c_267_p N_noxref_6_M20_noxref_g ) capacitor c=0.00672952f \
 //x=6.395 //y=7.4 //x2=6.26 //y2=6.02
cc_382 ( N_noxref_2_M20_noxref_d N_noxref_6_M20_noxref_g ) capacitor \
 c=0.015318f //x=6.335 //y=5.02 //x2=6.26 //y2=6.02
cc_383 ( N_noxref_2_c_384_p N_noxref_6_M31_noxref_g ) capacitor c=0.00726866f \
 //x=16.385 //y=7.4 //x2=15.81 //y2=6.02
cc_384 ( N_noxref_2_M31_noxref_s N_noxref_6_M31_noxref_g ) capacitor \
 c=0.054195f //x=15.455 //y=5.02 //x2=15.81 //y2=6.02
cc_385 ( N_noxref_2_c_384_p N_noxref_6_M32_noxref_g ) capacitor c=0.00672952f \
 //x=16.385 //y=7.4 //x2=16.25 //y2=6.02
cc_386 ( N_noxref_2_M32_noxref_d N_noxref_6_M32_noxref_g ) capacitor \
 c=0.015318f //x=16.325 //y=5.02 //x2=16.25 //y2=6.02
cc_387 ( N_noxref_2_c_260_n N_noxref_6_c_1190_n ) capacitor c=0.015293f \
 //x=4.81 //y=7.4 //x2=5.92 //y2=4.7
cc_388 ( N_noxref_2_c_263_n N_noxref_6_c_1191_n ) capacitor c=0.0149273f \
 //x=14.8 //y=7.4 //x2=15.91 //y2=4.7
cc_389 ( N_noxref_2_c_266_p N_noxref_6_M13_noxref_d ) capacitor c=0.00285091f \
 //x=21.09 //y=7.4 //x2=1.385 //y2=5.02
cc_390 ( N_noxref_2_c_366_p N_noxref_6_M13_noxref_d ) capacitor c=0.0141016f \
 //x=1.885 //y=7.4 //x2=1.385 //y2=5.02
cc_391 ( N_noxref_2_M14_noxref_d N_noxref_6_M13_noxref_d ) capacitor \
 c=0.0664752f //x=1.825 //y=5.02 //x2=1.385 //y2=5.02
cc_392 ( N_noxref_2_c_266_p N_noxref_6_M15_noxref_d ) capacitor c=0.00275186f \
 //x=21.09 //y=7.4 //x2=2.265 //y2=5.02
cc_393 ( N_noxref_2_c_355_p N_noxref_6_M15_noxref_d ) capacitor c=0.0140346f \
 //x=2.765 //y=7.4 //x2=2.265 //y2=5.02
cc_394 ( N_noxref_2_c_260_n N_noxref_6_M15_noxref_d ) capacitor c=4.9285e-19 \
 //x=4.81 //y=7.4 //x2=2.265 //y2=5.02
cc_395 ( N_noxref_2_M13_noxref_s N_noxref_6_M15_noxref_d ) capacitor \
 c=0.00130656f //x=0.955 //y=5.02 //x2=2.265 //y2=5.02
cc_396 ( N_noxref_2_M14_noxref_d N_noxref_6_M15_noxref_d ) capacitor \
 c=0.0664752f //x=1.825 //y=5.02 //x2=2.265 //y2=5.02
cc_397 ( N_noxref_2_M16_noxref_d N_noxref_6_M15_noxref_d ) capacitor \
 c=0.0664752f //x=2.705 //y=5.02 //x2=2.265 //y2=5.02
cc_398 ( N_noxref_2_c_266_p N_noxref_6_M17_noxref_d ) capacitor c=0.00275235f \
 //x=21.09 //y=7.4 //x2=3.145 //y2=5.02
cc_399 ( N_noxref_2_c_281_p N_noxref_6_M17_noxref_d ) capacitor c=0.0137384f \
 //x=3.645 //y=7.4 //x2=3.145 //y2=5.02
cc_400 ( N_noxref_2_c_260_n N_noxref_6_M17_noxref_d ) capacitor c=0.00939849f \
 //x=4.81 //y=7.4 //x2=3.145 //y2=5.02
cc_401 ( N_noxref_2_M16_noxref_d N_noxref_6_M17_noxref_d ) capacitor \
 c=0.0664752f //x=2.705 //y=5.02 //x2=3.145 //y2=5.02
cc_402 ( N_noxref_2_M18_noxref_d N_noxref_6_M17_noxref_d ) capacitor \
 c=0.0664752f //x=3.585 //y=5.02 //x2=3.145 //y2=5.02
cc_403 ( N_noxref_2_M19_noxref_s N_noxref_6_M17_noxref_d ) capacitor \
 c=4.52683e-19 //x=5.465 //y=5.02 //x2=3.145 //y2=5.02
cc_404 ( N_noxref_2_c_266_p N_noxref_7_c_1385_n ) capacitor c=0.035625f \
 //x=21.09 //y=7.4 //x2=9.875 //y2=4.07
cc_405 ( N_noxref_2_c_366_p N_noxref_7_c_1385_n ) capacitor c=0.00113322f \
 //x=1.885 //y=7.4 //x2=9.875 //y2=4.07
cc_406 ( N_noxref_2_c_260_n N_noxref_7_c_1385_n ) capacitor c=0.0140578f \
 //x=4.81 //y=7.4 //x2=9.875 //y2=4.07
cc_407 ( N_noxref_2_c_261_n N_noxref_7_c_1385_n ) capacitor c=0.0140578f \
 //x=8.14 //y=7.4 //x2=9.875 //y2=4.07
cc_408 ( N_noxref_2_c_266_p N_noxref_7_c_1386_n ) capacitor c=0.00189266f \
 //x=21.09 //y=7.4 //x2=1.225 //y2=4.07
cc_409 ( N_noxref_2_c_258_n N_noxref_7_c_1386_n ) capacitor c=0.0017219f \
 //x=0.74 //y=7.4 //x2=1.225 //y2=4.07
cc_410 ( N_noxref_2_M13_noxref_s N_noxref_7_c_1386_n ) capacitor c=0.00128242f \
 //x=0.955 //y=5.02 //x2=1.225 //y2=4.07
cc_411 ( N_noxref_2_c_266_p N_noxref_7_c_1416_n ) capacitor c=0.0158405f \
 //x=21.09 //y=7.4 //x2=13.945 //y2=4.07
cc_412 ( N_noxref_2_c_262_n N_noxref_7_c_1416_n ) capacitor c=0.0140578f \
 //x=11.47 //y=7.4 //x2=13.945 //y2=4.07
cc_413 ( N_noxref_2_c_266_p N_noxref_7_c_1387_n ) capacitor c=0.0403243f \
 //x=21.09 //y=7.4 //x2=19.865 //y2=4.07
cc_414 ( N_noxref_2_c_421_p N_noxref_7_c_1387_n ) capacitor c=0.00161566f \
 //x=14.63 //y=7.4 //x2=19.865 //y2=4.07
cc_415 ( N_noxref_2_c_422_p N_noxref_7_c_1387_n ) capacitor c=0.00172186f \
 //x=15.505 //y=7.4 //x2=19.865 //y2=4.07
cc_416 ( N_noxref_2_c_384_p N_noxref_7_c_1387_n ) capacitor c=6.61469e-19 \
 //x=16.385 //y=7.4 //x2=19.865 //y2=4.07
cc_417 ( N_noxref_2_c_424_p N_noxref_7_c_1387_n ) capacitor c=0.00168692f \
 //x=17.96 //y=7.4 //x2=19.865 //y2=4.07
cc_418 ( N_noxref_2_c_425_p N_noxref_7_c_1387_n ) capacitor c=0.00172186f \
 //x=18.835 //y=7.4 //x2=19.865 //y2=4.07
cc_419 ( N_noxref_2_c_426_p N_noxref_7_c_1387_n ) capacitor c=6.61469e-19 \
 //x=19.715 //y=7.4 //x2=19.865 //y2=4.07
cc_420 ( N_noxref_2_c_263_n N_noxref_7_c_1387_n ) capacitor c=0.0269494f \
 //x=14.8 //y=7.4 //x2=19.865 //y2=4.07
cc_421 ( N_noxref_2_c_264_n N_noxref_7_c_1387_n ) capacitor c=0.0301177f \
 //x=18.13 //y=7.4 //x2=19.865 //y2=4.07
cc_422 ( N_noxref_2_M31_noxref_s N_noxref_7_c_1387_n ) capacitor c=0.00363031f \
 //x=15.455 //y=5.02 //x2=19.865 //y2=4.07
cc_423 ( N_noxref_2_M34_noxref_d N_noxref_7_c_1387_n ) capacitor c=5.05307e-19 \
 //x=17.205 //y=5.02 //x2=19.865 //y2=4.07
cc_424 ( N_noxref_2_M35_noxref_s N_noxref_7_c_1387_n ) capacitor c=0.00351625f \
 //x=18.785 //y=5.02 //x2=19.865 //y2=4.07
cc_425 ( N_noxref_2_c_266_p N_noxref_7_c_1430_n ) capacitor c=0.00172491f \
 //x=21.09 //y=7.4 //x2=14.175 //y2=4.07
cc_426 ( N_noxref_2_c_263_n N_noxref_7_c_1430_n ) capacitor c=0.00104972f \
 //x=14.8 //y=7.4 //x2=14.175 //y2=4.07
cc_427 ( N_noxref_2_M30_noxref_d N_noxref_7_c_1430_n ) capacitor c=5.14736e-19 \
 //x=13.875 //y=5.02 //x2=14.175 //y2=4.07
cc_428 ( N_noxref_2_c_266_p N_noxref_7_c_1389_n ) capacitor c=9.2251e-19 \
 //x=21.09 //y=7.4 //x2=1.11 //y2=2.08
cc_429 ( N_noxref_2_c_258_n N_noxref_7_c_1389_n ) capacitor c=0.0159723f \
 //x=0.74 //y=7.4 //x2=1.11 //y2=2.08
cc_430 ( N_noxref_2_M13_noxref_s N_noxref_7_c_1389_n ) capacitor c=0.0122951f \
 //x=0.955 //y=5.02 //x2=1.11 //y2=2.08
cc_431 ( N_noxref_2_c_261_n N_noxref_7_c_1390_n ) capacitor c=4.57806e-19 \
 //x=8.14 //y=7.4 //x2=9.99 //y2=2.08
cc_432 ( N_noxref_2_c_262_n N_noxref_7_c_1390_n ) capacitor c=3.69525e-19 \
 //x=11.47 //y=7.4 //x2=9.99 //y2=2.08
cc_433 ( N_noxref_2_c_266_p N_noxref_7_c_1438_n ) capacitor c=0.00453473f \
 //x=21.09 //y=7.4 //x2=13.495 //y2=5.2
cc_434 ( N_noxref_2_c_314_p N_noxref_7_c_1438_n ) capacitor c=4.48391e-19 \
 //x=13.055 //y=7.4 //x2=13.495 //y2=5.2
cc_435 ( N_noxref_2_c_359_p N_noxref_7_c_1438_n ) capacitor c=4.48377e-19 \
 //x=13.935 //y=7.4 //x2=13.495 //y2=5.2
cc_436 ( N_noxref_2_M28_noxref_d N_noxref_7_c_1438_n ) capacitor c=0.0124506f \
 //x=12.995 //y=5.02 //x2=13.495 //y2=5.2
cc_437 ( N_noxref_2_c_262_n N_noxref_7_c_1442_n ) capacitor c=0.00985474f \
 //x=11.47 //y=7.4 //x2=12.785 //y2=5.2
cc_438 ( N_noxref_2_M27_noxref_s N_noxref_7_c_1442_n ) capacitor c=0.087833f \
 //x=12.125 //y=5.02 //x2=12.785 //y2=5.2
cc_439 ( N_noxref_2_c_266_p N_noxref_7_c_1444_n ) capacitor c=0.00307016f \
 //x=21.09 //y=7.4 //x2=13.975 //y2=5.2
cc_440 ( N_noxref_2_c_359_p N_noxref_7_c_1444_n ) capacitor c=7.73167e-19 \
 //x=13.935 //y=7.4 //x2=13.975 //y2=5.2
cc_441 ( N_noxref_2_M30_noxref_d N_noxref_7_c_1444_n ) capacitor c=0.016133f \
 //x=13.875 //y=5.02 //x2=13.975 //y2=5.2
cc_442 ( N_noxref_2_M31_noxref_s N_noxref_7_c_1444_n ) capacitor c=2.44532e-19 \
 //x=15.455 //y=5.02 //x2=13.975 //y2=5.2
cc_443 ( N_noxref_2_c_262_n N_noxref_7_c_1393_n ) capacitor c=0.00151618f \
 //x=11.47 //y=7.4 //x2=14.06 //y2=4.07
cc_444 ( N_noxref_2_c_263_n N_noxref_7_c_1393_n ) capacitor c=0.0451944f \
 //x=14.8 //y=7.4 //x2=14.06 //y2=4.07
cc_445 ( N_noxref_2_c_259_n N_noxref_7_c_1394_n ) capacitor c=6.61994e-19 \
 //x=21.09 //y=7.4 //x2=19.98 //y2=2.08
cc_446 ( N_noxref_2_c_264_n N_noxref_7_c_1394_n ) capacitor c=6.2696e-19 \
 //x=18.13 //y=7.4 //x2=19.98 //y2=2.08
cc_447 ( N_noxref_2_c_366_p N_noxref_7_M13_noxref_g ) capacitor c=0.00749687f \
 //x=1.885 //y=7.4 //x2=1.31 //y2=6.02
cc_448 ( N_noxref_2_M13_noxref_s N_noxref_7_M13_noxref_g ) capacitor \
 c=0.0477201f //x=0.955 //y=5.02 //x2=1.31 //y2=6.02
cc_449 ( N_noxref_2_c_366_p N_noxref_7_M14_noxref_g ) capacitor c=0.00675175f \
 //x=1.885 //y=7.4 //x2=1.75 //y2=6.02
cc_450 ( N_noxref_2_M14_noxref_d N_noxref_7_M14_noxref_g ) capacitor \
 c=0.015318f //x=1.825 //y=5.02 //x2=1.75 //y2=6.02
cc_451 ( N_noxref_2_c_303_p N_noxref_7_M25_noxref_g ) capacitor c=0.00673971f \
 //x=10.605 //y=7.4 //x2=10.03 //y2=6.02
cc_452 ( N_noxref_2_M24_noxref_d N_noxref_7_M25_noxref_g ) capacitor \
 c=0.015318f //x=9.665 //y=5.02 //x2=10.03 //y2=6.02
cc_453 ( N_noxref_2_c_303_p N_noxref_7_M26_noxref_g ) capacitor c=0.00672952f \
 //x=10.605 //y=7.4 //x2=10.47 //y2=6.02
cc_454 ( N_noxref_2_c_262_n N_noxref_7_M26_noxref_g ) capacitor c=0.00864163f \
 //x=11.47 //y=7.4 //x2=10.47 //y2=6.02
cc_455 ( N_noxref_2_M26_noxref_d N_noxref_7_M26_noxref_g ) capacitor \
 c=0.0430452f //x=10.545 //y=5.02 //x2=10.47 //y2=6.02
cc_456 ( N_noxref_2_c_463_p N_noxref_7_M37_noxref_g ) capacitor c=0.00673971f \
 //x=20.595 //y=7.4 //x2=20.02 //y2=6.02
cc_457 ( N_noxref_2_M36_noxref_d N_noxref_7_M37_noxref_g ) capacitor \
 c=0.015318f //x=19.655 //y=5.02 //x2=20.02 //y2=6.02
cc_458 ( N_noxref_2_c_463_p N_noxref_7_M38_noxref_g ) capacitor c=0.00672952f \
 //x=20.595 //y=7.4 //x2=20.46 //y2=6.02
cc_459 ( N_noxref_2_c_259_n N_noxref_7_M38_noxref_g ) capacitor c=0.024326f \
 //x=21.09 //y=7.4 //x2=20.46 //y2=6.02
cc_460 ( N_noxref_2_M38_noxref_d N_noxref_7_M38_noxref_g ) capacitor \
 c=0.0430452f //x=20.535 //y=5.02 //x2=20.46 //y2=6.02
cc_461 ( N_noxref_2_c_258_n N_noxref_7_c_1466_n ) capacitor c=0.00757682f \
 //x=0.74 //y=7.4 //x2=1.385 //y2=4.79
cc_462 ( N_noxref_2_M13_noxref_s N_noxref_7_c_1466_n ) capacitor c=0.00445117f \
 //x=0.955 //y=5.02 //x2=1.385 //y2=4.79
cc_463 ( N_noxref_2_c_266_p N_noxref_7_M27_noxref_d ) capacitor c=0.00275225f \
 //x=21.09 //y=7.4 //x2=12.555 //y2=5.02
cc_464 ( N_noxref_2_c_314_p N_noxref_7_M27_noxref_d ) capacitor c=0.0140317f \
 //x=13.055 //y=7.4 //x2=12.555 //y2=5.02
cc_465 ( N_noxref_2_c_263_n N_noxref_7_M27_noxref_d ) capacitor c=6.94454e-19 \
 //x=14.8 //y=7.4 //x2=12.555 //y2=5.02
cc_466 ( N_noxref_2_M28_noxref_d N_noxref_7_M27_noxref_d ) capacitor \
 c=0.0664752f //x=12.995 //y=5.02 //x2=12.555 //y2=5.02
cc_467 ( N_noxref_2_c_266_p N_noxref_7_M29_noxref_d ) capacitor c=0.00285083f \
 //x=21.09 //y=7.4 //x2=13.435 //y2=5.02
cc_468 ( N_noxref_2_c_359_p N_noxref_7_M29_noxref_d ) capacitor c=0.0140984f \
 //x=13.935 //y=7.4 //x2=13.435 //y2=5.02
cc_469 ( N_noxref_2_c_263_n N_noxref_7_M29_noxref_d ) capacitor c=0.0120541f \
 //x=14.8 //y=7.4 //x2=13.435 //y2=5.02
cc_470 ( N_noxref_2_M27_noxref_s N_noxref_7_M29_noxref_d ) capacitor \
 c=0.00111971f //x=12.125 //y=5.02 //x2=13.435 //y2=5.02
cc_471 ( N_noxref_2_M28_noxref_d N_noxref_7_M29_noxref_d ) capacitor \
 c=0.0664752f //x=12.995 //y=5.02 //x2=13.435 //y2=5.02
cc_472 ( N_noxref_2_M30_noxref_d N_noxref_7_M29_noxref_d ) capacitor \
 c=0.0664752f //x=13.875 //y=5.02 //x2=13.435 //y2=5.02
cc_473 ( N_noxref_2_M31_noxref_s N_noxref_7_M29_noxref_d ) capacitor \
 c=4.54516e-19 //x=15.455 //y=5.02 //x2=13.435 //y2=5.02
cc_474 ( N_noxref_2_c_260_n N_noxref_10_c_1841_n ) capacitor c=4.47073e-19 \
 //x=4.81 //y=7.4 //x2=6.66 //y2=2.08
cc_475 ( N_noxref_2_c_261_n N_noxref_10_c_1841_n ) capacitor c=3.37458e-19 \
 //x=8.14 //y=7.4 //x2=6.66 //y2=2.08
cc_476 ( N_noxref_2_c_268_p N_noxref_10_M21_noxref_g ) capacitor c=0.00673971f \
 //x=7.275 //y=7.4 //x2=6.7 //y2=6.02
cc_477 ( N_noxref_2_M20_noxref_d N_noxref_10_M21_noxref_g ) capacitor \
 c=0.015318f //x=6.335 //y=5.02 //x2=6.7 //y2=6.02
cc_478 ( N_noxref_2_c_268_p N_noxref_10_M22_noxref_g ) capacitor c=0.00672952f \
 //x=7.275 //y=7.4 //x2=7.14 //y2=6.02
cc_479 ( N_noxref_2_c_261_n N_noxref_10_M22_noxref_g ) capacitor c=0.00864163f \
 //x=8.14 //y=7.4 //x2=7.14 //y2=6.02
cc_480 ( N_noxref_2_M22_noxref_d N_noxref_10_M22_noxref_g ) capacitor \
 c=0.0430452f //x=7.215 //y=5.02 //x2=7.14 //y2=6.02
cc_481 ( N_noxref_2_c_263_n N_noxref_14_c_2072_n ) capacitor c=9.06385e-19 \
 //x=14.8 //y=7.4 //x2=16.65 //y2=2.08
cc_482 ( N_noxref_2_c_264_n N_noxref_14_c_2072_n ) capacitor c=5.81514e-19 \
 //x=18.13 //y=7.4 //x2=16.65 //y2=2.08
cc_483 ( N_noxref_2_c_490_p N_noxref_14_M33_noxref_g ) capacitor c=0.00673971f \
 //x=17.265 //y=7.4 //x2=16.69 //y2=6.02
cc_484 ( N_noxref_2_M32_noxref_d N_noxref_14_M33_noxref_g ) capacitor \
 c=0.015318f //x=16.325 //y=5.02 //x2=16.69 //y2=6.02
cc_485 ( N_noxref_2_c_490_p N_noxref_14_M34_noxref_g ) capacitor c=0.00672952f \
 //x=17.265 //y=7.4 //x2=17.13 //y2=6.02
cc_486 ( N_noxref_2_c_264_n N_noxref_14_M34_noxref_g ) capacitor c=0.00864163f \
 //x=18.13 //y=7.4 //x2=17.13 //y2=6.02
cc_487 ( N_noxref_2_M34_noxref_d N_noxref_14_M34_noxref_g ) capacitor \
 c=0.0430452f //x=17.205 //y=5.02 //x2=17.13 //y2=6.02
cc_488 ( N_noxref_2_c_266_p N_noxref_15_c_2146_n ) capacitor c=0.00460134f \
 //x=21.09 //y=7.4 //x2=16.825 //y2=5.2
cc_489 ( N_noxref_2_c_384_p N_noxref_15_c_2146_n ) capacitor c=4.48705e-19 \
 //x=16.385 //y=7.4 //x2=16.825 //y2=5.2
cc_490 ( N_noxref_2_c_490_p N_noxref_15_c_2146_n ) capacitor c=4.48705e-19 \
 //x=17.265 //y=7.4 //x2=16.825 //y2=5.2
cc_491 ( N_noxref_2_M32_noxref_d N_noxref_15_c_2146_n ) capacitor c=0.0126924f \
 //x=16.325 //y=5.02 //x2=16.825 //y2=5.2
cc_492 ( N_noxref_2_c_263_n N_noxref_15_c_2150_n ) capacitor c=0.00985474f \
 //x=14.8 //y=7.4 //x2=16.115 //y2=5.2
cc_493 ( N_noxref_2_M31_noxref_s N_noxref_15_c_2150_n ) capacitor c=0.087833f \
 //x=15.455 //y=5.02 //x2=16.115 //y2=5.2
cc_494 ( N_noxref_2_c_266_p N_noxref_15_c_2152_n ) capacitor c=0.00307195f \
 //x=21.09 //y=7.4 //x2=17.305 //y2=5.2
cc_495 ( N_noxref_2_c_490_p N_noxref_15_c_2152_n ) capacitor c=7.73167e-19 \
 //x=17.265 //y=7.4 //x2=17.305 //y2=5.2
cc_496 ( N_noxref_2_M34_noxref_d N_noxref_15_c_2152_n ) capacitor c=0.0161518f \
 //x=17.205 //y=5.02 //x2=17.305 //y2=5.2
cc_497 ( N_noxref_2_M35_noxref_s N_noxref_15_c_2152_n ) capacitor \
 c=2.44532e-19 //x=18.785 //y=5.02 //x2=17.305 //y2=5.2
cc_498 ( N_noxref_2_c_263_n N_noxref_15_c_2142_n ) capacitor c=0.00151618f \
 //x=14.8 //y=7.4 //x2=17.39 //y2=5.115
cc_499 ( N_noxref_2_c_264_n N_noxref_15_c_2142_n ) capacitor c=0.0455537f \
 //x=18.13 //y=7.4 //x2=17.39 //y2=5.115
cc_500 ( N_noxref_2_c_266_p N_noxref_15_M31_noxref_d ) capacitor c=0.00285083f \
 //x=21.09 //y=7.4 //x2=15.885 //y2=5.02
cc_501 ( N_noxref_2_c_384_p N_noxref_15_M31_noxref_d ) capacitor c=0.0140984f \
 //x=16.385 //y=7.4 //x2=15.885 //y2=5.02
cc_502 ( N_noxref_2_c_264_n N_noxref_15_M31_noxref_d ) capacitor c=6.94454e-19 \
 //x=18.13 //y=7.4 //x2=15.885 //y2=5.02
cc_503 ( N_noxref_2_M32_noxref_d N_noxref_15_M31_noxref_d ) capacitor \
 c=0.0664752f //x=16.325 //y=5.02 //x2=15.885 //y2=5.02
cc_504 ( N_noxref_2_c_266_p N_noxref_15_M33_noxref_d ) capacitor c=0.00285083f \
 //x=21.09 //y=7.4 //x2=16.765 //y2=5.02
cc_505 ( N_noxref_2_c_490_p N_noxref_15_M33_noxref_d ) capacitor c=0.0140984f \
 //x=17.265 //y=7.4 //x2=16.765 //y2=5.02
cc_506 ( N_noxref_2_c_264_n N_noxref_15_M33_noxref_d ) capacitor c=0.0120541f \
 //x=18.13 //y=7.4 //x2=16.765 //y2=5.02
cc_507 ( N_noxref_2_M31_noxref_s N_noxref_15_M33_noxref_d ) capacitor \
 c=0.00111971f //x=15.455 //y=5.02 //x2=16.765 //y2=5.02
cc_508 ( N_noxref_2_M32_noxref_d N_noxref_15_M33_noxref_d ) capacitor \
 c=0.0664752f //x=16.325 //y=5.02 //x2=16.765 //y2=5.02
cc_509 ( N_noxref_2_M34_noxref_d N_noxref_15_M33_noxref_d ) capacitor \
 c=0.0664752f //x=17.205 //y=5.02 //x2=16.765 //y2=5.02
cc_510 ( N_noxref_2_M35_noxref_s N_noxref_15_M33_noxref_d ) capacitor \
 c=4.54516e-19 //x=18.785 //y=5.02 //x2=16.765 //y2=5.02
cc_511 ( N_noxref_2_c_266_p N_noxref_17_c_2265_n ) capacitor c=0.00126216f \
 //x=21.09 //y=7.4 //x2=19.24 //y2=2.08
cc_512 ( N_noxref_2_c_426_p N_noxref_17_c_2265_n ) capacitor c=2.87813e-19 \
 //x=19.715 //y=7.4 //x2=19.24 //y2=2.08
cc_513 ( N_noxref_2_c_264_n N_noxref_17_c_2265_n ) capacitor c=0.0160121f \
 //x=18.13 //y=7.4 //x2=19.24 //y2=2.08
cc_514 ( N_noxref_2_c_426_p N_noxref_17_M35_noxref_g ) capacitor c=0.00726866f \
 //x=19.715 //y=7.4 //x2=19.14 //y2=6.02
cc_515 ( N_noxref_2_M35_noxref_s N_noxref_17_M35_noxref_g ) capacitor \
 c=0.054195f //x=18.785 //y=5.02 //x2=19.14 //y2=6.02
cc_516 ( N_noxref_2_c_426_p N_noxref_17_M36_noxref_g ) capacitor c=0.00672952f \
 //x=19.715 //y=7.4 //x2=19.58 //y2=6.02
cc_517 ( N_noxref_2_M36_noxref_d N_noxref_17_M36_noxref_g ) capacitor \
 c=0.015318f //x=19.655 //y=5.02 //x2=19.58 //y2=6.02
cc_518 ( N_noxref_2_c_264_n N_noxref_17_c_2283_n ) capacitor c=0.0150435f \
 //x=18.13 //y=7.4 //x2=19.24 //y2=4.7
cc_519 ( N_noxref_2_c_266_p N_noxref_18_c_2330_n ) capacitor c=0.00459955f \
 //x=21.09 //y=7.4 //x2=20.155 //y2=5.2
cc_520 ( N_noxref_2_c_426_p N_noxref_18_c_2330_n ) capacitor c=4.48705e-19 \
 //x=19.715 //y=7.4 //x2=20.155 //y2=5.2
cc_521 ( N_noxref_2_c_463_p N_noxref_18_c_2330_n ) capacitor c=4.48693e-19 \
 //x=20.595 //y=7.4 //x2=20.155 //y2=5.2
cc_522 ( N_noxref_2_M36_noxref_d N_noxref_18_c_2330_n ) capacitor c=0.01269f \
 //x=19.655 //y=5.02 //x2=20.155 //y2=5.2
cc_523 ( N_noxref_2_c_264_n N_noxref_18_c_2334_n ) capacitor c=0.00985474f \
 //x=18.13 //y=7.4 //x2=19.445 //y2=5.2
cc_524 ( N_noxref_2_M35_noxref_s N_noxref_18_c_2334_n ) capacitor c=0.087833f \
 //x=18.785 //y=5.02 //x2=19.445 //y2=5.2
cc_525 ( N_noxref_2_c_266_p N_noxref_18_c_2336_n ) capacitor c=0.00445413f \
 //x=21.09 //y=7.4 //x2=20.635 //y2=5.2
cc_526 ( N_noxref_2_c_463_p N_noxref_18_c_2336_n ) capacitor c=7.21492e-19 \
 //x=20.595 //y=7.4 //x2=20.635 //y2=5.2
cc_527 ( N_noxref_2_M38_noxref_d N_noxref_18_c_2336_n ) capacitor c=0.0165872f \
 //x=20.535 //y=5.02 //x2=20.635 //y2=5.2
cc_528 ( N_noxref_2_c_259_n N_noxref_18_c_2326_n ) capacitor c=0.0466813f \
 //x=21.09 //y=7.4 //x2=20.72 //y2=5.115
cc_529 ( N_noxref_2_c_264_n N_noxref_18_c_2326_n ) capacitor c=0.00151618f \
 //x=18.13 //y=7.4 //x2=20.72 //y2=5.115
cc_530 ( N_noxref_2_c_266_p N_noxref_18_M35_noxref_d ) capacitor c=0.00285083f \
 //x=21.09 //y=7.4 //x2=19.215 //y2=5.02
cc_531 ( N_noxref_2_c_426_p N_noxref_18_M35_noxref_d ) capacitor c=0.0140984f \
 //x=19.715 //y=7.4 //x2=19.215 //y2=5.02
cc_532 ( N_noxref_2_c_259_n N_noxref_18_M35_noxref_d ) capacitor c=6.94454e-19 \
 //x=21.09 //y=7.4 //x2=19.215 //y2=5.02
cc_533 ( N_noxref_2_M36_noxref_d N_noxref_18_M35_noxref_d ) capacitor \
 c=0.0664752f //x=19.655 //y=5.02 //x2=19.215 //y2=5.02
cc_534 ( N_noxref_2_c_266_p N_noxref_18_M37_noxref_d ) capacitor c=0.00706239f \
 //x=21.09 //y=7.4 //x2=20.095 //y2=5.02
cc_535 ( N_noxref_2_c_463_p N_noxref_18_M37_noxref_d ) capacitor c=0.0138379f \
 //x=20.595 //y=7.4 //x2=20.095 //y2=5.02
cc_536 ( N_noxref_2_c_259_n N_noxref_18_M37_noxref_d ) capacitor c=0.0123189f \
 //x=21.09 //y=7.4 //x2=20.095 //y2=5.02
cc_537 ( N_noxref_2_M35_noxref_s N_noxref_18_M37_noxref_d ) capacitor \
 c=0.00111971f //x=18.785 //y=5.02 //x2=20.095 //y2=5.02
cc_538 ( N_noxref_2_M36_noxref_d N_noxref_18_M37_noxref_d ) capacitor \
 c=0.0664752f //x=19.655 //y=5.02 //x2=20.095 //y2=5.02
cc_539 ( N_noxref_2_M38_noxref_d N_noxref_18_M37_noxref_d ) capacitor \
 c=0.0664752f //x=20.535 //y=5.02 //x2=20.095 //y2=5.02
cc_540 ( N_noxref_3_c_553_n N_noxref_4_c_783_n ) capacitor c=0.011463f \
 //x=9.135 //y=3.33 //x2=10.845 //y2=3.33
cc_541 ( N_noxref_3_M24_noxref_g N_noxref_4_c_800_n ) capacitor c=0.0169521f \
 //x=9.59 //y=6.02 //x2=10.165 //y2=5.2
cc_542 ( N_noxref_3_c_561_n N_noxref_4_c_804_n ) capacitor c=0.00539951f \
 //x=9.25 //y=2.08 //x2=9.455 //y2=5.2
cc_543 ( N_noxref_3_M23_noxref_g N_noxref_4_c_804_n ) capacitor c=0.0177326f \
 //x=9.15 //y=6.02 //x2=9.455 //y2=5.2
cc_544 ( N_noxref_3_c_599_n N_noxref_4_c_804_n ) capacitor c=0.00581252f \
 //x=9.25 //y=4.7 //x2=9.455 //y2=5.2
cc_545 ( N_noxref_3_c_560_n N_noxref_4_c_785_n ) capacitor c=3.49822e-19 \
 //x=7.4 //y=3.33 //x2=10.73 //y2=3.33
cc_546 ( N_noxref_3_c_561_n N_noxref_4_c_785_n ) capacitor c=0.00318783f \
 //x=9.25 //y=2.08 //x2=10.73 //y2=3.33
cc_547 ( N_noxref_3_M24_noxref_g N_noxref_4_M23_noxref_d ) capacitor \
 c=0.0173476f //x=9.59 //y=6.02 //x2=9.225 //y2=5.02
cc_548 ( N_noxref_3_c_547_n N_noxref_5_c_932_n ) capacitor c=0.00360213f \
 //x=7.285 //y=3.33 //x2=13.205 //y2=4.44
cc_549 ( N_noxref_3_c_552_n N_noxref_5_c_932_n ) capacitor c=4.49102e-19 \
 //x=3.445 //y=3.33 //x2=13.205 //y2=4.44
cc_550 ( N_noxref_3_c_558_n N_noxref_5_c_932_n ) capacitor c=0.0200057f \
 //x=3.33 //y=2.08 //x2=13.205 //y2=4.44
cc_551 ( N_noxref_3_c_576_n N_noxref_5_c_932_n ) capacitor c=0.0185297f \
 //x=6.835 //y=5.2 //x2=13.205 //y2=4.44
cc_552 ( N_noxref_3_c_580_n N_noxref_5_c_932_n ) capacitor c=0.0181237f \
 //x=6.125 //y=5.2 //x2=13.205 //y2=4.44
cc_553 ( N_noxref_3_c_560_n N_noxref_5_c_932_n ) capacitor c=0.0208321f \
 //x=7.4 //y=3.33 //x2=13.205 //y2=4.44
cc_554 ( N_noxref_3_c_561_n N_noxref_5_c_932_n ) capacitor c=0.0198304f \
 //x=9.25 //y=2.08 //x2=13.205 //y2=4.44
cc_555 ( N_noxref_3_c_626_p N_noxref_5_c_932_n ) capacitor c=0.0111881f \
 //x=3.33 //y=4.7 //x2=13.205 //y2=4.44
cc_556 ( N_noxref_3_c_599_n N_noxref_5_c_932_n ) capacitor c=0.0107057f \
 //x=9.25 //y=4.7 //x2=13.205 //y2=4.44
cc_557 ( N_noxref_3_c_558_n N_noxref_5_c_950_n ) capacitor c=0.00153281f \
 //x=3.33 //y=2.08 //x2=2.335 //y2=4.44
cc_558 ( N_noxref_3_c_552_n N_noxref_5_c_929_n ) capacitor c=0.00526349f \
 //x=3.445 //y=3.33 //x2=2.22 //y2=2.08
cc_559 ( N_noxref_3_c_558_n N_noxref_5_c_929_n ) capacitor c=0.0511464f \
 //x=3.33 //y=2.08 //x2=2.22 //y2=2.08
cc_560 ( N_noxref_3_c_631_p N_noxref_5_c_929_n ) capacitor c=0.00228632f \
 //x=3.33 //y=2.08 //x2=2.22 //y2=2.08
cc_561 ( N_noxref_3_c_626_p N_noxref_5_c_929_n ) capacitor c=0.00218014f \
 //x=3.33 //y=4.7 //x2=2.22 //y2=2.08
cc_562 ( N_noxref_3_M17_noxref_g N_noxref_5_M15_noxref_g ) capacitor \
 c=0.0101598f //x=3.07 //y=6.02 //x2=2.19 //y2=6.02
cc_563 ( N_noxref_3_M17_noxref_g N_noxref_5_M16_noxref_g ) capacitor \
 c=0.0602553f //x=3.07 //y=6.02 //x2=2.63 //y2=6.02
cc_564 ( N_noxref_3_M18_noxref_g N_noxref_5_M16_noxref_g ) capacitor \
 c=0.0101598f //x=3.51 //y=6.02 //x2=2.63 //y2=6.02
cc_565 ( N_noxref_3_c_636_p N_noxref_5_c_981_n ) capacitor c=0.00456962f \
 //x=3.32 //y=0.915 //x2=2.31 //y2=0.91
cc_566 ( N_noxref_3_c_637_p N_noxref_5_c_982_n ) capacitor c=0.00438372f \
 //x=3.32 //y=1.26 //x2=2.31 //y2=1.22
cc_567 ( N_noxref_3_c_638_p N_noxref_5_c_983_n ) capacitor c=0.00438372f \
 //x=3.32 //y=1.57 //x2=2.31 //y2=1.45
cc_568 ( N_noxref_3_c_558_n N_noxref_5_c_984_n ) capacitor c=0.0023343f \
 //x=3.33 //y=2.08 //x2=2.31 //y2=1.915
cc_569 ( N_noxref_3_c_631_p N_noxref_5_c_984_n ) capacitor c=0.00933826f \
 //x=3.33 //y=2.08 //x2=2.31 //y2=1.915
cc_570 ( N_noxref_3_c_641_p N_noxref_5_c_984_n ) capacitor c=0.00438372f \
 //x=3.33 //y=1.915 //x2=2.31 //y2=1.915
cc_571 ( N_noxref_3_c_626_p N_noxref_5_c_987_n ) capacitor c=0.0611812f \
 //x=3.33 //y=4.7 //x2=2.555 //y2=4.79
cc_572 ( N_noxref_3_c_558_n N_noxref_5_c_988_n ) capacitor c=0.00142741f \
 //x=3.33 //y=2.08 //x2=2.22 //y2=4.7
cc_573 ( N_noxref_3_c_626_p N_noxref_5_c_988_n ) capacitor c=0.00487508f \
 //x=3.33 //y=4.7 //x2=2.22 //y2=4.7
cc_574 ( N_noxref_3_c_547_n N_noxref_6_c_1207_n ) capacitor c=0.146341f \
 //x=7.285 //y=3.33 //x2=5.805 //y2=3.7
cc_575 ( N_noxref_3_c_547_n N_noxref_6_c_1208_n ) capacitor c=0.0294746f \
 //x=7.285 //y=3.33 //x2=4.185 //y2=3.7
cc_576 ( N_noxref_3_c_558_n N_noxref_6_c_1208_n ) capacitor c=0.00687545f \
 //x=3.33 //y=2.08 //x2=4.185 //y2=3.7
cc_577 ( N_noxref_3_c_547_n N_noxref_6_c_1134_n ) capacitor c=0.108749f \
 //x=7.285 //y=3.33 //x2=15.795 //y2=3.7
cc_578 ( N_noxref_3_c_553_n N_noxref_6_c_1134_n ) capacitor c=0.175696f \
 //x=9.135 //y=3.33 //x2=15.795 //y2=3.7
cc_579 ( N_noxref_3_c_557_n N_noxref_6_c_1134_n ) capacitor c=0.0267668f \
 //x=7.515 //y=3.33 //x2=15.795 //y2=3.7
cc_580 ( N_noxref_3_c_560_n N_noxref_6_c_1134_n ) capacitor c=0.0206034f \
 //x=7.4 //y=3.33 //x2=15.795 //y2=3.7
cc_581 ( N_noxref_3_c_561_n N_noxref_6_c_1134_n ) capacitor c=0.0205831f \
 //x=9.25 //y=2.08 //x2=15.795 //y2=3.7
cc_582 ( N_noxref_3_c_547_n N_noxref_6_c_1215_n ) capacitor c=0.0266674f \
 //x=7.285 //y=3.33 //x2=6.035 //y2=3.7
cc_583 ( N_noxref_3_M17_noxref_g N_noxref_6_c_1167_n ) capacitor c=0.01736f \
 //x=3.07 //y=6.02 //x2=3.205 //y2=5.155
cc_584 ( N_noxref_3_M18_noxref_g N_noxref_6_c_1171_n ) capacitor c=0.0194981f \
 //x=3.51 //y=6.02 //x2=3.985 //y2=5.155
cc_585 ( N_noxref_3_c_626_p N_noxref_6_c_1171_n ) capacitor c=0.00201851f \
 //x=3.33 //y=4.7 //x2=3.985 //y2=5.155
cc_586 ( N_noxref_3_c_657_p N_noxref_6_c_1136_n ) capacitor c=0.00359704f \
 //x=3.695 //y=1.415 //x2=3.985 //y2=1.665
cc_587 ( N_noxref_3_c_658_p N_noxref_6_c_1136_n ) capacitor c=0.00457401f \
 //x=3.85 //y=1.26 //x2=3.985 //y2=1.665
cc_588 ( N_noxref_3_c_547_n N_noxref_6_c_1221_n ) capacitor c=0.00628992f \
 //x=7.285 //y=3.33 //x2=3.67 //y2=1.665
cc_589 ( N_noxref_3_c_547_n N_noxref_6_c_1175_n ) capacitor c=0.0260398f \
 //x=7.285 //y=3.33 //x2=4.07 //y2=3.7
cc_590 ( N_noxref_3_c_552_n N_noxref_6_c_1175_n ) capacitor c=0.00117715f \
 //x=3.445 //y=3.33 //x2=4.07 //y2=3.7
cc_591 ( N_noxref_3_c_558_n N_noxref_6_c_1175_n ) capacitor c=0.0831612f \
 //x=3.33 //y=2.08 //x2=4.07 //y2=3.7
cc_592 ( N_noxref_3_c_560_n N_noxref_6_c_1175_n ) capacitor c=3.52729e-19 \
 //x=7.4 //y=3.33 //x2=4.07 //y2=3.7
cc_593 ( N_noxref_3_c_631_p N_noxref_6_c_1175_n ) capacitor c=0.00877984f \
 //x=3.33 //y=2.08 //x2=4.07 //y2=3.7
cc_594 ( N_noxref_3_c_641_p N_noxref_6_c_1175_n ) capacitor c=0.00283672f \
 //x=3.33 //y=1.915 //x2=4.07 //y2=3.7
cc_595 ( N_noxref_3_c_626_p N_noxref_6_c_1175_n ) capacitor c=0.013693f \
 //x=3.33 //y=4.7 //x2=4.07 //y2=3.7
cc_596 ( N_noxref_3_c_547_n N_noxref_6_c_1137_n ) capacitor c=0.0257693f \
 //x=7.285 //y=3.33 //x2=5.92 //y2=2.08
cc_597 ( N_noxref_3_c_558_n N_noxref_6_c_1137_n ) capacitor c=9.66956e-19 \
 //x=3.33 //y=2.08 //x2=5.92 //y2=2.08
cc_598 ( N_noxref_3_c_580_n N_noxref_6_c_1137_n ) capacitor c=0.00521572f \
 //x=6.125 //y=5.2 //x2=5.92 //y2=2.08
cc_599 ( N_noxref_3_c_560_n N_noxref_6_c_1137_n ) capacitor c=0.00319084f \
 //x=7.4 //y=3.33 //x2=5.92 //y2=2.08
cc_600 ( N_noxref_3_c_558_n N_noxref_6_c_1233_n ) capacitor c=0.0171303f \
 //x=3.33 //y=2.08 //x2=3.29 //y2=5.155
cc_601 ( N_noxref_3_c_626_p N_noxref_6_c_1233_n ) capacitor c=0.00475601f \
 //x=3.33 //y=4.7 //x2=3.29 //y2=5.155
cc_602 ( N_noxref_3_c_580_n N_noxref_6_M19_noxref_g ) capacitor c=0.0177326f \
 //x=6.125 //y=5.2 //x2=5.82 //y2=6.02
cc_603 ( N_noxref_3_c_576_n N_noxref_6_M20_noxref_g ) capacitor c=0.0169521f \
 //x=6.835 //y=5.2 //x2=6.26 //y2=6.02
cc_604 ( N_noxref_3_M19_noxref_d N_noxref_6_M20_noxref_g ) capacitor \
 c=0.0173476f //x=5.895 //y=5.02 //x2=6.26 //y2=6.02
cc_605 ( N_noxref_3_c_580_n N_noxref_6_c_1190_n ) capacitor c=0.00581252f \
 //x=6.125 //y=5.2 //x2=5.92 //y2=4.7
cc_606 ( N_noxref_3_c_636_p N_noxref_6_M2_noxref_d ) capacitor c=0.00217566f \
 //x=3.32 //y=0.915 //x2=3.395 //y2=0.915
cc_607 ( N_noxref_3_c_637_p N_noxref_6_M2_noxref_d ) capacitor c=0.0034598f \
 //x=3.32 //y=1.26 //x2=3.395 //y2=0.915
cc_608 ( N_noxref_3_c_638_p N_noxref_6_M2_noxref_d ) capacitor c=0.00544291f \
 //x=3.32 //y=1.57 //x2=3.395 //y2=0.915
cc_609 ( N_noxref_3_c_680_p N_noxref_6_M2_noxref_d ) capacitor c=0.00241102f \
 //x=3.695 //y=0.76 //x2=3.395 //y2=0.915
cc_610 ( N_noxref_3_c_657_p N_noxref_6_M2_noxref_d ) capacitor c=0.0140297f \
 //x=3.695 //y=1.415 //x2=3.395 //y2=0.915
cc_611 ( N_noxref_3_c_682_p N_noxref_6_M2_noxref_d ) capacitor c=0.00219619f \
 //x=3.85 //y=0.915 //x2=3.395 //y2=0.915
cc_612 ( N_noxref_3_c_658_p N_noxref_6_M2_noxref_d ) capacitor c=0.00603828f \
 //x=3.85 //y=1.26 //x2=3.395 //y2=0.915
cc_613 ( N_noxref_3_c_641_p N_noxref_6_M2_noxref_d ) capacitor c=0.00661782f \
 //x=3.33 //y=1.915 //x2=3.395 //y2=0.915
cc_614 ( N_noxref_3_M17_noxref_g N_noxref_6_M17_noxref_d ) capacitor \
 c=0.0180032f //x=3.07 //y=6.02 //x2=3.145 //y2=5.02
cc_615 ( N_noxref_3_M18_noxref_g N_noxref_6_M17_noxref_d ) capacitor \
 c=0.0194246f //x=3.51 //y=6.02 //x2=3.145 //y2=5.02
cc_616 ( N_noxref_3_c_547_n N_noxref_7_c_1385_n ) capacitor c=0.0428508f \
 //x=7.285 //y=3.33 //x2=9.875 //y2=4.07
cc_617 ( N_noxref_3_c_552_n N_noxref_7_c_1385_n ) capacitor c=0.0135672f \
 //x=3.445 //y=3.33 //x2=9.875 //y2=4.07
cc_618 ( N_noxref_3_c_553_n N_noxref_7_c_1385_n ) capacitor c=0.0110241f \
 //x=9.135 //y=3.33 //x2=9.875 //y2=4.07
cc_619 ( N_noxref_3_c_557_n N_noxref_7_c_1385_n ) capacitor c=5.70661e-19 \
 //x=7.515 //y=3.33 //x2=9.875 //y2=4.07
cc_620 ( N_noxref_3_c_558_n N_noxref_7_c_1385_n ) capacitor c=0.0206302f \
 //x=3.33 //y=2.08 //x2=9.875 //y2=4.07
cc_621 ( N_noxref_3_c_560_n N_noxref_7_c_1385_n ) capacitor c=0.0181936f \
 //x=7.4 //y=3.33 //x2=9.875 //y2=4.07
cc_622 ( N_noxref_3_c_561_n N_noxref_7_c_1385_n ) capacitor c=0.0184765f \
 //x=9.25 //y=2.08 //x2=9.875 //y2=4.07
cc_623 ( N_noxref_3_c_561_n N_noxref_7_c_1486_n ) capacitor c=0.00179385f \
 //x=9.25 //y=2.08 //x2=10.105 //y2=4.07
cc_624 ( N_noxref_3_c_558_n N_noxref_7_c_1389_n ) capacitor c=0.00175117f \
 //x=3.33 //y=2.08 //x2=1.11 //y2=2.08
cc_625 ( N_noxref_3_c_561_n N_noxref_7_c_1488_n ) capacitor c=0.00400249f \
 //x=9.25 //y=2.08 //x2=9.99 //y2=4.535
cc_626 ( N_noxref_3_c_599_n N_noxref_7_c_1488_n ) capacitor c=0.00417994f \
 //x=9.25 //y=4.7 //x2=9.99 //y2=4.535
cc_627 ( N_noxref_3_c_553_n N_noxref_7_c_1390_n ) capacitor c=0.00318578f \
 //x=9.135 //y=3.33 //x2=9.99 //y2=2.08
cc_628 ( N_noxref_3_c_560_n N_noxref_7_c_1390_n ) capacitor c=9.69022e-19 \
 //x=7.4 //y=3.33 //x2=9.99 //y2=2.08
cc_629 ( N_noxref_3_c_561_n N_noxref_7_c_1390_n ) capacitor c=0.0794726f \
 //x=9.25 //y=2.08 //x2=9.99 //y2=2.08
cc_630 ( N_noxref_3_c_566_n N_noxref_7_c_1390_n ) capacitor c=0.00308814f \
 //x=9.055 //y=1.915 //x2=9.99 //y2=2.08
cc_631 ( N_noxref_3_M23_noxref_g N_noxref_7_M25_noxref_g ) capacitor \
 c=0.0104611f //x=9.15 //y=6.02 //x2=10.03 //y2=6.02
cc_632 ( N_noxref_3_M24_noxref_g N_noxref_7_M25_noxref_g ) capacitor \
 c=0.106811f //x=9.59 //y=6.02 //x2=10.03 //y2=6.02
cc_633 ( N_noxref_3_M24_noxref_g N_noxref_7_M26_noxref_g ) capacitor \
 c=0.0100341f //x=9.59 //y=6.02 //x2=10.47 //y2=6.02
cc_634 ( N_noxref_3_c_562_n N_noxref_7_c_1497_n ) capacitor c=4.86506e-19 \
 //x=9.055 //y=0.865 //x2=10.025 //y2=0.905
cc_635 ( N_noxref_3_c_564_n N_noxref_7_c_1497_n ) capacitor c=0.00152104f \
 //x=9.055 //y=1.21 //x2=10.025 //y2=0.905
cc_636 ( N_noxref_3_c_569_n N_noxref_7_c_1497_n ) capacitor c=0.0151475f \
 //x=9.585 //y=0.865 //x2=10.025 //y2=0.905
cc_637 ( N_noxref_3_c_565_n N_noxref_7_c_1500_n ) capacitor c=0.00109982f \
 //x=9.055 //y=1.52 //x2=10.025 //y2=1.25
cc_638 ( N_noxref_3_c_571_n N_noxref_7_c_1500_n ) capacitor c=0.0111064f \
 //x=9.585 //y=1.21 //x2=10.025 //y2=1.25
cc_639 ( N_noxref_3_c_565_n N_noxref_7_c_1502_n ) capacitor c=9.57794e-19 \
 //x=9.055 //y=1.52 //x2=10.025 //y2=1.56
cc_640 ( N_noxref_3_c_566_n N_noxref_7_c_1502_n ) capacitor c=0.00662747f \
 //x=9.055 //y=1.915 //x2=10.025 //y2=1.56
cc_641 ( N_noxref_3_c_571_n N_noxref_7_c_1502_n ) capacitor c=0.00862358f \
 //x=9.585 //y=1.21 //x2=10.025 //y2=1.56
cc_642 ( N_noxref_3_c_569_n N_noxref_7_c_1505_n ) capacitor c=0.00124821f \
 //x=9.585 //y=0.865 //x2=10.555 //y2=0.905
cc_643 ( N_noxref_3_c_571_n N_noxref_7_c_1506_n ) capacitor c=0.00200715f \
 //x=9.585 //y=1.21 //x2=10.555 //y2=1.25
cc_644 ( N_noxref_3_c_561_n N_noxref_7_c_1507_n ) capacitor c=0.00307062f \
 //x=9.25 //y=2.08 //x2=9.99 //y2=2.08
cc_645 ( N_noxref_3_c_566_n N_noxref_7_c_1507_n ) capacitor c=0.0179092f \
 //x=9.055 //y=1.915 //x2=9.99 //y2=2.08
cc_646 ( N_noxref_3_c_561_n N_noxref_7_c_1509_n ) capacitor c=0.00344981f \
 //x=9.25 //y=2.08 //x2=10.02 //y2=4.7
cc_647 ( N_noxref_3_c_599_n N_noxref_7_c_1509_n ) capacitor c=0.0293367f \
 //x=9.25 //y=4.7 //x2=10.02 //y2=4.7
cc_648 ( N_noxref_3_c_547_n N_noxref_9_c_1793_n ) capacitor c=2.45218e-19 \
 //x=7.285 //y=3.33 //x2=3.985 //y2=0.54
cc_649 ( N_noxref_3_c_558_n N_noxref_9_c_1793_n ) capacitor c=0.00208521f \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_650 ( N_noxref_3_c_636_p N_noxref_9_c_1793_n ) capacitor c=0.0194423f \
 //x=3.32 //y=0.915 //x2=3.985 //y2=0.54
cc_651 ( N_noxref_3_c_682_p N_noxref_9_c_1793_n ) capacitor c=0.00656458f \
 //x=3.85 //y=0.915 //x2=3.985 //y2=0.54
cc_652 ( N_noxref_3_c_631_p N_noxref_9_c_1793_n ) capacitor c=2.20712e-19 \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_653 ( N_noxref_3_c_637_p N_noxref_9_c_1807_n ) capacitor c=0.00538829f \
 //x=3.32 //y=1.26 //x2=3.1 //y2=0.995
cc_654 ( N_noxref_3_c_636_p N_noxref_9_M2_noxref_s ) capacitor c=0.00538829f \
 //x=3.32 //y=0.915 //x2=2.965 //y2=0.375
cc_655 ( N_noxref_3_c_638_p N_noxref_9_M2_noxref_s ) capacitor c=0.00538829f \
 //x=3.32 //y=1.57 //x2=2.965 //y2=0.375
cc_656 ( N_noxref_3_c_682_p N_noxref_9_M2_noxref_s ) capacitor c=0.0143002f \
 //x=3.85 //y=0.915 //x2=2.965 //y2=0.375
cc_657 ( N_noxref_3_c_658_p N_noxref_9_M2_noxref_s ) capacitor c=0.00290153f \
 //x=3.85 //y=1.26 //x2=2.965 //y2=0.375
cc_658 ( N_noxref_3_c_576_n N_noxref_10_c_1850_n ) capacitor c=0.0127164f \
 //x=6.835 //y=5.2 //x2=6.66 //y2=4.535
cc_659 ( N_noxref_3_c_560_n N_noxref_10_c_1850_n ) capacitor c=0.0101284f \
 //x=7.4 //y=3.33 //x2=6.66 //y2=4.535
cc_660 ( N_noxref_3_c_547_n N_noxref_10_c_1841_n ) capacitor c=0.0222863f \
 //x=7.285 //y=3.33 //x2=6.66 //y2=2.08
cc_661 ( N_noxref_3_c_557_n N_noxref_10_c_1841_n ) capacitor c=0.00117715f \
 //x=7.515 //y=3.33 //x2=6.66 //y2=2.08
cc_662 ( N_noxref_3_c_560_n N_noxref_10_c_1841_n ) capacitor c=0.0730419f \
 //x=7.4 //y=3.33 //x2=6.66 //y2=2.08
cc_663 ( N_noxref_3_c_561_n N_noxref_10_c_1841_n ) capacitor c=7.76771e-19 \
 //x=9.25 //y=2.08 //x2=6.66 //y2=2.08
cc_664 ( N_noxref_3_c_576_n N_noxref_10_M21_noxref_g ) capacitor c=0.0166421f \
 //x=6.835 //y=5.2 //x2=6.7 //y2=6.02
cc_665 ( N_noxref_3_M21_noxref_d N_noxref_10_M21_noxref_g ) capacitor \
 c=0.0173476f //x=6.775 //y=5.02 //x2=6.7 //y2=6.02
cc_666 ( N_noxref_3_c_582_n N_noxref_10_M22_noxref_g ) capacitor c=0.018922f \
 //x=7.315 //y=5.2 //x2=7.14 //y2=6.02
cc_667 ( N_noxref_3_M21_noxref_d N_noxref_10_M22_noxref_g ) capacitor \
 c=0.0179769f //x=6.775 //y=5.02 //x2=7.14 //y2=6.02
cc_668 ( N_noxref_3_M4_noxref_d N_noxref_10_c_1860_n ) capacitor c=0.00217566f \
 //x=6.77 //y=0.905 //x2=6.695 //y2=0.905
cc_669 ( N_noxref_3_M4_noxref_d N_noxref_10_c_1861_n ) capacitor c=0.0034598f \
 //x=6.77 //y=0.905 //x2=6.695 //y2=1.25
cc_670 ( N_noxref_3_M4_noxref_d N_noxref_10_c_1862_n ) capacitor c=0.0065582f \
 //x=6.77 //y=0.905 //x2=6.695 //y2=1.56
cc_671 ( N_noxref_3_c_560_n N_noxref_10_c_1863_n ) capacitor c=0.0142673f \
 //x=7.4 //y=3.33 //x2=7.065 //y2=4.79
cc_672 ( N_noxref_3_c_743_p N_noxref_10_c_1863_n ) capacitor c=0.00407665f \
 //x=6.92 //y=5.2 //x2=7.065 //y2=4.79
cc_673 ( N_noxref_3_M4_noxref_d N_noxref_10_c_1865_n ) capacitor c=0.00241102f \
 //x=6.77 //y=0.905 //x2=7.07 //y2=0.75
cc_674 ( N_noxref_3_c_559_n N_noxref_10_c_1866_n ) capacitor c=0.00359704f \
 //x=7.315 //y=1.655 //x2=7.07 //y2=1.405
cc_675 ( N_noxref_3_M4_noxref_d N_noxref_10_c_1866_n ) capacitor c=0.0138845f \
 //x=6.77 //y=0.905 //x2=7.07 //y2=1.405
cc_676 ( N_noxref_3_M4_noxref_d N_noxref_10_c_1868_n ) capacitor c=0.00132245f \
 //x=6.77 //y=0.905 //x2=7.225 //y2=0.905
cc_677 ( N_noxref_3_c_559_n N_noxref_10_c_1869_n ) capacitor c=0.00457401f \
 //x=7.315 //y=1.655 //x2=7.225 //y2=1.25
cc_678 ( N_noxref_3_M4_noxref_d N_noxref_10_c_1869_n ) capacitor c=0.00566463f \
 //x=6.77 //y=0.905 //x2=7.225 //y2=1.25
cc_679 ( N_noxref_3_c_560_n N_noxref_10_c_1871_n ) capacitor c=0.00877984f \
 //x=7.4 //y=3.33 //x2=6.66 //y2=2.08
cc_680 ( N_noxref_3_c_560_n N_noxref_10_c_1872_n ) capacitor c=0.00306024f \
 //x=7.4 //y=3.33 //x2=6.66 //y2=1.915
cc_681 ( N_noxref_3_M4_noxref_d N_noxref_10_c_1872_n ) capacitor c=0.00660593f \
 //x=6.77 //y=0.905 //x2=6.66 //y2=1.915
cc_682 ( N_noxref_3_c_576_n N_noxref_10_c_1874_n ) capacitor c=0.00346527f \
 //x=6.835 //y=5.2 //x2=6.69 //y2=4.7
cc_683 ( N_noxref_3_c_560_n N_noxref_10_c_1874_n ) capacitor c=0.00533692f \
 //x=7.4 //y=3.33 //x2=6.69 //y2=4.7
cc_684 ( N_noxref_3_c_547_n N_noxref_11_c_1933_n ) capacitor c=0.00241565f \
 //x=7.285 //y=3.33 //x2=5.505 //y2=1.495
cc_685 ( N_noxref_3_c_756_p N_noxref_11_c_1933_n ) capacitor c=3.15806e-19 \
 //x=7.045 //y=1.655 //x2=5.505 //y2=1.495
cc_686 ( N_noxref_3_c_547_n N_noxref_11_c_1914_n ) capacitor c=0.010299f \
 //x=7.285 //y=3.33 //x2=6.39 //y2=1.58
cc_687 ( N_noxref_3_c_547_n N_noxref_11_c_1921_n ) capacitor c=0.00241565f \
 //x=7.285 //y=3.33 //x2=6.475 //y2=1.495
cc_688 ( N_noxref_3_c_756_p N_noxref_11_c_1921_n ) capacitor c=0.020324f \
 //x=7.045 //y=1.655 //x2=6.475 //y2=1.495
cc_689 ( N_noxref_3_c_547_n N_noxref_11_c_1922_n ) capacitor c=7.52304e-19 \
 //x=7.285 //y=3.33 //x2=7.36 //y2=0.53
cc_690 ( N_noxref_3_c_559_n N_noxref_11_c_1922_n ) capacitor c=0.00465965f \
 //x=7.315 //y=1.655 //x2=7.36 //y2=0.53
cc_691 ( N_noxref_3_M4_noxref_d N_noxref_11_c_1922_n ) capacitor c=0.0117692f \
 //x=6.77 //y=0.905 //x2=7.36 //y2=0.53
cc_692 ( N_noxref_3_c_557_n N_noxref_11_M3_noxref_s ) capacitor c=3.47564e-19 \
 //x=7.515 //y=3.33 //x2=5.37 //y2=0.365
cc_693 ( N_noxref_3_c_559_n N_noxref_11_M3_noxref_s ) capacitor c=0.0141735f \
 //x=7.315 //y=1.655 //x2=5.37 //y2=0.365
cc_694 ( N_noxref_3_M4_noxref_d N_noxref_11_M3_noxref_s ) capacitor \
 c=0.0439476f //x=6.77 //y=0.905 //x2=5.37 //y2=0.365
cc_695 ( N_noxref_3_c_553_n N_noxref_12_c_1985_n ) capacitor c=0.00241565f \
 //x=9.135 //y=3.33 //x2=8.835 //y2=1.495
cc_696 ( N_noxref_3_c_559_n N_noxref_12_c_1985_n ) capacitor c=3.22188e-19 \
 //x=7.315 //y=1.655 //x2=8.835 //y2=1.495
cc_697 ( N_noxref_3_c_566_n N_noxref_12_c_1985_n ) capacitor c=0.0034165f \
 //x=9.055 //y=1.915 //x2=8.835 //y2=1.495
cc_698 ( N_noxref_3_c_553_n N_noxref_12_c_1966_n ) capacitor c=0.00649414f \
 //x=9.135 //y=3.33 //x2=9.72 //y2=1.58
cc_699 ( N_noxref_3_c_561_n N_noxref_12_c_1966_n ) capacitor c=0.011692f \
 //x=9.25 //y=2.08 //x2=9.72 //y2=1.58
cc_700 ( N_noxref_3_c_565_n N_noxref_12_c_1966_n ) capacitor c=0.00703567f \
 //x=9.055 //y=1.52 //x2=9.72 //y2=1.58
cc_701 ( N_noxref_3_c_566_n N_noxref_12_c_1966_n ) capacitor c=0.0203514f \
 //x=9.055 //y=1.915 //x2=9.72 //y2=1.58
cc_702 ( N_noxref_3_c_568_n N_noxref_12_c_1966_n ) capacitor c=0.00780629f \
 //x=9.43 //y=1.365 //x2=9.72 //y2=1.58
cc_703 ( N_noxref_3_c_571_n N_noxref_12_c_1966_n ) capacitor c=0.00339872f \
 //x=9.585 //y=1.21 //x2=9.72 //y2=1.58
cc_704 ( N_noxref_3_c_566_n N_noxref_12_c_1973_n ) capacitor c=6.71402e-19 \
 //x=9.055 //y=1.915 //x2=9.805 //y2=1.495
cc_705 ( N_noxref_3_c_562_n N_noxref_12_M5_noxref_s ) capacitor c=0.0326577f \
 //x=9.055 //y=0.865 //x2=8.7 //y2=0.365
cc_706 ( N_noxref_3_c_565_n N_noxref_12_M5_noxref_s ) capacitor c=3.48408e-19 \
 //x=9.055 //y=1.52 //x2=8.7 //y2=0.365
cc_707 ( N_noxref_3_c_569_n N_noxref_12_M5_noxref_s ) capacitor c=0.0120759f \
 //x=9.585 //y=0.865 //x2=8.7 //y2=0.365
cc_708 ( N_noxref_4_c_800_n N_noxref_5_c_932_n ) capacitor c=0.0185297f \
 //x=10.165 //y=5.2 //x2=13.205 //y2=4.44
cc_709 ( N_noxref_4_c_804_n N_noxref_5_c_932_n ) capacitor c=0.018142f \
 //x=9.455 //y=5.2 //x2=13.205 //y2=4.44
cc_710 ( N_noxref_4_c_785_n N_noxref_5_c_932_n ) capacitor c=0.0208321f \
 //x=10.73 //y=3.33 //x2=13.205 //y2=4.44
cc_711 ( N_noxref_4_c_786_n N_noxref_5_c_932_n ) capacitor c=0.0215137f \
 //x=12.58 //y=2.08 //x2=13.205 //y2=4.44
cc_712 ( N_noxref_4_c_819_n N_noxref_5_c_932_n ) capacitor c=0.0109968f \
 //x=12.58 //y=4.7 //x2=13.205 //y2=4.44
cc_713 ( N_noxref_4_c_786_n N_noxref_5_c_995_n ) capacitor c=0.00400249f \
 //x=12.58 //y=2.08 //x2=13.32 //y2=4.535
cc_714 ( N_noxref_4_c_819_n N_noxref_5_c_995_n ) capacitor c=0.00415951f \
 //x=12.58 //y=4.7 //x2=13.32 //y2=4.535
cc_715 ( N_noxref_4_c_779_n N_noxref_5_c_930_n ) capacitor c=0.00720056f \
 //x=12.465 //y=3.33 //x2=13.32 //y2=2.08
cc_716 ( N_noxref_4_c_785_n N_noxref_5_c_930_n ) capacitor c=0.00102338f \
 //x=10.73 //y=3.33 //x2=13.32 //y2=2.08
cc_717 ( N_noxref_4_c_786_n N_noxref_5_c_930_n ) capacitor c=0.0785565f \
 //x=12.58 //y=2.08 //x2=13.32 //y2=2.08
cc_718 ( N_noxref_4_c_791_n N_noxref_5_c_930_n ) capacitor c=0.00308814f \
 //x=12.385 //y=1.915 //x2=13.32 //y2=2.08
cc_719 ( N_noxref_4_M27_noxref_g N_noxref_5_M29_noxref_g ) capacitor \
 c=0.0104611f //x=12.48 //y=6.02 //x2=13.36 //y2=6.02
cc_720 ( N_noxref_4_M28_noxref_g N_noxref_5_M29_noxref_g ) capacitor \
 c=0.106811f //x=12.92 //y=6.02 //x2=13.36 //y2=6.02
cc_721 ( N_noxref_4_M28_noxref_g N_noxref_5_M30_noxref_g ) capacitor \
 c=0.0100341f //x=12.92 //y=6.02 //x2=13.8 //y2=6.02
cc_722 ( N_noxref_4_c_787_n N_noxref_5_c_1004_n ) capacitor c=4.86506e-19 \
 //x=12.385 //y=0.865 //x2=13.355 //y2=0.905
cc_723 ( N_noxref_4_c_789_n N_noxref_5_c_1004_n ) capacitor c=0.00152104f \
 //x=12.385 //y=1.21 //x2=13.355 //y2=0.905
cc_724 ( N_noxref_4_c_794_n N_noxref_5_c_1004_n ) capacitor c=0.0151475f \
 //x=12.915 //y=0.865 //x2=13.355 //y2=0.905
cc_725 ( N_noxref_4_c_790_n N_noxref_5_c_1007_n ) capacitor c=0.00109982f \
 //x=12.385 //y=1.52 //x2=13.355 //y2=1.25
cc_726 ( N_noxref_4_c_796_n N_noxref_5_c_1007_n ) capacitor c=0.0111064f \
 //x=12.915 //y=1.21 //x2=13.355 //y2=1.25
cc_727 ( N_noxref_4_c_790_n N_noxref_5_c_1009_n ) capacitor c=9.57794e-19 \
 //x=12.385 //y=1.52 //x2=13.355 //y2=1.56
cc_728 ( N_noxref_4_c_791_n N_noxref_5_c_1009_n ) capacitor c=0.00662747f \
 //x=12.385 //y=1.915 //x2=13.355 //y2=1.56
cc_729 ( N_noxref_4_c_796_n N_noxref_5_c_1009_n ) capacitor c=0.00862358f \
 //x=12.915 //y=1.21 //x2=13.355 //y2=1.56
cc_730 ( N_noxref_4_c_794_n N_noxref_5_c_1012_n ) capacitor c=0.00124821f \
 //x=12.915 //y=0.865 //x2=13.885 //y2=0.905
cc_731 ( N_noxref_4_c_796_n N_noxref_5_c_1013_n ) capacitor c=0.00200715f \
 //x=12.915 //y=1.21 //x2=13.885 //y2=1.25
cc_732 ( N_noxref_4_c_786_n N_noxref_5_c_1014_n ) capacitor c=0.00307062f \
 //x=12.58 //y=2.08 //x2=13.32 //y2=2.08
cc_733 ( N_noxref_4_c_791_n N_noxref_5_c_1014_n ) capacitor c=0.0179092f \
 //x=12.385 //y=1.915 //x2=13.32 //y2=2.08
cc_734 ( N_noxref_4_c_786_n N_noxref_5_c_1016_n ) capacitor c=0.00342116f \
 //x=12.58 //y=2.08 //x2=13.35 //y2=4.7
cc_735 ( N_noxref_4_c_819_n N_noxref_5_c_1016_n ) capacitor c=0.0292158f \
 //x=12.58 //y=4.7 //x2=13.35 //y2=4.7
cc_736 ( N_noxref_4_c_779_n N_noxref_6_c_1134_n ) capacitor c=0.175696f \
 //x=12.465 //y=3.33 //x2=15.795 //y2=3.7
cc_737 ( N_noxref_4_c_783_n N_noxref_6_c_1134_n ) capacitor c=0.0293967f \
 //x=10.845 //y=3.33 //x2=15.795 //y2=3.7
cc_738 ( N_noxref_4_c_869_p N_noxref_6_c_1134_n ) capacitor c=0.0037701f \
 //x=10.375 //y=1.655 //x2=15.795 //y2=3.7
cc_739 ( N_noxref_4_c_785_n N_noxref_6_c_1134_n ) capacitor c=0.0206034f \
 //x=10.73 //y=3.33 //x2=15.795 //y2=3.7
cc_740 ( N_noxref_4_c_786_n N_noxref_6_c_1134_n ) capacitor c=0.0205831f \
 //x=12.58 //y=2.08 //x2=15.795 //y2=3.7
cc_741 ( N_noxref_4_c_779_n N_noxref_7_c_1416_n ) capacitor c=0.0110241f \
 //x=12.465 //y=3.33 //x2=13.945 //y2=4.07
cc_742 ( N_noxref_4_c_783_n N_noxref_7_c_1416_n ) capacitor c=8.88358e-19 \
 //x=10.845 //y=3.33 //x2=13.945 //y2=4.07
cc_743 ( N_noxref_4_c_785_n N_noxref_7_c_1416_n ) capacitor c=0.0181936f \
 //x=10.73 //y=3.33 //x2=13.945 //y2=4.07
cc_744 ( N_noxref_4_c_786_n N_noxref_7_c_1416_n ) capacitor c=0.0184765f \
 //x=12.58 //y=2.08 //x2=13.945 //y2=4.07
cc_745 ( N_noxref_4_c_785_n N_noxref_7_c_1486_n ) capacitor c=0.00117715f \
 //x=10.73 //y=3.33 //x2=10.105 //y2=4.07
cc_746 ( N_noxref_4_c_800_n N_noxref_7_c_1488_n ) capacitor c=0.0127164f \
 //x=10.165 //y=5.2 //x2=9.99 //y2=4.535
cc_747 ( N_noxref_4_c_785_n N_noxref_7_c_1488_n ) capacitor c=0.0101319f \
 //x=10.73 //y=3.33 //x2=9.99 //y2=4.535
cc_748 ( N_noxref_4_c_783_n N_noxref_7_c_1390_n ) capacitor c=0.00329059f \
 //x=10.845 //y=3.33 //x2=9.99 //y2=2.08
cc_749 ( N_noxref_4_c_785_n N_noxref_7_c_1390_n ) capacitor c=0.0742673f \
 //x=10.73 //y=3.33 //x2=9.99 //y2=2.08
cc_750 ( N_noxref_4_c_786_n N_noxref_7_c_1390_n ) capacitor c=9.69022e-19 \
 //x=12.58 //y=2.08 //x2=9.99 //y2=2.08
cc_751 ( N_noxref_4_M28_noxref_g N_noxref_7_c_1438_n ) capacitor c=0.0169521f \
 //x=12.92 //y=6.02 //x2=13.495 //y2=5.2
cc_752 ( N_noxref_4_c_786_n N_noxref_7_c_1442_n ) capacitor c=0.00539951f \
 //x=12.58 //y=2.08 //x2=12.785 //y2=5.2
cc_753 ( N_noxref_4_M27_noxref_g N_noxref_7_c_1442_n ) capacitor c=0.0177326f \
 //x=12.48 //y=6.02 //x2=12.785 //y2=5.2
cc_754 ( N_noxref_4_c_819_n N_noxref_7_c_1442_n ) capacitor c=0.00581252f \
 //x=12.58 //y=4.7 //x2=12.785 //y2=5.2
cc_755 ( N_noxref_4_c_785_n N_noxref_7_c_1393_n ) capacitor c=3.49822e-19 \
 //x=10.73 //y=3.33 //x2=14.06 //y2=4.07
cc_756 ( N_noxref_4_c_786_n N_noxref_7_c_1393_n ) capacitor c=0.00389543f \
 //x=12.58 //y=2.08 //x2=14.06 //y2=4.07
cc_757 ( N_noxref_4_c_800_n N_noxref_7_M25_noxref_g ) capacitor c=0.0166421f \
 //x=10.165 //y=5.2 //x2=10.03 //y2=6.02
cc_758 ( N_noxref_4_M25_noxref_d N_noxref_7_M25_noxref_g ) capacitor \
 c=0.0173476f //x=10.105 //y=5.02 //x2=10.03 //y2=6.02
cc_759 ( N_noxref_4_c_806_n N_noxref_7_M26_noxref_g ) capacitor c=0.018922f \
 //x=10.645 //y=5.2 //x2=10.47 //y2=6.02
cc_760 ( N_noxref_4_M25_noxref_d N_noxref_7_M26_noxref_g ) capacitor \
 c=0.0179769f //x=10.105 //y=5.02 //x2=10.47 //y2=6.02
cc_761 ( N_noxref_4_M6_noxref_d N_noxref_7_c_1497_n ) capacitor c=0.00217566f \
 //x=10.1 //y=0.905 //x2=10.025 //y2=0.905
cc_762 ( N_noxref_4_M6_noxref_d N_noxref_7_c_1500_n ) capacitor c=0.0034598f \
 //x=10.1 //y=0.905 //x2=10.025 //y2=1.25
cc_763 ( N_noxref_4_M6_noxref_d N_noxref_7_c_1502_n ) capacitor c=0.0065582f \
 //x=10.1 //y=0.905 //x2=10.025 //y2=1.56
cc_764 ( N_noxref_4_c_785_n N_noxref_7_c_1534_n ) capacitor c=0.0142673f \
 //x=10.73 //y=3.33 //x2=10.395 //y2=4.79
cc_765 ( N_noxref_4_c_896_p N_noxref_7_c_1534_n ) capacitor c=0.00407665f \
 //x=10.25 //y=5.2 //x2=10.395 //y2=4.79
cc_766 ( N_noxref_4_M6_noxref_d N_noxref_7_c_1536_n ) capacitor c=0.00241102f \
 //x=10.1 //y=0.905 //x2=10.4 //y2=0.75
cc_767 ( N_noxref_4_c_784_n N_noxref_7_c_1537_n ) capacitor c=0.00359704f \
 //x=10.645 //y=1.655 //x2=10.4 //y2=1.405
cc_768 ( N_noxref_4_M6_noxref_d N_noxref_7_c_1537_n ) capacitor c=0.0138845f \
 //x=10.1 //y=0.905 //x2=10.4 //y2=1.405
cc_769 ( N_noxref_4_M6_noxref_d N_noxref_7_c_1505_n ) capacitor c=0.00132245f \
 //x=10.1 //y=0.905 //x2=10.555 //y2=0.905
cc_770 ( N_noxref_4_c_784_n N_noxref_7_c_1506_n ) capacitor c=0.00457401f \
 //x=10.645 //y=1.655 //x2=10.555 //y2=1.25
cc_771 ( N_noxref_4_M6_noxref_d N_noxref_7_c_1506_n ) capacitor c=0.00566463f \
 //x=10.1 //y=0.905 //x2=10.555 //y2=1.25
cc_772 ( N_noxref_4_c_785_n N_noxref_7_c_1507_n ) capacitor c=0.00877984f \
 //x=10.73 //y=3.33 //x2=9.99 //y2=2.08
cc_773 ( N_noxref_4_c_785_n N_noxref_7_c_1543_n ) capacitor c=0.00306024f \
 //x=10.73 //y=3.33 //x2=9.99 //y2=1.915
cc_774 ( N_noxref_4_M6_noxref_d N_noxref_7_c_1543_n ) capacitor c=0.00660593f \
 //x=10.1 //y=0.905 //x2=9.99 //y2=1.915
cc_775 ( N_noxref_4_c_800_n N_noxref_7_c_1509_n ) capacitor c=0.00346527f \
 //x=10.165 //y=5.2 //x2=10.02 //y2=4.7
cc_776 ( N_noxref_4_c_785_n N_noxref_7_c_1509_n ) capacitor c=0.00517969f \
 //x=10.73 //y=3.33 //x2=10.02 //y2=4.7
cc_777 ( N_noxref_4_M28_noxref_g N_noxref_7_M27_noxref_d ) capacitor \
 c=0.0173476f //x=12.92 //y=6.02 //x2=12.555 //y2=5.02
cc_778 ( N_noxref_4_c_869_p N_noxref_12_c_1985_n ) capacitor c=3.15806e-19 \
 //x=10.375 //y=1.655 //x2=8.835 //y2=1.495
cc_779 ( N_noxref_4_c_869_p N_noxref_12_c_1973_n ) capacitor c=0.0203424f \
 //x=10.375 //y=1.655 //x2=9.805 //y2=1.495
cc_780 ( N_noxref_4_c_784_n N_noxref_12_c_1974_n ) capacitor c=0.0046686f \
 //x=10.645 //y=1.655 //x2=10.69 //y2=0.53
cc_781 ( N_noxref_4_M6_noxref_d N_noxref_12_c_1974_n ) capacitor c=0.0117932f \
 //x=10.1 //y=0.905 //x2=10.69 //y2=0.53
cc_782 ( N_noxref_4_c_783_n N_noxref_12_M5_noxref_s ) capacitor c=3.47564e-19 \
 //x=10.845 //y=3.33 //x2=8.7 //y2=0.365
cc_783 ( N_noxref_4_c_784_n N_noxref_12_M5_noxref_s ) capacitor c=0.0141735f \
 //x=10.645 //y=1.655 //x2=8.7 //y2=0.365
cc_784 ( N_noxref_4_M6_noxref_d N_noxref_12_M5_noxref_s ) capacitor \
 c=0.043966f //x=10.1 //y=0.905 //x2=8.7 //y2=0.365
cc_785 ( N_noxref_4_c_779_n N_noxref_13_c_2038_n ) capacitor c=0.00241565f \
 //x=12.465 //y=3.33 //x2=12.165 //y2=1.495
cc_786 ( N_noxref_4_c_784_n N_noxref_13_c_2038_n ) capacitor c=3.22188e-19 \
 //x=10.645 //y=1.655 //x2=12.165 //y2=1.495
cc_787 ( N_noxref_4_c_791_n N_noxref_13_c_2038_n ) capacitor c=0.0034165f \
 //x=12.385 //y=1.915 //x2=12.165 //y2=1.495
cc_788 ( N_noxref_4_c_779_n N_noxref_13_c_2019_n ) capacitor c=0.00649414f \
 //x=12.465 //y=3.33 //x2=13.05 //y2=1.58
cc_789 ( N_noxref_4_c_786_n N_noxref_13_c_2019_n ) capacitor c=0.011692f \
 //x=12.58 //y=2.08 //x2=13.05 //y2=1.58
cc_790 ( N_noxref_4_c_790_n N_noxref_13_c_2019_n ) capacitor c=0.00703567f \
 //x=12.385 //y=1.52 //x2=13.05 //y2=1.58
cc_791 ( N_noxref_4_c_791_n N_noxref_13_c_2019_n ) capacitor c=0.0203514f \
 //x=12.385 //y=1.915 //x2=13.05 //y2=1.58
cc_792 ( N_noxref_4_c_793_n N_noxref_13_c_2019_n ) capacitor c=0.00780629f \
 //x=12.76 //y=1.365 //x2=13.05 //y2=1.58
cc_793 ( N_noxref_4_c_796_n N_noxref_13_c_2019_n ) capacitor c=0.00339872f \
 //x=12.915 //y=1.21 //x2=13.05 //y2=1.58
cc_794 ( N_noxref_4_c_791_n N_noxref_13_c_2026_n ) capacitor c=6.71402e-19 \
 //x=12.385 //y=1.915 //x2=13.135 //y2=1.495
cc_795 ( N_noxref_4_c_787_n N_noxref_13_M7_noxref_s ) capacitor c=0.0326577f \
 //x=12.385 //y=0.865 //x2=12.03 //y2=0.365
cc_796 ( N_noxref_4_c_790_n N_noxref_13_M7_noxref_s ) capacitor c=3.48408e-19 \
 //x=12.385 //y=1.52 //x2=12.03 //y2=0.365
cc_797 ( N_noxref_4_c_794_n N_noxref_13_M7_noxref_s ) capacitor c=0.0120759f \
 //x=12.915 //y=0.865 //x2=12.03 //y2=0.365
cc_798 ( N_noxref_5_c_932_n N_noxref_6_c_1207_n ) capacitor c=0.00940379f \
 //x=13.205 //y=4.44 //x2=5.805 //y2=3.7
cc_799 ( N_noxref_5_c_932_n N_noxref_6_c_1208_n ) capacitor c=7.95009e-19 \
 //x=13.205 //y=4.44 //x2=4.185 //y2=3.7
cc_800 ( N_noxref_5_c_932_n N_noxref_6_c_1134_n ) capacitor c=0.0492712f \
 //x=13.205 //y=4.44 //x2=15.795 //y2=3.7
cc_801 ( N_noxref_5_c_930_n N_noxref_6_c_1134_n ) capacitor c=0.0225527f \
 //x=13.32 //y=2.08 //x2=15.795 //y2=3.7
cc_802 ( N_noxref_5_c_932_n N_noxref_6_c_1215_n ) capacitor c=6.59192e-19 \
 //x=13.205 //y=4.44 //x2=6.035 //y2=3.7
cc_803 ( N_noxref_5_c_950_n N_noxref_6_c_1161_n ) capacitor c=0.00330099f \
 //x=2.335 //y=4.44 //x2=2.325 //y2=5.155
cc_804 ( N_noxref_5_c_929_n N_noxref_6_c_1161_n ) capacitor c=0.014564f \
 //x=2.22 //y=2.08 //x2=2.325 //y2=5.155
cc_805 ( N_noxref_5_M15_noxref_g N_noxref_6_c_1161_n ) capacitor c=0.016514f \
 //x=2.19 //y=6.02 //x2=2.325 //y2=5.155
cc_806 ( N_noxref_5_c_988_n N_noxref_6_c_1161_n ) capacitor c=0.00322046f \
 //x=2.22 //y=4.7 //x2=2.325 //y2=5.155
cc_807 ( N_noxref_5_M16_noxref_g N_noxref_6_c_1167_n ) capacitor c=0.01736f \
 //x=2.63 //y=6.02 //x2=3.205 //y2=5.155
cc_808 ( N_noxref_5_c_932_n N_noxref_6_c_1171_n ) capacitor c=0.0183122f \
 //x=13.205 //y=4.44 //x2=3.985 //y2=5.155
cc_809 ( N_noxref_5_c_932_n N_noxref_6_c_1175_n ) capacitor c=0.0210274f \
 //x=13.205 //y=4.44 //x2=4.07 //y2=3.7
cc_810 ( N_noxref_5_c_929_n N_noxref_6_c_1175_n ) capacitor c=0.00319363f \
 //x=2.22 //y=2.08 //x2=4.07 //y2=3.7
cc_811 ( N_noxref_5_c_932_n N_noxref_6_c_1137_n ) capacitor c=0.0198304f \
 //x=13.205 //y=4.44 //x2=5.92 //y2=2.08
cc_812 ( N_noxref_5_c_930_n N_noxref_6_c_1138_n ) capacitor c=0.00101176f \
 //x=13.32 //y=2.08 //x2=15.91 //y2=2.08
cc_813 ( N_noxref_5_c_932_n N_noxref_6_c_1269_n ) capacitor c=0.0311227f \
 //x=13.205 //y=4.44 //x2=2.41 //y2=5.155
cc_814 ( N_noxref_5_c_987_n N_noxref_6_c_1269_n ) capacitor c=0.00426767f \
 //x=2.555 //y=4.79 //x2=2.41 //y2=5.155
cc_815 ( N_noxref_5_c_932_n N_noxref_6_c_1190_n ) capacitor c=0.0107057f \
 //x=13.205 //y=4.44 //x2=5.92 //y2=4.7
cc_816 ( N_noxref_5_M15_noxref_g N_noxref_6_M15_noxref_d ) capacitor \
 c=0.0180032f //x=2.19 //y=6.02 //x2=2.265 //y2=5.02
cc_817 ( N_noxref_5_M16_noxref_g N_noxref_6_M15_noxref_d ) capacitor \
 c=0.0180032f //x=2.63 //y=6.02 //x2=2.265 //y2=5.02
cc_818 ( N_noxref_5_c_932_n N_noxref_7_c_1385_n ) capacitor c=0.656956f \
 //x=13.205 //y=4.44 //x2=9.875 //y2=4.07
cc_819 ( N_noxref_5_c_950_n N_noxref_7_c_1385_n ) capacitor c=0.0291328f \
 //x=2.335 //y=4.44 //x2=9.875 //y2=4.07
cc_820 ( N_noxref_5_c_929_n N_noxref_7_c_1385_n ) capacitor c=0.0265867f \
 //x=2.22 //y=2.08 //x2=9.875 //y2=4.07
cc_821 ( N_noxref_5_c_988_n N_noxref_7_c_1385_n ) capacitor c=6.38735e-19 \
 //x=2.22 //y=4.7 //x2=9.875 //y2=4.07
cc_822 ( N_noxref_5_c_929_n N_noxref_7_c_1386_n ) capacitor c=0.00128547f \
 //x=2.22 //y=2.08 //x2=1.225 //y2=4.07
cc_823 ( N_noxref_5_c_932_n N_noxref_7_c_1416_n ) capacitor c=0.300301f \
 //x=13.205 //y=4.44 //x2=13.945 //y2=4.07
cc_824 ( N_noxref_5_c_930_n N_noxref_7_c_1416_n ) capacitor c=0.0187718f \
 //x=13.32 //y=2.08 //x2=13.945 //y2=4.07
cc_825 ( N_noxref_5_c_1045_p N_noxref_7_c_1416_n ) capacitor c=0.00756255f \
 //x=13.725 //y=4.79 //x2=13.945 //y2=4.07
cc_826 ( N_noxref_5_c_1016_n N_noxref_7_c_1416_n ) capacitor c=4.6185e-19 \
 //x=13.35 //y=4.7 //x2=13.945 //y2=4.07
cc_827 ( N_noxref_5_c_932_n N_noxref_7_c_1486_n ) capacitor c=0.0263375f \
 //x=13.205 //y=4.44 //x2=10.105 //y2=4.07
cc_828 ( N_noxref_5_c_930_n N_noxref_7_c_1430_n ) capacitor c=0.00117715f \
 //x=13.32 //y=2.08 //x2=14.175 //y2=4.07
cc_829 ( N_noxref_5_c_950_n N_noxref_7_c_1389_n ) capacitor c=0.00551083f \
 //x=2.335 //y=4.44 //x2=1.11 //y2=2.08
cc_830 ( N_noxref_5_c_929_n N_noxref_7_c_1389_n ) capacitor c=0.0535714f \
 //x=2.22 //y=2.08 //x2=1.11 //y2=2.08
cc_831 ( N_noxref_5_c_984_n N_noxref_7_c_1389_n ) capacitor c=0.00231304f \
 //x=2.31 //y=1.915 //x2=1.11 //y2=2.08
cc_832 ( N_noxref_5_c_988_n N_noxref_7_c_1389_n ) capacitor c=0.00183762f \
 //x=2.22 //y=4.7 //x2=1.11 //y2=2.08
cc_833 ( N_noxref_5_c_932_n N_noxref_7_c_1488_n ) capacitor c=0.0016972f \
 //x=13.205 //y=4.44 //x2=9.99 //y2=4.535
cc_834 ( N_noxref_5_c_932_n N_noxref_7_c_1390_n ) capacitor c=0.0207534f \
 //x=13.205 //y=4.44 //x2=9.99 //y2=2.08
cc_835 ( N_noxref_5_c_932_n N_noxref_7_c_1438_n ) capacitor c=0.00325337f \
 //x=13.205 //y=4.44 //x2=13.495 //y2=5.2
cc_836 ( N_noxref_5_c_995_n N_noxref_7_c_1438_n ) capacitor c=0.0126416f \
 //x=13.32 //y=4.535 //x2=13.495 //y2=5.2
cc_837 ( N_noxref_5_c_930_n N_noxref_7_c_1438_n ) capacitor c=3.74769e-19 \
 //x=13.32 //y=2.08 //x2=13.495 //y2=5.2
cc_838 ( N_noxref_5_M29_noxref_g N_noxref_7_c_1438_n ) capacitor c=0.0166421f \
 //x=13.36 //y=6.02 //x2=13.495 //y2=5.2
cc_839 ( N_noxref_5_c_1016_n N_noxref_7_c_1438_n ) capacitor c=0.00346519f \
 //x=13.35 //y=4.7 //x2=13.495 //y2=5.2
cc_840 ( N_noxref_5_c_932_n N_noxref_7_c_1442_n ) capacitor c=0.0172877f \
 //x=13.205 //y=4.44 //x2=12.785 //y2=5.2
cc_841 ( N_noxref_5_M30_noxref_g N_noxref_7_c_1444_n ) capacitor c=0.0199348f \
 //x=13.8 //y=6.02 //x2=13.975 //y2=5.2
cc_842 ( N_noxref_5_c_1062_p N_noxref_7_c_1392_n ) capacitor c=0.00359704f \
 //x=13.73 //y=1.405 //x2=13.975 //y2=1.655
cc_843 ( N_noxref_5_c_1013_n N_noxref_7_c_1392_n ) capacitor c=0.00457401f \
 //x=13.885 //y=1.25 //x2=13.975 //y2=1.655
cc_844 ( N_noxref_5_c_932_n N_noxref_7_c_1393_n ) capacitor c=0.00707546f \
 //x=13.205 //y=4.44 //x2=14.06 //y2=4.07
cc_845 ( N_noxref_5_c_995_n N_noxref_7_c_1393_n ) capacitor c=0.00923416f \
 //x=13.32 //y=4.535 //x2=14.06 //y2=4.07
cc_846 ( N_noxref_5_c_930_n N_noxref_7_c_1393_n ) capacitor c=0.0757812f \
 //x=13.32 //y=2.08 //x2=14.06 //y2=4.07
cc_847 ( N_noxref_5_c_1045_p N_noxref_7_c_1393_n ) capacitor c=0.0142673f \
 //x=13.725 //y=4.79 //x2=14.06 //y2=4.07
cc_848 ( N_noxref_5_c_1014_n N_noxref_7_c_1393_n ) capacitor c=0.00877984f \
 //x=13.32 //y=2.08 //x2=14.06 //y2=4.07
cc_849 ( N_noxref_5_c_1069_p N_noxref_7_c_1393_n ) capacitor c=0.00306024f \
 //x=13.32 //y=1.915 //x2=14.06 //y2=4.07
cc_850 ( N_noxref_5_c_1016_n N_noxref_7_c_1393_n ) capacitor c=0.00518077f \
 //x=13.35 //y=4.7 //x2=14.06 //y2=4.07
cc_851 ( N_noxref_5_c_1045_p N_noxref_7_c_1581_n ) capacitor c=0.00408717f \
 //x=13.725 //y=4.79 //x2=13.58 //y2=5.2
cc_852 ( N_noxref_5_M15_noxref_g N_noxref_7_M13_noxref_g ) capacitor \
 c=0.0105869f //x=2.19 //y=6.02 //x2=1.31 //y2=6.02
cc_853 ( N_noxref_5_M15_noxref_g N_noxref_7_M14_noxref_g ) capacitor \
 c=0.10632f //x=2.19 //y=6.02 //x2=1.75 //y2=6.02
cc_854 ( N_noxref_5_M16_noxref_g N_noxref_7_M14_noxref_g ) capacitor \
 c=0.0101598f //x=2.63 //y=6.02 //x2=1.75 //y2=6.02
cc_855 ( N_noxref_5_c_1075_p N_noxref_7_c_1396_n ) capacitor c=5.72482e-19 \
 //x=1.785 //y=0.91 //x2=0.81 //y2=0.875
cc_856 ( N_noxref_5_c_1075_p N_noxref_7_c_1398_n ) capacitor c=0.00149976f \
 //x=1.785 //y=0.91 //x2=0.81 //y2=1.22
cc_857 ( N_noxref_5_c_1077_p N_noxref_7_c_1399_n ) capacitor c=0.00111227f \
 //x=1.785 //y=1.22 //x2=0.81 //y2=1.53
cc_858 ( N_noxref_5_c_929_n N_noxref_7_c_1400_n ) capacitor c=0.00238338f \
 //x=2.22 //y=2.08 //x2=0.81 //y2=1.915
cc_859 ( N_noxref_5_c_984_n N_noxref_7_c_1400_n ) capacitor c=0.00964411f \
 //x=2.31 //y=1.915 //x2=0.81 //y2=1.915
cc_860 ( N_noxref_5_c_1075_p N_noxref_7_c_1403_n ) capacitor c=0.0160123f \
 //x=1.785 //y=0.91 //x2=1.34 //y2=0.875
cc_861 ( N_noxref_5_c_981_n N_noxref_7_c_1403_n ) capacitor c=0.00103227f \
 //x=2.31 //y=0.91 //x2=1.34 //y2=0.875
cc_862 ( N_noxref_5_c_1077_p N_noxref_7_c_1405_n ) capacitor c=0.0124075f \
 //x=1.785 //y=1.22 //x2=1.34 //y2=1.22
cc_863 ( N_noxref_5_c_982_n N_noxref_7_c_1405_n ) capacitor c=0.0010154f \
 //x=2.31 //y=1.22 //x2=1.34 //y2=1.22
cc_864 ( N_noxref_5_c_983_n N_noxref_7_c_1405_n ) capacitor c=9.23422e-19 \
 //x=2.31 //y=1.45 //x2=1.34 //y2=1.22
cc_865 ( N_noxref_5_c_929_n N_noxref_7_c_1595_n ) capacitor c=0.00147352f \
 //x=2.22 //y=2.08 //x2=1.675 //y2=4.79
cc_866 ( N_noxref_5_c_988_n N_noxref_7_c_1595_n ) capacitor c=0.0168581f \
 //x=2.22 //y=4.7 //x2=1.675 //y2=4.79
cc_867 ( N_noxref_5_c_929_n N_noxref_7_c_1466_n ) capacitor c=0.00141297f \
 //x=2.22 //y=2.08 //x2=1.385 //y2=4.79
cc_868 ( N_noxref_5_c_988_n N_noxref_7_c_1466_n ) capacitor c=0.00484466f \
 //x=2.22 //y=4.7 //x2=1.385 //y2=4.79
cc_869 ( N_noxref_5_c_932_n N_noxref_7_c_1534_n ) capacitor c=0.00960248f \
 //x=13.205 //y=4.44 //x2=10.395 //y2=4.79
cc_870 ( N_noxref_5_c_932_n N_noxref_7_c_1509_n ) capacitor c=0.00203982f \
 //x=13.205 //y=4.44 //x2=10.02 //y2=4.7
cc_871 ( N_noxref_5_c_1004_n N_noxref_7_M8_noxref_d ) capacitor c=0.00217566f \
 //x=13.355 //y=0.905 //x2=13.43 //y2=0.905
cc_872 ( N_noxref_5_c_1007_n N_noxref_7_M8_noxref_d ) capacitor c=0.0034598f \
 //x=13.355 //y=1.25 //x2=13.43 //y2=0.905
cc_873 ( N_noxref_5_c_1009_n N_noxref_7_M8_noxref_d ) capacitor c=0.0065582f \
 //x=13.355 //y=1.56 //x2=13.43 //y2=0.905
cc_874 ( N_noxref_5_c_1094_p N_noxref_7_M8_noxref_d ) capacitor c=0.00241102f \
 //x=13.73 //y=0.75 //x2=13.43 //y2=0.905
cc_875 ( N_noxref_5_c_1062_p N_noxref_7_M8_noxref_d ) capacitor c=0.0138845f \
 //x=13.73 //y=1.405 //x2=13.43 //y2=0.905
cc_876 ( N_noxref_5_c_1012_n N_noxref_7_M8_noxref_d ) capacitor c=0.00132245f \
 //x=13.885 //y=0.905 //x2=13.43 //y2=0.905
cc_877 ( N_noxref_5_c_1013_n N_noxref_7_M8_noxref_d ) capacitor c=0.00566463f \
 //x=13.885 //y=1.25 //x2=13.43 //y2=0.905
cc_878 ( N_noxref_5_c_1069_p N_noxref_7_M8_noxref_d ) capacitor c=0.00660593f \
 //x=13.32 //y=1.915 //x2=13.43 //y2=0.905
cc_879 ( N_noxref_5_M29_noxref_g N_noxref_7_M29_noxref_d ) capacitor \
 c=0.0173476f //x=13.36 //y=6.02 //x2=13.435 //y2=5.02
cc_880 ( N_noxref_5_M30_noxref_g N_noxref_7_M29_noxref_d ) capacitor \
 c=0.0179769f //x=13.8 //y=6.02 //x2=13.435 //y2=5.02
cc_881 ( N_noxref_5_c_1075_p N_noxref_8_c_1748_n ) capacitor c=0.0167228f \
 //x=1.785 //y=0.91 //x2=2.445 //y2=0.54
cc_882 ( N_noxref_5_c_981_n N_noxref_8_c_1748_n ) capacitor c=0.00534519f \
 //x=2.31 //y=0.91 //x2=2.445 //y2=0.54
cc_883 ( N_noxref_5_c_929_n N_noxref_8_c_1759_n ) capacitor c=0.012357f \
 //x=2.22 //y=2.08 //x2=2.445 //y2=1.59
cc_884 ( N_noxref_5_c_1077_p N_noxref_8_c_1759_n ) capacitor c=0.0153476f \
 //x=1.785 //y=1.22 //x2=2.445 //y2=1.59
cc_885 ( N_noxref_5_c_984_n N_noxref_8_c_1759_n ) capacitor c=0.0230663f \
 //x=2.31 //y=1.915 //x2=2.445 //y2=1.59
cc_886 ( N_noxref_5_c_1075_p N_noxref_8_M0_noxref_s ) capacitor c=0.00798959f \
 //x=1.785 //y=0.91 //x2=0.455 //y2=0.375
cc_887 ( N_noxref_5_c_983_n N_noxref_8_M0_noxref_s ) capacitor c=0.00212176f \
 //x=2.31 //y=1.45 //x2=0.455 //y2=0.375
cc_888 ( N_noxref_5_c_984_n N_noxref_8_M0_noxref_s ) capacitor c=0.00298115f \
 //x=2.31 //y=1.915 //x2=0.455 //y2=0.375
cc_889 ( N_noxref_5_c_1109_p N_noxref_9_c_1788_n ) capacitor c=2.14837e-19 \
 //x=2.155 //y=0.755 //x2=3.015 //y2=0.995
cc_890 ( N_noxref_5_c_981_n N_noxref_9_c_1788_n ) capacitor c=0.00123426f \
 //x=2.31 //y=0.91 //x2=3.015 //y2=0.995
cc_891 ( N_noxref_5_c_982_n N_noxref_9_c_1788_n ) capacitor c=0.0129288f \
 //x=2.31 //y=1.22 //x2=3.015 //y2=0.995
cc_892 ( N_noxref_5_c_983_n N_noxref_9_c_1788_n ) capacitor c=0.00142359f \
 //x=2.31 //y=1.45 //x2=3.015 //y2=0.995
cc_893 ( N_noxref_5_c_1075_p N_noxref_9_M1_noxref_d ) capacitor c=0.00223875f \
 //x=1.785 //y=0.91 //x2=1.86 //y2=0.91
cc_894 ( N_noxref_5_c_1077_p N_noxref_9_M1_noxref_d ) capacitor c=0.00262485f \
 //x=1.785 //y=1.22 //x2=1.86 //y2=0.91
cc_895 ( N_noxref_5_c_1109_p N_noxref_9_M1_noxref_d ) capacitor c=0.00220746f \
 //x=2.155 //y=0.755 //x2=1.86 //y2=0.91
cc_896 ( N_noxref_5_c_1116_p N_noxref_9_M1_noxref_d ) capacitor c=0.00194798f \
 //x=2.155 //y=1.375 //x2=1.86 //y2=0.91
cc_897 ( N_noxref_5_c_981_n N_noxref_9_M1_noxref_d ) capacitor c=0.00198465f \
 //x=2.31 //y=0.91 //x2=1.86 //y2=0.91
cc_898 ( N_noxref_5_c_982_n N_noxref_9_M1_noxref_d ) capacitor c=0.00128384f \
 //x=2.31 //y=1.22 //x2=1.86 //y2=0.91
cc_899 ( N_noxref_5_c_981_n N_noxref_9_M2_noxref_s ) capacitor c=7.21316e-19 \
 //x=2.31 //y=0.91 //x2=2.965 //y2=0.375
cc_900 ( N_noxref_5_c_982_n N_noxref_9_M2_noxref_s ) capacitor c=0.00348171f \
 //x=2.31 //y=1.22 //x2=2.965 //y2=0.375
cc_901 ( N_noxref_5_c_932_n N_noxref_10_c_1850_n ) capacitor c=0.0016972f \
 //x=13.205 //y=4.44 //x2=6.66 //y2=4.535
cc_902 ( N_noxref_5_c_932_n N_noxref_10_c_1841_n ) capacitor c=0.0189188f \
 //x=13.205 //y=4.44 //x2=6.66 //y2=2.08
cc_903 ( N_noxref_5_c_932_n N_noxref_10_c_1863_n ) capacitor c=0.00960248f \
 //x=13.205 //y=4.44 //x2=7.065 //y2=4.79
cc_904 ( N_noxref_5_c_932_n N_noxref_10_c_1874_n ) capacitor c=0.00203982f \
 //x=13.205 //y=4.44 //x2=6.69 //y2=4.7
cc_905 ( N_noxref_5_c_1009_n N_noxref_13_c_2026_n ) capacitor c=0.00623646f \
 //x=13.355 //y=1.56 //x2=13.135 //y2=1.495
cc_906 ( N_noxref_5_c_1014_n N_noxref_13_c_2026_n ) capacitor c=0.00176439f \
 //x=13.32 //y=2.08 //x2=13.135 //y2=1.495
cc_907 ( N_noxref_5_c_930_n N_noxref_13_c_2027_n ) capacitor c=0.0016032f \
 //x=13.32 //y=2.08 //x2=14.02 //y2=0.53
cc_908 ( N_noxref_5_c_1004_n N_noxref_13_c_2027_n ) capacitor c=0.0188655f \
 //x=13.355 //y=0.905 //x2=14.02 //y2=0.53
cc_909 ( N_noxref_5_c_1012_n N_noxref_13_c_2027_n ) capacitor c=0.00656458f \
 //x=13.885 //y=0.905 //x2=14.02 //y2=0.53
cc_910 ( N_noxref_5_c_1014_n N_noxref_13_c_2027_n ) capacitor c=2.1838e-19 \
 //x=13.32 //y=2.08 //x2=14.02 //y2=0.53
cc_911 ( N_noxref_5_c_1004_n N_noxref_13_M7_noxref_s ) capacitor c=0.00623646f \
 //x=13.355 //y=0.905 //x2=12.03 //y2=0.365
cc_912 ( N_noxref_5_c_1012_n N_noxref_13_M7_noxref_s ) capacitor c=0.0143002f \
 //x=13.885 //y=0.905 //x2=12.03 //y2=0.365
cc_913 ( N_noxref_5_c_1013_n N_noxref_13_M7_noxref_s ) capacitor c=0.00290153f \
 //x=13.885 //y=1.25 //x2=12.03 //y2=0.365
cc_914 ( N_noxref_6_c_1207_n N_noxref_7_c_1385_n ) capacitor c=0.147021f \
 //x=5.805 //y=3.7 //x2=9.875 //y2=4.07
cc_915 ( N_noxref_6_c_1208_n N_noxref_7_c_1385_n ) capacitor c=0.0294294f \
 //x=4.185 //y=3.7 //x2=9.875 //y2=4.07
cc_916 ( N_noxref_6_c_1134_n N_noxref_7_c_1385_n ) capacitor c=0.338937f \
 //x=15.795 //y=3.7 //x2=9.875 //y2=4.07
cc_917 ( N_noxref_6_c_1215_n N_noxref_7_c_1385_n ) capacitor c=0.0264478f \
 //x=6.035 //y=3.7 //x2=9.875 //y2=4.07
cc_918 ( N_noxref_6_c_1165_n N_noxref_7_c_1385_n ) capacitor c=0.0154449f \
 //x=1.615 //y=5.155 //x2=9.875 //y2=4.07
cc_919 ( N_noxref_6_c_1175_n N_noxref_7_c_1385_n ) capacitor c=0.0200328f \
 //x=4.07 //y=3.7 //x2=9.875 //y2=4.07
cc_920 ( N_noxref_6_c_1137_n N_noxref_7_c_1385_n ) capacitor c=0.0203111f \
 //x=5.92 //y=2.08 //x2=9.875 //y2=4.07
cc_921 ( N_noxref_6_c_1134_n N_noxref_7_c_1416_n ) capacitor c=0.339146f \
 //x=15.795 //y=3.7 //x2=13.945 //y2=4.07
cc_922 ( N_noxref_6_c_1134_n N_noxref_7_c_1486_n ) capacitor c=0.0267832f \
 //x=15.795 //y=3.7 //x2=10.105 //y2=4.07
cc_923 ( N_noxref_6_c_1134_n N_noxref_7_c_1387_n ) capacitor c=0.176049f \
 //x=15.795 //y=3.7 //x2=19.865 //y2=4.07
cc_924 ( N_noxref_6_c_1138_n N_noxref_7_c_1387_n ) capacitor c=0.0242341f \
 //x=15.91 //y=2.08 //x2=19.865 //y2=4.07
cc_925 ( N_noxref_6_c_1191_n N_noxref_7_c_1387_n ) capacitor c=0.00703556f \
 //x=15.91 //y=4.7 //x2=19.865 //y2=4.07
cc_926 ( N_noxref_6_c_1134_n N_noxref_7_c_1430_n ) capacitor c=0.0266833f \
 //x=15.795 //y=3.7 //x2=14.175 //y2=4.07
cc_927 ( N_noxref_6_c_1138_n N_noxref_7_c_1430_n ) capacitor c=3.50683e-19 \
 //x=15.91 //y=2.08 //x2=14.175 //y2=4.07
cc_928 ( N_noxref_6_c_1134_n N_noxref_7_c_1390_n ) capacitor c=0.0243898f \
 //x=15.795 //y=3.7 //x2=9.99 //y2=2.08
cc_929 ( N_noxref_6_c_1134_n N_noxref_7_c_1626_n ) capacitor c=0.00433945f \
 //x=15.795 //y=3.7 //x2=13.705 //y2=1.655
cc_930 ( N_noxref_6_c_1134_n N_noxref_7_c_1393_n ) capacitor c=0.0269561f \
 //x=15.795 //y=3.7 //x2=14.06 //y2=4.07
cc_931 ( N_noxref_6_c_1138_n N_noxref_7_c_1393_n ) capacitor c=0.0145678f \
 //x=15.91 //y=2.08 //x2=14.06 //y2=4.07
cc_932 ( N_noxref_6_c_1165_n N_noxref_7_M13_noxref_g ) capacitor c=0.0213876f \
 //x=1.615 //y=5.155 //x2=1.31 //y2=6.02
cc_933 ( N_noxref_6_c_1161_n N_noxref_7_M14_noxref_g ) capacitor c=0.0178794f \
 //x=2.325 //y=5.155 //x2=1.75 //y2=6.02
cc_934 ( N_noxref_6_M13_noxref_d N_noxref_7_M14_noxref_g ) capacitor \
 c=0.0180032f //x=1.385 //y=5.02 //x2=1.75 //y2=6.02
cc_935 ( N_noxref_6_c_1165_n N_noxref_7_c_1595_n ) capacitor c=0.00429591f \
 //x=1.615 //y=5.155 //x2=1.675 //y2=4.79
cc_936 ( N_noxref_6_M2_noxref_d N_noxref_8_M0_noxref_s ) capacitor \
 c=0.00309936f //x=3.395 //y=0.915 //x2=0.455 //y2=0.375
cc_937 ( N_noxref_6_c_1136_n N_noxref_9_c_1793_n ) capacitor c=0.00466084f \
 //x=3.985 //y=1.665 //x2=3.985 //y2=0.54
cc_938 ( N_noxref_6_M2_noxref_d N_noxref_9_c_1793_n ) capacitor c=0.0117786f \
 //x=3.395 //y=0.915 //x2=3.985 //y2=0.54
cc_939 ( N_noxref_6_c_1221_n N_noxref_9_c_1807_n ) capacitor c=0.020048f \
 //x=3.67 //y=1.665 //x2=3.1 //y2=0.995
cc_940 ( N_noxref_6_M2_noxref_d N_noxref_9_M1_noxref_d ) capacitor \
 c=5.27807e-19 //x=3.395 //y=0.915 //x2=1.86 //y2=0.91
cc_941 ( N_noxref_6_c_1136_n N_noxref_9_M2_noxref_s ) capacitor c=0.0207678f \
 //x=3.985 //y=1.665 //x2=2.965 //y2=0.375
cc_942 ( N_noxref_6_M2_noxref_d N_noxref_9_M2_noxref_s ) capacitor \
 c=0.0426444f //x=3.395 //y=0.915 //x2=2.965 //y2=0.375
cc_943 ( N_noxref_6_c_1137_n N_noxref_10_c_1850_n ) capacitor c=0.00400249f \
 //x=5.92 //y=2.08 //x2=6.66 //y2=4.535
cc_944 ( N_noxref_6_c_1190_n N_noxref_10_c_1850_n ) capacitor c=0.00417994f \
 //x=5.92 //y=4.7 //x2=6.66 //y2=4.535
cc_945 ( N_noxref_6_c_1134_n N_noxref_10_c_1841_n ) capacitor c=0.0169594f \
 //x=15.795 //y=3.7 //x2=6.66 //y2=2.08
cc_946 ( N_noxref_6_c_1215_n N_noxref_10_c_1841_n ) capacitor c=0.00131333f \
 //x=6.035 //y=3.7 //x2=6.66 //y2=2.08
cc_947 ( N_noxref_6_c_1175_n N_noxref_10_c_1841_n ) capacitor c=8.12815e-19 \
 //x=4.07 //y=3.7 //x2=6.66 //y2=2.08
cc_948 ( N_noxref_6_c_1137_n N_noxref_10_c_1841_n ) capacitor c=0.0781945f \
 //x=5.92 //y=2.08 //x2=6.66 //y2=2.08
cc_949 ( N_noxref_6_c_1143_n N_noxref_10_c_1841_n ) capacitor c=0.00308814f \
 //x=5.725 //y=1.915 //x2=6.66 //y2=2.08
cc_950 ( N_noxref_6_M19_noxref_g N_noxref_10_M21_noxref_g ) capacitor \
 c=0.0104611f //x=5.82 //y=6.02 //x2=6.7 //y2=6.02
cc_951 ( N_noxref_6_M20_noxref_g N_noxref_10_M21_noxref_g ) capacitor \
 c=0.106811f //x=6.26 //y=6.02 //x2=6.7 //y2=6.02
cc_952 ( N_noxref_6_M20_noxref_g N_noxref_10_M22_noxref_g ) capacitor \
 c=0.0100341f //x=6.26 //y=6.02 //x2=7.14 //y2=6.02
cc_953 ( N_noxref_6_c_1139_n N_noxref_10_c_1860_n ) capacitor c=4.86506e-19 \
 //x=5.725 //y=0.865 //x2=6.695 //y2=0.905
cc_954 ( N_noxref_6_c_1141_n N_noxref_10_c_1860_n ) capacitor c=0.00152104f \
 //x=5.725 //y=1.21 //x2=6.695 //y2=0.905
cc_955 ( N_noxref_6_c_1146_n N_noxref_10_c_1860_n ) capacitor c=0.0151475f \
 //x=6.255 //y=0.865 //x2=6.695 //y2=0.905
cc_956 ( N_noxref_6_c_1142_n N_noxref_10_c_1861_n ) capacitor c=0.00109982f \
 //x=5.725 //y=1.52 //x2=6.695 //y2=1.25
cc_957 ( N_noxref_6_c_1148_n N_noxref_10_c_1861_n ) capacitor c=0.0111064f \
 //x=6.255 //y=1.21 //x2=6.695 //y2=1.25
cc_958 ( N_noxref_6_c_1142_n N_noxref_10_c_1862_n ) capacitor c=9.57794e-19 \
 //x=5.725 //y=1.52 //x2=6.695 //y2=1.56
cc_959 ( N_noxref_6_c_1143_n N_noxref_10_c_1862_n ) capacitor c=0.00662747f \
 //x=5.725 //y=1.915 //x2=6.695 //y2=1.56
cc_960 ( N_noxref_6_c_1148_n N_noxref_10_c_1862_n ) capacitor c=0.00862358f \
 //x=6.255 //y=1.21 //x2=6.695 //y2=1.56
cc_961 ( N_noxref_6_c_1146_n N_noxref_10_c_1868_n ) capacitor c=0.00124821f \
 //x=6.255 //y=0.865 //x2=7.225 //y2=0.905
cc_962 ( N_noxref_6_c_1148_n N_noxref_10_c_1869_n ) capacitor c=0.00200715f \
 //x=6.255 //y=1.21 //x2=7.225 //y2=1.25
cc_963 ( N_noxref_6_c_1137_n N_noxref_10_c_1871_n ) capacitor c=0.00307062f \
 //x=5.92 //y=2.08 //x2=6.66 //y2=2.08
cc_964 ( N_noxref_6_c_1143_n N_noxref_10_c_1871_n ) capacitor c=0.0179092f \
 //x=5.725 //y=1.915 //x2=6.66 //y2=2.08
cc_965 ( N_noxref_6_c_1137_n N_noxref_10_c_1874_n ) capacitor c=0.00344981f \
 //x=5.92 //y=2.08 //x2=6.69 //y2=4.7
cc_966 ( N_noxref_6_c_1190_n N_noxref_10_c_1874_n ) capacitor c=0.0293367f \
 //x=5.92 //y=4.7 //x2=6.69 //y2=4.7
cc_967 ( N_noxref_6_c_1136_n N_noxref_11_c_1933_n ) capacitor c=3.04182e-19 \
 //x=3.985 //y=1.665 //x2=5.505 //y2=1.495
cc_968 ( N_noxref_6_c_1143_n N_noxref_11_c_1933_n ) capacitor c=0.0034165f \
 //x=5.725 //y=1.915 //x2=5.505 //y2=1.495
cc_969 ( N_noxref_6_c_1137_n N_noxref_11_c_1914_n ) capacitor c=0.0116993f \
 //x=5.92 //y=2.08 //x2=6.39 //y2=1.58
cc_970 ( N_noxref_6_c_1142_n N_noxref_11_c_1914_n ) capacitor c=0.00703567f \
 //x=5.725 //y=1.52 //x2=6.39 //y2=1.58
cc_971 ( N_noxref_6_c_1143_n N_noxref_11_c_1914_n ) capacitor c=0.0203514f \
 //x=5.725 //y=1.915 //x2=6.39 //y2=1.58
cc_972 ( N_noxref_6_c_1145_n N_noxref_11_c_1914_n ) capacitor c=0.00780629f \
 //x=6.1 //y=1.365 //x2=6.39 //y2=1.58
cc_973 ( N_noxref_6_c_1148_n N_noxref_11_c_1914_n ) capacitor c=0.00339872f \
 //x=6.255 //y=1.21 //x2=6.39 //y2=1.58
cc_974 ( N_noxref_6_c_1143_n N_noxref_11_c_1921_n ) capacitor c=6.71402e-19 \
 //x=5.725 //y=1.915 //x2=6.475 //y2=1.495
cc_975 ( N_noxref_6_c_1139_n N_noxref_11_M3_noxref_s ) capacitor c=0.0327502f \
 //x=5.725 //y=0.865 //x2=5.37 //y2=0.365
cc_976 ( N_noxref_6_c_1142_n N_noxref_11_M3_noxref_s ) capacitor c=3.48408e-19 \
 //x=5.725 //y=1.52 //x2=5.37 //y2=0.365
cc_977 ( N_noxref_6_c_1146_n N_noxref_11_M3_noxref_s ) capacitor c=0.0120759f \
 //x=6.255 //y=0.865 //x2=5.37 //y2=0.365
cc_978 ( N_noxref_6_c_1134_n N_noxref_12_c_1966_n ) capacitor c=0.00299723f \
 //x=15.795 //y=3.7 //x2=9.72 //y2=1.58
cc_979 ( N_noxref_6_c_1134_n N_noxref_12_c_1973_n ) capacitor c=0.00187232f \
 //x=15.795 //y=3.7 //x2=9.805 //y2=1.495
cc_980 ( N_noxref_6_c_1134_n N_noxref_12_c_1974_n ) capacitor c=4.7198e-19 \
 //x=15.795 //y=3.7 //x2=10.69 //y2=0.53
cc_981 ( N_noxref_6_c_1134_n N_noxref_13_c_2019_n ) capacitor c=0.00299723f \
 //x=15.795 //y=3.7 //x2=13.05 //y2=1.58
cc_982 ( N_noxref_6_c_1134_n N_noxref_13_c_2026_n ) capacitor c=0.00187232f \
 //x=15.795 //y=3.7 //x2=13.135 //y2=1.495
cc_983 ( N_noxref_6_c_1134_n N_noxref_13_c_2027_n ) capacitor c=4.7198e-19 \
 //x=15.795 //y=3.7 //x2=14.02 //y2=0.53
cc_984 ( N_noxref_6_c_1134_n N_noxref_13_M7_noxref_s ) capacitor c=3.97107e-19 \
 //x=15.795 //y=3.7 //x2=12.03 //y2=0.365
cc_985 ( N_noxref_6_c_1138_n N_noxref_14_c_2081_n ) capacitor c=0.00400249f \
 //x=15.91 //y=2.08 //x2=16.65 //y2=4.535
cc_986 ( N_noxref_6_c_1191_n N_noxref_14_c_2081_n ) capacitor c=0.00417994f \
 //x=15.91 //y=4.7 //x2=16.65 //y2=4.535
cc_987 ( N_noxref_6_c_1134_n N_noxref_14_c_2072_n ) capacitor c=0.00735597f \
 //x=15.795 //y=3.7 //x2=16.65 //y2=2.08
cc_988 ( N_noxref_6_c_1138_n N_noxref_14_c_2072_n ) capacitor c=0.0836795f \
 //x=15.91 //y=2.08 //x2=16.65 //y2=2.08
cc_989 ( N_noxref_6_c_1153_n N_noxref_14_c_2072_n ) capacitor c=0.00308814f \
 //x=15.715 //y=1.915 //x2=16.65 //y2=2.08
cc_990 ( N_noxref_6_M31_noxref_g N_noxref_14_M33_noxref_g ) capacitor \
 c=0.0104611f //x=15.81 //y=6.02 //x2=16.69 //y2=6.02
cc_991 ( N_noxref_6_M32_noxref_g N_noxref_14_M33_noxref_g ) capacitor \
 c=0.106811f //x=16.25 //y=6.02 //x2=16.69 //y2=6.02
cc_992 ( N_noxref_6_M32_noxref_g N_noxref_14_M34_noxref_g ) capacitor \
 c=0.0100341f //x=16.25 //y=6.02 //x2=17.13 //y2=6.02
cc_993 ( N_noxref_6_c_1149_n N_noxref_14_c_2089_n ) capacitor c=4.86506e-19 \
 //x=15.715 //y=0.865 //x2=16.685 //y2=0.905
cc_994 ( N_noxref_6_c_1151_n N_noxref_14_c_2089_n ) capacitor c=0.00152104f \
 //x=15.715 //y=1.21 //x2=16.685 //y2=0.905
cc_995 ( N_noxref_6_c_1156_n N_noxref_14_c_2089_n ) capacitor c=0.0151475f \
 //x=16.245 //y=0.865 //x2=16.685 //y2=0.905
cc_996 ( N_noxref_6_c_1152_n N_noxref_14_c_2092_n ) capacitor c=0.00109982f \
 //x=15.715 //y=1.52 //x2=16.685 //y2=1.25
cc_997 ( N_noxref_6_c_1158_n N_noxref_14_c_2092_n ) capacitor c=0.0111064f \
 //x=16.245 //y=1.21 //x2=16.685 //y2=1.25
cc_998 ( N_noxref_6_c_1152_n N_noxref_14_c_2094_n ) capacitor c=9.57794e-19 \
 //x=15.715 //y=1.52 //x2=16.685 //y2=1.56
cc_999 ( N_noxref_6_c_1153_n N_noxref_14_c_2094_n ) capacitor c=0.00662747f \
 //x=15.715 //y=1.915 //x2=16.685 //y2=1.56
cc_1000 ( N_noxref_6_c_1158_n N_noxref_14_c_2094_n ) capacitor c=0.00862358f \
 //x=16.245 //y=1.21 //x2=16.685 //y2=1.56
cc_1001 ( N_noxref_6_c_1156_n N_noxref_14_c_2097_n ) capacitor c=0.00124821f \
 //x=16.245 //y=0.865 //x2=17.215 //y2=0.905
cc_1002 ( N_noxref_6_c_1158_n N_noxref_14_c_2098_n ) capacitor c=0.00200715f \
 //x=16.245 //y=1.21 //x2=17.215 //y2=1.25
cc_1003 ( N_noxref_6_c_1138_n N_noxref_14_c_2099_n ) capacitor c=0.00307062f \
 //x=15.91 //y=2.08 //x2=16.65 //y2=2.08
cc_1004 ( N_noxref_6_c_1153_n N_noxref_14_c_2099_n ) capacitor c=0.0179092f \
 //x=15.715 //y=1.915 //x2=16.65 //y2=2.08
cc_1005 ( N_noxref_6_c_1138_n N_noxref_14_c_2101_n ) capacitor c=0.00344981f \
 //x=15.91 //y=2.08 //x2=16.68 //y2=4.7
cc_1006 ( N_noxref_6_c_1191_n N_noxref_14_c_2101_n ) capacitor c=0.0293367f \
 //x=15.91 //y=4.7 //x2=16.68 //y2=4.7
cc_1007 ( N_noxref_6_M32_noxref_g N_noxref_15_c_2146_n ) capacitor c=0.017965f \
 //x=16.25 //y=6.02 //x2=16.825 //y2=5.2
cc_1008 ( N_noxref_6_c_1138_n N_noxref_15_c_2150_n ) capacitor c=0.00530485f \
 //x=15.91 //y=2.08 //x2=16.115 //y2=5.2
cc_1009 ( N_noxref_6_M31_noxref_g N_noxref_15_c_2150_n ) capacitor \
 c=0.0177326f //x=15.81 //y=6.02 //x2=16.115 //y2=5.2
cc_1010 ( N_noxref_6_c_1191_n N_noxref_15_c_2150_n ) capacitor c=0.00582246f \
 //x=15.91 //y=4.7 //x2=16.115 //y2=5.2
cc_1011 ( N_noxref_6_c_1138_n N_noxref_15_c_2142_n ) capacitor c=0.00394392f \
 //x=15.91 //y=2.08 //x2=17.39 //y2=5.115
cc_1012 ( N_noxref_6_M32_noxref_g N_noxref_15_M31_noxref_d ) capacitor \
 c=0.0173476f //x=16.25 //y=6.02 //x2=15.885 //y2=5.02
cc_1013 ( N_noxref_6_c_1134_n N_noxref_16_c_2232_n ) capacitor c=0.00188872f \
 //x=15.795 //y=3.7 //x2=15.495 //y2=1.495
cc_1014 ( N_noxref_6_c_1153_n N_noxref_16_c_2232_n ) capacitor c=0.0034165f \
 //x=15.715 //y=1.915 //x2=15.495 //y2=1.495
cc_1015 ( N_noxref_6_c_1134_n N_noxref_16_c_2213_n ) capacitor c=0.0056636f \
 //x=15.795 //y=3.7 //x2=16.38 //y2=1.58
cc_1016 ( N_noxref_6_c_1138_n N_noxref_16_c_2213_n ) capacitor c=0.011766f \
 //x=15.91 //y=2.08 //x2=16.38 //y2=1.58
cc_1017 ( N_noxref_6_c_1152_n N_noxref_16_c_2213_n ) capacitor c=0.00703567f \
 //x=15.715 //y=1.52 //x2=16.38 //y2=1.58
cc_1018 ( N_noxref_6_c_1153_n N_noxref_16_c_2213_n ) capacitor c=0.0207598f \
 //x=15.715 //y=1.915 //x2=16.38 //y2=1.58
cc_1019 ( N_noxref_6_c_1155_n N_noxref_16_c_2213_n ) capacitor c=0.00780629f \
 //x=16.09 //y=1.365 //x2=16.38 //y2=1.58
cc_1020 ( N_noxref_6_c_1158_n N_noxref_16_c_2213_n ) capacitor c=0.00339872f \
 //x=16.245 //y=1.21 //x2=16.38 //y2=1.58
cc_1021 ( N_noxref_6_c_1153_n N_noxref_16_c_2220_n ) capacitor c=6.71402e-19 \
 //x=15.715 //y=1.915 //x2=16.465 //y2=1.495
cc_1022 ( N_noxref_6_c_1149_n N_noxref_16_M9_noxref_s ) capacitor c=0.0326577f \
 //x=15.715 //y=0.865 //x2=15.36 //y2=0.365
cc_1023 ( N_noxref_6_c_1152_n N_noxref_16_M9_noxref_s ) capacitor \
 c=3.48408e-19 //x=15.715 //y=1.52 //x2=15.36 //y2=0.365
cc_1024 ( N_noxref_6_c_1156_n N_noxref_16_M9_noxref_s ) capacitor c=0.0120759f \
 //x=16.245 //y=0.865 //x2=15.36 //y2=0.365
cc_1025 ( N_noxref_7_c_1400_n N_noxref_8_c_1766_n ) capacitor c=0.0034165f \
 //x=0.81 //y=1.915 //x2=0.59 //y2=1.505
cc_1026 ( N_noxref_7_c_1385_n N_noxref_8_c_1741_n ) capacitor c=0.00179505f \
 //x=9.875 //y=4.07 //x2=1.475 //y2=1.59
cc_1027 ( N_noxref_7_c_1386_n N_noxref_8_c_1741_n ) capacitor c=0.00102628f \
 //x=1.225 //y=4.07 //x2=1.475 //y2=1.59
cc_1028 ( N_noxref_7_c_1389_n N_noxref_8_c_1741_n ) capacitor c=0.0122033f \
 //x=1.11 //y=2.08 //x2=1.475 //y2=1.59
cc_1029 ( N_noxref_7_c_1399_n N_noxref_8_c_1741_n ) capacitor c=0.00703864f \
 //x=0.81 //y=1.53 //x2=1.475 //y2=1.59
cc_1030 ( N_noxref_7_c_1400_n N_noxref_8_c_1741_n ) capacitor c=0.0259045f \
 //x=0.81 //y=1.915 //x2=1.475 //y2=1.59
cc_1031 ( N_noxref_7_c_1402_n N_noxref_8_c_1741_n ) capacitor c=0.00708583f \
 //x=1.185 //y=1.375 //x2=1.475 //y2=1.59
cc_1032 ( N_noxref_7_c_1405_n N_noxref_8_c_1741_n ) capacitor c=0.00698822f \
 //x=1.34 //y=1.22 //x2=1.475 //y2=1.59
cc_1033 ( N_noxref_7_c_1385_n N_noxref_8_c_1759_n ) capacitor c=0.0058169f \
 //x=9.875 //y=4.07 //x2=2.445 //y2=1.59
cc_1034 ( N_noxref_7_c_1385_n N_noxref_8_M0_noxref_s ) capacitor c=0.00262629f \
 //x=9.875 //y=4.07 //x2=0.455 //y2=0.375
cc_1035 ( N_noxref_7_c_1396_n N_noxref_8_M0_noxref_s ) capacitor c=0.0327271f \
 //x=0.81 //y=0.875 //x2=0.455 //y2=0.375
cc_1036 ( N_noxref_7_c_1399_n N_noxref_8_M0_noxref_s ) capacitor c=7.99997e-19 \
 //x=0.81 //y=1.53 //x2=0.455 //y2=0.375
cc_1037 ( N_noxref_7_c_1400_n N_noxref_8_M0_noxref_s ) capacitor c=0.00122123f \
 //x=0.81 //y=1.915 //x2=0.455 //y2=0.375
cc_1038 ( N_noxref_7_c_1403_n N_noxref_8_M0_noxref_s ) capacitor c=0.0121427f \
 //x=1.34 //y=0.875 //x2=0.455 //y2=0.375
cc_1039 ( N_noxref_7_c_1385_n N_noxref_9_c_1788_n ) capacitor c=0.0020922f \
 //x=9.875 //y=4.07 //x2=3.015 //y2=0.995
cc_1040 ( N_noxref_7_c_1385_n N_noxref_9_M2_noxref_s ) capacitor c=0.00143334f \
 //x=9.875 //y=4.07 //x2=2.965 //y2=0.375
cc_1041 ( N_noxref_7_c_1385_n N_noxref_10_c_1841_n ) capacitor c=0.0169317f \
 //x=9.875 //y=4.07 //x2=6.66 //y2=2.08
cc_1042 ( N_noxref_7_c_1502_n N_noxref_12_c_1973_n ) capacitor c=0.00623646f \
 //x=10.025 //y=1.56 //x2=9.805 //y2=1.495
cc_1043 ( N_noxref_7_c_1507_n N_noxref_12_c_1973_n ) capacitor c=0.00176439f \
 //x=9.99 //y=2.08 //x2=9.805 //y2=1.495
cc_1044 ( N_noxref_7_c_1390_n N_noxref_12_c_1974_n ) capacitor c=0.0016032f \
 //x=9.99 //y=2.08 //x2=10.69 //y2=0.53
cc_1045 ( N_noxref_7_c_1497_n N_noxref_12_c_1974_n ) capacitor c=0.0188655f \
 //x=10.025 //y=0.905 //x2=10.69 //y2=0.53
cc_1046 ( N_noxref_7_c_1505_n N_noxref_12_c_1974_n ) capacitor c=0.00656458f \
 //x=10.555 //y=0.905 //x2=10.69 //y2=0.53
cc_1047 ( N_noxref_7_c_1507_n N_noxref_12_c_1974_n ) capacitor c=2.1838e-19 \
 //x=9.99 //y=2.08 //x2=10.69 //y2=0.53
cc_1048 ( N_noxref_7_c_1497_n N_noxref_12_M5_noxref_s ) capacitor \
 c=0.00623646f //x=10.025 //y=0.905 //x2=8.7 //y2=0.365
cc_1049 ( N_noxref_7_c_1505_n N_noxref_12_M5_noxref_s ) capacitor c=0.0143002f \
 //x=10.555 //y=0.905 //x2=8.7 //y2=0.365
cc_1050 ( N_noxref_7_c_1506_n N_noxref_12_M5_noxref_s ) capacitor \
 c=0.00290153f //x=10.555 //y=1.25 //x2=8.7 //y2=0.365
cc_1051 ( N_noxref_7_c_1626_n N_noxref_13_c_2038_n ) capacitor c=3.15806e-19 \
 //x=13.705 //y=1.655 //x2=12.165 //y2=1.495
cc_1052 ( N_noxref_7_c_1626_n N_noxref_13_c_2026_n ) capacitor c=0.0203424f \
 //x=13.705 //y=1.655 //x2=13.135 //y2=1.495
cc_1053 ( N_noxref_7_c_1392_n N_noxref_13_c_2027_n ) capacitor c=0.00467111f \
 //x=13.975 //y=1.655 //x2=14.02 //y2=0.53
cc_1054 ( N_noxref_7_M8_noxref_d N_noxref_13_c_2027_n ) capacitor c=0.0117932f \
 //x=13.43 //y=0.905 //x2=14.02 //y2=0.53
cc_1055 ( N_noxref_7_c_1392_n N_noxref_13_M7_noxref_s ) capacitor c=0.014284f \
 //x=13.975 //y=1.655 //x2=12.03 //y2=0.365
cc_1056 ( N_noxref_7_M8_noxref_d N_noxref_13_M7_noxref_s ) capacitor \
 c=0.043966f //x=13.43 //y=0.905 //x2=12.03 //y2=0.365
cc_1057 ( N_noxref_7_c_1387_n N_noxref_14_c_2081_n ) capacitor c=0.00135863f \
 //x=19.865 //y=4.07 //x2=16.65 //y2=4.535
cc_1058 ( N_noxref_7_c_1387_n N_noxref_14_c_2072_n ) capacitor c=0.0265817f \
 //x=19.865 //y=4.07 //x2=16.65 //y2=2.08
cc_1059 ( N_noxref_7_c_1393_n N_noxref_14_c_2072_n ) capacitor c=0.00116185f \
 //x=14.06 //y=4.07 //x2=16.65 //y2=2.08
cc_1060 ( N_noxref_7_c_1387_n N_noxref_14_c_2106_n ) capacitor c=0.00561113f \
 //x=19.865 //y=4.07 //x2=17.055 //y2=4.79
cc_1061 ( N_noxref_7_c_1387_n N_noxref_14_c_2101_n ) capacitor c=0.00127126f \
 //x=19.865 //y=4.07 //x2=16.68 //y2=4.7
cc_1062 ( N_noxref_7_c_1387_n N_noxref_15_c_2146_n ) capacitor c=0.0137325f \
 //x=19.865 //y=4.07 //x2=16.825 //y2=5.2
cc_1063 ( N_noxref_7_c_1387_n N_noxref_15_c_2150_n ) capacitor c=0.013479f \
 //x=19.865 //y=4.07 //x2=16.115 //y2=5.2
cc_1064 ( N_noxref_7_c_1387_n N_noxref_15_c_2177_n ) capacitor c=0.0034482f \
 //x=19.865 //y=4.07 //x2=17.035 //y2=1.655
cc_1065 ( N_noxref_7_c_1387_n N_noxref_15_c_2142_n ) capacitor c=0.0289918f \
 //x=19.865 //y=4.07 //x2=17.39 //y2=5.115
cc_1066 ( N_noxref_7_c_1393_n N_noxref_15_c_2142_n ) capacitor c=3.49822e-19 \
 //x=14.06 //y=4.07 //x2=17.39 //y2=5.115
cc_1067 ( N_noxref_7_c_1394_n N_noxref_15_c_2142_n ) capacitor c=8.97258e-19 \
 //x=19.98 //y=2.08 //x2=17.39 //y2=5.115
cc_1068 ( N_noxref_7_c_1392_n N_noxref_16_c_2232_n ) capacitor c=3.22188e-19 \
 //x=13.975 //y=1.655 //x2=15.495 //y2=1.495
cc_1069 ( N_noxref_7_c_1387_n N_noxref_16_c_2213_n ) capacitor c=0.00234538f \
 //x=19.865 //y=4.07 //x2=16.38 //y2=1.58
cc_1070 ( N_noxref_7_c_1387_n N_noxref_16_c_2220_n ) capacitor c=0.00121496f \
 //x=19.865 //y=4.07 //x2=16.465 //y2=1.495
cc_1071 ( N_noxref_7_c_1387_n N_noxref_16_M9_noxref_s ) capacitor \
 c=2.47199e-19 //x=19.865 //y=4.07 //x2=15.36 //y2=0.365
cc_1072 ( N_noxref_7_c_1387_n N_noxref_17_c_2265_n ) capacitor c=0.0299282f \
 //x=19.865 //y=4.07 //x2=19.24 //y2=2.08
cc_1073 ( N_noxref_7_c_1681_p N_noxref_17_c_2265_n ) capacitor c=0.00400249f \
 //x=19.98 //y=4.535 //x2=19.24 //y2=2.08
cc_1074 ( N_noxref_7_c_1394_n N_noxref_17_c_2265_n ) capacitor c=0.0858984f \
 //x=19.98 //y=2.08 //x2=19.24 //y2=2.08
cc_1075 ( N_noxref_7_c_1683_p N_noxref_17_c_2265_n ) capacitor c=0.00307062f \
 //x=19.98 //y=2.08 //x2=19.24 //y2=2.08
cc_1076 ( N_noxref_7_c_1684_p N_noxref_17_c_2265_n ) capacitor c=0.00344981f \
 //x=20.01 //y=4.7 //x2=19.24 //y2=2.08
cc_1077 ( N_noxref_7_M37_noxref_g N_noxref_17_M35_noxref_g ) capacitor \
 c=0.0104611f //x=20.02 //y=6.02 //x2=19.14 //y2=6.02
cc_1078 ( N_noxref_7_M37_noxref_g N_noxref_17_M36_noxref_g ) capacitor \
 c=0.106811f //x=20.02 //y=6.02 //x2=19.58 //y2=6.02
cc_1079 ( N_noxref_7_M38_noxref_g N_noxref_17_M36_noxref_g ) capacitor \
 c=0.0100341f //x=20.46 //y=6.02 //x2=19.58 //y2=6.02
cc_1080 ( N_noxref_7_c_1688_p N_noxref_17_c_2266_n ) capacitor c=4.86506e-19 \
 //x=20.015 //y=0.905 //x2=19.045 //y2=0.865
cc_1081 ( N_noxref_7_c_1688_p N_noxref_17_c_2268_n ) capacitor c=0.00152104f \
 //x=20.015 //y=0.905 //x2=19.045 //y2=1.21
cc_1082 ( N_noxref_7_c_1690_p N_noxref_17_c_2269_n ) capacitor c=0.00109982f \
 //x=20.015 //y=1.25 //x2=19.045 //y2=1.52
cc_1083 ( N_noxref_7_c_1691_p N_noxref_17_c_2269_n ) capacitor c=9.57794e-19 \
 //x=20.015 //y=1.56 //x2=19.045 //y2=1.52
cc_1084 ( N_noxref_7_c_1394_n N_noxref_17_c_2270_n ) capacitor c=0.00308814f \
 //x=19.98 //y=2.08 //x2=19.045 //y2=1.915
cc_1085 ( N_noxref_7_c_1691_p N_noxref_17_c_2270_n ) capacitor c=0.00662747f \
 //x=20.015 //y=1.56 //x2=19.045 //y2=1.915
cc_1086 ( N_noxref_7_c_1683_p N_noxref_17_c_2270_n ) capacitor c=0.0179092f \
 //x=19.98 //y=2.08 //x2=19.045 //y2=1.915
cc_1087 ( N_noxref_7_c_1688_p N_noxref_17_c_2273_n ) capacitor c=0.0151475f \
 //x=20.015 //y=0.905 //x2=19.575 //y2=0.865
cc_1088 ( N_noxref_7_c_1696_p N_noxref_17_c_2273_n ) capacitor c=0.00124821f \
 //x=20.545 //y=0.905 //x2=19.575 //y2=0.865
cc_1089 ( N_noxref_7_c_1690_p N_noxref_17_c_2275_n ) capacitor c=0.0111064f \
 //x=20.015 //y=1.25 //x2=19.575 //y2=1.21
cc_1090 ( N_noxref_7_c_1691_p N_noxref_17_c_2275_n ) capacitor c=0.00862358f \
 //x=20.015 //y=1.56 //x2=19.575 //y2=1.21
cc_1091 ( N_noxref_7_c_1699_p N_noxref_17_c_2275_n ) capacitor c=0.00200715f \
 //x=20.545 //y=1.25 //x2=19.575 //y2=1.21
cc_1092 ( N_noxref_7_c_1387_n N_noxref_17_c_2283_n ) capacitor c=0.00695432f \
 //x=19.865 //y=4.07 //x2=19.24 //y2=4.7
cc_1093 ( N_noxref_7_c_1681_p N_noxref_17_c_2283_n ) capacitor c=0.00417994f \
 //x=19.98 //y=4.535 //x2=19.24 //y2=4.7
cc_1094 ( N_noxref_7_c_1684_p N_noxref_17_c_2283_n ) capacitor c=0.0293367f \
 //x=20.01 //y=4.7 //x2=19.24 //y2=4.7
cc_1095 ( N_noxref_7_c_1387_n N_noxref_18_c_2330_n ) capacitor c=0.0020315f \
 //x=19.865 //y=4.07 //x2=20.155 //y2=5.2
cc_1096 ( N_noxref_7_c_1681_p N_noxref_18_c_2330_n ) capacitor c=0.0129794f \
 //x=19.98 //y=4.535 //x2=20.155 //y2=5.2
cc_1097 ( N_noxref_7_M37_noxref_g N_noxref_18_c_2330_n ) capacitor \
 c=0.0166421f //x=20.02 //y=6.02 //x2=20.155 //y2=5.2
cc_1098 ( N_noxref_7_c_1684_p N_noxref_18_c_2330_n ) capacitor c=0.00346627f \
 //x=20.01 //y=4.7 //x2=20.155 //y2=5.2
cc_1099 ( N_noxref_7_c_1387_n N_noxref_18_c_2334_n ) capacitor c=0.0128624f \
 //x=19.865 //y=4.07 //x2=19.445 //y2=5.2
cc_1100 ( N_noxref_7_M38_noxref_g N_noxref_18_c_2336_n ) capacitor \
 c=0.0223536f //x=20.46 //y=6.02 //x2=20.635 //y2=5.2
cc_1101 ( N_noxref_7_c_1709_p N_noxref_18_c_2325_n ) capacitor c=0.00359704f \
 //x=20.39 //y=1.405 //x2=20.635 //y2=1.655
cc_1102 ( N_noxref_7_c_1699_p N_noxref_18_c_2325_n ) capacitor c=0.00457401f \
 //x=20.545 //y=1.25 //x2=20.635 //y2=1.655
cc_1103 ( N_noxref_7_c_1387_n N_noxref_18_c_2326_n ) capacitor c=0.00642908f \
 //x=19.865 //y=4.07 //x2=20.72 //y2=5.115
cc_1104 ( N_noxref_7_c_1681_p N_noxref_18_c_2326_n ) capacitor c=0.0101115f \
 //x=19.98 //y=4.535 //x2=20.72 //y2=5.115
cc_1105 ( N_noxref_7_c_1394_n N_noxref_18_c_2326_n ) capacitor c=0.0819328f \
 //x=19.98 //y=2.08 //x2=20.72 //y2=5.115
cc_1106 ( N_noxref_7_c_1714_p N_noxref_18_c_2326_n ) capacitor c=0.0142673f \
 //x=20.385 //y=4.79 //x2=20.72 //y2=5.115
cc_1107 ( N_noxref_7_c_1683_p N_noxref_18_c_2326_n ) capacitor c=0.00877984f \
 //x=19.98 //y=2.08 //x2=20.72 //y2=5.115
cc_1108 ( N_noxref_7_c_1716_p N_noxref_18_c_2326_n ) capacitor c=0.00306024f \
 //x=19.98 //y=1.915 //x2=20.72 //y2=5.115
cc_1109 ( N_noxref_7_c_1684_p N_noxref_18_c_2326_n ) capacitor c=0.00533692f \
 //x=20.01 //y=4.7 //x2=20.72 //y2=5.115
cc_1110 ( N_noxref_7_c_1714_p N_noxref_18_c_2366_n ) capacitor c=0.00414324f \
 //x=20.385 //y=4.79 //x2=20.24 //y2=5.2
cc_1111 ( N_noxref_7_c_1688_p N_noxref_18_M12_noxref_d ) capacitor \
 c=0.00217566f //x=20.015 //y=0.905 //x2=20.09 //y2=0.905
cc_1112 ( N_noxref_7_c_1690_p N_noxref_18_M12_noxref_d ) capacitor \
 c=0.0034598f //x=20.015 //y=1.25 //x2=20.09 //y2=0.905
cc_1113 ( N_noxref_7_c_1691_p N_noxref_18_M12_noxref_d ) capacitor \
 c=0.0065582f //x=20.015 //y=1.56 //x2=20.09 //y2=0.905
cc_1114 ( N_noxref_7_c_1722_p N_noxref_18_M12_noxref_d ) capacitor \
 c=0.00241102f //x=20.39 //y=0.75 //x2=20.09 //y2=0.905
cc_1115 ( N_noxref_7_c_1709_p N_noxref_18_M12_noxref_d ) capacitor \
 c=0.0138845f //x=20.39 //y=1.405 //x2=20.09 //y2=0.905
cc_1116 ( N_noxref_7_c_1696_p N_noxref_18_M12_noxref_d ) capacitor \
 c=0.00132245f //x=20.545 //y=0.905 //x2=20.09 //y2=0.905
cc_1117 ( N_noxref_7_c_1699_p N_noxref_18_M12_noxref_d ) capacitor \
 c=0.00566463f //x=20.545 //y=1.25 //x2=20.09 //y2=0.905
cc_1118 ( N_noxref_7_c_1716_p N_noxref_18_M12_noxref_d ) capacitor \
 c=0.00660593f //x=19.98 //y=1.915 //x2=20.09 //y2=0.905
cc_1119 ( N_noxref_7_M37_noxref_g N_noxref_18_M37_noxref_d ) capacitor \
 c=0.0173476f //x=20.02 //y=6.02 //x2=20.095 //y2=5.02
cc_1120 ( N_noxref_7_M38_noxref_g N_noxref_18_M37_noxref_d ) capacitor \
 c=0.0179769f //x=20.46 //y=6.02 //x2=20.095 //y2=5.02
cc_1121 ( N_noxref_7_c_1387_n N_noxref_19_c_2407_n ) capacitor c=0.00121629f \
 //x=19.865 //y=4.07 //x2=18.825 //y2=1.495
cc_1122 ( N_noxref_7_c_1387_n N_noxref_19_c_2390_n ) capacitor c=0.00725714f \
 //x=19.865 //y=4.07 //x2=19.71 //y2=1.58
cc_1123 ( N_noxref_7_c_1387_n N_noxref_19_c_2397_n ) capacitor c=0.00122289f \
 //x=19.865 //y=4.07 //x2=19.795 //y2=1.495
cc_1124 ( N_noxref_7_c_1691_p N_noxref_19_c_2397_n ) capacitor c=0.00623646f \
 //x=20.015 //y=1.56 //x2=19.795 //y2=1.495
cc_1125 ( N_noxref_7_c_1683_p N_noxref_19_c_2397_n ) capacitor c=0.00176439f \
 //x=19.98 //y=2.08 //x2=19.795 //y2=1.495
cc_1126 ( N_noxref_7_c_1394_n N_noxref_19_c_2398_n ) capacitor c=0.00161845f \
 //x=19.98 //y=2.08 //x2=20.68 //y2=0.53
cc_1127 ( N_noxref_7_c_1688_p N_noxref_19_c_2398_n ) capacitor c=0.0186143f \
 //x=20.015 //y=0.905 //x2=20.68 //y2=0.53
cc_1128 ( N_noxref_7_c_1696_p N_noxref_19_c_2398_n ) capacitor c=0.00656458f \
 //x=20.545 //y=0.905 //x2=20.68 //y2=0.53
cc_1129 ( N_noxref_7_c_1683_p N_noxref_19_c_2398_n ) capacitor c=2.1838e-19 \
 //x=19.98 //y=2.08 //x2=20.68 //y2=0.53
cc_1130 ( N_noxref_7_c_1688_p N_noxref_19_M11_noxref_s ) capacitor \
 c=0.00623646f //x=20.015 //y=0.905 //x2=18.69 //y2=0.365
cc_1131 ( N_noxref_7_c_1696_p N_noxref_19_M11_noxref_s ) capacitor \
 c=0.0143002f //x=20.545 //y=0.905 //x2=18.69 //y2=0.365
cc_1132 ( N_noxref_7_c_1699_p N_noxref_19_M11_noxref_s ) capacitor \
 c=0.00290153f //x=20.545 //y=1.25 //x2=18.69 //y2=0.365
cc_1133 ( N_noxref_8_c_1748_n N_noxref_9_c_1788_n ) capacitor c=0.0136048f \
 //x=2.445 //y=0.54 //x2=3.015 //y2=0.995
cc_1134 ( N_noxref_8_c_1759_n N_noxref_9_c_1788_n ) capacitor c=0.0102225f \
 //x=2.445 //y=1.59 //x2=3.015 //y2=0.995
cc_1135 ( N_noxref_8_M0_noxref_s N_noxref_9_c_1788_n ) capacitor c=0.0228676f \
 //x=0.455 //y=0.375 //x2=3.015 //y2=0.995
cc_1136 ( N_noxref_8_M0_noxref_s N_noxref_9_c_1790_n ) capacitor c=0.0180035f \
 //x=0.455 //y=0.375 //x2=3.1 //y2=0.625
cc_1137 ( N_noxref_8_c_1748_n N_noxref_9_M1_noxref_d ) capacitor c=0.0129526f \
 //x=2.445 //y=0.54 //x2=1.86 //y2=0.91
cc_1138 ( N_noxref_8_c_1759_n N_noxref_9_M1_noxref_d ) capacitor c=0.00908243f \
 //x=2.445 //y=1.59 //x2=1.86 //y2=0.91
cc_1139 ( N_noxref_8_M0_noxref_s N_noxref_9_M1_noxref_d ) capacitor \
 c=0.0159202f //x=0.455 //y=0.375 //x2=1.86 //y2=0.91
cc_1140 ( N_noxref_8_M0_noxref_s N_noxref_9_M2_noxref_s ) capacitor \
 c=0.0213553f //x=0.455 //y=0.375 //x2=2.965 //y2=0.375
cc_1141 ( N_noxref_9_c_1796_n N_noxref_11_M3_noxref_s ) capacitor \
 c=0.00164795f //x=4.07 //y=0.625 //x2=5.37 //y2=0.365
cc_1142 ( N_noxref_10_c_1862_n N_noxref_11_c_1921_n ) capacitor c=0.00623646f \
 //x=6.695 //y=1.56 //x2=6.475 //y2=1.495
cc_1143 ( N_noxref_10_c_1871_n N_noxref_11_c_1921_n ) capacitor c=0.00176439f \
 //x=6.66 //y=2.08 //x2=6.475 //y2=1.495
cc_1144 ( N_noxref_10_c_1841_n N_noxref_11_c_1922_n ) capacitor c=0.00159897f \
 //x=6.66 //y=2.08 //x2=7.36 //y2=0.53
cc_1145 ( N_noxref_10_c_1860_n N_noxref_11_c_1922_n ) capacitor c=0.0188655f \
 //x=6.695 //y=0.905 //x2=7.36 //y2=0.53
cc_1146 ( N_noxref_10_c_1868_n N_noxref_11_c_1922_n ) capacitor c=0.00656458f \
 //x=7.225 //y=0.905 //x2=7.36 //y2=0.53
cc_1147 ( N_noxref_10_c_1871_n N_noxref_11_c_1922_n ) capacitor c=2.1838e-19 \
 //x=6.66 //y=2.08 //x2=7.36 //y2=0.53
cc_1148 ( N_noxref_10_c_1860_n N_noxref_11_M3_noxref_s ) capacitor \
 c=0.00623646f //x=6.695 //y=0.905 //x2=5.37 //y2=0.365
cc_1149 ( N_noxref_10_c_1868_n N_noxref_11_M3_noxref_s ) capacitor \
 c=0.0143002f //x=7.225 //y=0.905 //x2=5.37 //y2=0.365
cc_1150 ( N_noxref_10_c_1869_n N_noxref_11_M3_noxref_s ) capacitor \
 c=0.00290153f //x=7.225 //y=1.25 //x2=5.37 //y2=0.365
cc_1151 ( N_noxref_11_c_1925_n N_noxref_12_M5_noxref_s ) capacitor \
 c=0.00174327f //x=7.445 //y=0.615 //x2=8.7 //y2=0.365
cc_1152 ( N_noxref_12_c_1977_n N_noxref_13_M7_noxref_s ) capacitor \
 c=0.00174327f //x=10.775 //y=0.615 //x2=12.03 //y2=0.365
cc_1153 ( N_noxref_13_c_2030_n N_noxref_16_M9_noxref_s ) capacitor \
 c=0.00174327f //x=14.105 //y=0.615 //x2=15.36 //y2=0.365
cc_1154 ( N_noxref_14_c_2081_n N_noxref_15_c_2146_n ) capacitor c=0.0129927f \
 //x=16.65 //y=4.535 //x2=16.825 //y2=5.2
cc_1155 ( N_noxref_14_M33_noxref_g N_noxref_15_c_2146_n ) capacitor \
 c=0.0166421f //x=16.69 //y=6.02 //x2=16.825 //y2=5.2
cc_1156 ( N_noxref_14_c_2101_n N_noxref_15_c_2146_n ) capacitor c=0.00346635f \
 //x=16.68 //y=4.7 //x2=16.825 //y2=5.2
cc_1157 ( N_noxref_14_M34_noxref_g N_noxref_15_c_2152_n ) capacitor \
 c=0.0199348f //x=17.13 //y=6.02 //x2=17.305 //y2=5.2
cc_1158 ( N_noxref_14_c_2112_p N_noxref_15_c_2141_n ) capacitor c=0.00359704f \
 //x=17.06 //y=1.405 //x2=17.305 //y2=1.655
cc_1159 ( N_noxref_14_c_2098_n N_noxref_15_c_2141_n ) capacitor c=0.00457401f \
 //x=17.215 //y=1.25 //x2=17.305 //y2=1.655
cc_1160 ( N_noxref_14_c_2081_n N_noxref_15_c_2142_n ) capacitor c=0.0101284f \
 //x=16.65 //y=4.535 //x2=17.39 //y2=5.115
cc_1161 ( N_noxref_14_c_2072_n N_noxref_15_c_2142_n ) capacitor c=0.080318f \
 //x=16.65 //y=2.08 //x2=17.39 //y2=5.115
cc_1162 ( N_noxref_14_c_2106_n N_noxref_15_c_2142_n ) capacitor c=0.0142673f \
 //x=17.055 //y=4.79 //x2=17.39 //y2=5.115
cc_1163 ( N_noxref_14_c_2099_n N_noxref_15_c_2142_n ) capacitor c=0.00877984f \
 //x=16.65 //y=2.08 //x2=17.39 //y2=5.115
cc_1164 ( N_noxref_14_c_2118_p N_noxref_15_c_2142_n ) capacitor c=0.00306024f \
 //x=16.65 //y=1.915 //x2=17.39 //y2=5.115
cc_1165 ( N_noxref_14_c_2101_n N_noxref_15_c_2142_n ) capacitor c=0.00533692f \
 //x=16.68 //y=4.7 //x2=17.39 //y2=5.115
cc_1166 ( N_noxref_14_c_2106_n N_noxref_15_c_2193_n ) capacitor c=0.00408717f \
 //x=17.055 //y=4.79 //x2=16.91 //y2=5.2
cc_1167 ( N_noxref_14_c_2089_n N_noxref_15_M10_noxref_d ) capacitor \
 c=0.00217566f //x=16.685 //y=0.905 //x2=16.76 //y2=0.905
cc_1168 ( N_noxref_14_c_2092_n N_noxref_15_M10_noxref_d ) capacitor \
 c=0.0034598f //x=16.685 //y=1.25 //x2=16.76 //y2=0.905
cc_1169 ( N_noxref_14_c_2094_n N_noxref_15_M10_noxref_d ) capacitor \
 c=0.0065582f //x=16.685 //y=1.56 //x2=16.76 //y2=0.905
cc_1170 ( N_noxref_14_c_2124_p N_noxref_15_M10_noxref_d ) capacitor \
 c=0.00241102f //x=17.06 //y=0.75 //x2=16.76 //y2=0.905
cc_1171 ( N_noxref_14_c_2112_p N_noxref_15_M10_noxref_d ) capacitor \
 c=0.0138845f //x=17.06 //y=1.405 //x2=16.76 //y2=0.905
cc_1172 ( N_noxref_14_c_2097_n N_noxref_15_M10_noxref_d ) capacitor \
 c=0.00132245f //x=17.215 //y=0.905 //x2=16.76 //y2=0.905
cc_1173 ( N_noxref_14_c_2098_n N_noxref_15_M10_noxref_d ) capacitor \
 c=0.00566463f //x=17.215 //y=1.25 //x2=16.76 //y2=0.905
cc_1174 ( N_noxref_14_c_2118_p N_noxref_15_M10_noxref_d ) capacitor \
 c=0.00660593f //x=16.65 //y=1.915 //x2=16.76 //y2=0.905
cc_1175 ( N_noxref_14_M33_noxref_g N_noxref_15_M33_noxref_d ) capacitor \
 c=0.0173476f //x=16.69 //y=6.02 //x2=16.765 //y2=5.02
cc_1176 ( N_noxref_14_M34_noxref_g N_noxref_15_M33_noxref_d ) capacitor \
 c=0.0179769f //x=17.13 //y=6.02 //x2=16.765 //y2=5.02
cc_1177 ( N_noxref_14_c_2094_n N_noxref_16_c_2220_n ) capacitor c=0.00623646f \
 //x=16.685 //y=1.56 //x2=16.465 //y2=1.495
cc_1178 ( N_noxref_14_c_2099_n N_noxref_16_c_2220_n ) capacitor c=0.00176439f \
 //x=16.65 //y=2.08 //x2=16.465 //y2=1.495
cc_1179 ( N_noxref_14_c_2072_n N_noxref_16_c_2221_n ) capacitor c=0.00161845f \
 //x=16.65 //y=2.08 //x2=17.35 //y2=0.53
cc_1180 ( N_noxref_14_c_2089_n N_noxref_16_c_2221_n ) capacitor c=0.0186143f \
 //x=16.685 //y=0.905 //x2=17.35 //y2=0.53
cc_1181 ( N_noxref_14_c_2097_n N_noxref_16_c_2221_n ) capacitor c=0.00656458f \
 //x=17.215 //y=0.905 //x2=17.35 //y2=0.53
cc_1182 ( N_noxref_14_c_2099_n N_noxref_16_c_2221_n ) capacitor c=2.1838e-19 \
 //x=16.65 //y=2.08 //x2=17.35 //y2=0.53
cc_1183 ( N_noxref_14_c_2089_n N_noxref_16_M9_noxref_s ) capacitor \
 c=0.00623646f //x=16.685 //y=0.905 //x2=15.36 //y2=0.365
cc_1184 ( N_noxref_14_c_2097_n N_noxref_16_M9_noxref_s ) capacitor \
 c=0.0143002f //x=17.215 //y=0.905 //x2=15.36 //y2=0.365
cc_1185 ( N_noxref_14_c_2098_n N_noxref_16_M9_noxref_s ) capacitor \
 c=0.00290153f //x=17.215 //y=1.25 //x2=15.36 //y2=0.365
cc_1186 ( N_noxref_14_c_2072_n N_noxref_17_c_2265_n ) capacitor c=0.00105994f \
 //x=16.65 //y=2.08 //x2=19.24 //y2=2.08
cc_1187 ( N_noxref_15_c_2177_n N_noxref_16_c_2232_n ) capacitor c=3.15806e-19 \
 //x=17.035 //y=1.655 //x2=15.495 //y2=1.495
cc_1188 ( N_noxref_15_c_2177_n N_noxref_16_c_2220_n ) capacitor c=0.0203424f \
 //x=17.035 //y=1.655 //x2=16.465 //y2=1.495
cc_1189 ( N_noxref_15_c_2141_n N_noxref_16_c_2221_n ) capacitor c=0.00469114f \
 //x=17.305 //y=1.655 //x2=17.35 //y2=0.53
cc_1190 ( N_noxref_15_M10_noxref_d N_noxref_16_c_2221_n ) capacitor \
 c=0.0118355f //x=16.76 //y=0.905 //x2=17.35 //y2=0.53
cc_1191 ( N_noxref_15_c_2141_n N_noxref_16_M9_noxref_s ) capacitor \
 c=0.0143484f //x=17.305 //y=1.655 //x2=15.36 //y2=0.365
cc_1192 ( N_noxref_15_M10_noxref_d N_noxref_16_M9_noxref_s ) capacitor \
 c=0.043966f //x=16.76 //y=0.905 //x2=15.36 //y2=0.365
cc_1193 ( N_noxref_15_c_2142_n N_noxref_17_c_2265_n ) capacitor c=0.0166833f \
 //x=17.39 //y=5.115 //x2=19.24 //y2=2.08
cc_1194 ( N_noxref_15_c_2142_n N_noxref_18_c_2326_n ) capacitor c=3.49822e-19 \
 //x=17.39 //y=5.115 //x2=20.72 //y2=5.115
cc_1195 ( N_noxref_15_c_2141_n N_noxref_19_c_2407_n ) capacitor c=3.22188e-19 \
 //x=17.305 //y=1.655 //x2=18.825 //y2=1.495
cc_1196 ( N_noxref_16_c_2224_n N_noxref_19_M11_noxref_s ) capacitor \
 c=0.00174327f //x=17.435 //y=0.615 //x2=18.69 //y2=0.365
cc_1197 ( N_noxref_17_M36_noxref_g N_noxref_18_c_2330_n ) capacitor \
 c=0.017965f //x=19.58 //y=6.02 //x2=20.155 //y2=5.2
cc_1198 ( N_noxref_17_c_2265_n N_noxref_18_c_2334_n ) capacitor c=0.00549854f \
 //x=19.24 //y=2.08 //x2=19.445 //y2=5.2
cc_1199 ( N_noxref_17_M35_noxref_g N_noxref_18_c_2334_n ) capacitor \
 c=0.0177326f //x=19.14 //y=6.02 //x2=19.445 //y2=5.2
cc_1200 ( N_noxref_17_c_2283_n N_noxref_18_c_2334_n ) capacitor c=0.00569763f \
 //x=19.24 //y=4.7 //x2=19.445 //y2=5.2
cc_1201 ( N_noxref_17_c_2265_n N_noxref_18_c_2326_n ) capacitor c=0.00413825f \
 //x=19.24 //y=2.08 //x2=20.72 //y2=5.115
cc_1202 ( N_noxref_17_M36_noxref_g N_noxref_18_M35_noxref_d ) capacitor \
 c=0.0173476f //x=19.58 //y=6.02 //x2=19.215 //y2=5.02
cc_1203 ( N_noxref_17_c_2270_n N_noxref_19_c_2407_n ) capacitor c=0.0034165f \
 //x=19.045 //y=1.915 //x2=18.825 //y2=1.495
cc_1204 ( N_noxref_17_c_2265_n N_noxref_19_c_2390_n ) capacitor c=0.0123126f \
 //x=19.24 //y=2.08 //x2=19.71 //y2=1.58
cc_1205 ( N_noxref_17_c_2269_n N_noxref_19_c_2390_n ) capacitor c=0.00703567f \
 //x=19.045 //y=1.52 //x2=19.71 //y2=1.58
cc_1206 ( N_noxref_17_c_2270_n N_noxref_19_c_2390_n ) capacitor c=0.0210414f \
 //x=19.045 //y=1.915 //x2=19.71 //y2=1.58
cc_1207 ( N_noxref_17_c_2272_n N_noxref_19_c_2390_n ) capacitor c=0.00780629f \
 //x=19.42 //y=1.365 //x2=19.71 //y2=1.58
cc_1208 ( N_noxref_17_c_2275_n N_noxref_19_c_2390_n ) capacitor c=0.00339872f \
 //x=19.575 //y=1.21 //x2=19.71 //y2=1.58
cc_1209 ( N_noxref_17_c_2270_n N_noxref_19_c_2397_n ) capacitor c=6.71402e-19 \
 //x=19.045 //y=1.915 //x2=19.795 //y2=1.495
cc_1210 ( N_noxref_17_c_2266_n N_noxref_19_M11_noxref_s ) capacitor \
 c=0.0326577f //x=19.045 //y=0.865 //x2=18.69 //y2=0.365
cc_1211 ( N_noxref_17_c_2269_n N_noxref_19_M11_noxref_s ) capacitor \
 c=3.48408e-19 //x=19.045 //y=1.52 //x2=18.69 //y2=0.365
cc_1212 ( N_noxref_17_c_2273_n N_noxref_19_M11_noxref_s ) capacitor \
 c=0.0120759f //x=19.575 //y=0.865 //x2=18.69 //y2=0.365
cc_1213 ( N_noxref_18_c_2384_p N_noxref_19_c_2407_n ) capacitor c=3.15806e-19 \
 //x=20.365 //y=1.655 //x2=18.825 //y2=1.495
cc_1214 ( N_noxref_18_c_2384_p N_noxref_19_c_2397_n ) capacitor c=0.0203424f \
 //x=20.365 //y=1.655 //x2=19.795 //y2=1.495
cc_1215 ( N_noxref_18_c_2325_n N_noxref_19_c_2398_n ) capacitor c=0.00469114f \
 //x=20.635 //y=1.655 //x2=20.68 //y2=0.53
cc_1216 ( N_noxref_18_M12_noxref_d N_noxref_19_c_2398_n ) capacitor \
 c=0.0118355f //x=20.09 //y=0.905 //x2=20.68 //y2=0.53
cc_1217 ( N_noxref_18_c_2325_n N_noxref_19_M11_noxref_s ) capacitor \
 c=0.0144625f //x=20.635 //y=1.655 //x2=18.69 //y2=0.365
cc_1218 ( N_noxref_18_M12_noxref_d N_noxref_19_M11_noxref_s ) capacitor \
 c=0.043966f //x=20.09 //y=0.905 //x2=18.69 //y2=0.365
