VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AND3X1
  CLASS CORE ;
  FOREIGN AND3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.810 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.771900 ;
    PORT
      LAYER li1 ;
        RECT 5.840 4.665 6.010 7.020 ;
        RECT 5.840 4.495 6.375 4.665 ;
        RECT 6.205 2.165 6.375 4.495 ;
        RECT 5.835 1.995 6.375 2.165 ;
        RECT 5.835 0.840 6.005 1.995 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.915 1.195 4.865 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.014850 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.915 2.305 4.865 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 3.245 1.915 3.415 4.865 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 7.465 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 7.200 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.005 5.215 1.175 7.230 ;
        RECT 1.885 5.555 2.055 7.230 ;
        RECT 2.765 5.555 2.935 7.230 ;
        RECT 3.645 5.555 3.815 7.230 ;
        RECT 4.640 4.110 4.980 7.230 ;
        RECT 5.400 5.185 5.570 7.230 ;
        RECT 6.280 5.185 6.450 7.230 ;
        RECT 6.860 4.110 7.200 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 7.200 7.570 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 7.200 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.990 0.170 1.160 1.130 ;
        RECT 4.640 0.170 4.980 2.720 ;
        RECT 5.355 0.620 5.525 1.750 ;
        RECT 6.325 0.620 6.495 1.750 ;
        RECT 5.355 0.450 6.495 0.620 ;
        RECT 5.355 0.170 5.525 0.450 ;
        RECT 5.840 0.170 6.010 0.450 ;
        RECT 6.325 0.170 6.495 0.450 ;
        RECT 6.860 0.170 7.200 2.720 ;
        RECT -0.170 -0.170 7.200 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 7.200 0.170 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 1.445 5.240 1.615 7.020 ;
        RECT 2.325 5.240 2.495 7.020 ;
        RECT 3.205 5.240 3.375 7.020 ;
        RECT 1.445 5.070 4.155 5.240 ;
        RECT 0.505 1.675 0.675 1.755 ;
        RECT 1.475 1.675 1.645 1.755 ;
        RECT 2.445 1.675 2.615 1.755 ;
        RECT 0.505 1.505 2.615 1.675 ;
        RECT 0.505 0.375 0.675 1.505 ;
        RECT 1.475 0.625 1.645 1.505 ;
        RECT 2.445 1.425 2.615 1.505 ;
        RECT 1.965 1.080 2.135 1.160 ;
        RECT 3.015 1.080 3.185 1.755 ;
        RECT 3.985 1.750 4.155 5.070 ;
        RECT 5.465 1.920 5.635 4.865 ;
        RECT 1.965 0.910 3.185 1.080 ;
        RECT 1.965 0.830 2.135 0.910 ;
        RECT 2.445 0.625 2.615 0.705 ;
        RECT 1.475 0.455 2.615 0.625 ;
        RECT 1.475 0.375 1.645 0.455 ;
        RECT 2.445 0.375 2.615 0.455 ;
        RECT 3.015 0.625 3.185 0.910 ;
        RECT 3.500 1.580 4.155 1.750 ;
        RECT 3.500 0.845 3.670 1.580 ;
        RECT 3.985 0.625 4.155 1.395 ;
        RECT 3.015 0.455 4.155 0.625 ;
        RECT 3.015 0.375 3.185 0.455 ;
        RECT 3.985 0.375 4.155 0.455 ;
      LAYER mcon ;
        RECT 3.985 3.245 4.155 3.415 ;
        RECT 5.465 3.245 5.635 3.415 ;
      LAYER met1 ;
        RECT 3.955 3.415 4.185 3.445 ;
        RECT 5.435 3.415 5.665 3.445 ;
        RECT 3.925 3.245 5.695 3.415 ;
        RECT 3.955 3.215 4.185 3.245 ;
        RECT 5.435 3.215 5.665 3.245 ;
  END
END AND3X1
END LIBRARY

