magic
tech sky130A
magscale 1 2
timestamp 1652393989
<< nwell >>
rect 55 1463 89 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 1833 944 1867 979
rect 131 871 165 905
rect 871 871 905 905
rect 1167 871 1201 905
rect 1463 871 1497 905
rect 1685 871 1719 905
rect 1833 870 1867 905
rect 131 797 165 831
rect 353 797 387 831
rect 1685 797 1719 831
rect 1833 796 1867 831
rect 131 723 165 757
rect 353 723 387 757
rect 871 723 905 757
rect 1167 723 1201 757
rect 1463 723 1497 757
rect 1685 723 1719 757
rect 1833 722 1867 757
rect 131 649 165 683
rect 353 649 387 683
rect 871 649 905 683
rect 1167 649 1201 683
rect 1463 649 1497 683
rect 1685 649 1719 683
rect 1833 648 1867 683
rect 131 575 165 609
rect 353 575 387 609
rect 871 575 905 609
rect 1167 575 1201 609
rect 1463 575 1497 609
rect 1685 575 1719 609
rect 1833 574 1867 609
rect 131 501 165 535
rect 353 501 387 535
rect 871 501 905 535
rect 1167 501 1201 535
rect 1463 501 1497 535
rect 1685 501 1719 535
rect 1833 500 1867 535
rect 1833 426 1867 461
<< metal1 >>
rect -34 1446 2032 1514
rect -34 -34 2032 34
use votern3x1_pcell  votern3x1_pcell_0 pcells
timestamp 1652393950
transform 1 0 0 0 1 0
box -87 -34 2085 1550
<< labels >>
rlabel locali 1833 649 1867 683 1 YN
port 1 nsew signal output
rlabel locali 1833 723 1867 757 1 YN
port 1 nsew signal output
rlabel locali 1833 797 1867 831 1 YN
port 1 nsew signal output
rlabel locali 1833 871 1867 905 1 YN
port 1 nsew signal output
rlabel locali 1833 945 1867 979 1 YN
port 1 nsew signal output
rlabel locali 1833 575 1867 609 1 YN
port 1 nsew signal output
rlabel locali 1833 501 1867 535 1 YN
port 1 nsew signal output
rlabel locali 1833 427 1867 461 1 YN
port 1 nsew signal output
rlabel locali 353 723 387 757 1 A
port 2 nsew signal input
rlabel locali 353 797 387 831 1 A
port 2 nsew signal input
rlabel locali 353 649 387 683 1 A
port 2 nsew signal input
rlabel locali 353 575 387 609 1 A
port 2 nsew signal input
rlabel locali 353 501 387 535 1 A
port 2 nsew signal input
rlabel locali 1685 501 1719 535 1 A
port 2 nsew signal input
rlabel locali 1685 575 1719 609 1 A
port 2 nsew signal input
rlabel locali 1685 649 1719 683 1 A
port 2 nsew signal input
rlabel locali 1685 723 1719 757 1 A
port 2 nsew signal input
rlabel locali 1685 797 1719 831 1 A
port 2 nsew signal input
rlabel locali 1685 871 1719 905 1 A
port 2 nsew signal input
rlabel locali 131 797 165 831 1 B
port 3 nsew signal input
rlabel locali 131 723 165 757 1 B
port 3 nsew signal input
rlabel locali 131 649 165 683 1 B
port 3 nsew signal input
rlabel locali 131 575 165 609 1 B
port 3 nsew signal input
rlabel locali 131 501 165 535 1 B
port 3 nsew signal input
rlabel locali 871 723 905 757 1 B
port 3 nsew signal input
rlabel locali 871 649 905 683 1 B
port 3 nsew signal input
rlabel locali 871 575 905 609 1 B
port 3 nsew signal input
rlabel locali 871 501 905 535 1 B
port 3 nsew signal input
rlabel locali 131 871 165 905 1 B
port 3 nsew signal input
rlabel locali 871 871 905 905 1 B
port 3 nsew signal input
rlabel locali 1167 501 1201 535 1 C
port 4 nsew signal input
rlabel locali 1167 575 1201 609 1 C
port 4 nsew signal input
rlabel locali 1167 649 1201 683 1 C
port 4 nsew signal input
rlabel locali 1167 723 1201 757 1 C
port 4 nsew signal input
rlabel locali 1167 871 1201 905 1 C
port 4 nsew signal input
rlabel locali 1463 723 1497 757 1 C
port 4 nsew signal input
rlabel locali 1463 649 1497 683 1 C
port 4 nsew signal input
rlabel locali 1463 575 1497 609 1 C
port 4 nsew signal input
rlabel locali 1463 501 1497 535 1 C
port 4 nsew signal input
rlabel locali 1463 871 1497 905 1 C
port 4 nsew signal input
rlabel metal1 -34 1446 2032 1514 1 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 -34 -34 2032 34 1 VGND
port 5 nsew ground bidirectional abutment
rlabel nwell 55 1463 89 1497 1 VPB
port 5 nsew power bidirectional
rlabel pwell 57 -17 91 17 1 VNB
port 5 nsew ground bidirectional
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1998 1480
string LEFsymmetry X Y R90
<< end >>
