* SPICE3 file created from DFFRNX1.ext - technology: sky130A

.subckt DFFRNX1 Q QN D RN VPB VNB
M1000 QN Q a_3924_182.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1001 VPB.t26 a_147_159.t7 a_277_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_599_943.t4 a_1304_166# VPB.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t31 a_599_943.t7 a_2141_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPB.t17 RN a_277_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPB.t28 a_277_1004.t8 QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=1.74p ps=13.74u
M1006 a_599_943.t2 RN VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 QN Q VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_147_159.t5 RN VPB.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 Q QN VPB.t1 pshort w=2u l=0.15u
+  ad=1.16p pd=9.16u as=0p ps=0u
M1010 VNB QN a_4626_73.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1011 VNB a_147_159.t14 a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB.t7 a_599_943.t9 a_277_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPB.t24 a_147_159.t8 a_2141_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VNB a_599_943.t8 a_2036_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPB.t5 a_2141_1004.t6 a_147_159.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_147_159.t2 RN VPB.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 Q a_147_159.t9 VPB.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_277_1004.t6 a_147_159.t10 VPB.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VNB a_277_1004.t7 a_3643_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPB.t29 a_277_1004.t10 a_599_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPB.t18 RN a_599_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t3 Q QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VNB a_2141_1004.t5 a_2681_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_277_1004.t3 RN VPB.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_2141_1004.t0 a_599_943.t10 VPB.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 QN a_277_1004.t11 VPB.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPB.t20 a_1304_166# a_599_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPB.t10 RN QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 Q a_147_159.t11 a_4626_73.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1030 a_599_943.t5 a_277_1004.t12 VPB.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_277_1004.t1 a_599_943.t11 VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_2141_1004.t3 a_147_159.t13 VPB.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 QN RN VPB.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_147_159.t0 a_2141_1004.t7 VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 VNB a_277_1004.t9 a_1053_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPB.t13 RN a_147_159.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPB.t0 QN Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPB.t12 RN a_147_159.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPB.t21 a_147_159.t15 Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u








R0 a_147_159.n10 a_147_159.t7 512.525
R1 a_147_159.n8 a_147_159.t8 472.359
R2 a_147_159.n6 a_147_159.t15 472.359
R3 a_147_159.n8 a_147_159.t13 384.527
R4 a_147_159.n6 a_147_159.t9 384.527
R5 a_147_159.n10 a_147_159.t10 371.139
R6 a_147_159.n11 a_147_159.t14 324.268
R7 a_147_159.n9 a_147_159.t12 277.772
R8 a_147_159.n7 a_147_159.t11 277.772
R9 a_147_159.n16 a_147_159.n14 249.704
R10 a_147_159.n14 a_147_159.n5 127.74
R11 a_147_159.n11 a_147_159.n10 119.654
R12 a_147_159.n12 a_147_159.n11 83.572
R13 a_147_159.n13 a_147_159.n7 81.396
R14 a_147_159.n4 a_147_159.n3 79.232
R15 a_147_159.n12 a_147_159.n9 76
R16 a_147_159.n14 a_147_159.n13 76
R17 a_147_159.n9 a_147_159.n8 67.001
R18 a_147_159.n7 a_147_159.n6 67.001
R19 a_147_159.n5 a_147_159.n4 63.152
R20 a_147_159.n16 a_147_159.n15 30
R21 a_147_159.n17 a_147_159.n0 24.383
R22 a_147_159.n17 a_147_159.n16 23.684
R23 a_147_159.n5 a_147_159.n1 16.08
R24 a_147_159.n4 a_147_159.n2 16.08
R25 a_147_159.n1 a_147_159.t4 14.282
R26 a_147_159.n1 a_147_159.t2 14.282
R27 a_147_159.n2 a_147_159.t3 14.282
R28 a_147_159.n2 a_147_159.t5 14.282
R29 a_147_159.n3 a_147_159.t1 14.282
R30 a_147_159.n3 a_147_159.t0 14.282
R31 a_147_159.n13 a_147_159.n12 4.035
R32 a_277_1004.n7 a_277_1004.t10 512.525
R33 a_277_1004.n5 a_277_1004.t8 512.525
R34 a_277_1004.n7 a_277_1004.t12 371.139
R35 a_277_1004.n5 a_277_1004.t11 371.139
R36 a_277_1004.n8 a_277_1004.t9 297.715
R37 a_277_1004.n6 a_277_1004.t7 297.715
R38 a_277_1004.n12 a_277_1004.n10 229.673
R39 a_277_1004.n10 a_277_1004.n4 154.293
R40 a_277_1004.n8 a_277_1004.n7 146.207
R41 a_277_1004.n6 a_277_1004.n5 146.207
R42 a_277_1004.n9 a_277_1004.n6 85.476
R43 a_277_1004.n3 a_277_1004.n2 79.232
R44 a_277_1004.n10 a_277_1004.n9 77.315
R45 a_277_1004.n9 a_277_1004.n8 76
R46 a_277_1004.n4 a_277_1004.n3 63.152
R47 a_277_1004.n4 a_277_1004.n0 16.08
R48 a_277_1004.n3 a_277_1004.n1 16.08
R49 a_277_1004.n12 a_277_1004.n11 15.218
R50 a_277_1004.n0 a_277_1004.t2 14.282
R51 a_277_1004.n0 a_277_1004.t1 14.282
R52 a_277_1004.n1 a_277_1004.t4 14.282
R53 a_277_1004.n1 a_277_1004.t3 14.282
R54 a_277_1004.n2 a_277_1004.t5 14.282
R55 a_277_1004.n2 a_277_1004.t6 14.282
R56 a_277_1004.n13 a_277_1004.n12 12.014
R57 VPB VPB.n473 126.832
R58 VPB.n40 VPB.n38 94.117
R59 VPB.n395 VPB.n393 94.117
R60 VPB.n332 VPB.n330 94.117
R61 VPB.n129 VPB.n127 94.117
R62 VPB.n255 VPB.n253 94.117
R63 VPB.n268 VPB.n267 80.104
R64 VPB.n139 VPB.n138 80.104
R65 VPB.n408 VPB.n407 80.104
R66 VPB.n50 VPB.n49 80.104
R67 VPB.n216 VPB.n215 76
R68 VPB.n221 VPB.n220 76
R69 VPB.n226 VPB.n225 76
R70 VPB.n230 VPB.n229 76
R71 VPB.n257 VPB.n256 76
R72 VPB.n261 VPB.n260 76
R73 VPB.n266 VPB.n265 76
R74 VPB.n271 VPB.n270 76
R75 VPB.n278 VPB.n277 76
R76 VPB.n283 VPB.n282 76
R77 VPB.n288 VPB.n287 76
R78 VPB.n295 VPB.n294 76
R79 VPB.n300 VPB.n299 76
R80 VPB.n305 VPB.n304 76
R81 VPB.n309 VPB.n308 76
R82 VPB.n313 VPB.n312 76
R83 VPB.n328 VPB.n325 76
R84 VPB.n334 VPB.n333 76
R85 VPB.n339 VPB.n338 76
R86 VPB.n344 VPB.n343 76
R87 VPB.n351 VPB.n350 76
R88 VPB.n356 VPB.n355 76
R89 VPB.n361 VPB.n360 76
R90 VPB.n366 VPB.n365 76
R91 VPB.n370 VPB.n369 76
R92 VPB.n397 VPB.n396 76
R93 VPB.n401 VPB.n400 76
R94 VPB.n406 VPB.n405 76
R95 VPB.n411 VPB.n410 76
R96 VPB.n418 VPB.n417 76
R97 VPB.n423 VPB.n422 76
R98 VPB.n428 VPB.n427 76
R99 VPB.n435 VPB.n434 76
R100 VPB.n440 VPB.n439 76
R101 VPB.n445 VPB.n444 76
R102 VPB.n449 VPB.n448 76
R103 VPB.n453 VPB.n452 76
R104 VPB.n466 VPB.n465 76
R105 VPB.n297 VPB.n296 75.654
R106 VPB.n161 VPB.n160 75.654
R107 VPB.n437 VPB.n436 75.654
R108 VPB.n72 VPB.n71 75.654
R109 VPB.n22 VPB.n21 61.764
R110 VPB.n377 VPB.n376 61.764
R111 VPB.n88 VPB.n87 61.764
R112 VPB.n111 VPB.n110 61.764
R113 VPB.n237 VPB.n236 61.764
R114 VPB.n78 VPB.t25 55.106
R115 VPB.n441 VPB.t30 55.106
R116 VPB.n362 VPB.t8 55.106
R117 VPB.n167 VPB.t2 55.106
R118 VPB.n301 VPB.t27 55.106
R119 VPB.n222 VPB.t1 55.106
R120 VPB.n45 VPB.t7 55.106
R121 VPB.n402 VPB.t18 55.106
R122 VPB.n335 VPB.t24 55.106
R123 VPB.n134 VPB.t12 55.106
R124 VPB.n262 VPB.t3 55.106
R125 VPB.n205 VPB.t21 55.106
R126 VPB.n202 VPB.n201 48.952
R127 VPB.n275 VPB.n274 48.952
R128 VPB.n143 VPB.n142 48.952
R129 VPB.n341 VPB.n340 48.952
R130 VPB.n415 VPB.n414 48.952
R131 VPB.n54 VPB.n53 48.952
R132 VPB.n218 VPB.n217 44.502
R133 VPB.n292 VPB.n291 44.502
R134 VPB.n157 VPB.n156 44.502
R135 VPB.n358 VPB.n357 44.502
R136 VPB.n432 VPB.n431 44.502
R137 VPB.n68 VPB.n67 44.502
R138 VPB.n66 VPB.n14 40.824
R139 VPB.n57 VPB.n15 40.824
R140 VPB.n430 VPB.n429 40.824
R141 VPB.n413 VPB.n412 40.824
R142 VPB.n346 VPB.n345 40.824
R143 VPB.n155 VPB.n103 40.824
R144 VPB.n146 VPB.n104 40.824
R145 VPB.n290 VPB.n289 40.824
R146 VPB.n273 VPB.n272 40.824
R147 VPB.n196 VPB.n195 40.824
R148 VPB.n210 VPB.n209 35.118
R149 VPB.n470 VPB.n466 20.452
R150 VPB.n194 VPB.n191 20.452
R151 VPB.n198 VPB.n197 17.801
R152 VPB.n280 VPB.n279 17.801
R153 VPB.n148 VPB.n147 17.801
R154 VPB.n348 VPB.n347 17.801
R155 VPB.n420 VPB.n419 17.801
R156 VPB.n59 VPB.n58 17.801
R157 VPB.n14 VPB.t16 14.282
R158 VPB.n14 VPB.t26 14.282
R159 VPB.n15 VPB.t6 14.282
R160 VPB.n15 VPB.t17 14.282
R161 VPB.n429 VPB.t19 14.282
R162 VPB.n429 VPB.t29 14.282
R163 VPB.n412 VPB.t11 14.282
R164 VPB.n412 VPB.t20 14.282
R165 VPB.n345 VPB.t23 14.282
R166 VPB.n345 VPB.t31 14.282
R167 VPB.n103 VPB.t15 14.282
R168 VPB.n103 VPB.t5 14.282
R169 VPB.n104 VPB.t14 14.282
R170 VPB.n104 VPB.t13 14.282
R171 VPB.n289 VPB.t9 14.282
R172 VPB.n289 VPB.t28 14.282
R173 VPB.n272 VPB.t4 14.282
R174 VPB.n272 VPB.t10 14.282
R175 VPB.n195 VPB.t22 14.282
R176 VPB.n195 VPB.t0 14.282
R177 VPB.n194 VPB.n193 13.653
R178 VPB.n193 VPB.n192 13.653
R179 VPB.n208 VPB.n207 13.653
R180 VPB.n207 VPB.n206 13.653
R181 VPB.n204 VPB.n203 13.653
R182 VPB.n203 VPB.n202 13.653
R183 VPB.n200 VPB.n199 13.653
R184 VPB.n199 VPB.n198 13.653
R185 VPB.n215 VPB.n214 13.653
R186 VPB.n214 VPB.n213 13.653
R187 VPB.n220 VPB.n219 13.653
R188 VPB.n219 VPB.n218 13.653
R189 VPB.n225 VPB.n224 13.653
R190 VPB.n224 VPB.n223 13.653
R191 VPB.n229 VPB.n228 13.653
R192 VPB.n228 VPB.n227 13.653
R193 VPB.n256 VPB.n255 13.653
R194 VPB.n255 VPB.n254 13.653
R195 VPB.n260 VPB.n259 13.653
R196 VPB.n259 VPB.n258 13.653
R197 VPB.n265 VPB.n264 13.653
R198 VPB.n264 VPB.n263 13.653
R199 VPB.n270 VPB.n269 13.653
R200 VPB.n269 VPB.n268 13.653
R201 VPB.n277 VPB.n276 13.653
R202 VPB.n276 VPB.n275 13.653
R203 VPB.n282 VPB.n281 13.653
R204 VPB.n281 VPB.n280 13.653
R205 VPB.n287 VPB.n286 13.653
R206 VPB.n286 VPB.n285 13.653
R207 VPB.n294 VPB.n293 13.653
R208 VPB.n293 VPB.n292 13.653
R209 VPB.n299 VPB.n298 13.653
R210 VPB.n298 VPB.n297 13.653
R211 VPB.n304 VPB.n303 13.653
R212 VPB.n303 VPB.n302 13.653
R213 VPB.n308 VPB.n307 13.653
R214 VPB.n307 VPB.n306 13.653
R215 VPB.n312 VPB.n311 13.653
R216 VPB.n311 VPB.n310 13.653
R217 VPB.n130 VPB.n129 13.653
R218 VPB.n129 VPB.n128 13.653
R219 VPB.n133 VPB.n132 13.653
R220 VPB.n132 VPB.n131 13.653
R221 VPB.n137 VPB.n136 13.653
R222 VPB.n136 VPB.n135 13.653
R223 VPB.n141 VPB.n140 13.653
R224 VPB.n140 VPB.n139 13.653
R225 VPB.n145 VPB.n144 13.653
R226 VPB.n144 VPB.n143 13.653
R227 VPB.n150 VPB.n149 13.653
R228 VPB.n149 VPB.n148 13.653
R229 VPB.n154 VPB.n153 13.653
R230 VPB.n153 VPB.n152 13.653
R231 VPB.n159 VPB.n158 13.653
R232 VPB.n158 VPB.n157 13.653
R233 VPB.n163 VPB.n162 13.653
R234 VPB.n162 VPB.n161 13.653
R235 VPB.n166 VPB.n165 13.653
R236 VPB.n165 VPB.n164 13.653
R237 VPB.n170 VPB.n169 13.653
R238 VPB.n169 VPB.n168 13.653
R239 VPB.n328 VPB.n327 13.653
R240 VPB.n327 VPB.n326 13.653
R241 VPB.n333 VPB.n332 13.653
R242 VPB.n332 VPB.n331 13.653
R243 VPB.n338 VPB.n337 13.653
R244 VPB.n337 VPB.n336 13.653
R245 VPB.n343 VPB.n342 13.653
R246 VPB.n342 VPB.n341 13.653
R247 VPB.n350 VPB.n349 13.653
R248 VPB.n349 VPB.n348 13.653
R249 VPB.n355 VPB.n354 13.653
R250 VPB.n354 VPB.n353 13.653
R251 VPB.n360 VPB.n359 13.653
R252 VPB.n359 VPB.n358 13.653
R253 VPB.n365 VPB.n364 13.653
R254 VPB.n364 VPB.n363 13.653
R255 VPB.n369 VPB.n368 13.653
R256 VPB.n368 VPB.n367 13.653
R257 VPB.n396 VPB.n395 13.653
R258 VPB.n395 VPB.n394 13.653
R259 VPB.n400 VPB.n399 13.653
R260 VPB.n399 VPB.n398 13.653
R261 VPB.n405 VPB.n404 13.653
R262 VPB.n404 VPB.n403 13.653
R263 VPB.n410 VPB.n409 13.653
R264 VPB.n409 VPB.n408 13.653
R265 VPB.n417 VPB.n416 13.653
R266 VPB.n416 VPB.n415 13.653
R267 VPB.n422 VPB.n421 13.653
R268 VPB.n421 VPB.n420 13.653
R269 VPB.n427 VPB.n426 13.653
R270 VPB.n426 VPB.n425 13.653
R271 VPB.n434 VPB.n433 13.653
R272 VPB.n433 VPB.n432 13.653
R273 VPB.n439 VPB.n438 13.653
R274 VPB.n438 VPB.n437 13.653
R275 VPB.n444 VPB.n443 13.653
R276 VPB.n443 VPB.n442 13.653
R277 VPB.n448 VPB.n447 13.653
R278 VPB.n447 VPB.n446 13.653
R279 VPB.n452 VPB.n451 13.653
R280 VPB.n451 VPB.n450 13.653
R281 VPB.n41 VPB.n40 13.653
R282 VPB.n40 VPB.n39 13.653
R283 VPB.n44 VPB.n43 13.653
R284 VPB.n43 VPB.n42 13.653
R285 VPB.n48 VPB.n47 13.653
R286 VPB.n47 VPB.n46 13.653
R287 VPB.n52 VPB.n51 13.653
R288 VPB.n51 VPB.n50 13.653
R289 VPB.n56 VPB.n55 13.653
R290 VPB.n55 VPB.n54 13.653
R291 VPB.n61 VPB.n60 13.653
R292 VPB.n60 VPB.n59 13.653
R293 VPB.n65 VPB.n64 13.653
R294 VPB.n64 VPB.n63 13.653
R295 VPB.n70 VPB.n69 13.653
R296 VPB.n69 VPB.n68 13.653
R297 VPB.n74 VPB.n73 13.653
R298 VPB.n73 VPB.n72 13.653
R299 VPB.n77 VPB.n76 13.653
R300 VPB.n76 VPB.n75 13.653
R301 VPB.n81 VPB.n80 13.653
R302 VPB.n80 VPB.n79 13.653
R303 VPB.n466 VPB.n0 13.653
R304 VPB VPB.n0 13.653
R305 VPB.n213 VPB.n212 13.35
R306 VPB.n285 VPB.n284 13.35
R307 VPB.n152 VPB.n151 13.35
R308 VPB.n353 VPB.n352 13.35
R309 VPB.n425 VPB.n424 13.35
R310 VPB.n63 VPB.n62 13.35
R311 VPB.n470 VPB.n469 13.276
R312 VPB.n469 VPB.n467 13.276
R313 VPB.n36 VPB.n18 13.276
R314 VPB.n18 VPB.n16 13.276
R315 VPB.n391 VPB.n373 13.276
R316 VPB.n373 VPB.n371 13.276
R317 VPB.n102 VPB.n84 13.276
R318 VPB.n84 VPB.n82 13.276
R319 VPB.n125 VPB.n107 13.276
R320 VPB.n107 VPB.n105 13.276
R321 VPB.n251 VPB.n233 13.276
R322 VPB.n233 VPB.n231 13.276
R323 VPB.n204 VPB.n200 13.276
R324 VPB.n256 VPB.n252 13.276
R325 VPB.n130 VPB.n126 13.276
R326 VPB.n133 VPB.n130 13.276
R327 VPB.n141 VPB.n137 13.276
R328 VPB.n145 VPB.n141 13.276
R329 VPB.n154 VPB.n150 13.276
R330 VPB.n163 VPB.n159 13.276
R331 VPB.n166 VPB.n163 13.276
R332 VPB.n328 VPB.n170 13.276
R333 VPB.n329 VPB.n328 13.276
R334 VPB.n333 VPB.n329 13.276
R335 VPB.n396 VPB.n392 13.276
R336 VPB.n41 VPB.n37 13.276
R337 VPB.n44 VPB.n41 13.276
R338 VPB.n52 VPB.n48 13.276
R339 VPB.n56 VPB.n52 13.276
R340 VPB.n65 VPB.n61 13.276
R341 VPB.n74 VPB.n70 13.276
R342 VPB.n77 VPB.n74 13.276
R343 VPB.n466 VPB.n81 13.276
R344 VPB.n191 VPB.n173 13.276
R345 VPB.n173 VPB.n171 13.276
R346 VPB.n178 VPB.n176 12.796
R347 VPB.n178 VPB.n177 12.564
R348 VPB.n170 VPB.n167 12.558
R349 VPB.n81 VPB.n78 12.558
R350 VPB.n134 VPB.n133 12.2
R351 VPB.n45 VPB.n44 12.2
R352 VPB.n187 VPB.n186 12.198
R353 VPB.n184 VPB.n183 12.198
R354 VPB.n184 VPB.n181 12.198
R355 VPB.n205 VPB.n204 11.841
R356 VPB.n150 VPB.n146 9.329
R357 VPB.n61 VPB.n57 9.329
R358 VPB.n155 VPB.n154 8.97
R359 VPB.n66 VPB.n65 8.97
R360 VPB.n191 VPB.n190 7.5
R361 VPB.n176 VPB.n175 7.5
R362 VPB.n183 VPB.n182 7.5
R363 VPB.n181 VPB.n180 7.5
R364 VPB.n173 VPB.n172 7.5
R365 VPB.n188 VPB.n174 7.5
R366 VPB.n233 VPB.n232 7.5
R367 VPB.n246 VPB.n245 7.5
R368 VPB.n240 VPB.n239 7.5
R369 VPB.n242 VPB.n241 7.5
R370 VPB.n235 VPB.n234 7.5
R371 VPB.n251 VPB.n250 7.5
R372 VPB.n107 VPB.n106 7.5
R373 VPB.n120 VPB.n119 7.5
R374 VPB.n114 VPB.n113 7.5
R375 VPB.n116 VPB.n115 7.5
R376 VPB.n109 VPB.n108 7.5
R377 VPB.n125 VPB.n124 7.5
R378 VPB.n84 VPB.n83 7.5
R379 VPB.n97 VPB.n96 7.5
R380 VPB.n91 VPB.n90 7.5
R381 VPB.n93 VPB.n92 7.5
R382 VPB.n86 VPB.n85 7.5
R383 VPB.n102 VPB.n101 7.5
R384 VPB.n373 VPB.n372 7.5
R385 VPB.n386 VPB.n385 7.5
R386 VPB.n380 VPB.n379 7.5
R387 VPB.n382 VPB.n381 7.5
R388 VPB.n375 VPB.n374 7.5
R389 VPB.n391 VPB.n390 7.5
R390 VPB.n18 VPB.n17 7.5
R391 VPB.n31 VPB.n30 7.5
R392 VPB.n25 VPB.n24 7.5
R393 VPB.n27 VPB.n26 7.5
R394 VPB.n20 VPB.n19 7.5
R395 VPB.n36 VPB.n35 7.5
R396 VPB.n469 VPB.n468 7.5
R397 VPB.n12 VPB.n11 7.5
R398 VPB.n6 VPB.n5 7.5
R399 VPB.n8 VPB.n7 7.5
R400 VPB.n2 VPB.n1 7.5
R401 VPB.n471 VPB.n470 7.5
R402 VPB.n37 VPB.n36 7.176
R403 VPB.n392 VPB.n391 7.176
R404 VPB.n329 VPB.n102 7.176
R405 VPB.n126 VPB.n125 7.176
R406 VPB.n252 VPB.n251 7.176
R407 VPB.n247 VPB.n244 6.729
R408 VPB.n243 VPB.n240 6.729
R409 VPB.n238 VPB.n235 6.729
R410 VPB.n121 VPB.n118 6.729
R411 VPB.n117 VPB.n114 6.729
R412 VPB.n112 VPB.n109 6.729
R413 VPB.n98 VPB.n95 6.729
R414 VPB.n94 VPB.n91 6.729
R415 VPB.n89 VPB.n86 6.729
R416 VPB.n387 VPB.n384 6.729
R417 VPB.n383 VPB.n380 6.729
R418 VPB.n378 VPB.n375 6.729
R419 VPB.n32 VPB.n29 6.729
R420 VPB.n28 VPB.n25 6.729
R421 VPB.n23 VPB.n20 6.729
R422 VPB.n13 VPB.n10 6.729
R423 VPB.n9 VPB.n6 6.729
R424 VPB.n4 VPB.n2 6.729
R425 VPB.n238 VPB.n237 6.728
R426 VPB.n243 VPB.n242 6.728
R427 VPB.n247 VPB.n246 6.728
R428 VPB.n250 VPB.n249 6.728
R429 VPB.n112 VPB.n111 6.728
R430 VPB.n117 VPB.n116 6.728
R431 VPB.n121 VPB.n120 6.728
R432 VPB.n124 VPB.n123 6.728
R433 VPB.n89 VPB.n88 6.728
R434 VPB.n94 VPB.n93 6.728
R435 VPB.n98 VPB.n97 6.728
R436 VPB.n101 VPB.n100 6.728
R437 VPB.n378 VPB.n377 6.728
R438 VPB.n383 VPB.n382 6.728
R439 VPB.n387 VPB.n386 6.728
R440 VPB.n390 VPB.n389 6.728
R441 VPB.n23 VPB.n22 6.728
R442 VPB.n28 VPB.n27 6.728
R443 VPB.n32 VPB.n31 6.728
R444 VPB.n35 VPB.n34 6.728
R445 VPB.n4 VPB.n3 6.728
R446 VPB.n9 VPB.n8 6.728
R447 VPB.n13 VPB.n12 6.728
R448 VPB.n472 VPB.n471 6.728
R449 VPB.n200 VPB.n196 6.458
R450 VPB.n350 VPB.n346 6.458
R451 VPB.n190 VPB.n189 6.398
R452 VPB.n209 VPB.n194 6.112
R453 VPB.n209 VPB.n208 6.101
R454 VPB.n294 VPB.n290 4.305
R455 VPB.n159 VPB.n155 4.305
R456 VPB.n434 VPB.n430 4.305
R457 VPB.n70 VPB.n66 4.305
R458 VPB.n277 VPB.n273 3.947
R459 VPB.n146 VPB.n145 3.947
R460 VPB.n417 VPB.n413 3.947
R461 VPB.n57 VPB.n56 3.947
R462 VPB.n225 VPB.n222 1.794
R463 VPB.n365 VPB.n362 1.794
R464 VPB.n208 VPB.n205 1.435
R465 VPB.n338 VPB.n335 1.435
R466 VPB.n188 VPB.n179 1.402
R467 VPB.n188 VPB.n184 1.402
R468 VPB.n188 VPB.n185 1.402
R469 VPB.n188 VPB.n187 1.402
R470 VPB.n265 VPB.n262 1.076
R471 VPB.n137 VPB.n134 1.076
R472 VPB.n405 VPB.n402 1.076
R473 VPB.n48 VPB.n45 1.076
R474 VPB.n189 VPB.n188 0.735
R475 VPB.n188 VPB.n178 0.735
R476 VPB.n304 VPB.n301 0.717
R477 VPB.n167 VPB.n166 0.717
R478 VPB.n444 VPB.n441 0.717
R479 VPB.n78 VPB.n77 0.717
R480 VPB.n248 VPB.n247 0.387
R481 VPB.n248 VPB.n243 0.387
R482 VPB.n248 VPB.n238 0.387
R483 VPB.n249 VPB.n248 0.387
R484 VPB.n122 VPB.n121 0.387
R485 VPB.n122 VPB.n117 0.387
R486 VPB.n122 VPB.n112 0.387
R487 VPB.n123 VPB.n122 0.387
R488 VPB.n99 VPB.n98 0.387
R489 VPB.n99 VPB.n94 0.387
R490 VPB.n99 VPB.n89 0.387
R491 VPB.n100 VPB.n99 0.387
R492 VPB.n388 VPB.n387 0.387
R493 VPB.n388 VPB.n383 0.387
R494 VPB.n388 VPB.n378 0.387
R495 VPB.n389 VPB.n388 0.387
R496 VPB.n33 VPB.n32 0.387
R497 VPB.n33 VPB.n28 0.387
R498 VPB.n33 VPB.n23 0.387
R499 VPB.n34 VPB.n33 0.387
R500 VPB.n473 VPB.n13 0.387
R501 VPB.n473 VPB.n9 0.387
R502 VPB.n473 VPB.n4 0.387
R503 VPB.n473 VPB.n472 0.387
R504 VPB.n257 VPB.n230 0.272
R505 VPB.n314 VPB.n313 0.272
R506 VPB.n397 VPB.n370 0.272
R507 VPB.n454 VPB.n453 0.272
R508 VPB.n465 VPB 0.198
R509 VPB.n211 VPB.n210 0.136
R510 VPB.n216 VPB.n211 0.136
R511 VPB.n221 VPB.n216 0.136
R512 VPB.n226 VPB.n221 0.136
R513 VPB.n230 VPB.n226 0.136
R514 VPB.n261 VPB.n257 0.136
R515 VPB.n266 VPB.n261 0.136
R516 VPB.n271 VPB.n266 0.136
R517 VPB.n278 VPB.n271 0.136
R518 VPB.n283 VPB.n278 0.136
R519 VPB.n288 VPB.n283 0.136
R520 VPB.n295 VPB.n288 0.136
R521 VPB.n300 VPB.n295 0.136
R522 VPB.n305 VPB.n300 0.136
R523 VPB.n309 VPB.n305 0.136
R524 VPB.n313 VPB.n309 0.136
R525 VPB.n315 VPB.n314 0.136
R526 VPB.n316 VPB.n315 0.136
R527 VPB.n317 VPB.n316 0.136
R528 VPB.n318 VPB.n317 0.136
R529 VPB.n319 VPB.n318 0.136
R530 VPB.n320 VPB.n319 0.136
R531 VPB.n321 VPB.n320 0.136
R532 VPB.n322 VPB.n321 0.136
R533 VPB.n323 VPB.n322 0.136
R534 VPB.n324 VPB.n323 0.136
R535 VPB.n325 VPB.n324 0.136
R536 VPB.n325 VPB 0.136
R537 VPB.n334 VPB 0.136
R538 VPB.n339 VPB.n334 0.136
R539 VPB.n344 VPB.n339 0.136
R540 VPB.n351 VPB.n344 0.136
R541 VPB.n356 VPB.n351 0.136
R542 VPB.n361 VPB.n356 0.136
R543 VPB.n366 VPB.n361 0.136
R544 VPB.n370 VPB.n366 0.136
R545 VPB.n401 VPB.n397 0.136
R546 VPB.n406 VPB.n401 0.136
R547 VPB.n411 VPB.n406 0.136
R548 VPB.n418 VPB.n411 0.136
R549 VPB.n423 VPB.n418 0.136
R550 VPB.n428 VPB.n423 0.136
R551 VPB.n435 VPB.n428 0.136
R552 VPB.n440 VPB.n435 0.136
R553 VPB.n445 VPB.n440 0.136
R554 VPB.n449 VPB.n445 0.136
R555 VPB.n453 VPB.n449 0.136
R556 VPB.n455 VPB.n454 0.136
R557 VPB.n456 VPB.n455 0.136
R558 VPB.n457 VPB.n456 0.136
R559 VPB.n458 VPB.n457 0.136
R560 VPB.n459 VPB.n458 0.136
R561 VPB.n460 VPB.n459 0.136
R562 VPB.n461 VPB.n460 0.136
R563 VPB.n462 VPB.n461 0.136
R564 VPB.n463 VPB.n462 0.136
R565 VPB.n464 VPB.n463 0.136
R566 VPB.n465 VPB.n464 0.136
R567 a_599_943.n6 a_599_943.t7 480.392
R568 a_599_943.n8 a_599_943.t11 454.685
R569 a_599_943.n8 a_599_943.t9 428.979
R570 a_599_943.n6 a_599_943.t10 403.272
R571 a_599_943.n7 a_599_943.t8 266.974
R572 a_599_943.n9 a_599_943.t12 221.453
R573 a_599_943.n13 a_599_943.n11 196.598
R574 a_599_943.n11 a_599_943.n5 180.846
R575 a_599_943.n9 a_599_943.n8 108.494
R576 a_599_943.n7 a_599_943.n6 108.494
R577 a_599_943.n10 a_599_943.n9 80.035
R578 a_599_943.n4 a_599_943.n3 79.232
R579 a_599_943.n10 a_599_943.n7 77.315
R580 a_599_943.n11 a_599_943.n10 76
R581 a_599_943.n5 a_599_943.n4 63.152
R582 a_599_943.n13 a_599_943.n12 30
R583 a_599_943.n14 a_599_943.n0 24.383
R584 a_599_943.n14 a_599_943.n13 23.684
R585 a_599_943.n5 a_599_943.n1 16.08
R586 a_599_943.n4 a_599_943.n2 16.08
R587 a_599_943.n1 a_599_943.t1 14.282
R588 a_599_943.n1 a_599_943.t2 14.282
R589 a_599_943.n2 a_599_943.t3 14.282
R590 a_599_943.n2 a_599_943.t4 14.282
R591 a_599_943.n3 a_599_943.t6 14.282
R592 a_599_943.n3 a_599_943.t5 14.282
R593 a_91_75.t0 a_91_75.n0 117.777
R594 a_91_75.n2 a_91_75.n1 55.228
R595 a_91_75.n4 a_91_75.n3 9.111
R596 a_91_75.n8 a_91_75.n6 7.859
R597 a_91_75.t0 a_91_75.n2 4.04
R598 a_91_75.t0 a_91_75.n8 3.034
R599 a_91_75.n6 a_91_75.n4 1.964
R600 a_91_75.n6 a_91_75.n5 1.964
R601 a_91_75.n8 a_91_75.n7 0.443
R602 a_372_182.n10 a_372_182.n8 82.852
R603 a_372_182.n11 a_372_182.n0 49.6
R604 a_372_182.n7 a_372_182.n6 32.833
R605 a_372_182.n8 a_372_182.t1 32.416
R606 a_372_182.n10 a_372_182.n9 27.2
R607 a_372_182.n3 a_372_182.n2 23.284
R608 a_372_182.n11 a_372_182.n10 22.4
R609 a_372_182.n7 a_372_182.n4 19.017
R610 a_372_182.n6 a_372_182.n5 13.494
R611 a_372_182.t1 a_372_182.n1 7.04
R612 a_372_182.t1 a_372_182.n3 5.727
R613 a_372_182.n8 a_372_182.n7 1.435
R614 a_3643_75.t0 a_3643_75.n0 117.777
R615 a_3643_75.n2 a_3643_75.n1 55.228
R616 a_3643_75.n4 a_3643_75.n3 9.111
R617 a_3643_75.n8 a_3643_75.n6 7.859
R618 a_3643_75.t0 a_3643_75.n2 4.04
R619 a_3643_75.t0 a_3643_75.n8 3.034
R620 a_3643_75.n6 a_3643_75.n4 1.964
R621 a_3643_75.n6 a_3643_75.n5 1.964
R622 a_3643_75.n8 a_3643_75.n7 0.443
R623 VNB.n136 VNB.n135 199.897
R624 VNB.n27 VNB.n26 199.897
R625 VNB.n10 VNB.n9 199.897
R626 VNB.n260 VNB.n259 199.897
R627 VNB.n335 VNB.n334 199.897
R628 VNB.n36 VNB.n34 154.509
R629 VNB.n145 VNB.n143 154.509
R630 VNB.n269 VNB.n267 154.509
R631 VNB.n210 VNB.n208 154.509
R632 VNB.n344 VNB.n342 154.509
R633 VNB.n301 VNB.n300 147.75
R634 VNB.n102 VNB.n101 121.366
R635 VNB.n226 VNB.n225 121.366
R636 VNB.n308 VNB.n305 121.366
R637 VNB.n183 VNB.n182 85.559
R638 VNB.n65 VNB.n16 85.559
R639 VNB.n382 VNB.n381 85.559
R640 VNB.n408 VNB.n407 76
R641 VNB.n106 VNB.n105 76
R642 VNB.n117 VNB.n116 76
R643 VNB.n121 VNB.n120 76
R644 VNB.n125 VNB.n124 76
R645 VNB.n147 VNB.n146 76
R646 VNB.n151 VNB.n150 76
R647 VNB.n155 VNB.n154 76
R648 VNB.n159 VNB.n158 76
R649 VNB.n163 VNB.n162 76
R650 VNB.n167 VNB.n166 76
R651 VNB.n171 VNB.n170 76
R652 VNB.n175 VNB.n174 76
R653 VNB.n179 VNB.n178 76
R654 VNB.n185 VNB.n184 76
R655 VNB.n189 VNB.n188 76
R656 VNB.n193 VNB.n192 76
R657 VNB.n206 VNB.n205 76
R658 VNB.n212 VNB.n211 76
R659 VNB.n216 VNB.n215 76
R660 VNB.n220 VNB.n219 76
R661 VNB.n224 VNB.n223 76
R662 VNB.n230 VNB.n229 76
R663 VNB.n241 VNB.n240 76
R664 VNB.n245 VNB.n244 76
R665 VNB.n249 VNB.n248 76
R666 VNB.n271 VNB.n270 76
R667 VNB.n275 VNB.n274 76
R668 VNB.n279 VNB.n278 76
R669 VNB.n283 VNB.n282 76
R670 VNB.n287 VNB.n286 76
R671 VNB.n291 VNB.n290 76
R672 VNB.n295 VNB.n294 76
R673 VNB.n299 VNB.n298 76
R674 VNB.n304 VNB.n303 76
R675 VNB.n316 VNB.n315 76
R676 VNB.n320 VNB.n319 76
R677 VNB.n324 VNB.n323 76
R678 VNB.n346 VNB.n345 76
R679 VNB.n350 VNB.n349 76
R680 VNB.n354 VNB.n353 76
R681 VNB.n358 VNB.n357 76
R682 VNB.n362 VNB.n361 76
R683 VNB.n366 VNB.n365 76
R684 VNB.n370 VNB.n369 76
R685 VNB.n374 VNB.n373 76
R686 VNB.n378 VNB.n377 76
R687 VNB.n384 VNB.n383 76
R688 VNB.n388 VNB.n387 76
R689 VNB.n314 VNB.n313 64.552
R690 VNB.n111 VNB.n110 63.835
R691 VNB.n235 VNB.n234 63.835
R692 VNB.n181 VNB.n180 41.971
R693 VNB.n63 VNB.n62 41.971
R694 VNB.n380 VNB.n379 41.971
R695 VNB.n103 VNB.n102 36.937
R696 VNB.n227 VNB.n226 36.937
R697 VNB.n308 VNB.n307 36.937
R698 VNB.n99 VNB.n98 35.118
R699 VNB.n307 VNB.n306 29.844
R700 VNB.n110 VNB.n109 28.421
R701 VNB.n234 VNB.n233 28.421
R702 VNB.n313 VNB.n312 28.421
R703 VNB.n114 VNB.n113 27.855
R704 VNB.n238 VNB.n237 27.855
R705 VNB.n110 VNB.n108 25.263
R706 VNB.n234 VNB.n232 25.263
R707 VNB.n313 VNB.n311 25.263
R708 VNB.n108 VNB.n107 24.383
R709 VNB.n232 VNB.n231 24.383
R710 VNB.n311 VNB.n310 24.383
R711 VNB.n88 VNB.n85 20.452
R712 VNB.n407 VNB.n404 20.452
R713 VNB.n115 VNB.n114 16.721
R714 VNB.n239 VNB.n238 16.721
R715 VNB.n407 VNB.n406 13.653
R716 VNB.n406 VNB.n405 13.653
R717 VNB.n387 VNB.n386 13.653
R718 VNB.n386 VNB.n385 13.653
R719 VNB.n383 VNB.n380 13.653
R720 VNB.n377 VNB.n376 13.653
R721 VNB.n376 VNB.n375 13.653
R722 VNB.n373 VNB.n372 13.653
R723 VNB.n372 VNB.n371 13.653
R724 VNB.n369 VNB.n368 13.653
R725 VNB.n368 VNB.n367 13.653
R726 VNB.n365 VNB.n364 13.653
R727 VNB.n364 VNB.n363 13.653
R728 VNB.n361 VNB.n360 13.653
R729 VNB.n360 VNB.n359 13.653
R730 VNB.n357 VNB.n356 13.653
R731 VNB.n356 VNB.n355 13.653
R732 VNB.n353 VNB.n352 13.653
R733 VNB.n352 VNB.n351 13.653
R734 VNB.n349 VNB.n348 13.653
R735 VNB.n348 VNB.n347 13.653
R736 VNB.n345 VNB.n344 13.653
R737 VNB.n344 VNB.n343 13.653
R738 VNB.n323 VNB.n322 13.653
R739 VNB.n322 VNB.n321 13.653
R740 VNB.n319 VNB.n318 13.653
R741 VNB.n318 VNB.n317 13.653
R742 VNB.n315 VNB.n309 13.653
R743 VNB.n309 VNB.n308 13.653
R744 VNB.n303 VNB.n302 13.653
R745 VNB.n302 VNB.n301 13.653
R746 VNB.n298 VNB.n297 13.653
R747 VNB.n297 VNB.n296 13.653
R748 VNB.n294 VNB.n293 13.653
R749 VNB.n293 VNB.n292 13.653
R750 VNB.n290 VNB.n289 13.653
R751 VNB.n289 VNB.n288 13.653
R752 VNB.n286 VNB.n285 13.653
R753 VNB.n285 VNB.n284 13.653
R754 VNB.n282 VNB.n281 13.653
R755 VNB.n281 VNB.n280 13.653
R756 VNB.n278 VNB.n277 13.653
R757 VNB.n277 VNB.n276 13.653
R758 VNB.n274 VNB.n273 13.653
R759 VNB.n273 VNB.n272 13.653
R760 VNB.n270 VNB.n269 13.653
R761 VNB.n269 VNB.n268 13.653
R762 VNB.n248 VNB.n247 13.653
R763 VNB.n247 VNB.n246 13.653
R764 VNB.n244 VNB.n243 13.653
R765 VNB.n243 VNB.n242 13.653
R766 VNB.n240 VNB.n239 13.653
R767 VNB.n229 VNB.n228 13.653
R768 VNB.n228 VNB.n227 13.653
R769 VNB.n223 VNB.n222 13.653
R770 VNB.n222 VNB.n221 13.653
R771 VNB.n219 VNB.n218 13.653
R772 VNB.n218 VNB.n217 13.653
R773 VNB.n215 VNB.n214 13.653
R774 VNB.n214 VNB.n213 13.653
R775 VNB.n211 VNB.n210 13.653
R776 VNB.n210 VNB.n209 13.653
R777 VNB.n206 VNB.n70 13.653
R778 VNB.n70 VNB.n69 13.653
R779 VNB.n68 VNB.n67 13.653
R780 VNB.n67 VNB.n66 13.653
R781 VNB.n64 VNB.n63 13.653
R782 VNB.n61 VNB.n60 13.653
R783 VNB.n60 VNB.n59 13.653
R784 VNB.n58 VNB.n57 13.653
R785 VNB.n57 VNB.n56 13.653
R786 VNB.n55 VNB.n54 13.653
R787 VNB.n54 VNB.n53 13.653
R788 VNB.n52 VNB.n51 13.653
R789 VNB.n51 VNB.n50 13.653
R790 VNB.n49 VNB.n48 13.653
R791 VNB.n48 VNB.n47 13.653
R792 VNB.n46 VNB.n45 13.653
R793 VNB.n45 VNB.n44 13.653
R794 VNB.n43 VNB.n42 13.653
R795 VNB.n42 VNB.n41 13.653
R796 VNB.n40 VNB.n39 13.653
R797 VNB.n39 VNB.n38 13.653
R798 VNB.n37 VNB.n36 13.653
R799 VNB.n36 VNB.n35 13.653
R800 VNB.n192 VNB.n191 13.653
R801 VNB.n191 VNB.n190 13.653
R802 VNB.n188 VNB.n187 13.653
R803 VNB.n187 VNB.n186 13.653
R804 VNB.n184 VNB.n181 13.653
R805 VNB.n178 VNB.n177 13.653
R806 VNB.n177 VNB.n176 13.653
R807 VNB.n174 VNB.n173 13.653
R808 VNB.n173 VNB.n172 13.653
R809 VNB.n170 VNB.n169 13.653
R810 VNB.n169 VNB.n168 13.653
R811 VNB.n166 VNB.n165 13.653
R812 VNB.n165 VNB.n164 13.653
R813 VNB.n162 VNB.n161 13.653
R814 VNB.n161 VNB.n160 13.653
R815 VNB.n158 VNB.n157 13.653
R816 VNB.n157 VNB.n156 13.653
R817 VNB.n154 VNB.n153 13.653
R818 VNB.n153 VNB.n152 13.653
R819 VNB.n150 VNB.n149 13.653
R820 VNB.n149 VNB.n148 13.653
R821 VNB.n146 VNB.n145 13.653
R822 VNB.n145 VNB.n144 13.653
R823 VNB.n124 VNB.n123 13.653
R824 VNB.n123 VNB.n122 13.653
R825 VNB.n120 VNB.n119 13.653
R826 VNB.n119 VNB.n118 13.653
R827 VNB.n116 VNB.n115 13.653
R828 VNB.n105 VNB.n104 13.653
R829 VNB.n104 VNB.n103 13.653
R830 VNB.n95 VNB.n94 13.653
R831 VNB.n94 VNB.n93 13.653
R832 VNB.n96 VNB.n92 13.653
R833 VNB.n92 VNB.n91 13.653
R834 VNB.n97 VNB.n90 13.653
R835 VNB.n90 VNB.n89 13.653
R836 VNB.n88 VNB.n87 13.653
R837 VNB.n87 VNB.n86 13.653
R838 VNB.n396 VNB.n393 13.577
R839 VNB.n327 VNB.n325 13.276
R840 VNB.n340 VNB.n327 13.276
R841 VNB.n252 VNB.n250 13.276
R842 VNB.n265 VNB.n252 13.276
R843 VNB.n2 VNB.n0 13.276
R844 VNB.n15 VNB.n2 13.276
R845 VNB.n19 VNB.n17 13.276
R846 VNB.n32 VNB.n19 13.276
R847 VNB.n128 VNB.n126 13.276
R848 VNB.n141 VNB.n128 13.276
R849 VNB.n73 VNB.n71 13.276
R850 VNB.n85 VNB.n73 13.276
R851 VNB.n391 VNB.n389 13.276
R852 VNB.n404 VNB.n391 13.276
R853 VNB.n97 VNB.n96 13.276
R854 VNB.n96 VNB.n95 13.276
R855 VNB.n146 VNB.n142 13.276
R856 VNB.n37 VNB.n33 13.276
R857 VNB.n40 VNB.n37 13.276
R858 VNB.n43 VNB.n40 13.276
R859 VNB.n46 VNB.n43 13.276
R860 VNB.n49 VNB.n46 13.276
R861 VNB.n52 VNB.n49 13.276
R862 VNB.n55 VNB.n52 13.276
R863 VNB.n58 VNB.n55 13.276
R864 VNB.n61 VNB.n58 13.276
R865 VNB.n64 VNB.n61 13.276
R866 VNB.n206 VNB.n68 13.276
R867 VNB.n207 VNB.n206 13.276
R868 VNB.n211 VNB.n207 13.276
R869 VNB.n270 VNB.n266 13.276
R870 VNB.n345 VNB.n341 13.276
R871 VNB.n68 VNB.n65 12.02
R872 VNB.n85 VNB.n84 7.5
R873 VNB.n76 VNB.n75 7.5
R874 VNB.n79 VNB.n78 7.5
R875 VNB.n73 VNB.n72 7.5
R876 VNB.n141 VNB.n140 7.5
R877 VNB.n134 VNB.n133 7.5
R878 VNB.n130 VNB.n129 7.5
R879 VNB.n128 VNB.n127 7.5
R880 VNB.n32 VNB.n31 7.5
R881 VNB.n25 VNB.n24 7.5
R882 VNB.n21 VNB.n20 7.5
R883 VNB.n19 VNB.n18 7.5
R884 VNB.n15 VNB.n14 7.5
R885 VNB.n8 VNB.n7 7.5
R886 VNB.n4 VNB.n3 7.5
R887 VNB.n2 VNB.n1 7.5
R888 VNB.n265 VNB.n264 7.5
R889 VNB.n258 VNB.n257 7.5
R890 VNB.n254 VNB.n253 7.5
R891 VNB.n252 VNB.n251 7.5
R892 VNB.n340 VNB.n339 7.5
R893 VNB.n333 VNB.n332 7.5
R894 VNB.n329 VNB.n328 7.5
R895 VNB.n327 VNB.n326 7.5
R896 VNB.n398 VNB.n397 7.5
R897 VNB.n404 VNB.n403 7.5
R898 VNB.n391 VNB.n390 7.5
R899 VNB.n395 VNB.n394 7.5
R900 VNB.n341 VNB.n340 7.176
R901 VNB.n266 VNB.n265 7.176
R902 VNB.n207 VNB.n15 7.176
R903 VNB.n33 VNB.n32 7.176
R904 VNB.n142 VNB.n141 7.176
R905 VNB.n137 VNB.n134 7.011
R906 VNB.n132 VNB.n130 7.011
R907 VNB.n28 VNB.n25 7.011
R908 VNB.n23 VNB.n21 7.011
R909 VNB.n11 VNB.n8 7.011
R910 VNB.n6 VNB.n4 7.011
R911 VNB.n261 VNB.n258 7.011
R912 VNB.n256 VNB.n254 7.011
R913 VNB.n336 VNB.n333 7.011
R914 VNB.n331 VNB.n329 7.011
R915 VNB.n400 VNB.n398 7.011
R916 VNB.n140 VNB.n139 7.01
R917 VNB.n132 VNB.n131 7.01
R918 VNB.n137 VNB.n136 7.01
R919 VNB.n31 VNB.n30 7.01
R920 VNB.n23 VNB.n22 7.01
R921 VNB.n28 VNB.n27 7.01
R922 VNB.n14 VNB.n13 7.01
R923 VNB.n6 VNB.n5 7.01
R924 VNB.n11 VNB.n10 7.01
R925 VNB.n264 VNB.n263 7.01
R926 VNB.n256 VNB.n255 7.01
R927 VNB.n261 VNB.n260 7.01
R928 VNB.n339 VNB.n338 7.01
R929 VNB.n331 VNB.n330 7.01
R930 VNB.n336 VNB.n335 7.01
R931 VNB.n400 VNB.n399 7.01
R932 VNB.n77 VNB.n74 7.01
R933 VNB.n81 VNB.n79 7.01
R934 VNB.n84 VNB.n83 7.01
R935 VNB.n81 VNB.n80 7.01
R936 VNB.n77 VNB.n76 7.01
R937 VNB.n396 VNB.n395 6.788
R938 VNB.n403 VNB.n402 6.788
R939 VNB.n98 VNB.n88 6.111
R940 VNB.n98 VNB.n97 6.1
R941 VNB.n116 VNB.n111 2.511
R942 VNB.n240 VNB.n235 2.511
R943 VNB.n114 VNB.n112 1.99
R944 VNB.n238 VNB.n236 1.99
R945 VNB.n184 VNB.n183 1.255
R946 VNB.n65 VNB.n64 1.255
R947 VNB.n315 VNB.n314 1.255
R948 VNB.n383 VNB.n382 1.255
R949 VNB.n401 VNB.n392 0.921
R950 VNB.n401 VNB.n396 0.476
R951 VNB.n402 VNB.n401 0.475
R952 VNB.n147 VNB.n125 0.272
R953 VNB.n194 VNB.n193 0.272
R954 VNB.n271 VNB.n249 0.272
R955 VNB.n346 VNB.n324 0.272
R956 VNB.n138 VNB.n132 0.246
R957 VNB.n139 VNB.n138 0.246
R958 VNB.n138 VNB.n137 0.246
R959 VNB.n29 VNB.n23 0.246
R960 VNB.n30 VNB.n29 0.246
R961 VNB.n29 VNB.n28 0.246
R962 VNB.n12 VNB.n6 0.246
R963 VNB.n13 VNB.n12 0.246
R964 VNB.n12 VNB.n11 0.246
R965 VNB.n262 VNB.n256 0.246
R966 VNB.n263 VNB.n262 0.246
R967 VNB.n262 VNB.n261 0.246
R968 VNB.n337 VNB.n331 0.246
R969 VNB.n338 VNB.n337 0.246
R970 VNB.n337 VNB.n336 0.246
R971 VNB.n401 VNB.n400 0.246
R972 VNB.n83 VNB.n82 0.246
R973 VNB.n82 VNB.n81 0.246
R974 VNB.n82 VNB.n77 0.246
R975 VNB.n100 VNB.n99 0.136
R976 VNB.n106 VNB.n100 0.136
R977 VNB.n117 VNB.n106 0.136
R978 VNB.n121 VNB.n117 0.136
R979 VNB.n125 VNB.n121 0.136
R980 VNB.n151 VNB.n147 0.136
R981 VNB.n155 VNB.n151 0.136
R982 VNB.n159 VNB.n155 0.136
R983 VNB.n163 VNB.n159 0.136
R984 VNB.n167 VNB.n163 0.136
R985 VNB.n171 VNB.n167 0.136
R986 VNB.n175 VNB.n171 0.136
R987 VNB.n179 VNB.n175 0.136
R988 VNB.n185 VNB.n179 0.136
R989 VNB.n189 VNB.n185 0.136
R990 VNB.n193 VNB.n189 0.136
R991 VNB.n195 VNB.n194 0.136
R992 VNB.n196 VNB.n195 0.136
R993 VNB.n197 VNB.n196 0.136
R994 VNB.n198 VNB.n197 0.136
R995 VNB.n199 VNB.n198 0.136
R996 VNB.n200 VNB.n199 0.136
R997 VNB.n201 VNB.n200 0.136
R998 VNB.n202 VNB.n201 0.136
R999 VNB.n203 VNB.n202 0.136
R1000 VNB.n204 VNB.n203 0.136
R1001 VNB.n205 VNB.n204 0.136
R1002 VNB.n205 VNB 0.136
R1003 VNB.n212 VNB 0.136
R1004 VNB.n216 VNB.n212 0.136
R1005 VNB.n220 VNB.n216 0.136
R1006 VNB.n224 VNB.n220 0.136
R1007 VNB.n230 VNB.n224 0.136
R1008 VNB.n241 VNB.n230 0.136
R1009 VNB.n245 VNB.n241 0.136
R1010 VNB.n249 VNB.n245 0.136
R1011 VNB.n275 VNB.n271 0.136
R1012 VNB.n279 VNB.n275 0.136
R1013 VNB.n283 VNB.n279 0.136
R1014 VNB.n287 VNB.n283 0.136
R1015 VNB.n291 VNB.n287 0.136
R1016 VNB.n295 VNB.n291 0.136
R1017 VNB.n299 VNB.n295 0.136
R1018 VNB.n304 VNB.n299 0.136
R1019 VNB.n316 VNB.n304 0.136
R1020 VNB.n320 VNB.n316 0.136
R1021 VNB.n324 VNB.n320 0.136
R1022 VNB.n350 VNB.n346 0.136
R1023 VNB.n354 VNB.n350 0.136
R1024 VNB.n358 VNB.n354 0.136
R1025 VNB.n362 VNB.n358 0.136
R1026 VNB.n366 VNB.n362 0.136
R1027 VNB.n370 VNB.n366 0.136
R1028 VNB.n374 VNB.n370 0.136
R1029 VNB.n378 VNB.n374 0.136
R1030 VNB.n384 VNB.n378 0.136
R1031 VNB.n388 VNB.n384 0.136
R1032 VNB.n408 VNB.n388 0.136
R1033 VNB.n408 VNB 0.031
R1034 a_2141_1004.n4 a_2141_1004.t6 512.525
R1035 a_2141_1004.n4 a_2141_1004.t7 371.139
R1036 a_2141_1004.n5 a_2141_1004.t5 271.162
R1037 a_2141_1004.n8 a_2141_1004.n6 194.086
R1038 a_2141_1004.n5 a_2141_1004.n4 172.76
R1039 a_2141_1004.n6 a_2141_1004.n3 162.547
R1040 a_2141_1004.n6 a_2141_1004.n5 153.315
R1041 a_2141_1004.n3 a_2141_1004.n2 76.002
R1042 a_2141_1004.n8 a_2141_1004.n7 30
R1043 a_2141_1004.n9 a_2141_1004.n0 24.383
R1044 a_2141_1004.n9 a_2141_1004.n8 23.684
R1045 a_2141_1004.n1 a_2141_1004.t4 14.282
R1046 a_2141_1004.n1 a_2141_1004.t3 14.282
R1047 a_2141_1004.n2 a_2141_1004.t1 14.282
R1048 a_2141_1004.n2 a_2141_1004.t0 14.282
R1049 a_2141_1004.n3 a_2141_1004.n1 12.85
R1050 a_4626_73.n12 a_4626_73.n11 26.811
R1051 a_4626_73.n6 a_4626_73.n5 24.977
R1052 a_4626_73.n2 a_4626_73.n1 24.877
R1053 a_4626_73.t0 a_4626_73.n2 12.677
R1054 a_4626_73.t0 a_4626_73.n3 11.595
R1055 a_4626_73.t1 a_4626_73.n8 8.137
R1056 a_4626_73.t0 a_4626_73.n4 7.273
R1057 a_4626_73.t0 a_4626_73.n0 6.109
R1058 a_4626_73.t1 a_4626_73.n7 4.864
R1059 a_4626_73.t0 a_4626_73.n12 2.074
R1060 a_4626_73.n7 a_4626_73.n6 1.13
R1061 a_4626_73.n12 a_4626_73.t1 0.937
R1062 a_4626_73.t1 a_4626_73.n10 0.804
R1063 a_4626_73.n10 a_4626_73.n9 0.136
R1064 a_1334_182.n9 a_1334_182.n7 82.852
R1065 a_1334_182.n3 a_1334_182.n1 44.628
R1066 a_1334_182.t0 a_1334_182.n9 32.417
R1067 a_1334_182.n7 a_1334_182.n6 27.2
R1068 a_1334_182.n5 a_1334_182.n4 23.498
R1069 a_1334_182.n3 a_1334_182.n2 23.284
R1070 a_1334_182.n7 a_1334_182.n5 22.4
R1071 a_1334_182.t0 a_1334_182.n11 20.241
R1072 a_1334_182.n11 a_1334_182.n10 13.494
R1073 a_1334_182.t0 a_1334_182.n0 8.137
R1074 a_1334_182.t0 a_1334_182.n3 5.727
R1075 a_1334_182.n9 a_1334_182.n8 1.435
R1076 a_2036_73.n12 a_2036_73.n11 26.811
R1077 a_2036_73.n6 a_2036_73.n5 24.977
R1078 a_2036_73.n2 a_2036_73.n1 24.877
R1079 a_2036_73.t0 a_2036_73.n2 12.677
R1080 a_2036_73.t0 a_2036_73.n3 11.595
R1081 a_2036_73.t1 a_2036_73.n8 8.137
R1082 a_2036_73.t0 a_2036_73.n4 7.273
R1083 a_2036_73.t0 a_2036_73.n0 6.109
R1084 a_2036_73.t1 a_2036_73.n7 4.864
R1085 a_2036_73.t0 a_2036_73.n12 2.074
R1086 a_2036_73.n7 a_2036_73.n6 1.13
R1087 a_2036_73.n12 a_2036_73.t1 0.937
R1088 a_2036_73.t1 a_2036_73.n10 0.804
R1089 a_2036_73.n10 a_2036_73.n9 0.136
R1090 a_2681_75.n4 a_2681_75.n3 19.724
R1091 a_2681_75.t0 a_2681_75.n5 11.595
R1092 a_2681_75.t0 a_2681_75.n4 9.207
R1093 a_2681_75.n2 a_2681_75.n0 8.543
R1094 a_2681_75.t0 a_2681_75.n2 3.034
R1095 a_2681_75.n2 a_2681_75.n1 0.443
R1096 a_3924_182.n8 a_3924_182.n6 96.467
R1097 a_3924_182.n3 a_3924_182.n1 44.628
R1098 a_3924_182.t0 a_3924_182.n8 32.417
R1099 a_3924_182.n3 a_3924_182.n2 23.284
R1100 a_3924_182.n6 a_3924_182.n5 22.349
R1101 a_3924_182.t0 a_3924_182.n10 20.241
R1102 a_3924_182.n10 a_3924_182.n9 13.494
R1103 a_3924_182.n6 a_3924_182.n4 8.443
R1104 a_3924_182.t0 a_3924_182.n0 8.137
R1105 a_3924_182.t0 a_3924_182.n3 5.727
R1106 a_3924_182.n8 a_3924_182.n7 1.435
R1107 a_1053_75.n1 a_1053_75.n0 25.576
R1108 a_1053_75.n3 a_1053_75.n2 9.111
R1109 a_1053_75.n7 a_1053_75.n6 2.455
R1110 a_1053_75.n5 a_1053_75.n3 1.964
R1111 a_1053_75.n5 a_1053_75.n4 1.964
R1112 a_1053_75.t0 a_1053_75.n1 1.871
R1113 a_1053_75.n7 a_1053_75.n5 0.636
R1114 a_1053_75.t0 a_1053_75.n7 0.246
R1115 a_2962_182.n10 a_2962_182.n8 82.852
R1116 a_2962_182.n11 a_2962_182.n0 49.6
R1117 a_2962_182.n7 a_2962_182.n6 32.833
R1118 a_2962_182.n8 a_2962_182.t1 32.416
R1119 a_2962_182.n10 a_2962_182.n9 27.2
R1120 a_2962_182.n3 a_2962_182.n2 23.284
R1121 a_2962_182.n11 a_2962_182.n10 22.4
R1122 a_2962_182.n7 a_2962_182.n4 19.017
R1123 a_2962_182.n6 a_2962_182.n5 13.494
R1124 a_2962_182.t1 a_2962_182.n1 7.04
R1125 a_2962_182.t1 a_2962_182.n3 5.727
R1126 a_2962_182.n8 a_2962_182.n7 1.435



































































































































































































































































































































































































































































































































































































































.ends
