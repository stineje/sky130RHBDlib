// File: dffx1_pcell.spi.pex
// Created: Tue Oct 15 15:56:33 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_DFFX1_PCELL\%noxref_1 ( 37 41 44 49 59 67 75 81 87 95 103 111 119 \
 130 134 136 139 141 143 146 147 148 149 150 151 )
c257 ( 151 0 ) capacitor c=0.0208202f //x=19.12 //y=0.865
c258 ( 150 0 ) capacitor c=0.0208124f //x=15.79 //y=0.865
c259 ( 149 0 ) capacitor c=0.0208017f //x=12.46 //y=0.865
c260 ( 148 0 ) capacitor c=0.0208017f //x=9.13 //y=0.865
c261 ( 147 0 ) capacitor c=0.0208019f //x=5.8 //y=0.865
c262 ( 146 0 ) capacitor c=0.022675f //x=0.885 //y=0.875
c263 ( 145 0 ) capacitor c=0.00440095f //x=19.24 //y=0
c264 ( 143 0 ) capacitor c=0.108011f //x=18.13 //y=0
c265 ( 142 0 ) capacitor c=0.00440095f //x=15.98 //y=0
c266 ( 141 0 ) capacitor c=0.107594f //x=14.8 //y=0
c267 ( 140 0 ) capacitor c=0.00440095f //x=12.65 //y=0
c268 ( 139 0 ) capacitor c=0.107063f //x=11.47 //y=0
c269 ( 138 0 ) capacitor c=0.00440095f //x=9.25 //y=0
c270 ( 136 0 ) capacitor c=0.107063f //x=8.14 //y=0
c271 ( 135 0 ) capacitor c=0.00440095f //x=5.99 //y=0
c272 ( 134 0 ) capacitor c=0.109996f //x=4.81 //y=0
c273 ( 133 0 ) capacitor c=0.00440144f //x=1.075 //y=0
c274 ( 130 0 ) capacitor c=0.25934f //x=21.09 //y=0
c275 ( 119 0 ) capacitor c=0.0426751f //x=19.225 //y=0
c276 ( 111 0 ) capacitor c=0.0751168f //x=17.96 //y=0
c277 ( 103 0 ) capacitor c=0.0426751f //x=15.895 //y=0
c278 ( 95 0 ) capacitor c=0.0751168f //x=14.63 //y=0
c279 ( 87 0 ) capacitor c=0.0389288f //x=12.565 //y=0
c280 ( 81 0 ) capacitor c=0.0720403f //x=11.3 //y=0
c281 ( 75 0 ) capacitor c=0.0389288f //x=9.235 //y=0
c282 ( 67 0 ) capacitor c=0.0720423f //x=7.97 //y=0
c283 ( 59 0 ) capacitor c=0.0389288f //x=5.905 //y=0
c284 ( 49 0 ) capacitor c=0.131745f //x=4.64 //y=0
c285 ( 44 0 ) capacitor c=0.178285f //x=0.74 //y=0
c286 ( 41 0 ) capacitor c=0.0367385f //x=0.99 //y=0
c287 ( 37 0 ) capacitor c=0.713f //x=21.09 //y=0
r288 (  128 130 ) resistor r=26.5322 //w=0.357 //l=0.74 //layer=li \
 //thickness=0.1 //x=20.35 //y=0 //x2=21.09 //y2=0
r289 (  126 145 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.395 //y=0 //x2=19.31 //y2=0
r290 (  126 128 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=19.395 //y=0 //x2=20.35 //y2=0
r291 (  121 145 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.31 //y=0.17 //x2=19.31 //y2=0
r292 (  121 151 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=19.31 //y=0.17 //x2=19.31 //y2=0.955
r293 (  120 143 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.3 //y=0 //x2=18.13 //y2=0
r294 (  119 145 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.225 //y=0 //x2=19.31 //y2=0
r295 (  119 120 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=19.225 //y=0 //x2=18.3 //y2=0
r296 (  114 116 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=16.65 //y=0 //x2=17.76 //y2=0
r297 (  112 142 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.065 //y=0 //x2=15.98 //y2=0
r298 (  112 114 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=16.065 //y=0 //x2=16.65 //y2=0
r299 (  111 143 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.96 //y=0 //x2=18.13 //y2=0
r300 (  111 116 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=17.96 //y=0 //x2=17.76 //y2=0
r301 (  107 142 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.98 //y=0.17 //x2=15.98 //y2=0
r302 (  107 150 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=15.98 //y=0.17 //x2=15.98 //y2=0.955
r303 (  104 141 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.97 //y=0 //x2=14.8 //y2=0
r304 (  104 106 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.97 //y=0 //x2=15.54 //y2=0
r305 (  103 142 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.895 //y=0 //x2=15.98 //y2=0
r306 (  103 106 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=15.895 //y=0 //x2=15.54 //y2=0
r307 (  98 100 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=12.95 //y=0 //x2=14.06 //y2=0
r308 (  96 140 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.735 //y=0 //x2=12.65 //y2=0
r309 (  96 98 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=12.735 //y=0 //x2=12.95 //y2=0
r310 (  95 141 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.63 //y=0 //x2=14.8 //y2=0
r311 (  95 100 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.63 //y=0 //x2=14.06 //y2=0
r312 (  91 140 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.65 //y=0.17 //x2=12.65 //y2=0
r313 (  91 149 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=12.65 //y=0.17 //x2=12.65 //y2=0.955
r314 (  88 139 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.64 //y=0 //x2=11.47 //y2=0
r315 (  88 90 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=11.64 //y=0 //x2=11.84 //y2=0
r316 (  87 140 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.565 //y=0 //x2=12.65 //y2=0
r317 (  87 90 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=12.565 //y=0 //x2=11.84 //y2=0
r318 (  82 138 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.405 //y=0 //x2=9.32 //y2=0
r319 (  82 84 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=9.405 //y=0 //x2=10.36 //y2=0
r320 (  81 139 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.3 //y=0 //x2=11.47 //y2=0
r321 (  81 84 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=11.3 //y=0 //x2=10.36 //y2=0
r322 (  77 138 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.32 //y=0.17 //x2=9.32 //y2=0
r323 (  77 148 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=9.32 //y=0.17 //x2=9.32 //y2=0.955
r324 (  76 136 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=0 //x2=8.14 //y2=0
r325 (  75 138 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.235 //y=0 //x2=9.32 //y2=0
r326 (  75 76 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=9.235 //y=0 //x2=8.31 //y2=0
r327 (  70 72 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r328 (  68 135 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.075 //y=0 //x2=5.99 //y2=0
r329 (  68 70 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=6.075 //y=0 //x2=6.66 //y2=0
r330 (  67 136 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=8.14 //y2=0
r331 (  67 72 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=7.77 //y2=0
r332 (  63 135 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.99 //y=0.17 //x2=5.99 //y2=0
r333 (  63 147 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=5.99 //y=0.17 //x2=5.99 //y2=0.955
r334 (  60 134 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=4.81 //y2=0
r335 (  60 62 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=5.55 //y2=0
r336 (  59 135 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.905 //y=0 //x2=5.99 //y2=0
r337 (  59 62 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=5.905 //y=0 //x2=5.55 //y2=0
r338 (  54 56 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=0 //x2=4.07 //y2=0
r339 (  52 54 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r340 (  50 133 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.075 //y2=0
r341 (  50 52 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.85 //y2=0
r342 (  49 134 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.81 //y2=0
r343 (  49 56 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.07 //y2=0
r344 (  45 133 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0
r345 (  45 146 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0.965
r346 (  41 133 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=1.075 //y2=0
r347 (  41 44 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=0.74 //y2=0
r348 (  37 130 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.09 //y=0 //x2=21.09 //y2=0
r349 (  35 128 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=0 //x2=20.35 //y2=0
r350 (  35 37 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=0 //x2=21.09 //y2=0
r351 (  33 145 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.24 //y=0 //x2=19.24 //y2=0
r352 (  33 35 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.24 //y=0 //x2=20.35 //y2=0
r353 (  31 116 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=0 //x2=17.76 //y2=0
r354 (  31 33 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=0 //x2=19.24 //y2=0
r355 (  29 114 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=0 //x2=16.65 //y2=0
r356 (  29 31 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=0 //x2=17.76 //y2=0
r357 (  27 106 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.54 //y=0 //x2=15.54 //y2=0
r358 (  27 29 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.54 //y=0 //x2=16.65 //y2=0
r359 (  25 100 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=0 //x2=14.06 //y2=0
r360 (  25 27 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=0 //x2=15.54 //y2=0
r361 (  23 98 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.95 //y=0 //x2=12.95 //y2=0
r362 (  23 25 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.95 //y=0 //x2=14.06 //y2=0
r363 (  21 90 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.84 //y=0 //x2=11.84 //y2=0
r364 (  21 23 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.84 //y=0 //x2=12.95 //y2=0
r365 (  19 84 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r366 (  19 21 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=0 //x2=11.84 //y2=0
r367 (  17 138 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=0 //x2=9.25 //y2=0
r368 (  17 19 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=0 //x2=10.36 //y2=0
r369 (  15 72 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r370 (  15 17 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=9.25 //y2=0
r371 (  13 70 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r372 (  13 15 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r373 (  11 62 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r374 (  11 13 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r375 (  9 56 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r376 (  9 11 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=0 //x2=5.55 //y2=0
r377 (  7 54 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r378 (  7 9 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.07 //y2=0
r379 (  5 52 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r380 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r381 (  2 44 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r382 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
ends PM_DFFX1_PCELL\%noxref_1

subckt PM_DFFX1_PCELL\%noxref_2 ( 37 44 51 61 69 79 85 93 101 111 117 125 135 \
 145 149 159 169 177 181 189 197 207 213 221 231 244 251 256 260 265 270 274 \
 275 276 277 278 279 280 281 282 283 284 285 286 287 288 289 290 291 292 )
c289 ( 292 0 ) capacitor c=0.0383753f //x=20.535 //y=5.02
c290 ( 291 0 ) capacitor c=0.0240874f //x=19.655 //y=5.02
c291 ( 290 0 ) capacitor c=0.0493657f //x=18.785 //y=5.02
c292 ( 289 0 ) capacitor c=0.0381505f //x=17.205 //y=5.02
c293 ( 288 0 ) capacitor c=0.0240879f //x=16.325 //y=5.02
c294 ( 287 0 ) capacitor c=0.0493657f //x=15.455 //y=5.02
c295 ( 286 0 ) capacitor c=0.038145f //x=13.875 //y=5.02
c296 ( 285 0 ) capacitor c=0.0240074f //x=12.995 //y=5.02
c297 ( 284 0 ) capacitor c=0.0490303f //x=12.125 //y=5.02
c298 ( 283 0 ) capacitor c=0.0380679f //x=10.545 //y=5.02
c299 ( 282 0 ) capacitor c=0.024008f //x=9.665 //y=5.02
c300 ( 281 0 ) capacitor c=0.0490303f //x=8.795 //y=5.02
c301 ( 280 0 ) capacitor c=0.0380679f //x=7.215 //y=5.02
c302 ( 279 0 ) capacitor c=0.024008f //x=6.335 //y=5.02
c303 ( 278 0 ) capacitor c=0.049209f //x=5.465 //y=5.02
c304 ( 277 0 ) capacitor c=0.0452179f //x=3.585 //y=5.02
c305 ( 276 0 ) capacitor c=0.024152f //x=2.705 //y=5.02
c306 ( 275 0 ) capacitor c=0.02424f //x=1.825 //y=5.02
c307 ( 274 0 ) capacitor c=0.0531407f //x=0.955 //y=5.02
c308 ( 273 0 ) capacitor c=0.00591168f //x=20.68 //y=7.4
c309 ( 272 0 ) capacitor c=0.00591168f //x=19.8 //y=7.4
c310 ( 271 0 ) capacitor c=0.00591168f //x=18.92 //y=7.4
c311 ( 270 0 ) capacitor c=0.116788f //x=18.13 //y=7.4
c312 ( 269 0 ) capacitor c=0.00591168f //x=17.35 //y=7.4
c313 ( 268 0 ) capacitor c=0.00591168f //x=16.47 //y=7.4
c314 ( 267 0 ) capacitor c=0.00591168f //x=15.54 //y=7.4
c315 ( 265 0 ) capacitor c=0.116163f //x=14.8 //y=7.4
c316 ( 264 0 ) capacitor c=0.00591168f //x=14.06 //y=7.4
c317 ( 262 0 ) capacitor c=0.00591168f //x=13.14 //y=7.4
c318 ( 261 0 ) capacitor c=0.00591168f //x=12.26 //y=7.4
c319 ( 260 0 ) capacitor c=0.114361f //x=11.47 //y=7.4
c320 ( 259 0 ) capacitor c=0.00591168f //x=10.69 //y=7.4
c321 ( 258 0 ) capacitor c=0.00591168f //x=9.81 //y=7.4
c322 ( 257 0 ) capacitor c=0.00591168f //x=8.93 //y=7.4
c323 ( 256 0 ) capacitor c=0.11449f //x=8.14 //y=7.4
c324 ( 255 0 ) capacitor c=0.00591168f //x=7.36 //y=7.4
c325 ( 254 0 ) capacitor c=0.00591168f //x=6.48 //y=7.4
c326 ( 253 0 ) capacitor c=0.00591168f //x=5.55 //y=7.4
c327 ( 251 0 ) capacitor c=0.13457f //x=4.81 //y=7.4
c328 ( 250 0 ) capacitor c=0.00591168f //x=3.73 //y=7.4
c329 ( 249 0 ) capacitor c=0.00591168f //x=2.85 //y=7.4
c330 ( 248 0 ) capacitor c=0.00591168f //x=1.97 //y=7.4
c331 ( 247 0 ) capacitor c=0.00591168f //x=1.09 //y=7.4
c332 ( 244 0 ) capacitor c=0.237727f //x=21.09 //y=7.4
c333 ( 231 0 ) capacitor c=0.0284327f //x=20.595 //y=7.4
c334 ( 221 0 ) capacitor c=0.0288633f //x=19.715 //y=7.4
c335 ( 213 0 ) capacitor c=0.0240981f //x=18.835 //y=7.4
c336 ( 207 0 ) capacitor c=0.0236224f //x=17.96 //y=7.4
c337 ( 197 0 ) capacitor c=0.0288639f //x=17.265 //y=7.4
c338 ( 189 0 ) capacitor c=0.0288633f //x=16.385 //y=7.4
c339 ( 181 0 ) capacitor c=0.0240981f //x=15.505 //y=7.4
c340 ( 177 0 ) capacitor c=0.0236947f //x=14.63 //y=7.4
c341 ( 169 0 ) capacitor c=0.0288598f //x=13.935 //y=7.4
c342 ( 159 0 ) capacitor c=0.0288369f //x=13.055 //y=7.4
c343 ( 149 0 ) capacitor c=0.0240981f //x=12.175 //y=7.4
c344 ( 145 0 ) capacitor c=0.0236224f //x=11.3 //y=7.4
c345 ( 135 0 ) capacitor c=0.0288359f //x=10.605 //y=7.4
c346 ( 125 0 ) capacitor c=0.0288369f //x=9.725 //y=7.4
c347 ( 117 0 ) capacitor c=0.0240981f //x=8.845 //y=7.4
c348 ( 111 0 ) capacitor c=0.0236224f //x=7.97 //y=7.4
c349 ( 101 0 ) capacitor c=0.0288359f //x=7.275 //y=7.4
c350 ( 93 0 ) capacitor c=0.0288369f //x=6.395 //y=7.4
c351 ( 85 0 ) capacitor c=0.0240981f //x=5.515 //y=7.4
c352 ( 79 0 ) capacitor c=0.0394667f //x=4.64 //y=7.4
c353 ( 69 0 ) capacitor c=0.0288488f //x=3.645 //y=7.4
c354 ( 61 0 ) capacitor c=0.0287505f //x=2.765 //y=7.4
c355 ( 51 0 ) capacitor c=0.028511f //x=1.885 //y=7.4
c356 ( 44 0 ) capacitor c=0.234426f //x=0.74 //y=7.4
c357 ( 41 0 ) capacitor c=0.0452081f //x=1.005 //y=7.4
c358 ( 37 0 ) capacitor c=0.747675f //x=21.09 //y=7.4
r359 (  242 273 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.765 //y=7.4 //x2=20.68 //y2=7.4
r360 (  242 244 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=20.765 //y=7.4 //x2=21.09 //y2=7.4
r361 (  235 273 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.68 //y=7.23 //x2=20.68 //y2=7.4
r362 (  235 292 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.68 //y=7.23 //x2=20.68 //y2=6.745
r363 (  232 272 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.885 //y=7.4 //x2=19.8 //y2=7.4
r364 (  232 234 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=19.885 //y=7.4 //x2=20.35 //y2=7.4
r365 (  231 273 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.595 //y=7.4 //x2=20.68 //y2=7.4
r366 (  231 234 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=20.595 //y=7.4 //x2=20.35 //y2=7.4
r367 (  225 272 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.8 //y=7.23 //x2=19.8 //y2=7.4
r368 (  225 291 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=19.8 //y=7.23 //x2=19.8 //y2=6.745
r369 (  222 271 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.005 //y=7.4 //x2=18.92 //y2=7.4
r370 (  222 224 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=19.005 //y=7.4 //x2=19.24 //y2=7.4
r371 (  221 272 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.715 //y=7.4 //x2=19.8 //y2=7.4
r372 (  221 224 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=19.715 //y=7.4 //x2=19.24 //y2=7.4
r373 (  215 271 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.92 //y=7.23 //x2=18.92 //y2=7.4
r374 (  215 290 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=18.92 //y=7.23 //x2=18.92 //y2=6.405
r375 (  214 270 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.3 //y=7.4 //x2=18.13 //y2=7.4
r376 (  213 271 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.835 //y=7.4 //x2=18.92 //y2=7.4
r377 (  213 214 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=18.835 //y=7.4 //x2=18.3 //y2=7.4
r378 (  208 269 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.435 //y=7.4 //x2=17.35 //y2=7.4
r379 (  208 210 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=17.435 //y=7.4 //x2=17.76 //y2=7.4
r380 (  207 270 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.96 //y=7.4 //x2=18.13 //y2=7.4
r381 (  207 210 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=17.96 //y=7.4 //x2=17.76 //y2=7.4
r382 (  201 269 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.35 //y=7.23 //x2=17.35 //y2=7.4
r383 (  201 289 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.35 //y=7.23 //x2=17.35 //y2=6.745
r384 (  198 268 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.555 //y=7.4 //x2=16.47 //y2=7.4
r385 (  198 200 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=16.555 //y=7.4 //x2=16.65 //y2=7.4
r386 (  197 269 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.265 //y=7.4 //x2=17.35 //y2=7.4
r387 (  197 200 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=17.265 //y=7.4 //x2=16.65 //y2=7.4
r388 (  191 268 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.47 //y=7.23 //x2=16.47 //y2=7.4
r389 (  191 288 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.47 //y=7.23 //x2=16.47 //y2=6.745
r390 (  190 267 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.675 //y=7.4 //x2=15.59 //y2=7.4
r391 (  189 268 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.385 //y=7.4 //x2=16.47 //y2=7.4
r392 (  189 190 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=16.385 //y=7.4 //x2=15.675 //y2=7.4
r393 (  183 267 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.59 //y=7.23 //x2=15.59 //y2=7.4
r394 (  183 287 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=15.59 //y=7.23 //x2=15.59 //y2=6.405
r395 (  182 265 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.97 //y=7.4 //x2=14.8 //y2=7.4
r396 (  181 267 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.505 //y=7.4 //x2=15.59 //y2=7.4
r397 (  181 182 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=15.505 //y=7.4 //x2=14.97 //y2=7.4
r398 (  178 264 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.105 //y=7.4 //x2=14.02 //y2=7.4
r399 (  177 265 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.63 //y=7.4 //x2=14.8 //y2=7.4
r400 (  177 178 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=14.63 //y=7.4 //x2=14.105 //y2=7.4
r401 (  171 264 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.02 //y=7.23 //x2=14.02 //y2=7.4
r402 (  171 286 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.02 //y=7.23 //x2=14.02 //y2=6.745
r403 (  170 262 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.225 //y=7.4 //x2=13.14 //y2=7.4
r404 (  169 264 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.935 //y=7.4 //x2=14.02 //y2=7.4
r405 (  169 170 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=13.935 //y=7.4 //x2=13.225 //y2=7.4
r406 (  163 262 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.14 //y=7.23 //x2=13.14 //y2=7.4
r407 (  163 285 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=13.14 //y=7.23 //x2=13.14 //y2=6.745
r408 (  160 261 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.345 //y=7.4 //x2=12.26 //y2=7.4
r409 (  160 162 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=12.345 //y=7.4 //x2=12.95 //y2=7.4
r410 (  159 262 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.055 //y=7.4 //x2=13.14 //y2=7.4
r411 (  159 162 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=13.055 //y=7.4 //x2=12.95 //y2=7.4
r412 (  153 261 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.26 //y=7.23 //x2=12.26 //y2=7.4
r413 (  153 284 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=12.26 //y=7.23 //x2=12.26 //y2=6.405
r414 (  150 260 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.64 //y=7.4 //x2=11.47 //y2=7.4
r415 (  150 152 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=11.64 //y=7.4 //x2=11.84 //y2=7.4
r416 (  149 261 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.175 //y=7.4 //x2=12.26 //y2=7.4
r417 (  149 152 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=12.175 //y=7.4 //x2=11.84 //y2=7.4
r418 (  146 259 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.775 //y=7.4 //x2=10.69 //y2=7.4
r419 (  145 260 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.3 //y=7.4 //x2=11.47 //y2=7.4
r420 (  145 146 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=11.3 //y=7.4 //x2=10.775 //y2=7.4
r421 (  139 259 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.69 //y=7.23 //x2=10.69 //y2=7.4
r422 (  139 283 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.69 //y=7.23 //x2=10.69 //y2=6.745
r423 (  136 258 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.895 //y=7.4 //x2=9.81 //y2=7.4
r424 (  136 138 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=9.895 //y=7.4 //x2=10.36 //y2=7.4
r425 (  135 259 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.605 //y=7.4 //x2=10.69 //y2=7.4
r426 (  135 138 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=10.605 //y=7.4 //x2=10.36 //y2=7.4
r427 (  129 258 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.81 //y=7.23 //x2=9.81 //y2=7.4
r428 (  129 282 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=9.81 //y=7.23 //x2=9.81 //y2=6.745
r429 (  126 257 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.015 //y=7.4 //x2=8.93 //y2=7.4
r430 (  126 128 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=9.015 //y=7.4 //x2=9.25 //y2=7.4
r431 (  125 258 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.725 //y=7.4 //x2=9.81 //y2=7.4
r432 (  125 128 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=9.725 //y=7.4 //x2=9.25 //y2=7.4
r433 (  119 257 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.93 //y=7.23 //x2=8.93 //y2=7.4
r434 (  119 281 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=8.93 //y=7.23 //x2=8.93 //y2=6.405
r435 (  118 256 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=7.4 //x2=8.14 //y2=7.4
r436 (  117 257 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.845 //y=7.4 //x2=8.93 //y2=7.4
r437 (  117 118 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=8.845 //y=7.4 //x2=8.31 //y2=7.4
r438 (  112 255 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.445 //y=7.4 //x2=7.36 //y2=7.4
r439 (  112 114 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=7.445 //y=7.4 //x2=7.77 //y2=7.4
r440 (  111 256 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=8.14 //y2=7.4
r441 (  111 114 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=7.77 //y2=7.4
r442 (  105 255 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.36 //y=7.23 //x2=7.36 //y2=7.4
r443 (  105 280 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.36 //y=7.23 //x2=7.36 //y2=6.745
r444 (  102 254 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.565 //y=7.4 //x2=6.48 //y2=7.4
r445 (  102 104 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=6.565 //y=7.4 //x2=6.66 //y2=7.4
r446 (  101 255 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.275 //y=7.4 //x2=7.36 //y2=7.4
r447 (  101 104 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=7.275 //y=7.4 //x2=6.66 //y2=7.4
r448 (  95 254 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.48 //y=7.23 //x2=6.48 //y2=7.4
r449 (  95 279 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.48 //y=7.23 //x2=6.48 //y2=6.745
r450 (  94 253 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.685 //y=7.4 //x2=5.6 //y2=7.4
r451 (  93 254 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.395 //y=7.4 //x2=6.48 //y2=7.4
r452 (  93 94 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=6.395 //y=7.4 //x2=5.685 //y2=7.4
r453 (  87 253 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.6 //y=7.23 //x2=5.6 //y2=7.4
r454 (  87 278 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=5.6 //y=7.23 //x2=5.6 //y2=6.405
r455 (  86 251 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=4.81 //y2=7.4
r456 (  85 253 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.515 //y=7.4 //x2=5.6 //y2=7.4
r457 (  85 86 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=5.515 //y=7.4 //x2=4.98 //y2=7.4
r458 (  80 250 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=3.73 //y2=7.4
r459 (  80 82 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=4.07 //y2=7.4
r460 (  79 251 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.81 //y2=7.4
r461 (  79 82 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.07 //y2=7.4
r462 (  73 250 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=7.4
r463 (  73 277 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=6.745
r464 (  70 249 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.85 //y2=7.4
r465 (  70 72 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.96 //y2=7.4
r466 (  69 250 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=3.73 //y2=7.4
r467 (  69 72 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=2.96 //y2=7.4
r468 (  63 249 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=7.4
r469 (  63 276 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=6.745
r470 (  62 248 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.055 //y=7.4 //x2=1.97 //y2=7.4
r471 (  61 249 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.85 //y2=7.4
r472 (  61 62 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.055 //y2=7.4
r473 (  55 248 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=7.4
r474 (  55 275 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=6.745
r475 (  52 247 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.09 //y2=7.4
r476 (  52 54 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.85 //y2=7.4
r477 (  51 248 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.97 //y2=7.4
r478 (  51 54 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.85 //y2=7.4
r479 (  45 247 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=7.4
r480 (  45 274 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=6.405
r481 (  41 247 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=1.09 //y2=7.4
r482 (  41 44 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=0.74 //y2=7.4
r483 (  37 244 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.09 //y=7.4 //x2=21.09 //y2=7.4
r484 (  35 234 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=7.4 //x2=20.35 //y2=7.4
r485 (  35 37 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=7.4 //x2=21.09 //y2=7.4
r486 (  33 224 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.24 //y=7.4 //x2=19.24 //y2=7.4
r487 (  33 35 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.24 //y=7.4 //x2=20.35 //y2=7.4
r488 (  31 210 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=7.4 //x2=17.76 //y2=7.4
r489 (  31 33 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=7.4 //x2=19.24 //y2=7.4
r490 (  29 200 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=7.4 //x2=16.65 //y2=7.4
r491 (  29 31 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=7.4 //x2=17.76 //y2=7.4
r492 (  27 267 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.54 //y=7.4 //x2=15.54 //y2=7.4
r493 (  27 29 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.54 //y=7.4 //x2=16.65 //y2=7.4
r494 (  25 264 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=7.4 //x2=14.06 //y2=7.4
r495 (  25 27 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=7.4 //x2=15.54 //y2=7.4
r496 (  23 162 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.95 //y=7.4 //x2=12.95 //y2=7.4
r497 (  23 25 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.95 //y=7.4 //x2=14.06 //y2=7.4
r498 (  21 152 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.84 //y=7.4 //x2=11.84 //y2=7.4
r499 (  21 23 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.84 //y=7.4 //x2=12.95 //y2=7.4
r500 (  19 138 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r501 (  19 21 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=7.4 //x2=11.84 //y2=7.4
r502 (  17 128 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=7.4 //x2=9.25 //y2=7.4
r503 (  17 19 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=7.4 //x2=10.36 //y2=7.4
r504 (  15 114 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=7.4 //x2=7.77 //y2=7.4
r505 (  15 17 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=7.4 //x2=9.25 //y2=7.4
r506 (  13 104 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r507 (  13 15 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.4 //x2=7.77 //y2=7.4
r508 (  11 253 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r509 (  11 13 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.66 //y2=7.4
r510 (  9 82 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=7.4 //x2=4.07 //y2=7.4
r511 (  9 11 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=7.4 //x2=5.55 //y2=7.4
r512 (  7 72 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r513 (  7 9 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r514 (  5 54 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r515 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r516 (  2 44 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r517 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_DFFX1_PCELL\%noxref_2

subckt PM_DFFX1_PCELL\%noxref_3 ( 1 2 3 4 12 25 26 37 39 40 44 46 53 54 55 56 \
 57 58 59 63 64 65 70 72 75 76 77 78 79 80 84 86 89 90 95 96 101 110 113 115 \
 116 )
c232 ( 116 0 ) capacitor c=0.0220291f //x=6.775 //y=5.02
c233 ( 115 0 ) capacitor c=0.0217503f //x=5.895 //y=5.02
c234 ( 113 0 ) capacitor c=0.00866655f //x=6.77 //y=0.905
c235 ( 110 0 ) capacitor c=0.0588816f //x=9.25 //y=4.7
c236 ( 101 0 ) capacitor c=0.058931f //x=3.33 //y=4.7
c237 ( 96 0 ) capacitor c=0.0273931f //x=3.33 //y=1.915
c238 ( 95 0 ) capacitor c=0.0464411f //x=3.33 //y=2.08
c239 ( 90 0 ) capacitor c=0.0318948f //x=9.585 //y=1.21
c240 ( 89 0 ) capacitor c=0.0187384f //x=9.585 //y=0.865
c241 ( 86 0 ) capacitor c=0.0141798f //x=9.43 //y=1.365
c242 ( 84 0 ) capacitor c=0.0149844f //x=9.43 //y=0.71
c243 ( 80 0 ) capacitor c=0.0853292f //x=9.055 //y=1.915
c244 ( 79 0 ) capacitor c=0.0229722f //x=9.055 //y=1.52
c245 ( 78 0 ) capacitor c=0.0234352f //x=9.055 //y=1.21
c246 ( 77 0 ) capacitor c=0.0199343f //x=9.055 //y=0.865
c247 ( 76 0 ) capacitor c=0.0432517f //x=3.85 //y=1.26
c248 ( 75 0 ) capacitor c=0.0200379f //x=3.85 //y=0.915
c249 ( 72 0 ) capacitor c=0.0158629f //x=3.695 //y=1.415
c250 ( 70 0 ) capacitor c=0.0157803f //x=3.695 //y=0.76
c251 ( 65 0 ) capacitor c=0.0218028f //x=3.32 //y=1.57
c252 ( 64 0 ) capacitor c=0.0207459f //x=3.32 //y=1.26
c253 ( 63 0 ) capacitor c=0.0194308f //x=3.32 //y=0.915
c254 ( 59 0 ) capacitor c=0.110275f //x=9.59 //y=6.02
c255 ( 58 0 ) capacitor c=0.154305f //x=9.15 //y=6.02
c256 ( 57 0 ) capacitor c=0.158794f //x=3.51 //y=6.02
c257 ( 56 0 ) capacitor c=0.110114f //x=3.07 //y=6.02
c258 ( 53 0 ) capacitor c=0.00211606f //x=6.92 //y=5.2
c259 ( 46 0 ) capacitor c=0.0917424f //x=9.25 //y=2.08
c260 ( 44 0 ) capacitor c=0.108359f //x=7.4 //y=3.33
c261 ( 40 0 ) capacitor c=0.00498573f //x=7.045 //y=1.655
c262 ( 39 0 ) capacitor c=0.0136303f //x=7.315 //y=1.655
c263 ( 37 0 ) capacitor c=0.0137522f //x=7.315 //y=5.2
c264 ( 26 0 ) capacitor c=0.00251635f //x=6.125 //y=5.2
c265 ( 25 0 ) capacitor c=0.0142423f //x=6.835 //y=5.2
c266 ( 12 0 ) capacitor c=0.0883349f //x=3.33 //y=2.08
c267 ( 4 0 ) capacitor c=0.0042919f //x=7.515 //y=3.33
c268 ( 3 0 ) capacitor c=0.0617718f //x=9.135 //y=3.33
c269 ( 2 0 ) capacitor c=0.0149802f //x=3.445 //y=3.33
c270 ( 1 0 ) capacitor c=0.108369f //x=7.285 //y=3.33
r271 (  108 110 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=9.15 //y=4.7 //x2=9.25 //y2=4.7
r272 (  95 96 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.33 //y=2.08 //x2=3.33 //y2=1.915
r273 (  91 110 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=9.59 //y=4.865 //x2=9.25 //y2=4.7
r274 (  90 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.585 //y=1.21 //x2=9.545 //y2=1.365
r275 (  89 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.585 //y=0.865 //x2=9.545 //y2=0.71
r276 (  89 90 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.585 //y=0.865 //x2=9.585 //y2=1.21
r277 (  87 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.21 //y=1.365 //x2=9.095 //y2=1.365
r278 (  86 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.43 //y=1.365 //x2=9.545 //y2=1.365
r279 (  85 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.21 //y=0.71 //x2=9.095 //y2=0.71
r280 (  84 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.43 //y=0.71 //x2=9.545 //y2=0.71
r281 (  84 85 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=9.43 //y=0.71 //x2=9.21 //y2=0.71
r282 (  81 108 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=9.15 //y=4.865 //x2=9.15 //y2=4.7
r283 (  80 105 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=9.055 //y=1.915 //x2=9.25 //y2=2.08
r284 (  79 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.055 //y=1.52 //x2=9.095 //y2=1.365
r285 (  79 80 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=9.055 //y=1.52 //x2=9.055 //y2=1.915
r286 (  78 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.055 //y=1.21 //x2=9.095 //y2=1.365
r287 (  77 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.055 //y=0.865 //x2=9.095 //y2=0.71
r288 (  77 78 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.055 //y=0.865 //x2=9.055 //y2=1.21
r289 (  76 103 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=1.26 //x2=3.81 //y2=1.415
r290 (  75 102 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.81 //y2=0.76
r291 (  75 76 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.85 //y2=1.26
r292 (  73 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=1.415 //x2=3.36 //y2=1.415
r293 (  72 103 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=1.415 //x2=3.81 //y2=1.415
r294 (  71 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=0.76 //x2=3.36 //y2=0.76
r295 (  70 102 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.81 //y2=0.76
r296 (  70 71 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.475 //y2=0.76
r297 (  67 101 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=3.51 //y=4.865 //x2=3.33 //y2=4.7
r298 (  65 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.36 //y2=1.415
r299 (  65 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.32 //y2=1.915
r300 (  64 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.26 //x2=3.36 //y2=1.415
r301 (  63 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.36 //y2=0.76
r302 (  63 64 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.32 //y2=1.26
r303 (  60 101 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=3.07 //y=4.865 //x2=3.33 //y2=4.7
r304 (  59 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.59 //y=6.02 //x2=9.59 //y2=4.865
r305 (  58 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.15 //y=6.02 //x2=9.15 //y2=4.865
r306 (  57 67 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.51 //y=6.02 //x2=3.51 //y2=4.865
r307 (  56 60 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.07 //y=6.02 //x2=3.07 //y2=4.865
r308 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.32 //y=1.365 //x2=9.43 //y2=1.365
r309 (  55 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.32 //y=1.365 //x2=9.21 //y2=1.365
r310 (  54 72 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.695 //y2=1.415
r311 (  54 73 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.475 //y2=1.415
r312 (  51 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=4.7 //x2=9.25 //y2=4.7
r313 (  49 51 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=9.25 //y=3.33 //x2=9.25 //y2=4.7
r314 (  46 105 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=2.08 //x2=9.25 //y2=2.08
r315 (  46 49 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=9.25 //y=2.08 //x2=9.25 //y2=3.33
r316 (  42 44 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=7.4 //y=5.115 //x2=7.4 //y2=3.33
r317 (  41 44 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=7.4 //y=1.74 //x2=7.4 //y2=3.33
r318 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.655 //x2=7.4 //y2=1.74
r319 (  39 40 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.655 //x2=7.045 //y2=1.655
r320 (  38 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.005 //y=5.2 //x2=6.92 //y2=5.2
r321 (  37 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.2 //x2=7.4 //y2=5.115
r322 (  37 38 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.2 //x2=7.005 //y2=5.2
r323 (  33 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.96 //y=1.57 //x2=7.045 //y2=1.655
r324 (  33 113 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=6.96 //y=1.57 //x2=6.96 //y2=1
r325 (  27 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.92 //y=5.285 //x2=6.92 //y2=5.2
r326 (  27 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=6.92 //y=5.285 //x2=6.92 //y2=5.725
r327 (  25 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.835 //y=5.2 //x2=6.92 //y2=5.2
r328 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=6.835 //y=5.2 //x2=6.125 //y2=5.2
r329 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.04 //y=5.285 //x2=6.125 //y2=5.2
r330 (  19 115 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=6.04 //y=5.285 //x2=6.04 //y2=5.725
r331 (  17 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r332 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=3.33 //x2=3.33 //y2=4.7
r333 (  12 95 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r334 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.08 //x2=3.33 //y2=3.33
r335 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.25 //y=3.33 //x2=9.25 //y2=3.33
r336 (  8 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=7.4 \
 //y=3.33 //x2=7.4 //y2=3.33
r337 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=3.33 //x2=3.33 //y2=3.33
r338 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.515 //y=3.33 //x2=7.4 //y2=3.33
r339 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.135 //y=3.33 //x2=9.25 //y2=3.33
r340 (  3 4 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=9.135 //y=3.33 //x2=7.515 //y2=3.33
r341 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.445 //y=3.33 //x2=3.33 //y2=3.33
r342 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.285 //y=3.33 //x2=7.4 //y2=3.33
r343 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=7.285 //y=3.33 //x2=3.445 //y2=3.33
ends PM_DFFX1_PCELL\%noxref_3

subckt PM_DFFX1_PCELL\%noxref_4 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 \
 47 48 52 54 57 58 68 71 73 74 )
c150 ( 74 0 ) capacitor c=0.0220291f //x=10.105 //y=5.02
c151 ( 73 0 ) capacitor c=0.0217503f //x=9.225 //y=5.02
c152 ( 71 0 ) capacitor c=0.00866655f //x=10.1 //y=0.905
c153 ( 68 0 ) capacitor c=0.0588816f //x=12.58 //y=4.7
c154 ( 58 0 ) capacitor c=0.0318948f //x=12.915 //y=1.21
c155 ( 57 0 ) capacitor c=0.0187384f //x=12.915 //y=0.865
c156 ( 54 0 ) capacitor c=0.0141798f //x=12.76 //y=1.365
c157 ( 52 0 ) capacitor c=0.0149844f //x=12.76 //y=0.71
c158 ( 48 0 ) capacitor c=0.0853292f //x=12.385 //y=1.915
c159 ( 47 0 ) capacitor c=0.0229722f //x=12.385 //y=1.52
c160 ( 46 0 ) capacitor c=0.0234352f //x=12.385 //y=1.21
c161 ( 45 0 ) capacitor c=0.0199343f //x=12.385 //y=0.865
c162 ( 44 0 ) capacitor c=0.110275f //x=12.92 //y=6.02
c163 ( 43 0 ) capacitor c=0.154305f //x=12.48 //y=6.02
c164 ( 41 0 ) capacitor c=0.00211606f //x=10.25 //y=5.2
c165 ( 34 0 ) capacitor c=0.0911845f //x=12.58 //y=2.08
c166 ( 32 0 ) capacitor c=0.108686f //x=10.73 //y=3.33
c167 ( 28 0 ) capacitor c=0.00525782f //x=10.375 //y=1.655
c168 ( 27 0 ) capacitor c=0.0139525f //x=10.645 //y=1.655
c169 ( 25 0 ) capacitor c=0.0137522f //x=10.645 //y=5.2
c170 ( 14 0 ) capacitor c=0.00251459f //x=9.455 //y=5.2
c171 ( 13 0 ) capacitor c=0.0143649f //x=10.165 //y=5.2
c172 ( 2 0 ) capacitor c=0.00861293f //x=10.845 //y=3.33
c173 ( 1 0 ) capacitor c=0.067133f //x=12.465 //y=3.33
r174 (  66 68 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=12.48 //y=4.7 //x2=12.58 //y2=4.7
r175 (  59 68 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=12.92 //y=4.865 //x2=12.58 //y2=4.7
r176 (  58 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.915 //y=1.21 //x2=12.875 //y2=1.365
r177 (  57 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.915 //y=0.865 //x2=12.875 //y2=0.71
r178 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.915 //y=0.865 //x2=12.915 //y2=1.21
r179 (  55 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.54 //y=1.365 //x2=12.425 //y2=1.365
r180 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.76 //y=1.365 //x2=12.875 //y2=1.365
r181 (  53 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.54 //y=0.71 //x2=12.425 //y2=0.71
r182 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.76 //y=0.71 //x2=12.875 //y2=0.71
r183 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=12.76 //y=0.71 //x2=12.54 //y2=0.71
r184 (  49 66 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=12.48 //y=4.865 //x2=12.48 //y2=4.7
r185 (  48 63 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=12.385 //y=1.915 //x2=12.58 //y2=2.08
r186 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.385 //y=1.52 //x2=12.425 //y2=1.365
r187 (  47 48 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=12.385 //y=1.52 //x2=12.385 //y2=1.915
r188 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.385 //y=1.21 //x2=12.425 //y2=1.365
r189 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.385 //y=0.865 //x2=12.425 //y2=0.71
r190 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.385 //y=0.865 //x2=12.385 //y2=1.21
r191 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.92 //y=6.02 //x2=12.92 //y2=4.865
r192 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.48 //y=6.02 //x2=12.48 //y2=4.865
r193 (  42 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.65 //y=1.365 //x2=12.76 //y2=1.365
r194 (  42 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.65 //y=1.365 //x2=12.54 //y2=1.365
r195 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.58 //y=4.7 //x2=12.58 //y2=4.7
r196 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=12.58 //y=3.33 //x2=12.58 //y2=4.7
r197 (  34 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.58 //y=2.08 //x2=12.58 //y2=2.08
r198 (  34 37 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=12.58 //y=2.08 //x2=12.58 //y2=3.33
r199 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=10.73 //y=5.115 //x2=10.73 //y2=3.33
r200 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=10.73 //y=1.74 //x2=10.73 //y2=3.33
r201 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.645 //y=1.655 //x2=10.73 //y2=1.74
r202 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=10.645 //y=1.655 //x2=10.375 //y2=1.655
r203 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.335 //y=5.2 //x2=10.25 //y2=5.2
r204 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.645 //y=5.2 //x2=10.73 //y2=5.115
r205 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=10.645 //y=5.2 //x2=10.335 //y2=5.2
r206 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.29 //y=1.57 //x2=10.375 //y2=1.655
r207 (  21 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=10.29 //y=1.57 //x2=10.29 //y2=1
r208 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.25 //y=5.285 //x2=10.25 //y2=5.2
r209 (  15 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=10.25 //y=5.285 //x2=10.25 //y2=5.725
r210 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.165 //y=5.2 //x2=10.25 //y2=5.2
r211 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.165 //y=5.2 //x2=9.455 //y2=5.2
r212 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.37 //y=5.285 //x2=9.455 //y2=5.2
r213 (  7 73 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=9.37 //y=5.285 //x2=9.37 //y2=5.725
r214 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.58 //y=3.33 //x2=12.58 //y2=3.33
r215 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.73 //y=3.33 //x2=10.73 //y2=3.33
r216 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.845 //y=3.33 //x2=10.73 //y2=3.33
r217 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.465 //y=3.33 //x2=12.58 //y2=3.33
r218 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=12.465 //y=3.33 //x2=10.845 //y2=3.33
ends PM_DFFX1_PCELL\%noxref_4

subckt PM_DFFX1_PCELL\%noxref_5 ( 1 2 8 15 17 23 24 25 26 27 28 29 30 31 33 39 \
 40 41 42 43 48 49 50 55 57 59 65 66 70 79 80 83 )
c205 ( 83 0 ) capacitor c=0.0331838f //x=13.35 //y=4.7
c206 ( 80 0 ) capacitor c=0.0279499f //x=13.32 //y=1.915
c207 ( 79 0 ) capacitor c=0.0437302f //x=13.32 //y=2.08
c208 ( 70 0 ) capacitor c=0.0334842f //x=2.22 //y=4.7
c209 ( 66 0 ) capacitor c=0.0429696f //x=13.885 //y=1.25
c210 ( 65 0 ) capacitor c=0.0192208f //x=13.885 //y=0.905
c211 ( 59 0 ) capacitor c=0.0158629f //x=13.73 //y=1.405
c212 ( 57 0 ) capacitor c=0.0157803f //x=13.73 //y=0.75
c213 ( 55 0 ) capacitor c=0.0299681f //x=13.725 //y=4.79
c214 ( 50 0 ) capacitor c=0.0205163f //x=13.355 //y=1.56
c215 ( 49 0 ) capacitor c=0.0168481f //x=13.355 //y=1.25
c216 ( 48 0 ) capacitor c=0.0174783f //x=13.355 //y=0.905
c217 ( 43 0 ) capacitor c=0.0245352f //x=2.555 //y=4.79
c218 ( 42 0 ) capacitor c=0.0850619f //x=2.31 //y=1.915
c219 ( 41 0 ) capacitor c=0.0170266f //x=2.31 //y=1.45
c220 ( 40 0 ) capacitor c=0.018609f //x=2.31 //y=1.22
c221 ( 39 0 ) capacitor c=0.0187309f //x=2.31 //y=0.91
c222 ( 33 0 ) capacitor c=0.014725f //x=2.155 //y=1.375
c223 ( 31 0 ) capacitor c=0.0146567f //x=2.155 //y=0.755
c224 ( 30 0 ) capacitor c=0.0335408f //x=1.785 //y=1.22
c225 ( 29 0 ) capacitor c=0.0173761f //x=1.785 //y=0.91
c226 ( 28 0 ) capacitor c=0.15358f //x=13.8 //y=6.02
c227 ( 27 0 ) capacitor c=0.110281f //x=13.36 //y=6.02
c228 ( 26 0 ) capacitor c=0.110114f //x=2.63 //y=6.02
c229 ( 25 0 ) capacitor c=0.11012f //x=2.19 //y=6.02
c230 ( 17 0 ) capacitor c=0.0746615f //x=13.32 //y=2.08
c231 ( 15 0 ) capacitor c=0.00369614f //x=13.32 //y=4.535
c232 ( 8 0 ) capacitor c=0.100158f //x=2.22 //y=2.08
c233 ( 2 0 ) capacitor c=0.0154455f //x=2.335 //y=4.44
c234 ( 1 0 ) capacitor c=0.257146f //x=13.205 //y=4.44
r235 (  85 86 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=13.35 //y=4.79 //x2=13.35 //y2=4.865
r236 (  83 85 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=13.35 //y=4.7 //x2=13.35 //y2=4.79
r237 (  79 80 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=13.32 //y=2.08 //x2=13.32 //y2=1.915
r238 (  72 73 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.79 //x2=2.22 //y2=4.865
r239 (  70 72 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.7 //x2=2.22 //y2=4.79
r240 (  66 90 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.885 //y=1.25 //x2=13.845 //y2=1.405
r241 (  65 89 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.885 //y=0.905 //x2=13.845 //y2=0.75
r242 (  65 66 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.885 //y=0.905 //x2=13.885 //y2=1.25
r243 (  60 88 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.51 //y=1.405 //x2=13.395 //y2=1.405
r244 (  59 90 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.73 //y=1.405 //x2=13.845 //y2=1.405
r245 (  58 87 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.51 //y=0.75 //x2=13.395 //y2=0.75
r246 (  57 89 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.73 //y=0.75 //x2=13.845 //y2=0.75
r247 (  57 58 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=13.73 //y=0.75 //x2=13.51 //y2=0.75
r248 (  56 85 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=13.485 //y=4.79 //x2=13.35 //y2=4.79
r249 (  55 62 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=13.725 //y=4.79 //x2=13.8 //y2=4.865
r250 (  55 56 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=13.725 //y=4.79 //x2=13.485 //y2=4.79
r251 (  50 88 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.355 //y=1.56 //x2=13.395 //y2=1.405
r252 (  50 80 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=13.355 //y=1.56 //x2=13.355 //y2=1.915
r253 (  49 88 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.355 //y=1.25 //x2=13.395 //y2=1.405
r254 (  48 87 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.355 //y=0.905 //x2=13.395 //y2=0.75
r255 (  48 49 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.355 //y=0.905 //x2=13.355 //y2=1.25
r256 (  44 72 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.355 //y=4.79 //x2=2.22 //y2=4.79
r257 (  43 45 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.63 //y2=4.865
r258 (  43 44 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.355 //y2=4.79
r259 (  42 77 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.915 //x2=2.235 //y2=2.08
r260 (  41 75 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.27 //y2=1.375
r261 (  41 42 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.31 //y2=1.915
r262 (  40 75 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.22 //x2=2.27 //y2=1.375
r263 (  39 74 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.27 //y2=0.755
r264 (  39 40 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.31 //y2=1.22
r265 (  34 68 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=1.375 //x2=1.825 //y2=1.375
r266 (  33 75 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=1.375 //x2=2.27 //y2=1.375
r267 (  32 67 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=0.755 //x2=1.825 //y2=0.755
r268 (  31 74 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=2.27 //y2=0.755
r269 (  31 32 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=1.94 //y2=0.755
r270 (  30 68 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=1.22 //x2=1.825 //y2=1.375
r271 (  29 67 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.825 //y2=0.755
r272 (  29 30 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.785 //y2=1.22
r273 (  28 62 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.8 //y=6.02 //x2=13.8 //y2=4.865
r274 (  27 86 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.36 //y=6.02 //x2=13.36 //y2=4.865
r275 (  26 45 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.63 //y=6.02 //x2=2.63 //y2=4.865
r276 (  25 73 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.19 //y=6.02 //x2=2.19 //y2=4.865
r277 (  24 59 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.62 //y=1.405 //x2=13.73 //y2=1.405
r278 (  24 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.62 //y=1.405 //x2=13.51 //y2=1.405
r279 (  23 33 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=2.155 //y2=1.375
r280 (  23 34 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=1.94 //y2=1.375
r281 (  22 83 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=13.35 //y=4.7 //x2=13.35 //y2=4.7
r282 (  17 79 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=13.32 //y=2.08 //x2=13.32 //y2=2.08
r283 (  17 20 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=13.32 //y=2.08 //x2=13.32 //y2=4.44
r284 (  15 22 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=13.32 //y=4.535 //x2=13.335 //y2=4.7
r285 (  15 20 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=13.32 //y=4.535 //x2=13.32 //y2=4.44
r286 (  13 70 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=4.7 //x2=2.22 //y2=4.7
r287 (  11 13 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=2.22 //y=4.44 //x2=2.22 //y2=4.7
r288 (  8 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=2.08
r289 (  8 11 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li //thickness=0.1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=4.44
r290 (  6 20 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=13.32 //y=4.44 //x2=13.32 //y2=4.44
r291 (  4 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.22 //y=4.44 //x2=2.22 //y2=4.44
r292 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.335 //y=4.44 //x2=2.22 //y2=4.44
r293 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.205 //y=4.44 //x2=13.32 //y2=4.44
r294 (  1 2 ) resistor r=10.3721 //w=0.131 //l=10.87 //layer=m1 \
 //thickness=0.36 //x=13.205 //y=4.44 //x2=2.335 //y2=4.44
ends PM_DFFX1_PCELL\%noxref_5

subckt PM_DFFX1_PCELL\%noxref_6 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 63 \
 64 65 66 67 68 69 70 71 72 76 78 81 82 86 87 88 89 93 95 98 99 109 118 121 \
 123 124 125 )
c251 ( 125 0 ) capacitor c=0.023087f //x=3.145 //y=5.02
c252 ( 124 0 ) capacitor c=0.023519f //x=2.265 //y=5.02
c253 ( 123 0 ) capacitor c=0.0224735f //x=1.385 //y=5.02
c254 ( 121 0 ) capacitor c=0.00872971f //x=3.395 //y=0.915
c255 ( 118 0 ) capacitor c=0.0593152f //x=15.91 //y=4.7
c256 ( 109 0 ) capacitor c=0.0588816f //x=5.92 //y=4.7
c257 ( 99 0 ) capacitor c=0.0318948f //x=16.245 //y=1.21
c258 ( 98 0 ) capacitor c=0.0187384f //x=16.245 //y=0.865
c259 ( 95 0 ) capacitor c=0.0141798f //x=16.09 //y=1.365
c260 ( 93 0 ) capacitor c=0.0149844f //x=16.09 //y=0.71
c261 ( 89 0 ) capacitor c=0.0860049f //x=15.715 //y=1.915
c262 ( 88 0 ) capacitor c=0.0229722f //x=15.715 //y=1.52
c263 ( 87 0 ) capacitor c=0.0234352f //x=15.715 //y=1.21
c264 ( 86 0 ) capacitor c=0.0199343f //x=15.715 //y=0.865
c265 ( 82 0 ) capacitor c=0.0318948f //x=6.255 //y=1.21
c266 ( 81 0 ) capacitor c=0.0187384f //x=6.255 //y=0.865
c267 ( 78 0 ) capacitor c=0.0141798f //x=6.1 //y=1.365
c268 ( 76 0 ) capacitor c=0.0149844f //x=6.1 //y=0.71
c269 ( 72 0 ) capacitor c=0.0860049f //x=5.725 //y=1.915
c270 ( 71 0 ) capacitor c=0.0229722f //x=5.725 //y=1.52
c271 ( 70 0 ) capacitor c=0.0234352f //x=5.725 //y=1.21
c272 ( 69 0 ) capacitor c=0.0199343f //x=5.725 //y=0.865
c273 ( 68 0 ) capacitor c=0.110275f //x=16.25 //y=6.02
c274 ( 67 0 ) capacitor c=0.154305f //x=15.81 //y=6.02
c275 ( 66 0 ) capacitor c=0.110275f //x=6.26 //y=6.02
c276 ( 65 0 ) capacitor c=0.154305f //x=5.82 //y=6.02
c277 ( 62 0 ) capacitor c=0.00106608f //x=3.29 //y=5.155
c278 ( 61 0 ) capacitor c=0.00207162f //x=2.41 //y=5.155
c279 ( 54 0 ) capacitor c=0.0963543f //x=15.91 //y=2.08
c280 ( 46 0 ) capacitor c=0.0913801f //x=5.92 //y=2.08
c281 ( 44 0 ) capacitor c=0.109654f //x=4.07 //y=3.7
c282 ( 40 0 ) capacitor c=0.00493499f //x=3.67 //y=1.665
c283 ( 39 0 ) capacitor c=0.0154052f //x=3.985 //y=1.665
c284 ( 33 0 ) capacitor c=0.0284988f //x=3.985 //y=5.155
c285 ( 25 0 ) capacitor c=0.0176454f //x=3.205 //y=5.155
c286 ( 18 0 ) capacitor c=0.00351598f //x=1.615 //y=5.155
c287 ( 17 0 ) capacitor c=0.0154196f //x=2.325 //y=5.155
c288 ( 4 0 ) capacitor c=0.00424317f //x=6.035 //y=3.7
c289 ( 3 0 ) capacitor c=0.222674f //x=15.795 //y=3.7
c290 ( 2 0 ) capacitor c=0.0125346f //x=4.185 //y=3.7
c291 ( 1 0 ) capacitor c=0.0285004f //x=5.805 //y=3.7
r292 (  116 118 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=15.81 //y=4.7 //x2=15.91 //y2=4.7
r293 (  107 109 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=5.82 //y=4.7 //x2=5.92 //y2=4.7
r294 (  100 118 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=16.25 //y=4.865 //x2=15.91 //y2=4.7
r295 (  99 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.245 //y=1.21 //x2=16.205 //y2=1.365
r296 (  98 119 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.245 //y=0.865 //x2=16.205 //y2=0.71
r297 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.245 //y=0.865 //x2=16.245 //y2=1.21
r298 (  96 115 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.87 //y=1.365 //x2=15.755 //y2=1.365
r299 (  95 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.09 //y=1.365 //x2=16.205 //y2=1.365
r300 (  94 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.87 //y=0.71 //x2=15.755 //y2=0.71
r301 (  93 119 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.09 //y=0.71 //x2=16.205 //y2=0.71
r302 (  93 94 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=16.09 //y=0.71 //x2=15.87 //y2=0.71
r303 (  90 116 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=15.81 //y=4.865 //x2=15.81 //y2=4.7
r304 (  89 113 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=15.715 //y=1.915 //x2=15.91 //y2=2.08
r305 (  88 115 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.715 //y=1.52 //x2=15.755 //y2=1.365
r306 (  88 89 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=15.715 //y=1.52 //x2=15.715 //y2=1.915
r307 (  87 115 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.715 //y=1.21 //x2=15.755 //y2=1.365
r308 (  86 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.715 //y=0.865 //x2=15.755 //y2=0.71
r309 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.715 //y=0.865 //x2=15.715 //y2=1.21
r310 (  83 109 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=6.26 //y=4.865 //x2=5.92 //y2=4.7
r311 (  82 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.255 //y=1.21 //x2=6.215 //y2=1.365
r312 (  81 110 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.255 //y=0.865 //x2=6.215 //y2=0.71
r313 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.255 //y=0.865 //x2=6.255 //y2=1.21
r314 (  79 106 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.88 //y=1.365 //x2=5.765 //y2=1.365
r315 (  78 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.1 //y=1.365 //x2=6.215 //y2=1.365
r316 (  77 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.88 //y=0.71 //x2=5.765 //y2=0.71
r317 (  76 110 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.1 //y=0.71 //x2=6.215 //y2=0.71
r318 (  76 77 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=6.1 //y=0.71 //x2=5.88 //y2=0.71
r319 (  73 107 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=5.82 //y=4.865 //x2=5.82 //y2=4.7
r320 (  72 104 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=5.725 //y=1.915 //x2=5.92 //y2=2.08
r321 (  71 106 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.725 //y=1.52 //x2=5.765 //y2=1.365
r322 (  71 72 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=5.725 //y=1.52 //x2=5.725 //y2=1.915
r323 (  70 106 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.725 //y=1.21 //x2=5.765 //y2=1.365
r324 (  69 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.725 //y=0.865 //x2=5.765 //y2=0.71
r325 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.725 //y=0.865 //x2=5.725 //y2=1.21
r326 (  68 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.25 //y=6.02 //x2=16.25 //y2=4.865
r327 (  67 90 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.81 //y=6.02 //x2=15.81 //y2=4.865
r328 (  66 83 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.26 //y=6.02 //x2=6.26 //y2=4.865
r329 (  65 73 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.82 //y=6.02 //x2=5.82 //y2=4.865
r330 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.98 //y=1.365 //x2=16.09 //y2=1.365
r331 (  64 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.98 //y=1.365 //x2=15.87 //y2=1.365
r332 (  63 78 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.99 //y=1.365 //x2=6.1 //y2=1.365
r333 (  63 79 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.99 //y=1.365 //x2=5.88 //y2=1.365
r334 (  59 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.91 //y=4.7 //x2=15.91 //y2=4.7
r335 (  57 59 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=15.91 //y=3.7 //x2=15.91 //y2=4.7
r336 (  54 113 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.91 //y=2.08 //x2=15.91 //y2=2.08
r337 (  54 57 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=15.91 //y=2.08 //x2=15.91 //y2=3.7
r338 (  51 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=4.7 //x2=5.92 //y2=4.7
r339 (  49 51 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=5.92 //y=3.7 //x2=5.92 //y2=4.7
r340 (  46 104 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=2.08 //x2=5.92 //y2=2.08
r341 (  46 49 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.08 //x2=5.92 //y2=3.7
r342 (  42 44 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=4.07 //y=5.07 //x2=4.07 //y2=3.7
r343 (  41 44 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=4.07 //y=1.75 //x2=4.07 //y2=3.7
r344 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=4.07 //y2=1.75
r345 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=3.67 //y2=1.665
r346 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.67 //y2=1.665
r347 (  35 121 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.585 //y2=1.01
r348 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.375 //y=5.155 //x2=3.29 //y2=5.155
r349 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=4.07 //y2=5.07
r350 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=3.375 //y2=5.155
r351 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.155
r352 (  27 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.725
r353 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.495 //y=5.155 //x2=2.41 //y2=5.155
r354 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=3.29 //y2=5.155
r355 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=2.495 //y2=5.155
r356 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.155
r357 (  19 124 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.725
r358 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=2.41 //y2=5.155
r359 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=1.615 //y2=5.155
r360 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.615 //y2=5.155
r361 (  11 123 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.53 //y2=5.725
r362 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.91 //y=3.7 //x2=15.91 //y2=3.7
r363 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.92 //y=3.7 //x2=5.92 //y2=3.7
r364 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=3.7 //x2=4.07 //y2=3.7
r365 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.035 //y=3.7 //x2=5.92 //y2=3.7
r366 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.795 //y=3.7 //x2=15.91 //y2=3.7
r367 (  3 4 ) resistor r=9.31298 //w=0.131 //l=9.76 //layer=m1 \
 //thickness=0.36 //x=15.795 //y=3.7 //x2=6.035 //y2=3.7
r368 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.185 //y=3.7 //x2=4.07 //y2=3.7
r369 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.805 //y=3.7 //x2=5.92 //y2=3.7
r370 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=5.805 //y=3.7 //x2=4.185 //y2=3.7
ends PM_DFFX1_PCELL\%noxref_6

subckt PM_DFFX1_PCELL\%noxref_7 ( 1 2 3 4 5 6 16 23 25 35 36 47 49 50 54 55 57 \
 63 66 67 68 69 70 71 72 73 74 75 76 77 78 79 81 87 88 89 90 94 95 96 101 103 \
 105 111 112 113 114 115 120 122 124 130 131 141 142 145 154 155 158 166 168 \
 169 )
c356 ( 169 0 ) capacitor c=0.0220291f //x=13.435 //y=5.02
c357 ( 168 0 ) capacitor c=0.0217503f //x=12.555 //y=5.02
c358 ( 166 0 ) capacitor c=0.00866655f //x=13.43 //y=0.905
c359 ( 158 0 ) capacitor c=0.0335797f //x=20.01 //y=4.7
c360 ( 155 0 ) capacitor c=0.0279499f //x=19.98 //y=1.915
c361 ( 154 0 ) capacitor c=0.0437302f //x=19.98 //y=2.08
c362 ( 145 0 ) capacitor c=0.0331095f //x=10.02 //y=4.7
c363 ( 142 0 ) capacitor c=0.0279499f //x=9.99 //y=1.915
c364 ( 141 0 ) capacitor c=0.0437302f //x=9.99 //y=2.08
c365 ( 131 0 ) capacitor c=0.0429696f //x=20.545 //y=1.25
c366 ( 130 0 ) capacitor c=0.0192208f //x=20.545 //y=0.905
c367 ( 124 0 ) capacitor c=0.0158629f //x=20.39 //y=1.405
c368 ( 122 0 ) capacitor c=0.0157803f //x=20.39 //y=0.75
c369 ( 120 0 ) capacitor c=0.0366192f //x=20.385 //y=4.79
c370 ( 115 0 ) capacitor c=0.0205163f //x=20.015 //y=1.56
c371 ( 114 0 ) capacitor c=0.0168481f //x=20.015 //y=1.25
c372 ( 113 0 ) capacitor c=0.0174783f //x=20.015 //y=0.905
c373 ( 112 0 ) capacitor c=0.0429696f //x=10.555 //y=1.25
c374 ( 111 0 ) capacitor c=0.0192208f //x=10.555 //y=0.905
c375 ( 105 0 ) capacitor c=0.0158629f //x=10.4 //y=1.405
c376 ( 103 0 ) capacitor c=0.0157803f //x=10.4 //y=0.75
c377 ( 101 0 ) capacitor c=0.0295235f //x=10.395 //y=4.79
c378 ( 96 0 ) capacitor c=0.0205163f //x=10.025 //y=1.56
c379 ( 95 0 ) capacitor c=0.0168481f //x=10.025 //y=1.25
c380 ( 94 0 ) capacitor c=0.0174783f //x=10.025 //y=0.905
c381 ( 90 0 ) capacitor c=0.0559896f //x=1.385 //y=4.79
c382 ( 89 0 ) capacitor c=0.0298189f //x=1.675 //y=4.79
c383 ( 88 0 ) capacitor c=0.0347816f //x=1.34 //y=1.22
c384 ( 87 0 ) capacitor c=0.0187487f //x=1.34 //y=0.875
c385 ( 81 0 ) capacitor c=0.0137055f //x=1.185 //y=1.375
c386 ( 79 0 ) capacitor c=0.0149861f //x=1.185 //y=0.72
c387 ( 78 0 ) capacitor c=0.102158f //x=0.81 //y=1.915
c388 ( 77 0 ) capacitor c=0.0229444f //x=0.81 //y=1.53
c389 ( 76 0 ) capacitor c=0.0234352f //x=0.81 //y=1.22
c390 ( 75 0 ) capacitor c=0.0198724f //x=0.81 //y=0.875
c391 ( 74 0 ) capacitor c=0.15358f //x=20.46 //y=6.02
c392 ( 73 0 ) capacitor c=0.110281f //x=20.02 //y=6.02
c393 ( 72 0 ) capacitor c=0.15358f //x=10.47 //y=6.02
c394 ( 71 0 ) capacitor c=0.110281f //x=10.03 //y=6.02
c395 ( 70 0 ) capacitor c=0.110114f //x=1.75 //y=6.02
c396 ( 69 0 ) capacitor c=0.158956f //x=1.31 //y=6.02
c397 ( 63 0 ) capacitor c=0.0023043f //x=13.58 //y=5.2
c398 ( 57 0 ) capacitor c=0.0796561f //x=19.98 //y=2.08
c399 ( 55 0 ) capacitor c=0.00453889f //x=19.98 //y=4.535
c400 ( 54 0 ) capacitor c=0.111855f //x=14.06 //y=4.07
c401 ( 50 0 ) capacitor c=0.00525782f //x=13.705 //y=1.655
c402 ( 49 0 ) capacitor c=0.0140405f //x=13.975 //y=1.655
c403 ( 47 0 ) capacitor c=0.0140419f //x=13.975 //y=5.2
c404 ( 36 0 ) capacitor c=0.00251459f //x=12.785 //y=5.2
c405 ( 35 0 ) capacitor c=0.0143111f //x=13.495 //y=5.2
c406 ( 25 0 ) capacitor c=0.0739568f //x=9.99 //y=2.08
c407 ( 23 0 ) capacitor c=0.00453889f //x=9.99 //y=4.535
c408 ( 16 0 ) capacitor c=0.124161f //x=1.11 //y=2.08
c409 ( 6 0 ) capacitor c=0.00579158f //x=14.175 //y=4.07
c410 ( 5 0 ) capacitor c=0.23267f //x=19.865 //y=4.07
c411 ( 4 0 ) capacitor c=0.00412846f //x=10.105 //y=4.07
c412 ( 3 0 ) capacitor c=0.0575173f //x=13.945 //y=4.07
c413 ( 2 0 ) capacitor c=0.0160831f //x=1.225 //y=4.07
c414 ( 1 0 ) capacitor c=0.163286f //x=9.875 //y=4.07
r415 (  160 161 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=20.01 //y=4.79 //x2=20.01 //y2=4.865
r416 (  158 160 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=20.01 //y=4.7 //x2=20.01 //y2=4.79
r417 (  154 155 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=19.98 //y=2.08 //x2=19.98 //y2=1.915
r418 (  147 148 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=10.02 //y=4.79 //x2=10.02 //y2=4.865
r419 (  145 147 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=10.02 //y=4.7 //x2=10.02 //y2=4.79
r420 (  141 142 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=9.99 //y=2.08 //x2=9.99 //y2=1.915
r421 (  131 165 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.545 //y=1.25 //x2=20.505 //y2=1.405
r422 (  130 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.545 //y=0.905 //x2=20.505 //y2=0.75
r423 (  130 131 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.545 //y=0.905 //x2=20.545 //y2=1.25
r424 (  125 163 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.17 //y=1.405 //x2=20.055 //y2=1.405
r425 (  124 165 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.39 //y=1.405 //x2=20.505 //y2=1.405
r426 (  123 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.17 //y=0.75 //x2=20.055 //y2=0.75
r427 (  122 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.39 //y=0.75 //x2=20.505 //y2=0.75
r428 (  122 123 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=20.39 //y=0.75 //x2=20.17 //y2=0.75
r429 (  121 160 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=20.145 //y=4.79 //x2=20.01 //y2=4.79
r430 (  120 127 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.385 //y=4.79 //x2=20.46 //y2=4.865
r431 (  120 121 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=20.385 //y=4.79 //x2=20.145 //y2=4.79
r432 (  115 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.015 //y=1.56 //x2=20.055 //y2=1.405
r433 (  115 155 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=20.015 //y=1.56 //x2=20.015 //y2=1.915
r434 (  114 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.015 //y=1.25 //x2=20.055 //y2=1.405
r435 (  113 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.015 //y=0.905 //x2=20.055 //y2=0.75
r436 (  113 114 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.015 //y=0.905 //x2=20.015 //y2=1.25
r437 (  112 152 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.555 //y=1.25 //x2=10.515 //y2=1.405
r438 (  111 151 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.555 //y=0.905 //x2=10.515 //y2=0.75
r439 (  111 112 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.555 //y=0.905 //x2=10.555 //y2=1.25
r440 (  106 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.18 //y=1.405 //x2=10.065 //y2=1.405
r441 (  105 152 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.4 //y=1.405 //x2=10.515 //y2=1.405
r442 (  104 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.18 //y=0.75 //x2=10.065 //y2=0.75
r443 (  103 151 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.4 //y=0.75 //x2=10.515 //y2=0.75
r444 (  103 104 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.4 //y=0.75 //x2=10.18 //y2=0.75
r445 (  102 147 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=10.155 //y=4.79 //x2=10.02 //y2=4.79
r446 (  101 108 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.395 //y=4.79 //x2=10.47 //y2=4.865
r447 (  101 102 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=10.395 //y=4.79 //x2=10.155 //y2=4.79
r448 (  96 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.025 //y=1.56 //x2=10.065 //y2=1.405
r449 (  96 142 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=10.025 //y=1.56 //x2=10.025 //y2=1.915
r450 (  95 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.025 //y=1.25 //x2=10.065 //y2=1.405
r451 (  94 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.025 //y=0.905 //x2=10.065 //y2=0.75
r452 (  94 95 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.025 //y=0.905 //x2=10.025 //y2=1.25
r453 (  89 91 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.75 //y2=4.865
r454 (  89 90 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.385 //y2=4.79
r455 (  88 139 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=1.22 //x2=1.3 //y2=1.375
r456 (  87 138 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.3 //y2=0.72
r457 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.34 //y2=1.22
r458 (  84 90 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.385 //y2=4.79
r459 (  84 137 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.11 //y2=4.7
r460 (  82 133 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=1.375 //x2=0.85 //y2=1.375
r461 (  81 139 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=1.375 //x2=1.3 //y2=1.375
r462 (  80 132 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=0.72 //x2=0.85 //y2=0.72
r463 (  79 138 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=1.3 //y2=0.72
r464 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=0.965 //y2=0.72
r465 (  78 135 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.915 //x2=1.11 //y2=2.08
r466 (  77 133 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.85 //y2=1.375
r467 (  77 78 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.81 //y2=1.915
r468 (  76 133 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.22 //x2=0.85 //y2=1.375
r469 (  75 132 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.85 //y2=0.72
r470 (  75 76 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.81 //y2=1.22
r471 (  74 127 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.46 //y=6.02 //x2=20.46 //y2=4.865
r472 (  73 161 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.02 //y=6.02 //x2=20.02 //y2=4.865
r473 (  72 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.47 //y=6.02 //x2=10.47 //y2=4.865
r474 (  71 148 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.03 //y=6.02 //x2=10.03 //y2=4.865
r475 (  70 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.75 //y=6.02 //x2=1.75 //y2=4.865
r476 (  69 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.31 //y=6.02 //x2=1.31 //y2=4.865
r477 (  68 124 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.28 //y=1.405 //x2=20.39 //y2=1.405
r478 (  68 125 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.28 //y=1.405 //x2=20.17 //y2=1.405
r479 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.29 //y=1.405 //x2=10.4 //y2=1.405
r480 (  67 106 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.29 //y=1.405 //x2=10.18 //y2=1.405
r481 (  66 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=1.185 //y2=1.375
r482 (  66 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=0.965 //y2=1.375
r483 (  65 158 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.01 //y=4.7 //x2=20.01 //y2=4.7
r484 (  62 145 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.02 //y=4.7 //x2=10.02 //y2=4.7
r485 (  57 154 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.98 //y=2.08 //x2=19.98 //y2=2.08
r486 (  57 60 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.08 //x2=19.98 //y2=4.07
r487 (  55 65 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=19.98 //y=4.535 //x2=19.995 //y2=4.7
r488 (  55 60 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=19.98 //y=4.535 //x2=19.98 //y2=4.07
r489 (  52 54 ) resistor r=71.5294 //w=0.187 //l=1.045 //layer=li \
 //thickness=0.1 //x=14.06 //y=5.115 //x2=14.06 //y2=4.07
r490 (  51 54 ) resistor r=159.487 //w=0.187 //l=2.33 //layer=li \
 //thickness=0.1 //x=14.06 //y=1.74 //x2=14.06 //y2=4.07
r491 (  49 51 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.975 //y=1.655 //x2=14.06 //y2=1.74
r492 (  49 50 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=13.975 //y=1.655 //x2=13.705 //y2=1.655
r493 (  48 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.665 //y=5.2 //x2=13.58 //y2=5.2
r494 (  47 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.975 //y=5.2 //x2=14.06 //y2=5.115
r495 (  47 48 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=13.975 //y=5.2 //x2=13.665 //y2=5.2
r496 (  43 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.62 //y=1.57 //x2=13.705 //y2=1.655
r497 (  43 166 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=13.62 //y=1.57 //x2=13.62 //y2=1
r498 (  37 63 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.58 //y=5.285 //x2=13.58 //y2=5.2
r499 (  37 169 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=13.58 //y=5.285 //x2=13.58 //y2=5.725
r500 (  35 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.495 //y=5.2 //x2=13.58 //y2=5.2
r501 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=13.495 //y=5.2 //x2=12.785 //y2=5.2
r502 (  29 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.7 //y=5.285 //x2=12.785 //y2=5.2
r503 (  29 168 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=12.7 //y=5.285 //x2=12.7 //y2=5.725
r504 (  25 141 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.99 //y=2.08 //x2=9.99 //y2=2.08
r505 (  25 28 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=9.99 //y=2.08 //x2=9.99 //y2=4.07
r506 (  23 62 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=9.99 //y=4.535 //x2=10.005 //y2=4.7
r507 (  23 28 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=9.99 //y=4.535 //x2=9.99 //y2=4.07
r508 (  21 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r509 (  19 21 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.07 //x2=1.11 //y2=4.7
r510 (  16 135 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r511 (  16 19 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.08 //x2=1.11 //y2=4.07
r512 (  14 60 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=19.98 //y=4.07 //x2=19.98 //y2=4.07
r513 (  12 54 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.06 //y=4.07 //x2=14.06 //y2=4.07
r514 (  10 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.99 //y=4.07 //x2=9.99 //y2=4.07
r515 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.07
r516 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=14.175 //y=4.07 //x2=14.06 //y2=4.07
r517 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=19.865 //y=4.07 //x2=19.98 //y2=4.07
r518 (  5 6 ) resistor r=5.42939 //w=0.131 //l=5.69 //layer=m1 \
 //thickness=0.36 //x=19.865 //y=4.07 //x2=14.175 //y2=4.07
r519 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.105 //y=4.07 //x2=9.99 //y2=4.07
r520 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=4.07 //x2=14.06 //y2=4.07
r521 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=4.07 //x2=10.105 //y2=4.07
r522 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.225 //y=4.07 //x2=1.11 //y2=4.07
r523 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.875 //y=4.07 //x2=9.99 //y2=4.07
r524 (  1 2 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=9.875 //y=4.07 //x2=1.225 //y2=4.07
ends PM_DFFX1_PCELL\%noxref_7

subckt PM_DFFX1_PCELL\%noxref_8 ( 1 5 9 13 17 35 )
c47 ( 35 0 ) capacitor c=0.0703709f //x=0.455 //y=0.375
c48 ( 17 0 ) capacitor c=0.0221229f //x=2.445 //y=1.59
c49 ( 13 0 ) capacitor c=0.0156939f //x=2.445 //y=0.54
c50 ( 9 0 ) capacitor c=0.00678203f //x=1.56 //y=0.625
c51 ( 5 0 ) capacitor c=0.0206412f //x=1.475 //y=1.59
c52 ( 1 0 ) capacitor c=0.0109947f //x=0.59 //y=1.505
r53 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=1.59 //x2=1.56 //y2=1.63
r54 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=1.59 //x2=2.045 //y2=1.59
r55 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=1.59 //x2=2.53 //y2=1.59
r56 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=1.59 //x2=2.045 //y2=1.59
r57 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=0.54 //x2=1.56 //y2=0.5
r58 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=0.54 //x2=2.045 //y2=0.54
r59 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=0.54 //x2=2.53 //y2=0.54
r60 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=0.54 //x2=2.045 //y2=0.54
r61 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=1.63
r62 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=0.89
r63 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.5
r64 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.89
r65 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.675 //y=1.59 //x2=0.59 //y2=1.63
r66 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.675 //y=1.59 //x2=1.075 //y2=1.59
r67 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.475 //y=1.59 //x2=1.56 //y2=1.63
r68 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.475 //y=1.59 //x2=1.075 //y2=1.59
r69 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.59 //y=1.505 //x2=0.59 //y2=1.63
r70 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.59 //y=1.505 //x2=0.59 //y2=0.89
ends PM_DFFX1_PCELL\%noxref_8

subckt PM_DFFX1_PCELL\%noxref_9 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.043074f //x=2.965 //y=0.375
c54 ( 28 0 ) capacitor c=0.00465142f //x=1.86 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=3.1 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=4.07 //y=0.625
c57 ( 11 0 ) capacitor c=0.0149771f //x=3.985 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=3.1 //y=0.625
c59 ( 1 0 ) capacitor c=0.0253322f //x=3.015 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.185 //y=0.54 //x2=3.1 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.185 //y=0.54 //x2=3.585 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.985 //y=0.54 //x2=4.07 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.985 //y=0.54 //x2=3.585 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.135 //y=0.995 //x2=2.05 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=3.1 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=2.135 //y2=0.995
ends PM_DFFX1_PCELL\%noxref_9

subckt PM_DFFX1_PCELL\%noxref_10 ( 1 3 7 8 9 10 11 12 17 19 21 27 28 30 31 34 )
c73 ( 34 0 ) capacitor c=0.0331095f //x=6.69 //y=4.7
c74 ( 31 0 ) capacitor c=0.0279499f //x=6.66 //y=1.915
c75 ( 30 0 ) capacitor c=0.0437302f //x=6.66 //y=2.08
c76 ( 28 0 ) capacitor c=0.0429696f //x=7.225 //y=1.25
c77 ( 27 0 ) capacitor c=0.0192208f //x=7.225 //y=0.905
c78 ( 21 0 ) capacitor c=0.0158629f //x=7.07 //y=1.405
c79 ( 19 0 ) capacitor c=0.0157803f //x=7.07 //y=0.75
c80 ( 17 0 ) capacitor c=0.0295235f //x=7.065 //y=4.79
c81 ( 12 0 ) capacitor c=0.0205163f //x=6.695 //y=1.56
c82 ( 11 0 ) capacitor c=0.0168481f //x=6.695 //y=1.25
c83 ( 10 0 ) capacitor c=0.0174783f //x=6.695 //y=0.905
c84 ( 9 0 ) capacitor c=0.15358f //x=7.14 //y=6.02
c85 ( 8 0 ) capacitor c=0.110281f //x=6.7 //y=6.02
c86 ( 3 0 ) capacitor c=0.0737925f //x=6.66 //y=2.08
c87 ( 1 0 ) capacitor c=0.00453889f //x=6.66 //y=4.535
r88 (  36 37 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=6.69 //y=4.79 //x2=6.69 //y2=4.865
r89 (  34 36 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=6.69 //y=4.7 //x2=6.69 //y2=4.79
r90 (  30 31 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.66 //y=2.08 //x2=6.66 //y2=1.915
r91 (  28 41 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.225 //y=1.25 //x2=7.185 //y2=1.405
r92 (  27 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.225 //y=0.905 //x2=7.185 //y2=0.75
r93 (  27 28 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.225 //y=0.905 //x2=7.225 //y2=1.25
r94 (  22 39 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.85 //y=1.405 //x2=6.735 //y2=1.405
r95 (  21 41 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.07 //y=1.405 //x2=7.185 //y2=1.405
r96 (  20 38 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.85 //y=0.75 //x2=6.735 //y2=0.75
r97 (  19 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.07 //y=0.75 //x2=7.185 //y2=0.75
r98 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.07 //y=0.75 //x2=6.85 //y2=0.75
r99 (  18 36 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=6.825 //y=4.79 //x2=6.69 //y2=4.79
r100 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.065 //y=4.79 //x2=7.14 //y2=4.865
r101 (  17 18 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=7.065 //y=4.79 //x2=6.825 //y2=4.79
r102 (  12 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.695 //y=1.56 //x2=6.735 //y2=1.405
r103 (  12 31 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=6.695 //y=1.56 //x2=6.695 //y2=1.915
r104 (  11 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.695 //y=1.25 //x2=6.735 //y2=1.405
r105 (  10 38 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.695 //y=0.905 //x2=6.735 //y2=0.75
r106 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.695 //y=0.905 //x2=6.695 //y2=1.25
r107 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.14 //y=6.02 //x2=7.14 //y2=4.865
r108 (  8 37 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.7 //y=6.02 //x2=6.7 //y2=4.865
r109 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.96 //y=1.405 //x2=7.07 //y2=1.405
r110 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.96 //y=1.405 //x2=6.85 //y2=1.405
r111 (  6 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.69 //y=4.7 //x2=6.69 //y2=4.7
r112 (  3 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=2.08 //x2=6.66 //y2=2.08
r113 (  1 6 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=6.66 //y=4.535 //x2=6.675 //y2=4.7
r114 (  1 3 ) resistor r=168.043 //w=0.187 //l=2.455 //layer=li \
 //thickness=0.1 //x=6.66 //y=4.535 //x2=6.66 //y2=2.08
ends PM_DFFX1_PCELL\%noxref_10

subckt PM_DFFX1_PCELL\%noxref_11 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0638069f //x=5.37 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=7.445 //y=0.615
c54 ( 13 0 ) capacitor c=0.0148848f //x=7.36 //y=0.53
c55 ( 10 0 ) capacitor c=0.00664066f //x=6.475 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=6.475 //y=0.615
c57 ( 5 0 ) capacitor c=0.0196287f //x=6.39 //y=1.58
c58 ( 1 0 ) capacitor c=0.00828748f //x=5.505 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=7.445 //y=0.615 //x2=7.445 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=7.445 //y=0.615 //x2=7.445 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.56 //y=0.53 //x2=6.475 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.56 //y=0.53 //x2=6.96 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.36 //y=0.53 //x2=7.445 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.36 //y=0.53 //x2=6.96 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=6.475 //y=1.495 //x2=6.475 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.475 //y=1.495 //x2=6.475 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.475 //y=0.615 //x2=6.475 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.475 //y=0.615 //x2=6.475 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.59 //y=1.58 //x2=5.505 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.59 //y=1.58 //x2=5.99 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.39 //y=1.58 //x2=6.475 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.39 //y=1.58 //x2=5.99 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=5.505 //y=1.495 //x2=5.505 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=5.505 //y=1.495 //x2=5.505 //y2=0.88
ends PM_DFFX1_PCELL\%noxref_11

subckt PM_DFFX1_PCELL\%noxref_12 ( 1 5 9 10 13 17 29 )
c53 ( 29 0 ) capacitor c=0.0638071f //x=8.7 //y=0.365
c54 ( 17 0 ) capacitor c=0.00722223f //x=10.775 //y=0.615
c55 ( 13 0 ) capacitor c=0.0149613f //x=10.69 //y=0.53
c56 ( 10 0 ) capacitor c=0.00687696f //x=9.805 //y=1.495
c57 ( 9 0 ) capacitor c=0.006761f //x=9.805 //y=0.615
c58 ( 5 0 ) capacitor c=0.0201208f //x=9.72 //y=1.58
c59 ( 1 0 ) capacitor c=0.00828748f //x=8.835 //y=1.495
r60 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=10.775 //y=0.615 //x2=10.775 //y2=0.49
r61 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=10.775 //y=0.615 //x2=10.775 //y2=0.88
r62 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.89 //y=0.53 //x2=9.805 //y2=0.49
r63 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.89 //y=0.53 //x2=10.29 //y2=0.53
r64 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.69 //y=0.53 //x2=10.775 //y2=0.49
r65 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.69 //y=0.53 //x2=10.29 //y2=0.53
r66 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=9.805 //y=1.495 //x2=9.805 //y2=1.62
r67 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=9.805 //y=1.495 //x2=9.805 //y2=0.88
r68 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=9.805 //y=0.615 //x2=9.805 //y2=0.49
r69 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=9.805 //y=0.615 //x2=9.805 //y2=0.88
r70 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.92 //y=1.58 //x2=8.835 //y2=1.62
r71 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.92 //y=1.58 //x2=9.32 //y2=1.58
r72 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.72 //y=1.58 //x2=9.805 //y2=1.62
r73 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.72 //y=1.58 //x2=9.32 //y2=1.58
r74 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=8.835 //y=1.495 //x2=8.835 //y2=1.62
r75 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=8.835 //y=1.495 //x2=8.835 //y2=0.88
ends PM_DFFX1_PCELL\%noxref_12

subckt PM_DFFX1_PCELL\%noxref_13 ( 1 5 9 10 13 17 29 )
c53 ( 29 0 ) capacitor c=0.0637486f //x=12.03 //y=0.365
c54 ( 17 0 ) capacitor c=0.00722223f //x=14.105 //y=0.615
c55 ( 13 0 ) capacitor c=0.0149666f //x=14.02 //y=0.53
c56 ( 10 0 ) capacitor c=0.00687696f //x=13.135 //y=1.495
c57 ( 9 0 ) capacitor c=0.006761f //x=13.135 //y=0.615
c58 ( 5 0 ) capacitor c=0.0201208f //x=13.05 //y=1.58
c59 ( 1 0 ) capacitor c=0.00828748f //x=12.165 //y=1.495
r60 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=14.105 //y=0.615 //x2=14.105 //y2=0.49
r61 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=14.105 //y=0.615 //x2=14.105 //y2=0.88
r62 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.22 //y=0.53 //x2=13.135 //y2=0.49
r63 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.22 //y=0.53 //x2=13.62 //y2=0.53
r64 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.02 //y=0.53 //x2=14.105 //y2=0.49
r65 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.02 //y=0.53 //x2=13.62 //y2=0.53
r66 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=13.135 //y=1.495 //x2=13.135 //y2=1.62
r67 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=13.135 //y=1.495 //x2=13.135 //y2=0.88
r68 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=13.135 //y=0.615 //x2=13.135 //y2=0.49
r69 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=13.135 //y=0.615 //x2=13.135 //y2=0.88
r70 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.25 //y=1.58 //x2=12.165 //y2=1.62
r71 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.25 //y=1.58 //x2=12.65 //y2=1.58
r72 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.05 //y=1.58 //x2=13.135 //y2=1.62
r73 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.05 //y=1.58 //x2=12.65 //y2=1.58
r74 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=12.165 //y=1.495 //x2=12.165 //y2=1.62
r75 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=12.165 //y=1.495 //x2=12.165 //y2=0.88
ends PM_DFFX1_PCELL\%noxref_13

subckt PM_DFFX1_PCELL\%noxref_14 ( 1 3 7 8 9 10 11 12 17 19 21 27 28 30 31 34 )
c69 ( 34 0 ) capacitor c=0.0331552f //x=16.68 //y=4.7
c70 ( 31 0 ) capacitor c=0.0279499f //x=16.65 //y=1.915
c71 ( 30 0 ) capacitor c=0.0437302f //x=16.65 //y=2.08
c72 ( 28 0 ) capacitor c=0.0429696f //x=17.215 //y=1.25
c73 ( 27 0 ) capacitor c=0.0192208f //x=17.215 //y=0.905
c74 ( 21 0 ) capacitor c=0.0158629f //x=17.06 //y=1.405
c75 ( 19 0 ) capacitor c=0.0157803f //x=17.06 //y=0.75
c76 ( 17 0 ) capacitor c=0.0299681f //x=17.055 //y=4.79
c77 ( 12 0 ) capacitor c=0.0205163f //x=16.685 //y=1.56
c78 ( 11 0 ) capacitor c=0.0168481f //x=16.685 //y=1.25
c79 ( 10 0 ) capacitor c=0.0174783f //x=16.685 //y=0.905
c80 ( 9 0 ) capacitor c=0.15358f //x=17.13 //y=6.02
c81 ( 8 0 ) capacitor c=0.110281f //x=16.69 //y=6.02
c82 ( 3 0 ) capacitor c=0.079216f //x=16.65 //y=2.08
c83 ( 1 0 ) capacitor c=0.00453889f //x=16.65 //y=4.535
r84 (  36 37 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=16.68 //y=4.79 //x2=16.68 //y2=4.865
r85 (  34 36 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=16.68 //y=4.7 //x2=16.68 //y2=4.79
r86 (  30 31 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=16.65 //y=2.08 //x2=16.65 //y2=1.915
r87 (  28 41 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.215 //y=1.25 //x2=17.175 //y2=1.405
r88 (  27 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.215 //y=0.905 //x2=17.175 //y2=0.75
r89 (  27 28 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.215 //y=0.905 //x2=17.215 //y2=1.25
r90 (  22 39 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.84 //y=1.405 //x2=16.725 //y2=1.405
r91 (  21 41 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.06 //y=1.405 //x2=17.175 //y2=1.405
r92 (  20 38 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.84 //y=0.75 //x2=16.725 //y2=0.75
r93 (  19 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.06 //y=0.75 //x2=17.175 //y2=0.75
r94 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=17.06 //y=0.75 //x2=16.84 //y2=0.75
r95 (  18 36 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=16.815 //y=4.79 //x2=16.68 //y2=4.79
r96 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=17.055 //y=4.79 //x2=17.13 //y2=4.865
r97 (  17 18 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=17.055 //y=4.79 //x2=16.815 //y2=4.79
r98 (  12 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.685 //y=1.56 //x2=16.725 //y2=1.405
r99 (  12 31 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=16.685 //y=1.56 //x2=16.685 //y2=1.915
r100 (  11 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.685 //y=1.25 //x2=16.725 //y2=1.405
r101 (  10 38 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.685 //y=0.905 //x2=16.725 //y2=0.75
r102 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.685 //y=0.905 //x2=16.685 //y2=1.25
r103 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.13 //y=6.02 //x2=17.13 //y2=4.865
r104 (  8 37 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.69 //y=6.02 //x2=16.69 //y2=4.865
r105 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=16.95 //y=1.405 //x2=17.06 //y2=1.405
r106 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=16.95 //y=1.405 //x2=16.84 //y2=1.405
r107 (  6 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.68 //y=4.7 //x2=16.68 //y2=4.7
r108 (  3 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.65 //y=2.08 //x2=16.65 //y2=2.08
r109 (  1 6 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=16.65 //y=4.535 //x2=16.665 //y2=4.7
r110 (  1 3 ) resistor r=168.043 //w=0.187 //l=2.455 //layer=li \
 //thickness=0.1 //x=16.65 //y=4.535 //x2=16.65 //y2=2.08
ends PM_DFFX1_PCELL\%noxref_14

subckt PM_DFFX1_PCELL\%noxref_15 ( 7 8 19 21 22 24 25 26 28 29 )
c72 ( 29 0 ) capacitor c=0.0220291f //x=16.765 //y=5.02
c73 ( 28 0 ) capacitor c=0.0217503f //x=15.885 //y=5.02
c74 ( 26 0 ) capacitor c=0.00866655f //x=16.76 //y=0.905
c75 ( 25 0 ) capacitor c=0.0023043f //x=16.91 //y=5.2
c76 ( 24 0 ) capacitor c=0.116717f //x=17.39 //y=5.115
c77 ( 22 0 ) capacitor c=0.00550359f //x=17.035 //y=1.655
c78 ( 21 0 ) capacitor c=0.0144081f //x=17.305 //y=1.655
c79 ( 19 0 ) capacitor c=0.0140462f //x=17.305 //y=5.2
c80 ( 8 0 ) capacitor c=0.00265417f //x=16.115 //y=5.2
c81 ( 7 0 ) capacitor c=0.0149089f //x=16.825 //y=5.2
r82 (  23 24 ) resistor r=231.016 //w=0.187 //l=3.375 //layer=li \
 //thickness=0.1 //x=17.39 //y=1.74 //x2=17.39 //y2=5.115
r83 (  21 23 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.305 //y=1.655 //x2=17.39 //y2=1.74
r84 (  21 22 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=17.305 //y=1.655 //x2=17.035 //y2=1.655
r85 (  20 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=16.995 //y=5.2 //x2=16.91 //y2=5.2
r86 (  19 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.305 //y=5.2 //x2=17.39 //y2=5.115
r87 (  19 20 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=17.305 //y=5.2 //x2=16.995 //y2=5.2
r88 (  15 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.95 //y=1.57 //x2=17.035 //y2=1.655
r89 (  15 26 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=16.95 //y=1.57 //x2=16.95 //y2=1
r90 (  9 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=16.91 //y=5.285 //x2=16.91 //y2=5.2
r91 (  9 29 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li //thickness=0.1 \
 //x=16.91 //y=5.285 //x2=16.91 //y2=5.725
r92 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=16.825 //y=5.2 //x2=16.91 //y2=5.2
r93 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=16.825 //y=5.2 //x2=16.115 //y2=5.2
r94 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.03 //y=5.285 //x2=16.115 //y2=5.2
r95 (  1 28 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li //thickness=0.1 \
 //x=16.03 //y=5.285 //x2=16.03 //y2=5.725
ends PM_DFFX1_PCELL\%noxref_15

subckt PM_DFFX1_PCELL\%noxref_16 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0638269f //x=15.36 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=17.435 //y=0.615
c54 ( 13 0 ) capacitor c=0.0154622f //x=17.35 //y=0.53
c55 ( 10 0 ) capacitor c=0.00709043f //x=16.465 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=16.465 //y=0.615
c57 ( 5 0 ) capacitor c=0.0207245f //x=16.38 //y=1.58
c58 ( 1 0 ) capacitor c=0.00856252f //x=15.495 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=17.435 //y=0.615 //x2=17.435 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=17.435 //y=0.615 //x2=17.435 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.55 //y=0.53 //x2=16.465 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.55 //y=0.53 //x2=16.95 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.35 //y=0.53 //x2=17.435 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.35 //y=0.53 //x2=16.95 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=16.465 //y=1.495 //x2=16.465 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=16.465 //y=1.495 //x2=16.465 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=16.465 //y=0.615 //x2=16.465 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=16.465 //y=0.615 //x2=16.465 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.58 //y=1.58 //x2=15.495 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.58 //y=1.58 //x2=15.98 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.38 //y=1.58 //x2=16.465 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.38 //y=1.58 //x2=15.98 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=15.495 //y=1.495 //x2=15.495 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=15.495 //y=1.495 //x2=15.495 //y2=0.88
ends PM_DFFX1_PCELL\%noxref_16

subckt PM_DFFX1_PCELL\%noxref_17 ( 2 7 8 9 10 11 12 13 17 19 22 23 33 )
c60 ( 33 0 ) capacitor c=0.0593152f //x=19.24 //y=4.7
c61 ( 23 0 ) capacitor c=0.0318948f //x=19.575 //y=1.21
c62 ( 22 0 ) capacitor c=0.0187384f //x=19.575 //y=0.865
c63 ( 19 0 ) capacitor c=0.0141798f //x=19.42 //y=1.365
c64 ( 17 0 ) capacitor c=0.0149844f //x=19.42 //y=0.71
c65 ( 13 0 ) capacitor c=0.0860049f //x=19.045 //y=1.915
c66 ( 12 0 ) capacitor c=0.0229722f //x=19.045 //y=1.52
c67 ( 11 0 ) capacitor c=0.0234352f //x=19.045 //y=1.21
c68 ( 10 0 ) capacitor c=0.0199343f //x=19.045 //y=0.865
c69 ( 9 0 ) capacitor c=0.110275f //x=19.58 //y=6.02
c70 ( 8 0 ) capacitor c=0.154305f //x=19.14 //y=6.02
c71 ( 2 0 ) capacitor c=0.100185f //x=19.24 //y=2.08
r72 (  31 33 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=19.14 //y=4.7 //x2=19.24 //y2=4.7
r73 (  24 33 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=19.58 //y=4.865 //x2=19.24 //y2=4.7
r74 (  23 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.575 //y=1.21 //x2=19.535 //y2=1.365
r75 (  22 34 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.575 //y=0.865 //x2=19.535 //y2=0.71
r76 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=19.575 //y=0.865 //x2=19.575 //y2=1.21
r77 (  20 30 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.2 //y=1.365 //x2=19.085 //y2=1.365
r78 (  19 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.42 //y=1.365 //x2=19.535 //y2=1.365
r79 (  18 29 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.2 //y=0.71 //x2=19.085 //y2=0.71
r80 (  17 34 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.42 //y=0.71 //x2=19.535 //y2=0.71
r81 (  17 18 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=19.42 //y=0.71 //x2=19.2 //y2=0.71
r82 (  14 31 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=19.14 //y=4.865 //x2=19.14 //y2=4.7
r83 (  13 28 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=19.045 //y=1.915 //x2=19.24 //y2=2.08
r84 (  12 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.045 //y=1.52 //x2=19.085 //y2=1.365
r85 (  12 13 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=19.045 //y=1.52 //x2=19.045 //y2=1.915
r86 (  11 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.045 //y=1.21 //x2=19.085 //y2=1.365
r87 (  10 29 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.045 //y=0.865 //x2=19.085 //y2=0.71
r88 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=19.045 //y=0.865 //x2=19.045 //y2=1.21
r89 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.58 //y=6.02 //x2=19.58 //y2=4.865
r90 (  8 14 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.14 //y=6.02 //x2=19.14 //y2=4.865
r91 (  7 19 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=19.31 //y=1.365 //x2=19.42 //y2=1.365
r92 (  7 20 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=19.31 //y=1.365 //x2=19.2 //y2=1.365
r93 (  5 33 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.24 //y=4.7 //x2=19.24 //y2=4.7
r94 (  2 28 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.24 //y=2.08 //x2=19.24 //y2=2.08
r95 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=19.24 //y=2.08 //x2=19.24 //y2=4.7
ends PM_DFFX1_PCELL\%noxref_17

subckt PM_DFFX1_PCELL\%noxref_18 ( 7 8 19 21 22 24 25 26 28 29 )
c65 ( 29 0 ) capacitor c=0.0220291f //x=20.095 //y=5.02
c66 ( 28 0 ) capacitor c=0.0217503f //x=19.215 //y=5.02
c67 ( 26 0 ) capacitor c=0.0084702f //x=20.09 //y=0.905
c68 ( 25 0 ) capacitor c=0.00427536f //x=20.24 //y=5.2
c69 ( 24 0 ) capacitor c=0.132738f //x=20.72 //y=5.115
c70 ( 22 0 ) capacitor c=0.00781917f //x=20.365 //y=1.655
c71 ( 21 0 ) capacitor c=0.0167625f //x=20.635 //y=1.655
c72 ( 19 0 ) capacitor c=0.0162757f //x=20.635 //y=5.2
c73 ( 8 0 ) capacitor c=0.00265417f //x=19.445 //y=5.2
c74 ( 7 0 ) capacitor c=0.0157611f //x=20.155 //y=5.2
r75 (  23 24 ) resistor r=231.016 //w=0.187 //l=3.375 //layer=li \
 //thickness=0.1 //x=20.72 //y=1.74 //x2=20.72 //y2=5.115
r76 (  21 23 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.635 //y=1.655 //x2=20.72 //y2=1.74
r77 (  21 22 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=20.635 //y=1.655 //x2=20.365 //y2=1.655
r78 (  20 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.325 //y=5.2 //x2=20.24 //y2=5.2
r79 (  19 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.635 //y=5.2 //x2=20.72 //y2=5.115
r80 (  19 20 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=20.635 //y=5.2 //x2=20.325 //y2=5.2
r81 (  15 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.28 //y=1.57 //x2=20.365 //y2=1.655
r82 (  15 26 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=20.28 //y=1.57 //x2=20.28 //y2=1
r83 (  9 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.24 //y=5.285 //x2=20.24 //y2=5.2
r84 (  9 29 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li //thickness=0.1 \
 //x=20.24 //y=5.285 //x2=20.24 //y2=5.725
r85 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.155 //y=5.2 //x2=20.24 //y2=5.2
r86 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=20.155 //y=5.2 //x2=19.445 //y2=5.2
r87 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=19.36 //y=5.285 //x2=19.445 //y2=5.2
r88 (  1 28 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li //thickness=0.1 \
 //x=19.36 //y=5.285 //x2=19.36 //y2=5.725
ends PM_DFFX1_PCELL\%noxref_18

subckt PM_DFFX1_PCELL\%noxref_19 ( 1 5 9 10 13 17 29 )
c47 ( 29 0 ) capacitor c=0.0644508f //x=18.69 //y=0.365
c48 ( 17 0 ) capacitor c=0.00722223f //x=20.765 //y=0.615
c49 ( 13 0 ) capacitor c=0.0154622f //x=20.68 //y=0.53
c50 ( 10 0 ) capacitor c=0.00708989f //x=19.795 //y=1.495
c51 ( 9 0 ) capacitor c=0.006761f //x=19.795 //y=0.615
c52 ( 5 0 ) capacitor c=0.0208654f //x=19.71 //y=1.58
c53 ( 1 0 ) capacitor c=0.00881098f //x=18.825 //y=1.495
r54 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=20.765 //y=0.615 //x2=20.765 //y2=0.49
r55 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=20.765 //y=0.615 //x2=20.765 //y2=0.88
r56 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.88 //y=0.53 //x2=19.795 //y2=0.49
r57 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.88 //y=0.53 //x2=20.28 //y2=0.53
r58 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.68 //y=0.53 //x2=20.765 //y2=0.49
r59 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.68 //y=0.53 //x2=20.28 //y2=0.53
r60 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=19.795 //y=1.495 //x2=19.795 //y2=1.62
r61 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=19.795 //y=1.495 //x2=19.795 //y2=0.88
r62 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=19.795 //y=0.615 //x2=19.795 //y2=0.49
r63 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=19.795 //y=0.615 //x2=19.795 //y2=0.88
r64 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.91 //y=1.58 //x2=18.825 //y2=1.62
r65 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.91 //y=1.58 //x2=19.31 //y2=1.58
r66 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.71 //y=1.58 //x2=19.795 //y2=1.62
r67 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.71 //y=1.58 //x2=19.31 //y2=1.58
r68 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=18.825 //y=1.495 //x2=18.825 //y2=1.62
r69 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=18.825 //y=1.495 //x2=18.825 //y2=0.88
ends PM_DFFX1_PCELL\%noxref_19

