* SPICE3 file created from BUFX1.ext - technology: sky130A

.subckt BUFX1 Y A VDD GND
X0 VDD a_185_182 Y VDD pshort w=2 l=0.15 M=2
X1 a_185_182 A GND GND nshort w=3 l=0.15
X2 VDD A a_185_182 VDD pshort w=2 l=0.15 M=2
X3 Y a_185_182 GND GND nshort w=3 l=0.15
C0 VDD GND 2.50fF
.ends
