// File: TMRDFFQNX1.spi.pex
// Created: Tue Oct 15 15:51:34 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_TMRDFFQNX1\%GND ( 1 123 127 130 135 145 153 161 167 173 181 189 197 \
 205 211 217 225 235 243 251 259 267 273 279 287 295 303 311 317 327 333 339 \
 347 355 363 371 377 383 391 399 407 415 421 427 440 444 446 449 451 453 456 \
 458 460 462 465 467 469 472 475 477 479 482 484 486 489 491 492 493 494 495 \
 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510 511 )
c936 ( 511 0 ) capacitor c=0.0215012f //x=72.03 //y=0.865
c937 ( 510 0 ) capacitor c=0.0215012f //x=68.7 //y=0.865
c938 ( 509 0 ) capacitor c=0.0207058f //x=65.37 //y=0.865
c939 ( 508 0 ) capacitor c=0.0207407f //x=62.04 //y=0.865
c940 ( 507 0 ) capacitor c=0.0207407f //x=58.71 //y=0.865
c941 ( 506 0 ) capacitor c=0.0207407f //x=55.38 //y=0.865
c942 ( 505 0 ) capacitor c=0.0207407f //x=52.05 //y=0.865
c943 ( 504 0 ) capacitor c=0.0207407f //x=48.72 //y=0.865
c944 ( 503 0 ) capacitor c=0.0226075f //x=43.805 //y=0.875
c945 ( 502 0 ) capacitor c=0.0207407f //x=40.58 //y=0.865
c946 ( 501 0 ) capacitor c=0.0207675f //x=37.25 //y=0.865
c947 ( 500 0 ) capacitor c=0.0207675f //x=33.92 //y=0.865
c948 ( 499 0 ) capacitor c=0.0207675f //x=30.59 //y=0.865
c949 ( 498 0 ) capacitor c=0.0207675f //x=27.26 //y=0.865
c950 ( 497 0 ) capacitor c=0.0226344f //x=22.345 //y=0.875
c951 ( 496 0 ) capacitor c=0.0207675f //x=19.12 //y=0.865
c952 ( 495 0 ) capacitor c=0.0207675f //x=15.79 //y=0.865
c953 ( 494 0 ) capacitor c=0.0207675f //x=12.46 //y=0.865
c954 ( 493 0 ) capacitor c=0.0207675f //x=9.13 //y=0.865
c955 ( 492 0 ) capacitor c=0.0208019f //x=5.8 //y=0.865
c956 ( 491 0 ) capacitor c=0.022675f //x=0.885 //y=0.875
c957 ( 490 0 ) capacitor c=0.00440095f //x=72.22 //y=0
c958 ( 489 0 ) capacitor c=0.101477f //x=71.04 //y=0
c959 ( 488 0 ) capacitor c=0.00440095f //x=68.82 //y=0
c960 ( 486 0 ) capacitor c=0.115716f //x=67.71 //y=0
c961 ( 485 0 ) capacitor c=0.00440095f //x=65.56 //y=0
c962 ( 484 0 ) capacitor c=0.10307f //x=64.38 //y=0
c963 ( 483 0 ) capacitor c=0.00440095f //x=62.23 //y=0
c964 ( 482 0 ) capacitor c=0.105373f //x=61.05 //y=0
c965 ( 481 0 ) capacitor c=0.00440095f //x=58.83 //y=0
c966 ( 479 0 ) capacitor c=0.105373f //x=57.72 //y=0
c967 ( 478 0 ) capacitor c=0.00440095f //x=55.57 //y=0
c968 ( 477 0 ) capacitor c=0.105373f //x=54.39 //y=0
c969 ( 476 0 ) capacitor c=0.00440095f //x=52.24 //y=0
c970 ( 475 0 ) capacitor c=0.104903f //x=51.06 //y=0
c971 ( 474 0 ) capacitor c=0.00440095f //x=48.84 //y=0
c972 ( 472 0 ) capacitor c=0.108614f //x=47.73 //y=0
c973 ( 471 0 ) capacitor c=0.00440144f //x=44.03 //y=0
c974 ( 469 0 ) capacitor c=0.104362f //x=42.92 //y=0
c975 ( 468 0 ) capacitor c=0.00440095f //x=40.77 //y=0
c976 ( 467 0 ) capacitor c=0.105632f //x=39.59 //y=0
c977 ( 466 0 ) capacitor c=0.00440095f //x=37.44 //y=0
c978 ( 465 0 ) capacitor c=0.106656f //x=36.26 //y=0
c979 ( 464 0 ) capacitor c=0.00440095f //x=34.04 //y=0
c980 ( 462 0 ) capacitor c=0.106969f //x=32.93 //y=0
c981 ( 461 0 ) capacitor c=0.00440095f //x=30.78 //y=0
c982 ( 460 0 ) capacitor c=0.106848f //x=29.6 //y=0
c983 ( 459 0 ) capacitor c=0.00440095f //x=27.45 //y=0
c984 ( 458 0 ) capacitor c=0.109784f //x=26.27 //y=0
c985 ( 457 0 ) capacitor c=0.00440144f //x=22.535 //y=0
c986 ( 456 0 ) capacitor c=0.10575f //x=21.46 //y=0
c987 ( 455 0 ) capacitor c=0.00440095f //x=19.24 //y=0
c988 ( 453 0 ) capacitor c=0.106969f //x=18.13 //y=0
c989 ( 452 0 ) capacitor c=0.00440095f //x=15.98 //y=0
c990 ( 451 0 ) capacitor c=0.106969f //x=14.8 //y=0
c991 ( 450 0 ) capacitor c=0.00440095f //x=12.65 //y=0
c992 ( 449 0 ) capacitor c=0.106969f //x=11.47 //y=0
c993 ( 448 0 ) capacitor c=0.00440095f //x=9.25 //y=0
c994 ( 446 0 ) capacitor c=0.106848f //x=8.14 //y=0
c995 ( 445 0 ) capacitor c=0.00440095f //x=5.99 //y=0
c996 ( 444 0 ) capacitor c=0.109537f //x=4.81 //y=0
c997 ( 443 0 ) capacitor c=0.00440144f //x=1.075 //y=0
c998 ( 440 0 ) capacitor c=0.258637f //x=73.63 //y=0
c999 ( 427 0 ) capacitor c=0.0389876f //x=72.135 //y=0
c1000 ( 421 0 ) capacitor c=0.0716428f //x=70.87 //y=0
c1001 ( 415 0 ) capacitor c=0.0388276f //x=68.805 //y=0
c1002 ( 407 0 ) capacitor c=0.0717268f //x=67.54 //y=0
c1003 ( 399 0 ) capacitor c=0.039094f //x=65.475 //y=0
c1004 ( 391 0 ) capacitor c=0.0718026f //x=64.21 //y=0
c1005 ( 383 0 ) capacitor c=0.0388888f //x=62.145 //y=0
c1006 ( 377 0 ) capacitor c=0.0718026f //x=60.88 //y=0
c1007 ( 371 0 ) capacitor c=0.0388888f //x=58.815 //y=0
c1008 ( 363 0 ) capacitor c=0.0718026f //x=57.55 //y=0
c1009 ( 355 0 ) capacitor c=0.0388888f //x=55.485 //y=0
c1010 ( 347 0 ) capacitor c=0.0718026f //x=54.22 //y=0
c1011 ( 339 0 ) capacitor c=0.0388888f //x=52.155 //y=0
c1012 ( 333 0 ) capacitor c=0.0718026f //x=50.89 //y=0
c1013 ( 327 0 ) capacitor c=0.0388888f //x=48.825 //y=0
c1014 ( 317 0 ) capacitor c=0.133362f //x=47.56 //y=0
c1015 ( 311 0 ) capacitor c=0.0339325f //x=43.91 //y=0
c1016 ( 303 0 ) capacitor c=0.0718011f //x=42.75 //y=0
c1017 ( 295 0 ) capacitor c=0.0388888f //x=40.685 //y=0
c1018 ( 287 0 ) capacitor c=0.0718137f //x=39.42 //y=0
c1019 ( 279 0 ) capacitor c=0.0389039f //x=37.355 //y=0
c1020 ( 273 0 ) capacitor c=0.0718422f //x=36.09 //y=0
c1021 ( 267 0 ) capacitor c=0.0389039f //x=34.025 //y=0
c1022 ( 259 0 ) capacitor c=0.0718422f //x=32.76 //y=0
c1023 ( 251 0 ) capacitor c=0.0389039f //x=30.695 //y=0
c1024 ( 243 0 ) capacitor c=0.0718417f //x=29.43 //y=0
c1025 ( 235 0 ) capacitor c=0.0389039f //x=27.365 //y=0
c1026 ( 225 0 ) capacitor c=0.133515f //x=26.1 //y=0
c1027 ( 217 0 ) capacitor c=0.0339482f //x=22.45 //y=0
c1028 ( 211 0 ) capacitor c=0.0718422f //x=21.29 //y=0
c1029 ( 205 0 ) capacitor c=0.0389039f //x=19.225 //y=0
c1030 ( 197 0 ) capacitor c=0.0718422f //x=17.96 //y=0
c1031 ( 189 0 ) capacitor c=0.0389039f //x=15.895 //y=0
c1032 ( 181 0 ) capacitor c=0.0718422f //x=14.63 //y=0
c1033 ( 173 0 ) capacitor c=0.0389039f //x=12.565 //y=0
c1034 ( 167 0 ) capacitor c=0.0718422f //x=11.3 //y=0
c1035 ( 161 0 ) capacitor c=0.0389039f //x=9.235 //y=0
c1036 ( 153 0 ) capacitor c=0.0718609f //x=7.97 //y=0
c1037 ( 145 0 ) capacitor c=0.0389288f //x=5.905 //y=0
c1038 ( 135 0 ) capacitor c=0.131745f //x=4.64 //y=0
c1039 ( 130 0 ) capacitor c=0.178285f //x=0.74 //y=0
c1040 ( 127 0 ) capacitor c=0.0367385f //x=0.99 //y=0
c1041 ( 123 0 ) capacitor c=2.29191f //x=73.63 //y=0
r1042 (  438 440 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=72.52 //y=0 //x2=73.63 //y2=0
r1043 (  436 490 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.305 //y=0 //x2=72.22 //y2=0
r1044 (  436 438 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=72.305 //y=0 //x2=72.52 //y2=0
r1045 (  431 490 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=72.22 //y=0.17 //x2=72.22 //y2=0
r1046 (  431 511 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=72.22 //y=0.17 //x2=72.22 //y2=0.955
r1047 (  428 489 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=71.21 //y=0 //x2=71.04 //y2=0
r1048 (  428 430 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=71.21 //y=0 //x2=71.41 //y2=0
r1049 (  427 490 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.135 //y=0 //x2=72.22 //y2=0
r1050 (  427 430 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=72.135 //y=0 //x2=71.41 //y2=0
r1051 (  422 488 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.975 //y=0 //x2=68.89 //y2=0
r1052 (  422 424 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=68.975 //y=0 //x2=69.93 //y2=0
r1053 (  421 489 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=70.87 //y=0 //x2=71.04 //y2=0
r1054 (  421 424 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=70.87 //y=0 //x2=69.93 //y2=0
r1055 (  417 488 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.89 //y=0.17 //x2=68.89 //y2=0
r1056 (  417 510 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=68.89 //y=0.17 //x2=68.89 //y2=0.955
r1057 (  416 486 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.88 //y=0 //x2=67.71 //y2=0
r1058 (  415 488 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.805 //y=0 //x2=68.89 //y2=0
r1059 (  415 416 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=68.805 //y=0 //x2=67.88 //y2=0
r1060 (  410 412 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=66.23 //y=0 //x2=67.34 //y2=0
r1061 (  408 485 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.645 //y=0 //x2=65.56 //y2=0
r1062 (  408 410 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=65.645 //y=0 //x2=66.23 //y2=0
r1063 (  407 486 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.54 //y=0 //x2=67.71 //y2=0
r1064 (  407 412 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=67.54 //y=0 //x2=67.34 //y2=0
r1065 (  403 485 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=65.56 //y=0.17 //x2=65.56 //y2=0
r1066 (  403 509 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=65.56 //y=0.17 //x2=65.56 //y2=0.955
r1067 (  400 484 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.55 //y=0 //x2=64.38 //y2=0
r1068 (  400 402 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=64.55 //y=0 //x2=65.12 //y2=0
r1069 (  399 485 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.475 //y=0 //x2=65.56 //y2=0
r1070 (  399 402 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=65.475 //y=0 //x2=65.12 //y2=0
r1071 (  394 396 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=62.53 //y=0 //x2=63.64 //y2=0
r1072 (  392 483 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.315 //y=0 //x2=62.23 //y2=0
r1073 (  392 394 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=62.315 //y=0 //x2=62.53 //y2=0
r1074 (  391 484 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.21 //y=0 //x2=64.38 //y2=0
r1075 (  391 396 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=64.21 //y=0 //x2=63.64 //y2=0
r1076 (  387 483 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.23 //y=0.17 //x2=62.23 //y2=0
r1077 (  387 508 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=62.23 //y=0.17 //x2=62.23 //y2=0.955
r1078 (  384 482 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.22 //y=0 //x2=61.05 //y2=0
r1079 (  384 386 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=61.22 //y=0 //x2=61.42 //y2=0
r1080 (  383 483 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.145 //y=0 //x2=62.23 //y2=0
r1081 (  383 386 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=62.145 //y=0 //x2=61.42 //y2=0
r1082 (  378 481 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.985 //y=0 //x2=58.9 //y2=0
r1083 (  378 380 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=58.985 //y=0 //x2=59.94 //y2=0
r1084 (  377 482 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=60.88 //y=0 //x2=61.05 //y2=0
r1085 (  377 380 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=60.88 //y=0 //x2=59.94 //y2=0
r1086 (  373 481 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.9 //y=0.17 //x2=58.9 //y2=0
r1087 (  373 507 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=58.9 //y=0.17 //x2=58.9 //y2=0.955
r1088 (  372 479 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.89 //y=0 //x2=57.72 //y2=0
r1089 (  371 481 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.815 //y=0 //x2=58.9 //y2=0
r1090 (  371 372 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=58.815 //y=0 //x2=57.89 //y2=0
r1091 (  366 368 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=56.24 //y=0 //x2=57.35 //y2=0
r1092 (  364 478 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.655 //y=0 //x2=55.57 //y2=0
r1093 (  364 366 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=55.655 //y=0 //x2=56.24 //y2=0
r1094 (  363 479 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.55 //y=0 //x2=57.72 //y2=0
r1095 (  363 368 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=57.55 //y=0 //x2=57.35 //y2=0
r1096 (  359 478 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=55.57 //y=0.17 //x2=55.57 //y2=0
r1097 (  359 506 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=55.57 //y=0.17 //x2=55.57 //y2=0.955
r1098 (  356 477 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=54.56 //y=0 //x2=54.39 //y2=0
r1099 (  356 358 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=54.56 //y=0 //x2=55.13 //y2=0
r1100 (  355 478 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.485 //y=0 //x2=55.57 //y2=0
r1101 (  355 358 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=55.485 //y=0 //x2=55.13 //y2=0
r1102 (  350 352 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=52.54 //y=0 //x2=53.65 //y2=0
r1103 (  348 476 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=52.325 //y=0 //x2=52.24 //y2=0
r1104 (  348 350 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=52.325 //y=0 //x2=52.54 //y2=0
r1105 (  347 477 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=54.22 //y=0 //x2=54.39 //y2=0
r1106 (  347 352 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=54.22 //y=0 //x2=53.65 //y2=0
r1107 (  343 476 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=52.24 //y=0.17 //x2=52.24 //y2=0
r1108 (  343 505 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=52.24 //y=0.17 //x2=52.24 //y2=0.955
r1109 (  340 475 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=51.23 //y=0 //x2=51.06 //y2=0
r1110 (  340 342 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=51.23 //y=0 //x2=51.43 //y2=0
r1111 (  339 476 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=52.155 //y=0 //x2=52.24 //y2=0
r1112 (  339 342 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=52.155 //y=0 //x2=51.43 //y2=0
r1113 (  334 474 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=48.995 //y=0 //x2=48.91 //y2=0
r1114 (  334 336 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=48.995 //y=0 //x2=49.95 //y2=0
r1115 (  333 475 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=50.89 //y=0 //x2=51.06 //y2=0
r1116 (  333 336 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=50.89 //y=0 //x2=49.95 //y2=0
r1117 (  329 474 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.91 //y=0.17 //x2=48.91 //y2=0
r1118 (  329 504 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=48.91 //y=0.17 //x2=48.91 //y2=0.955
r1119 (  328 472 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.9 //y=0 //x2=47.73 //y2=0
r1120 (  327 474 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=48.825 //y=0 //x2=48.91 //y2=0
r1121 (  327 328 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=48.825 //y=0 //x2=47.9 //y2=0
r1122 (  322 324 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=46.25 //y=0 //x2=47.36 //y2=0
r1123 (  320 322 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=45.14 //y=0 //x2=46.25 //y2=0
r1124 (  318 471 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.08 //y=0 //x2=43.995 //y2=0
r1125 (  318 320 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=44.08 //y=0 //x2=45.14 //y2=0
r1126 (  317 472 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.56 //y=0 //x2=47.73 //y2=0
r1127 (  317 324 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=47.56 //y=0 //x2=47.36 //y2=0
r1128 (  313 471 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.995 //y=0.17 //x2=43.995 //y2=0
r1129 (  313 503 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=43.995 //y=0.17 //x2=43.995 //y2=0.965
r1130 (  312 469 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.09 //y=0 //x2=42.92 //y2=0
r1131 (  311 471 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=43.91 //y=0 //x2=43.995 //y2=0
r1132 (  311 312 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=43.91 //y=0 //x2=43.09 //y2=0
r1133 (  306 308 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=41.44 //y=0 //x2=42.55 //y2=0
r1134 (  304 468 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.855 //y=0 //x2=40.77 //y2=0
r1135 (  304 306 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=40.855 //y=0 //x2=41.44 //y2=0
r1136 (  303 469 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=42.75 //y=0 //x2=42.92 //y2=0
r1137 (  303 308 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=42.75 //y=0 //x2=42.55 //y2=0
r1138 (  299 468 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.77 //y=0.17 //x2=40.77 //y2=0
r1139 (  299 502 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=40.77 //y=0.17 //x2=40.77 //y2=0.955
r1140 (  296 467 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.76 //y=0 //x2=39.59 //y2=0
r1141 (  296 298 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=39.76 //y=0 //x2=40.33 //y2=0
r1142 (  295 468 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.685 //y=0 //x2=40.77 //y2=0
r1143 (  295 298 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=40.685 //y=0 //x2=40.33 //y2=0
r1144 (  290 292 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=37.74 //y=0 //x2=38.85 //y2=0
r1145 (  288 466 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.525 //y=0 //x2=37.44 //y2=0
r1146 (  288 290 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=37.525 //y=0 //x2=37.74 //y2=0
r1147 (  287 467 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.42 //y=0 //x2=39.59 //y2=0
r1148 (  287 292 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=39.42 //y=0 //x2=38.85 //y2=0
r1149 (  283 466 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.44 //y=0.17 //x2=37.44 //y2=0
r1150 (  283 501 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=37.44 //y=0.17 //x2=37.44 //y2=0.955
r1151 (  280 465 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.43 //y=0 //x2=36.26 //y2=0
r1152 (  280 282 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=36.43 //y=0 //x2=36.63 //y2=0
r1153 (  279 466 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.355 //y=0 //x2=37.44 //y2=0
r1154 (  279 282 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=37.355 //y=0 //x2=36.63 //y2=0
r1155 (  274 464 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.195 //y=0 //x2=34.11 //y2=0
r1156 (  274 276 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=34.195 //y=0 //x2=35.15 //y2=0
r1157 (  273 465 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.09 //y=0 //x2=36.26 //y2=0
r1158 (  273 276 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=36.09 //y=0 //x2=35.15 //y2=0
r1159 (  269 464 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=34.11 //y=0.17 //x2=34.11 //y2=0
r1160 (  269 500 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=34.11 //y=0.17 //x2=34.11 //y2=0.955
r1161 (  268 462 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.1 //y=0 //x2=32.93 //y2=0
r1162 (  267 464 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.025 //y=0 //x2=34.11 //y2=0
r1163 (  267 268 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=34.025 //y=0 //x2=33.1 //y2=0
r1164 (  262 264 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=31.45 //y=0 //x2=32.56 //y2=0
r1165 (  260 461 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.865 //y=0 //x2=30.78 //y2=0
r1166 (  260 262 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=30.865 //y=0 //x2=31.45 //y2=0
r1167 (  259 462 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.76 //y=0 //x2=32.93 //y2=0
r1168 (  259 264 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=32.76 //y=0 //x2=32.56 //y2=0
r1169 (  255 461 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.78 //y=0.17 //x2=30.78 //y2=0
r1170 (  255 499 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=30.78 //y=0.17 //x2=30.78 //y2=0.955
r1171 (  252 460 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.77 //y=0 //x2=29.6 //y2=0
r1172 (  252 254 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=29.77 //y=0 //x2=30.34 //y2=0
r1173 (  251 461 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.695 //y=0 //x2=30.78 //y2=0
r1174 (  251 254 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=30.695 //y=0 //x2=30.34 //y2=0
r1175 (  246 248 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=27.75 //y=0 //x2=28.86 //y2=0
r1176 (  244 459 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.535 //y=0 //x2=27.45 //y2=0
r1177 (  244 246 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=27.535 //y=0 //x2=27.75 //y2=0
r1178 (  243 460 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.43 //y=0 //x2=29.6 //y2=0
r1179 (  243 248 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=29.43 //y=0 //x2=28.86 //y2=0
r1180 (  239 459 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.45 //y=0.17 //x2=27.45 //y2=0
r1181 (  239 498 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=27.45 //y=0.17 //x2=27.45 //y2=0.955
r1182 (  236 458 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.44 //y=0 //x2=26.27 //y2=0
r1183 (  236 238 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=26.44 //y=0 //x2=26.64 //y2=0
r1184 (  235 459 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.365 //y=0 //x2=27.45 //y2=0
r1185 (  235 238 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=27.365 //y=0 //x2=26.64 //y2=0
r1186 (  230 232 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=24.05 //y=0 //x2=25.16 //y2=0
r1187 (  228 230 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=22.94 //y=0 //x2=24.05 //y2=0
r1188 (  226 457 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.62 //y=0 //x2=22.535 //y2=0
r1189 (  226 228 ) resistor r=11.4734 //w=0.357 //l=0.32 //layer=li \
 //thickness=0.1 //x=22.62 //y=0 //x2=22.94 //y2=0
r1190 (  225 458 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.1 //y=0 //x2=26.27 //y2=0
r1191 (  225 232 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=26.1 //y=0 //x2=25.16 //y2=0
r1192 (  221 457 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.535 //y=0.17 //x2=22.535 //y2=0
r1193 (  221 497 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=22.535 //y=0.17 //x2=22.535 //y2=0.965
r1194 (  218 456 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.63 //y=0 //x2=21.46 //y2=0
r1195 (  218 220 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=21.63 //y=0 //x2=21.83 //y2=0
r1196 (  217 457 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.45 //y=0 //x2=22.535 //y2=0
r1197 (  217 220 ) resistor r=22.2297 //w=0.357 //l=0.62 //layer=li \
 //thickness=0.1 //x=22.45 //y=0 //x2=21.83 //y2=0
r1198 (  212 455 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.395 //y=0 //x2=19.31 //y2=0
r1199 (  212 214 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=19.395 //y=0 //x2=20.35 //y2=0
r1200 (  211 456 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.29 //y=0 //x2=21.46 //y2=0
r1201 (  211 214 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=21.29 //y=0 //x2=20.35 //y2=0
r1202 (  207 455 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.31 //y=0.17 //x2=19.31 //y2=0
r1203 (  207 496 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=19.31 //y=0.17 //x2=19.31 //y2=0.955
r1204 (  206 453 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.3 //y=0 //x2=18.13 //y2=0
r1205 (  205 455 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.225 //y=0 //x2=19.31 //y2=0
r1206 (  205 206 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=19.225 //y=0 //x2=18.3 //y2=0
r1207 (  200 202 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=16.65 //y=0 //x2=17.76 //y2=0
r1208 (  198 452 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.065 //y=0 //x2=15.98 //y2=0
r1209 (  198 200 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=16.065 //y=0 //x2=16.65 //y2=0
r1210 (  197 453 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.96 //y=0 //x2=18.13 //y2=0
r1211 (  197 202 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=17.96 //y=0 //x2=17.76 //y2=0
r1212 (  193 452 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.98 //y=0.17 //x2=15.98 //y2=0
r1213 (  193 495 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=15.98 //y=0.17 //x2=15.98 //y2=0.955
r1214 (  190 451 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.97 //y=0 //x2=14.8 //y2=0
r1215 (  190 192 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.97 //y=0 //x2=15.54 //y2=0
r1216 (  189 452 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.895 //y=0 //x2=15.98 //y2=0
r1217 (  189 192 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=15.895 //y=0 //x2=15.54 //y2=0
r1218 (  184 186 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=12.95 //y=0 //x2=14.06 //y2=0
r1219 (  182 450 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.735 //y=0 //x2=12.65 //y2=0
r1220 (  182 184 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=12.735 //y=0 //x2=12.95 //y2=0
r1221 (  181 451 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.63 //y=0 //x2=14.8 //y2=0
r1222 (  181 186 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.63 //y=0 //x2=14.06 //y2=0
r1223 (  177 450 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.65 //y=0.17 //x2=12.65 //y2=0
r1224 (  177 494 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=12.65 //y=0.17 //x2=12.65 //y2=0.955
r1225 (  174 449 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.64 //y=0 //x2=11.47 //y2=0
r1226 (  174 176 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=11.64 //y=0 //x2=11.84 //y2=0
r1227 (  173 450 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.565 //y=0 //x2=12.65 //y2=0
r1228 (  173 176 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=12.565 //y=0 //x2=11.84 //y2=0
r1229 (  168 448 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.405 //y=0 //x2=9.32 //y2=0
r1230 (  168 170 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=9.405 //y=0 //x2=10.36 //y2=0
r1231 (  167 449 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.3 //y=0 //x2=11.47 //y2=0
r1232 (  167 170 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=11.3 //y=0 //x2=10.36 //y2=0
r1233 (  163 448 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.32 //y=0.17 //x2=9.32 //y2=0
r1234 (  163 493 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=9.32 //y=0.17 //x2=9.32 //y2=0.955
r1235 (  162 446 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=0 //x2=8.14 //y2=0
r1236 (  161 448 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.235 //y=0 //x2=9.32 //y2=0
r1237 (  161 162 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=9.235 //y=0 //x2=8.31 //y2=0
r1238 (  156 158 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r1239 (  154 445 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.075 //y=0 //x2=5.99 //y2=0
r1240 (  154 156 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=6.075 //y=0 //x2=6.66 //y2=0
r1241 (  153 446 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=8.14 //y2=0
r1242 (  153 158 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=7.77 //y2=0
r1243 (  149 445 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.99 //y=0.17 //x2=5.99 //y2=0
r1244 (  149 492 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=5.99 //y=0.17 //x2=5.99 //y2=0.955
r1245 (  146 444 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=4.81 //y2=0
r1246 (  146 148 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=5.55 //y2=0
r1247 (  145 445 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.905 //y=0 //x2=5.99 //y2=0
r1248 (  145 148 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=5.905 //y=0 //x2=5.55 //y2=0
r1249 (  140 142 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=0 //x2=4.07 //y2=0
r1250 (  138 140 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r1251 (  136 443 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.075 //y2=0
r1252 (  136 138 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.85 //y2=0
r1253 (  135 444 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.81 //y2=0
r1254 (  135 142 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.07 //y2=0
r1255 (  131 443 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0
r1256 (  131 491 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0.965
r1257 (  127 443 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=1.075 //y2=0
r1258 (  127 130 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=0.74 //y2=0
r1259 (  123 440 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=73.63 //y=0 //x2=73.63 //y2=0
r1260 (  121 438 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=72.52 //y=0 //x2=72.52 //y2=0
r1261 (  121 123 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=72.52 //y=0 //x2=73.63 //y2=0
r1262 (  119 430 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=71.41 //y=0 //x2=71.41 //y2=0
r1263 (  119 121 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=71.41 //y=0 //x2=72.52 //y2=0
r1264 (  117 424 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=69.93 //y=0 //x2=69.93 //y2=0
r1265 (  117 119 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=69.93 //y=0 //x2=71.41 //y2=0
r1266 (  115 488 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=68.82 //y=0 //x2=68.82 //y2=0
r1267 (  115 117 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=68.82 //y=0 //x2=69.93 //y2=0
r1268 (  113 412 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=67.34 //y=0 //x2=67.34 //y2=0
r1269 (  113 115 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=67.34 //y=0 //x2=68.82 //y2=0
r1270 (  111 410 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=66.23 //y=0 //x2=66.23 //y2=0
r1271 (  111 113 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=66.23 //y=0 //x2=67.34 //y2=0
r1272 (  109 402 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=65.12 //y=0 //x2=65.12 //y2=0
r1273 (  109 111 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=65.12 //y=0 //x2=66.23 //y2=0
r1274 (  107 396 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=63.64 //y=0 //x2=63.64 //y2=0
r1275 (  107 109 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=63.64 //y=0 //x2=65.12 //y2=0
r1276 (  105 394 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=62.53 //y=0 //x2=62.53 //y2=0
r1277 (  105 107 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=62.53 //y=0 //x2=63.64 //y2=0
r1278 (  103 386 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=61.42 //y=0 //x2=61.42 //y2=0
r1279 (  103 105 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=61.42 //y=0 //x2=62.53 //y2=0
r1280 (  101 380 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=59.94 //y=0 //x2=59.94 //y2=0
r1281 (  101 103 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=59.94 //y=0 //x2=61.42 //y2=0
r1282 (  99 481 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=58.83 //y=0 //x2=58.83 //y2=0
r1283 (  99 101 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=58.83 //y=0 //x2=59.94 //y2=0
r1284 (  97 368 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=57.35 //y=0 //x2=57.35 //y2=0
r1285 (  97 99 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=57.35 //y=0 //x2=58.83 //y2=0
r1286 (  95 366 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=56.24 //y=0 //x2=56.24 //y2=0
r1287 (  95 97 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=56.24 //y=0 //x2=57.35 //y2=0
r1288 (  93 358 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=55.13 //y=0 //x2=55.13 //y2=0
r1289 (  93 95 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=55.13 //y=0 //x2=56.24 //y2=0
r1290 (  91 352 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=53.65 //y=0 //x2=53.65 //y2=0
r1291 (  91 93 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=53.65 //y=0 //x2=55.13 //y2=0
r1292 (  89 350 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=52.54 //y=0 //x2=52.54 //y2=0
r1293 (  89 91 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=52.54 //y=0 //x2=53.65 //y2=0
r1294 (  87 342 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=51.43 //y=0 //x2=51.43 //y2=0
r1295 (  87 89 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=51.43 //y=0 //x2=52.54 //y2=0
r1296 (  85 336 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=49.95 //y=0 //x2=49.95 //y2=0
r1297 (  85 87 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=49.95 //y=0 //x2=51.43 //y2=0
r1298 (  83 474 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=48.84 //y=0 //x2=48.84 //y2=0
r1299 (  83 85 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=48.84 //y=0 //x2=49.95 //y2=0
r1300 (  81 324 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=47.36 //y=0 //x2=47.36 //y2=0
r1301 (  81 83 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=47.36 //y=0 //x2=48.84 //y2=0
r1302 (  79 322 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=46.25 //y=0 //x2=46.25 //y2=0
r1303 (  79 81 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=46.25 //y=0 //x2=47.36 //y2=0
r1304 (  77 320 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=45.14 //y=0 //x2=45.14 //y2=0
r1305 (  77 79 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=45.14 //y=0 //x2=46.25 //y2=0
r1306 (  75 471 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=44.03 //y=0 //x2=44.03 //y2=0
r1307 (  75 77 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=44.03 //y=0 //x2=45.14 //y2=0
r1308 (  73 308 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=42.55 //y=0 //x2=42.55 //y2=0
r1309 (  73 75 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=42.55 //y=0 //x2=44.03 //y2=0
r1310 (  71 306 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=41.44 //y=0 //x2=41.44 //y2=0
r1311 (  71 73 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=41.44 //y=0 //x2=42.55 //y2=0
r1312 (  69 298 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=40.33 //y=0 //x2=40.33 //y2=0
r1313 (  69 71 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=40.33 //y=0 //x2=41.44 //y2=0
r1314 (  67 292 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=38.85 //y=0 //x2=38.85 //y2=0
r1315 (  67 69 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=38.85 //y=0 //x2=40.33 //y2=0
r1316 (  65 290 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37.74 //y=0 //x2=37.74 //y2=0
r1317 (  65 67 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=37.74 //y=0 //x2=38.85 //y2=0
r1318 (  62 282 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=36.63 //y=0 //x2=36.63 //y2=0
r1319 (  60 276 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.15 //y=0 //x2=35.15 //y2=0
r1320 (  60 62 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=35.15 //y=0 //x2=36.63 //y2=0
r1321 (  58 464 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.04 //y=0 //x2=34.04 //y2=0
r1322 (  58 60 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=34.04 //y=0 //x2=35.15 //y2=0
r1323 (  56 264 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.56 //y=0 //x2=32.56 //y2=0
r1324 (  56 58 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=32.56 //y=0 //x2=34.04 //y2=0
r1325 (  54 262 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.45 //y=0 //x2=31.45 //y2=0
r1326 (  54 56 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.45 //y=0 //x2=32.56 //y2=0
r1327 (  52 254 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=30.34 //y=0 //x2=30.34 //y2=0
r1328 (  52 54 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=30.34 //y=0 //x2=31.45 //y2=0
r1329 (  50 248 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.86 //y=0 //x2=28.86 //y2=0
r1330 (  50 52 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=28.86 //y=0 //x2=30.34 //y2=0
r1331 (  48 246 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.75 //y=0 //x2=27.75 //y2=0
r1332 (  48 50 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=27.75 //y=0 //x2=28.86 //y2=0
r1333 (  46 238 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=26.64 //y=0 //x2=26.64 //y2=0
r1334 (  46 48 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=26.64 //y=0 //x2=27.75 //y2=0
r1335 (  44 232 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.16 //y=0 //x2=25.16 //y2=0
r1336 (  44 46 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=25.16 //y=0 //x2=26.64 //y2=0
r1337 (  42 230 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.05 //y=0 //x2=24.05 //y2=0
r1338 (  42 44 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=24.05 //y=0 //x2=25.16 //y2=0
r1339 (  40 228 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.94 //y=0 //x2=22.94 //y2=0
r1340 (  40 42 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.94 //y=0 //x2=24.05 //y2=0
r1341 (  38 220 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.83 //y=0 //x2=21.83 //y2=0
r1342 (  38 40 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.83 //y=0 //x2=22.94 //y2=0
r1343 (  36 214 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=0 //x2=20.35 //y2=0
r1344 (  36 38 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=0 //x2=21.83 //y2=0
r1345 (  34 455 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.24 //y=0 //x2=19.24 //y2=0
r1346 (  34 36 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.24 //y=0 //x2=20.35 //y2=0
r1347 (  32 202 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=0 //x2=17.76 //y2=0
r1348 (  32 34 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=0 //x2=19.24 //y2=0
r1349 (  30 200 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=0 //x2=16.65 //y2=0
r1350 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=0 //x2=17.76 //y2=0
r1351 (  28 192 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.54 //y=0 //x2=15.54 //y2=0
r1352 (  28 30 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.54 //y=0 //x2=16.65 //y2=0
r1353 (  26 186 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=0 //x2=14.06 //y2=0
r1354 (  26 28 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=0 //x2=15.54 //y2=0
r1355 (  24 184 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.95 //y=0 //x2=12.95 //y2=0
r1356 (  24 26 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.95 //y=0 //x2=14.06 //y2=0
r1357 (  22 176 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.84 //y=0 //x2=11.84 //y2=0
r1358 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.84 //y=0 //x2=12.95 //y2=0
r1359 (  20 170 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r1360 (  20 22 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=0 //x2=11.84 //y2=0
r1361 (  18 448 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=0 //x2=9.25 //y2=0
r1362 (  18 20 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=0 //x2=10.36 //y2=0
r1363 (  16 158 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r1364 (  16 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=9.25 //y2=0
r1365 (  14 156 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r1366 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r1367 (  12 148 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r1368 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r1369 (  10 142 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r1370 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=0 //x2=5.55 //y2=0
r1371 (  8 140 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r1372 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.07 //y2=0
r1373 (  6 138 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r1374 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r1375 (  3 130 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r1376 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r1377 (  1 65 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=37.185 //y=0 //x2=37.74 //y2=0
r1378 (  1 62 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=37.185 //y=0 //x2=36.63 //y2=0
ends PM_TMRDFFQNX1\%GND

subckt PM_TMRDFFQNX1\%VDD ( 1 123 130 137 147 155 165 171 179 187 197 203 211 \
 221 231 235 245 255 263 267 275 283 293 299 307 317 327 331 341 351 361 369 \
 373 383 393 401 405 413 421 431 437 445 455 465 469 479 489 497 501 509 517 \
 527 533 541 549 559 569 575 583 593 603 607 617 627 635 639 647 655 665 671 \
 679 689 699 703 713 723 735 743 751 761 767 782 789 794 798 803 808 812 818 \
 823 828 832 837 842 848 852 857 862 866 871 876 877 878 879 880 881 882 883 \
 884 885 886 887 888 889 890 891 892 893 894 895 896 897 898 899 900 901 902 \
 903 904 905 906 907 908 909 910 911 912 913 914 915 916 917 918 919 920 921 \
 922 923 924 925 926 927 928 929 930 931 932 933 934 935 936 937 )
c998 ( 937 0 ) capacitor c=0.0476806f //x=66.785 //y=5.025
c999 ( 936 0 ) capacitor c=0.0241714f //x=65.905 //y=5.025
c1000 ( 935 0 ) capacitor c=0.0467094f //x=65.035 //y=5.025
c1001 ( 934 0 ) capacitor c=0.0382077f //x=63.455 //y=5.02
c1002 ( 933 0 ) capacitor c=0.0240874f //x=62.575 //y=5.02
c1003 ( 932 0 ) capacitor c=0.0490303f //x=61.705 //y=5.02
c1004 ( 931 0 ) capacitor c=0.0381674f //x=60.125 //y=5.02
c1005 ( 930 0 ) capacitor c=0.0240879f //x=59.245 //y=5.02
c1006 ( 929 0 ) capacitor c=0.0493657f //x=58.375 //y=5.02
c1007 ( 928 0 ) capacitor c=0.038145f //x=56.795 //y=5.02
c1008 ( 927 0 ) capacitor c=0.0240074f //x=55.915 //y=5.02
c1009 ( 926 0 ) capacitor c=0.0490303f //x=55.045 //y=5.02
c1010 ( 925 0 ) capacitor c=0.0380679f //x=53.465 //y=5.02
c1011 ( 924 0 ) capacitor c=0.024008f //x=52.585 //y=5.02
c1012 ( 923 0 ) capacitor c=0.0490303f //x=51.715 //y=5.02
c1013 ( 922 0 ) capacitor c=0.0380679f //x=50.135 //y=5.02
c1014 ( 921 0 ) capacitor c=0.024008f //x=49.255 //y=5.02
c1015 ( 920 0 ) capacitor c=0.049209f //x=48.385 //y=5.02
c1016 ( 919 0 ) capacitor c=0.0452179f //x=46.505 //y=5.02
c1017 ( 918 0 ) capacitor c=0.024152f //x=45.625 //y=5.02
c1018 ( 917 0 ) capacitor c=0.024152f //x=44.745 //y=5.02
c1019 ( 916 0 ) capacitor c=0.0531894f //x=43.875 //y=5.02
c1020 ( 915 0 ) capacitor c=0.0380679f //x=41.995 //y=5.02
c1021 ( 914 0 ) capacitor c=0.024008f //x=41.115 //y=5.02
c1022 ( 913 0 ) capacitor c=0.0490303f //x=40.245 //y=5.02
c1023 ( 912 0 ) capacitor c=0.0380679f //x=38.665 //y=5.02
c1024 ( 911 0 ) capacitor c=0.024008f //x=37.785 //y=5.02
c1025 ( 910 0 ) capacitor c=0.0490303f //x=36.915 //y=5.02
c1026 ( 909 0 ) capacitor c=0.0380679f //x=35.335 //y=5.02
c1027 ( 908 0 ) capacitor c=0.0240074f //x=34.455 //y=5.02
c1028 ( 907 0 ) capacitor c=0.0490303f //x=33.585 //y=5.02
c1029 ( 906 0 ) capacitor c=0.0380679f //x=32.005 //y=5.02
c1030 ( 905 0 ) capacitor c=0.024008f //x=31.125 //y=5.02
c1031 ( 904 0 ) capacitor c=0.0490303f //x=30.255 //y=5.02
c1032 ( 903 0 ) capacitor c=0.0380679f //x=28.675 //y=5.02
c1033 ( 902 0 ) capacitor c=0.024008f //x=27.795 //y=5.02
c1034 ( 901 0 ) capacitor c=0.049209f //x=26.925 //y=5.02
c1035 ( 900 0 ) capacitor c=0.0452179f //x=25.045 //y=5.02
c1036 ( 899 0 ) capacitor c=0.024152f //x=24.165 //y=5.02
c1037 ( 898 0 ) capacitor c=0.024152f //x=23.285 //y=5.02
c1038 ( 897 0 ) capacitor c=0.0531894f //x=22.415 //y=5.02
c1039 ( 896 0 ) capacitor c=0.0380679f //x=20.535 //y=5.02
c1040 ( 895 0 ) capacitor c=0.024008f //x=19.655 //y=5.02
c1041 ( 894 0 ) capacitor c=0.0490303f //x=18.785 //y=5.02
c1042 ( 893 0 ) capacitor c=0.0380679f //x=17.205 //y=5.02
c1043 ( 892 0 ) capacitor c=0.0240093f //x=16.325 //y=5.02
c1044 ( 891 0 ) capacitor c=0.0490349f //x=15.455 //y=5.02
c1045 ( 890 0 ) capacitor c=0.0380692f //x=13.875 //y=5.02
c1046 ( 889 0 ) capacitor c=0.0240074f //x=12.995 //y=5.02
c1047 ( 888 0 ) capacitor c=0.0490303f //x=12.125 //y=5.02
c1048 ( 887 0 ) capacitor c=0.0380679f //x=10.545 //y=5.02
c1049 ( 886 0 ) capacitor c=0.024008f //x=9.665 //y=5.02
c1050 ( 885 0 ) capacitor c=0.0490303f //x=8.795 //y=5.02
c1051 ( 884 0 ) capacitor c=0.0380679f //x=7.215 //y=5.02
c1052 ( 883 0 ) capacitor c=0.024008f //x=6.335 //y=5.02
c1053 ( 882 0 ) capacitor c=0.049209f //x=5.465 //y=5.02
c1054 ( 881 0 ) capacitor c=0.0452179f //x=3.585 //y=5.02
c1055 ( 880 0 ) capacitor c=0.024152f //x=2.705 //y=5.02
c1056 ( 879 0 ) capacitor c=0.02424f //x=1.825 //y=5.02
c1057 ( 878 0 ) capacitor c=0.0531407f //x=0.955 //y=5.02
c1058 ( 877 0 ) capacitor c=0.113329f //x=71.04 //y=7.4
c1059 ( 876 0 ) capacitor c=0.121198f //x=67.71 //y=7.4
c1060 ( 875 0 ) capacitor c=0.00591168f //x=66.93 //y=7.4
c1061 ( 874 0 ) capacitor c=0.00591168f //x=66.05 //y=7.4
c1062 ( 873 0 ) capacitor c=0.00591168f //x=65.12 //y=7.4
c1063 ( 871 0 ) capacitor c=0.115257f //x=64.38 //y=7.4
c1064 ( 870 0 ) capacitor c=0.00591168f //x=63.64 //y=7.4
c1065 ( 868 0 ) capacitor c=0.00591168f //x=62.72 //y=7.4
c1066 ( 867 0 ) capacitor c=0.00591168f //x=61.84 //y=7.4
c1067 ( 866 0 ) capacitor c=0.114092f //x=61.05 //y=7.4
c1068 ( 865 0 ) capacitor c=0.00591168f //x=60.27 //y=7.4
c1069 ( 864 0 ) capacitor c=0.00591168f //x=59.39 //y=7.4
c1070 ( 863 0 ) capacitor c=0.00591168f //x=58.51 //y=7.4
c1071 ( 862 0 ) capacitor c=0.115932f //x=57.72 //y=7.4
c1072 ( 861 0 ) capacitor c=0.00591168f //x=56.94 //y=7.4
c1073 ( 860 0 ) capacitor c=0.00591168f //x=56.06 //y=7.4
c1074 ( 859 0 ) capacitor c=0.00591168f //x=55.13 //y=7.4
c1075 ( 857 0 ) capacitor c=0.114361f //x=54.39 //y=7.4
c1076 ( 856 0 ) capacitor c=0.00591168f //x=53.65 //y=7.4
c1077 ( 854 0 ) capacitor c=0.00591168f //x=52.73 //y=7.4
c1078 ( 853 0 ) capacitor c=0.00591168f //x=51.85 //y=7.4
c1079 ( 852 0 ) capacitor c=0.11449f //x=51.06 //y=7.4
c1080 ( 851 0 ) capacitor c=0.00591168f //x=50.28 //y=7.4
c1081 ( 850 0 ) capacitor c=0.00591168f //x=49.4 //y=7.4
c1082 ( 849 0 ) capacitor c=0.00591168f //x=48.52 //y=7.4
c1083 ( 848 0 ) capacitor c=0.13457f //x=47.73 //y=7.4
c1084 ( 847 0 ) capacitor c=0.00591168f //x=46.65 //y=7.4
c1085 ( 846 0 ) capacitor c=0.00591168f //x=45.77 //y=7.4
c1086 ( 845 0 ) capacitor c=0.00591168f //x=44.89 //y=7.4
c1087 ( 844 0 ) capacitor c=0.00591168f //x=44.03 //y=7.4
c1088 ( 842 0 ) capacitor c=0.139223f //x=42.92 //y=7.4
c1089 ( 841 0 ) capacitor c=0.00591168f //x=42.14 //y=7.4
c1090 ( 840 0 ) capacitor c=0.00591168f //x=41.26 //y=7.4
c1091 ( 839 0 ) capacitor c=0.00591168f //x=40.33 //y=7.4
c1092 ( 837 0 ) capacitor c=0.11449f //x=39.59 //y=7.4
c1093 ( 836 0 ) capacitor c=0.00591168f //x=38.85 //y=7.4
c1094 ( 834 0 ) capacitor c=0.00591168f //x=37.93 //y=7.4
c1095 ( 833 0 ) capacitor c=0.00591168f //x=37.05 //y=7.4
c1096 ( 832 0 ) capacitor c=0.11432f //x=36.26 //y=7.4
c1097 ( 831 0 ) capacitor c=0.00591168f //x=35.48 //y=7.4
c1098 ( 830 0 ) capacitor c=0.00591168f //x=34.6 //y=7.4
c1099 ( 829 0 ) capacitor c=0.00591168f //x=33.72 //y=7.4
c1100 ( 828 0 ) capacitor c=0.114361f //x=32.93 //y=7.4
c1101 ( 827 0 ) capacitor c=0.00591168f //x=32.15 //y=7.4
c1102 ( 826 0 ) capacitor c=0.00591168f //x=31.27 //y=7.4
c1103 ( 825 0 ) capacitor c=0.00591168f //x=30.34 //y=7.4
c1104 ( 823 0 ) capacitor c=0.11449f //x=29.6 //y=7.4
c1105 ( 822 0 ) capacitor c=0.00591168f //x=28.86 //y=7.4
c1106 ( 820 0 ) capacitor c=0.00591168f //x=27.94 //y=7.4
c1107 ( 819 0 ) capacitor c=0.00591168f //x=27.06 //y=7.4
c1108 ( 818 0 ) capacitor c=0.13457f //x=26.27 //y=7.4
c1109 ( 817 0 ) capacitor c=0.00591168f //x=25.16 //y=7.4
c1110 ( 815 0 ) capacitor c=0.00591168f //x=24.31 //y=7.4
c1111 ( 814 0 ) capacitor c=0.00591168f //x=23.43 //y=7.4
c1112 ( 813 0 ) capacitor c=0.00591168f //x=22.55 //y=7.4
c1113 ( 812 0 ) capacitor c=0.139223f //x=21.46 //y=7.4
c1114 ( 811 0 ) capacitor c=0.00591168f //x=20.68 //y=7.4
c1115 ( 810 0 ) capacitor c=0.00591168f //x=19.8 //y=7.4
c1116 ( 809 0 ) capacitor c=0.00591168f //x=18.92 //y=7.4
c1117 ( 808 0 ) capacitor c=0.11449f //x=18.13 //y=7.4
c1118 ( 807 0 ) capacitor c=0.00591168f //x=17.35 //y=7.4
c1119 ( 806 0 ) capacitor c=0.00591168f //x=16.47 //y=7.4
c1120 ( 805 0 ) capacitor c=0.00591168f //x=15.54 //y=7.4
c1121 ( 803 0 ) capacitor c=0.114458f //x=14.8 //y=7.4
c1122 ( 802 0 ) capacitor c=0.00591168f //x=14.06 //y=7.4
c1123 ( 800 0 ) capacitor c=0.00591168f //x=13.14 //y=7.4
c1124 ( 799 0 ) capacitor c=0.00591168f //x=12.26 //y=7.4
c1125 ( 798 0 ) capacitor c=0.114361f //x=11.47 //y=7.4
c1126 ( 797 0 ) capacitor c=0.00591168f //x=10.69 //y=7.4
c1127 ( 796 0 ) capacitor c=0.00591168f //x=9.81 //y=7.4
c1128 ( 795 0 ) capacitor c=0.00591168f //x=8.93 //y=7.4
c1129 ( 794 0 ) capacitor c=0.11449f //x=8.14 //y=7.4
c1130 ( 793 0 ) capacitor c=0.00591168f //x=7.36 //y=7.4
c1131 ( 792 0 ) capacitor c=0.00591168f //x=6.48 //y=7.4
c1132 ( 791 0 ) capacitor c=0.00591168f //x=5.55 //y=7.4
c1133 ( 789 0 ) capacitor c=0.13457f //x=4.81 //y=7.4
c1134 ( 788 0 ) capacitor c=0.00591168f //x=3.73 //y=7.4
c1135 ( 787 0 ) capacitor c=0.00591168f //x=2.85 //y=7.4
c1136 ( 786 0 ) capacitor c=0.00591168f //x=1.97 //y=7.4
c1137 ( 785 0 ) capacitor c=0.00591168f //x=1.09 //y=7.4
c1138 ( 782 0 ) capacitor c=0.334471f //x=73.63 //y=7.4
c1139 ( 767 0 ) capacitor c=0.120978f //x=70.87 //y=7.4
c1140 ( 761 0 ) capacitor c=0.0236224f //x=67.54 //y=7.4
c1141 ( 751 0 ) capacitor c=0.028539f //x=66.845 //y=7.4
c1142 ( 743 0 ) capacitor c=0.0285075f //x=65.965 //y=7.4
c1143 ( 735 0 ) capacitor c=0.0275884f //x=65.085 //y=7.4
c1144 ( 731 0 ) capacitor c=0.0275781f //x=64.21 //y=7.4
c1145 ( 723 0 ) capacitor c=0.0284327f //x=63.515 //y=7.4
c1146 ( 713 0 ) capacitor c=0.0288431f //x=62.635 //y=7.4
c1147 ( 703 0 ) capacitor c=0.0240981f //x=61.755 //y=7.4
c1148 ( 699 0 ) capacitor c=0.0237088f //x=60.88 //y=7.4
c1149 ( 689 0 ) capacitor c=0.0288639f //x=60.185 //y=7.4
c1150 ( 679 0 ) capacitor c=0.0288633f //x=59.305 //y=7.4
c1151 ( 671 0 ) capacitor c=0.0240981f //x=58.425 //y=7.4
c1152 ( 665 0 ) capacitor c=0.0236947f //x=57.55 //y=7.4
c1153 ( 655 0 ) capacitor c=0.0288598f //x=56.855 //y=7.4
c1154 ( 647 0 ) capacitor c=0.0288369f //x=55.975 //y=7.4
c1155 ( 639 0 ) capacitor c=0.0240981f //x=55.095 //y=7.4
c1156 ( 635 0 ) capacitor c=0.0236224f //x=54.22 //y=7.4
c1157 ( 627 0 ) capacitor c=0.0288359f //x=53.525 //y=7.4
c1158 ( 617 0 ) capacitor c=0.0288369f //x=52.645 //y=7.4
c1159 ( 607 0 ) capacitor c=0.0240981f //x=51.765 //y=7.4
c1160 ( 603 0 ) capacitor c=0.0236224f //x=50.89 //y=7.4
c1161 ( 593 0 ) capacitor c=0.0288359f //x=50.195 //y=7.4
c1162 ( 583 0 ) capacitor c=0.0288369f //x=49.315 //y=7.4
c1163 ( 575 0 ) capacitor c=0.0240981f //x=48.435 //y=7.4
c1164 ( 569 0 ) capacitor c=0.0394667f //x=47.56 //y=7.4
c1165 ( 559 0 ) capacitor c=0.0288488f //x=46.565 //y=7.4
c1166 ( 549 0 ) capacitor c=0.0287505f //x=45.685 //y=7.4
c1167 ( 541 0 ) capacitor c=0.0284966f //x=44.805 //y=7.4
c1168 ( 533 0 ) capacitor c=0.0383672f //x=43.925 //y=7.4
c1169 ( 527 0 ) capacitor c=0.0236224f //x=42.75 //y=7.4
c1170 ( 517 0 ) capacitor c=0.0288359f //x=42.055 //y=7.4
c1171 ( 509 0 ) capacitor c=0.0288369f //x=41.175 //y=7.4
c1172 ( 501 0 ) capacitor c=0.0240981f //x=40.295 //y=7.4
c1173 ( 497 0 ) capacitor c=0.0236224f //x=39.42 //y=7.4
c1174 ( 489 0 ) capacitor c=0.0288359f //x=38.725 //y=7.4
c1175 ( 479 0 ) capacitor c=0.0288369f //x=37.845 //y=7.4
c1176 ( 469 0 ) capacitor c=0.0240981f //x=36.965 //y=7.4
c1177 ( 465 0 ) capacitor c=0.0236224f //x=36.09 //y=7.4
c1178 ( 455 0 ) capacitor c=0.0288357f //x=35.395 //y=7.4
c1179 ( 445 0 ) capacitor c=0.0288369f //x=34.515 //y=7.4
c1180 ( 437 0 ) capacitor c=0.0240981f //x=33.635 //y=7.4
c1181 ( 431 0 ) capacitor c=0.0236224f //x=32.76 //y=7.4
c1182 ( 421 0 ) capacitor c=0.0288359f //x=32.065 //y=7.4
c1183 ( 413 0 ) capacitor c=0.0288369f //x=31.185 //y=7.4
c1184 ( 405 0 ) capacitor c=0.0240981f //x=30.305 //y=7.4
c1185 ( 401 0 ) capacitor c=0.0236224f //x=29.43 //y=7.4
c1186 ( 393 0 ) capacitor c=0.0288359f //x=28.735 //y=7.4
c1187 ( 383 0 ) capacitor c=0.0288369f //x=27.855 //y=7.4
c1188 ( 373 0 ) capacitor c=0.0240981f //x=26.975 //y=7.4
c1189 ( 369 0 ) capacitor c=0.0394667f //x=26.1 //y=7.4
c1190 ( 361 0 ) capacitor c=0.0288488f //x=25.105 //y=7.4
c1191 ( 351 0 ) capacitor c=0.0287505f //x=24.225 //y=7.4
c1192 ( 341 0 ) capacitor c=0.0284966f //x=23.345 //y=7.4
c1193 ( 331 0 ) capacitor c=0.0383672f //x=22.465 //y=7.4
c1194 ( 327 0 ) capacitor c=0.0236224f //x=21.29 //y=7.4
c1195 ( 317 0 ) capacitor c=0.0288359f //x=20.595 //y=7.4
c1196 ( 307 0 ) capacitor c=0.0288369f //x=19.715 //y=7.4
c1197 ( 299 0 ) capacitor c=0.0240981f //x=18.835 //y=7.4
c1198 ( 293 0 ) capacitor c=0.0236224f //x=17.96 //y=7.4
c1199 ( 283 0 ) capacitor c=0.0288359f //x=17.265 //y=7.4
c1200 ( 275 0 ) capacitor c=0.0288373f //x=16.385 //y=7.4
c1201 ( 267 0 ) capacitor c=0.0240981f //x=15.505 //y=7.4
c1202 ( 263 0 ) capacitor c=0.0236224f //x=14.63 //y=7.4
c1203 ( 255 0 ) capacitor c=0.0288361f //x=13.935 //y=7.4
c1204 ( 245 0 ) capacitor c=0.0288369f //x=13.055 //y=7.4
c1205 ( 235 0 ) capacitor c=0.0240981f //x=12.175 //y=7.4
c1206 ( 231 0 ) capacitor c=0.0236224f //x=11.3 //y=7.4
c1207 ( 221 0 ) capacitor c=0.0288359f //x=10.605 //y=7.4
c1208 ( 211 0 ) capacitor c=0.0288369f //x=9.725 //y=7.4
c1209 ( 203 0 ) capacitor c=0.0240981f //x=8.845 //y=7.4
c1210 ( 197 0 ) capacitor c=0.0236224f //x=7.97 //y=7.4
c1211 ( 187 0 ) capacitor c=0.0288359f //x=7.275 //y=7.4
c1212 ( 179 0 ) capacitor c=0.0288369f //x=6.395 //y=7.4
c1213 ( 171 0 ) capacitor c=0.0240981f //x=5.515 //y=7.4
c1214 ( 165 0 ) capacitor c=0.0394667f //x=4.64 //y=7.4
c1215 ( 155 0 ) capacitor c=0.0288488f //x=3.645 //y=7.4
c1216 ( 147 0 ) capacitor c=0.0287505f //x=2.765 //y=7.4
c1217 ( 137 0 ) capacitor c=0.028511f //x=1.885 //y=7.4
c1218 ( 130 0 ) capacitor c=0.234426f //x=0.74 //y=7.4
c1219 ( 127 0 ) capacitor c=0.0452081f //x=1.005 //y=7.4
c1220 ( 123 0 ) capacitor c=2.44404f //x=73.63 //y=7.4
r1221 (  780 782 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=72.52 //y=7.4 //x2=73.63 //y2=7.4
r1222 (  778 780 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=71.41 //y=7.4 //x2=72.52 //y2=7.4
r1223 (  776 877 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=71.21 //y=7.4 //x2=71.04 //y2=7.4
r1224 (  776 778 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=71.21 //y=7.4 //x2=71.41 //y2=7.4
r1225 (  770 772 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=68.82 //y=7.4 //x2=69.93 //y2=7.4
r1226 (  768 876 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.88 //y=7.4 //x2=67.71 //y2=7.4
r1227 (  768 770 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=67.88 //y=7.4 //x2=68.82 //y2=7.4
r1228 (  767 877 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=70.87 //y=7.4 //x2=71.04 //y2=7.4
r1229 (  767 772 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=70.87 //y=7.4 //x2=69.93 //y2=7.4
r1230 (  762 875 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.015 //y=7.4 //x2=66.93 //y2=7.4
r1231 (  762 764 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=67.015 //y=7.4 //x2=67.34 //y2=7.4
r1232 (  761 876 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.54 //y=7.4 //x2=67.71 //y2=7.4
r1233 (  761 764 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=67.54 //y=7.4 //x2=67.34 //y2=7.4
r1234 (  755 875 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=66.93 //y=7.23 //x2=66.93 //y2=7.4
r1235 (  755 937 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=66.93 //y=7.23 //x2=66.93 //y2=6.4
r1236 (  752 874 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.135 //y=7.4 //x2=66.05 //y2=7.4
r1237 (  752 754 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=66.135 //y=7.4 //x2=66.23 //y2=7.4
r1238 (  751 875 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.845 //y=7.4 //x2=66.93 //y2=7.4
r1239 (  751 754 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=66.845 //y=7.4 //x2=66.23 //y2=7.4
r1240 (  745 874 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=66.05 //y=7.23 //x2=66.05 //y2=7.4
r1241 (  745 936 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=66.05 //y=7.23 //x2=66.05 //y2=6.74
r1242 (  744 873 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.255 //y=7.4 //x2=65.17 //y2=7.4
r1243 (  743 874 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.965 //y=7.4 //x2=66.05 //y2=7.4
r1244 (  743 744 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=65.965 //y=7.4 //x2=65.255 //y2=7.4
r1245 (  737 873 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=65.17 //y=7.23 //x2=65.17 //y2=7.4
r1246 (  737 935 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=65.17 //y=7.23 //x2=65.17 //y2=6.4
r1247 (  736 871 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.55 //y=7.4 //x2=64.38 //y2=7.4
r1248 (  735 873 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.085 //y=7.4 //x2=65.17 //y2=7.4
r1249 (  735 736 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=65.085 //y=7.4 //x2=64.55 //y2=7.4
r1250 (  732 870 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.685 //y=7.4 //x2=63.6 //y2=7.4
r1251 (  731 871 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.21 //y=7.4 //x2=64.38 //y2=7.4
r1252 (  731 732 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=64.21 //y=7.4 //x2=63.685 //y2=7.4
r1253 (  725 870 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=63.6 //y=7.23 //x2=63.6 //y2=7.4
r1254 (  725 934 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=63.6 //y=7.23 //x2=63.6 //y2=6.745
r1255 (  724 868 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.805 //y=7.4 //x2=62.72 //y2=7.4
r1256 (  723 870 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.515 //y=7.4 //x2=63.6 //y2=7.4
r1257 (  723 724 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=63.515 //y=7.4 //x2=62.805 //y2=7.4
r1258 (  717 868 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.72 //y=7.23 //x2=62.72 //y2=7.4
r1259 (  717 933 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=62.72 //y=7.23 //x2=62.72 //y2=6.745
r1260 (  714 867 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=61.925 //y=7.4 //x2=61.84 //y2=7.4
r1261 (  714 716 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=61.925 //y=7.4 //x2=62.53 //y2=7.4
r1262 (  713 868 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.635 //y=7.4 //x2=62.72 //y2=7.4
r1263 (  713 716 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=62.635 //y=7.4 //x2=62.53 //y2=7.4
r1264 (  707 867 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.84 //y=7.23 //x2=61.84 //y2=7.4
r1265 (  707 932 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=61.84 //y=7.23 //x2=61.84 //y2=6.405
r1266 (  704 866 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.22 //y=7.4 //x2=61.05 //y2=7.4
r1267 (  704 706 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=61.22 //y=7.4 //x2=61.42 //y2=7.4
r1268 (  703 867 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=61.755 //y=7.4 //x2=61.84 //y2=7.4
r1269 (  703 706 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=61.755 //y=7.4 //x2=61.42 //y2=7.4
r1270 (  700 865 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.355 //y=7.4 //x2=60.27 //y2=7.4
r1271 (  699 866 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=60.88 //y=7.4 //x2=61.05 //y2=7.4
r1272 (  699 700 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=60.88 //y=7.4 //x2=60.355 //y2=7.4
r1273 (  693 865 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=60.27 //y=7.23 //x2=60.27 //y2=7.4
r1274 (  693 931 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=60.27 //y=7.23 //x2=60.27 //y2=6.745
r1275 (  690 864 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.475 //y=7.4 //x2=59.39 //y2=7.4
r1276 (  690 692 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=59.475 //y=7.4 //x2=59.94 //y2=7.4
r1277 (  689 865 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.185 //y=7.4 //x2=60.27 //y2=7.4
r1278 (  689 692 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=60.185 //y=7.4 //x2=59.94 //y2=7.4
r1279 (  683 864 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=59.39 //y=7.23 //x2=59.39 //y2=7.4
r1280 (  683 930 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=59.39 //y=7.23 //x2=59.39 //y2=6.745
r1281 (  680 863 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.595 //y=7.4 //x2=58.51 //y2=7.4
r1282 (  680 682 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=58.595 //y=7.4 //x2=58.83 //y2=7.4
r1283 (  679 864 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.305 //y=7.4 //x2=59.39 //y2=7.4
r1284 (  679 682 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=59.305 //y=7.4 //x2=58.83 //y2=7.4
r1285 (  673 863 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.51 //y=7.23 //x2=58.51 //y2=7.4
r1286 (  673 929 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=58.51 //y=7.23 //x2=58.51 //y2=6.405
r1287 (  672 862 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.89 //y=7.4 //x2=57.72 //y2=7.4
r1288 (  671 863 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.425 //y=7.4 //x2=58.51 //y2=7.4
r1289 (  671 672 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=58.425 //y=7.4 //x2=57.89 //y2=7.4
r1290 (  666 861 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=57.025 //y=7.4 //x2=56.94 //y2=7.4
r1291 (  666 668 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=57.025 //y=7.4 //x2=57.35 //y2=7.4
r1292 (  665 862 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.55 //y=7.4 //x2=57.72 //y2=7.4
r1293 (  665 668 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=57.55 //y=7.4 //x2=57.35 //y2=7.4
r1294 (  659 861 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=56.94 //y=7.23 //x2=56.94 //y2=7.4
r1295 (  659 928 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=56.94 //y=7.23 //x2=56.94 //y2=6.745
r1296 (  656 860 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.145 //y=7.4 //x2=56.06 //y2=7.4
r1297 (  656 658 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=56.145 //y=7.4 //x2=56.24 //y2=7.4
r1298 (  655 861 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.855 //y=7.4 //x2=56.94 //y2=7.4
r1299 (  655 658 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=56.855 //y=7.4 //x2=56.24 //y2=7.4
r1300 (  649 860 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=56.06 //y=7.23 //x2=56.06 //y2=7.4
r1301 (  649 927 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=56.06 //y=7.23 //x2=56.06 //y2=6.745
r1302 (  648 859 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.265 //y=7.4 //x2=55.18 //y2=7.4
r1303 (  647 860 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.975 //y=7.4 //x2=56.06 //y2=7.4
r1304 (  647 648 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=55.975 //y=7.4 //x2=55.265 //y2=7.4
r1305 (  641 859 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=55.18 //y=7.23 //x2=55.18 //y2=7.4
r1306 (  641 926 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=55.18 //y=7.23 //x2=55.18 //y2=6.405
r1307 (  640 857 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=54.56 //y=7.4 //x2=54.39 //y2=7.4
r1308 (  639 859 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.095 //y=7.4 //x2=55.18 //y2=7.4
r1309 (  639 640 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=55.095 //y=7.4 //x2=54.56 //y2=7.4
r1310 (  636 856 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.695 //y=7.4 //x2=53.61 //y2=7.4
r1311 (  635 857 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=54.22 //y=7.4 //x2=54.39 //y2=7.4
r1312 (  635 636 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=54.22 //y=7.4 //x2=53.695 //y2=7.4
r1313 (  629 856 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=53.61 //y=7.23 //x2=53.61 //y2=7.4
r1314 (  629 925 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=53.61 //y=7.23 //x2=53.61 //y2=6.745
r1315 (  628 854 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=52.815 //y=7.4 //x2=52.73 //y2=7.4
r1316 (  627 856 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.525 //y=7.4 //x2=53.61 //y2=7.4
r1317 (  627 628 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=53.525 //y=7.4 //x2=52.815 //y2=7.4
r1318 (  621 854 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=52.73 //y=7.23 //x2=52.73 //y2=7.4
r1319 (  621 924 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=52.73 //y=7.23 //x2=52.73 //y2=6.745
r1320 (  618 853 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.935 //y=7.4 //x2=51.85 //y2=7.4
r1321 (  618 620 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=51.935 //y=7.4 //x2=52.54 //y2=7.4
r1322 (  617 854 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=52.645 //y=7.4 //x2=52.73 //y2=7.4
r1323 (  617 620 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=52.645 //y=7.4 //x2=52.54 //y2=7.4
r1324 (  611 853 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=51.85 //y=7.23 //x2=51.85 //y2=7.4
r1325 (  611 923 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=51.85 //y=7.23 //x2=51.85 //y2=6.405
r1326 (  608 852 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=51.23 //y=7.4 //x2=51.06 //y2=7.4
r1327 (  608 610 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=51.23 //y=7.4 //x2=51.43 //y2=7.4
r1328 (  607 853 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.765 //y=7.4 //x2=51.85 //y2=7.4
r1329 (  607 610 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=51.765 //y=7.4 //x2=51.43 //y2=7.4
r1330 (  604 851 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.365 //y=7.4 //x2=50.28 //y2=7.4
r1331 (  603 852 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=50.89 //y=7.4 //x2=51.06 //y2=7.4
r1332 (  603 604 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=50.89 //y=7.4 //x2=50.365 //y2=7.4
r1333 (  597 851 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=50.28 //y=7.23 //x2=50.28 //y2=7.4
r1334 (  597 922 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=50.28 //y=7.23 //x2=50.28 //y2=6.745
r1335 (  594 850 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.485 //y=7.4 //x2=49.4 //y2=7.4
r1336 (  594 596 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=49.485 //y=7.4 //x2=49.95 //y2=7.4
r1337 (  593 851 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.195 //y=7.4 //x2=50.28 //y2=7.4
r1338 (  593 596 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=50.195 //y=7.4 //x2=49.95 //y2=7.4
r1339 (  587 850 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.4 //y=7.23 //x2=49.4 //y2=7.4
r1340 (  587 921 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=49.4 //y=7.23 //x2=49.4 //y2=6.745
r1341 (  584 849 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=48.605 //y=7.4 //x2=48.52 //y2=7.4
r1342 (  584 586 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=48.605 //y=7.4 //x2=48.84 //y2=7.4
r1343 (  583 850 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.315 //y=7.4 //x2=49.4 //y2=7.4
r1344 (  583 586 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=49.315 //y=7.4 //x2=48.84 //y2=7.4
r1345 (  577 849 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.52 //y=7.23 //x2=48.52 //y2=7.4
r1346 (  577 920 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=48.52 //y=7.23 //x2=48.52 //y2=6.405
r1347 (  576 848 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.9 //y=7.4 //x2=47.73 //y2=7.4
r1348 (  575 849 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=48.435 //y=7.4 //x2=48.52 //y2=7.4
r1349 (  575 576 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=48.435 //y=7.4 //x2=47.9 //y2=7.4
r1350 (  570 847 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.735 //y=7.4 //x2=46.65 //y2=7.4
r1351 (  570 572 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=46.735 //y=7.4 //x2=47.36 //y2=7.4
r1352 (  569 848 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.56 //y=7.4 //x2=47.73 //y2=7.4
r1353 (  569 572 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=47.56 //y=7.4 //x2=47.36 //y2=7.4
r1354 (  563 847 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=46.65 //y=7.23 //x2=46.65 //y2=7.4
r1355 (  563 919 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.65 //y=7.23 //x2=46.65 //y2=6.745
r1356 (  560 846 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.855 //y=7.4 //x2=45.77 //y2=7.4
r1357 (  560 562 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=45.855 //y=7.4 //x2=46.25 //y2=7.4
r1358 (  559 847 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.565 //y=7.4 //x2=46.65 //y2=7.4
r1359 (  559 562 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=46.565 //y=7.4 //x2=46.25 //y2=7.4
r1360 (  553 846 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=45.77 //y=7.23 //x2=45.77 //y2=7.4
r1361 (  553 918 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=45.77 //y=7.23 //x2=45.77 //y2=6.745
r1362 (  550 845 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.975 //y=7.4 //x2=44.89 //y2=7.4
r1363 (  550 552 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=44.975 //y=7.4 //x2=45.14 //y2=7.4
r1364 (  549 846 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.685 //y=7.4 //x2=45.77 //y2=7.4
r1365 (  549 552 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=45.685 //y=7.4 //x2=45.14 //y2=7.4
r1366 (  543 845 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=44.89 //y=7.23 //x2=44.89 //y2=7.4
r1367 (  543 917 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=44.89 //y=7.23 //x2=44.89 //y2=6.745
r1368 (  542 844 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.095 //y=7.4 //x2=44.01 //y2=7.4
r1369 (  541 845 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.805 //y=7.4 //x2=44.89 //y2=7.4
r1370 (  541 542 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=44.805 //y=7.4 //x2=44.095 //y2=7.4
r1371 (  535 844 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=44.01 //y=7.23 //x2=44.01 //y2=7.4
r1372 (  535 916 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=44.01 //y=7.23 //x2=44.01 //y2=6.405
r1373 (  534 842 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.09 //y=7.4 //x2=42.92 //y2=7.4
r1374 (  533 844 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=43.925 //y=7.4 //x2=44.01 //y2=7.4
r1375 (  533 534 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=43.925 //y=7.4 //x2=43.09 //y2=7.4
r1376 (  528 841 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.225 //y=7.4 //x2=42.14 //y2=7.4
r1377 (  528 530 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=42.225 //y=7.4 //x2=42.55 //y2=7.4
r1378 (  527 842 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=42.75 //y=7.4 //x2=42.92 //y2=7.4
r1379 (  527 530 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=42.75 //y=7.4 //x2=42.55 //y2=7.4
r1380 (  521 841 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=42.14 //y=7.23 //x2=42.14 //y2=7.4
r1381 (  521 915 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=42.14 //y=7.23 //x2=42.14 //y2=6.745
r1382 (  518 840 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.345 //y=7.4 //x2=41.26 //y2=7.4
r1383 (  518 520 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=41.345 //y=7.4 //x2=41.44 //y2=7.4
r1384 (  517 841 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.055 //y=7.4 //x2=42.14 //y2=7.4
r1385 (  517 520 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=42.055 //y=7.4 //x2=41.44 //y2=7.4
r1386 (  511 840 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=41.26 //y=7.23 //x2=41.26 //y2=7.4
r1387 (  511 914 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=41.26 //y=7.23 //x2=41.26 //y2=6.745
r1388 (  510 839 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.465 //y=7.4 //x2=40.38 //y2=7.4
r1389 (  509 840 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.175 //y=7.4 //x2=41.26 //y2=7.4
r1390 (  509 510 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=41.175 //y=7.4 //x2=40.465 //y2=7.4
r1391 (  503 839 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.38 //y=7.23 //x2=40.38 //y2=7.4
r1392 (  503 913 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=40.38 //y=7.23 //x2=40.38 //y2=6.405
r1393 (  502 837 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.76 //y=7.4 //x2=39.59 //y2=7.4
r1394 (  501 839 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.295 //y=7.4 //x2=40.38 //y2=7.4
r1395 (  501 502 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=40.295 //y=7.4 //x2=39.76 //y2=7.4
r1396 (  498 836 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.895 //y=7.4 //x2=38.81 //y2=7.4
r1397 (  497 837 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.42 //y=7.4 //x2=39.59 //y2=7.4
r1398 (  497 498 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=39.42 //y=7.4 //x2=38.895 //y2=7.4
r1399 (  491 836 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.81 //y=7.23 //x2=38.81 //y2=7.4
r1400 (  491 912 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=38.81 //y=7.23 //x2=38.81 //y2=6.745
r1401 (  490 834 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.015 //y=7.4 //x2=37.93 //y2=7.4
r1402 (  489 836 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.725 //y=7.4 //x2=38.81 //y2=7.4
r1403 (  489 490 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=38.725 //y=7.4 //x2=38.015 //y2=7.4
r1404 (  483 834 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.93 //y=7.23 //x2=37.93 //y2=7.4
r1405 (  483 911 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=37.93 //y=7.23 //x2=37.93 //y2=6.745
r1406 (  480 833 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.135 //y=7.4 //x2=37.05 //y2=7.4
r1407 (  480 482 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=37.135 //y=7.4 //x2=37.74 //y2=7.4
r1408 (  479 834 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.845 //y=7.4 //x2=37.93 //y2=7.4
r1409 (  479 482 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=37.845 //y=7.4 //x2=37.74 //y2=7.4
r1410 (  473 833 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.05 //y=7.23 //x2=37.05 //y2=7.4
r1411 (  473 910 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=37.05 //y=7.23 //x2=37.05 //y2=6.405
r1412 (  470 832 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.43 //y=7.4 //x2=36.26 //y2=7.4
r1413 (  470 472 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=36.43 //y=7.4 //x2=36.63 //y2=7.4
r1414 (  469 833 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.965 //y=7.4 //x2=37.05 //y2=7.4
r1415 (  469 472 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=36.965 //y=7.4 //x2=36.63 //y2=7.4
r1416 (  466 831 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.565 //y=7.4 //x2=35.48 //y2=7.4
r1417 (  465 832 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.09 //y=7.4 //x2=36.26 //y2=7.4
r1418 (  465 466 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=36.09 //y=7.4 //x2=35.565 //y2=7.4
r1419 (  459 831 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=35.48 //y=7.23 //x2=35.48 //y2=7.4
r1420 (  459 909 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=35.48 //y=7.23 //x2=35.48 //y2=6.745
r1421 (  456 830 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.685 //y=7.4 //x2=34.6 //y2=7.4
r1422 (  456 458 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=34.685 //y=7.4 //x2=35.15 //y2=7.4
r1423 (  455 831 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.395 //y=7.4 //x2=35.48 //y2=7.4
r1424 (  455 458 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=35.395 //y=7.4 //x2=35.15 //y2=7.4
r1425 (  449 830 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=34.6 //y=7.23 //x2=34.6 //y2=7.4
r1426 (  449 908 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=34.6 //y=7.23 //x2=34.6 //y2=6.745
r1427 (  446 829 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.805 //y=7.4 //x2=33.72 //y2=7.4
r1428 (  446 448 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=33.805 //y=7.4 //x2=34.04 //y2=7.4
r1429 (  445 830 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.515 //y=7.4 //x2=34.6 //y2=7.4
r1430 (  445 448 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=34.515 //y=7.4 //x2=34.04 //y2=7.4
r1431 (  439 829 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.72 //y=7.23 //x2=33.72 //y2=7.4
r1432 (  439 907 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=33.72 //y=7.23 //x2=33.72 //y2=6.405
r1433 (  438 828 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.1 //y=7.4 //x2=32.93 //y2=7.4
r1434 (  437 829 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.635 //y=7.4 //x2=33.72 //y2=7.4
r1435 (  437 438 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=33.635 //y=7.4 //x2=33.1 //y2=7.4
r1436 (  432 827 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.235 //y=7.4 //x2=32.15 //y2=7.4
r1437 (  432 434 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=32.235 //y=7.4 //x2=32.56 //y2=7.4
r1438 (  431 828 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.76 //y=7.4 //x2=32.93 //y2=7.4
r1439 (  431 434 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=32.76 //y=7.4 //x2=32.56 //y2=7.4
r1440 (  425 827 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.15 //y=7.23 //x2=32.15 //y2=7.4
r1441 (  425 906 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=32.15 //y=7.23 //x2=32.15 //y2=6.745
r1442 (  422 826 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.355 //y=7.4 //x2=31.27 //y2=7.4
r1443 (  422 424 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=31.355 //y=7.4 //x2=31.45 //y2=7.4
r1444 (  421 827 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.065 //y=7.4 //x2=32.15 //y2=7.4
r1445 (  421 424 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=32.065 //y=7.4 //x2=31.45 //y2=7.4
r1446 (  415 826 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=31.27 //y=7.23 //x2=31.27 //y2=7.4
r1447 (  415 905 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=31.27 //y=7.23 //x2=31.27 //y2=6.745
r1448 (  414 825 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.475 //y=7.4 //x2=30.39 //y2=7.4
r1449 (  413 826 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.185 //y=7.4 //x2=31.27 //y2=7.4
r1450 (  413 414 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=31.185 //y=7.4 //x2=30.475 //y2=7.4
r1451 (  407 825 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.39 //y=7.23 //x2=30.39 //y2=7.4
r1452 (  407 904 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=30.39 //y=7.23 //x2=30.39 //y2=6.405
r1453 (  406 823 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.77 //y=7.4 //x2=29.6 //y2=7.4
r1454 (  405 825 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.305 //y=7.4 //x2=30.39 //y2=7.4
r1455 (  405 406 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=30.305 //y=7.4 //x2=29.77 //y2=7.4
r1456 (  402 822 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.905 //y=7.4 //x2=28.82 //y2=7.4
r1457 (  401 823 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.43 //y=7.4 //x2=29.6 //y2=7.4
r1458 (  401 402 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=29.43 //y=7.4 //x2=28.905 //y2=7.4
r1459 (  395 822 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=28.82 //y=7.23 //x2=28.82 //y2=7.4
r1460 (  395 903 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=28.82 //y=7.23 //x2=28.82 //y2=6.745
r1461 (  394 820 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.025 //y=7.4 //x2=27.94 //y2=7.4
r1462 (  393 822 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.735 //y=7.4 //x2=28.82 //y2=7.4
r1463 (  393 394 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=28.735 //y=7.4 //x2=28.025 //y2=7.4
r1464 (  387 820 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.94 //y=7.23 //x2=27.94 //y2=7.4
r1465 (  387 902 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=27.94 //y=7.23 //x2=27.94 //y2=6.745
r1466 (  384 819 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.145 //y=7.4 //x2=27.06 //y2=7.4
r1467 (  384 386 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=27.145 //y=7.4 //x2=27.75 //y2=7.4
r1468 (  383 820 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.855 //y=7.4 //x2=27.94 //y2=7.4
r1469 (  383 386 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=27.855 //y=7.4 //x2=27.75 //y2=7.4
r1470 (  377 819 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.06 //y=7.23 //x2=27.06 //y2=7.4
r1471 (  377 901 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=27.06 //y=7.23 //x2=27.06 //y2=6.405
r1472 (  374 818 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.44 //y=7.4 //x2=26.27 //y2=7.4
r1473 (  374 376 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=26.44 //y=7.4 //x2=26.64 //y2=7.4
r1474 (  373 819 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.975 //y=7.4 //x2=27.06 //y2=7.4
r1475 (  373 376 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=26.975 //y=7.4 //x2=26.64 //y2=7.4
r1476 (  370 817 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.275 //y=7.4 //x2=25.19 //y2=7.4
r1477 (  369 818 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.1 //y=7.4 //x2=26.27 //y2=7.4
r1478 (  369 370 ) resistor r=29.5798 //w=0.357 //l=0.825 //layer=li \
 //thickness=0.1 //x=26.1 //y=7.4 //x2=25.275 //y2=7.4
r1479 (  363 817 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.19 //y=7.23 //x2=25.19 //y2=7.4
r1480 (  363 900 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=25.19 //y=7.23 //x2=25.19 //y2=6.745
r1481 (  362 815 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.395 //y=7.4 //x2=24.31 //y2=7.4
r1482 (  361 817 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.105 //y=7.4 //x2=25.19 //y2=7.4
r1483 (  361 362 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=25.105 //y=7.4 //x2=24.395 //y2=7.4
r1484 (  355 815 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.31 //y=7.23 //x2=24.31 //y2=7.4
r1485 (  355 899 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=24.31 //y=7.23 //x2=24.31 //y2=6.745
r1486 (  352 814 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.515 //y=7.4 //x2=23.43 //y2=7.4
r1487 (  352 354 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=23.515 //y=7.4 //x2=24.05 //y2=7.4
r1488 (  351 815 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.225 //y=7.4 //x2=24.31 //y2=7.4
r1489 (  351 354 ) resistor r=6.27451 //w=0.357 //l=0.175 //layer=li \
 //thickness=0.1 //x=24.225 //y=7.4 //x2=24.05 //y2=7.4
r1490 (  345 814 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.43 //y=7.23 //x2=23.43 //y2=7.4
r1491 (  345 898 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=23.43 //y=7.23 //x2=23.43 //y2=6.745
r1492 (  342 813 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.635 //y=7.4 //x2=22.55 //y2=7.4
r1493 (  342 344 ) resistor r=10.9356 //w=0.357 //l=0.305 //layer=li \
 //thickness=0.1 //x=22.635 //y=7.4 //x2=22.94 //y2=7.4
r1494 (  341 814 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.345 //y=7.4 //x2=23.43 //y2=7.4
r1495 (  341 344 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=23.345 //y=7.4 //x2=22.94 //y2=7.4
r1496 (  335 813 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.55 //y=7.23 //x2=22.55 //y2=7.4
r1497 (  335 897 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=22.55 //y=7.23 //x2=22.55 //y2=6.405
r1498 (  332 812 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.63 //y=7.4 //x2=21.46 //y2=7.4
r1499 (  332 334 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=21.63 //y=7.4 //x2=21.83 //y2=7.4
r1500 (  331 813 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.465 //y=7.4 //x2=22.55 //y2=7.4
r1501 (  331 334 ) resistor r=22.7675 //w=0.357 //l=0.635 //layer=li \
 //thickness=0.1 //x=22.465 //y=7.4 //x2=21.83 //y2=7.4
r1502 (  328 811 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.765 //y=7.4 //x2=20.68 //y2=7.4
r1503 (  327 812 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.29 //y=7.4 //x2=21.46 //y2=7.4
r1504 (  327 328 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=21.29 //y=7.4 //x2=20.765 //y2=7.4
r1505 (  321 811 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.68 //y=7.23 //x2=20.68 //y2=7.4
r1506 (  321 896 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.68 //y=7.23 //x2=20.68 //y2=6.745
r1507 (  318 810 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.885 //y=7.4 //x2=19.8 //y2=7.4
r1508 (  318 320 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=19.885 //y=7.4 //x2=20.35 //y2=7.4
r1509 (  317 811 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.595 //y=7.4 //x2=20.68 //y2=7.4
r1510 (  317 320 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=20.595 //y=7.4 //x2=20.35 //y2=7.4
r1511 (  311 810 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.8 //y=7.23 //x2=19.8 //y2=7.4
r1512 (  311 895 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=19.8 //y=7.23 //x2=19.8 //y2=6.745
r1513 (  308 809 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.005 //y=7.4 //x2=18.92 //y2=7.4
r1514 (  308 310 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=19.005 //y=7.4 //x2=19.24 //y2=7.4
r1515 (  307 810 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.715 //y=7.4 //x2=19.8 //y2=7.4
r1516 (  307 310 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=19.715 //y=7.4 //x2=19.24 //y2=7.4
r1517 (  301 809 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.92 //y=7.23 //x2=18.92 //y2=7.4
r1518 (  301 894 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=18.92 //y=7.23 //x2=18.92 //y2=6.405
r1519 (  300 808 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.3 //y=7.4 //x2=18.13 //y2=7.4
r1520 (  299 809 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.835 //y=7.4 //x2=18.92 //y2=7.4
r1521 (  299 300 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=18.835 //y=7.4 //x2=18.3 //y2=7.4
r1522 (  294 807 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.435 //y=7.4 //x2=17.35 //y2=7.4
r1523 (  294 296 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=17.435 //y=7.4 //x2=17.76 //y2=7.4
r1524 (  293 808 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.96 //y=7.4 //x2=18.13 //y2=7.4
r1525 (  293 296 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=17.96 //y=7.4 //x2=17.76 //y2=7.4
r1526 (  287 807 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.35 //y=7.23 //x2=17.35 //y2=7.4
r1527 (  287 893 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.35 //y=7.23 //x2=17.35 //y2=6.745
r1528 (  284 806 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.555 //y=7.4 //x2=16.47 //y2=7.4
r1529 (  284 286 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=16.555 //y=7.4 //x2=16.65 //y2=7.4
r1530 (  283 807 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.265 //y=7.4 //x2=17.35 //y2=7.4
r1531 (  283 286 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=17.265 //y=7.4 //x2=16.65 //y2=7.4
r1532 (  277 806 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.47 //y=7.23 //x2=16.47 //y2=7.4
r1533 (  277 892 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.47 //y=7.23 //x2=16.47 //y2=6.745
r1534 (  276 805 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.675 //y=7.4 //x2=15.59 //y2=7.4
r1535 (  275 806 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.385 //y=7.4 //x2=16.47 //y2=7.4
r1536 (  275 276 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=16.385 //y=7.4 //x2=15.675 //y2=7.4
r1537 (  269 805 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.59 //y=7.23 //x2=15.59 //y2=7.4
r1538 (  269 891 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=15.59 //y=7.23 //x2=15.59 //y2=6.405
r1539 (  268 803 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.97 //y=7.4 //x2=14.8 //y2=7.4
r1540 (  267 805 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.505 //y=7.4 //x2=15.59 //y2=7.4
r1541 (  267 268 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=15.505 //y=7.4 //x2=14.97 //y2=7.4
r1542 (  264 802 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.105 //y=7.4 //x2=14.02 //y2=7.4
r1543 (  263 803 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.63 //y=7.4 //x2=14.8 //y2=7.4
r1544 (  263 264 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=14.63 //y=7.4 //x2=14.105 //y2=7.4
r1545 (  257 802 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.02 //y=7.23 //x2=14.02 //y2=7.4
r1546 (  257 890 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.02 //y=7.23 //x2=14.02 //y2=6.745
r1547 (  256 800 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.225 //y=7.4 //x2=13.14 //y2=7.4
r1548 (  255 802 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.935 //y=7.4 //x2=14.02 //y2=7.4
r1549 (  255 256 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=13.935 //y=7.4 //x2=13.225 //y2=7.4
r1550 (  249 800 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.14 //y=7.23 //x2=13.14 //y2=7.4
r1551 (  249 889 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=13.14 //y=7.23 //x2=13.14 //y2=6.745
r1552 (  246 799 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.345 //y=7.4 //x2=12.26 //y2=7.4
r1553 (  246 248 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=12.345 //y=7.4 //x2=12.95 //y2=7.4
r1554 (  245 800 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.055 //y=7.4 //x2=13.14 //y2=7.4
r1555 (  245 248 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=13.055 //y=7.4 //x2=12.95 //y2=7.4
r1556 (  239 799 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.26 //y=7.23 //x2=12.26 //y2=7.4
r1557 (  239 888 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=12.26 //y=7.23 //x2=12.26 //y2=6.405
r1558 (  236 798 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.64 //y=7.4 //x2=11.47 //y2=7.4
r1559 (  236 238 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=11.64 //y=7.4 //x2=11.84 //y2=7.4
r1560 (  235 799 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.175 //y=7.4 //x2=12.26 //y2=7.4
r1561 (  235 238 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=12.175 //y=7.4 //x2=11.84 //y2=7.4
r1562 (  232 797 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.775 //y=7.4 //x2=10.69 //y2=7.4
r1563 (  231 798 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.3 //y=7.4 //x2=11.47 //y2=7.4
r1564 (  231 232 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=11.3 //y=7.4 //x2=10.775 //y2=7.4
r1565 (  225 797 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.69 //y=7.23 //x2=10.69 //y2=7.4
r1566 (  225 887 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.69 //y=7.23 //x2=10.69 //y2=6.745
r1567 (  222 796 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.895 //y=7.4 //x2=9.81 //y2=7.4
r1568 (  222 224 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=9.895 //y=7.4 //x2=10.36 //y2=7.4
r1569 (  221 797 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.605 //y=7.4 //x2=10.69 //y2=7.4
r1570 (  221 224 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=10.605 //y=7.4 //x2=10.36 //y2=7.4
r1571 (  215 796 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.81 //y=7.23 //x2=9.81 //y2=7.4
r1572 (  215 886 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=9.81 //y=7.23 //x2=9.81 //y2=6.745
r1573 (  212 795 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.015 //y=7.4 //x2=8.93 //y2=7.4
r1574 (  212 214 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=9.015 //y=7.4 //x2=9.25 //y2=7.4
r1575 (  211 796 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.725 //y=7.4 //x2=9.81 //y2=7.4
r1576 (  211 214 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=9.725 //y=7.4 //x2=9.25 //y2=7.4
r1577 (  205 795 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.93 //y=7.23 //x2=8.93 //y2=7.4
r1578 (  205 885 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=8.93 //y=7.23 //x2=8.93 //y2=6.405
r1579 (  204 794 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=7.4 //x2=8.14 //y2=7.4
r1580 (  203 795 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.845 //y=7.4 //x2=8.93 //y2=7.4
r1581 (  203 204 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=8.845 //y=7.4 //x2=8.31 //y2=7.4
r1582 (  198 793 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.445 //y=7.4 //x2=7.36 //y2=7.4
r1583 (  198 200 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=7.445 //y=7.4 //x2=7.77 //y2=7.4
r1584 (  197 794 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=8.14 //y2=7.4
r1585 (  197 200 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=7.77 //y2=7.4
r1586 (  191 793 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.36 //y=7.23 //x2=7.36 //y2=7.4
r1587 (  191 884 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.36 //y=7.23 //x2=7.36 //y2=6.745
r1588 (  188 792 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.565 //y=7.4 //x2=6.48 //y2=7.4
r1589 (  188 190 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=6.565 //y=7.4 //x2=6.66 //y2=7.4
r1590 (  187 793 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.275 //y=7.4 //x2=7.36 //y2=7.4
r1591 (  187 190 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=7.275 //y=7.4 //x2=6.66 //y2=7.4
r1592 (  181 792 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.48 //y=7.23 //x2=6.48 //y2=7.4
r1593 (  181 883 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.48 //y=7.23 //x2=6.48 //y2=6.745
r1594 (  180 791 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.685 //y=7.4 //x2=5.6 //y2=7.4
r1595 (  179 792 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.395 //y=7.4 //x2=6.48 //y2=7.4
r1596 (  179 180 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=6.395 //y=7.4 //x2=5.685 //y2=7.4
r1597 (  173 791 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.6 //y=7.23 //x2=5.6 //y2=7.4
r1598 (  173 882 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=5.6 //y=7.23 //x2=5.6 //y2=6.405
r1599 (  172 789 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=4.81 //y2=7.4
r1600 (  171 791 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.515 //y=7.4 //x2=5.6 //y2=7.4
r1601 (  171 172 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=5.515 //y=7.4 //x2=4.98 //y2=7.4
r1602 (  166 788 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=3.73 //y2=7.4
r1603 (  166 168 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=4.07 //y2=7.4
r1604 (  165 789 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.81 //y2=7.4
r1605 (  165 168 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.07 //y2=7.4
r1606 (  159 788 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=7.4
r1607 (  159 881 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=6.745
r1608 (  156 787 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.85 //y2=7.4
r1609 (  156 158 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.96 //y2=7.4
r1610 (  155 788 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=3.73 //y2=7.4
r1611 (  155 158 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=2.96 //y2=7.4
r1612 (  149 787 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=7.4
r1613 (  149 880 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=6.745
r1614 (  148 786 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.055 //y=7.4 //x2=1.97 //y2=7.4
r1615 (  147 787 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.85 //y2=7.4
r1616 (  147 148 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.055 //y2=7.4
r1617 (  141 786 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=7.4
r1618 (  141 879 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=6.745
r1619 (  138 785 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.09 //y2=7.4
r1620 (  138 140 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.85 //y2=7.4
r1621 (  137 786 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.97 //y2=7.4
r1622 (  137 140 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.85 //y2=7.4
r1623 (  131 785 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=7.4
r1624 (  131 878 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=6.405
r1625 (  127 785 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=1.09 //y2=7.4
r1626 (  127 130 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=0.74 //y2=7.4
r1627 (  123 782 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=73.63 //y=7.4 //x2=73.63 //y2=7.4
r1628 (  121 780 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=72.52 //y=7.4 //x2=72.52 //y2=7.4
r1629 (  121 123 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=72.52 //y=7.4 //x2=73.63 //y2=7.4
r1630 (  119 778 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=71.41 //y=7.4 //x2=71.41 //y2=7.4
r1631 (  119 121 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=71.41 //y=7.4 //x2=72.52 //y2=7.4
r1632 (  117 772 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=69.93 //y=7.4 //x2=69.93 //y2=7.4
r1633 (  117 119 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=69.93 //y=7.4 //x2=71.41 //y2=7.4
r1634 (  115 770 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=68.82 //y=7.4 //x2=68.82 //y2=7.4
r1635 (  115 117 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=68.82 //y=7.4 //x2=69.93 //y2=7.4
r1636 (  113 764 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=67.34 //y=7.4 //x2=67.34 //y2=7.4
r1637 (  113 115 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=67.34 //y=7.4 //x2=68.82 //y2=7.4
r1638 (  111 754 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=66.23 //y=7.4 //x2=66.23 //y2=7.4
r1639 (  111 113 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=66.23 //y=7.4 //x2=67.34 //y2=7.4
r1640 (  109 873 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=65.12 //y=7.4 //x2=65.12 //y2=7.4
r1641 (  109 111 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=65.12 //y=7.4 //x2=66.23 //y2=7.4
r1642 (  107 870 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=63.64 //y=7.4 //x2=63.64 //y2=7.4
r1643 (  107 109 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=63.64 //y=7.4 //x2=65.12 //y2=7.4
r1644 (  105 716 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=62.53 //y=7.4 //x2=62.53 //y2=7.4
r1645 (  105 107 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=62.53 //y=7.4 //x2=63.64 //y2=7.4
r1646 (  103 706 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=61.42 //y=7.4 //x2=61.42 //y2=7.4
r1647 (  103 105 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=61.42 //y=7.4 //x2=62.53 //y2=7.4
r1648 (  101 692 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=59.94 //y=7.4 //x2=59.94 //y2=7.4
r1649 (  101 103 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=59.94 //y=7.4 //x2=61.42 //y2=7.4
r1650 (  99 682 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=58.83 //y=7.4 //x2=58.83 //y2=7.4
r1651 (  99 101 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=58.83 //y=7.4 //x2=59.94 //y2=7.4
r1652 (  97 668 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=57.35 //y=7.4 //x2=57.35 //y2=7.4
r1653 (  97 99 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=57.35 //y=7.4 //x2=58.83 //y2=7.4
r1654 (  95 658 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=56.24 //y=7.4 //x2=56.24 //y2=7.4
r1655 (  95 97 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=56.24 //y=7.4 //x2=57.35 //y2=7.4
r1656 (  93 859 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=55.13 //y=7.4 //x2=55.13 //y2=7.4
r1657 (  93 95 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=55.13 //y=7.4 //x2=56.24 //y2=7.4
r1658 (  91 856 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=53.65 //y=7.4 //x2=53.65 //y2=7.4
r1659 (  91 93 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=53.65 //y=7.4 //x2=55.13 //y2=7.4
r1660 (  89 620 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=52.54 //y=7.4 //x2=52.54 //y2=7.4
r1661 (  89 91 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=52.54 //y=7.4 //x2=53.65 //y2=7.4
r1662 (  87 610 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=51.43 //y=7.4 //x2=51.43 //y2=7.4
r1663 (  87 89 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=51.43 //y=7.4 //x2=52.54 //y2=7.4
r1664 (  85 596 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=49.95 //y=7.4 //x2=49.95 //y2=7.4
r1665 (  85 87 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=49.95 //y=7.4 //x2=51.43 //y2=7.4
r1666 (  83 586 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=48.84 //y=7.4 //x2=48.84 //y2=7.4
r1667 (  83 85 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=48.84 //y=7.4 //x2=49.95 //y2=7.4
r1668 (  81 572 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=47.36 //y=7.4 //x2=47.36 //y2=7.4
r1669 (  81 83 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=47.36 //y=7.4 //x2=48.84 //y2=7.4
r1670 (  79 562 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=46.25 //y=7.4 //x2=46.25 //y2=7.4
r1671 (  79 81 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=46.25 //y=7.4 //x2=47.36 //y2=7.4
r1672 (  77 552 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=45.14 //y=7.4 //x2=45.14 //y2=7.4
r1673 (  77 79 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=45.14 //y=7.4 //x2=46.25 //y2=7.4
r1674 (  75 844 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=44.03 //y=7.4 //x2=44.03 //y2=7.4
r1675 (  75 77 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=44.03 //y=7.4 //x2=45.14 //y2=7.4
r1676 (  73 530 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=42.55 //y=7.4 //x2=42.55 //y2=7.4
r1677 (  73 75 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=42.55 //y=7.4 //x2=44.03 //y2=7.4
r1678 (  71 520 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=41.44 //y=7.4 //x2=41.44 //y2=7.4
r1679 (  71 73 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=41.44 //y=7.4 //x2=42.55 //y2=7.4
r1680 (  69 839 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=40.33 //y=7.4 //x2=40.33 //y2=7.4
r1681 (  69 71 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=40.33 //y=7.4 //x2=41.44 //y2=7.4
r1682 (  67 836 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=38.85 //y=7.4 //x2=38.85 //y2=7.4
r1683 (  67 69 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=38.85 //y=7.4 //x2=40.33 //y2=7.4
r1684 (  65 482 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37.74 //y=7.4 //x2=37.74 //y2=7.4
r1685 (  65 67 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=37.74 //y=7.4 //x2=38.85 //y2=7.4
r1686 (  62 472 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=36.63 //y=7.4 //x2=36.63 //y2=7.4
r1687 (  60 458 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.15 //y=7.4 //x2=35.15 //y2=7.4
r1688 (  60 62 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=35.15 //y=7.4 //x2=36.63 //y2=7.4
r1689 (  58 448 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.04 //y=7.4 //x2=34.04 //y2=7.4
r1690 (  58 60 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=34.04 //y=7.4 //x2=35.15 //y2=7.4
r1691 (  56 434 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.56 //y=7.4 //x2=32.56 //y2=7.4
r1692 (  56 58 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=32.56 //y=7.4 //x2=34.04 //y2=7.4
r1693 (  54 424 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.45 //y=7.4 //x2=31.45 //y2=7.4
r1694 (  54 56 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.45 //y=7.4 //x2=32.56 //y2=7.4
r1695 (  52 825 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=30.34 //y=7.4 //x2=30.34 //y2=7.4
r1696 (  52 54 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=30.34 //y=7.4 //x2=31.45 //y2=7.4
r1697 (  50 822 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.86 //y=7.4 //x2=28.86 //y2=7.4
r1698 (  50 52 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=28.86 //y=7.4 //x2=30.34 //y2=7.4
r1699 (  48 386 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.75 //y=7.4 //x2=27.75 //y2=7.4
r1700 (  48 50 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=27.75 //y=7.4 //x2=28.86 //y2=7.4
r1701 (  46 376 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=26.64 //y=7.4 //x2=26.64 //y2=7.4
r1702 (  46 48 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=26.64 //y=7.4 //x2=27.75 //y2=7.4
r1703 (  44 817 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.16 //y=7.4 //x2=25.16 //y2=7.4
r1704 (  44 46 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=25.16 //y=7.4 //x2=26.64 //y2=7.4
r1705 (  42 354 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.05 //y=7.4 //x2=24.05 //y2=7.4
r1706 (  42 44 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=24.05 //y=7.4 //x2=25.16 //y2=7.4
r1707 (  40 344 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.94 //y=7.4 //x2=22.94 //y2=7.4
r1708 (  40 42 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.94 //y=7.4 //x2=24.05 //y2=7.4
r1709 (  38 334 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.83 //y=7.4 //x2=21.83 //y2=7.4
r1710 (  38 40 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.83 //y=7.4 //x2=22.94 //y2=7.4
r1711 (  36 320 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=7.4 //x2=20.35 //y2=7.4
r1712 (  36 38 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=7.4 //x2=21.83 //y2=7.4
r1713 (  34 310 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.24 //y=7.4 //x2=19.24 //y2=7.4
r1714 (  34 36 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.24 //y=7.4 //x2=20.35 //y2=7.4
r1715 (  32 296 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=7.4 //x2=17.76 //y2=7.4
r1716 (  32 34 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=7.4 //x2=19.24 //y2=7.4
r1717 (  30 286 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=7.4 //x2=16.65 //y2=7.4
r1718 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=7.4 //x2=17.76 //y2=7.4
r1719 (  28 805 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.54 //y=7.4 //x2=15.54 //y2=7.4
r1720 (  28 30 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.54 //y=7.4 //x2=16.65 //y2=7.4
r1721 (  26 802 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=7.4 //x2=14.06 //y2=7.4
r1722 (  26 28 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=7.4 //x2=15.54 //y2=7.4
r1723 (  24 248 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.95 //y=7.4 //x2=12.95 //y2=7.4
r1724 (  24 26 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.95 //y=7.4 //x2=14.06 //y2=7.4
r1725 (  22 238 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.84 //y=7.4 //x2=11.84 //y2=7.4
r1726 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.84 //y=7.4 //x2=12.95 //y2=7.4
r1727 (  20 224 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r1728 (  20 22 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=7.4 //x2=11.84 //y2=7.4
r1729 (  18 214 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=7.4 //x2=9.25 //y2=7.4
r1730 (  18 20 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=7.4 //x2=10.36 //y2=7.4
r1731 (  16 200 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=7.4 //x2=7.77 //y2=7.4
r1732 (  16 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=7.4 //x2=9.25 //y2=7.4
r1733 (  14 190 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r1734 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.4 //x2=7.77 //y2=7.4
r1735 (  12 791 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r1736 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.66 //y2=7.4
r1737 (  10 168 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=7.4 //x2=4.07 //y2=7.4
r1738 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=7.4 //x2=5.55 //y2=7.4
r1739 (  8 158 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r1740 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r1741 (  6 140 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r1742 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r1743 (  3 130 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r1744 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r1745 (  1 65 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=37.185 //y=7.4 //x2=37.74 //y2=7.4
r1746 (  1 62 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=37.185 //y=7.4 //x2=36.63 //y2=7.4
ends PM_TMRDFFQNX1\%VDD

subckt PM_TMRDFFQNX1\%noxref_3 ( 1 2 3 4 12 25 26 37 39 40 44 46 53 54 55 56 \
 57 58 59 63 64 65 70 72 75 76 77 78 79 80 84 86 89 90 95 96 101 110 113 115 \
 116 )
c232 ( 116 0 ) capacitor c=0.0220291f //x=6.775 //y=5.02
c233 ( 115 0 ) capacitor c=0.0217503f //x=5.895 //y=5.02
c234 ( 113 0 ) capacitor c=0.00866655f //x=6.77 //y=0.905
c235 ( 110 0 ) capacitor c=0.0588816f //x=9.25 //y=4.7
c236 ( 101 0 ) capacitor c=0.058931f //x=3.33 //y=4.7
c237 ( 96 0 ) capacitor c=0.0273931f //x=3.33 //y=1.915
c238 ( 95 0 ) capacitor c=0.0464411f //x=3.33 //y=2.08
c239 ( 90 0 ) capacitor c=0.0318948f //x=9.585 //y=1.21
c240 ( 89 0 ) capacitor c=0.0187384f //x=9.585 //y=0.865
c241 ( 86 0 ) capacitor c=0.0141798f //x=9.43 //y=1.365
c242 ( 84 0 ) capacitor c=0.0149844f //x=9.43 //y=0.71
c243 ( 80 0 ) capacitor c=0.0816311f //x=9.055 //y=1.915
c244 ( 79 0 ) capacitor c=0.0229722f //x=9.055 //y=1.52
c245 ( 78 0 ) capacitor c=0.0234352f //x=9.055 //y=1.21
c246 ( 77 0 ) capacitor c=0.0199343f //x=9.055 //y=0.865
c247 ( 76 0 ) capacitor c=0.0432517f //x=3.85 //y=1.26
c248 ( 75 0 ) capacitor c=0.0200379f //x=3.85 //y=0.915
c249 ( 72 0 ) capacitor c=0.0158629f //x=3.695 //y=1.415
c250 ( 70 0 ) capacitor c=0.0157803f //x=3.695 //y=0.76
c251 ( 65 0 ) capacitor c=0.0218028f //x=3.32 //y=1.57
c252 ( 64 0 ) capacitor c=0.0207459f //x=3.32 //y=1.26
c253 ( 63 0 ) capacitor c=0.0194308f //x=3.32 //y=0.915
c254 ( 59 0 ) capacitor c=0.110275f //x=9.59 //y=6.02
c255 ( 58 0 ) capacitor c=0.154305f //x=9.15 //y=6.02
c256 ( 57 0 ) capacitor c=0.158794f //x=3.51 //y=6.02
c257 ( 56 0 ) capacitor c=0.110114f //x=3.07 //y=6.02
c258 ( 53 0 ) capacitor c=0.00211606f //x=6.92 //y=5.2
c259 ( 46 0 ) capacitor c=0.0894554f //x=9.25 //y=2.08
c260 ( 44 0 ) capacitor c=0.106205f //x=7.4 //y=3.33
c261 ( 40 0 ) capacitor c=0.00436419f //x=7.045 //y=1.655
c262 ( 39 0 ) capacitor c=0.0127039f //x=7.315 //y=1.655
c263 ( 37 0 ) capacitor c=0.0137522f //x=7.315 //y=5.2
c264 ( 26 0 ) capacitor c=0.00251635f //x=6.125 //y=5.2
c265 ( 25 0 ) capacitor c=0.0142423f //x=6.835 //y=5.2
c266 ( 12 0 ) capacitor c=0.0882402f //x=3.33 //y=2.08
c267 ( 4 0 ) capacitor c=0.00305824f //x=7.515 //y=3.33
c268 ( 3 0 ) capacitor c=0.0402189f //x=9.135 //y=3.33
c269 ( 2 0 ) capacitor c=0.0149802f //x=3.445 //y=3.33
c270 ( 1 0 ) capacitor c=0.100545f //x=7.285 //y=3.33
r271 (  108 110 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=9.15 //y=4.7 //x2=9.25 //y2=4.7
r272 (  95 96 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.33 //y=2.08 //x2=3.33 //y2=1.915
r273 (  91 110 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=9.59 //y=4.865 //x2=9.25 //y2=4.7
r274 (  90 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.585 //y=1.21 //x2=9.545 //y2=1.365
r275 (  89 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.585 //y=0.865 //x2=9.545 //y2=0.71
r276 (  89 90 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.585 //y=0.865 //x2=9.585 //y2=1.21
r277 (  87 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.21 //y=1.365 //x2=9.095 //y2=1.365
r278 (  86 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.43 //y=1.365 //x2=9.545 //y2=1.365
r279 (  85 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.21 //y=0.71 //x2=9.095 //y2=0.71
r280 (  84 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.43 //y=0.71 //x2=9.545 //y2=0.71
r281 (  84 85 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=9.43 //y=0.71 //x2=9.21 //y2=0.71
r282 (  81 108 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=9.15 //y=4.865 //x2=9.15 //y2=4.7
r283 (  80 105 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=9.055 //y=1.915 //x2=9.25 //y2=2.08
r284 (  79 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.055 //y=1.52 //x2=9.095 //y2=1.365
r285 (  79 80 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=9.055 //y=1.52 //x2=9.055 //y2=1.915
r286 (  78 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.055 //y=1.21 //x2=9.095 //y2=1.365
r287 (  77 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.055 //y=0.865 //x2=9.095 //y2=0.71
r288 (  77 78 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.055 //y=0.865 //x2=9.055 //y2=1.21
r289 (  76 103 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=1.26 //x2=3.81 //y2=1.415
r290 (  75 102 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.81 //y2=0.76
r291 (  75 76 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.85 //y2=1.26
r292 (  73 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=1.415 //x2=3.36 //y2=1.415
r293 (  72 103 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=1.415 //x2=3.81 //y2=1.415
r294 (  71 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=0.76 //x2=3.36 //y2=0.76
r295 (  70 102 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.81 //y2=0.76
r296 (  70 71 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.475 //y2=0.76
r297 (  67 101 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=3.51 //y=4.865 //x2=3.33 //y2=4.7
r298 (  65 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.36 //y2=1.415
r299 (  65 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.32 //y2=1.915
r300 (  64 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.26 //x2=3.36 //y2=1.415
r301 (  63 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.36 //y2=0.76
r302 (  63 64 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.32 //y2=1.26
r303 (  60 101 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=3.07 //y=4.865 //x2=3.33 //y2=4.7
r304 (  59 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.59 //y=6.02 //x2=9.59 //y2=4.865
r305 (  58 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.15 //y=6.02 //x2=9.15 //y2=4.865
r306 (  57 67 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.51 //y=6.02 //x2=3.51 //y2=4.865
r307 (  56 60 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.07 //y=6.02 //x2=3.07 //y2=4.865
r308 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.32 //y=1.365 //x2=9.43 //y2=1.365
r309 (  55 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.32 //y=1.365 //x2=9.21 //y2=1.365
r310 (  54 72 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.695 //y2=1.415
r311 (  54 73 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.475 //y2=1.415
r312 (  51 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=4.7 //x2=9.25 //y2=4.7
r313 (  49 51 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=9.25 //y=3.33 //x2=9.25 //y2=4.7
r314 (  46 105 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=2.08 //x2=9.25 //y2=2.08
r315 (  46 49 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=9.25 //y=2.08 //x2=9.25 //y2=3.33
r316 (  42 44 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=7.4 //y=5.115 //x2=7.4 //y2=3.33
r317 (  41 44 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=7.4 //y=1.74 //x2=7.4 //y2=3.33
r318 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.655 //x2=7.4 //y2=1.74
r319 (  39 40 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.655 //x2=7.045 //y2=1.655
r320 (  38 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.005 //y=5.2 //x2=6.92 //y2=5.2
r321 (  37 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.2 //x2=7.4 //y2=5.115
r322 (  37 38 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.2 //x2=7.005 //y2=5.2
r323 (  33 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.96 //y=1.57 //x2=7.045 //y2=1.655
r324 (  33 113 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=6.96 //y=1.57 //x2=6.96 //y2=1
r325 (  27 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.92 //y=5.285 //x2=6.92 //y2=5.2
r326 (  27 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=6.92 //y=5.285 //x2=6.92 //y2=5.725
r327 (  25 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.835 //y=5.2 //x2=6.92 //y2=5.2
r328 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=6.835 //y=5.2 //x2=6.125 //y2=5.2
r329 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.04 //y=5.285 //x2=6.125 //y2=5.2
r330 (  19 115 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=6.04 //y=5.285 //x2=6.04 //y2=5.725
r331 (  17 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r332 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=3.33 //x2=3.33 //y2=4.7
r333 (  12 95 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r334 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.08 //x2=3.33 //y2=3.33
r335 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.25 //y=3.33 //x2=9.25 //y2=3.33
r336 (  8 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=7.4 \
 //y=3.33 //x2=7.4 //y2=3.33
r337 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=3.33 //x2=3.33 //y2=3.33
r338 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.515 //y=3.33 //x2=7.4 //y2=3.33
r339 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.135 //y=3.33 //x2=9.25 //y2=3.33
r340 (  3 4 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=9.135 //y=3.33 //x2=7.515 //y2=3.33
r341 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.445 //y=3.33 //x2=3.33 //y2=3.33
r342 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.285 //y=3.33 //x2=7.4 //y2=3.33
r343 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=7.285 //y=3.33 //x2=3.445 //y2=3.33
ends PM_TMRDFFQNX1\%noxref_3

subckt PM_TMRDFFQNX1\%noxref_4 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 \
 48 52 54 57 58 68 71 73 74 )
c150 ( 74 0 ) capacitor c=0.0220291f //x=10.105 //y=5.02
c151 ( 73 0 ) capacitor c=0.0217503f //x=9.225 //y=5.02
c152 ( 71 0 ) capacitor c=0.00866655f //x=10.1 //y=0.905
c153 ( 68 0 ) capacitor c=0.0588816f //x=12.58 //y=4.7
c154 ( 58 0 ) capacitor c=0.0318948f //x=12.915 //y=1.21
c155 ( 57 0 ) capacitor c=0.0187384f //x=12.915 //y=0.865
c156 ( 54 0 ) capacitor c=0.0141798f //x=12.76 //y=1.365
c157 ( 52 0 ) capacitor c=0.0149844f //x=12.76 //y=0.71
c158 ( 48 0 ) capacitor c=0.0816311f //x=12.385 //y=1.915
c159 ( 47 0 ) capacitor c=0.0229722f //x=12.385 //y=1.52
c160 ( 46 0 ) capacitor c=0.0234352f //x=12.385 //y=1.21
c161 ( 45 0 ) capacitor c=0.0199343f //x=12.385 //y=0.865
c162 ( 44 0 ) capacitor c=0.110275f //x=12.92 //y=6.02
c163 ( 43 0 ) capacitor c=0.154305f //x=12.48 //y=6.02
c164 ( 41 0 ) capacitor c=0.00211606f //x=10.25 //y=5.2
c165 ( 34 0 ) capacitor c=0.0889544f //x=12.58 //y=2.08
c166 ( 32 0 ) capacitor c=0.106752f //x=10.73 //y=3.33
c167 ( 28 0 ) capacitor c=0.00436419f //x=10.375 //y=1.655
c168 ( 27 0 ) capacitor c=0.0127039f //x=10.645 //y=1.655
c169 ( 25 0 ) capacitor c=0.0137522f //x=10.645 //y=5.2
c170 ( 14 0 ) capacitor c=0.00251459f //x=9.455 //y=5.2
c171 ( 13 0 ) capacitor c=0.0143649f //x=10.165 //y=5.2
c172 ( 2 0 ) capacitor c=0.00703116f //x=10.845 //y=3.33
c173 ( 1 0 ) capacitor c=0.0455801f //x=12.465 //y=3.33
r174 (  66 68 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=12.48 //y=4.7 //x2=12.58 //y2=4.7
r175 (  59 68 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=12.92 //y=4.865 //x2=12.58 //y2=4.7
r176 (  58 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.915 //y=1.21 //x2=12.875 //y2=1.365
r177 (  57 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.915 //y=0.865 //x2=12.875 //y2=0.71
r178 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.915 //y=0.865 //x2=12.915 //y2=1.21
r179 (  55 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.54 //y=1.365 //x2=12.425 //y2=1.365
r180 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.76 //y=1.365 //x2=12.875 //y2=1.365
r181 (  53 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.54 //y=0.71 //x2=12.425 //y2=0.71
r182 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.76 //y=0.71 //x2=12.875 //y2=0.71
r183 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=12.76 //y=0.71 //x2=12.54 //y2=0.71
r184 (  49 66 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=12.48 //y=4.865 //x2=12.48 //y2=4.7
r185 (  48 63 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=12.385 //y=1.915 //x2=12.58 //y2=2.08
r186 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.385 //y=1.52 //x2=12.425 //y2=1.365
r187 (  47 48 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=12.385 //y=1.52 //x2=12.385 //y2=1.915
r188 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.385 //y=1.21 //x2=12.425 //y2=1.365
r189 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.385 //y=0.865 //x2=12.425 //y2=0.71
r190 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.385 //y=0.865 //x2=12.385 //y2=1.21
r191 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.92 //y=6.02 //x2=12.92 //y2=4.865
r192 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.48 //y=6.02 //x2=12.48 //y2=4.865
r193 (  42 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.65 //y=1.365 //x2=12.76 //y2=1.365
r194 (  42 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.65 //y=1.365 //x2=12.54 //y2=1.365
r195 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.58 //y=4.7 //x2=12.58 //y2=4.7
r196 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=12.58 //y=3.33 //x2=12.58 //y2=4.7
r197 (  34 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.58 //y=2.08 //x2=12.58 //y2=2.08
r198 (  34 37 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=12.58 //y=2.08 //x2=12.58 //y2=3.33
r199 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=10.73 //y=5.115 //x2=10.73 //y2=3.33
r200 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=10.73 //y=1.74 //x2=10.73 //y2=3.33
r201 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.645 //y=1.655 //x2=10.73 //y2=1.74
r202 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=10.645 //y=1.655 //x2=10.375 //y2=1.655
r203 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.335 //y=5.2 //x2=10.25 //y2=5.2
r204 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.645 //y=5.2 //x2=10.73 //y2=5.115
r205 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=10.645 //y=5.2 //x2=10.335 //y2=5.2
r206 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.29 //y=1.57 //x2=10.375 //y2=1.655
r207 (  21 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=10.29 //y=1.57 //x2=10.29 //y2=1
r208 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.25 //y=5.285 //x2=10.25 //y2=5.2
r209 (  15 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=10.25 //y=5.285 //x2=10.25 //y2=5.725
r210 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.165 //y=5.2 //x2=10.25 //y2=5.2
r211 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.165 //y=5.2 //x2=9.455 //y2=5.2
r212 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.37 //y=5.285 //x2=9.455 //y2=5.2
r213 (  7 73 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=9.37 //y=5.285 //x2=9.37 //y2=5.725
r214 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.58 //y=3.33 //x2=12.58 //y2=3.33
r215 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.73 //y=3.33 //x2=10.73 //y2=3.33
r216 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.845 //y=3.33 //x2=10.73 //y2=3.33
r217 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.465 //y=3.33 //x2=12.58 //y2=3.33
r218 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=12.465 //y=3.33 //x2=10.845 //y2=3.33
ends PM_TMRDFFQNX1\%noxref_4

subckt PM_TMRDFFQNX1\%noxref_5 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 63 \
 64 65 66 67 68 69 70 71 72 76 78 81 82 86 87 88 89 93 95 98 99 109 118 121 \
 123 124 125 )
c248 ( 125 0 ) capacitor c=0.023087f //x=3.145 //y=5.02
c249 ( 124 0 ) capacitor c=0.023519f //x=2.265 //y=5.02
c250 ( 123 0 ) capacitor c=0.0224735f //x=1.385 //y=5.02
c251 ( 121 0 ) capacitor c=0.00872971f //x=3.395 //y=0.915
c252 ( 118 0 ) capacitor c=0.0588845f //x=15.91 //y=4.7
c253 ( 109 0 ) capacitor c=0.0588816f //x=5.92 //y=4.7
c254 ( 99 0 ) capacitor c=0.0318948f //x=16.245 //y=1.21
c255 ( 98 0 ) capacitor c=0.0187384f //x=16.245 //y=0.865
c256 ( 95 0 ) capacitor c=0.0141798f //x=16.09 //y=1.365
c257 ( 93 0 ) capacitor c=0.0149844f //x=16.09 //y=0.71
c258 ( 89 0 ) capacitor c=0.0816311f //x=15.715 //y=1.915
c259 ( 88 0 ) capacitor c=0.0229722f //x=15.715 //y=1.52
c260 ( 87 0 ) capacitor c=0.0234352f //x=15.715 //y=1.21
c261 ( 86 0 ) capacitor c=0.0199343f //x=15.715 //y=0.865
c262 ( 82 0 ) capacitor c=0.0318948f //x=6.255 //y=1.21
c263 ( 81 0 ) capacitor c=0.0187384f //x=6.255 //y=0.865
c264 ( 78 0 ) capacitor c=0.0141798f //x=6.1 //y=1.365
c265 ( 76 0 ) capacitor c=0.0149844f //x=6.1 //y=0.71
c266 ( 72 0 ) capacitor c=0.0860049f //x=5.725 //y=1.915
c267 ( 71 0 ) capacitor c=0.0229722f //x=5.725 //y=1.52
c268 ( 70 0 ) capacitor c=0.0234352f //x=5.725 //y=1.21
c269 ( 69 0 ) capacitor c=0.0199343f //x=5.725 //y=0.865
c270 ( 68 0 ) capacitor c=0.110275f //x=16.25 //y=6.02
c271 ( 67 0 ) capacitor c=0.154305f //x=15.81 //y=6.02
c272 ( 66 0 ) capacitor c=0.110275f //x=6.26 //y=6.02
c273 ( 65 0 ) capacitor c=0.154305f //x=5.82 //y=6.02
c274 ( 62 0 ) capacitor c=0.00106608f //x=3.29 //y=5.155
c275 ( 61 0 ) capacitor c=0.00207162f //x=2.41 //y=5.155
c276 ( 54 0 ) capacitor c=0.0918023f //x=15.91 //y=2.08
c277 ( 46 0 ) capacitor c=0.0905231f //x=5.92 //y=2.08
c278 ( 44 0 ) capacitor c=0.109488f //x=4.07 //y=3.7
c279 ( 40 0 ) capacitor c=0.00493499f //x=3.67 //y=1.665
c280 ( 39 0 ) capacitor c=0.0154052f //x=3.985 //y=1.665
c281 ( 33 0 ) capacitor c=0.0284988f //x=3.985 //y=5.155
c282 ( 25 0 ) capacitor c=0.0176454f //x=3.205 //y=5.155
c283 ( 18 0 ) capacitor c=0.00351598f //x=1.615 //y=5.155
c284 ( 17 0 ) capacitor c=0.0154196f //x=2.325 //y=5.155
c285 ( 4 0 ) capacitor c=0.00424317f //x=6.035 //y=3.7
c286 ( 3 0 ) capacitor c=0.173045f //x=15.795 //y=3.7
c287 ( 2 0 ) capacitor c=0.0125346f //x=4.185 //y=3.7
c288 ( 1 0 ) capacitor c=0.0285004f //x=5.805 //y=3.7
r289 (  116 118 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=15.81 //y=4.7 //x2=15.91 //y2=4.7
r290 (  107 109 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=5.82 //y=4.7 //x2=5.92 //y2=4.7
r291 (  100 118 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=16.25 //y=4.865 //x2=15.91 //y2=4.7
r292 (  99 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.245 //y=1.21 //x2=16.205 //y2=1.365
r293 (  98 119 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.245 //y=0.865 //x2=16.205 //y2=0.71
r294 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.245 //y=0.865 //x2=16.245 //y2=1.21
r295 (  96 115 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.87 //y=1.365 //x2=15.755 //y2=1.365
r296 (  95 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.09 //y=1.365 //x2=16.205 //y2=1.365
r297 (  94 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.87 //y=0.71 //x2=15.755 //y2=0.71
r298 (  93 119 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.09 //y=0.71 //x2=16.205 //y2=0.71
r299 (  93 94 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=16.09 //y=0.71 //x2=15.87 //y2=0.71
r300 (  90 116 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=15.81 //y=4.865 //x2=15.81 //y2=4.7
r301 (  89 113 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=15.715 //y=1.915 //x2=15.91 //y2=2.08
r302 (  88 115 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.715 //y=1.52 //x2=15.755 //y2=1.365
r303 (  88 89 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=15.715 //y=1.52 //x2=15.715 //y2=1.915
r304 (  87 115 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.715 //y=1.21 //x2=15.755 //y2=1.365
r305 (  86 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.715 //y=0.865 //x2=15.755 //y2=0.71
r306 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.715 //y=0.865 //x2=15.715 //y2=1.21
r307 (  83 109 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=6.26 //y=4.865 //x2=5.92 //y2=4.7
r308 (  82 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.255 //y=1.21 //x2=6.215 //y2=1.365
r309 (  81 110 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.255 //y=0.865 //x2=6.215 //y2=0.71
r310 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.255 //y=0.865 //x2=6.255 //y2=1.21
r311 (  79 106 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.88 //y=1.365 //x2=5.765 //y2=1.365
r312 (  78 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.1 //y=1.365 //x2=6.215 //y2=1.365
r313 (  77 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.88 //y=0.71 //x2=5.765 //y2=0.71
r314 (  76 110 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.1 //y=0.71 //x2=6.215 //y2=0.71
r315 (  76 77 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=6.1 //y=0.71 //x2=5.88 //y2=0.71
r316 (  73 107 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=5.82 //y=4.865 //x2=5.82 //y2=4.7
r317 (  72 104 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=5.725 //y=1.915 //x2=5.92 //y2=2.08
r318 (  71 106 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.725 //y=1.52 //x2=5.765 //y2=1.365
r319 (  71 72 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=5.725 //y=1.52 //x2=5.725 //y2=1.915
r320 (  70 106 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.725 //y=1.21 //x2=5.765 //y2=1.365
r321 (  69 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.725 //y=0.865 //x2=5.765 //y2=0.71
r322 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.725 //y=0.865 //x2=5.725 //y2=1.21
r323 (  68 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.25 //y=6.02 //x2=16.25 //y2=4.865
r324 (  67 90 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.81 //y=6.02 //x2=15.81 //y2=4.865
r325 (  66 83 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.26 //y=6.02 //x2=6.26 //y2=4.865
r326 (  65 73 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.82 //y=6.02 //x2=5.82 //y2=4.865
r327 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.98 //y=1.365 //x2=16.09 //y2=1.365
r328 (  64 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.98 //y=1.365 //x2=15.87 //y2=1.365
r329 (  63 78 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.99 //y=1.365 //x2=6.1 //y2=1.365
r330 (  63 79 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.99 //y=1.365 //x2=5.88 //y2=1.365
r331 (  59 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.91 //y=4.7 //x2=15.91 //y2=4.7
r332 (  57 59 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=15.91 //y=3.7 //x2=15.91 //y2=4.7
r333 (  54 113 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.91 //y=2.08 //x2=15.91 //y2=2.08
r334 (  54 57 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=15.91 //y=2.08 //x2=15.91 //y2=3.7
r335 (  51 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=4.7 //x2=5.92 //y2=4.7
r336 (  49 51 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=5.92 //y=3.7 //x2=5.92 //y2=4.7
r337 (  46 104 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=2.08 //x2=5.92 //y2=2.08
r338 (  46 49 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.08 //x2=5.92 //y2=3.7
r339 (  42 44 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=4.07 //y=5.07 //x2=4.07 //y2=3.7
r340 (  41 44 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=4.07 //y=1.75 //x2=4.07 //y2=3.7
r341 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=4.07 //y2=1.75
r342 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=3.67 //y2=1.665
r343 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.67 //y2=1.665
r344 (  35 121 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.585 //y2=1.01
r345 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.375 //y=5.155 //x2=3.29 //y2=5.155
r346 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=4.07 //y2=5.07
r347 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=3.375 //y2=5.155
r348 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.155
r349 (  27 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.725
r350 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.495 //y=5.155 //x2=2.41 //y2=5.155
r351 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=3.29 //y2=5.155
r352 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=2.495 //y2=5.155
r353 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.155
r354 (  19 124 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.725
r355 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=2.41 //y2=5.155
r356 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=1.615 //y2=5.155
r357 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.615 //y2=5.155
r358 (  11 123 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.53 //y2=5.725
r359 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.91 //y=3.7 //x2=15.91 //y2=3.7
r360 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.92 //y=3.7 //x2=5.92 //y2=3.7
r361 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=3.7 //x2=4.07 //y2=3.7
r362 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.035 //y=3.7 //x2=5.92 //y2=3.7
r363 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.795 //y=3.7 //x2=15.91 //y2=3.7
r364 (  3 4 ) resistor r=9.31298 //w=0.131 //l=9.76 //layer=m1 \
 //thickness=0.36 //x=15.795 //y=3.7 //x2=6.035 //y2=3.7
r365 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.185 //y=3.7 //x2=4.07 //y2=3.7
r366 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.805 //y=3.7 //x2=5.92 //y2=3.7
r367 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=5.805 //y=3.7 //x2=4.185 //y2=3.7
ends PM_TMRDFFQNX1\%noxref_5

subckt PM_TMRDFFQNX1\%noxref_6 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 \
 48 52 54 57 58 68 71 73 74 )
c150 ( 74 0 ) capacitor c=0.0220291f //x=16.765 //y=5.02
c151 ( 73 0 ) capacitor c=0.0217503f //x=15.885 //y=5.02
c152 ( 71 0 ) capacitor c=0.00866655f //x=16.76 //y=0.905
c153 ( 68 0 ) capacitor c=0.0588816f //x=19.24 //y=4.7
c154 ( 58 0 ) capacitor c=0.0318948f //x=19.575 //y=1.21
c155 ( 57 0 ) capacitor c=0.0187384f //x=19.575 //y=0.865
c156 ( 54 0 ) capacitor c=0.0141798f //x=19.42 //y=1.365
c157 ( 52 0 ) capacitor c=0.0149844f //x=19.42 //y=0.71
c158 ( 48 0 ) capacitor c=0.0816311f //x=19.045 //y=1.915
c159 ( 47 0 ) capacitor c=0.0229722f //x=19.045 //y=1.52
c160 ( 46 0 ) capacitor c=0.0234352f //x=19.045 //y=1.21
c161 ( 45 0 ) capacitor c=0.0199343f //x=19.045 //y=0.865
c162 ( 44 0 ) capacitor c=0.110275f //x=19.58 //y=6.02
c163 ( 43 0 ) capacitor c=0.154305f //x=19.14 //y=6.02
c164 ( 41 0 ) capacitor c=0.00211606f //x=16.91 //y=5.2
c165 ( 34 0 ) capacitor c=0.0889334f //x=19.24 //y=2.08
c166 ( 32 0 ) capacitor c=0.10676f //x=17.39 //y=3.7
c167 ( 28 0 ) capacitor c=0.00436419f //x=17.035 //y=1.655
c168 ( 27 0 ) capacitor c=0.0127039f //x=17.305 //y=1.655
c169 ( 25 0 ) capacitor c=0.0137522f //x=17.305 //y=5.2
c170 ( 14 0 ) capacitor c=0.0025165f //x=16.115 //y=5.2
c171 ( 13 0 ) capacitor c=0.0142497f //x=16.825 //y=5.2
c172 ( 2 0 ) capacitor c=0.00701934f //x=17.505 //y=3.7
c173 ( 1 0 ) capacitor c=0.0472012f //x=19.125 //y=3.7
r174 (  66 68 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=19.14 //y=4.7 //x2=19.24 //y2=4.7
r175 (  59 68 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=19.58 //y=4.865 //x2=19.24 //y2=4.7
r176 (  58 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.575 //y=1.21 //x2=19.535 //y2=1.365
r177 (  57 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.575 //y=0.865 //x2=19.535 //y2=0.71
r178 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=19.575 //y=0.865 //x2=19.575 //y2=1.21
r179 (  55 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.2 //y=1.365 //x2=19.085 //y2=1.365
r180 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.42 //y=1.365 //x2=19.535 //y2=1.365
r181 (  53 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.2 //y=0.71 //x2=19.085 //y2=0.71
r182 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.42 //y=0.71 //x2=19.535 //y2=0.71
r183 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=19.42 //y=0.71 //x2=19.2 //y2=0.71
r184 (  49 66 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=19.14 //y=4.865 //x2=19.14 //y2=4.7
r185 (  48 63 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=19.045 //y=1.915 //x2=19.24 //y2=2.08
r186 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.045 //y=1.52 //x2=19.085 //y2=1.365
r187 (  47 48 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=19.045 //y=1.52 //x2=19.045 //y2=1.915
r188 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.045 //y=1.21 //x2=19.085 //y2=1.365
r189 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.045 //y=0.865 //x2=19.085 //y2=0.71
r190 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=19.045 //y=0.865 //x2=19.045 //y2=1.21
r191 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.58 //y=6.02 //x2=19.58 //y2=4.865
r192 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.14 //y=6.02 //x2=19.14 //y2=4.865
r193 (  42 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=19.31 //y=1.365 //x2=19.42 //y2=1.365
r194 (  42 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=19.31 //y=1.365 //x2=19.2 //y2=1.365
r195 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.24 //y=4.7 //x2=19.24 //y2=4.7
r196 (  37 39 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=19.24 //y=3.7 //x2=19.24 //y2=4.7
r197 (  34 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.24 //y=2.08 //x2=19.24 //y2=2.08
r198 (  34 37 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=19.24 //y=2.08 //x2=19.24 //y2=3.7
r199 (  30 32 ) resistor r=96.8556 //w=0.187 //l=1.415 //layer=li \
 //thickness=0.1 //x=17.39 //y=5.115 //x2=17.39 //y2=3.7
r200 (  29 32 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=17.39 //y=1.74 //x2=17.39 //y2=3.7
r201 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.305 //y=1.655 //x2=17.39 //y2=1.74
r202 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=17.305 //y=1.655 //x2=17.035 //y2=1.655
r203 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.995 //y=5.2 //x2=16.91 //y2=5.2
r204 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.305 //y=5.2 //x2=17.39 //y2=5.115
r205 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=17.305 //y=5.2 //x2=16.995 //y2=5.2
r206 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.95 //y=1.57 //x2=17.035 //y2=1.655
r207 (  21 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=16.95 //y=1.57 //x2=16.95 //y2=1
r208 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.91 //y=5.285 //x2=16.91 //y2=5.2
r209 (  15 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=16.91 //y=5.285 //x2=16.91 //y2=5.725
r210 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.825 //y=5.2 //x2=16.91 //y2=5.2
r211 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=16.825 //y=5.2 //x2=16.115 //y2=5.2
r212 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.03 //y=5.285 //x2=16.115 //y2=5.2
r213 (  7 73 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=16.03 //y=5.285 //x2=16.03 //y2=5.725
r214 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=19.24 //y=3.7 //x2=19.24 //y2=3.7
r215 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.39 //y=3.7 //x2=17.39 //y2=3.7
r216 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.505 //y=3.7 //x2=17.39 //y2=3.7
r217 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=19.125 //y=3.7 //x2=19.24 //y2=3.7
r218 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=19.125 //y=3.7 //x2=17.505 //y2=3.7
ends PM_TMRDFFQNX1\%noxref_6

subckt PM_TMRDFFQNX1\%noxref_7 ( 1 2 3 4 5 6 16 23 25 35 36 47 49 50 54 55 57 \
 63 66 67 68 69 70 71 72 73 74 75 76 77 78 79 81 87 88 89 90 94 95 96 101 103 \
 105 111 112 113 114 115 120 122 124 130 131 141 142 145 154 155 158 166 168 \
 169 )
c353 ( 169 0 ) capacitor c=0.0220291f //x=13.435 //y=5.02
c354 ( 168 0 ) capacitor c=0.0217503f //x=12.555 //y=5.02
c355 ( 166 0 ) capacitor c=0.00866655f //x=13.43 //y=0.905
c356 ( 158 0 ) capacitor c=0.0331095f //x=20.01 //y=4.7
c357 ( 155 0 ) capacitor c=0.0279499f //x=19.98 //y=1.915
c358 ( 154 0 ) capacitor c=0.0421302f //x=19.98 //y=2.08
c359 ( 145 0 ) capacitor c=0.0331095f //x=10.02 //y=4.7
c360 ( 142 0 ) capacitor c=0.0279499f //x=9.99 //y=1.915
c361 ( 141 0 ) capacitor c=0.0421302f //x=9.99 //y=2.08
c362 ( 131 0 ) capacitor c=0.0429696f //x=20.545 //y=1.25
c363 ( 130 0 ) capacitor c=0.0192208f //x=20.545 //y=0.905
c364 ( 124 0 ) capacitor c=0.0158629f //x=20.39 //y=1.405
c365 ( 122 0 ) capacitor c=0.0157803f //x=20.39 //y=0.75
c366 ( 120 0 ) capacitor c=0.0295235f //x=20.385 //y=4.79
c367 ( 115 0 ) capacitor c=0.0204188f //x=20.015 //y=1.56
c368 ( 114 0 ) capacitor c=0.0168481f //x=20.015 //y=1.25
c369 ( 113 0 ) capacitor c=0.0174783f //x=20.015 //y=0.905
c370 ( 112 0 ) capacitor c=0.0429696f //x=10.555 //y=1.25
c371 ( 111 0 ) capacitor c=0.0192208f //x=10.555 //y=0.905
c372 ( 105 0 ) capacitor c=0.0158629f //x=10.4 //y=1.405
c373 ( 103 0 ) capacitor c=0.0157803f //x=10.4 //y=0.75
c374 ( 101 0 ) capacitor c=0.0295235f //x=10.395 //y=4.79
c375 ( 96 0 ) capacitor c=0.0204188f //x=10.025 //y=1.56
c376 ( 95 0 ) capacitor c=0.0168481f //x=10.025 //y=1.25
c377 ( 94 0 ) capacitor c=0.0174783f //x=10.025 //y=0.905
c378 ( 90 0 ) capacitor c=0.0559896f //x=1.385 //y=4.79
c379 ( 89 0 ) capacitor c=0.0298189f //x=1.675 //y=4.79
c380 ( 88 0 ) capacitor c=0.0347816f //x=1.34 //y=1.22
c381 ( 87 0 ) capacitor c=0.0187487f //x=1.34 //y=0.875
c382 ( 81 0 ) capacitor c=0.0137055f //x=1.185 //y=1.375
c383 ( 79 0 ) capacitor c=0.0149861f //x=1.185 //y=0.72
c384 ( 78 0 ) capacitor c=0.102158f //x=0.81 //y=1.915
c385 ( 77 0 ) capacitor c=0.0229444f //x=0.81 //y=1.53
c386 ( 76 0 ) capacitor c=0.0234352f //x=0.81 //y=1.22
c387 ( 75 0 ) capacitor c=0.0198724f //x=0.81 //y=0.875
c388 ( 74 0 ) capacitor c=0.15358f //x=20.46 //y=6.02
c389 ( 73 0 ) capacitor c=0.110281f //x=20.02 //y=6.02
c390 ( 72 0 ) capacitor c=0.15358f //x=10.47 //y=6.02
c391 ( 71 0 ) capacitor c=0.110281f //x=10.03 //y=6.02
c392 ( 70 0 ) capacitor c=0.110114f //x=1.75 //y=6.02
c393 ( 69 0 ) capacitor c=0.158956f //x=1.31 //y=6.02
c394 ( 63 0 ) capacitor c=0.0021186f //x=13.58 //y=5.2
c395 ( 57 0 ) capacitor c=0.0729826f //x=19.98 //y=2.08
c396 ( 55 0 ) capacitor c=0.00453889f //x=19.98 //y=4.535
c397 ( 54 0 ) capacitor c=0.108418f //x=14.06 //y=4.07
c398 ( 50 0 ) capacitor c=0.00436419f //x=13.705 //y=1.655
c399 ( 49 0 ) capacitor c=0.0127039f //x=13.975 //y=1.655
c400 ( 47 0 ) capacitor c=0.0137562f //x=13.975 //y=5.2
c401 ( 36 0 ) capacitor c=0.00251459f //x=12.785 //y=5.2
c402 ( 35 0 ) capacitor c=0.0142537f //x=13.495 //y=5.2
c403 ( 25 0 ) capacitor c=0.0719497f //x=9.99 //y=2.08
c404 ( 23 0 ) capacitor c=0.00453889f //x=9.99 //y=4.535
c405 ( 16 0 ) capacitor c=0.124161f //x=1.11 //y=2.08
c406 ( 6 0 ) capacitor c=0.00408661f //x=14.175 //y=4.07
c407 ( 5 0 ) capacitor c=0.100584f //x=19.865 //y=4.07
c408 ( 4 0 ) capacitor c=0.00412846f //x=10.105 //y=4.07
c409 ( 3 0 ) capacitor c=0.0519595f //x=13.945 //y=4.07
c410 ( 2 0 ) capacitor c=0.0160831f //x=1.225 //y=4.07
c411 ( 1 0 ) capacitor c=0.163286f //x=9.875 //y=4.07
r412 (  160 161 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=20.01 //y=4.79 //x2=20.01 //y2=4.865
r413 (  158 160 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=20.01 //y=4.7 //x2=20.01 //y2=4.79
r414 (  154 155 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=19.98 //y=2.08 //x2=19.98 //y2=1.915
r415 (  147 148 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=10.02 //y=4.79 //x2=10.02 //y2=4.865
r416 (  145 147 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=10.02 //y=4.7 //x2=10.02 //y2=4.79
r417 (  141 142 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=9.99 //y=2.08 //x2=9.99 //y2=1.915
r418 (  131 165 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.545 //y=1.25 //x2=20.505 //y2=1.405
r419 (  130 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.545 //y=0.905 //x2=20.505 //y2=0.75
r420 (  130 131 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.545 //y=0.905 //x2=20.545 //y2=1.25
r421 (  125 163 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.17 //y=1.405 //x2=20.055 //y2=1.405
r422 (  124 165 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.39 //y=1.405 //x2=20.505 //y2=1.405
r423 (  123 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.17 //y=0.75 //x2=20.055 //y2=0.75
r424 (  122 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.39 //y=0.75 //x2=20.505 //y2=0.75
r425 (  122 123 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=20.39 //y=0.75 //x2=20.17 //y2=0.75
r426 (  121 160 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=20.145 //y=4.79 //x2=20.01 //y2=4.79
r427 (  120 127 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.385 //y=4.79 //x2=20.46 //y2=4.865
r428 (  120 121 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=20.385 //y=4.79 //x2=20.145 //y2=4.79
r429 (  115 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.015 //y=1.56 //x2=20.055 //y2=1.405
r430 (  115 155 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=20.015 //y=1.56 //x2=20.015 //y2=1.915
r431 (  114 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.015 //y=1.25 //x2=20.055 //y2=1.405
r432 (  113 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.015 //y=0.905 //x2=20.055 //y2=0.75
r433 (  113 114 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.015 //y=0.905 //x2=20.015 //y2=1.25
r434 (  112 152 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.555 //y=1.25 //x2=10.515 //y2=1.405
r435 (  111 151 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.555 //y=0.905 //x2=10.515 //y2=0.75
r436 (  111 112 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.555 //y=0.905 //x2=10.555 //y2=1.25
r437 (  106 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.18 //y=1.405 //x2=10.065 //y2=1.405
r438 (  105 152 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.4 //y=1.405 //x2=10.515 //y2=1.405
r439 (  104 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.18 //y=0.75 //x2=10.065 //y2=0.75
r440 (  103 151 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.4 //y=0.75 //x2=10.515 //y2=0.75
r441 (  103 104 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.4 //y=0.75 //x2=10.18 //y2=0.75
r442 (  102 147 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=10.155 //y=4.79 //x2=10.02 //y2=4.79
r443 (  101 108 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.395 //y=4.79 //x2=10.47 //y2=4.865
r444 (  101 102 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=10.395 //y=4.79 //x2=10.155 //y2=4.79
r445 (  96 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.025 //y=1.56 //x2=10.065 //y2=1.405
r446 (  96 142 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=10.025 //y=1.56 //x2=10.025 //y2=1.915
r447 (  95 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.025 //y=1.25 //x2=10.065 //y2=1.405
r448 (  94 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.025 //y=0.905 //x2=10.065 //y2=0.75
r449 (  94 95 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.025 //y=0.905 //x2=10.025 //y2=1.25
r450 (  89 91 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.75 //y2=4.865
r451 (  89 90 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.385 //y2=4.79
r452 (  88 139 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=1.22 //x2=1.3 //y2=1.375
r453 (  87 138 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.3 //y2=0.72
r454 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.34 //y2=1.22
r455 (  84 90 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.385 //y2=4.79
r456 (  84 137 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.11 //y2=4.7
r457 (  82 133 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=1.375 //x2=0.85 //y2=1.375
r458 (  81 139 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=1.375 //x2=1.3 //y2=1.375
r459 (  80 132 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=0.72 //x2=0.85 //y2=0.72
r460 (  79 138 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=1.3 //y2=0.72
r461 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=0.965 //y2=0.72
r462 (  78 135 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.915 //x2=1.11 //y2=2.08
r463 (  77 133 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.85 //y2=1.375
r464 (  77 78 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.81 //y2=1.915
r465 (  76 133 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.22 //x2=0.85 //y2=1.375
r466 (  75 132 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.85 //y2=0.72
r467 (  75 76 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.81 //y2=1.22
r468 (  74 127 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.46 //y=6.02 //x2=20.46 //y2=4.865
r469 (  73 161 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.02 //y=6.02 //x2=20.02 //y2=4.865
r470 (  72 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.47 //y=6.02 //x2=10.47 //y2=4.865
r471 (  71 148 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.03 //y=6.02 //x2=10.03 //y2=4.865
r472 (  70 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.75 //y=6.02 //x2=1.75 //y2=4.865
r473 (  69 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.31 //y=6.02 //x2=1.31 //y2=4.865
r474 (  68 124 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.28 //y=1.405 //x2=20.39 //y2=1.405
r475 (  68 125 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.28 //y=1.405 //x2=20.17 //y2=1.405
r476 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.29 //y=1.405 //x2=10.4 //y2=1.405
r477 (  67 106 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.29 //y=1.405 //x2=10.18 //y2=1.405
r478 (  66 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=1.185 //y2=1.375
r479 (  66 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=0.965 //y2=1.375
r480 (  65 158 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.01 //y=4.7 //x2=20.01 //y2=4.7
r481 (  62 145 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.02 //y=4.7 //x2=10.02 //y2=4.7
r482 (  57 154 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.98 //y=2.08 //x2=19.98 //y2=2.08
r483 (  57 60 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.08 //x2=19.98 //y2=4.07
r484 (  55 65 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=19.98 //y=4.535 //x2=19.995 //y2=4.7
r485 (  55 60 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=19.98 //y=4.535 //x2=19.98 //y2=4.07
r486 (  52 54 ) resistor r=71.5294 //w=0.187 //l=1.045 //layer=li \
 //thickness=0.1 //x=14.06 //y=5.115 //x2=14.06 //y2=4.07
r487 (  51 54 ) resistor r=159.487 //w=0.187 //l=2.33 //layer=li \
 //thickness=0.1 //x=14.06 //y=1.74 //x2=14.06 //y2=4.07
r488 (  49 51 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.975 //y=1.655 //x2=14.06 //y2=1.74
r489 (  49 50 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=13.975 //y=1.655 //x2=13.705 //y2=1.655
r490 (  48 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.665 //y=5.2 //x2=13.58 //y2=5.2
r491 (  47 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.975 //y=5.2 //x2=14.06 //y2=5.115
r492 (  47 48 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=13.975 //y=5.2 //x2=13.665 //y2=5.2
r493 (  43 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.62 //y=1.57 //x2=13.705 //y2=1.655
r494 (  43 166 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=13.62 //y=1.57 //x2=13.62 //y2=1
r495 (  37 63 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.58 //y=5.285 //x2=13.58 //y2=5.2
r496 (  37 169 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=13.58 //y=5.285 //x2=13.58 //y2=5.725
r497 (  35 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.495 //y=5.2 //x2=13.58 //y2=5.2
r498 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=13.495 //y=5.2 //x2=12.785 //y2=5.2
r499 (  29 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.7 //y=5.285 //x2=12.785 //y2=5.2
r500 (  29 168 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=12.7 //y=5.285 //x2=12.7 //y2=5.725
r501 (  25 141 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.99 //y=2.08 //x2=9.99 //y2=2.08
r502 (  25 28 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=9.99 //y=2.08 //x2=9.99 //y2=4.07
r503 (  23 62 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=9.99 //y=4.535 //x2=10.005 //y2=4.7
r504 (  23 28 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=9.99 //y=4.535 //x2=9.99 //y2=4.07
r505 (  21 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r506 (  19 21 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.07 //x2=1.11 //y2=4.7
r507 (  16 135 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r508 (  16 19 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.08 //x2=1.11 //y2=4.07
r509 (  14 60 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=19.98 //y=4.07 //x2=19.98 //y2=4.07
r510 (  12 54 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.06 //y=4.07 //x2=14.06 //y2=4.07
r511 (  10 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.99 //y=4.07 //x2=9.99 //y2=4.07
r512 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.07
r513 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=14.175 //y=4.07 //x2=14.06 //y2=4.07
r514 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=19.865 //y=4.07 //x2=19.98 //y2=4.07
r515 (  5 6 ) resistor r=5.42939 //w=0.131 //l=5.69 //layer=m1 \
 //thickness=0.36 //x=19.865 //y=4.07 //x2=14.175 //y2=4.07
r516 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.105 //y=4.07 //x2=9.99 //y2=4.07
r517 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=4.07 //x2=14.06 //y2=4.07
r518 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=4.07 //x2=10.105 //y2=4.07
r519 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.225 //y=4.07 //x2=1.11 //y2=4.07
r520 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.875 //y=4.07 //x2=9.99 //y2=4.07
r521 (  1 2 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=9.875 //y=4.07 //x2=1.225 //y2=4.07
ends PM_TMRDFFQNX1\%noxref_7

subckt PM_TMRDFFQNX1\%noxref_8 ( 1 2 3 4 12 25 26 37 39 40 44 46 53 54 55 56 \
 57 58 59 63 64 65 70 72 75 76 77 78 79 80 84 86 89 90 95 96 101 110 113 115 \
 116 )
c232 ( 116 0 ) capacitor c=0.0220291f //x=28.235 //y=5.02
c233 ( 115 0 ) capacitor c=0.0217503f //x=27.355 //y=5.02
c234 ( 113 0 ) capacitor c=0.00866655f //x=28.23 //y=0.905
c235 ( 110 0 ) capacitor c=0.0588816f //x=30.71 //y=4.7
c236 ( 101 0 ) capacitor c=0.058931f //x=24.79 //y=4.7
c237 ( 96 0 ) capacitor c=0.0273931f //x=24.79 //y=1.915
c238 ( 95 0 ) capacitor c=0.0457054f //x=24.79 //y=2.08
c239 ( 90 0 ) capacitor c=0.0318948f //x=31.045 //y=1.21
c240 ( 89 0 ) capacitor c=0.0187384f //x=31.045 //y=0.865
c241 ( 86 0 ) capacitor c=0.0141798f //x=30.89 //y=1.365
c242 ( 84 0 ) capacitor c=0.0149844f //x=30.89 //y=0.71
c243 ( 80 0 ) capacitor c=0.0816311f //x=30.515 //y=1.915
c244 ( 79 0 ) capacitor c=0.0229722f //x=30.515 //y=1.52
c245 ( 78 0 ) capacitor c=0.0234352f //x=30.515 //y=1.21
c246 ( 77 0 ) capacitor c=0.0199343f //x=30.515 //y=0.865
c247 ( 76 0 ) capacitor c=0.0432517f //x=25.31 //y=1.26
c248 ( 75 0 ) capacitor c=0.0200379f //x=25.31 //y=0.915
c249 ( 72 0 ) capacitor c=0.0158629f //x=25.155 //y=1.415
c250 ( 70 0 ) capacitor c=0.0157803f //x=25.155 //y=0.76
c251 ( 65 0 ) capacitor c=0.0218028f //x=24.78 //y=1.57
c252 ( 64 0 ) capacitor c=0.0207459f //x=24.78 //y=1.26
c253 ( 63 0 ) capacitor c=0.0194308f //x=24.78 //y=0.915
c254 ( 59 0 ) capacitor c=0.110275f //x=31.05 //y=6.02
c255 ( 58 0 ) capacitor c=0.154305f //x=30.61 //y=6.02
c256 ( 57 0 ) capacitor c=0.158794f //x=24.97 //y=6.02
c257 ( 56 0 ) capacitor c=0.110114f //x=24.53 //y=6.02
c258 ( 53 0 ) capacitor c=0.00211606f //x=28.38 //y=5.2
c259 ( 46 0 ) capacitor c=0.0864117f //x=30.71 //y=2.08
c260 ( 44 0 ) capacitor c=0.103161f //x=28.86 //y=3.33
c261 ( 40 0 ) capacitor c=0.00436419f //x=28.505 //y=1.655
c262 ( 39 0 ) capacitor c=0.0127039f //x=28.775 //y=1.655
c263 ( 37 0 ) capacitor c=0.0137522f //x=28.775 //y=5.2
c264 ( 26 0 ) capacitor c=0.00251635f //x=27.585 //y=5.2
c265 ( 25 0 ) capacitor c=0.0142423f //x=28.295 //y=5.2
c266 ( 12 0 ) capacitor c=0.0836809f //x=24.79 //y=2.08
c267 ( 4 0 ) capacitor c=0.00280195f //x=28.975 //y=3.33
c268 ( 3 0 ) capacitor c=0.0346903f //x=30.595 //y=3.33
c269 ( 2 0 ) capacitor c=0.0127233f //x=24.905 //y=3.33
c270 ( 1 0 ) capacitor c=0.0559579f //x=28.745 //y=3.33
r271 (  108 110 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=30.61 //y=4.7 //x2=30.71 //y2=4.7
r272 (  95 96 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=24.79 //y=2.08 //x2=24.79 //y2=1.915
r273 (  91 110 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=31.05 //y=4.865 //x2=30.71 //y2=4.7
r274 (  90 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.045 //y=1.21 //x2=31.005 //y2=1.365
r275 (  89 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.045 //y=0.865 //x2=31.005 //y2=0.71
r276 (  89 90 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=31.045 //y=0.865 //x2=31.045 //y2=1.21
r277 (  87 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.67 //y=1.365 //x2=30.555 //y2=1.365
r278 (  86 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.89 //y=1.365 //x2=31.005 //y2=1.365
r279 (  85 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.67 //y=0.71 //x2=30.555 //y2=0.71
r280 (  84 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.89 //y=0.71 //x2=31.005 //y2=0.71
r281 (  84 85 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=30.89 //y=0.71 //x2=30.67 //y2=0.71
r282 (  81 108 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=30.61 //y=4.865 //x2=30.61 //y2=4.7
r283 (  80 105 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=30.515 //y=1.915 //x2=30.71 //y2=2.08
r284 (  79 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.515 //y=1.52 //x2=30.555 //y2=1.365
r285 (  79 80 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=30.515 //y=1.52 //x2=30.515 //y2=1.915
r286 (  78 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.515 //y=1.21 //x2=30.555 //y2=1.365
r287 (  77 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.515 //y=0.865 //x2=30.555 //y2=0.71
r288 (  77 78 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=30.515 //y=0.865 //x2=30.515 //y2=1.21
r289 (  76 103 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.31 //y=1.26 //x2=25.27 //y2=1.415
r290 (  75 102 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.31 //y=0.915 //x2=25.27 //y2=0.76
r291 (  75 76 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=25.31 //y=0.915 //x2=25.31 //y2=1.26
r292 (  73 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.935 //y=1.415 //x2=24.82 //y2=1.415
r293 (  72 103 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.155 //y=1.415 //x2=25.27 //y2=1.415
r294 (  71 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.935 //y=0.76 //x2=24.82 //y2=0.76
r295 (  70 102 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.155 //y=0.76 //x2=25.27 //y2=0.76
r296 (  70 71 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=25.155 //y=0.76 //x2=24.935 //y2=0.76
r297 (  67 101 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=24.97 //y=4.865 //x2=24.79 //y2=4.7
r298 (  65 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.78 //y=1.57 //x2=24.82 //y2=1.415
r299 (  65 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.78 //y=1.57 //x2=24.78 //y2=1.915
r300 (  64 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.78 //y=1.26 //x2=24.82 //y2=1.415
r301 (  63 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.78 //y=0.915 //x2=24.82 //y2=0.76
r302 (  63 64 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.78 //y=0.915 //x2=24.78 //y2=1.26
r303 (  60 101 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=24.53 //y=4.865 //x2=24.79 //y2=4.7
r304 (  59 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=31.05 //y=6.02 //x2=31.05 //y2=4.865
r305 (  58 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=30.61 //y=6.02 //x2=30.61 //y2=4.865
r306 (  57 67 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=24.97 //y=6.02 //x2=24.97 //y2=4.865
r307 (  56 60 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=24.53 //y=6.02 //x2=24.53 //y2=4.865
r308 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=30.78 //y=1.365 //x2=30.89 //y2=1.365
r309 (  55 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=30.78 //y=1.365 //x2=30.67 //y2=1.365
r310 (  54 72 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.045 //y=1.415 //x2=25.155 //y2=1.415
r311 (  54 73 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.045 //y=1.415 //x2=24.935 //y2=1.415
r312 (  51 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=30.71 //y=4.7 //x2=30.71 //y2=4.7
r313 (  49 51 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=30.71 //y=3.33 //x2=30.71 //y2=4.7
r314 (  46 105 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=30.71 //y=2.08 //x2=30.71 //y2=2.08
r315 (  46 49 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=30.71 //y=2.08 //x2=30.71 //y2=3.33
r316 (  42 44 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=28.86 //y=5.115 //x2=28.86 //y2=3.33
r317 (  41 44 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=28.86 //y=1.74 //x2=28.86 //y2=3.33
r318 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=28.775 //y=1.655 //x2=28.86 //y2=1.74
r319 (  39 40 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=28.775 //y=1.655 //x2=28.505 //y2=1.655
r320 (  38 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.465 //y=5.2 //x2=28.38 //y2=5.2
r321 (  37 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=28.775 //y=5.2 //x2=28.86 //y2=5.115
r322 (  37 38 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=28.775 //y=5.2 //x2=28.465 //y2=5.2
r323 (  33 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=28.42 //y=1.57 //x2=28.505 //y2=1.655
r324 (  33 113 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=28.42 //y=1.57 //x2=28.42 //y2=1
r325 (  27 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.38 //y=5.285 //x2=28.38 //y2=5.2
r326 (  27 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=28.38 //y=5.285 //x2=28.38 //y2=5.725
r327 (  25 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.295 //y=5.2 //x2=28.38 //y2=5.2
r328 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=28.295 //y=5.2 //x2=27.585 //y2=5.2
r329 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=27.5 //y=5.285 //x2=27.585 //y2=5.2
r330 (  19 115 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=27.5 //y=5.285 //x2=27.5 //y2=5.725
r331 (  17 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=24.79 //y=4.7 //x2=24.79 //y2=4.7
r332 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=24.79 //y=3.33 //x2=24.79 //y2=4.7
r333 (  12 95 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=24.79 //y=2.08 //x2=24.79 //y2=2.08
r334 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=24.79 //y=2.08 //x2=24.79 //y2=3.33
r335 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=30.71 //y=3.33 //x2=30.71 //y2=3.33
r336 (  8 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=28.86 //y=3.33 //x2=28.86 //y2=3.33
r337 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=24.79 //y=3.33 //x2=24.79 //y2=3.33
r338 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=28.975 //y=3.33 //x2=28.86 //y2=3.33
r339 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=30.595 //y=3.33 //x2=30.71 //y2=3.33
r340 (  3 4 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=30.595 //y=3.33 //x2=28.975 //y2=3.33
r341 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=24.905 //y=3.33 //x2=24.79 //y2=3.33
r342 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=28.745 //y=3.33 //x2=28.86 //y2=3.33
r343 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=28.745 //y=3.33 //x2=24.905 //y2=3.33
ends PM_TMRDFFQNX1\%noxref_8

subckt PM_TMRDFFQNX1\%noxref_9 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 \
 48 52 54 57 58 68 71 73 74 )
c153 ( 74 0 ) capacitor c=0.0220291f //x=31.565 //y=5.02
c154 ( 73 0 ) capacitor c=0.0217503f //x=30.685 //y=5.02
c155 ( 71 0 ) capacitor c=0.00866655f //x=31.56 //y=0.905
c156 ( 68 0 ) capacitor c=0.0588816f //x=34.04 //y=4.7
c157 ( 58 0 ) capacitor c=0.0318948f //x=34.375 //y=1.21
c158 ( 57 0 ) capacitor c=0.0187384f //x=34.375 //y=0.865
c159 ( 54 0 ) capacitor c=0.0141798f //x=34.22 //y=1.365
c160 ( 52 0 ) capacitor c=0.0149844f //x=34.22 //y=0.71
c161 ( 48 0 ) capacitor c=0.0816311f //x=33.845 //y=1.915
c162 ( 47 0 ) capacitor c=0.0229722f //x=33.845 //y=1.52
c163 ( 46 0 ) capacitor c=0.0234352f //x=33.845 //y=1.21
c164 ( 45 0 ) capacitor c=0.0199343f //x=33.845 //y=0.865
c165 ( 44 0 ) capacitor c=0.110275f //x=34.38 //y=6.02
c166 ( 43 0 ) capacitor c=0.154305f //x=33.94 //y=6.02
c167 ( 41 0 ) capacitor c=0.00211606f //x=31.71 //y=5.2
c168 ( 34 0 ) capacitor c=0.0859106f //x=34.04 //y=2.08
c169 ( 32 0 ) capacitor c=0.103708f //x=32.19 //y=3.33
c170 ( 28 0 ) capacitor c=0.00436419f //x=31.835 //y=1.655
c171 ( 27 0 ) capacitor c=0.0127039f //x=32.105 //y=1.655
c172 ( 25 0 ) capacitor c=0.0137522f //x=32.105 //y=5.2
c173 ( 14 0 ) capacitor c=0.00251459f //x=30.915 //y=5.2
c174 ( 13 0 ) capacitor c=0.0143649f //x=31.625 //y=5.2
c175 ( 2 0 ) capacitor c=0.00668619f //x=32.305 //y=3.33
c176 ( 1 0 ) capacitor c=0.0400514f //x=33.925 //y=3.33
r177 (  66 68 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=33.94 //y=4.7 //x2=34.04 //y2=4.7
r178 (  59 68 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=34.38 //y=4.865 //x2=34.04 //y2=4.7
r179 (  58 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.375 //y=1.21 //x2=34.335 //y2=1.365
r180 (  57 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.375 //y=0.865 //x2=34.335 //y2=0.71
r181 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=34.375 //y=0.865 //x2=34.375 //y2=1.21
r182 (  55 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34 //y=1.365 //x2=33.885 //y2=1.365
r183 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.22 //y=1.365 //x2=34.335 //y2=1.365
r184 (  53 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34 //y=0.71 //x2=33.885 //y2=0.71
r185 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.22 //y=0.71 //x2=34.335 //y2=0.71
r186 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=34.22 //y=0.71 //x2=34 //y2=0.71
r187 (  49 66 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=33.94 //y=4.865 //x2=33.94 //y2=4.7
r188 (  48 63 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=33.845 //y=1.915 //x2=34.04 //y2=2.08
r189 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.845 //y=1.52 //x2=33.885 //y2=1.365
r190 (  47 48 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=33.845 //y=1.52 //x2=33.845 //y2=1.915
r191 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.845 //y=1.21 //x2=33.885 //y2=1.365
r192 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.845 //y=0.865 //x2=33.885 //y2=0.71
r193 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=33.845 //y=0.865 //x2=33.845 //y2=1.21
r194 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=34.38 //y=6.02 //x2=34.38 //y2=4.865
r195 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=33.94 //y=6.02 //x2=33.94 //y2=4.865
r196 (  42 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=34.11 //y=1.365 //x2=34.22 //y2=1.365
r197 (  42 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=34.11 //y=1.365 //x2=34 //y2=1.365
r198 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.04 //y=4.7 //x2=34.04 //y2=4.7
r199 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=34.04 //y=3.33 //x2=34.04 //y2=4.7
r200 (  34 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.04 //y=2.08 //x2=34.04 //y2=2.08
r201 (  34 37 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=34.04 //y=2.08 //x2=34.04 //y2=3.33
r202 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=32.19 //y=5.115 //x2=32.19 //y2=3.33
r203 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=32.19 //y=1.74 //x2=32.19 //y2=3.33
r204 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.105 //y=1.655 //x2=32.19 //y2=1.74
r205 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=32.105 //y=1.655 //x2=31.835 //y2=1.655
r206 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.795 //y=5.2 //x2=31.71 //y2=5.2
r207 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.105 //y=5.2 //x2=32.19 //y2=5.115
r208 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=32.105 //y=5.2 //x2=31.795 //y2=5.2
r209 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=31.75 //y=1.57 //x2=31.835 //y2=1.655
r210 (  21 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=31.75 //y=1.57 //x2=31.75 //y2=1
r211 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.71 //y=5.285 //x2=31.71 //y2=5.2
r212 (  15 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=31.71 //y=5.285 //x2=31.71 //y2=5.725
r213 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.625 //y=5.2 //x2=31.71 //y2=5.2
r214 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=31.625 //y=5.2 //x2=30.915 //y2=5.2
r215 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=30.83 //y=5.285 //x2=30.915 //y2=5.2
r216 (  7 73 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=30.83 //y=5.285 //x2=30.83 //y2=5.725
r217 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=34.04 //y=3.33 //x2=34.04 //y2=3.33
r218 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=32.19 //y=3.33 //x2=32.19 //y2=3.33
r219 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=32.305 //y=3.33 //x2=32.19 //y2=3.33
r220 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=33.925 //y=3.33 //x2=34.04 //y2=3.33
r221 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=33.925 //y=3.33 //x2=32.305 //y2=3.33
ends PM_TMRDFFQNX1\%noxref_9

subckt PM_TMRDFFQNX1\%noxref_10 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 63 \
 64 65 66 67 68 69 70 71 72 76 78 81 82 86 87 88 89 93 95 98 99 109 118 121 \
 123 124 125 )
c258 ( 125 0 ) capacitor c=0.023087f //x=24.605 //y=5.02
c259 ( 124 0 ) capacitor c=0.023519f //x=23.725 //y=5.02
c260 ( 123 0 ) capacitor c=0.0224735f //x=22.845 //y=5.02
c261 ( 121 0 ) capacitor c=0.00872971f //x=24.855 //y=0.915
c262 ( 118 0 ) capacitor c=0.0588816f //x=37.37 //y=4.7
c263 ( 109 0 ) capacitor c=0.0588816f //x=27.38 //y=4.7
c264 ( 99 0 ) capacitor c=0.0318948f //x=37.705 //y=1.21
c265 ( 98 0 ) capacitor c=0.0187384f //x=37.705 //y=0.865
c266 ( 95 0 ) capacitor c=0.0141798f //x=37.55 //y=1.365
c267 ( 93 0 ) capacitor c=0.0149844f //x=37.55 //y=0.71
c268 ( 89 0 ) capacitor c=0.0816311f //x=37.175 //y=1.915
c269 ( 88 0 ) capacitor c=0.0229722f //x=37.175 //y=1.52
c270 ( 87 0 ) capacitor c=0.0234352f //x=37.175 //y=1.21
c271 ( 86 0 ) capacitor c=0.0199343f //x=37.175 //y=0.865
c272 ( 82 0 ) capacitor c=0.0318948f //x=27.715 //y=1.21
c273 ( 81 0 ) capacitor c=0.0187384f //x=27.715 //y=0.865
c274 ( 78 0 ) capacitor c=0.0141798f //x=27.56 //y=1.365
c275 ( 76 0 ) capacitor c=0.0149844f //x=27.56 //y=0.71
c276 ( 72 0 ) capacitor c=0.0816311f //x=27.185 //y=1.915
c277 ( 71 0 ) capacitor c=0.0229722f //x=27.185 //y=1.52
c278 ( 70 0 ) capacitor c=0.0234352f //x=27.185 //y=1.21
c279 ( 69 0 ) capacitor c=0.0199343f //x=27.185 //y=0.865
c280 ( 68 0 ) capacitor c=0.110275f //x=37.71 //y=6.02
c281 ( 67 0 ) capacitor c=0.154305f //x=37.27 //y=6.02
c282 ( 66 0 ) capacitor c=0.110275f //x=27.72 //y=6.02
c283 ( 65 0 ) capacitor c=0.154305f //x=27.28 //y=6.02
c284 ( 62 0 ) capacitor c=0.00106608f //x=24.75 //y=5.155
c285 ( 61 0 ) capacitor c=0.00207162f //x=23.87 //y=5.155
c286 ( 54 0 ) capacitor c=0.0890863f //x=37.37 //y=2.08
c287 ( 46 0 ) capacitor c=0.0858897f //x=27.38 //y=2.08
c288 ( 44 0 ) capacitor c=0.104635f //x=25.53 //y=3.7
c289 ( 40 0 ) capacitor c=0.00431225f //x=25.13 //y=1.665
c290 ( 39 0 ) capacitor c=0.0143009f //x=25.445 //y=1.665
c291 ( 33 0 ) capacitor c=0.0284988f //x=25.445 //y=5.155
c292 ( 25 0 ) capacitor c=0.0176454f //x=24.665 //y=5.155
c293 ( 18 0 ) capacitor c=0.00332903f //x=23.075 //y=5.155
c294 ( 17 0 ) capacitor c=0.014837f //x=23.785 //y=5.155
c295 ( 4 0 ) capacitor c=0.00424317f //x=27.495 //y=3.7
c296 ( 3 0 ) capacitor c=0.161586f //x=37.255 //y=3.7
c297 ( 2 0 ) capacitor c=0.0125346f //x=25.645 //y=3.7
c298 ( 1 0 ) capacitor c=0.0285004f //x=27.265 //y=3.7
r299 (  116 118 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=37.27 //y=4.7 //x2=37.37 //y2=4.7
r300 (  107 109 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=27.28 //y=4.7 //x2=27.38 //y2=4.7
r301 (  100 118 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=37.71 //y=4.865 //x2=37.37 //y2=4.7
r302 (  99 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.705 //y=1.21 //x2=37.665 //y2=1.365
r303 (  98 119 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.705 //y=0.865 //x2=37.665 //y2=0.71
r304 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=37.705 //y=0.865 //x2=37.705 //y2=1.21
r305 (  96 115 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.33 //y=1.365 //x2=37.215 //y2=1.365
r306 (  95 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.55 //y=1.365 //x2=37.665 //y2=1.365
r307 (  94 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.33 //y=0.71 //x2=37.215 //y2=0.71
r308 (  93 119 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.55 //y=0.71 //x2=37.665 //y2=0.71
r309 (  93 94 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=37.55 //y=0.71 //x2=37.33 //y2=0.71
r310 (  90 116 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=37.27 //y=4.865 //x2=37.27 //y2=4.7
r311 (  89 113 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=37.175 //y=1.915 //x2=37.37 //y2=2.08
r312 (  88 115 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.175 //y=1.52 //x2=37.215 //y2=1.365
r313 (  88 89 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=37.175 //y=1.52 //x2=37.175 //y2=1.915
r314 (  87 115 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.175 //y=1.21 //x2=37.215 //y2=1.365
r315 (  86 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.175 //y=0.865 //x2=37.215 //y2=0.71
r316 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=37.175 //y=0.865 //x2=37.175 //y2=1.21
r317 (  83 109 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=27.72 //y=4.865 //x2=27.38 //y2=4.7
r318 (  82 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.715 //y=1.21 //x2=27.675 //y2=1.365
r319 (  81 110 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.715 //y=0.865 //x2=27.675 //y2=0.71
r320 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.715 //y=0.865 //x2=27.715 //y2=1.21
r321 (  79 106 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.34 //y=1.365 //x2=27.225 //y2=1.365
r322 (  78 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.56 //y=1.365 //x2=27.675 //y2=1.365
r323 (  77 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.34 //y=0.71 //x2=27.225 //y2=0.71
r324 (  76 110 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.56 //y=0.71 //x2=27.675 //y2=0.71
r325 (  76 77 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=27.56 //y=0.71 //x2=27.34 //y2=0.71
r326 (  73 107 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=27.28 //y=4.865 //x2=27.28 //y2=4.7
r327 (  72 104 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=27.185 //y=1.915 //x2=27.38 //y2=2.08
r328 (  71 106 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.185 //y=1.52 //x2=27.225 //y2=1.365
r329 (  71 72 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=27.185 //y=1.52 //x2=27.185 //y2=1.915
r330 (  70 106 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.185 //y=1.21 //x2=27.225 //y2=1.365
r331 (  69 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.185 //y=0.865 //x2=27.225 //y2=0.71
r332 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.185 //y=0.865 //x2=27.185 //y2=1.21
r333 (  68 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=37.71 //y=6.02 //x2=37.71 //y2=4.865
r334 (  67 90 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=37.27 //y=6.02 //x2=37.27 //y2=4.865
r335 (  66 83 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=27.72 //y=6.02 //x2=27.72 //y2=4.865
r336 (  65 73 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=27.28 //y=6.02 //x2=27.28 //y2=4.865
r337 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=37.44 //y=1.365 //x2=37.55 //y2=1.365
r338 (  64 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=37.44 //y=1.365 //x2=37.33 //y2=1.365
r339 (  63 78 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=27.45 //y=1.365 //x2=27.56 //y2=1.365
r340 (  63 79 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=27.45 //y=1.365 //x2=27.34 //y2=1.365
r341 (  59 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=37.37 //y=4.7 //x2=37.37 //y2=4.7
r342 (  57 59 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=37.37 //y=3.7 //x2=37.37 //y2=4.7
r343 (  54 113 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=37.37 //y=2.08 //x2=37.37 //y2=2.08
r344 (  54 57 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=37.37 //y=2.08 //x2=37.37 //y2=3.7
r345 (  51 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=27.38 //y=4.7 //x2=27.38 //y2=4.7
r346 (  49 51 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=27.38 //y=3.7 //x2=27.38 //y2=4.7
r347 (  46 104 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=27.38 //y=2.08 //x2=27.38 //y2=2.08
r348 (  46 49 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=27.38 //y=2.08 //x2=27.38 //y2=3.7
r349 (  42 44 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=25.53 //y=5.07 //x2=25.53 //y2=3.7
r350 (  41 44 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=25.53 //y=1.75 //x2=25.53 //y2=3.7
r351 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.445 //y=1.665 //x2=25.53 //y2=1.75
r352 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=25.445 //y=1.665 //x2=25.13 //y2=1.665
r353 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.045 //y=1.58 //x2=25.13 //y2=1.665
r354 (  35 121 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=25.045 //y=1.58 //x2=25.045 //y2=1.01
r355 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.835 //y=5.155 //x2=24.75 //y2=5.155
r356 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.445 //y=5.155 //x2=25.53 //y2=5.07
r357 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=25.445 //y=5.155 //x2=24.835 //y2=5.155
r358 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.75 //y=5.24 //x2=24.75 //y2=5.155
r359 (  27 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=24.75 //y=5.24 //x2=24.75 //y2=5.725
r360 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.955 //y=5.155 //x2=23.87 //y2=5.155
r361 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.665 //y=5.155 //x2=24.75 //y2=5.155
r362 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=24.665 //y=5.155 //x2=23.955 //y2=5.155
r363 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.87 //y=5.24 //x2=23.87 //y2=5.155
r364 (  19 124 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=23.87 //y=5.24 //x2=23.87 //y2=5.725
r365 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.785 //y=5.155 //x2=23.87 //y2=5.155
r366 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=23.785 //y=5.155 //x2=23.075 //y2=5.155
r367 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=22.99 //y=5.24 //x2=23.075 //y2=5.155
r368 (  11 123 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.99 //y=5.24 //x2=22.99 //y2=5.725
r369 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=37.37 //y=3.7 //x2=37.37 //y2=3.7
r370 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=27.38 //y=3.7 //x2=27.38 //y2=3.7
r371 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=25.53 //y=3.7 //x2=25.53 //y2=3.7
r372 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=27.495 //y=3.7 //x2=27.38 //y2=3.7
r373 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=37.255 //y=3.7 //x2=37.37 //y2=3.7
r374 (  3 4 ) resistor r=9.31298 //w=0.131 //l=9.76 //layer=m1 \
 //thickness=0.36 //x=37.255 //y=3.7 //x2=27.495 //y2=3.7
r375 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=25.645 //y=3.7 //x2=25.53 //y2=3.7
r376 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=27.265 //y=3.7 //x2=27.38 //y2=3.7
r377 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=27.265 //y=3.7 //x2=25.645 //y2=3.7
ends PM_TMRDFFQNX1\%noxref_10

subckt PM_TMRDFFQNX1\%noxref_11 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 \
 47 48 52 54 57 58 68 71 73 74 )
c151 ( 74 0 ) capacitor c=0.0220291f //x=38.225 //y=5.02
c152 ( 73 0 ) capacitor c=0.0217503f //x=37.345 //y=5.02
c153 ( 71 0 ) capacitor c=0.00866655f //x=38.22 //y=0.905
c154 ( 68 0 ) capacitor c=0.0588816f //x=40.7 //y=4.7
c155 ( 58 0 ) capacitor c=0.0318948f //x=41.035 //y=1.21
c156 ( 57 0 ) capacitor c=0.0187384f //x=41.035 //y=0.865
c157 ( 54 0 ) capacitor c=0.0141798f //x=40.88 //y=1.365
c158 ( 52 0 ) capacitor c=0.0149844f //x=40.88 //y=0.71
c159 ( 48 0 ) capacitor c=0.0813322f //x=40.505 //y=1.915
c160 ( 47 0 ) capacitor c=0.0229267f //x=40.505 //y=1.52
c161 ( 46 0 ) capacitor c=0.0234352f //x=40.505 //y=1.21
c162 ( 45 0 ) capacitor c=0.0199343f //x=40.505 //y=0.865
c163 ( 44 0 ) capacitor c=0.110275f //x=41.04 //y=6.02
c164 ( 43 0 ) capacitor c=0.154305f //x=40.6 //y=6.02
c165 ( 41 0 ) capacitor c=0.00211606f //x=38.37 //y=5.2
c166 ( 34 0 ) capacitor c=0.0867306f //x=40.7 //y=2.08
c167 ( 32 0 ) capacitor c=0.105846f //x=38.85 //y=3.7
c168 ( 28 0 ) capacitor c=0.00404073f //x=38.495 //y=1.655
c169 ( 27 0 ) capacitor c=0.0122201f //x=38.765 //y=1.655
c170 ( 25 0 ) capacitor c=0.0137522f //x=38.765 //y=5.2
c171 ( 14 0 ) capacitor c=0.00251459f //x=37.575 //y=5.2
c172 ( 13 0 ) capacitor c=0.0142423f //x=38.285 //y=5.2
c173 ( 2 0 ) capacitor c=0.00701934f //x=38.965 //y=3.7
c174 ( 1 0 ) capacitor c=0.0472012f //x=40.585 //y=3.7
r175 (  66 68 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=40.6 //y=4.7 //x2=40.7 //y2=4.7
r176 (  59 68 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=41.04 //y=4.865 //x2=40.7 //y2=4.7
r177 (  58 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.035 //y=1.21 //x2=40.995 //y2=1.365
r178 (  57 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.035 //y=0.865 //x2=40.995 //y2=0.71
r179 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=41.035 //y=0.865 //x2=41.035 //y2=1.21
r180 (  55 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.66 //y=1.365 //x2=40.545 //y2=1.365
r181 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.88 //y=1.365 //x2=40.995 //y2=1.365
r182 (  53 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.66 //y=0.71 //x2=40.545 //y2=0.71
r183 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.88 //y=0.71 //x2=40.995 //y2=0.71
r184 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=40.88 //y=0.71 //x2=40.66 //y2=0.71
r185 (  49 66 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=40.6 //y=4.865 //x2=40.6 //y2=4.7
r186 (  48 63 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=40.505 //y=1.915 //x2=40.7 //y2=2.08
r187 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.505 //y=1.52 //x2=40.545 //y2=1.365
r188 (  47 48 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=40.505 //y=1.52 //x2=40.505 //y2=1.915
r189 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.505 //y=1.21 //x2=40.545 //y2=1.365
r190 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.505 //y=0.865 //x2=40.545 //y2=0.71
r191 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=40.505 //y=0.865 //x2=40.505 //y2=1.21
r192 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.04 //y=6.02 //x2=41.04 //y2=4.865
r193 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=40.6 //y=6.02 //x2=40.6 //y2=4.865
r194 (  42 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=40.77 //y=1.365 //x2=40.88 //y2=1.365
r195 (  42 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=40.77 //y=1.365 //x2=40.66 //y2=1.365
r196 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=40.7 //y=4.7 //x2=40.7 //y2=4.7
r197 (  37 39 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=40.7 //y=3.7 //x2=40.7 //y2=4.7
r198 (  34 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=40.7 //y=2.08 //x2=40.7 //y2=2.08
r199 (  34 37 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=40.7 //y=2.08 //x2=40.7 //y2=3.7
r200 (  30 32 ) resistor r=96.8556 //w=0.187 //l=1.415 //layer=li \
 //thickness=0.1 //x=38.85 //y=5.115 //x2=38.85 //y2=3.7
r201 (  29 32 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=38.85 //y=1.74 //x2=38.85 //y2=3.7
r202 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=38.765 //y=1.655 //x2=38.85 //y2=1.74
r203 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=38.765 //y=1.655 //x2=38.495 //y2=1.655
r204 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.455 //y=5.2 //x2=38.37 //y2=5.2
r205 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=38.765 //y=5.2 //x2=38.85 //y2=5.115
r206 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=38.765 //y=5.2 //x2=38.455 //y2=5.2
r207 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=38.41 //y=1.57 //x2=38.495 //y2=1.655
r208 (  21 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=38.41 //y=1.57 //x2=38.41 //y2=1
r209 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.37 //y=5.285 //x2=38.37 //y2=5.2
r210 (  15 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=38.37 //y=5.285 //x2=38.37 //y2=5.725
r211 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.285 //y=5.2 //x2=38.37 //y2=5.2
r212 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=38.285 //y=5.2 //x2=37.575 //y2=5.2
r213 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=37.49 //y=5.285 //x2=37.575 //y2=5.2
r214 (  7 73 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=37.49 //y=5.285 //x2=37.49 //y2=5.725
r215 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=40.7 //y=3.7 //x2=40.7 //y2=3.7
r216 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=38.85 //y=3.7 //x2=38.85 //y2=3.7
r217 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=38.965 //y=3.7 //x2=38.85 //y2=3.7
r218 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=40.585 //y=3.7 //x2=40.7 //y2=3.7
r219 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=40.585 //y=3.7 //x2=38.965 //y2=3.7
ends PM_TMRDFFQNX1\%noxref_11

subckt PM_TMRDFFQNX1\%noxref_12 ( 1 2 3 4 5 6 16 23 25 35 36 47 49 50 54 55 57 \
 63 66 67 68 69 70 71 72 73 74 75 76 77 78 79 81 87 88 89 90 94 95 96 101 103 \
 105 111 112 113 114 115 120 122 124 130 131 141 142 145 154 155 158 166 168 \
 169 )
c355 ( 169 0 ) capacitor c=0.0220291f //x=34.895 //y=5.02
c356 ( 168 0 ) capacitor c=0.0217503f //x=34.015 //y=5.02
c357 ( 166 0 ) capacitor c=0.00866655f //x=34.89 //y=0.905
c358 ( 158 0 ) capacitor c=0.0331095f //x=41.47 //y=4.7
c359 ( 155 0 ) capacitor c=0.0279499f //x=41.44 //y=1.915
c360 ( 154 0 ) capacitor c=0.0421676f //x=41.44 //y=2.08
c361 ( 145 0 ) capacitor c=0.0331095f //x=31.48 //y=4.7
c362 ( 142 0 ) capacitor c=0.0279499f //x=31.45 //y=1.915
c363 ( 141 0 ) capacitor c=0.0421302f //x=31.45 //y=2.08
c364 ( 131 0 ) capacitor c=0.0429696f //x=42.005 //y=1.25
c365 ( 130 0 ) capacitor c=0.0192208f //x=42.005 //y=0.905
c366 ( 124 0 ) capacitor c=0.0148884f //x=41.85 //y=1.405
c367 ( 122 0 ) capacitor c=0.0157803f //x=41.85 //y=0.75
c368 ( 120 0 ) capacitor c=0.0295235f //x=41.845 //y=4.79
c369 ( 115 0 ) capacitor c=0.0204188f //x=41.475 //y=1.56
c370 ( 114 0 ) capacitor c=0.0168481f //x=41.475 //y=1.25
c371 ( 113 0 ) capacitor c=0.0174783f //x=41.475 //y=0.905
c372 ( 112 0 ) capacitor c=0.0429696f //x=32.015 //y=1.25
c373 ( 111 0 ) capacitor c=0.0192208f //x=32.015 //y=0.905
c374 ( 105 0 ) capacitor c=0.0158629f //x=31.86 //y=1.405
c375 ( 103 0 ) capacitor c=0.0157803f //x=31.86 //y=0.75
c376 ( 101 0 ) capacitor c=0.0295235f //x=31.855 //y=4.79
c377 ( 96 0 ) capacitor c=0.0204188f //x=31.485 //y=1.56
c378 ( 95 0 ) capacitor c=0.0168481f //x=31.485 //y=1.25
c379 ( 94 0 ) capacitor c=0.0174783f //x=31.485 //y=0.905
c380 ( 90 0 ) capacitor c=0.0556143f //x=22.845 //y=4.79
c381 ( 89 0 ) capacitor c=0.0293157f //x=23.135 //y=4.79
c382 ( 88 0 ) capacitor c=0.0347816f //x=22.8 //y=1.22
c383 ( 87 0 ) capacitor c=0.0187487f //x=22.8 //y=0.875
c384 ( 81 0 ) capacitor c=0.0137055f //x=22.645 //y=1.375
c385 ( 79 0 ) capacitor c=0.0149861f //x=22.645 //y=0.72
c386 ( 78 0 ) capacitor c=0.0965296f //x=22.27 //y=1.915
c387 ( 77 0 ) capacitor c=0.0229444f //x=22.27 //y=1.53
c388 ( 76 0 ) capacitor c=0.0234352f //x=22.27 //y=1.22
c389 ( 75 0 ) capacitor c=0.0198724f //x=22.27 //y=0.875
c390 ( 74 0 ) capacitor c=0.15358f //x=41.92 //y=6.02
c391 ( 73 0 ) capacitor c=0.110281f //x=41.48 //y=6.02
c392 ( 72 0 ) capacitor c=0.15358f //x=31.93 //y=6.02
c393 ( 71 0 ) capacitor c=0.110281f //x=31.49 //y=6.02
c394 ( 70 0 ) capacitor c=0.110114f //x=23.21 //y=6.02
c395 ( 69 0 ) capacitor c=0.158956f //x=22.77 //y=6.02
c396 ( 63 0 ) capacitor c=0.00211606f //x=35.04 //y=5.2
c397 ( 57 0 ) capacitor c=0.0711385f //x=41.44 //y=2.08
c398 ( 55 0 ) capacitor c=0.00453889f //x=41.44 //y=4.535
c399 ( 54 0 ) capacitor c=0.105358f //x=35.52 //y=4.07
c400 ( 50 0 ) capacitor c=0.00436419f //x=35.165 //y=1.655
c401 ( 49 0 ) capacitor c=0.0127039f //x=35.435 //y=1.655
c402 ( 47 0 ) capacitor c=0.0137522f //x=35.435 //y=5.2
c403 ( 36 0 ) capacitor c=0.00251459f //x=34.245 //y=5.2
c404 ( 35 0 ) capacitor c=0.0142529f //x=34.955 //y=5.2
c405 ( 25 0 ) capacitor c=0.0699667f //x=31.45 //y=2.08
c406 ( 23 0 ) capacitor c=0.00453889f //x=31.45 //y=4.535
c407 ( 16 0 ) capacitor c=0.103259f //x=22.57 //y=2.08
c408 ( 6 0 ) capacitor c=0.00407792f //x=35.635 //y=4.07
c409 ( 5 0 ) capacitor c=0.0992605f //x=41.325 //y=4.07
c410 ( 4 0 ) capacitor c=0.00412846f //x=31.565 //y=4.07
c411 ( 3 0 ) capacitor c=0.0519266f //x=35.405 //y=4.07
c412 ( 2 0 ) capacitor c=0.0101712f //x=22.685 //y=4.07
c413 ( 1 0 ) capacitor c=0.130427f //x=31.335 //y=4.07
r414 (  160 161 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=41.47 //y=4.79 //x2=41.47 //y2=4.865
r415 (  158 160 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=41.47 //y=4.7 //x2=41.47 //y2=4.79
r416 (  154 155 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=41.44 //y=2.08 //x2=41.44 //y2=1.915
r417 (  147 148 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=31.48 //y=4.79 //x2=31.48 //y2=4.865
r418 (  145 147 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=31.48 //y=4.7 //x2=31.48 //y2=4.79
r419 (  141 142 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=31.45 //y=2.08 //x2=31.45 //y2=1.915
r420 (  131 165 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.005 //y=1.25 //x2=41.965 //y2=1.405
r421 (  130 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.005 //y=0.905 //x2=41.965 //y2=0.75
r422 (  130 131 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=42.005 //y=0.905 //x2=42.005 //y2=1.25
r423 (  125 163 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.63 //y=1.405 //x2=41.515 //y2=1.405
r424 (  124 165 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.85 //y=1.405 //x2=41.965 //y2=1.405
r425 (  123 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.63 //y=0.75 //x2=41.515 //y2=0.75
r426 (  122 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.85 //y=0.75 //x2=41.965 //y2=0.75
r427 (  122 123 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=41.85 //y=0.75 //x2=41.63 //y2=0.75
r428 (  121 160 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=41.605 //y=4.79 //x2=41.47 //y2=4.79
r429 (  120 127 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=41.845 //y=4.79 //x2=41.92 //y2=4.865
r430 (  120 121 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=41.845 //y=4.79 //x2=41.605 //y2=4.79
r431 (  115 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.475 //y=1.56 //x2=41.515 //y2=1.405
r432 (  115 155 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=41.475 //y=1.56 //x2=41.475 //y2=1.915
r433 (  114 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.475 //y=1.25 //x2=41.515 //y2=1.405
r434 (  113 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.475 //y=0.905 //x2=41.515 //y2=0.75
r435 (  113 114 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=41.475 //y=0.905 //x2=41.475 //y2=1.25
r436 (  112 152 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.015 //y=1.25 //x2=31.975 //y2=1.405
r437 (  111 151 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.015 //y=0.905 //x2=31.975 //y2=0.75
r438 (  111 112 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=32.015 //y=0.905 //x2=32.015 //y2=1.25
r439 (  106 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.64 //y=1.405 //x2=31.525 //y2=1.405
r440 (  105 152 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.86 //y=1.405 //x2=31.975 //y2=1.405
r441 (  104 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.64 //y=0.75 //x2=31.525 //y2=0.75
r442 (  103 151 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.86 //y=0.75 //x2=31.975 //y2=0.75
r443 (  103 104 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=31.86 //y=0.75 //x2=31.64 //y2=0.75
r444 (  102 147 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=31.615 //y=4.79 //x2=31.48 //y2=4.79
r445 (  101 108 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=31.855 //y=4.79 //x2=31.93 //y2=4.865
r446 (  101 102 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=31.855 //y=4.79 //x2=31.615 //y2=4.79
r447 (  96 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.485 //y=1.56 //x2=31.525 //y2=1.405
r448 (  96 142 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=31.485 //y=1.56 //x2=31.485 //y2=1.915
r449 (  95 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.485 //y=1.25 //x2=31.525 //y2=1.405
r450 (  94 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.485 //y=0.905 //x2=31.525 //y2=0.75
r451 (  94 95 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=31.485 //y=0.905 //x2=31.485 //y2=1.25
r452 (  89 91 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=23.135 //y=4.79 //x2=23.21 //y2=4.865
r453 (  89 90 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=23.135 //y=4.79 //x2=22.845 //y2=4.79
r454 (  88 139 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.8 //y=1.22 //x2=22.76 //y2=1.375
r455 (  87 138 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.8 //y=0.875 //x2=22.76 //y2=0.72
r456 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.8 //y=0.875 //x2=22.8 //y2=1.22
r457 (  84 90 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=22.77 //y=4.865 //x2=22.845 //y2=4.79
r458 (  84 137 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=22.77 //y=4.865 //x2=22.57 //y2=4.7
r459 (  82 133 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.425 //y=1.375 //x2=22.31 //y2=1.375
r460 (  81 139 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.645 //y=1.375 //x2=22.76 //y2=1.375
r461 (  80 132 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.425 //y=0.72 //x2=22.31 //y2=0.72
r462 (  79 138 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.645 //y=0.72 //x2=22.76 //y2=0.72
r463 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=22.645 //y=0.72 //x2=22.425 //y2=0.72
r464 (  78 135 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=22.27 //y=1.915 //x2=22.57 //y2=2.08
r465 (  77 133 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.27 //y=1.53 //x2=22.31 //y2=1.375
r466 (  77 78 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=22.27 //y=1.53 //x2=22.27 //y2=1.915
r467 (  76 133 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.27 //y=1.22 //x2=22.31 //y2=1.375
r468 (  75 132 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.27 //y=0.875 //x2=22.31 //y2=0.72
r469 (  75 76 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.27 //y=0.875 //x2=22.27 //y2=1.22
r470 (  74 127 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.92 //y=6.02 //x2=41.92 //y2=4.865
r471 (  73 161 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.48 //y=6.02 //x2=41.48 //y2=4.865
r472 (  72 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=31.93 //y=6.02 //x2=31.93 //y2=4.865
r473 (  71 148 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=31.49 //y=6.02 //x2=31.49 //y2=4.865
r474 (  70 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=23.21 //y=6.02 //x2=23.21 //y2=4.865
r475 (  69 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.77 //y=6.02 //x2=22.77 //y2=4.865
r476 (  68 124 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=41.74 //y=1.405 //x2=41.85 //y2=1.405
r477 (  68 125 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=41.74 //y=1.405 //x2=41.63 //y2=1.405
r478 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=31.75 //y=1.405 //x2=31.86 //y2=1.405
r479 (  67 106 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=31.75 //y=1.405 //x2=31.64 //y2=1.405
r480 (  66 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=22.535 //y=1.375 //x2=22.645 //y2=1.375
r481 (  66 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=22.535 //y=1.375 //x2=22.425 //y2=1.375
r482 (  65 158 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=41.47 //y=4.7 //x2=41.47 //y2=4.7
r483 (  62 145 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.48 //y=4.7 //x2=31.48 //y2=4.7
r484 (  57 154 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=41.44 //y=2.08 //x2=41.44 //y2=2.08
r485 (  57 60 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=41.44 //y=2.08 //x2=41.44 //y2=4.07
r486 (  55 65 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=41.44 //y=4.535 //x2=41.455 //y2=4.7
r487 (  55 60 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=41.44 //y=4.535 //x2=41.44 //y2=4.07
r488 (  52 54 ) resistor r=71.5294 //w=0.187 //l=1.045 //layer=li \
 //thickness=0.1 //x=35.52 //y=5.115 //x2=35.52 //y2=4.07
r489 (  51 54 ) resistor r=159.487 //w=0.187 //l=2.33 //layer=li \
 //thickness=0.1 //x=35.52 //y=1.74 //x2=35.52 //y2=4.07
r490 (  49 51 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=35.435 //y=1.655 //x2=35.52 //y2=1.74
r491 (  49 50 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=35.435 //y=1.655 //x2=35.165 //y2=1.655
r492 (  48 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.125 //y=5.2 //x2=35.04 //y2=5.2
r493 (  47 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=35.435 //y=5.2 //x2=35.52 //y2=5.115
r494 (  47 48 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=35.435 //y=5.2 //x2=35.125 //y2=5.2
r495 (  43 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=35.08 //y=1.57 //x2=35.165 //y2=1.655
r496 (  43 166 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=35.08 //y=1.57 //x2=35.08 //y2=1
r497 (  37 63 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.04 //y=5.285 //x2=35.04 //y2=5.2
r498 (  37 169 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=35.04 //y=5.285 //x2=35.04 //y2=5.725
r499 (  35 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.955 //y=5.2 //x2=35.04 //y2=5.2
r500 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=34.955 //y=5.2 //x2=34.245 //y2=5.2
r501 (  29 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=34.16 //y=5.285 //x2=34.245 //y2=5.2
r502 (  29 168 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=34.16 //y=5.285 //x2=34.16 //y2=5.725
r503 (  25 141 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.45 //y=2.08 //x2=31.45 //y2=2.08
r504 (  25 28 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=31.45 //y=2.08 //x2=31.45 //y2=4.07
r505 (  23 62 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=31.45 //y=4.535 //x2=31.465 //y2=4.7
r506 (  23 28 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=31.45 //y=4.535 //x2=31.45 //y2=4.07
r507 (  21 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.57 //y=4.7 //x2=22.57 //y2=4.7
r508 (  19 21 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=22.57 //y=4.07 //x2=22.57 //y2=4.7
r509 (  16 135 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.57 //y=2.08 //x2=22.57 //y2=2.08
r510 (  16 19 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=22.57 //y=2.08 //x2=22.57 //y2=4.07
r511 (  14 60 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=41.44 //y=4.07 //x2=41.44 //y2=4.07
r512 (  12 54 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=35.52 //y=4.07 //x2=35.52 //y2=4.07
r513 (  10 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=31.45 //y=4.07 //x2=31.45 //y2=4.07
r514 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=22.57 //y=4.07 //x2=22.57 //y2=4.07
r515 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=35.635 //y=4.07 //x2=35.52 //y2=4.07
r516 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=41.325 //y=4.07 //x2=41.44 //y2=4.07
r517 (  5 6 ) resistor r=5.42939 //w=0.131 //l=5.69 //layer=m1 \
 //thickness=0.36 //x=41.325 //y=4.07 //x2=35.635 //y2=4.07
r518 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.565 //y=4.07 //x2=31.45 //y2=4.07
r519 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=35.405 //y=4.07 //x2=35.52 //y2=4.07
r520 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=35.405 //y=4.07 //x2=31.565 //y2=4.07
r521 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=22.685 //y=4.07 //x2=22.57 //y2=4.07
r522 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.335 //y=4.07 //x2=31.45 //y2=4.07
r523 (  1 2 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=31.335 //y=4.07 //x2=22.685 //y2=4.07
ends PM_TMRDFFQNX1\%noxref_12

subckt PM_TMRDFFQNX1\%D ( 1 2 3 4 11 12 13 14 15 17 22 24 28 30 40 41 42 43 44 \
 45 46 47 48 49 50 51 56 58 60 66 67 68 69 70 75 77 79 85 86 87 88 89 94 96 98 \
 104 105 107 108 111 120 121 124 133 134 137 )
c424 ( 137 0 ) capacitor c=0.0331095f //x=49.61 //y=4.7
c425 ( 134 0 ) capacitor c=0.0279499f //x=49.58 //y=1.915
c426 ( 133 0 ) capacitor c=0.0421676f //x=49.58 //y=2.08
c427 ( 124 0 ) capacitor c=0.0331095f //x=28.15 //y=4.7
c428 ( 121 0 ) capacitor c=0.0279499f //x=28.12 //y=1.915
c429 ( 120 0 ) capacitor c=0.0421262f //x=28.12 //y=2.08
c430 ( 111 0 ) capacitor c=0.0331095f //x=6.69 //y=4.7
c431 ( 108 0 ) capacitor c=0.0279499f //x=6.66 //y=1.915
c432 ( 107 0 ) capacitor c=0.0421262f //x=6.66 //y=2.08
c433 ( 105 0 ) capacitor c=0.0429696f //x=50.145 //y=1.25
c434 ( 104 0 ) capacitor c=0.0192208f //x=50.145 //y=0.905
c435 ( 98 0 ) capacitor c=0.0148884f //x=49.99 //y=1.405
c436 ( 96 0 ) capacitor c=0.0157803f //x=49.99 //y=0.75
c437 ( 94 0 ) capacitor c=0.0295235f //x=49.985 //y=4.79
c438 ( 89 0 ) capacitor c=0.0204188f //x=49.615 //y=1.56
c439 ( 88 0 ) capacitor c=0.0168481f //x=49.615 //y=1.25
c440 ( 87 0 ) capacitor c=0.0174783f //x=49.615 //y=0.905
c441 ( 86 0 ) capacitor c=0.0429696f //x=28.685 //y=1.25
c442 ( 85 0 ) capacitor c=0.0192208f //x=28.685 //y=0.905
c443 ( 79 0 ) capacitor c=0.0158629f //x=28.53 //y=1.405
c444 ( 77 0 ) capacitor c=0.0157803f //x=28.53 //y=0.75
c445 ( 75 0 ) capacitor c=0.0295235f //x=28.525 //y=4.79
c446 ( 70 0 ) capacitor c=0.0204188f //x=28.155 //y=1.56
c447 ( 69 0 ) capacitor c=0.0168481f //x=28.155 //y=1.25
c448 ( 68 0 ) capacitor c=0.0174783f //x=28.155 //y=0.905
c449 ( 67 0 ) capacitor c=0.0429696f //x=7.225 //y=1.25
c450 ( 66 0 ) capacitor c=0.0192208f //x=7.225 //y=0.905
c451 ( 60 0 ) capacitor c=0.0158629f //x=7.07 //y=1.405
c452 ( 58 0 ) capacitor c=0.0157803f //x=7.07 //y=0.75
c453 ( 56 0 ) capacitor c=0.0295235f //x=7.065 //y=4.79
c454 ( 51 0 ) capacitor c=0.0204188f //x=6.695 //y=1.56
c455 ( 50 0 ) capacitor c=0.0168481f //x=6.695 //y=1.25
c456 ( 49 0 ) capacitor c=0.0174783f //x=6.695 //y=0.905
c457 ( 48 0 ) capacitor c=0.15358f //x=50.06 //y=6.02
c458 ( 47 0 ) capacitor c=0.110281f //x=49.62 //y=6.02
c459 ( 46 0 ) capacitor c=0.15358f //x=28.6 //y=6.02
c460 ( 45 0 ) capacitor c=0.110281f //x=28.16 //y=6.02
c461 ( 44 0 ) capacitor c=0.15358f //x=7.14 //y=6.02
c462 ( 43 0 ) capacitor c=0.110281f //x=6.7 //y=6.02
c463 ( 30 0 ) capacitor c=0.0671606f //x=49.58 //y=2.08
c464 ( 28 0 ) capacitor c=0.00453889f //x=49.58 //y=4.535
c465 ( 24 0 ) capacitor c=0.069138f //x=28.12 //y=2.08
c466 ( 22 0 ) capacitor c=0.00453889f //x=28.12 //y=4.535
c467 ( 17 0 ) capacitor c=0.0711209f //x=6.66 //y=2.08
c468 ( 15 0 ) capacitor c=0.00453889f //x=6.66 //y=4.535
c469 ( 4 0 ) capacitor c=0.0070827f //x=28.235 //y=2.59
c470 ( 3 0 ) capacitor c=0.371601f //x=49.465 //y=2.59
c471 ( 2 0 ) capacitor c=0.0159421f //x=6.775 //y=2.59
c472 ( 1 0 ) capacitor c=0.508623f //x=28.005 //y=2.59
r473 (  139 140 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=49.61 //y=4.79 //x2=49.61 //y2=4.865
r474 (  137 139 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=49.61 //y=4.7 //x2=49.61 //y2=4.79
r475 (  133 134 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=49.58 //y=2.08 //x2=49.58 //y2=1.915
r476 (  126 127 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=28.15 //y=4.79 //x2=28.15 //y2=4.865
r477 (  124 126 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=28.15 //y=4.7 //x2=28.15 //y2=4.79
r478 (  120 121 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=28.12 //y=2.08 //x2=28.12 //y2=1.915
r479 (  113 114 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=6.69 //y=4.79 //x2=6.69 //y2=4.865
r480 (  111 113 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=6.69 //y=4.7 //x2=6.69 //y2=4.79
r481 (  107 108 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.66 //y=2.08 //x2=6.66 //y2=1.915
r482 (  105 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.145 //y=1.25 //x2=50.105 //y2=1.405
r483 (  104 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.145 //y=0.905 //x2=50.105 //y2=0.75
r484 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=50.145 //y=0.905 //x2=50.145 //y2=1.25
r485 (  99 142 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.77 //y=1.405 //x2=49.655 //y2=1.405
r486 (  98 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.99 //y=1.405 //x2=50.105 //y2=1.405
r487 (  97 141 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.77 //y=0.75 //x2=49.655 //y2=0.75
r488 (  96 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.99 //y=0.75 //x2=50.105 //y2=0.75
r489 (  96 97 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=49.99 //y=0.75 //x2=49.77 //y2=0.75
r490 (  95 139 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=49.745 //y=4.79 //x2=49.61 //y2=4.79
r491 (  94 101 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=49.985 //y=4.79 //x2=50.06 //y2=4.865
r492 (  94 95 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=49.985 //y=4.79 //x2=49.745 //y2=4.79
r493 (  89 142 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.615 //y=1.56 //x2=49.655 //y2=1.405
r494 (  89 134 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=49.615 //y=1.56 //x2=49.615 //y2=1.915
r495 (  88 142 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.615 //y=1.25 //x2=49.655 //y2=1.405
r496 (  87 141 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.615 //y=0.905 //x2=49.655 //y2=0.75
r497 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=49.615 //y=0.905 //x2=49.615 //y2=1.25
r498 (  86 131 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.685 //y=1.25 //x2=28.645 //y2=1.405
r499 (  85 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.685 //y=0.905 //x2=28.645 //y2=0.75
r500 (  85 86 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=28.685 //y=0.905 //x2=28.685 //y2=1.25
r501 (  80 129 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.31 //y=1.405 //x2=28.195 //y2=1.405
r502 (  79 131 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.53 //y=1.405 //x2=28.645 //y2=1.405
r503 (  78 128 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.31 //y=0.75 //x2=28.195 //y2=0.75
r504 (  77 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.53 //y=0.75 //x2=28.645 //y2=0.75
r505 (  77 78 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=28.53 //y=0.75 //x2=28.31 //y2=0.75
r506 (  76 126 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=28.285 //y=4.79 //x2=28.15 //y2=4.79
r507 (  75 82 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=28.525 //y=4.79 //x2=28.6 //y2=4.865
r508 (  75 76 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=28.525 //y=4.79 //x2=28.285 //y2=4.79
r509 (  70 129 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.155 //y=1.56 //x2=28.195 //y2=1.405
r510 (  70 121 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=28.155 //y=1.56 //x2=28.155 //y2=1.915
r511 (  69 129 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.155 //y=1.25 //x2=28.195 //y2=1.405
r512 (  68 128 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.155 //y=0.905 //x2=28.195 //y2=0.75
r513 (  68 69 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=28.155 //y=0.905 //x2=28.155 //y2=1.25
r514 (  67 118 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.225 //y=1.25 //x2=7.185 //y2=1.405
r515 (  66 117 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.225 //y=0.905 //x2=7.185 //y2=0.75
r516 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.225 //y=0.905 //x2=7.225 //y2=1.25
r517 (  61 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.85 //y=1.405 //x2=6.735 //y2=1.405
r518 (  60 118 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.07 //y=1.405 //x2=7.185 //y2=1.405
r519 (  59 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.85 //y=0.75 //x2=6.735 //y2=0.75
r520 (  58 117 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.07 //y=0.75 //x2=7.185 //y2=0.75
r521 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.07 //y=0.75 //x2=6.85 //y2=0.75
r522 (  57 113 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=6.825 //y=4.79 //x2=6.69 //y2=4.79
r523 (  56 63 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.065 //y=4.79 //x2=7.14 //y2=4.865
r524 (  56 57 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=7.065 //y=4.79 //x2=6.825 //y2=4.79
r525 (  51 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.695 //y=1.56 //x2=6.735 //y2=1.405
r526 (  51 108 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=6.695 //y=1.56 //x2=6.695 //y2=1.915
r527 (  50 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.695 //y=1.25 //x2=6.735 //y2=1.405
r528 (  49 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.695 //y=0.905 //x2=6.735 //y2=0.75
r529 (  49 50 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.695 //y=0.905 //x2=6.695 //y2=1.25
r530 (  48 101 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=50.06 //y=6.02 //x2=50.06 //y2=4.865
r531 (  47 140 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=49.62 //y=6.02 //x2=49.62 //y2=4.865
r532 (  46 82 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=28.6 //y=6.02 //x2=28.6 //y2=4.865
r533 (  45 127 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=28.16 //y=6.02 //x2=28.16 //y2=4.865
r534 (  44 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.14 //y=6.02 //x2=7.14 //y2=4.865
r535 (  43 114 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.7 //y=6.02 //x2=6.7 //y2=4.865
r536 (  42 98 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=49.88 //y=1.405 //x2=49.99 //y2=1.405
r537 (  42 99 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=49.88 //y=1.405 //x2=49.77 //y2=1.405
r538 (  41 79 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=28.42 //y=1.405 //x2=28.53 //y2=1.405
r539 (  41 80 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=28.42 //y=1.405 //x2=28.31 //y2=1.405
r540 (  40 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.96 //y=1.405 //x2=7.07 //y2=1.405
r541 (  40 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.96 //y=1.405 //x2=6.85 //y2=1.405
r542 (  39 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=49.61 //y=4.7 //x2=49.61 //y2=4.7
r543 (  37 124 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=28.15 //y=4.7 //x2=28.15 //y2=4.7
r544 (  35 111 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.69 //y=4.7 //x2=6.69 //y2=4.7
r545 (  30 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=49.58 //y=2.08 //x2=49.58 //y2=2.08
r546 (  28 39 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=49.58 //y=4.535 //x2=49.595 //y2=4.7
r547 (  24 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=28.12 //y=2.08 //x2=28.12 //y2=2.08
r548 (  22 37 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=28.12 //y=4.535 //x2=28.135 //y2=4.7
r549 (  17 107 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=2.08 //x2=6.66 //y2=2.08
r550 (  15 35 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=6.66 //y=4.535 //x2=6.675 //y2=4.7
r551 (  14 28 ) resistor r=133.134 //w=0.187 //l=1.945 //layer=li \
 //thickness=0.1 //x=49.58 //y=2.59 //x2=49.58 //y2=4.535
r552 (  14 30 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=49.58 //y=2.59 //x2=49.58 //y2=2.08
r553 (  13 22 ) resistor r=133.134 //w=0.187 //l=1.945 //layer=li \
 //thickness=0.1 //x=28.12 //y=2.59 //x2=28.12 //y2=4.535
r554 (  13 24 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=28.12 //y=2.59 //x2=28.12 //y2=2.08
r555 (  12 15 ) resistor r=107.807 //w=0.187 //l=1.575 //layer=li \
 //thickness=0.1 //x=6.66 //y=2.96 //x2=6.66 //y2=4.535
r556 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=6.66 //y=2.59 //x2=6.66 //y2=2.96
r557 (  11 17 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=6.66 //y=2.59 //x2=6.66 //y2=2.08
r558 (  10 14 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=49.58 //y=2.59 //x2=49.58 //y2=2.59
r559 (  8 13 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=28.12 //y=2.59 //x2=28.12 //y2=2.59
r560 (  6 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.66 //y=2.59 //x2=6.66 //y2=2.59
r561 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=28.235 //y=2.59 //x2=28.12 //y2=2.59
r562 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=49.465 //y=2.59 //x2=49.58 //y2=2.59
r563 (  3 4 ) resistor r=20.2576 //w=0.131 //l=21.23 //layer=m1 \
 //thickness=0.36 //x=49.465 //y=2.59 //x2=28.235 //y2=2.59
r564 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.775 //y=2.59 //x2=6.66 //y2=2.59
r565 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=28.005 //y=2.59 //x2=28.12 //y2=2.59
r566 (  1 2 ) resistor r=20.2576 //w=0.131 //l=21.23 //layer=m1 \
 //thickness=0.36 //x=28.005 //y=2.59 //x2=6.775 //y2=2.59
ends PM_TMRDFFQNX1\%D

subckt PM_TMRDFFQNX1\%noxref_14 ( 1 2 3 4 12 25 26 37 39 40 44 46 53 54 55 56 \
 57 58 59 63 64 65 70 72 75 76 77 78 79 80 84 86 89 90 95 96 101 110 113 115 \
 116 )
c233 ( 116 0 ) capacitor c=0.0220291f //x=49.695 //y=5.02
c234 ( 115 0 ) capacitor c=0.0217503f //x=48.815 //y=5.02
c235 ( 113 0 ) capacitor c=0.00866655f //x=49.69 //y=0.905
c236 ( 110 0 ) capacitor c=0.0588816f //x=52.17 //y=4.7
c237 ( 101 0 ) capacitor c=0.058931f //x=46.25 //y=4.7
c238 ( 96 0 ) capacitor c=0.0273931f //x=46.25 //y=1.915
c239 ( 95 0 ) capacitor c=0.0456313f //x=46.25 //y=2.08
c240 ( 90 0 ) capacitor c=0.0318948f //x=52.505 //y=1.21
c241 ( 89 0 ) capacitor c=0.0187384f //x=52.505 //y=0.865
c242 ( 86 0 ) capacitor c=0.0141798f //x=52.35 //y=1.365
c243 ( 84 0 ) capacitor c=0.0149844f //x=52.35 //y=0.71
c244 ( 80 0 ) capacitor c=0.0813322f //x=51.975 //y=1.915
c245 ( 79 0 ) capacitor c=0.0229267f //x=51.975 //y=1.52
c246 ( 78 0 ) capacitor c=0.0234352f //x=51.975 //y=1.21
c247 ( 77 0 ) capacitor c=0.0199343f //x=51.975 //y=0.865
c248 ( 76 0 ) capacitor c=0.0432517f //x=46.77 //y=1.26
c249 ( 75 0 ) capacitor c=0.0200379f //x=46.77 //y=0.915
c250 ( 72 0 ) capacitor c=0.0148873f //x=46.615 //y=1.415
c251 ( 70 0 ) capacitor c=0.0157803f //x=46.615 //y=0.76
c252 ( 65 0 ) capacitor c=0.0218028f //x=46.24 //y=1.57
c253 ( 64 0 ) capacitor c=0.0207459f //x=46.24 //y=1.26
c254 ( 63 0 ) capacitor c=0.0194308f //x=46.24 //y=0.915
c255 ( 59 0 ) capacitor c=0.110275f //x=52.51 //y=6.02
c256 ( 58 0 ) capacitor c=0.154305f //x=52.07 //y=6.02
c257 ( 57 0 ) capacitor c=0.158794f //x=46.43 //y=6.02
c258 ( 56 0 ) capacitor c=0.110114f //x=45.99 //y=6.02
c259 ( 53 0 ) capacitor c=0.00211606f //x=49.84 //y=5.2
c260 ( 46 0 ) capacitor c=0.0862378f //x=52.17 //y=2.08
c261 ( 44 0 ) capacitor c=0.103497f //x=50.32 //y=3.33
c262 ( 40 0 ) capacitor c=0.00404073f //x=49.965 //y=1.655
c263 ( 39 0 ) capacitor c=0.0122201f //x=50.235 //y=1.655
c264 ( 37 0 ) capacitor c=0.0137522f //x=50.235 //y=5.2
c265 ( 26 0 ) capacitor c=0.00251635f //x=49.045 //y=5.2
c266 ( 25 0 ) capacitor c=0.0142423f //x=49.755 //y=5.2
c267 ( 12 0 ) capacitor c=0.0813598f //x=46.25 //y=2.08
c268 ( 4 0 ) capacitor c=0.00280195f //x=50.435 //y=3.33
c269 ( 3 0 ) capacitor c=0.0346903f //x=52.055 //y=3.33
c270 ( 2 0 ) capacitor c=0.0127233f //x=46.365 //y=3.33
c271 ( 1 0 ) capacitor c=0.0559579f //x=50.205 //y=3.33
r272 (  108 110 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=52.07 //y=4.7 //x2=52.17 //y2=4.7
r273 (  95 96 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=46.25 //y=2.08 //x2=46.25 //y2=1.915
r274 (  91 110 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=52.51 //y=4.865 //x2=52.17 //y2=4.7
r275 (  90 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.505 //y=1.21 //x2=52.465 //y2=1.365
r276 (  89 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.505 //y=0.865 //x2=52.465 //y2=0.71
r277 (  89 90 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=52.505 //y=0.865 //x2=52.505 //y2=1.21
r278 (  87 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=52.13 //y=1.365 //x2=52.015 //y2=1.365
r279 (  86 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=52.35 //y=1.365 //x2=52.465 //y2=1.365
r280 (  85 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=52.13 //y=0.71 //x2=52.015 //y2=0.71
r281 (  84 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=52.35 //y=0.71 //x2=52.465 //y2=0.71
r282 (  84 85 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=52.35 //y=0.71 //x2=52.13 //y2=0.71
r283 (  81 108 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=52.07 //y=4.865 //x2=52.07 //y2=4.7
r284 (  80 105 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=51.975 //y=1.915 //x2=52.17 //y2=2.08
r285 (  79 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.975 //y=1.52 //x2=52.015 //y2=1.365
r286 (  79 80 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=51.975 //y=1.52 //x2=51.975 //y2=1.915
r287 (  78 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.975 //y=1.21 //x2=52.015 //y2=1.365
r288 (  77 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.975 //y=0.865 //x2=52.015 //y2=0.71
r289 (  77 78 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=51.975 //y=0.865 //x2=51.975 //y2=1.21
r290 (  76 103 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.77 //y=1.26 //x2=46.73 //y2=1.415
r291 (  75 102 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.77 //y=0.915 //x2=46.73 //y2=0.76
r292 (  75 76 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=46.77 //y=0.915 //x2=46.77 //y2=1.26
r293 (  73 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.395 //y=1.415 //x2=46.28 //y2=1.415
r294 (  72 103 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.615 //y=1.415 //x2=46.73 //y2=1.415
r295 (  71 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.395 //y=0.76 //x2=46.28 //y2=0.76
r296 (  70 102 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.615 //y=0.76 //x2=46.73 //y2=0.76
r297 (  70 71 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=46.615 //y=0.76 //x2=46.395 //y2=0.76
r298 (  67 101 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=46.43 //y=4.865 //x2=46.25 //y2=4.7
r299 (  65 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.24 //y=1.57 //x2=46.28 //y2=1.415
r300 (  65 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=46.24 //y=1.57 //x2=46.24 //y2=1.915
r301 (  64 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.24 //y=1.26 //x2=46.28 //y2=1.415
r302 (  63 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.24 //y=0.915 //x2=46.28 //y2=0.76
r303 (  63 64 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=46.24 //y=0.915 //x2=46.24 //y2=1.26
r304 (  60 101 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=45.99 //y=4.865 //x2=46.25 //y2=4.7
r305 (  59 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=52.51 //y=6.02 //x2=52.51 //y2=4.865
r306 (  58 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=52.07 //y=6.02 //x2=52.07 //y2=4.865
r307 (  57 67 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=46.43 //y=6.02 //x2=46.43 //y2=4.865
r308 (  56 60 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.99 //y=6.02 //x2=45.99 //y2=4.865
r309 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=52.24 //y=1.365 //x2=52.35 //y2=1.365
r310 (  55 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=52.24 //y=1.365 //x2=52.13 //y2=1.365
r311 (  54 72 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=46.505 //y=1.415 //x2=46.615 //y2=1.415
r312 (  54 73 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=46.505 //y=1.415 //x2=46.395 //y2=1.415
r313 (  51 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=52.17 //y=4.7 //x2=52.17 //y2=4.7
r314 (  49 51 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=52.17 //y=3.33 //x2=52.17 //y2=4.7
r315 (  46 105 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=52.17 //y=2.08 //x2=52.17 //y2=2.08
r316 (  46 49 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=52.17 //y=2.08 //x2=52.17 //y2=3.33
r317 (  42 44 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=50.32 //y=5.115 //x2=50.32 //y2=3.33
r318 (  41 44 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=50.32 //y=1.74 //x2=50.32 //y2=3.33
r319 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=50.235 //y=1.655 //x2=50.32 //y2=1.74
r320 (  39 40 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=50.235 //y=1.655 //x2=49.965 //y2=1.655
r321 (  38 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.925 //y=5.2 //x2=49.84 //y2=5.2
r322 (  37 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=50.235 //y=5.2 //x2=50.32 //y2=5.115
r323 (  37 38 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=50.235 //y=5.2 //x2=49.925 //y2=5.2
r324 (  33 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=49.88 //y=1.57 //x2=49.965 //y2=1.655
r325 (  33 113 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=49.88 //y=1.57 //x2=49.88 //y2=1
r326 (  27 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.84 //y=5.285 //x2=49.84 //y2=5.2
r327 (  27 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=49.84 //y=5.285 //x2=49.84 //y2=5.725
r328 (  25 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.755 //y=5.2 //x2=49.84 //y2=5.2
r329 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=49.755 //y=5.2 //x2=49.045 //y2=5.2
r330 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=48.96 //y=5.285 //x2=49.045 //y2=5.2
r331 (  19 115 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=48.96 //y=5.285 //x2=48.96 //y2=5.725
r332 (  17 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=46.25 //y=4.7 //x2=46.25 //y2=4.7
r333 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=46.25 //y=3.33 //x2=46.25 //y2=4.7
r334 (  12 95 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=46.25 //y=2.08 //x2=46.25 //y2=2.08
r335 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=46.25 //y=2.08 //x2=46.25 //y2=3.33
r336 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=52.17 //y=3.33 //x2=52.17 //y2=3.33
r337 (  8 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=50.32 //y=3.33 //x2=50.32 //y2=3.33
r338 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=46.25 //y=3.33 //x2=46.25 //y2=3.33
r339 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=50.435 //y=3.33 //x2=50.32 //y2=3.33
r340 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=52.055 //y=3.33 //x2=52.17 //y2=3.33
r341 (  3 4 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=52.055 //y=3.33 //x2=50.435 //y2=3.33
r342 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=46.365 //y=3.33 //x2=46.25 //y2=3.33
r343 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=50.205 //y=3.33 //x2=50.32 //y2=3.33
r344 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=50.205 //y=3.33 //x2=46.365 //y2=3.33
ends PM_TMRDFFQNX1\%noxref_14

subckt PM_TMRDFFQNX1\%noxref_15 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 \
 47 48 52 54 57 58 68 71 73 74 )
c151 ( 74 0 ) capacitor c=0.0220291f //x=53.025 //y=5.02
c152 ( 73 0 ) capacitor c=0.0217503f //x=52.145 //y=5.02
c153 ( 71 0 ) capacitor c=0.00866655f //x=53.02 //y=0.905
c154 ( 68 0 ) capacitor c=0.0588816f //x=55.5 //y=4.7
c155 ( 58 0 ) capacitor c=0.0318948f //x=55.835 //y=1.21
c156 ( 57 0 ) capacitor c=0.0187384f //x=55.835 //y=0.865
c157 ( 54 0 ) capacitor c=0.0141798f //x=55.68 //y=1.365
c158 ( 52 0 ) capacitor c=0.0149844f //x=55.68 //y=0.71
c159 ( 48 0 ) capacitor c=0.0813322f //x=55.305 //y=1.915
c160 ( 47 0 ) capacitor c=0.0229267f //x=55.305 //y=1.52
c161 ( 46 0 ) capacitor c=0.0234352f //x=55.305 //y=1.21
c162 ( 45 0 ) capacitor c=0.0199343f //x=55.305 //y=0.865
c163 ( 44 0 ) capacitor c=0.110275f //x=55.84 //y=6.02
c164 ( 43 0 ) capacitor c=0.154305f //x=55.4 //y=6.02
c165 ( 41 0 ) capacitor c=0.00211606f //x=53.17 //y=5.2
c166 ( 34 0 ) capacitor c=0.0859022f //x=55.5 //y=2.08
c167 ( 32 0 ) capacitor c=0.104682f //x=53.65 //y=3.33
c168 ( 28 0 ) capacitor c=0.00404073f //x=53.295 //y=1.655
c169 ( 27 0 ) capacitor c=0.0122201f //x=53.565 //y=1.655
c170 ( 25 0 ) capacitor c=0.0137522f //x=53.565 //y=5.2
c171 ( 14 0 ) capacitor c=0.00251459f //x=52.375 //y=5.2
c172 ( 13 0 ) capacitor c=0.0143649f //x=53.085 //y=5.2
c173 ( 2 0 ) capacitor c=0.00668619f //x=53.765 //y=3.33
c174 ( 1 0 ) capacitor c=0.0400514f //x=55.385 //y=3.33
r175 (  66 68 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=55.4 //y=4.7 //x2=55.5 //y2=4.7
r176 (  59 68 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=55.84 //y=4.865 //x2=55.5 //y2=4.7
r177 (  58 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.835 //y=1.21 //x2=55.795 //y2=1.365
r178 (  57 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.835 //y=0.865 //x2=55.795 //y2=0.71
r179 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=55.835 //y=0.865 //x2=55.835 //y2=1.21
r180 (  55 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.46 //y=1.365 //x2=55.345 //y2=1.365
r181 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.68 //y=1.365 //x2=55.795 //y2=1.365
r182 (  53 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.46 //y=0.71 //x2=55.345 //y2=0.71
r183 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.68 //y=0.71 //x2=55.795 //y2=0.71
r184 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=55.68 //y=0.71 //x2=55.46 //y2=0.71
r185 (  49 66 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=55.4 //y=4.865 //x2=55.4 //y2=4.7
r186 (  48 63 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=55.305 //y=1.915 //x2=55.5 //y2=2.08
r187 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.305 //y=1.52 //x2=55.345 //y2=1.365
r188 (  47 48 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=55.305 //y=1.52 //x2=55.305 //y2=1.915
r189 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.305 //y=1.21 //x2=55.345 //y2=1.365
r190 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.305 //y=0.865 //x2=55.345 //y2=0.71
r191 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=55.305 //y=0.865 //x2=55.305 //y2=1.21
r192 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.84 //y=6.02 //x2=55.84 //y2=4.865
r193 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.4 //y=6.02 //x2=55.4 //y2=4.865
r194 (  42 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=55.57 //y=1.365 //x2=55.68 //y2=1.365
r195 (  42 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=55.57 //y=1.365 //x2=55.46 //y2=1.365
r196 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=55.5 //y=4.7 //x2=55.5 //y2=4.7
r197 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=55.5 //y=3.33 //x2=55.5 //y2=4.7
r198 (  34 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=55.5 //y=2.08 //x2=55.5 //y2=2.08
r199 (  34 37 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=55.5 //y=2.08 //x2=55.5 //y2=3.33
r200 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=53.65 //y=5.115 //x2=53.65 //y2=3.33
r201 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=53.65 //y=1.74 //x2=53.65 //y2=3.33
r202 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=53.565 //y=1.655 //x2=53.65 //y2=1.74
r203 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=53.565 //y=1.655 //x2=53.295 //y2=1.655
r204 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.255 //y=5.2 //x2=53.17 //y2=5.2
r205 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=53.565 //y=5.2 //x2=53.65 //y2=5.115
r206 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=53.565 //y=5.2 //x2=53.255 //y2=5.2
r207 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=53.21 //y=1.57 //x2=53.295 //y2=1.655
r208 (  21 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=53.21 //y=1.57 //x2=53.21 //y2=1
r209 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.17 //y=5.285 //x2=53.17 //y2=5.2
r210 (  15 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=53.17 //y=5.285 //x2=53.17 //y2=5.725
r211 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.085 //y=5.2 //x2=53.17 //y2=5.2
r212 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=53.085 //y=5.2 //x2=52.375 //y2=5.2
r213 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=52.29 //y=5.285 //x2=52.375 //y2=5.2
r214 (  7 73 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=52.29 //y=5.285 //x2=52.29 //y2=5.725
r215 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=55.5 //y=3.33 //x2=55.5 //y2=3.33
r216 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=53.65 //y=3.33 //x2=53.65 //y2=3.33
r217 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=53.765 //y=3.33 //x2=53.65 //y2=3.33
r218 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=55.385 //y=3.33 //x2=55.5 //y2=3.33
r219 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=55.385 //y=3.33 //x2=53.765 //y2=3.33
ends PM_TMRDFFQNX1\%noxref_15

subckt PM_TMRDFFQNX1\%CLK ( 1 2 3 4 5 6 7 8 9 10 23 24 25 26 27 28 29 30 31 32 \
 33 34 35 36 37 38 39 40 41 43 54 56 63 72 74 80 89 91 103 104 105 106 107 108 \
 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 125 131 132 133 \
 134 135 140 141 142 147 149 151 157 158 159 160 161 163 169 170 171 172 173 \
 178 179 180 185 187 189 195 196 197 198 199 201 207 208 209 210 211 216 217 \
 218 223 225 227 233 234 238 247 248 251 262 271 272 275 286 295 296 299 )
c752 ( 299 0 ) capacitor c=0.0331838f //x=56.27 //y=4.7
c753 ( 296 0 ) capacitor c=0.0279499f //x=56.24 //y=1.915
c754 ( 295 0 ) capacitor c=0.0421676f //x=56.24 //y=2.08
c755 ( 286 0 ) capacitor c=0.0334842f //x=45.14 //y=4.7
c756 ( 275 0 ) capacitor c=0.0331706f //x=34.81 //y=4.7
c757 ( 272 0 ) capacitor c=0.0279499f //x=34.78 //y=1.915
c758 ( 271 0 ) capacitor c=0.0421302f //x=34.78 //y=2.08
c759 ( 262 0 ) capacitor c=0.0334842f //x=23.68 //y=4.7
c760 ( 251 0 ) capacitor c=0.0331706f //x=13.35 //y=4.7
c761 ( 248 0 ) capacitor c=0.0279499f //x=13.32 //y=1.915
c762 ( 247 0 ) capacitor c=0.0421302f //x=13.32 //y=2.08
c763 ( 238 0 ) capacitor c=0.0334842f //x=2.22 //y=4.7
c764 ( 234 0 ) capacitor c=0.0429696f //x=56.805 //y=1.25
c765 ( 233 0 ) capacitor c=0.0192208f //x=56.805 //y=0.905
c766 ( 227 0 ) capacitor c=0.0148884f //x=56.65 //y=1.405
c767 ( 225 0 ) capacitor c=0.0157803f //x=56.65 //y=0.75
c768 ( 223 0 ) capacitor c=0.0299681f //x=56.645 //y=4.79
c769 ( 218 0 ) capacitor c=0.0205163f //x=56.275 //y=1.56
c770 ( 217 0 ) capacitor c=0.0168481f //x=56.275 //y=1.25
c771 ( 216 0 ) capacitor c=0.0174783f //x=56.275 //y=0.905
c772 ( 211 0 ) capacitor c=0.0245352f //x=45.475 //y=4.79
c773 ( 210 0 ) capacitor c=0.0825763f //x=45.23 //y=1.915
c774 ( 209 0 ) capacitor c=0.0170266f //x=45.23 //y=1.45
c775 ( 208 0 ) capacitor c=0.018609f //x=45.23 //y=1.22
c776 ( 207 0 ) capacitor c=0.0187309f //x=45.23 //y=0.91
c777 ( 201 0 ) capacitor c=0.014725f //x=45.075 //y=1.375
c778 ( 199 0 ) capacitor c=0.0146567f //x=45.075 //y=0.755
c779 ( 198 0 ) capacitor c=0.0335408f //x=44.705 //y=1.22
c780 ( 197 0 ) capacitor c=0.0173761f //x=44.705 //y=0.91
c781 ( 196 0 ) capacitor c=0.0429696f //x=35.345 //y=1.25
c782 ( 195 0 ) capacitor c=0.0192208f //x=35.345 //y=0.905
c783 ( 189 0 ) capacitor c=0.0158629f //x=35.19 //y=1.405
c784 ( 187 0 ) capacitor c=0.0157803f //x=35.19 //y=0.75
c785 ( 185 0 ) capacitor c=0.0295235f //x=35.185 //y=4.79
c786 ( 180 0 ) capacitor c=0.0204188f //x=34.815 //y=1.56
c787 ( 179 0 ) capacitor c=0.0168481f //x=34.815 //y=1.25
c788 ( 178 0 ) capacitor c=0.0174783f //x=34.815 //y=0.905
c789 ( 173 0 ) capacitor c=0.0245352f //x=24.015 //y=4.79
c790 ( 172 0 ) capacitor c=0.0826403f //x=23.77 //y=1.915
c791 ( 171 0 ) capacitor c=0.0170266f //x=23.77 //y=1.45
c792 ( 170 0 ) capacitor c=0.018609f //x=23.77 //y=1.22
c793 ( 169 0 ) capacitor c=0.0187309f //x=23.77 //y=0.91
c794 ( 163 0 ) capacitor c=0.014725f //x=23.615 //y=1.375
c795 ( 161 0 ) capacitor c=0.0146567f //x=23.615 //y=0.755
c796 ( 160 0 ) capacitor c=0.0335408f //x=23.245 //y=1.22
c797 ( 159 0 ) capacitor c=0.0173761f //x=23.245 //y=0.91
c798 ( 158 0 ) capacitor c=0.0429696f //x=13.885 //y=1.25
c799 ( 157 0 ) capacitor c=0.0192208f //x=13.885 //y=0.905
c800 ( 151 0 ) capacitor c=0.0158629f //x=13.73 //y=1.405
c801 ( 149 0 ) capacitor c=0.0157803f //x=13.73 //y=0.75
c802 ( 147 0 ) capacitor c=0.0295269f //x=13.725 //y=4.79
c803 ( 142 0 ) capacitor c=0.0204188f //x=13.355 //y=1.56
c804 ( 141 0 ) capacitor c=0.0168481f //x=13.355 //y=1.25
c805 ( 140 0 ) capacitor c=0.0174783f //x=13.355 //y=0.905
c806 ( 135 0 ) capacitor c=0.0245352f //x=2.555 //y=4.79
c807 ( 134 0 ) capacitor c=0.0850619f //x=2.31 //y=1.915
c808 ( 133 0 ) capacitor c=0.0170266f //x=2.31 //y=1.45
c809 ( 132 0 ) capacitor c=0.018609f //x=2.31 //y=1.22
c810 ( 131 0 ) capacitor c=0.0187309f //x=2.31 //y=0.91
c811 ( 125 0 ) capacitor c=0.014725f //x=2.155 //y=1.375
c812 ( 123 0 ) capacitor c=0.0146567f //x=2.155 //y=0.755
c813 ( 122 0 ) capacitor c=0.0335408f //x=1.785 //y=1.22
c814 ( 121 0 ) capacitor c=0.0173761f //x=1.785 //y=0.91
c815 ( 120 0 ) capacitor c=0.15358f //x=56.72 //y=6.02
c816 ( 119 0 ) capacitor c=0.110281f //x=56.28 //y=6.02
c817 ( 118 0 ) capacitor c=0.110114f //x=45.55 //y=6.02
c818 ( 117 0 ) capacitor c=0.11012f //x=45.11 //y=6.02
c819 ( 116 0 ) capacitor c=0.15358f //x=35.26 //y=6.02
c820 ( 115 0 ) capacitor c=0.110281f //x=34.82 //y=6.02
c821 ( 114 0 ) capacitor c=0.110114f //x=24.09 //y=6.02
c822 ( 113 0 ) capacitor c=0.11012f //x=23.65 //y=6.02
c823 ( 112 0 ) capacitor c=0.15358f //x=13.8 //y=6.02
c824 ( 111 0 ) capacitor c=0.110281f //x=13.36 //y=6.02
c825 ( 110 0 ) capacitor c=0.110114f //x=2.63 //y=6.02
c826 ( 109 0 ) capacitor c=0.11012f //x=2.19 //y=6.02
c827 ( 91 0 ) capacitor c=0.0707124f //x=56.24 //y=2.08
c828 ( 89 0 ) capacitor c=0.00369614f //x=56.24 //y=4.535
c829 ( 80 0 ) capacitor c=0.0921731f //x=45.14 //y=2.08
c830 ( 74 0 ) capacitor c=0.0706586f //x=34.78 //y=2.08
c831 ( 72 0 ) capacitor c=0.00369614f //x=34.78 //y=4.535
c832 ( 63 0 ) capacitor c=0.0948276f //x=23.68 //y=2.08
c833 ( 56 0 ) capacitor c=0.0725839f //x=13.32 //y=2.08
c834 ( 54 0 ) capacitor c=0.00369614f //x=13.32 //y=4.535
c835 ( 43 0 ) capacitor c=0.100158f //x=2.22 //y=2.08
c836 ( 10 0 ) capacitor c=0.00697397f //x=45.255 //y=4.44
c837 ( 9 0 ) capacitor c=0.25424f //x=56.125 //y=4.44
c838 ( 8 0 ) capacitor c=0.00680508f //x=34.895 //y=4.44
c839 ( 7 0 ) capacitor c=0.250892f //x=45.025 //y=4.44
c840 ( 6 0 ) capacitor c=0.184244f //x=23.795 //y=4.44
c841 ( 5 0 ) capacitor c=0.241824f //x=34.665 //y=4.44
c842 ( 4 0 ) capacitor c=0.00759515f //x=13.465 //y=4.442
c843 ( 3 0 ) capacitor c=0.0725822f //x=16.745 //y=4.442
c844 ( 2 0 ) capacitor c=0.0154455f //x=2.335 //y=4.44
c845 ( 1 0 ) capacitor c=0.241824f //x=13.205 //y=4.44
r846 (  301 302 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=56.27 //y=4.79 //x2=56.27 //y2=4.865
r847 (  299 301 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=56.27 //y=4.7 //x2=56.27 //y2=4.79
r848 (  295 296 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=56.24 //y=2.08 //x2=56.24 //y2=1.915
r849 (  288 289 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=45.14 //y=4.79 //x2=45.14 //y2=4.865
r850 (  286 288 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=45.14 //y=4.7 //x2=45.14 //y2=4.79
r851 (  277 278 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=34.81 //y=4.79 //x2=34.81 //y2=4.865
r852 (  275 277 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=34.81 //y=4.7 //x2=34.81 //y2=4.79
r853 (  271 272 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=34.78 //y=2.08 //x2=34.78 //y2=1.915
r854 (  264 265 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=23.68 //y=4.79 //x2=23.68 //y2=4.865
r855 (  262 264 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=23.68 //y=4.7 //x2=23.68 //y2=4.79
r856 (  253 254 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=13.35 //y=4.79 //x2=13.35 //y2=4.865
r857 (  251 253 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=13.35 //y=4.7 //x2=13.35 //y2=4.79
r858 (  247 248 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=13.32 //y=2.08 //x2=13.32 //y2=1.915
r859 (  240 241 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.79 //x2=2.22 //y2=4.865
r860 (  238 240 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.7 //x2=2.22 //y2=4.79
r861 (  234 306 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.805 //y=1.25 //x2=56.765 //y2=1.405
r862 (  233 305 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.805 //y=0.905 //x2=56.765 //y2=0.75
r863 (  233 234 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=56.805 //y=0.905 //x2=56.805 //y2=1.25
r864 (  228 304 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=56.43 //y=1.405 //x2=56.315 //y2=1.405
r865 (  227 306 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=56.65 //y=1.405 //x2=56.765 //y2=1.405
r866 (  226 303 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=56.43 //y=0.75 //x2=56.315 //y2=0.75
r867 (  225 305 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=56.65 //y=0.75 //x2=56.765 //y2=0.75
r868 (  225 226 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=56.65 //y=0.75 //x2=56.43 //y2=0.75
r869 (  224 301 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=56.405 //y=4.79 //x2=56.27 //y2=4.79
r870 (  223 230 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=56.645 //y=4.79 //x2=56.72 //y2=4.865
r871 (  223 224 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=56.645 //y=4.79 //x2=56.405 //y2=4.79
r872 (  218 304 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.275 //y=1.56 //x2=56.315 //y2=1.405
r873 (  218 296 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=56.275 //y=1.56 //x2=56.275 //y2=1.915
r874 (  217 304 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.275 //y=1.25 //x2=56.315 //y2=1.405
r875 (  216 303 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.275 //y=0.905 //x2=56.315 //y2=0.75
r876 (  216 217 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=56.275 //y=0.905 //x2=56.275 //y2=1.25
r877 (  212 288 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=45.275 //y=4.79 //x2=45.14 //y2=4.79
r878 (  211 213 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=45.475 //y=4.79 //x2=45.55 //y2=4.865
r879 (  211 212 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=45.475 //y=4.79 //x2=45.275 //y2=4.79
r880 (  210 293 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=45.23 //y=1.915 //x2=45.155 //y2=2.08
r881 (  209 291 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=45.23 //y=1.45 //x2=45.19 //y2=1.375
r882 (  209 210 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=45.23 //y=1.45 //x2=45.23 //y2=1.915
r883 (  208 291 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.23 //y=1.22 //x2=45.19 //y2=1.375
r884 (  207 290 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.23 //y=0.91 //x2=45.19 //y2=0.755
r885 (  207 208 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=45.23 //y=0.91 //x2=45.23 //y2=1.22
r886 (  202 284 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.86 //y=1.375 //x2=44.745 //y2=1.375
r887 (  201 291 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.075 //y=1.375 //x2=45.19 //y2=1.375
r888 (  200 283 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.86 //y=0.755 //x2=44.745 //y2=0.755
r889 (  199 290 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.075 //y=0.755 //x2=45.19 //y2=0.755
r890 (  199 200 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=45.075 //y=0.755 //x2=44.86 //y2=0.755
r891 (  198 284 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.705 //y=1.22 //x2=44.745 //y2=1.375
r892 (  197 283 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.705 //y=0.91 //x2=44.745 //y2=0.755
r893 (  197 198 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=44.705 //y=0.91 //x2=44.705 //y2=1.22
r894 (  196 282 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.345 //y=1.25 //x2=35.305 //y2=1.405
r895 (  195 281 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.345 //y=0.905 //x2=35.305 //y2=0.75
r896 (  195 196 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=35.345 //y=0.905 //x2=35.345 //y2=1.25
r897 (  190 280 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.97 //y=1.405 //x2=34.855 //y2=1.405
r898 (  189 282 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.19 //y=1.405 //x2=35.305 //y2=1.405
r899 (  188 279 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.97 //y=0.75 //x2=34.855 //y2=0.75
r900 (  187 281 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.19 //y=0.75 //x2=35.305 //y2=0.75
r901 (  187 188 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=35.19 //y=0.75 //x2=34.97 //y2=0.75
r902 (  186 277 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=34.945 //y=4.79 //x2=34.81 //y2=4.79
r903 (  185 192 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=35.185 //y=4.79 //x2=35.26 //y2=4.865
r904 (  185 186 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=35.185 //y=4.79 //x2=34.945 //y2=4.79
r905 (  180 280 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.815 //y=1.56 //x2=34.855 //y2=1.405
r906 (  180 272 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=34.815 //y=1.56 //x2=34.815 //y2=1.915
r907 (  179 280 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.815 //y=1.25 //x2=34.855 //y2=1.405
r908 (  178 279 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.815 //y=0.905 //x2=34.855 //y2=0.75
r909 (  178 179 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=34.815 //y=0.905 //x2=34.815 //y2=1.25
r910 (  174 264 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=23.815 //y=4.79 //x2=23.68 //y2=4.79
r911 (  173 175 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=24.015 //y=4.79 //x2=24.09 //y2=4.865
r912 (  173 174 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=24.015 //y=4.79 //x2=23.815 //y2=4.79
r913 (  172 269 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=23.77 //y=1.915 //x2=23.695 //y2=2.08
r914 (  171 267 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=23.77 //y=1.45 //x2=23.73 //y2=1.375
r915 (  171 172 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=23.77 //y=1.45 //x2=23.77 //y2=1.915
r916 (  170 267 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.77 //y=1.22 //x2=23.73 //y2=1.375
r917 (  169 266 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.77 //y=0.91 //x2=23.73 //y2=0.755
r918 (  169 170 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=23.77 //y=0.91 //x2=23.77 //y2=1.22
r919 (  164 260 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.4 //y=1.375 //x2=23.285 //y2=1.375
r920 (  163 267 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.615 //y=1.375 //x2=23.73 //y2=1.375
r921 (  162 259 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.4 //y=0.755 //x2=23.285 //y2=0.755
r922 (  161 266 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.615 //y=0.755 //x2=23.73 //y2=0.755
r923 (  161 162 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=23.615 //y=0.755 //x2=23.4 //y2=0.755
r924 (  160 260 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.245 //y=1.22 //x2=23.285 //y2=1.375
r925 (  159 259 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.245 //y=0.91 //x2=23.285 //y2=0.755
r926 (  159 160 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=23.245 //y=0.91 //x2=23.245 //y2=1.22
r927 (  158 258 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.885 //y=1.25 //x2=13.845 //y2=1.405
r928 (  157 257 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.885 //y=0.905 //x2=13.845 //y2=0.75
r929 (  157 158 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.885 //y=0.905 //x2=13.885 //y2=1.25
r930 (  152 256 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.51 //y=1.405 //x2=13.395 //y2=1.405
r931 (  151 258 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.73 //y=1.405 //x2=13.845 //y2=1.405
r932 (  150 255 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.51 //y=0.75 //x2=13.395 //y2=0.75
r933 (  149 257 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.73 //y=0.75 //x2=13.845 //y2=0.75
r934 (  149 150 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=13.73 //y=0.75 //x2=13.51 //y2=0.75
r935 (  148 253 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=13.485 //y=4.79 //x2=13.35 //y2=4.79
r936 (  147 154 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=13.725 //y=4.79 //x2=13.8 //y2=4.865
r937 (  147 148 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=13.725 //y=4.79 //x2=13.485 //y2=4.79
r938 (  142 256 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.355 //y=1.56 //x2=13.395 //y2=1.405
r939 (  142 248 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=13.355 //y=1.56 //x2=13.355 //y2=1.915
r940 (  141 256 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.355 //y=1.25 //x2=13.395 //y2=1.405
r941 (  140 255 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.355 //y=0.905 //x2=13.395 //y2=0.75
r942 (  140 141 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.355 //y=0.905 //x2=13.355 //y2=1.25
r943 (  136 240 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.355 //y=4.79 //x2=2.22 //y2=4.79
r944 (  135 137 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.63 //y2=4.865
r945 (  135 136 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.355 //y2=4.79
r946 (  134 245 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.915 //x2=2.235 //y2=2.08
r947 (  133 243 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.27 //y2=1.375
r948 (  133 134 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.31 //y2=1.915
r949 (  132 243 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.22 //x2=2.27 //y2=1.375
r950 (  131 242 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.27 //y2=0.755
r951 (  131 132 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.31 //y2=1.22
r952 (  126 236 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=1.375 //x2=1.825 //y2=1.375
r953 (  125 243 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=1.375 //x2=2.27 //y2=1.375
r954 (  124 235 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=0.755 //x2=1.825 //y2=0.755
r955 (  123 242 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=2.27 //y2=0.755
r956 (  123 124 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=1.94 //y2=0.755
r957 (  122 236 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=1.22 //x2=1.825 //y2=1.375
r958 (  121 235 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.825 //y2=0.755
r959 (  121 122 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.785 //y2=1.22
r960 (  120 230 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=56.72 //y=6.02 //x2=56.72 //y2=4.865
r961 (  119 302 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=56.28 //y=6.02 //x2=56.28 //y2=4.865
r962 (  118 213 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.55 //y=6.02 //x2=45.55 //y2=4.865
r963 (  117 289 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.11 //y=6.02 //x2=45.11 //y2=4.865
r964 (  116 192 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=35.26 //y=6.02 //x2=35.26 //y2=4.865
r965 (  115 278 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=34.82 //y=6.02 //x2=34.82 //y2=4.865
r966 (  114 175 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=24.09 //y=6.02 //x2=24.09 //y2=4.865
r967 (  113 265 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=23.65 //y=6.02 //x2=23.65 //y2=4.865
r968 (  112 154 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.8 //y=6.02 //x2=13.8 //y2=4.865
r969 (  111 254 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.36 //y=6.02 //x2=13.36 //y2=4.865
r970 (  110 137 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.63 //y=6.02 //x2=2.63 //y2=4.865
r971 (  109 241 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.19 //y=6.02 //x2=2.19 //y2=4.865
r972 (  108 227 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=56.54 //y=1.405 //x2=56.65 //y2=1.405
r973 (  108 228 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=56.54 //y=1.405 //x2=56.43 //y2=1.405
r974 (  107 201 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=44.967 //y=1.375 //x2=45.075 //y2=1.375
r975 (  107 202 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=44.967 //y=1.375 //x2=44.86 //y2=1.375
r976 (  106 189 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=35.08 //y=1.405 //x2=35.19 //y2=1.405
r977 (  106 190 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=35.08 //y=1.405 //x2=34.97 //y2=1.405
r978 (  105 163 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=23.507 //y=1.375 //x2=23.615 //y2=1.375
r979 (  105 164 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=23.507 //y=1.375 //x2=23.4 //y2=1.375
r980 (  104 151 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.62 //y=1.405 //x2=13.73 //y2=1.405
r981 (  104 152 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.62 //y=1.405 //x2=13.51 //y2=1.405
r982 (  103 125 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=2.155 //y2=1.375
r983 (  103 126 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=1.94 //y2=1.375
r984 (  102 299 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=56.27 //y=4.7 //x2=56.27 //y2=4.7
r985 (  100 275 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.81 //y=4.7 //x2=34.81 //y2=4.7
r986 (  98 251 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=13.35 //y=4.7 //x2=13.35 //y2=4.7
r987 (  91 295 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=56.24 //y=2.08 //x2=56.24 //y2=2.08
r988 (  89 102 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=56.24 //y=4.535 //x2=56.255 //y2=4.7
r989 (  87 286 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=45.14 //y=4.7 //x2=45.14 //y2=4.7
r990 (  80 293 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=45.14 //y=2.08 //x2=45.14 //y2=2.08
r991 (  74 271 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.78 //y=2.08 //x2=34.78 //y2=2.08
r992 (  72 100 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=34.78 //y=4.535 //x2=34.795 //y2=4.7
r993 (  70 262 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=23.68 //y=4.7 //x2=23.68 //y2=4.7
r994 (  63 269 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=23.68 //y=2.08 //x2=23.68 //y2=2.08
r995 (  56 247 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=13.32 //y=2.08 //x2=13.32 //y2=2.08
r996 (  54 98 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=13.32 //y=4.535 //x2=13.335 //y2=4.7
r997 (  52 238 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=4.7 //x2=2.22 //y2=4.7
r998 (  43 245 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=2.08
r999 (  41 89 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=56.24 //y=4.44 //x2=56.24 //y2=4.535
r1000 (  40 41 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=56.24 //y=3.33 //x2=56.24 //y2=4.44
r1001 (  39 40 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=56.24 //y=2.59 //x2=56.24 //y2=3.33
r1002 (  39 91 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=56.24 //y=2.59 //x2=56.24 //y2=2.08
r1003 (  38 87 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=45.14 //y=4.44 //x2=45.14 //y2=4.7
r1004 (  37 38 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=45.14 //y=3.7 //x2=45.14 //y2=4.44
r1005 (  36 37 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=45.14 //y=3.33 //x2=45.14 //y2=3.7
r1006 (  36 80 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=45.14 //y=3.33 //x2=45.14 //y2=2.08
r1007 (  35 72 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=34.78 //y=4.44 //x2=34.78 //y2=4.535
r1008 (  34 35 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=34.78 //y=3.33 //x2=34.78 //y2=4.44
r1009 (  34 74 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=34.78 //y=3.33 //x2=34.78 //y2=2.08
r1010 (  33 70 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=23.68 //y=4.44 //x2=23.68 //y2=4.7
r1011 (  32 33 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=23.68 //y=3.7 //x2=23.68 //y2=4.44
r1012 (  31 32 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.68 //y=3.33 //x2=23.68 //y2=3.7
r1013 (  31 63 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=23.68 //y=3.33 //x2=23.68 //y2=2.08
r1014 (  30 54 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=13.32 //y=4.44 //x2=13.32 //y2=4.535
r1015 (  29 30 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=13.32 //y=3.33 //x2=13.32 //y2=4.44
r1016 (  28 29 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=13.32 //y=2.96 //x2=13.32 //y2=3.33
r1017 (  28 56 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=13.32 //y=2.96 //x2=13.32 //y2=2.08
r1018 (  27 52 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=2.22 //y=4.44 //x2=2.22 //y2=4.7
r1019 (  26 27 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.7 //x2=2.22 //y2=4.44
r1020 (  25 26 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.33 //x2=2.22 //y2=3.7
r1021 (  24 25 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.96 //x2=2.22 //y2=3.33
r1022 (  23 24 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.59 //x2=2.22 //y2=2.96
r1023 (  23 43 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.59 //x2=2.22 //y2=2.08
r1024 (  22 41 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=56.24 //y=4.44 //x2=56.24 //y2=4.44
r1025 (  20 38 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=45.14 //y=4.44 //x2=45.14 //y2=4.44
r1026 (  18 35 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=34.78 //y=4.44 //x2=34.78 //y2=4.44
r1027 (  16 33 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=23.68 //y=4.44 //x2=23.68 //y2=4.44
r1028 (  14 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=13.32 //y=4.44 //x2=13.32 //y2=4.44
r1029 (  12 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.22 //y=4.44 //x2=2.22 //y2=4.44
r1030 (  10 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=45.255 //y=4.44 //x2=45.14 //y2=4.44
r1031 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=56.125 //y=4.44 //x2=56.24 //y2=4.44
r1032 (  9 10 ) resistor r=10.3721 //w=0.131 //l=10.87 //layer=m1 \
 //thickness=0.36 //x=56.125 //y=4.44 //x2=45.255 //y2=4.44
r1033 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.895 //y=4.44 //x2=34.78 //y2=4.44
r1034 (  7 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=45.025 //y=4.44 //x2=45.14 //y2=4.44
r1035 (  7 8 ) resistor r=9.66603 //w=0.131 //l=10.13 //layer=m1 \
 //thickness=0.36 //x=45.025 //y=4.44 //x2=34.895 //y2=4.44
r1036 (  6 16 ) resistor r=0.0835756 //w=0.172 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.795 //y=4.44 //x2=23.68 //y2=4.44
r1037 (  5 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.665 //y=4.44 //x2=34.78 //y2=4.44
r1038 (  5 6 ) resistor r=10.3721 //w=0.131 //l=10.87 //layer=m1 \
 //thickness=0.36 //x=34.665 //y=4.44 //x2=23.795 //y2=4.44
r1039 (  4 14 ) resistor r=0.0928915 //w=0.224 //l=0.145997 //layer=m1 \
 //thickness=0.36 //x=13.465 //y=4.442 //x2=13.32 //y2=4.44
r1040 (  3 16 ) resistor r=5.04146 //w=0.172 //l=6.936 //layer=m1 \
 //thickness=0.36 //x=16.745 //y=4.442 //x2=23.68 //y2=4.44
r1041 (  3 4 ) resistor r=3.53448 //w=0.116 //l=3.28 //layer=m1 \
 //thickness=0.36 //x=16.745 //y=4.442 //x2=13.465 //y2=4.442
r1042 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.335 //y=4.44 //x2=2.22 //y2=4.44
r1043 (  1 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.205 //y=4.44 //x2=13.32 //y2=4.44
r1044 (  1 2 ) resistor r=10.3721 //w=0.131 //l=10.87 //layer=m1 \
 //thickness=0.36 //x=13.205 //y=4.44 //x2=2.335 //y2=4.44
ends PM_TMRDFFQNX1\%CLK

subckt PM_TMRDFFQNX1\%noxref_17 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 63 \
 64 65 66 67 68 69 70 71 72 76 78 81 82 86 87 88 89 93 95 98 99 109 118 121 \
 123 124 125 )
c255 ( 125 0 ) capacitor c=0.023087f //x=46.065 //y=5.02
c256 ( 124 0 ) capacitor c=0.023519f //x=45.185 //y=5.02
c257 ( 123 0 ) capacitor c=0.0224735f //x=44.305 //y=5.02
c258 ( 121 0 ) capacitor c=0.00872971f //x=46.315 //y=0.915
c259 ( 118 0 ) capacitor c=0.0593152f //x=58.83 //y=4.7
c260 ( 109 0 ) capacitor c=0.0588816f //x=48.84 //y=4.7
c261 ( 99 0 ) capacitor c=0.0318948f //x=59.165 //y=1.21
c262 ( 98 0 ) capacitor c=0.0187384f //x=59.165 //y=0.865
c263 ( 95 0 ) capacitor c=0.0141798f //x=59.01 //y=1.365
c264 ( 93 0 ) capacitor c=0.0149844f //x=59.01 //y=0.71
c265 ( 89 0 ) capacitor c=0.0813322f //x=58.635 //y=1.915
c266 ( 88 0 ) capacitor c=0.0229267f //x=58.635 //y=1.52
c267 ( 87 0 ) capacitor c=0.0234352f //x=58.635 //y=1.21
c268 ( 86 0 ) capacitor c=0.0199343f //x=58.635 //y=0.865
c269 ( 82 0 ) capacitor c=0.0318948f //x=49.175 //y=1.21
c270 ( 81 0 ) capacitor c=0.0187384f //x=49.175 //y=0.865
c271 ( 78 0 ) capacitor c=0.0141798f //x=49.02 //y=1.365
c272 ( 76 0 ) capacitor c=0.0149844f //x=49.02 //y=0.71
c273 ( 72 0 ) capacitor c=0.0813322f //x=48.645 //y=1.915
c274 ( 71 0 ) capacitor c=0.0229267f //x=48.645 //y=1.52
c275 ( 70 0 ) capacitor c=0.0234352f //x=48.645 //y=1.21
c276 ( 69 0 ) capacitor c=0.0199343f //x=48.645 //y=0.865
c277 ( 68 0 ) capacitor c=0.110275f //x=59.17 //y=6.02
c278 ( 67 0 ) capacitor c=0.154305f //x=58.73 //y=6.02
c279 ( 66 0 ) capacitor c=0.110275f //x=49.18 //y=6.02
c280 ( 65 0 ) capacitor c=0.154305f //x=48.74 //y=6.02
c281 ( 62 0 ) capacitor c=0.00106608f //x=46.21 //y=5.155
c282 ( 61 0 ) capacitor c=0.00207162f //x=45.33 //y=5.155
c283 ( 54 0 ) capacitor c=0.0907958f //x=58.83 //y=2.08
c284 ( 46 0 ) capacitor c=0.0836545f //x=48.84 //y=2.08
c285 ( 44 0 ) capacitor c=0.103675f //x=46.99 //y=3.7
c286 ( 40 0 ) capacitor c=0.00398962f //x=46.59 //y=1.665
c287 ( 39 0 ) capacitor c=0.0137288f //x=46.905 //y=1.665
c288 ( 33 0 ) capacitor c=0.0284988f //x=46.905 //y=5.155
c289 ( 25 0 ) capacitor c=0.0176454f //x=46.125 //y=5.155
c290 ( 18 0 ) capacitor c=0.00332903f //x=44.535 //y=5.155
c291 ( 17 0 ) capacitor c=0.014837f //x=45.245 //y=5.155
c292 ( 4 0 ) capacitor c=0.00424317f //x=48.955 //y=3.7
c293 ( 3 0 ) capacitor c=0.159775f //x=58.715 //y=3.7
c294 ( 2 0 ) capacitor c=0.0125346f //x=47.105 //y=3.7
c295 ( 1 0 ) capacitor c=0.0285004f //x=48.725 //y=3.7
r296 (  116 118 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=58.73 //y=4.7 //x2=58.83 //y2=4.7
r297 (  107 109 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=48.74 //y=4.7 //x2=48.84 //y2=4.7
r298 (  100 118 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=59.17 //y=4.865 //x2=58.83 //y2=4.7
r299 (  99 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.165 //y=1.21 //x2=59.125 //y2=1.365
r300 (  98 119 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.165 //y=0.865 //x2=59.125 //y2=0.71
r301 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=59.165 //y=0.865 //x2=59.165 //y2=1.21
r302 (  96 115 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.79 //y=1.365 //x2=58.675 //y2=1.365
r303 (  95 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.01 //y=1.365 //x2=59.125 //y2=1.365
r304 (  94 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.79 //y=0.71 //x2=58.675 //y2=0.71
r305 (  93 119 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.01 //y=0.71 //x2=59.125 //y2=0.71
r306 (  93 94 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=59.01 //y=0.71 //x2=58.79 //y2=0.71
r307 (  90 116 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=58.73 //y=4.865 //x2=58.73 //y2=4.7
r308 (  89 113 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=58.635 //y=1.915 //x2=58.83 //y2=2.08
r309 (  88 115 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.635 //y=1.52 //x2=58.675 //y2=1.365
r310 (  88 89 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=58.635 //y=1.52 //x2=58.635 //y2=1.915
r311 (  87 115 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.635 //y=1.21 //x2=58.675 //y2=1.365
r312 (  86 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.635 //y=0.865 //x2=58.675 //y2=0.71
r313 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=58.635 //y=0.865 //x2=58.635 //y2=1.21
r314 (  83 109 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=49.18 //y=4.865 //x2=48.84 //y2=4.7
r315 (  82 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.175 //y=1.21 //x2=49.135 //y2=1.365
r316 (  81 110 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.175 //y=0.865 //x2=49.135 //y2=0.71
r317 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=49.175 //y=0.865 //x2=49.175 //y2=1.21
r318 (  79 106 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=48.8 //y=1.365 //x2=48.685 //y2=1.365
r319 (  78 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.02 //y=1.365 //x2=49.135 //y2=1.365
r320 (  77 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=48.8 //y=0.71 //x2=48.685 //y2=0.71
r321 (  76 110 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.02 //y=0.71 //x2=49.135 //y2=0.71
r322 (  76 77 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=49.02 //y=0.71 //x2=48.8 //y2=0.71
r323 (  73 107 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=48.74 //y=4.865 //x2=48.74 //y2=4.7
r324 (  72 104 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=48.645 //y=1.915 //x2=48.84 //y2=2.08
r325 (  71 106 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=48.645 //y=1.52 //x2=48.685 //y2=1.365
r326 (  71 72 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=48.645 //y=1.52 //x2=48.645 //y2=1.915
r327 (  70 106 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=48.645 //y=1.21 //x2=48.685 //y2=1.365
r328 (  69 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=48.645 //y=0.865 //x2=48.685 //y2=0.71
r329 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=48.645 //y=0.865 //x2=48.645 //y2=1.21
r330 (  68 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.17 //y=6.02 //x2=59.17 //y2=4.865
r331 (  67 90 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=58.73 //y=6.02 //x2=58.73 //y2=4.865
r332 (  66 83 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=49.18 //y=6.02 //x2=49.18 //y2=4.865
r333 (  65 73 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=48.74 //y=6.02 //x2=48.74 //y2=4.865
r334 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=58.9 //y=1.365 //x2=59.01 //y2=1.365
r335 (  64 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=58.9 //y=1.365 //x2=58.79 //y2=1.365
r336 (  63 78 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=48.91 //y=1.365 //x2=49.02 //y2=1.365
r337 (  63 79 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=48.91 //y=1.365 //x2=48.8 //y2=1.365
r338 (  59 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=58.83 //y=4.7 //x2=58.83 //y2=4.7
r339 (  57 59 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=58.83 //y=3.7 //x2=58.83 //y2=4.7
r340 (  54 113 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=58.83 //y=2.08 //x2=58.83 //y2=2.08
r341 (  54 57 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=58.83 //y=2.08 //x2=58.83 //y2=3.7
r342 (  51 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=48.84 //y=4.7 //x2=48.84 //y2=4.7
r343 (  49 51 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=48.84 //y=3.7 //x2=48.84 //y2=4.7
r344 (  46 104 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=48.84 //y=2.08 //x2=48.84 //y2=2.08
r345 (  46 49 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=48.84 //y=2.08 //x2=48.84 //y2=3.7
r346 (  42 44 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=46.99 //y=5.07 //x2=46.99 //y2=3.7
r347 (  41 44 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=46.99 //y=1.75 //x2=46.99 //y2=3.7
r348 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=46.905 //y=1.665 //x2=46.99 //y2=1.75
r349 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=46.905 //y=1.665 //x2=46.59 //y2=1.665
r350 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=46.505 //y=1.58 //x2=46.59 //y2=1.665
r351 (  35 121 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=46.505 //y=1.58 //x2=46.505 //y2=1.01
r352 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.295 //y=5.155 //x2=46.21 //y2=5.155
r353 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=46.905 //y=5.155 //x2=46.99 //y2=5.07
r354 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=46.905 //y=5.155 //x2=46.295 //y2=5.155
r355 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.21 //y=5.24 //x2=46.21 //y2=5.155
r356 (  27 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.21 //y=5.24 //x2=46.21 //y2=5.725
r357 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.415 //y=5.155 //x2=45.33 //y2=5.155
r358 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.125 //y=5.155 //x2=46.21 //y2=5.155
r359 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=46.125 //y=5.155 //x2=45.415 //y2=5.155
r360 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.33 //y=5.24 //x2=45.33 //y2=5.155
r361 (  19 124 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=45.33 //y=5.24 //x2=45.33 //y2=5.725
r362 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.245 //y=5.155 //x2=45.33 //y2=5.155
r363 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=45.245 //y=5.155 //x2=44.535 //y2=5.155
r364 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=44.45 //y=5.24 //x2=44.535 //y2=5.155
r365 (  11 123 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=44.45 //y=5.24 //x2=44.45 //y2=5.725
r366 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=58.83 //y=3.7 //x2=58.83 //y2=3.7
r367 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=48.84 //y=3.7 //x2=48.84 //y2=3.7
r368 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=46.99 //y=3.7 //x2=46.99 //y2=3.7
r369 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=48.955 //y=3.7 //x2=48.84 //y2=3.7
r370 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=58.715 //y=3.7 //x2=58.83 //y2=3.7
r371 (  3 4 ) resistor r=9.31298 //w=0.131 //l=9.76 //layer=m1 \
 //thickness=0.36 //x=58.715 //y=3.7 //x2=48.955 //y2=3.7
r372 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=47.105 //y=3.7 //x2=46.99 //y2=3.7
r373 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=48.725 //y=3.7 //x2=48.84 //y2=3.7
r374 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=48.725 //y=3.7 //x2=47.105 //y2=3.7
ends PM_TMRDFFQNX1\%noxref_17

subckt PM_TMRDFFQNX1\%noxref_18 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 \
 47 48 52 54 57 58 68 71 73 74 )
c158 ( 74 0 ) capacitor c=0.0220291f //x=59.685 //y=5.02
c159 ( 73 0 ) capacitor c=0.0217503f //x=58.805 //y=5.02
c160 ( 71 0 ) capacitor c=0.00866655f //x=59.68 //y=0.905
c161 ( 68 0 ) capacitor c=0.0591178f //x=62.16 //y=4.7
c162 ( 58 0 ) capacitor c=0.0318948f //x=62.495 //y=1.21
c163 ( 57 0 ) capacitor c=0.0187384f //x=62.495 //y=0.865
c164 ( 54 0 ) capacitor c=0.0141798f //x=62.34 //y=1.365
c165 ( 52 0 ) capacitor c=0.0149844f //x=62.34 //y=0.71
c166 ( 48 0 ) capacitor c=0.0813322f //x=61.965 //y=1.915
c167 ( 47 0 ) capacitor c=0.0229267f //x=61.965 //y=1.52
c168 ( 46 0 ) capacitor c=0.0234352f //x=61.965 //y=1.21
c169 ( 45 0 ) capacitor c=0.0199343f //x=61.965 //y=0.865
c170 ( 44 0 ) capacitor c=0.110275f //x=62.5 //y=6.02
c171 ( 43 0 ) capacitor c=0.154305f //x=62.06 //y=6.02
c172 ( 41 0 ) capacitor c=0.0023043f //x=59.83 //y=5.2
c173 ( 34 0 ) capacitor c=0.0895062f //x=62.16 //y=2.08
c174 ( 32 0 ) capacitor c=0.107504f //x=60.31 //y=4.44
c175 ( 28 0 ) capacitor c=0.00404073f //x=59.955 //y=1.655
c176 ( 27 0 ) capacitor c=0.0122201f //x=60.225 //y=1.655
c177 ( 25 0 ) capacitor c=0.013932f //x=60.225 //y=5.2
c178 ( 14 0 ) capacitor c=0.00265417f //x=59.035 //y=5.2
c179 ( 13 0 ) capacitor c=0.0149571f //x=59.745 //y=5.2
c180 ( 2 0 ) capacitor c=0.0110675f //x=60.425 //y=4.44
c181 ( 1 0 ) capacitor c=0.0525534f //x=62.045 //y=4.44
r182 (  66 68 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=62.06 //y=4.7 //x2=62.16 //y2=4.7
r183 (  59 68 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=62.5 //y=4.865 //x2=62.16 //y2=4.7
r184 (  58 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.495 //y=1.21 //x2=62.455 //y2=1.365
r185 (  57 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.495 //y=0.865 //x2=62.455 //y2=0.71
r186 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=62.495 //y=0.865 //x2=62.495 //y2=1.21
r187 (  55 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=62.12 //y=1.365 //x2=62.005 //y2=1.365
r188 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=62.34 //y=1.365 //x2=62.455 //y2=1.365
r189 (  53 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=62.12 //y=0.71 //x2=62.005 //y2=0.71
r190 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=62.34 //y=0.71 //x2=62.455 //y2=0.71
r191 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=62.34 //y=0.71 //x2=62.12 //y2=0.71
r192 (  49 66 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=62.06 //y=4.865 //x2=62.06 //y2=4.7
r193 (  48 63 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=61.965 //y=1.915 //x2=62.16 //y2=2.08
r194 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.965 //y=1.52 //x2=62.005 //y2=1.365
r195 (  47 48 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=61.965 //y=1.52 //x2=61.965 //y2=1.915
r196 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.965 //y=1.21 //x2=62.005 //y2=1.365
r197 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=61.965 //y=0.865 //x2=62.005 //y2=0.71
r198 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=61.965 //y=0.865 //x2=61.965 //y2=1.21
r199 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=62.5 //y=6.02 //x2=62.5 //y2=4.865
r200 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=62.06 //y=6.02 //x2=62.06 //y2=4.865
r201 (  42 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=62.23 //y=1.365 //x2=62.34 //y2=1.365
r202 (  42 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=62.23 //y=1.365 //x2=62.12 //y2=1.365
r203 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=62.16 //y=4.7 //x2=62.16 //y2=4.7
r204 (  37 39 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=62.16 //y=4.44 //x2=62.16 //y2=4.7
r205 (  34 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=62.16 //y=2.08 //x2=62.16 //y2=2.08
r206 (  34 37 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=62.16 //y=2.08 //x2=62.16 //y2=4.44
r207 (  30 32 ) resistor r=46.2032 //w=0.187 //l=0.675 //layer=li \
 //thickness=0.1 //x=60.31 //y=5.115 //x2=60.31 //y2=4.44
r208 (  29 32 ) resistor r=184.813 //w=0.187 //l=2.7 //layer=li \
 //thickness=0.1 //x=60.31 //y=1.74 //x2=60.31 //y2=4.44
r209 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=60.225 //y=1.655 //x2=60.31 //y2=1.74
r210 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=60.225 //y=1.655 //x2=59.955 //y2=1.655
r211 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.915 //y=5.2 //x2=59.83 //y2=5.2
r212 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=60.225 //y=5.2 //x2=60.31 //y2=5.115
r213 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=60.225 //y=5.2 //x2=59.915 //y2=5.2
r214 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=59.87 //y=1.57 //x2=59.955 //y2=1.655
r215 (  21 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=59.87 //y=1.57 //x2=59.87 //y2=1
r216 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.83 //y=5.285 //x2=59.83 //y2=5.2
r217 (  15 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=59.83 //y=5.285 //x2=59.83 //y2=5.725
r218 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.745 //y=5.2 //x2=59.83 //y2=5.2
r219 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=59.745 //y=5.2 //x2=59.035 //y2=5.2
r220 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=58.95 //y=5.285 //x2=59.035 //y2=5.2
r221 (  7 73 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=58.95 //y=5.285 //x2=58.95 //y2=5.725
r222 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=62.16 //y=4.44 //x2=62.16 //y2=4.44
r223 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=60.31 //y=4.44 //x2=60.31 //y2=4.44
r224 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=60.425 //y=4.44 //x2=60.31 //y2=4.44
r225 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=62.045 //y=4.44 //x2=62.16 //y2=4.44
r226 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=62.045 //y=4.44 //x2=60.425 //y2=4.44
ends PM_TMRDFFQNX1\%noxref_18

subckt PM_TMRDFFQNX1\%noxref_19 ( 1 2 3 4 5 6 16 23 25 35 36 47 49 50 54 55 57 \
 63 66 67 68 69 70 71 72 73 74 75 76 77 78 79 81 87 88 89 90 94 95 96 101 103 \
 105 111 112 113 114 115 120 122 124 130 131 141 142 145 154 155 158 166 168 \
 169 )
c370 ( 169 0 ) capacitor c=0.0220291f //x=56.355 //y=5.02
c371 ( 168 0 ) capacitor c=0.0217503f //x=55.475 //y=5.02
c372 ( 166 0 ) capacitor c=0.00866655f //x=56.35 //y=0.905
c373 ( 158 0 ) capacitor c=0.0333434f //x=62.93 //y=4.7
c374 ( 155 0 ) capacitor c=0.0279499f //x=62.9 //y=1.915
c375 ( 154 0 ) capacitor c=0.0421676f //x=62.9 //y=2.08
c376 ( 145 0 ) capacitor c=0.0331095f //x=52.94 //y=4.7
c377 ( 142 0 ) capacitor c=0.0279499f //x=52.91 //y=1.915
c378 ( 141 0 ) capacitor c=0.0421676f //x=52.91 //y=2.08
c379 ( 131 0 ) capacitor c=0.0429696f //x=63.465 //y=1.25
c380 ( 130 0 ) capacitor c=0.0192208f //x=63.465 //y=0.905
c381 ( 124 0 ) capacitor c=0.0148884f //x=63.31 //y=1.405
c382 ( 122 0 ) capacitor c=0.0157803f //x=63.31 //y=0.75
c383 ( 120 0 ) capacitor c=0.0307199f //x=63.305 //y=4.79
c384 ( 115 0 ) capacitor c=0.0205163f //x=62.935 //y=1.56
c385 ( 114 0 ) capacitor c=0.0168481f //x=62.935 //y=1.25
c386 ( 113 0 ) capacitor c=0.0174783f //x=62.935 //y=0.905
c387 ( 112 0 ) capacitor c=0.0429696f //x=53.475 //y=1.25
c388 ( 111 0 ) capacitor c=0.0192208f //x=53.475 //y=0.905
c389 ( 105 0 ) capacitor c=0.0148884f //x=53.32 //y=1.405
c390 ( 103 0 ) capacitor c=0.0157803f //x=53.32 //y=0.75
c391 ( 101 0 ) capacitor c=0.0295235f //x=53.315 //y=4.79
c392 ( 96 0 ) capacitor c=0.0205163f //x=52.945 //y=1.56
c393 ( 95 0 ) capacitor c=0.0168481f //x=52.945 //y=1.25
c394 ( 94 0 ) capacitor c=0.0174783f //x=52.945 //y=0.905
c395 ( 90 0 ) capacitor c=0.0557698f //x=44.305 //y=4.79
c396 ( 89 0 ) capacitor c=0.0293157f //x=44.595 //y=4.79
c397 ( 88 0 ) capacitor c=0.0347816f //x=44.26 //y=1.22
c398 ( 87 0 ) capacitor c=0.0187487f //x=44.26 //y=0.875
c399 ( 81 0 ) capacitor c=0.0137055f //x=44.105 //y=1.375
c400 ( 79 0 ) capacitor c=0.0149861f //x=44.105 //y=0.72
c401 ( 78 0 ) capacitor c=0.096037f //x=43.73 //y=1.915
c402 ( 77 0 ) capacitor c=0.0228993f //x=43.73 //y=1.53
c403 ( 76 0 ) capacitor c=0.0234352f //x=43.73 //y=1.22
c404 ( 75 0 ) capacitor c=0.0198724f //x=43.73 //y=0.875
c405 ( 74 0 ) capacitor c=0.15358f //x=63.38 //y=6.02
c406 ( 73 0 ) capacitor c=0.110281f //x=62.94 //y=6.02
c407 ( 72 0 ) capacitor c=0.15358f //x=53.39 //y=6.02
c408 ( 71 0 ) capacitor c=0.110281f //x=52.95 //y=6.02
c409 ( 70 0 ) capacitor c=0.110114f //x=44.67 //y=6.02
c410 ( 69 0 ) capacitor c=0.158956f //x=44.23 //y=6.02
c411 ( 63 0 ) capacitor c=0.0023043f //x=56.5 //y=5.2
c412 ( 57 0 ) capacitor c=0.0728897f //x=62.9 //y=2.08
c413 ( 55 0 ) capacitor c=0.00453889f //x=62.9 //y=4.535
c414 ( 54 0 ) capacitor c=0.107708f //x=56.98 //y=4.07
c415 ( 50 0 ) capacitor c=0.00404073f //x=56.625 //y=1.655
c416 ( 49 0 ) capacitor c=0.0122201f //x=56.895 //y=1.655
c417 ( 47 0 ) capacitor c=0.0140419f //x=56.895 //y=5.2
c418 ( 36 0 ) capacitor c=0.00251459f //x=55.705 //y=5.2
c419 ( 35 0 ) capacitor c=0.0143111f //x=56.415 //y=5.2
c420 ( 25 0 ) capacitor c=0.0699131f //x=52.91 //y=2.08
c421 ( 23 0 ) capacitor c=0.00453889f //x=52.91 //y=4.535
c422 ( 16 0 ) capacitor c=0.100766f //x=44.03 //y=2.08
c423 ( 6 0 ) capacitor c=0.00579158f //x=57.095 //y=4.07
c424 ( 5 0 ) capacitor c=0.136665f //x=62.785 //y=4.07
c425 ( 4 0 ) capacitor c=0.00412846f //x=53.025 //y=4.07
c426 ( 3 0 ) capacitor c=0.0575173f //x=56.865 //y=4.07
c427 ( 2 0 ) capacitor c=0.0101712f //x=44.145 //y=4.07
c428 ( 1 0 ) capacitor c=0.130427f //x=52.795 //y=4.07
r429 (  160 161 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=62.93 //y=4.79 //x2=62.93 //y2=4.865
r430 (  158 160 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=62.93 //y=4.7 //x2=62.93 //y2=4.79
r431 (  154 155 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=62.9 //y=2.08 //x2=62.9 //y2=1.915
r432 (  147 148 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=52.94 //y=4.79 //x2=52.94 //y2=4.865
r433 (  145 147 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=52.94 //y=4.7 //x2=52.94 //y2=4.79
r434 (  141 142 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=52.91 //y=2.08 //x2=52.91 //y2=1.915
r435 (  131 165 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.465 //y=1.25 //x2=63.425 //y2=1.405
r436 (  130 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.465 //y=0.905 //x2=63.425 //y2=0.75
r437 (  130 131 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=63.465 //y=0.905 //x2=63.465 //y2=1.25
r438 (  125 163 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.09 //y=1.405 //x2=62.975 //y2=1.405
r439 (  124 165 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.31 //y=1.405 //x2=63.425 //y2=1.405
r440 (  123 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.09 //y=0.75 //x2=62.975 //y2=0.75
r441 (  122 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.31 //y=0.75 //x2=63.425 //y2=0.75
r442 (  122 123 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=63.31 //y=0.75 //x2=63.09 //y2=0.75
r443 (  121 160 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=63.065 //y=4.79 //x2=62.93 //y2=4.79
r444 (  120 127 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=63.305 //y=4.79 //x2=63.38 //y2=4.865
r445 (  120 121 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=63.305 //y=4.79 //x2=63.065 //y2=4.79
r446 (  115 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.935 //y=1.56 //x2=62.975 //y2=1.405
r447 (  115 155 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=62.935 //y=1.56 //x2=62.935 //y2=1.915
r448 (  114 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.935 //y=1.25 //x2=62.975 //y2=1.405
r449 (  113 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.935 //y=0.905 //x2=62.975 //y2=0.75
r450 (  113 114 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=62.935 //y=0.905 //x2=62.935 //y2=1.25
r451 (  112 152 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.475 //y=1.25 //x2=53.435 //y2=1.405
r452 (  111 151 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.475 //y=0.905 //x2=53.435 //y2=0.75
r453 (  111 112 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=53.475 //y=0.905 //x2=53.475 //y2=1.25
r454 (  106 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.1 //y=1.405 //x2=52.985 //y2=1.405
r455 (  105 152 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.32 //y=1.405 //x2=53.435 //y2=1.405
r456 (  104 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.1 //y=0.75 //x2=52.985 //y2=0.75
r457 (  103 151 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.32 //y=0.75 //x2=53.435 //y2=0.75
r458 (  103 104 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=53.32 //y=0.75 //x2=53.1 //y2=0.75
r459 (  102 147 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=53.075 //y=4.79 //x2=52.94 //y2=4.79
r460 (  101 108 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=53.315 //y=4.79 //x2=53.39 //y2=4.865
r461 (  101 102 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=53.315 //y=4.79 //x2=53.075 //y2=4.79
r462 (  96 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.945 //y=1.56 //x2=52.985 //y2=1.405
r463 (  96 142 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=52.945 //y=1.56 //x2=52.945 //y2=1.915
r464 (  95 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.945 //y=1.25 //x2=52.985 //y2=1.405
r465 (  94 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.945 //y=0.905 //x2=52.985 //y2=0.75
r466 (  94 95 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=52.945 //y=0.905 //x2=52.945 //y2=1.25
r467 (  89 91 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=44.595 //y=4.79 //x2=44.67 //y2=4.865
r468 (  89 90 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=44.595 //y=4.79 //x2=44.305 //y2=4.79
r469 (  88 139 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.26 //y=1.22 //x2=44.22 //y2=1.375
r470 (  87 138 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.26 //y=0.875 //x2=44.22 //y2=0.72
r471 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=44.26 //y=0.875 //x2=44.26 //y2=1.22
r472 (  84 90 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=44.23 //y=4.865 //x2=44.305 //y2=4.79
r473 (  84 137 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=44.23 //y=4.865 //x2=44.03 //y2=4.7
r474 (  82 133 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=43.885 //y=1.375 //x2=43.77 //y2=1.375
r475 (  81 139 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.105 //y=1.375 //x2=44.22 //y2=1.375
r476 (  80 132 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=43.885 //y=0.72 //x2=43.77 //y2=0.72
r477 (  79 138 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.105 //y=0.72 //x2=44.22 //y2=0.72
r478 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=44.105 //y=0.72 //x2=43.885 //y2=0.72
r479 (  78 135 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=43.73 //y=1.915 //x2=44.03 //y2=2.08
r480 (  77 133 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=43.73 //y=1.53 //x2=43.77 //y2=1.375
r481 (  77 78 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=43.73 //y=1.53 //x2=43.73 //y2=1.915
r482 (  76 133 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=43.73 //y=1.22 //x2=43.77 //y2=1.375
r483 (  75 132 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=43.73 //y=0.875 //x2=43.77 //y2=0.72
r484 (  75 76 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=43.73 //y=0.875 //x2=43.73 //y2=1.22
r485 (  74 127 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=63.38 //y=6.02 //x2=63.38 //y2=4.865
r486 (  73 161 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=62.94 //y=6.02 //x2=62.94 //y2=4.865
r487 (  72 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=53.39 //y=6.02 //x2=53.39 //y2=4.865
r488 (  71 148 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=52.95 //y=6.02 //x2=52.95 //y2=4.865
r489 (  70 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=44.67 //y=6.02 //x2=44.67 //y2=4.865
r490 (  69 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=44.23 //y=6.02 //x2=44.23 //y2=4.865
r491 (  68 124 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=63.2 //y=1.405 //x2=63.31 //y2=1.405
r492 (  68 125 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=63.2 //y=1.405 //x2=63.09 //y2=1.405
r493 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=53.21 //y=1.405 //x2=53.32 //y2=1.405
r494 (  67 106 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=53.21 //y=1.405 //x2=53.1 //y2=1.405
r495 (  66 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=43.995 //y=1.375 //x2=44.105 //y2=1.375
r496 (  66 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=43.995 //y=1.375 //x2=43.885 //y2=1.375
r497 (  65 158 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=62.93 //y=4.7 //x2=62.93 //y2=4.7
r498 (  62 145 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=52.94 //y=4.7 //x2=52.94 //y2=4.7
r499 (  57 154 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=62.9 //y=2.08 //x2=62.9 //y2=2.08
r500 (  57 60 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=62.9 //y=2.08 //x2=62.9 //y2=4.07
r501 (  55 65 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=62.9 //y=4.535 //x2=62.915 //y2=4.7
r502 (  55 60 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=62.9 //y=4.535 //x2=62.9 //y2=4.07
r503 (  52 54 ) resistor r=71.5294 //w=0.187 //l=1.045 //layer=li \
 //thickness=0.1 //x=56.98 //y=5.115 //x2=56.98 //y2=4.07
r504 (  51 54 ) resistor r=159.487 //w=0.187 //l=2.33 //layer=li \
 //thickness=0.1 //x=56.98 //y=1.74 //x2=56.98 //y2=4.07
r505 (  49 51 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.895 //y=1.655 //x2=56.98 //y2=1.74
r506 (  49 50 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=56.895 //y=1.655 //x2=56.625 //y2=1.655
r507 (  48 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.585 //y=5.2 //x2=56.5 //y2=5.2
r508 (  47 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.895 //y=5.2 //x2=56.98 //y2=5.115
r509 (  47 48 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=56.895 //y=5.2 //x2=56.585 //y2=5.2
r510 (  43 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.54 //y=1.57 //x2=56.625 //y2=1.655
r511 (  43 166 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=56.54 //y=1.57 //x2=56.54 //y2=1
r512 (  37 63 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.5 //y=5.285 //x2=56.5 //y2=5.2
r513 (  37 169 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=56.5 //y=5.285 //x2=56.5 //y2=5.725
r514 (  35 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=56.415 //y=5.2 //x2=56.5 //y2=5.2
r515 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=56.415 //y=5.2 //x2=55.705 //y2=5.2
r516 (  29 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=55.62 //y=5.285 //x2=55.705 //y2=5.2
r517 (  29 168 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=55.62 //y=5.285 //x2=55.62 //y2=5.725
r518 (  25 141 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=52.91 //y=2.08 //x2=52.91 //y2=2.08
r519 (  25 28 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=52.91 //y=2.08 //x2=52.91 //y2=4.07
r520 (  23 62 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=52.91 //y=4.535 //x2=52.925 //y2=4.7
r521 (  23 28 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=52.91 //y=4.535 //x2=52.91 //y2=4.07
r522 (  21 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=44.03 //y=4.7 //x2=44.03 //y2=4.7
r523 (  19 21 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=44.03 //y=4.07 //x2=44.03 //y2=4.7
r524 (  16 135 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=44.03 //y=2.08 //x2=44.03 //y2=2.08
r525 (  16 19 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=44.03 //y=2.08 //x2=44.03 //y2=4.07
r526 (  14 60 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=62.9 //y=4.07 //x2=62.9 //y2=4.07
r527 (  12 54 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=56.98 //y=4.07 //x2=56.98 //y2=4.07
r528 (  10 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=52.91 //y=4.07 //x2=52.91 //y2=4.07
r529 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=44.03 //y=4.07 //x2=44.03 //y2=4.07
r530 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=57.095 //y=4.07 //x2=56.98 //y2=4.07
r531 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=62.785 //y=4.07 //x2=62.9 //y2=4.07
r532 (  5 6 ) resistor r=5.42939 //w=0.131 //l=5.69 //layer=m1 \
 //thickness=0.36 //x=62.785 //y=4.07 //x2=57.095 //y2=4.07
r533 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=53.025 //y=4.07 //x2=52.91 //y2=4.07
r534 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=56.865 //y=4.07 //x2=56.98 //y2=4.07
r535 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=56.865 //y=4.07 //x2=53.025 //y2=4.07
r536 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=44.145 //y=4.07 //x2=44.03 //y2=4.07
r537 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=52.795 //y=4.07 //x2=52.91 //y2=4.07
r538 (  1 2 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=52.795 //y=4.07 //x2=44.145 //y2=4.07
ends PM_TMRDFFQNX1\%noxref_19

subckt PM_TMRDFFQNX1\%noxref_20 ( 1 2 3 4 5 6 17 19 29 30 41 43 44 48 50 60 69 \
 70 71 72 73 74 75 76 77 78 79 80 81 86 88 90 96 97 98 99 100 101 105 107 110 \
 111 112 113 117 118 119 120 124 126 132 133 135 136 139 148 161 164 166 167 )
c344 ( 167 0 ) capacitor c=0.0220235f //x=63.015 //y=5.02
c345 ( 166 0 ) capacitor c=0.0217503f //x=62.135 //y=5.02
c346 ( 164 0 ) capacitor c=0.00864721f //x=63.01 //y=0.905
c347 ( 161 0 ) capacitor c=0.0655948f //x=68.82 //y=4.705
c348 ( 148 0 ) capacitor c=0.0540823f //x=65.12 //y=2.08
c349 ( 139 0 ) capacitor c=0.0331552f //x=59.6 //y=4.7
c350 ( 136 0 ) capacitor c=0.0279499f //x=59.57 //y=1.915
c351 ( 135 0 ) capacitor c=0.0421676f //x=59.57 //y=2.08
c352 ( 133 0 ) capacitor c=0.0342409f //x=69.155 //y=1.21
c353 ( 132 0 ) capacitor c=0.0187384f //x=69.155 //y=0.865
c354 ( 126 0 ) capacitor c=0.0141797f //x=69 //y=1.365
c355 ( 124 0 ) capacitor c=0.0149844f //x=69 //y=0.71
c356 ( 120 0 ) capacitor c=0.0979048f //x=68.625 //y=1.915
c357 ( 119 0 ) capacitor c=0.0225105f //x=68.625 //y=1.52
c358 ( 118 0 ) capacitor c=0.0234376f //x=68.625 //y=1.21
c359 ( 117 0 ) capacitor c=0.0199343f //x=68.625 //y=0.865
c360 ( 113 0 ) capacitor c=0.0318948f //x=65.825 //y=1.21
c361 ( 112 0 ) capacitor c=0.0187384f //x=65.825 //y=0.865
c362 ( 111 0 ) capacitor c=0.0606536f //x=65.465 //y=4.795
c363 ( 110 0 ) capacitor c=0.0292043f //x=65.755 //y=4.795
c364 ( 107 0 ) capacitor c=0.0157913f //x=65.67 //y=1.365
c365 ( 105 0 ) capacitor c=0.0149844f //x=65.67 //y=0.71
c366 ( 101 0 ) capacitor c=0.0302441f //x=65.295 //y=1.915
c367 ( 100 0 ) capacitor c=0.0237559f //x=65.295 //y=1.52
c368 ( 99 0 ) capacitor c=0.0234352f //x=65.295 //y=1.21
c369 ( 98 0 ) capacitor c=0.0199931f //x=65.295 //y=0.865
c370 ( 97 0 ) capacitor c=0.0429696f //x=60.135 //y=1.25
c371 ( 96 0 ) capacitor c=0.0192208f //x=60.135 //y=0.905
c372 ( 90 0 ) capacitor c=0.0148884f //x=59.98 //y=1.405
c373 ( 88 0 ) capacitor c=0.0157803f //x=59.98 //y=0.75
c374 ( 86 0 ) capacitor c=0.0299681f //x=59.975 //y=4.79
c375 ( 81 0 ) capacitor c=0.0205163f //x=59.605 //y=1.56
c376 ( 80 0 ) capacitor c=0.0168481f //x=59.605 //y=1.25
c377 ( 79 0 ) capacitor c=0.0174783f //x=59.605 //y=0.905
c378 ( 78 0 ) capacitor c=0.110336f //x=69.15 //y=6.025
c379 ( 77 0 ) capacitor c=0.154049f //x=68.71 //y=6.025
c380 ( 76 0 ) capacitor c=0.110003f //x=65.83 //y=6.025
c381 ( 75 0 ) capacitor c=0.15424f //x=65.39 //y=6.025
c382 ( 74 0 ) capacitor c=0.15358f //x=60.05 //y=6.02
c383 ( 73 0 ) capacitor c=0.110281f //x=59.61 //y=6.02
c384 ( 69 0 ) capacitor c=0.0024826f //x=63.16 //y=5.2
c385 ( 60 0 ) capacitor c=0.117774f //x=68.82 //y=2.08
c386 ( 50 0 ) capacitor c=0.0959619f //x=65.12 //y=2.08
c387 ( 48 0 ) capacitor c=0.107292f //x=63.64 //y=3.7
c388 ( 44 0 ) capacitor c=0.00404073f //x=63.285 //y=1.655
c389 ( 43 0 ) capacitor c=0.0122201f //x=63.555 //y=1.655
c390 ( 41 0 ) capacitor c=0.0141743f //x=63.555 //y=5.2
c391 ( 30 0 ) capacitor c=0.0025891f //x=62.365 //y=5.2
c392 ( 29 0 ) capacitor c=0.0150834f //x=63.075 //y=5.2
c393 ( 19 0 ) capacitor c=0.0728369f //x=59.57 //y=2.08
c394 ( 17 0 ) capacitor c=0.00453889f //x=59.57 //y=4.535
c395 ( 6 0 ) capacitor c=0.0112191f //x=65.235 //y=4.44
c396 ( 5 0 ) capacitor c=0.0875589f //x=68.705 //y=4.44
c397 ( 4 0 ) capacitor c=0.00444525f //x=63.755 //y=3.7
c398 ( 3 0 ) capacitor c=0.0607201f //x=65.005 //y=3.7
c399 ( 2 0 ) capacitor c=0.00514884f //x=59.685 //y=3.7
c400 ( 1 0 ) capacitor c=0.0734822f //x=63.525 //y=3.7
r401 (  159 161 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=68.71 //y=4.705 //x2=68.82 //y2=4.705
r402 (  141 142 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=59.6 //y=4.79 //x2=59.6 //y2=4.865
r403 (  139 141 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=59.6 //y=4.7 //x2=59.6 //y2=4.79
r404 (  135 136 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=59.57 //y=2.08 //x2=59.57 //y2=1.915
r405 (  133 163 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.155 //y=1.21 //x2=69.115 //y2=1.365
r406 (  132 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.155 //y=0.865 //x2=69.115 //y2=0.71
r407 (  132 133 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=69.155 //y=0.865 //x2=69.155 //y2=1.21
r408 (  129 161 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=69.15 //y=4.87 //x2=68.82 //y2=4.705
r409 (  127 158 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.78 //y=1.365 //x2=68.665 //y2=1.365
r410 (  126 163 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69 //y=1.365 //x2=69.115 //y2=1.365
r411 (  125 157 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.78 //y=0.71 //x2=68.665 //y2=0.71
r412 (  124 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69 //y=0.71 //x2=69.115 //y2=0.71
r413 (  124 125 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=69 //y=0.71 //x2=68.78 //y2=0.71
r414 (  121 159 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=68.71 //y=4.87 //x2=68.71 //y2=4.705
r415 (  120 156 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=68.625 //y=1.915 //x2=68.82 //y2=2.08
r416 (  119 158 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.625 //y=1.52 //x2=68.665 //y2=1.365
r417 (  119 120 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=68.625 //y=1.52 //x2=68.625 //y2=1.915
r418 (  118 158 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.625 //y=1.21 //x2=68.665 //y2=1.365
r419 (  117 157 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.625 //y=0.865 //x2=68.665 //y2=0.71
r420 (  117 118 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=68.625 //y=0.865 //x2=68.625 //y2=1.21
r421 (  113 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.825 //y=1.21 //x2=65.785 //y2=1.365
r422 (  112 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.825 //y=0.865 //x2=65.785 //y2=0.71
r423 (  112 113 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=65.825 //y=0.865 //x2=65.825 //y2=1.21
r424 (  110 114 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=65.755 //y=4.795 //x2=65.83 //y2=4.87
r425 (  110 111 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=65.755 //y=4.795 //x2=65.465 //y2=4.795
r426 (  108 152 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=65.45 //y=1.365 //x2=65.335 //y2=1.365
r427 (  107 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=65.67 //y=1.365 //x2=65.785 //y2=1.365
r428 (  106 151 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=65.45 //y=0.71 //x2=65.335 //y2=0.71
r429 (  105 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=65.67 //y=0.71 //x2=65.785 //y2=0.71
r430 (  105 106 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=65.67 //y=0.71 //x2=65.45 //y2=0.71
r431 (  102 111 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=65.39 //y=4.87 //x2=65.465 //y2=4.795
r432 (  102 150 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=65.39 //y=4.87 //x2=65.12 //y2=4.705
r433 (  101 148 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=65.295 //y=1.915 //x2=65.12 //y2=2.08
r434 (  100 152 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.295 //y=1.52 //x2=65.335 //y2=1.365
r435 (  100 101 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=65.295 //y=1.52 //x2=65.295 //y2=1.915
r436 (  99 152 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.295 //y=1.21 //x2=65.335 //y2=1.365
r437 (  98 151 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.295 //y=0.865 //x2=65.335 //y2=0.71
r438 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=65.295 //y=0.865 //x2=65.295 //y2=1.21
r439 (  97 146 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.135 //y=1.25 //x2=60.095 //y2=1.405
r440 (  96 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.135 //y=0.905 //x2=60.095 //y2=0.75
r441 (  96 97 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=60.135 //y=0.905 //x2=60.135 //y2=1.25
r442 (  91 144 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.76 //y=1.405 //x2=59.645 //y2=1.405
r443 (  90 146 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.98 //y=1.405 //x2=60.095 //y2=1.405
r444 (  89 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.76 //y=0.75 //x2=59.645 //y2=0.75
r445 (  88 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.98 //y=0.75 //x2=60.095 //y2=0.75
r446 (  88 89 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=59.98 //y=0.75 //x2=59.76 //y2=0.75
r447 (  87 141 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=59.735 //y=4.79 //x2=59.6 //y2=4.79
r448 (  86 93 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=59.975 //y=4.79 //x2=60.05 //y2=4.865
r449 (  86 87 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=59.975 //y=4.79 //x2=59.735 //y2=4.79
r450 (  81 144 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.605 //y=1.56 //x2=59.645 //y2=1.405
r451 (  81 136 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=59.605 //y=1.56 //x2=59.605 //y2=1.915
r452 (  80 144 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.605 //y=1.25 //x2=59.645 //y2=1.405
r453 (  79 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.605 //y=0.905 //x2=59.645 //y2=0.75
r454 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=59.605 //y=0.905 //x2=59.605 //y2=1.25
r455 (  78 129 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=69.15 //y=6.025 //x2=69.15 //y2=4.87
r456 (  77 121 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=68.71 //y=6.025 //x2=68.71 //y2=4.87
r457 (  76 114 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=65.83 //y=6.025 //x2=65.83 //y2=4.87
r458 (  75 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=65.39 //y=6.025 //x2=65.39 //y2=4.87
r459 (  74 93 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=60.05 //y=6.02 //x2=60.05 //y2=4.865
r460 (  73 142 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.61 //y=6.02 //x2=59.61 //y2=4.865
r461 (  72 126 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=68.89 //y=1.365 //x2=69 //y2=1.365
r462 (  72 127 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=68.89 //y=1.365 //x2=68.78 //y2=1.365
r463 (  71 107 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=65.56 //y=1.365 //x2=65.67 //y2=1.365
r464 (  71 108 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=65.56 //y=1.365 //x2=65.45 //y2=1.365
r465 (  70 90 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=59.87 //y=1.405 //x2=59.98 //y2=1.405
r466 (  70 91 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=59.87 //y=1.405 //x2=59.76 //y2=1.405
r467 (  68 139 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=59.6 //y=4.7 //x2=59.6 //y2=4.7
r468 (  65 161 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=68.82 //y=4.705 //x2=68.82 //y2=4.705
r469 (  63 65 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=68.82 //y=4.44 //x2=68.82 //y2=4.705
r470 (  60 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=68.82 //y=2.08 //x2=68.82 //y2=2.08
r471 (  60 63 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=68.82 //y=2.08 //x2=68.82 //y2=4.44
r472 (  57 150 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=65.12 //y=4.705 //x2=65.12 //y2=4.705
r473 (  55 57 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=65.12 //y=4.44 //x2=65.12 //y2=4.705
r474 (  53 55 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=65.12 //y=3.7 //x2=65.12 //y2=4.44
r475 (  50 148 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=65.12 //y=2.08 //x2=65.12 //y2=2.08
r476 (  50 53 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=65.12 //y=2.08 //x2=65.12 //y2=3.7
r477 (  46 48 ) resistor r=96.8556 //w=0.187 //l=1.415 //layer=li \
 //thickness=0.1 //x=63.64 //y=5.115 //x2=63.64 //y2=3.7
r478 (  45 48 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=63.64 //y=1.74 //x2=63.64 //y2=3.7
r479 (  43 45 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=63.555 //y=1.655 //x2=63.64 //y2=1.74
r480 (  43 44 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=63.555 //y=1.655 //x2=63.285 //y2=1.655
r481 (  42 69 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.245 //y=5.2 //x2=63.16 //y2=5.2
r482 (  41 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=63.555 //y=5.2 //x2=63.64 //y2=5.115
r483 (  41 42 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=63.555 //y=5.2 //x2=63.245 //y2=5.2
r484 (  37 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=63.2 //y=1.57 //x2=63.285 //y2=1.655
r485 (  37 164 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=63.2 //y=1.57 //x2=63.2 //y2=1
r486 (  31 69 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.16 //y=5.285 //x2=63.16 //y2=5.2
r487 (  31 167 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=63.16 //y=5.285 //x2=63.16 //y2=5.725
r488 (  29 69 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.075 //y=5.2 //x2=63.16 //y2=5.2
r489 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=63.075 //y=5.2 //x2=62.365 //y2=5.2
r490 (  23 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=62.28 //y=5.285 //x2=62.365 //y2=5.2
r491 (  23 166 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=62.28 //y=5.285 //x2=62.28 //y2=5.725
r492 (  19 135 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=59.57 //y=2.08 //x2=59.57 //y2=2.08
r493 (  19 22 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=59.57 //y=2.08 //x2=59.57 //y2=3.7
r494 (  17 68 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=59.57 //y=4.535 //x2=59.585 //y2=4.7
r495 (  17 22 ) resistor r=57.1551 //w=0.187 //l=0.835 //layer=li \
 //thickness=0.1 //x=59.57 //y=4.535 //x2=59.57 //y2=3.7
r496 (  16 63 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=68.82 //y=4.44 //x2=68.82 //y2=4.44
r497 (  14 53 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=65.12 //y=3.7 //x2=65.12 //y2=3.7
r498 (  12 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=65.12 //y=4.44 //x2=65.12 //y2=4.44
r499 (  10 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=63.64 //y=3.7 //x2=63.64 //y2=3.7
r500 (  8 22 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=59.57 //y=3.7 //x2=59.57 //y2=3.7
r501 (  6 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=65.235 //y=4.44 //x2=65.12 //y2=4.44
r502 (  5 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=68.705 //y=4.44 //x2=68.82 //y2=4.44
r503 (  5 6 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=68.705 //y=4.44 //x2=65.235 //y2=4.44
r504 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=63.755 //y=3.7 //x2=63.64 //y2=3.7
r505 (  3 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=65.005 //y=3.7 //x2=65.12 //y2=3.7
r506 (  3 4 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=65.005 //y=3.7 //x2=63.755 //y2=3.7
r507 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=59.685 //y=3.7 //x2=59.57 //y2=3.7
r508 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=63.525 //y=3.7 //x2=63.64 //y2=3.7
r509 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=63.525 //y=3.7 //x2=59.685 //y2=3.7
ends PM_TMRDFFQNX1\%noxref_20

subckt PM_TMRDFFQNX1\%noxref_21 ( 1 2 3 4 5 6 17 19 29 30 41 43 44 48 49 51 59 \
 65 69 72 73 74 75 76 77 78 79 80 81 82 83 88 90 92 98 99 100 101 102 107 109 \
 111 117 118 119 120 121 126 128 130 136 137 139 140 143 152 153 156 164 165 \
 168 176 178 179 )
c502 ( 179 0 ) capacitor c=0.0220291f //x=41.555 //y=5.02
c503 ( 178 0 ) capacitor c=0.0217503f //x=40.675 //y=5.02
c504 ( 176 0 ) capacitor c=0.0084702f //x=41.55 //y=0.905
c505 ( 168 0 ) capacitor c=0.0352016f //x=72.91 //y=4.705
c506 ( 165 0 ) capacitor c=0.0279733f //x=72.89 //y=1.915
c507 ( 164 0 ) capacitor c=0.0467621f //x=72.89 //y=2.08
c508 ( 156 0 ) capacitor c=0.03845f //x=66.27 //y=4.705
c509 ( 153 0 ) capacitor c=0.0300885f //x=66.23 //y=1.915
c510 ( 152 0 ) capacitor c=0.050087f //x=66.23 //y=2.08
c511 ( 143 0 ) capacitor c=0.0331095f //x=38.14 //y=4.7
c512 ( 140 0 ) capacitor c=0.0279499f //x=38.11 //y=1.915
c513 ( 139 0 ) capacitor c=0.0420383f //x=38.11 //y=2.08
c514 ( 137 0 ) capacitor c=0.0237734f //x=73.455 //y=1.255
c515 ( 136 0 ) capacitor c=0.0191782f //x=73.455 //y=0.905
c516 ( 130 0 ) capacitor c=0.0351663f //x=73.3 //y=1.405
c517 ( 128 0 ) capacitor c=0.0157803f //x=73.3 //y=0.75
c518 ( 126 0 ) capacitor c=0.0373879f //x=73.295 //y=4.795
c519 ( 121 0 ) capacitor c=0.0200628f //x=72.925 //y=1.56
c520 ( 120 0 ) capacitor c=0.0168575f //x=72.925 //y=1.255
c521 ( 119 0 ) capacitor c=0.0174993f //x=72.925 //y=0.905
c522 ( 118 0 ) capacitor c=0.0447087f //x=66.795 //y=1.25
c523 ( 117 0 ) capacitor c=0.019286f //x=66.795 //y=0.905
c524 ( 111 0 ) capacitor c=0.0187932f //x=66.64 //y=1.405
c525 ( 109 0 ) capacitor c=0.0157795f //x=66.64 //y=0.75
c526 ( 107 0 ) capacitor c=0.029531f //x=66.635 //y=4.795
c527 ( 102 0 ) capacitor c=0.0206178f //x=66.265 //y=1.56
c528 ( 101 0 ) capacitor c=0.016848f //x=66.265 //y=1.25
c529 ( 100 0 ) capacitor c=0.0174777f //x=66.265 //y=0.905
c530 ( 99 0 ) capacitor c=0.0429696f //x=38.675 //y=1.25
c531 ( 98 0 ) capacitor c=0.0192208f //x=38.675 //y=0.905
c532 ( 92 0 ) capacitor c=0.0148884f //x=38.52 //y=1.405
c533 ( 90 0 ) capacitor c=0.0157803f //x=38.52 //y=0.75
c534 ( 88 0 ) capacitor c=0.0295235f //x=38.515 //y=4.79
c535 ( 83 0 ) capacitor c=0.0204188f //x=38.145 //y=1.56
c536 ( 82 0 ) capacitor c=0.0168481f //x=38.145 //y=1.25
c537 ( 81 0 ) capacitor c=0.0174783f //x=38.145 //y=0.905
c538 ( 80 0 ) capacitor c=0.15325f //x=73.37 //y=6.025
c539 ( 79 0 ) capacitor c=0.110411f //x=72.93 //y=6.025
c540 ( 78 0 ) capacitor c=0.154236f //x=66.71 //y=6.025
c541 ( 77 0 ) capacitor c=0.110294f //x=66.27 //y=6.025
c542 ( 76 0 ) capacitor c=0.15358f //x=38.59 //y=6.02
c543 ( 75 0 ) capacitor c=0.110281f //x=38.15 //y=6.02
c544 ( 69 0 ) capacitor c=0.00501304f //x=72.91 //y=4.705
c545 ( 65 0 ) capacitor c=0.00211606f //x=41.7 //y=5.2
c546 ( 59 0 ) capacitor c=0.0899745f //x=72.89 //y=2.08
c547 ( 51 0 ) capacitor c=0.106138f //x=66.23 //y=2.08
c548 ( 49 0 ) capacitor c=0.00669947f //x=66.23 //y=4.54
c549 ( 48 0 ) capacitor c=0.109862f //x=42.18 //y=2.22
c550 ( 44 0 ) capacitor c=0.00404073f //x=41.825 //y=1.655
c551 ( 43 0 ) capacitor c=0.0122167f //x=42.095 //y=1.655
c552 ( 41 0 ) capacitor c=0.0137995f //x=42.095 //y=5.2
c553 ( 30 0 ) capacitor c=0.00251459f //x=40.905 //y=5.2
c554 ( 29 0 ) capacitor c=0.0143649f //x=41.615 //y=5.2
c555 ( 19 0 ) capacitor c=0.0699202f //x=38.11 //y=2.08
c556 ( 17 0 ) capacitor c=0.00453889f //x=38.11 //y=4.535
c557 ( 6 0 ) capacitor c=0.0111493f //x=66.345 //y=4.07
c558 ( 5 0 ) capacitor c=0.20155f //x=72.775 //y=4.07
c559 ( 4 0 ) capacitor c=0.0053389f //x=42.295 //y=2.22
c560 ( 3 0 ) capacitor c=0.528702f //x=66.115 //y=2.22
c561 ( 2 0 ) capacitor c=0.0141371f //x=38.225 //y=2.22
c562 ( 1 0 ) capacitor c=0.0738364f //x=42.065 //y=2.22
r563 (  170 171 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=72.91 //y=4.795 //x2=72.91 //y2=4.87
r564 (  168 170 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=72.91 //y=4.705 //x2=72.91 //y2=4.795
r565 (  164 165 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=72.89 //y=2.08 //x2=72.89 //y2=1.915
r566 (  156 158 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=66.27 //y=4.705 //x2=66.27 //y2=4.795
r567 (  152 153 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=66.23 //y=2.08 //x2=66.23 //y2=1.915
r568 (  145 146 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=38.14 //y=4.79 //x2=38.14 //y2=4.865
r569 (  143 145 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=38.14 //y=4.7 //x2=38.14 //y2=4.79
r570 (  139 140 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=38.11 //y=2.08 //x2=38.11 //y2=1.915
r571 (  137 175 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=73.455 //y=1.255 //x2=73.455 //y2=1.367
r572 (  136 174 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=73.455 //y=0.905 //x2=73.415 //y2=0.75
r573 (  136 137 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=73.455 //y=0.905 //x2=73.455 //y2=1.255
r574 (  131 173 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.08 //y=1.405 //x2=72.965 //y2=1.405
r575 (  130 175 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=73.3 //y=1.405 //x2=73.455 //y2=1.367
r576 (  129 172 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.08 //y=0.75 //x2=72.965 //y2=0.75
r577 (  128 174 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.3 //y=0.75 //x2=73.415 //y2=0.75
r578 (  128 129 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=73.3 //y=0.75 //x2=73.08 //y2=0.75
r579 (  127 170 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=73.045 //y=4.795 //x2=72.91 //y2=4.795
r580 (  126 133 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=73.295 //y=4.795 //x2=73.37 //y2=4.87
r581 (  126 127 ) resistor r=128.191 //w=0.094 //l=0.25 //layer=ply \
 //thickness=0.18 //x=73.295 //y=4.795 //x2=73.045 //y2=4.795
r582 (  121 173 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.925 //y=1.56 //x2=72.965 //y2=1.405
r583 (  121 165 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=72.925 //y=1.56 //x2=72.925 //y2=1.915
r584 (  120 173 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=72.925 //y=1.255 //x2=72.965 //y2=1.405
r585 (  119 172 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.925 //y=0.905 //x2=72.965 //y2=0.75
r586 (  119 120 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=72.925 //y=0.905 //x2=72.925 //y2=1.255
r587 (  118 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.795 //y=1.25 //x2=66.755 //y2=1.405
r588 (  117 161 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.795 //y=0.905 //x2=66.755 //y2=0.75
r589 (  117 118 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=66.795 //y=0.905 //x2=66.795 //y2=1.25
r590 (  112 160 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.42 //y=1.405 //x2=66.305 //y2=1.405
r591 (  111 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.64 //y=1.405 //x2=66.755 //y2=1.405
r592 (  110 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.42 //y=0.75 //x2=66.305 //y2=0.75
r593 (  109 161 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.64 //y=0.75 //x2=66.755 //y2=0.75
r594 (  109 110 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=66.64 //y=0.75 //x2=66.42 //y2=0.75
r595 (  108 158 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=66.405 //y=4.795 //x2=66.27 //y2=4.795
r596 (  107 114 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=66.635 //y=4.795 //x2=66.71 //y2=4.87
r597 (  107 108 ) resistor r=117.936 //w=0.094 //l=0.23 //layer=ply \
 //thickness=0.18 //x=66.635 //y=4.795 //x2=66.405 //y2=4.795
r598 (  104 158 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=66.27 //y=4.87 //x2=66.27 //y2=4.795
r599 (  102 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.265 //y=1.56 //x2=66.305 //y2=1.405
r600 (  102 153 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=66.265 //y=1.56 //x2=66.265 //y2=1.915
r601 (  101 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.265 //y=1.25 //x2=66.305 //y2=1.405
r602 (  100 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.265 //y=0.905 //x2=66.305 //y2=0.75
r603 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=66.265 //y=0.905 //x2=66.265 //y2=1.25
r604 (  99 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.675 //y=1.25 //x2=38.635 //y2=1.405
r605 (  98 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.675 //y=0.905 //x2=38.635 //y2=0.75
r606 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=38.675 //y=0.905 //x2=38.675 //y2=1.25
r607 (  93 148 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=38.3 //y=1.405 //x2=38.185 //y2=1.405
r608 (  92 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=38.52 //y=1.405 //x2=38.635 //y2=1.405
r609 (  91 147 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=38.3 //y=0.75 //x2=38.185 //y2=0.75
r610 (  90 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=38.52 //y=0.75 //x2=38.635 //y2=0.75
r611 (  90 91 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=38.52 //y=0.75 //x2=38.3 //y2=0.75
r612 (  89 145 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=38.275 //y=4.79 //x2=38.14 //y2=4.79
r613 (  88 95 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=38.515 //y=4.79 //x2=38.59 //y2=4.865
r614 (  88 89 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=38.515 //y=4.79 //x2=38.275 //y2=4.79
r615 (  83 148 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.145 //y=1.56 //x2=38.185 //y2=1.405
r616 (  83 140 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=38.145 //y=1.56 //x2=38.145 //y2=1.915
r617 (  82 148 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.145 //y=1.25 //x2=38.185 //y2=1.405
r618 (  81 147 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.145 //y=0.905 //x2=38.185 //y2=0.75
r619 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=38.145 //y=0.905 //x2=38.145 //y2=1.25
r620 (  80 133 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=73.37 //y=6.025 //x2=73.37 //y2=4.87
r621 (  79 171 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=72.93 //y=6.025 //x2=72.93 //y2=4.87
r622 (  78 114 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=66.71 //y=6.025 //x2=66.71 //y2=4.87
r623 (  77 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=66.27 //y=6.025 //x2=66.27 //y2=4.87
r624 (  76 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=38.59 //y=6.02 //x2=38.59 //y2=4.865
r625 (  75 146 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=38.15 //y=6.02 //x2=38.15 //y2=4.865
r626 (  74 130 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=73.19 //y=1.405 //x2=73.3 //y2=1.405
r627 (  74 131 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=73.19 //y=1.405 //x2=73.08 //y2=1.405
r628 (  73 111 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=66.53 //y=1.405 //x2=66.64 //y2=1.405
r629 (  73 112 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=66.53 //y=1.405 //x2=66.42 //y2=1.405
r630 (  72 92 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=38.41 //y=1.405 //x2=38.52 //y2=1.405
r631 (  72 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=38.41 //y=1.405 //x2=38.3 //y2=1.405
r632 (  69 168 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=72.91 //y=4.705 //x2=72.91 //y2=4.705
r633 (  69 70 ) resistor r=10.3507 //w=0.207 //l=0.165 //layer=li \
 //thickness=0.1 //x=72.9 //y=4.705 //x2=72.9 //y2=4.54
r634 (  67 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=66.27 //y=4.705 //x2=66.27 //y2=4.705
r635 (  64 143 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=38.14 //y=4.7 //x2=38.14 //y2=4.7
r636 (  62 70 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=72.89 //y=4.07 //x2=72.89 //y2=4.54
r637 (  59 164 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=72.89 //y=2.08 //x2=72.89 //y2=2.08
r638 (  59 62 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=72.89 //y=2.08 //x2=72.89 //y2=4.07
r639 (  54 56 ) resistor r=126.631 //w=0.187 //l=1.85 //layer=li \
 //thickness=0.1 //x=66.23 //y=2.22 //x2=66.23 //y2=4.07
r640 (  51 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=66.23 //y=2.08 //x2=66.23 //y2=2.08
r641 (  51 54 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=66.23 //y=2.08 //x2=66.23 //y2=2.22
r642 (  49 67 ) resistor r=11.2426 //w=0.191 //l=0.174714 //layer=li \
 //thickness=0.1 //x=66.23 //y=4.54 //x2=66.25 //y2=4.705
r643 (  49 56 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=66.23 //y=4.54 //x2=66.23 //y2=4.07
r644 (  46 48 ) resistor r=198.16 //w=0.187 //l=2.895 //layer=li \
 //thickness=0.1 //x=42.18 //y=5.115 //x2=42.18 //y2=2.22
r645 (  45 48 ) resistor r=32.8556 //w=0.187 //l=0.48 //layer=li \
 //thickness=0.1 //x=42.18 //y=1.74 //x2=42.18 //y2=2.22
r646 (  43 45 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.095 //y=1.655 //x2=42.18 //y2=1.74
r647 (  43 44 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=42.095 //y=1.655 //x2=41.825 //y2=1.655
r648 (  42 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.785 //y=5.2 //x2=41.7 //y2=5.2
r649 (  41 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.095 //y=5.2 //x2=42.18 //y2=5.115
r650 (  41 42 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=42.095 //y=5.2 //x2=41.785 //y2=5.2
r651 (  37 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=41.74 //y=1.57 //x2=41.825 //y2=1.655
r652 (  37 176 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=41.74 //y=1.57 //x2=41.74 //y2=1
r653 (  31 65 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.7 //y=5.285 //x2=41.7 //y2=5.2
r654 (  31 179 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=41.7 //y=5.285 //x2=41.7 //y2=5.725
r655 (  29 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.615 //y=5.2 //x2=41.7 //y2=5.2
r656 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=41.615 //y=5.2 //x2=40.905 //y2=5.2
r657 (  23 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=40.82 //y=5.285 //x2=40.905 //y2=5.2
r658 (  23 178 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=40.82 //y=5.285 //x2=40.82 //y2=5.725
r659 (  19 139 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=38.11 //y=2.08 //x2=38.11 //y2=2.08
r660 (  19 22 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=38.11 //y=2.08 //x2=38.11 //y2=2.22
r661 (  17 64 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=38.11 //y=4.535 //x2=38.125 //y2=4.7
r662 (  17 22 ) resistor r=158.46 //w=0.187 //l=2.315 //layer=li \
 //thickness=0.1 //x=38.11 //y=4.535 //x2=38.11 //y2=2.22
r663 (  16 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=72.89 //y=4.07 //x2=72.89 //y2=4.07
r664 (  14 54 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=66.23 //y=2.22 //x2=66.23 //y2=2.22
r665 (  12 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=66.23 //y=4.07 //x2=66.23 //y2=4.07
r666 (  10 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=42.18 //y=2.22 //x2=42.18 //y2=2.22
r667 (  8 22 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=38.11 //y=2.22 //x2=38.11 //y2=2.22
r668 (  6 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=66.345 //y=4.07 //x2=66.23 //y2=4.07
r669 (  5 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=72.775 //y=4.07 //x2=72.89 //y2=4.07
r670 (  5 6 ) resistor r=6.1355 //w=0.131 //l=6.43 //layer=m1 //thickness=0.36 \
 //x=72.775 //y=4.07 //x2=66.345 //y2=4.07
r671 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=42.295 //y=2.22 //x2=42.18 //y2=2.22
r672 (  3 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=66.115 //y=2.22 //x2=66.23 //y2=2.22
r673 (  3 4 ) resistor r=22.729 //w=0.131 //l=23.82 //layer=m1 \
 //thickness=0.36 //x=66.115 //y=2.22 //x2=42.295 //y2=2.22
r674 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=38.225 //y=2.22 //x2=38.11 //y2=2.22
r675 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=42.065 //y=2.22 //x2=42.18 //y2=2.22
r676 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=42.065 //y=2.22 //x2=38.225 //y2=2.22
ends PM_TMRDFFQNX1\%noxref_21

subckt PM_TMRDFFQNX1\%noxref_22 ( 1 2 13 14 15 23 29 30 37 50 51 52 53 54 )
c91 ( 54 0 ) capacitor c=0.034295f //x=70.105 //y=5.025
c92 ( 53 0 ) capacitor c=0.0174957f //x=69.225 //y=5.025
c93 ( 51 0 ) capacitor c=0.0214849f //x=66.345 //y=5.025
c94 ( 50 0 ) capacitor c=0.0217161f //x=65.465 //y=5.025
c95 ( 49 0 ) capacitor c=0.00115294f //x=69.37 //y=6.91
c96 ( 37 0 ) capacitor c=0.0131238f //x=70.165 //y=6.91
c97 ( 30 0 ) capacitor c=0.00386507f //x=68.575 //y=6.91
c98 ( 29 0 ) capacitor c=0.00951687f //x=69.285 //y=6.91
c99 ( 23 0 ) capacitor c=0.0455351f //x=68.49 //y=5.21
c100 ( 15 0 ) capacitor c=0.00869404f //x=66.49 //y=5.295
c101 ( 14 0 ) capacitor c=0.00290434f //x=65.695 //y=5.21
c102 ( 13 0 ) capacitor c=0.0139202f //x=66.405 //y=5.21
c103 ( 2 0 ) capacitor c=0.0091252f //x=66.605 //y=5.21
c104 ( 1 0 ) capacitor c=0.0484159f //x=68.375 //y=5.21
r105 (  39 54 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.25 //y=6.825 //x2=70.25 //y2=6.74
r106 (  38 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.455 //y=6.91 //x2=69.37 //y2=6.91
r107 (  37 39 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=70.165 //y=6.91 //x2=70.25 //y2=6.825
r108 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=70.165 //y=6.91 //x2=69.455 //y2=6.91
r109 (  31 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.37 //y=6.825 //x2=69.37 //y2=6.91
r110 (  31 53 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.37 //y=6.825 //x2=69.37 //y2=6.74
r111 (  29 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.285 //y=6.91 //x2=69.37 //y2=6.91
r112 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=69.285 //y=6.91 //x2=68.575 //y2=6.91
r113 (  23 52 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=68.49 //y=5.21 //x2=68.49 //y2=6.06
r114 (  21 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=68.49 //y=6.825 //x2=68.575 //y2=6.91
r115 (  21 52 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.49 //y=6.825 //x2=68.49 //y2=6.74
r116 (  15 48 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=66.49 //y=5.295 //x2=66.49 //y2=5.17
r117 (  15 51 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=66.49 //y=5.295 //x2=66.49 //y2=6.06
r118 (  13 48 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=66.405 //y=5.21 //x2=66.49 //y2=5.17
r119 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=66.405 //y=5.21 //x2=65.695 //y2=5.21
r120 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=65.61 //y=5.295 //x2=65.695 //y2=5.21
r121 (  7 50 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=65.61 //y=5.295 //x2=65.61 //y2=5.72
r122 (  6 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=68.49 //y=5.21 //x2=68.49 //y2=5.21
r123 (  4 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=66.49 //y=5.21 //x2=66.49 //y2=5.21
r124 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=66.605 //y=5.21 //x2=66.49 //y2=5.21
r125 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=68.375 //y=5.21 //x2=68.49 //y2=5.21
r126 (  1 2 ) resistor r=1.68893 //w=0.131 //l=1.77 //layer=m1 \
 //thickness=0.36 //x=68.375 //y=5.21 //x2=66.605 //y2=5.21
ends PM_TMRDFFQNX1\%noxref_22

subckt PM_TMRDFFQNX1\%noxref_23 ( 1 2 3 4 5 6 17 19 29 30 41 43 44 48 50 59 67 \
 68 69 70 71 72 73 74 75 76 77 78 79 84 86 88 94 95 99 100 101 102 103 105 108 \
 111 112 113 114 115 116 117 118 122 124 127 128 129 130 135 136 139 156 163 \
 165 166 )
c459 ( 166 0 ) capacitor c=0.0220291f //x=20.095 //y=5.02
c460 ( 165 0 ) capacitor c=0.0217503f //x=19.215 //y=5.02
c461 ( 163 0 ) capacitor c=0.0084702f //x=20.09 //y=0.905
c462 ( 156 0 ) capacitor c=0.0583848f //x=71.78 //y=2.08
c463 ( 139 0 ) capacitor c=0.0331095f //x=16.68 //y=4.7
c464 ( 136 0 ) capacitor c=0.0279499f //x=16.65 //y=1.915
c465 ( 135 0 ) capacitor c=0.0421302f //x=16.65 //y=2.08
c466 ( 130 0 ) capacitor c=0.0316774f //x=72.485 //y=1.21
c467 ( 129 0 ) capacitor c=0.0187384f //x=72.485 //y=0.865
c468 ( 128 0 ) capacitor c=0.0590362f //x=72.125 //y=4.795
c469 ( 127 0 ) capacitor c=0.0296075f //x=72.415 //y=4.795
c470 ( 124 0 ) capacitor c=0.0157912f //x=72.33 //y=1.365
c471 ( 122 0 ) capacitor c=0.0149844f //x=72.33 //y=0.71
c472 ( 118 0 ) capacitor c=0.0302441f //x=71.955 //y=1.915
c473 ( 117 0 ) capacitor c=0.0234157f //x=71.955 //y=1.52
c474 ( 116 0 ) capacitor c=0.0234376f //x=71.955 //y=1.21
c475 ( 115 0 ) capacitor c=0.0199931f //x=71.955 //y=0.865
c476 ( 114 0 ) capacitor c=0.093437f //x=70.125 //y=1.915
c477 ( 113 0 ) capacitor c=0.0249466f //x=70.125 //y=1.56
c478 ( 112 0 ) capacitor c=0.0234397f //x=70.125 //y=1.25
c479 ( 111 0 ) capacitor c=0.0193195f //x=70.125 //y=0.905
c480 ( 108 0 ) capacitor c=0.0631944f //x=70.03 //y=4.87
c481 ( 105 0 ) capacitor c=0.0187941f //x=69.97 //y=1.405
c482 ( 103 0 ) capacitor c=0.0157803f //x=69.97 //y=0.75
c483 ( 102 0 ) capacitor c=0.010629f //x=69.665 //y=4.795
c484 ( 101 0 ) capacitor c=0.0194269f //x=69.955 //y=4.795
c485 ( 100 0 ) capacitor c=0.0365717f //x=69.595 //y=1.25
c486 ( 99 0 ) capacitor c=0.0175988f //x=69.595 //y=0.905
c487 ( 95 0 ) capacitor c=0.0429696f //x=17.215 //y=1.25
c488 ( 94 0 ) capacitor c=0.0192208f //x=17.215 //y=0.905
c489 ( 88 0 ) capacitor c=0.0158629f //x=17.06 //y=1.405
c490 ( 86 0 ) capacitor c=0.0157803f //x=17.06 //y=0.75
c491 ( 84 0 ) capacitor c=0.0295235f //x=17.055 //y=4.79
c492 ( 79 0 ) capacitor c=0.0204188f //x=16.685 //y=1.56
c493 ( 78 0 ) capacitor c=0.0168481f //x=16.685 //y=1.25
c494 ( 77 0 ) capacitor c=0.0174783f //x=16.685 //y=0.905
c495 ( 76 0 ) capacitor c=0.110622f //x=72.49 //y=6.025
c496 ( 75 0 ) capacitor c=0.154068f //x=72.05 //y=6.025
c497 ( 74 0 ) capacitor c=0.154291f //x=70.03 //y=6.025
c498 ( 73 0 ) capacitor c=0.110404f //x=69.59 //y=6.025
c499 ( 72 0 ) capacitor c=0.15358f //x=17.13 //y=6.02
c500 ( 71 0 ) capacitor c=0.110281f //x=16.69 //y=6.02
c501 ( 67 0 ) capacitor c=0.00211606f //x=20.24 //y=5.2
c502 ( 59 0 ) capacitor c=0.100881f //x=71.78 //y=2.08
c503 ( 50 0 ) capacitor c=0.105664f //x=70.3 //y=2.08
c504 ( 48 0 ) capacitor c=0.110619f //x=20.72 //y=2.96
c505 ( 44 0 ) capacitor c=0.00436419f //x=20.365 //y=1.655
c506 ( 43 0 ) capacitor c=0.0127039f //x=20.635 //y=1.655
c507 ( 41 0 ) capacitor c=0.0137995f //x=20.635 //y=5.2
c508 ( 30 0 ) capacitor c=0.00251459f //x=19.445 //y=5.2
c509 ( 29 0 ) capacitor c=0.0143649f //x=20.155 //y=5.2
c510 ( 19 0 ) capacitor c=0.0718857f //x=16.65 //y=2.08
c511 ( 17 0 ) capacitor c=0.00453889f //x=16.65 //y=4.535
c512 ( 6 0 ) capacitor c=0.0100496f //x=70.415 //y=2.08
c513 ( 5 0 ) capacitor c=0.0462526f //x=71.665 //y=2.08
c514 ( 4 0 ) capacitor c=0.00475948f //x=20.835 //y=2.96
c515 ( 3 0 ) capacitor c=0.950065f //x=70.185 //y=2.96
c516 ( 2 0 ) capacitor c=0.0130562f //x=16.765 //y=2.96
c517 ( 1 0 ) capacitor c=0.0719815f //x=20.605 //y=2.96
r518 (  141 142 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=16.68 //y=4.79 //x2=16.68 //y2=4.865
r519 (  139 141 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=16.68 //y=4.7 //x2=16.68 //y2=4.79
r520 (  135 136 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=16.65 //y=2.08 //x2=16.65 //y2=1.915
r521 (  130 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.485 //y=1.21 //x2=72.445 //y2=1.365
r522 (  129 161 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.485 //y=0.865 //x2=72.445 //y2=0.71
r523 (  129 130 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=72.485 //y=0.865 //x2=72.485 //y2=1.21
r524 (  127 131 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=72.415 //y=4.795 //x2=72.49 //y2=4.87
r525 (  127 128 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=72.415 //y=4.795 //x2=72.125 //y2=4.795
r526 (  125 160 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=72.11 //y=1.365 //x2=71.995 //y2=1.365
r527 (  124 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=72.33 //y=1.365 //x2=72.445 //y2=1.365
r528 (  123 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=72.11 //y=0.71 //x2=71.995 //y2=0.71
r529 (  122 161 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=72.33 //y=0.71 //x2=72.445 //y2=0.71
r530 (  122 123 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=72.33 //y=0.71 //x2=72.11 //y2=0.71
r531 (  119 128 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=72.05 //y=4.87 //x2=72.125 //y2=4.795
r532 (  119 158 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=72.05 //y=4.87 //x2=71.78 //y2=4.705
r533 (  118 156 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=71.955 //y=1.915 //x2=71.78 //y2=2.08
r534 (  117 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.955 //y=1.52 //x2=71.995 //y2=1.365
r535 (  117 118 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=71.955 //y=1.52 //x2=71.955 //y2=1.915
r536 (  116 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.955 //y=1.21 //x2=71.995 //y2=1.365
r537 (  115 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.955 //y=0.865 //x2=71.995 //y2=0.71
r538 (  115 116 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=71.955 //y=0.865 //x2=71.955 //y2=1.21
r539 (  114 152 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=70.125 //y=1.915 //x2=70.3 //y2=2.08
r540 (  113 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.125 //y=1.56 //x2=70.085 //y2=1.405
r541 (  113 114 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=70.125 //y=1.56 //x2=70.125 //y2=1.915
r542 (  112 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.125 //y=1.25 //x2=70.085 //y2=1.405
r543 (  111 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.125 //y=0.905 //x2=70.085 //y2=0.75
r544 (  111 112 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=70.125 //y=0.905 //x2=70.125 //y2=1.25
r545 (  108 154 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=70.03 //y=4.87 //x2=70.3 //y2=4.705
r546 (  106 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.75 //y=1.405 //x2=69.635 //y2=1.405
r547 (  105 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.97 //y=1.405 //x2=70.085 //y2=1.405
r548 (  104 147 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.75 //y=0.75 //x2=69.635 //y2=0.75
r549 (  103 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.97 //y=0.75 //x2=70.085 //y2=0.75
r550 (  103 104 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=69.97 //y=0.75 //x2=69.75 //y2=0.75
r551 (  101 108 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=69.955 //y=4.795 //x2=70.03 //y2=4.87
r552 (  101 102 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=69.955 //y=4.795 //x2=69.665 //y2=4.795
r553 (  100 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.595 //y=1.25 //x2=69.635 //y2=1.405
r554 (  99 147 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.595 //y=0.905 //x2=69.635 //y2=0.75
r555 (  99 100 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=69.595 //y=0.905 //x2=69.595 //y2=1.25
r556 (  96 102 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=69.59 //y=4.87 //x2=69.665 //y2=4.795
r557 (  95 146 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.215 //y=1.25 //x2=17.175 //y2=1.405
r558 (  94 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.215 //y=0.905 //x2=17.175 //y2=0.75
r559 (  94 95 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.215 //y=0.905 //x2=17.215 //y2=1.25
r560 (  89 144 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.84 //y=1.405 //x2=16.725 //y2=1.405
r561 (  88 146 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.06 //y=1.405 //x2=17.175 //y2=1.405
r562 (  87 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.84 //y=0.75 //x2=16.725 //y2=0.75
r563 (  86 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.06 //y=0.75 //x2=17.175 //y2=0.75
r564 (  86 87 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=17.06 //y=0.75 //x2=16.84 //y2=0.75
r565 (  85 141 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=16.815 //y=4.79 //x2=16.68 //y2=4.79
r566 (  84 91 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=17.055 //y=4.79 //x2=17.13 //y2=4.865
r567 (  84 85 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=17.055 //y=4.79 //x2=16.815 //y2=4.79
r568 (  79 144 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.685 //y=1.56 //x2=16.725 //y2=1.405
r569 (  79 136 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=16.685 //y=1.56 //x2=16.685 //y2=1.915
r570 (  78 144 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.685 //y=1.25 //x2=16.725 //y2=1.405
r571 (  77 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.685 //y=0.905 //x2=16.725 //y2=0.75
r572 (  77 78 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.685 //y=0.905 //x2=16.685 //y2=1.25
r573 (  76 131 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=72.49 //y=6.025 //x2=72.49 //y2=4.87
r574 (  75 119 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=72.05 //y=6.025 //x2=72.05 //y2=4.87
r575 (  74 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=70.03 //y=6.025 //x2=70.03 //y2=4.87
r576 (  73 96 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=69.59 //y=6.025 //x2=69.59 //y2=4.87
r577 (  72 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.13 //y=6.02 //x2=17.13 //y2=4.865
r578 (  71 142 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.69 //y=6.02 //x2=16.69 //y2=4.865
r579 (  70 124 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=72.22 //y=1.365 //x2=72.33 //y2=1.365
r580 (  70 125 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=72.22 //y=1.365 //x2=72.11 //y2=1.365
r581 (  69 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=69.86 //y=1.405 //x2=69.97 //y2=1.405
r582 (  69 106 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=69.86 //y=1.405 //x2=69.75 //y2=1.405
r583 (  68 88 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=16.95 //y=1.405 //x2=17.06 //y2=1.405
r584 (  68 89 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=16.95 //y=1.405 //x2=16.84 //y2=1.405
r585 (  66 139 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.68 //y=4.7 //x2=16.68 //y2=4.7
r586 (  63 158 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=71.78 //y=4.705 //x2=71.78 //y2=4.705
r587 (  59 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=71.78 //y=2.08 //x2=71.78 //y2=2.08
r588 (  59 63 ) resistor r=179.679 //w=0.187 //l=2.625 //layer=li \
 //thickness=0.1 //x=71.78 //y=2.08 //x2=71.78 //y2=4.705
r589 (  56 154 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=70.3 //y=4.705 //x2=70.3 //y2=4.705
r590 (  54 56 ) resistor r=119.444 //w=0.187 //l=1.745 //layer=li \
 //thickness=0.1 //x=70.3 //y=2.96 //x2=70.3 //y2=4.705
r591 (  50 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=70.3 //y=2.08 //x2=70.3 //y2=2.08
r592 (  50 54 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=70.3 //y=2.08 //x2=70.3 //y2=2.96
r593 (  46 48 ) resistor r=147.508 //w=0.187 //l=2.155 //layer=li \
 //thickness=0.1 //x=20.72 //y=5.115 //x2=20.72 //y2=2.96
r594 (  45 48 ) resistor r=83.508 //w=0.187 //l=1.22 //layer=li \
 //thickness=0.1 //x=20.72 //y=1.74 //x2=20.72 //y2=2.96
r595 (  43 45 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.635 //y=1.655 //x2=20.72 //y2=1.74
r596 (  43 44 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=20.635 //y=1.655 //x2=20.365 //y2=1.655
r597 (  42 67 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.325 //y=5.2 //x2=20.24 //y2=5.2
r598 (  41 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.635 //y=5.2 //x2=20.72 //y2=5.115
r599 (  41 42 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=20.635 //y=5.2 //x2=20.325 //y2=5.2
r600 (  37 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.28 //y=1.57 //x2=20.365 //y2=1.655
r601 (  37 163 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=20.28 //y=1.57 //x2=20.28 //y2=1
r602 (  31 67 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.24 //y=5.285 //x2=20.24 //y2=5.2
r603 (  31 166 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=20.24 //y=5.285 //x2=20.24 //y2=5.725
r604 (  29 67 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.155 //y=5.2 //x2=20.24 //y2=5.2
r605 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=20.155 //y=5.2 //x2=19.445 //y2=5.2
r606 (  23 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=19.36 //y=5.285 //x2=19.445 //y2=5.2
r607 (  23 165 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=19.36 //y=5.285 //x2=19.36 //y2=5.725
r608 (  19 135 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.65 //y=2.08 //x2=16.65 //y2=2.08
r609 (  19 22 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=16.65 //y=2.08 //x2=16.65 //y2=2.96
r610 (  17 66 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=16.65 //y=4.535 //x2=16.665 //y2=4.7
r611 (  17 22 ) resistor r=107.807 //w=0.187 //l=1.575 //layer=li \
 //thickness=0.1 //x=16.65 //y=4.535 //x2=16.65 //y2=2.96
r612 (  16 59 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=71.78 //y=2.08 //x2=71.78 //y2=2.08
r613 (  14 54 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=70.3 //y=2.96 //x2=70.3 //y2=2.96
r614 (  12 50 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=70.3 //y=2.08 //x2=70.3 //y2=2.08
r615 (  10 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=20.72 //y=2.96 //x2=20.72 //y2=2.96
r616 (  8 22 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=16.65 //y=2.96 //x2=16.65 //y2=2.96
r617 (  6 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=70.415 //y=2.08 //x2=70.3 //y2=2.08
r618 (  5 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=71.665 //y=2.08 //x2=71.78 //y2=2.08
r619 (  5 6 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=71.665 //y=2.08 //x2=70.415 //y2=2.08
r620 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.835 //y=2.96 //x2=20.72 //y2=2.96
r621 (  3 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=70.185 //y=2.96 //x2=70.3 //y2=2.96
r622 (  3 4 ) resistor r=47.0897 //w=0.131 //l=49.35 //layer=m1 \
 //thickness=0.36 //x=70.185 //y=2.96 //x2=20.835 //y2=2.96
r623 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.765 //y=2.96 //x2=16.65 //y2=2.96
r624 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=2.96 //x2=20.72 //y2=2.96
r625 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=2.96 //x2=16.765 //y2=2.96
ends PM_TMRDFFQNX1\%noxref_23

subckt PM_TMRDFFQNX1\%noxref_24 ( 1 2 13 14 15 21 27 28 35 46 47 48 49 50 )
c89 ( 50 0 ) capacitor c=0.0308836f //x=73.445 //y=5.025
c90 ( 49 0 ) capacitor c=0.0173945f //x=72.565 //y=5.025
c91 ( 47 0 ) capacitor c=0.0169278f //x=69.665 //y=5.025
c92 ( 46 0 ) capacitor c=0.0166762f //x=68.785 //y=5.025
c93 ( 45 0 ) capacitor c=0.00115294f //x=72.71 //y=6.91
c94 ( 35 0 ) capacitor c=0.0132983f //x=73.505 //y=6.91
c95 ( 28 0 ) capacitor c=0.00388794f //x=71.915 //y=6.91
c96 ( 27 0 ) capacitor c=0.00985708f //x=72.625 //y=6.91
c97 ( 21 0 ) capacitor c=0.0442221f //x=71.83 //y=5.21
c98 ( 15 0 ) capacitor c=0.0105083f //x=69.81 //y=5.295
c99 ( 14 0 ) capacitor c=0.00227812f //x=69.015 //y=5.21
c100 ( 13 0 ) capacitor c=0.0174384f //x=69.725 //y=5.21
c101 ( 2 0 ) capacitor c=0.00682032f //x=69.925 //y=5.21
c102 ( 1 0 ) capacitor c=0.0574911f //x=71.715 //y=5.21
r103 (  37 50 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.59 //y=6.825 //x2=73.59 //y2=6.74
r104 (  36 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.795 //y=6.91 //x2=72.71 //y2=6.91
r105 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=73.505 //y=6.91 //x2=73.59 //y2=6.825
r106 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=73.505 //y=6.91 //x2=72.795 //y2=6.91
r107 (  29 45 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.71 //y=6.825 //x2=72.71 //y2=6.91
r108 (  29 49 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.71 //y=6.825 //x2=72.71 //y2=6.74
r109 (  27 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.625 //y=6.91 //x2=72.71 //y2=6.91
r110 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=72.625 //y=6.91 //x2=71.915 //y2=6.91
r111 (  21 48 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=71.83 //y=5.21 //x2=71.83 //y2=6.06
r112 (  19 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=71.83 //y=6.825 //x2=71.915 //y2=6.91
r113 (  19 48 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.83 //y=6.825 //x2=71.83 //y2=6.74
r114 (  15 44 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=69.81 //y=5.295 //x2=69.81 //y2=5.17
r115 (  15 47 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=69.81 //y=5.295 //x2=69.81 //y2=6.06
r116 (  13 44 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=69.725 //y=5.21 //x2=69.81 //y2=5.17
r117 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=69.725 //y=5.21 //x2=69.015 //y2=5.21
r118 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=68.93 //y=5.295 //x2=69.015 //y2=5.21
r119 (  7 46 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=68.93 //y=5.295 //x2=68.93 //y2=5.72
r120 (  6 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=71.83 //y=5.21 //x2=71.83 //y2=5.21
r121 (  4 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=69.81 //y=5.21 //x2=69.81 //y2=5.21
r122 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=69.925 //y=5.21 //x2=69.81 //y2=5.21
r123 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=71.715 //y=5.21 //x2=71.83 //y2=5.21
r124 (  1 2 ) resistor r=1.70802 //w=0.131 //l=1.79 //layer=m1 \
 //thickness=0.36 //x=71.715 //y=5.21 //x2=69.925 //y2=5.21
ends PM_TMRDFFQNX1\%noxref_24

subckt PM_TMRDFFQNX1\%QN ( 1 2 3 4 11 12 13 14 15 16 17 18 31 32 45 47 48 63 \
 64 65 66 70 71 )
c169 ( 71 0 ) capacitor c=0.0167617f //x=73.005 //y=5.025
c170 ( 70 0 ) capacitor c=0.0164812f //x=72.125 //y=5.025
c171 ( 66 0 ) capacitor c=0.0108176f //x=73 //y=0.905
c172 ( 65 0 ) capacitor c=0.0131637f //x=69.67 //y=0.905
c173 ( 64 0 ) capacitor c=0.0131367f //x=66.34 //y=0.905
c174 ( 63 0 ) capacitor c=0.00421476f //x=73.15 //y=5.21
c175 ( 48 0 ) capacitor c=0.00775877f //x=73.275 //y=1.645
c176 ( 47 0 ) capacitor c=0.0165978f //x=73.545 //y=1.645
c177 ( 45 0 ) capacitor c=0.0160142f //x=73.545 //y=5.21
c178 ( 32 0 ) capacitor c=0.0029383f //x=72.355 //y=5.21
c179 ( 31 0 ) capacitor c=0.0155464f //x=73.065 //y=5.21
c180 ( 11 0 ) capacitor c=0.133166f //x=73.63 //y=2.22
c181 ( 4 0 ) capacitor c=0.00511584f //x=69.975 //y=1.18
c182 ( 3 0 ) capacitor c=0.0702096f //x=73.075 //y=1.18
c183 ( 2 0 ) capacitor c=0.0150174f //x=66.645 //y=1.18
c184 ( 1 0 ) capacitor c=0.0604206f //x=69.745 //y=1.18
r185 (  62 64 ) resistor r=13.3953 //w=0.172 //l=0.18 //layer=li \
 //thickness=0.1 //x=66.527 //y=1.18 //x2=66.527 //y2=1
r186 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=73.545 //y=1.645 //x2=73.63 //y2=1.73
r187 (  47 48 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=73.545 //y=1.645 //x2=73.275 //y2=1.645
r188 (  46 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.235 //y=5.21 //x2=73.15 //y2=5.21
r189 (  45 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=73.545 //y=5.21 //x2=73.63 //y2=5.125
r190 (  45 46 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=73.545 //y=5.21 //x2=73.235 //y2=5.21
r191 (  44 66 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=73.19 //y=1.18 //x2=73.19 //y2=1
r192 (  39 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=73.19 //y=1.56 //x2=73.275 //y2=1.645
r193 (  39 44 ) resistor r=26.0107 //w=0.187 //l=0.38 //layer=li \
 //thickness=0.1 //x=73.19 //y=1.56 //x2=73.19 //y2=1.18
r194 (  33 63 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.15 //y=5.295 //x2=73.15 //y2=5.21
r195 (  33 71 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=73.15 //y=5.295 //x2=73.15 //y2=5.72
r196 (  31 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.065 //y=5.21 //x2=73.15 //y2=5.21
r197 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=73.065 //y=5.21 //x2=72.355 //y2=5.21
r198 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=72.27 //y=5.295 //x2=72.355 //y2=5.21
r199 (  25 70 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=72.27 //y=5.295 //x2=72.27 //y2=5.72
r200 (  23 65 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=69.86 //y=1.18 //x2=69.86 //y2=1
r201 (  18 50 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=73.63 //y=4.81 //x2=73.63 //y2=5.125
r202 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=73.63 //y=4.44 //x2=73.63 //y2=4.81
r203 (  16 17 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=73.63 //y=4.07 //x2=73.63 //y2=4.44
r204 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=73.63 //y=3.7 //x2=73.63 //y2=4.07
r205 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=73.63 //y=3.33 //x2=73.63 //y2=3.7
r206 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=73.63 //y=2.96 //x2=73.63 //y2=3.33
r207 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=73.63 //y=2.59 //x2=73.63 //y2=2.96
r208 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=73.63 //y=2.22 //x2=73.63 //y2=2.59
r209 (  11 49 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=73.63 //y=2.22 //x2=73.63 //y2=1.73
r210 (  10 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=73.19 //y=1.18 //x2=73.19 //y2=1.18
r211 (  8 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=69.86 //y=1.18 //x2=69.86 //y2=1.18
r212 (  6 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=66.53 //y=1.18 //x2=66.53 //y2=1.18
r213 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=69.975 //y=1.18 //x2=69.86 //y2=1.18
r214 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=73.075 //y=1.18 //x2=73.19 //y2=1.18
r215 (  3 4 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=73.075 //y=1.18 //x2=69.975 //y2=1.18
r216 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=66.645 //y=1.18 //x2=66.53 //y2=1.18
r217 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=69.745 //y=1.18 //x2=69.86 //y2=1.18
r218 (  1 2 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=69.745 //y=1.18 //x2=66.645 //y2=1.18
ends PM_TMRDFFQNX1\%QN

subckt PM_TMRDFFQNX1\%noxref_26 ( 1 5 9 13 17 35 )
c47 ( 35 0 ) capacitor c=0.0703709f //x=0.455 //y=0.375
c48 ( 17 0 ) capacitor c=0.0221229f //x=2.445 //y=1.59
c49 ( 13 0 ) capacitor c=0.0156939f //x=2.445 //y=0.54
c50 ( 9 0 ) capacitor c=0.00678203f //x=1.56 //y=0.625
c51 ( 5 0 ) capacitor c=0.0206412f //x=1.475 //y=1.59
c52 ( 1 0 ) capacitor c=0.0109947f //x=0.59 //y=1.505
r53 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=1.59 //x2=1.56 //y2=1.63
r54 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=1.59 //x2=2.045 //y2=1.59
r55 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=1.59 //x2=2.53 //y2=1.59
r56 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=1.59 //x2=2.045 //y2=1.59
r57 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=0.54 //x2=1.56 //y2=0.5
r58 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=0.54 //x2=2.045 //y2=0.54
r59 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=0.54 //x2=2.53 //y2=0.54
r60 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=0.54 //x2=2.045 //y2=0.54
r61 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=1.63
r62 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=0.89
r63 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.5
r64 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.89
r65 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.675 //y=1.59 //x2=0.59 //y2=1.63
r66 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.675 //y=1.59 //x2=1.075 //y2=1.59
r67 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.475 //y=1.59 //x2=1.56 //y2=1.63
r68 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.475 //y=1.59 //x2=1.075 //y2=1.59
r69 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.59 //y=1.505 //x2=0.59 //y2=1.63
r70 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.59 //y=1.505 //x2=0.59 //y2=0.89
ends PM_TMRDFFQNX1\%noxref_26

subckt PM_TMRDFFQNX1\%noxref_27 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.043074f //x=2.965 //y=0.375
c54 ( 28 0 ) capacitor c=0.00465142f //x=1.86 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=3.1 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=4.07 //y=0.625
c57 ( 11 0 ) capacitor c=0.0149771f //x=3.985 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=3.1 //y=0.625
c59 ( 1 0 ) capacitor c=0.0251532f //x=3.015 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.185 //y=0.54 //x2=3.1 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.185 //y=0.54 //x2=3.585 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.985 //y=0.54 //x2=4.07 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.985 //y=0.54 //x2=3.585 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.135 //y=0.995 //x2=2.05 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=3.1 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=2.135 //y2=0.995
ends PM_TMRDFFQNX1\%noxref_27

subckt PM_TMRDFFQNX1\%noxref_28 ( 1 5 9 10 13 17 29 )
c54 ( 29 0 ) capacitor c=0.0634189f //x=5.37 //y=0.365
c55 ( 17 0 ) capacitor c=0.00722223f //x=7.445 //y=0.615
c56 ( 13 0 ) capacitor c=0.0146588f //x=7.36 //y=0.53
c57 ( 10 0 ) capacitor c=0.00656209f //x=6.475 //y=1.495
c58 ( 9 0 ) capacitor c=0.006761f //x=6.475 //y=0.615
c59 ( 5 0 ) capacitor c=0.0196287f //x=6.39 //y=1.58
c60 ( 1 0 ) capacitor c=0.00828748f //x=5.505 //y=1.495
r61 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=7.445 //y=0.615 //x2=7.445 //y2=0.49
r62 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=7.445 //y=0.615 //x2=7.445 //y2=0.88
r63 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.56 //y=0.53 //x2=6.475 //y2=0.49
r64 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.56 //y=0.53 //x2=6.96 //y2=0.53
r65 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.36 //y=0.53 //x2=7.445 //y2=0.49
r66 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.36 //y=0.53 //x2=6.96 //y2=0.53
r67 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=6.475 //y=1.495 //x2=6.475 //y2=1.62
r68 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.475 //y=1.495 //x2=6.475 //y2=0.88
r69 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.475 //y=0.615 //x2=6.475 //y2=0.49
r70 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.475 //y=0.615 //x2=6.475 //y2=0.88
r71 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.59 //y=1.58 //x2=5.505 //y2=1.62
r72 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.59 //y=1.58 //x2=5.99 //y2=1.58
r73 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.39 //y=1.58 //x2=6.475 //y2=1.62
r74 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.39 //y=1.58 //x2=5.99 //y2=1.58
r75 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=5.505 //y=1.495 //x2=5.505 //y2=1.62
r76 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=5.505 //y=1.495 //x2=5.505 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_28

subckt PM_TMRDFFQNX1\%noxref_29 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0634191f //x=8.7 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=10.775 //y=0.615
c54 ( 13 0 ) capacitor c=0.014662f //x=10.69 //y=0.53
c55 ( 10 0 ) capacitor c=0.00610102f //x=9.805 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=9.805 //y=0.615
c57 ( 5 0 ) capacitor c=0.0181202f //x=9.72 //y=1.58
c58 ( 1 0 ) capacitor c=0.00765941f //x=8.835 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=10.775 //y=0.615 //x2=10.775 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=10.775 //y=0.615 //x2=10.775 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.89 //y=0.53 //x2=9.805 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.89 //y=0.53 //x2=10.29 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.69 //y=0.53 //x2=10.775 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.69 //y=0.53 //x2=10.29 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=9.805 //y=1.495 //x2=9.805 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=9.805 //y=1.495 //x2=9.805 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=9.805 //y=0.615 //x2=9.805 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=9.805 //y=0.615 //x2=9.805 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.92 //y=1.58 //x2=8.835 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.92 //y=1.58 //x2=9.32 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.72 //y=1.58 //x2=9.805 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.72 //y=1.58 //x2=9.32 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=8.835 //y=1.495 //x2=8.835 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=8.835 //y=1.495 //x2=8.835 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_29

subckt PM_TMRDFFQNX1\%noxref_30 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0634191f //x=12.03 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=14.105 //y=0.615
c54 ( 13 0 ) capacitor c=0.014662f //x=14.02 //y=0.53
c55 ( 10 0 ) capacitor c=0.00610102f //x=13.135 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=13.135 //y=0.615
c57 ( 5 0 ) capacitor c=0.0181202f //x=13.05 //y=1.58
c58 ( 1 0 ) capacitor c=0.00765941f //x=12.165 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=14.105 //y=0.615 //x2=14.105 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=14.105 //y=0.615 //x2=14.105 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.22 //y=0.53 //x2=13.135 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.22 //y=0.53 //x2=13.62 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.02 //y=0.53 //x2=14.105 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.02 //y=0.53 //x2=13.62 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=13.135 //y=1.495 //x2=13.135 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=13.135 //y=1.495 //x2=13.135 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=13.135 //y=0.615 //x2=13.135 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=13.135 //y=0.615 //x2=13.135 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.25 //y=1.58 //x2=12.165 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.25 //y=1.58 //x2=12.65 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.05 //y=1.58 //x2=13.135 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.05 //y=1.58 //x2=12.65 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=12.165 //y=1.495 //x2=12.165 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=12.165 //y=1.495 //x2=12.165 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_30

subckt PM_TMRDFFQNX1\%noxref_31 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0634191f //x=15.36 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=17.435 //y=0.615
c54 ( 13 0 ) capacitor c=0.014662f //x=17.35 //y=0.53
c55 ( 10 0 ) capacitor c=0.00610102f //x=16.465 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=16.465 //y=0.615
c57 ( 5 0 ) capacitor c=0.0181202f //x=16.38 //y=1.58
c58 ( 1 0 ) capacitor c=0.00765941f //x=15.495 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=17.435 //y=0.615 //x2=17.435 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=17.435 //y=0.615 //x2=17.435 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.55 //y=0.53 //x2=16.465 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.55 //y=0.53 //x2=16.95 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.35 //y=0.53 //x2=17.435 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.35 //y=0.53 //x2=16.95 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=16.465 //y=1.495 //x2=16.465 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=16.465 //y=1.495 //x2=16.465 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=16.465 //y=0.615 //x2=16.465 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=16.465 //y=0.615 //x2=16.465 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.58 //y=1.58 //x2=15.495 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.58 //y=1.58 //x2=15.98 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.38 //y=1.58 //x2=16.465 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.38 //y=1.58 //x2=15.98 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=15.495 //y=1.495 //x2=15.495 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=15.495 //y=1.495 //x2=15.495 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_31

subckt PM_TMRDFFQNX1\%noxref_32 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0634191f //x=18.69 //y=0.365
c53 ( 17 0 ) capacitor c=0.0072343f //x=20.765 //y=0.615
c54 ( 13 0 ) capacitor c=0.014662f //x=20.68 //y=0.53
c55 ( 10 0 ) capacitor c=0.00610102f //x=19.795 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=19.795 //y=0.615
c57 ( 5 0 ) capacitor c=0.0181202f //x=19.71 //y=1.58
c58 ( 1 0 ) capacitor c=0.00765941f //x=18.825 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=20.765 //y=0.615 //x2=20.765 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=20.765 //y=0.615 //x2=20.765 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.88 //y=0.53 //x2=19.795 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.88 //y=0.53 //x2=20.28 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.68 //y=0.53 //x2=20.765 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.68 //y=0.53 //x2=20.28 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=19.795 //y=1.495 //x2=19.795 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=19.795 //y=1.495 //x2=19.795 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=19.795 //y=0.615 //x2=19.795 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=19.795 //y=0.615 //x2=19.795 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.91 //y=1.58 //x2=18.825 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.91 //y=1.58 //x2=19.31 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.71 //y=1.58 //x2=19.795 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.71 //y=1.58 //x2=19.31 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=18.825 //y=1.495 //x2=18.825 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=18.825 //y=1.495 //x2=18.825 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_32

subckt PM_TMRDFFQNX1\%noxref_33 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0679963f //x=21.915 //y=0.375
c51 ( 17 0 ) capacitor c=0.018806f //x=23.905 //y=1.59
c52 ( 13 0 ) capacitor c=0.0155484f //x=23.905 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=23.02 //y=0.625
c54 ( 5 0 ) capacitor c=0.0170872f //x=22.935 //y=1.59
c55 ( 1 0 ) capacitor c=0.00729042f //x=22.05 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.105 //y=1.59 //x2=23.02 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.105 //y=1.59 //x2=23.505 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.905 //y=1.59 //x2=23.99 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.905 //y=1.59 //x2=23.505 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.105 //y=0.54 //x2=23.02 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.105 //y=0.54 //x2=23.505 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.905 //y=0.54 //x2=23.99 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.905 //y=0.54 //x2=23.505 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=23.02 //y=1.505 //x2=23.02 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=23.02 //y=1.505 //x2=23.02 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=23.02 //y=0.625 //x2=23.02 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=23.02 //y=0.625 //x2=23.02 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=22.135 //y=1.59 //x2=22.05 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.135 //y=1.59 //x2=22.535 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=22.935 //y=1.59 //x2=23.02 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.935 //y=1.59 //x2=22.535 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=22.05 //y=1.505 //x2=22.05 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=22.05 //y=1.505 //x2=22.05 //y2=0.89
ends PM_TMRDFFQNX1\%noxref_33

subckt PM_TMRDFFQNX1\%noxref_34 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0418028f //x=24.425 //y=0.375
c54 ( 28 0 ) capacitor c=0.00460056f //x=23.32 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=24.56 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=25.53 //y=0.625
c57 ( 11 0 ) capacitor c=0.0145763f //x=25.445 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=24.56 //y=0.625
c59 ( 1 0 ) capacitor c=0.022715f //x=24.475 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=25.53 //y=0.625 //x2=25.53 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=25.53 //y=0.625 //x2=25.53 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=24.645 //y=0.54 //x2=24.56 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=24.645 //y=0.54 //x2=25.045 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.445 //y=0.54 //x2=25.53 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.445 //y=0.54 //x2=25.045 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=24.56 //y=1.08 //x2=24.56 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=24.56 //y=1.08 //x2=24.56 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=24.56 //y=0.91 //x2=24.56 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=24.56 //y=0.91 //x2=24.56 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=24.56 //y=0.625 //x2=24.56 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=24.56 //y=0.625 //x2=24.56 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.595 //y=0.995 //x2=23.51 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=24.475 //y=0.995 //x2=24.56 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=24.475 //y=0.995 //x2=23.595 //y2=0.995
ends PM_TMRDFFQNX1\%noxref_34

subckt PM_TMRDFFQNX1\%noxref_35 ( 1 5 9 10 13 17 29 )
c54 ( 29 0 ) capacitor c=0.0634189f //x=26.83 //y=0.365
c55 ( 17 0 ) capacitor c=0.00722223f //x=28.905 //y=0.615
c56 ( 13 0 ) capacitor c=0.0146588f //x=28.82 //y=0.53
c57 ( 10 0 ) capacitor c=0.00610027f //x=27.935 //y=1.495
c58 ( 9 0 ) capacitor c=0.006761f //x=27.935 //y=0.615
c59 ( 5 0 ) capacitor c=0.0181202f //x=27.85 //y=1.58
c60 ( 1 0 ) capacitor c=0.00765941f //x=26.965 //y=1.495
r61 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=28.905 //y=0.615 //x2=28.905 //y2=0.49
r62 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=28.905 //y=0.615 //x2=28.905 //y2=0.88
r63 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=28.02 //y=0.53 //x2=27.935 //y2=0.49
r64 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=28.02 //y=0.53 //x2=28.42 //y2=0.53
r65 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=28.82 //y=0.53 //x2=28.905 //y2=0.49
r66 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=28.82 //y=0.53 //x2=28.42 //y2=0.53
r67 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=27.935 //y=1.495 //x2=27.935 //y2=1.62
r68 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=27.935 //y=1.495 //x2=27.935 //y2=0.88
r69 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=27.935 //y=0.615 //x2=27.935 //y2=0.49
r70 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=27.935 //y=0.615 //x2=27.935 //y2=0.88
r71 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=27.05 //y=1.58 //x2=26.965 //y2=1.62
r72 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=27.05 //y=1.58 //x2=27.45 //y2=1.58
r73 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=27.85 //y=1.58 //x2=27.935 //y2=1.62
r74 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=27.85 //y=1.58 //x2=27.45 //y2=1.58
r75 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=26.965 //y=1.495 //x2=26.965 //y2=1.62
r76 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=26.965 //y=1.495 //x2=26.965 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_35

subckt PM_TMRDFFQNX1\%noxref_36 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0634191f //x=30.16 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=32.235 //y=0.615
c54 ( 13 0 ) capacitor c=0.014662f //x=32.15 //y=0.53
c55 ( 10 0 ) capacitor c=0.00610102f //x=31.265 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=31.265 //y=0.615
c57 ( 5 0 ) capacitor c=0.0181202f //x=31.18 //y=1.58
c58 ( 1 0 ) capacitor c=0.00765941f //x=30.295 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=32.235 //y=0.615 //x2=32.235 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=32.235 //y=0.615 //x2=32.235 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=31.35 //y=0.53 //x2=31.265 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=31.35 //y=0.53 //x2=31.75 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=32.15 //y=0.53 //x2=32.235 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=32.15 //y=0.53 //x2=31.75 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=31.265 //y=1.495 //x2=31.265 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=31.265 //y=1.495 //x2=31.265 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=31.265 //y=0.615 //x2=31.265 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=31.265 //y=0.615 //x2=31.265 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=30.38 //y=1.58 //x2=30.295 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.38 //y=1.58 //x2=30.78 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=31.18 //y=1.58 //x2=31.265 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=31.18 //y=1.58 //x2=30.78 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=30.295 //y=1.495 //x2=30.295 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=30.295 //y=1.495 //x2=30.295 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_36

subckt PM_TMRDFFQNX1\%noxref_37 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0634191f //x=33.49 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=35.565 //y=0.615
c54 ( 13 0 ) capacitor c=0.014662f //x=35.48 //y=0.53
c55 ( 10 0 ) capacitor c=0.00610102f //x=34.595 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=34.595 //y=0.615
c57 ( 5 0 ) capacitor c=0.0181202f //x=34.51 //y=1.58
c58 ( 1 0 ) capacitor c=0.00765941f //x=33.625 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=35.565 //y=0.615 //x2=35.565 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=35.565 //y=0.615 //x2=35.565 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=34.68 //y=0.53 //x2=34.595 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=34.68 //y=0.53 //x2=35.08 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=35.48 //y=0.53 //x2=35.565 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.48 //y=0.53 //x2=35.08 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=34.595 //y=1.495 //x2=34.595 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=34.595 //y=1.495 //x2=34.595 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=34.595 //y=0.615 //x2=34.595 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=34.595 //y=0.615 //x2=34.595 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=33.71 //y=1.58 //x2=33.625 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=33.71 //y=1.58 //x2=34.11 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=34.51 //y=1.58 //x2=34.595 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=34.51 //y=1.58 //x2=34.11 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=33.625 //y=1.495 //x2=33.625 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=33.625 //y=1.495 //x2=33.625 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_37

subckt PM_TMRDFFQNX1\%noxref_38 ( 1 5 9 10 13 17 29 )
c54 ( 29 0 ) capacitor c=0.0632684f //x=36.82 //y=0.365
c55 ( 17 0 ) capacitor c=0.00722223f //x=38.895 //y=0.615
c56 ( 13 0 ) capacitor c=0.0145042f //x=38.81 //y=0.53
c57 ( 10 0 ) capacitor c=0.00605993f //x=37.925 //y=1.495
c58 ( 9 0 ) capacitor c=0.006761f //x=37.925 //y=0.615
c59 ( 5 0 ) capacitor c=0.0181202f //x=37.84 //y=1.58
c60 ( 1 0 ) capacitor c=0.00765941f //x=36.955 //y=1.495
r61 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=38.895 //y=0.615 //x2=38.895 //y2=0.49
r62 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=38.895 //y=0.615 //x2=38.895 //y2=0.88
r63 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=38.01 //y=0.53 //x2=37.925 //y2=0.49
r64 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=38.01 //y=0.53 //x2=38.41 //y2=0.53
r65 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=38.81 //y=0.53 //x2=38.895 //y2=0.49
r66 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=38.81 //y=0.53 //x2=38.41 //y2=0.53
r67 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=37.925 //y=1.495 //x2=37.925 //y2=1.62
r68 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=37.925 //y=1.495 //x2=37.925 //y2=0.88
r69 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=37.925 //y=0.615 //x2=37.925 //y2=0.49
r70 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=37.925 //y=0.615 //x2=37.925 //y2=0.88
r71 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=37.04 //y=1.58 //x2=36.955 //y2=1.62
r72 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=37.04 //y=1.58 //x2=37.44 //y2=1.58
r73 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=37.84 //y=1.58 //x2=37.925 //y2=1.62
r74 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=37.84 //y=1.58 //x2=37.44 //y2=1.58
r75 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=36.955 //y=1.495 //x2=36.955 //y2=1.62
r76 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=36.955 //y=1.495 //x2=36.955 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_38

subckt PM_TMRDFFQNX1\%noxref_39 ( 1 5 9 10 13 17 29 )
c54 ( 29 0 ) capacitor c=0.0632577f //x=40.15 //y=0.365
c55 ( 17 0 ) capacitor c=0.0072343f //x=42.225 //y=0.615
c56 ( 13 0 ) capacitor c=0.0145076f //x=42.14 //y=0.53
c57 ( 10 0 ) capacitor c=0.00582081f //x=41.255 //y=1.495
c58 ( 9 0 ) capacitor c=0.006761f //x=41.255 //y=0.615
c59 ( 5 0 ) capacitor c=0.0173046f //x=41.17 //y=1.58
c60 ( 1 0 ) capacitor c=0.00733328f //x=40.285 //y=1.495
r61 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=42.225 //y=0.615 //x2=42.225 //y2=0.49
r62 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=42.225 //y=0.615 //x2=42.225 //y2=0.88
r63 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=41.34 //y=0.53 //x2=41.255 //y2=0.49
r64 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=41.34 //y=0.53 //x2=41.74 //y2=0.53
r65 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=42.14 //y=0.53 //x2=42.225 //y2=0.49
r66 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=42.14 //y=0.53 //x2=41.74 //y2=0.53
r67 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=41.255 //y=1.495 //x2=41.255 //y2=1.62
r68 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=41.255 //y=1.495 //x2=41.255 //y2=0.88
r69 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=41.255 //y=0.615 //x2=41.255 //y2=0.49
r70 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=41.255 //y=0.615 //x2=41.255 //y2=0.88
r71 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=40.37 //y=1.58 //x2=40.285 //y2=1.62
r72 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=40.37 //y=1.58 //x2=40.77 //y2=1.58
r73 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=41.17 //y=1.58 //x2=41.255 //y2=1.62
r74 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=41.17 //y=1.58 //x2=40.77 //y2=1.58
r75 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=40.285 //y=1.495 //x2=40.285 //y2=1.62
r76 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=40.285 //y=1.495 //x2=40.285 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_39

subckt PM_TMRDFFQNX1\%noxref_40 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0673029f //x=43.375 //y=0.375
c51 ( 17 0 ) capacitor c=0.0178317f //x=45.365 //y=1.59
c52 ( 13 0 ) capacitor c=0.0154936f //x=45.365 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=44.48 //y=0.625
c54 ( 5 0 ) capacitor c=0.0164013f //x=44.395 //y=1.59
c55 ( 1 0 ) capacitor c=0.00696517f //x=43.51 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=44.565 //y=1.59 //x2=44.48 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=44.565 //y=1.59 //x2=44.965 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.365 //y=1.59 //x2=45.45 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.365 //y=1.59 //x2=44.965 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=44.565 //y=0.54 //x2=44.48 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=44.565 //y=0.54 //x2=44.965 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.365 //y=0.54 //x2=45.45 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.365 //y=0.54 //x2=44.965 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=44.48 //y=1.505 //x2=44.48 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=44.48 //y=1.505 //x2=44.48 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=44.48 //y=0.625 //x2=44.48 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=44.48 //y=0.625 //x2=44.48 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=43.595 //y=1.59 //x2=43.51 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=43.595 //y=1.59 //x2=43.995 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=44.395 //y=1.59 //x2=44.48 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=44.395 //y=1.59 //x2=43.995 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=43.51 //y=1.505 //x2=43.51 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=43.51 //y=1.505 //x2=43.51 //y2=0.89
ends PM_TMRDFFQNX1\%noxref_40

subckt PM_TMRDFFQNX1\%noxref_41 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0413887f //x=45.885 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=44.78 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=46.02 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=46.99 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144274f //x=46.905 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=46.02 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=45.935 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=46.99 //y=0.625 //x2=46.99 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=46.99 //y=0.625 //x2=46.99 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=46.105 //y=0.54 //x2=46.02 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=46.105 //y=0.54 //x2=46.505 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=46.905 //y=0.54 //x2=46.99 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=46.905 //y=0.54 //x2=46.505 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=46.02 //y=1.08 //x2=46.02 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=46.02 //y=1.08 //x2=46.02 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=46.02 //y=0.91 //x2=46.02 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=46.02 //y=0.91 //x2=46.02 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=46.02 //y=0.625 //x2=46.02 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=46.02 //y=0.625 //x2=46.02 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.055 //y=0.995 //x2=44.97 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=45.935 //y=0.995 //x2=46.02 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=45.935 //y=0.995 //x2=45.055 //y2=0.995
ends PM_TMRDFFQNX1\%noxref_41

subckt PM_TMRDFFQNX1\%noxref_42 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0632682f //x=48.29 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=50.365 //y=0.615
c54 ( 13 0 ) capacitor c=0.0145084f //x=50.28 //y=0.53
c55 ( 10 0 ) capacitor c=0.00582081f //x=49.395 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=49.395 //y=0.615
c57 ( 5 0 ) capacitor c=0.0173046f //x=49.31 //y=1.58
c58 ( 1 0 ) capacitor c=0.00733328f //x=48.425 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=50.365 //y=0.615 //x2=50.365 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=50.365 //y=0.615 //x2=50.365 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=49.48 //y=0.53 //x2=49.395 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=49.48 //y=0.53 //x2=49.88 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=50.28 //y=0.53 //x2=50.365 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=50.28 //y=0.53 //x2=49.88 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=49.395 //y=1.495 //x2=49.395 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=49.395 //y=1.495 //x2=49.395 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=49.395 //y=0.615 //x2=49.395 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=49.395 //y=0.615 //x2=49.395 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=48.51 //y=1.58 //x2=48.425 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=48.51 //y=1.58 //x2=48.91 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=49.31 //y=1.58 //x2=49.395 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=49.31 //y=1.58 //x2=48.91 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=48.425 //y=1.495 //x2=48.425 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=48.425 //y=1.495 //x2=48.425 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_42

subckt PM_TMRDFFQNX1\%noxref_43 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0632684f //x=51.62 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=53.695 //y=0.615
c54 ( 13 0 ) capacitor c=0.0145084f //x=53.61 //y=0.53
c55 ( 10 0 ) capacitor c=0.00582081f //x=52.725 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=52.725 //y=0.615
c57 ( 5 0 ) capacitor c=0.0173046f //x=52.64 //y=1.58
c58 ( 1 0 ) capacitor c=0.00733328f //x=51.755 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=53.695 //y=0.615 //x2=53.695 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=53.695 //y=0.615 //x2=53.695 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=52.81 //y=0.53 //x2=52.725 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=52.81 //y=0.53 //x2=53.21 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=53.61 //y=0.53 //x2=53.695 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=53.61 //y=0.53 //x2=53.21 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=52.725 //y=1.495 //x2=52.725 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=52.725 //y=1.495 //x2=52.725 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=52.725 //y=0.615 //x2=52.725 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=52.725 //y=0.615 //x2=52.725 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=51.84 //y=1.58 //x2=51.755 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=51.84 //y=1.58 //x2=52.24 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=52.64 //y=1.58 //x2=52.725 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=52.64 //y=1.58 //x2=52.24 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=51.755 //y=1.495 //x2=51.755 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=51.755 //y=1.495 //x2=51.755 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_43

subckt PM_TMRDFFQNX1\%noxref_44 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0632684f //x=54.95 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=57.025 //y=0.615
c54 ( 13 0 ) capacitor c=0.0145084f //x=56.94 //y=0.53
c55 ( 10 0 ) capacitor c=0.00582081f //x=56.055 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=56.055 //y=0.615
c57 ( 5 0 ) capacitor c=0.0173046f //x=55.97 //y=1.58
c58 ( 1 0 ) capacitor c=0.00733328f //x=55.085 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=57.025 //y=0.615 //x2=57.025 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=57.025 //y=0.615 //x2=57.025 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=56.14 //y=0.53 //x2=56.055 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=56.14 //y=0.53 //x2=56.54 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=56.94 //y=0.53 //x2=57.025 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=56.94 //y=0.53 //x2=56.54 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=56.055 //y=1.495 //x2=56.055 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=56.055 //y=1.495 //x2=56.055 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=56.055 //y=0.615 //x2=56.055 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=56.055 //y=0.615 //x2=56.055 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=55.17 //y=1.58 //x2=55.085 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=55.17 //y=1.58 //x2=55.57 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=55.97 //y=1.58 //x2=56.055 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=55.97 //y=1.58 //x2=55.57 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=55.085 //y=1.495 //x2=55.085 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=55.085 //y=1.495 //x2=55.085 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_44

subckt PM_TMRDFFQNX1\%noxref_45 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0632684f //x=58.28 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=60.355 //y=0.615
c54 ( 13 0 ) capacitor c=0.0145084f //x=60.27 //y=0.53
c55 ( 10 0 ) capacitor c=0.00582081f //x=59.385 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=59.385 //y=0.615
c57 ( 5 0 ) capacitor c=0.0173046f //x=59.3 //y=1.58
c58 ( 1 0 ) capacitor c=0.00733328f //x=58.415 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=60.355 //y=0.615 //x2=60.355 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=60.355 //y=0.615 //x2=60.355 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=59.47 //y=0.53 //x2=59.385 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.47 //y=0.53 //x2=59.87 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=60.27 //y=0.53 //x2=60.355 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=60.27 //y=0.53 //x2=59.87 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=59.385 //y=1.495 //x2=59.385 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=59.385 //y=1.495 //x2=59.385 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=59.385 //y=0.615 //x2=59.385 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=59.385 //y=0.615 //x2=59.385 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=58.5 //y=1.58 //x2=58.415 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=58.5 //y=1.58 //x2=58.9 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=59.3 //y=1.58 //x2=59.385 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.3 //y=1.58 //x2=58.9 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=58.415 //y=1.495 //x2=58.415 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=58.415 //y=1.495 //x2=58.415 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_45

subckt PM_TMRDFFQNX1\%noxref_46 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0631409f //x=61.61 //y=0.365
c53 ( 17 0 ) capacitor c=0.00722223f //x=63.685 //y=0.615
c54 ( 13 0 ) capacitor c=0.0145084f //x=63.6 //y=0.53
c55 ( 10 0 ) capacitor c=0.00582081f //x=62.715 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=62.715 //y=0.615
c57 ( 5 0 ) capacitor c=0.0173046f //x=62.63 //y=1.58
c58 ( 1 0 ) capacitor c=0.00733328f //x=61.745 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=63.685 //y=0.615 //x2=63.685 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=63.685 //y=0.615 //x2=63.685 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=62.8 //y=0.53 //x2=62.715 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=62.8 //y=0.53 //x2=63.2 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=63.6 //y=0.53 //x2=63.685 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=63.6 //y=0.53 //x2=63.2 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=62.715 //y=1.495 //x2=62.715 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=62.715 //y=1.495 //x2=62.715 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=62.715 //y=0.615 //x2=62.715 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=62.715 //y=0.615 //x2=62.715 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=61.83 //y=1.58 //x2=61.745 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=61.83 //y=1.58 //x2=62.23 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=62.63 //y=1.58 //x2=62.715 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=62.63 //y=1.58 //x2=62.23 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=61.745 //y=1.495 //x2=61.745 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=61.745 //y=1.495 //x2=61.745 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_46

subckt PM_TMRDFFQNX1\%noxref_47 ( 1 5 9 10 13 17 29 )
c58 ( 29 0 ) capacitor c=0.0758145f //x=64.94 //y=0.365
c59 ( 17 0 ) capacitor c=0.0072249f //x=67.015 //y=0.615
c60 ( 13 0 ) capacitor c=0.0153113f //x=66.93 //y=0.53
c61 ( 10 0 ) capacitor c=0.00698223f //x=66.045 //y=1.495
c62 ( 9 0 ) capacitor c=0.006761f //x=66.045 //y=0.615
c63 ( 5 0 ) capacitor c=0.0191191f //x=65.96 //y=1.58
c64 ( 1 0 ) capacitor c=0.00483164f //x=65.075 //y=1.495
r65 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=67.015 //y=0.615 //x2=67.015 //y2=0.49
r66 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=67.015 //y=0.615 //x2=67.015 //y2=1.22
r67 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=66.13 //y=0.53 //x2=66.045 //y2=0.49
r68 (  14 29 ) resistor r=27.0374 //w=0.187 //l=0.395 //layer=li \
 //thickness=0.1 //x=66.13 //y=0.53 //x2=66.525 //y2=0.53
r69 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=66.93 //y=0.53 //x2=67.015 //y2=0.49
r70 (  13 29 ) resistor r=27.7219 //w=0.187 //l=0.405 //layer=li \
 //thickness=0.1 //x=66.93 //y=0.53 //x2=66.525 //y2=0.53
r71 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=66.045 //y=1.495 //x2=66.045 //y2=1.62
r72 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=66.045 //y=1.495 //x2=66.045 //y2=0.88
r73 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=66.045 //y=0.615 //x2=66.045 //y2=0.49
r74 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=66.045 //y=0.615 //x2=66.045 //y2=0.88
r75 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=65.16 //y=1.58 //x2=65.075 //y2=1.62
r76 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=65.16 //y=1.58 //x2=65.56 //y2=1.58
r77 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=65.96 //y=1.58 //x2=66.045 //y2=1.62
r78 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=65.96 //y=1.58 //x2=65.56 //y2=1.58
r79 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=65.075 //y=1.495 //x2=65.075 //y2=1.62
r80 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=65.075 //y=1.495 //x2=65.075 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_47

subckt PM_TMRDFFQNX1\%noxref_48 ( 1 5 9 10 13 17 29 )
c56 ( 29 0 ) capacitor c=0.0723103f //x=68.27 //y=0.365
c57 ( 17 0 ) capacitor c=0.0072249f //x=70.345 //y=0.615
c58 ( 13 0 ) capacitor c=0.0155051f //x=70.26 //y=0.53
c59 ( 10 0 ) capacitor c=0.00876912f //x=69.375 //y=1.495
c60 ( 9 0 ) capacitor c=0.006761f //x=69.375 //y=0.615
c61 ( 5 0 ) capacitor c=0.0182818f //x=69.29 //y=1.58
c62 ( 1 0 ) capacitor c=0.00857722f //x=68.405 //y=1.495
r63 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=70.345 //y=0.615 //x2=70.345 //y2=0.49
r64 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=70.345 //y=0.615 //x2=70.345 //y2=1.22
r65 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=69.46 //y=0.53 //x2=69.375 //y2=0.49
r66 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=69.46 //y=0.53 //x2=69.86 //y2=0.53
r67 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=70.26 //y=0.53 //x2=70.345 //y2=0.49
r68 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=70.26 //y=0.53 //x2=69.86 //y2=0.53
r69 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=69.375 //y=1.495 //x2=69.375 //y2=1.62
r70 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=69.375 //y=1.495 //x2=69.375 //y2=0.88
r71 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=69.375 //y=0.615 //x2=69.375 //y2=0.49
r72 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=69.375 //y=0.615 //x2=69.375 //y2=0.88
r73 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=68.49 //y=1.58 //x2=68.405 //y2=1.62
r74 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=68.49 //y=1.58 //x2=68.89 //y2=1.58
r75 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=69.29 //y=1.58 //x2=69.375 //y2=1.62
r76 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=69.29 //y=1.58 //x2=68.89 //y2=1.58
r77 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=68.405 //y=1.495 //x2=68.405 //y2=1.62
r78 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=68.405 //y=1.495 //x2=68.405 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_48

subckt PM_TMRDFFQNX1\%noxref_49 ( 1 5 9 10 13 17 29 )
c53 ( 29 0 ) capacitor c=0.0643725f //x=71.6 //y=0.365
c54 ( 17 0 ) capacitor c=0.00722228f //x=73.675 //y=0.615
c55 ( 13 0 ) capacitor c=0.0141607f //x=73.59 //y=0.53
c56 ( 10 0 ) capacitor c=0.00712138f //x=72.705 //y=1.495
c57 ( 9 0 ) capacitor c=0.006761f //x=72.705 //y=0.615
c58 ( 5 0 ) capacitor c=0.0233454f //x=72.62 //y=1.58
c59 ( 1 0 ) capacitor c=0.00481264f //x=71.735 //y=1.495
r60 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=73.675 //y=0.615 //x2=73.675 //y2=0.49
r61 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=73.675 //y=0.615 //x2=73.675 //y2=0.88
r62 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=72.79 //y=0.53 //x2=72.705 //y2=0.49
r63 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=72.79 //y=0.53 //x2=73.19 //y2=0.53
r64 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=73.59 //y=0.53 //x2=73.675 //y2=0.49
r65 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=73.59 //y=0.53 //x2=73.19 //y2=0.53
r66 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=72.705 //y=1.495 //x2=72.705 //y2=1.62
r67 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=72.705 //y=1.495 //x2=72.705 //y2=0.88
r68 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=72.705 //y=0.615 //x2=72.705 //y2=0.49
r69 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=72.705 //y=0.615 //x2=72.705 //y2=0.88
r70 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=71.82 //y=1.58 //x2=71.735 //y2=1.62
r71 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=71.82 //y=1.58 //x2=72.22 //y2=1.58
r72 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=72.62 //y=1.58 //x2=72.705 //y2=1.62
r73 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=72.62 //y=1.58 //x2=72.22 //y2=1.58
r74 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=71.735 //y=1.495 //x2=71.735 //y2=1.62
r75 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=71.735 //y=1.495 //x2=71.735 //y2=0.88
ends PM_TMRDFFQNX1\%noxref_49

