magic
tech sky130A
magscale 1 2
timestamp 1652395794
<< metal1 >>
rect 427 871 2651 905
rect 258 797 2793 831
rect 2841 797 3990 831
rect 833 723 1132 757
rect 1213 723 3163 757
rect 685 649 1427 683
rect 1509 649 1797 683
rect 2165 649 2478 683
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 814 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 666 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform -1 0 444 0 -1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 222 0 -1 814
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_0
timestamp 1652319931
transform 1 0 0 0 1 0
box -87 -34 1049 1550
use nand2x1_pcell  nand2x1_pcell_0
timestamp 1652323009
transform 1 0 962 0 1 0
box -87 -34 753 1550
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform -1 0 2146 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 1998 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 1850 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform 1 0 1480 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform 1 0 1184 0 1 740
box -53 -33 29 33
use nand2x1_pcell  nand2x1_pcell_1
timestamp 1652323009
transform 1 0 1628 0 1 0
box -87 -34 753 1550
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 3182 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 2812 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_18
timestamp 1648061256
transform 1 0 2664 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform 1 0 2516 0 1 666
box -53 -33 29 33
use nand2x1_pcell  nand2x1_pcell_2
timestamp 1652323009
transform 1 0 2294 0 1 0
box -87 -34 753 1550
use nand2x1_pcell  nand2x1_pcell_3
timestamp 1652323009
transform 1 0 2960 0 1 0
box -87 -34 753 1550
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform 1 0 3996 0 1 814
box -53 -33 29 33
use nand2x1_pcell  nand2x1_pcell_4
timestamp 1652323009
transform 1 0 3626 0 1 0
box -87 -34 753 1550
<< end >>
