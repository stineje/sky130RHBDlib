magic
tech sky130A
magscale 1 2
timestamp 1652328347
<< metal1 >>
rect 315 501 569 535
use invx1_pcell  invx1_pcell_1
timestamp 1652321374
transform 1 0 444 0 1 0
box -87 -34 531 1550
use invx1_pcell  invx1_pcell_0
timestamp 1652321374
transform 1 0 0 0 1 0
box -87 -34 531 1550
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 592 0 1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 296 0 -1 518
box -53 -33 29 33
<< end >>
