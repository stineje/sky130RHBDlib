* SPICE3 file created from MUX2X1.ext - technology: sky130A

.subckt MUX2X1 Y A0 A1 S VPB VNB
X0 a_661_1004# a_787_383# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6.14e+12p ps=5.014e+07u w=2e+06u l=150000u M=2
X1 VPB a_1453_383# a_1327_1004# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X2 a_185_182# S VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.6781e+12p ps=1.281e+07u w=3e+06u l=150000u
X3 a_661_1004# a_787_383# a_556_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4 a_661_1004# S VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X5 VPB S a_185_182# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X6 a_1327_1004# a_185_182# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X7 VPB a_1327_1004# a_1993_1004# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X8 VPB a_661_1004# a_1993_1004# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X9 VNB a_661_1004# a_1888_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X10 VNB a_185_182# a_1222_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X11 a_1993_1004# a_1327_1004# a_1888_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X12 VNB S a_556_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X13 a_1327_1004# a_1453_383# a_1222_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
.ends
