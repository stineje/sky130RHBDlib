* SPICE3 file created from DLATCH.ext - technology: sky130A

.subckt DLATCH Q D GATE VDD GND
X0 a_661_1004 GATE VDD VDD pshort w=2 l=0.15 M=2
X1 a_1771_1004 D VDD VDD pshort w=2 l=0.15 M=2
X2 a_2405_182 a_1771_1004 VDD VDD pshort w=2 l=0.15 M=2
X3 Q a_3007_383 a_2795_1005 VDD pshort w=2 l=0.15 M=2
X4 a_185_182 D GND GND nshort w=3 l=0.15
X5 a_3461_1005 a_2405_182 a_3007_383 VDD pshort w=2 l=0.15 M=2
X6 a_661_1004 GATE a_556_73 GND nshort w=3 l=0.15
X7 a_661_1004 a_185_182 VDD VDD pshort w=2 l=0.15 M=2
X8 a_1771_1004 GATE VDD VDD pshort w=2 l=0.15 M=2
X9 a_2795_1005 a_1295_182 VDD VDD pshort w=2 l=0.15 M=2
X10 VDD Q a_3461_1005 VDD pshort w=2 l=0.15 M=2
X11 VDD D a_185_182 VDD pshort w=2 l=0.15 M=2
X12 VDD a_661_1004 a_1295_182 VDD pshort w=2 l=0.15 M=2
X13 GND GATE a_1666_73 GND nshort w=3 l=0.15
X14 a_3007_383 a_2405_182 GND GND nshort w=3 l=0.15
X15 Q a_1295_182 GND GND nshort w=3 l=0.15
X16 Q a_3007_383 GND GND nshort w=3 l=0.15
X17 a_1295_182 a_661_1004 GND GND nshort w=3 l=0.15
X18 a_1771_1004 D a_1666_73 GND nshort w=3 l=0.15
X19 GND a_185_182 a_556_73 GND nshort w=3 l=0.15
X20 a_2405_182 a_1771_1004 GND GND nshort w=3 l=0.15
X21 a_3007_383 Q GND GND nshort w=3 l=0.15
C0 VDD GND 9.82fF
.ends
