magic
tech sky130A
magscale 1 2
timestamp 1669500663
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 2055 945 2089 979
rect 2721 945 2755 979
rect 205 871 239 905
rect 353 871 387 905
rect 945 871 979 905
rect 1241 871 1275 905
rect 1759 871 1793 905
rect 1907 871 1941 905
rect 2425 871 2459 905
rect 3165 871 3199 905
rect 205 797 239 831
rect 1241 797 1275 831
rect 1759 797 1793 831
rect 1907 773 1941 855
rect 3165 797 3199 831
rect 205 723 239 757
rect 353 723 387 757
rect 1907 723 1941 757
rect 2055 723 2089 757
rect 2721 723 2755 757
rect 3165 723 3199 757
rect 205 649 239 683
rect 353 649 387 683
rect 945 649 979 683
rect 1241 649 1275 683
rect 1759 649 1793 683
rect 2055 649 2089 683
rect 3165 649 3199 683
rect 205 575 239 609
rect 353 575 387 609
rect 945 575 979 609
rect 1241 575 1275 609
rect 1759 575 1793 609
rect 1981 575 2015 609
rect 3165 575 3199 609
rect 205 501 239 535
rect 353 501 387 535
rect 945 501 979 535
rect 1241 501 1275 535
rect 2721 501 2755 535
rect 3165 501 3199 535
rect 945 427 979 461
rect 2055 427 2089 461
rect 2721 427 2755 461
<< metal1 >>
rect -34 1446 3364 1514
rect 1977 871 2413 905
rect 275 797 1229 831
rect 423 723 1871 757
rect -34 -34 3364 34
use and2x1_pcell  and2x1_pcell_0 pcells
timestamp 1669500627
transform 1 0 0 0 1 0
box -87 -34 1197 1550
use li1_M1_contact  li1_M1_contact_0 pcells
timestamp 1648061256
transform -1 0 370 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 222 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 1924 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 1924 0 -1 888
box -53 -33 29 33
use xor2X1_pcell  xor2X1_pcell_0 pcells
timestamp 1669500627
transform 1 0 1110 0 1 0
box -87 -34 2307 1550
<< labels >>
rlabel locali 2721 723 2755 757 1 SUM
port 1 nsew signal output
rlabel locali 2055 723 2089 757 1 SUM
port 1 nsew signal output
rlabel locali 2721 427 2755 461 1 SUM
port 1 nsew signal output
rlabel locali 2721 501 2755 535 1 SUM
port 1 nsew signal output
rlabel locali 2721 945 2755 979 1 SUM
port 1 nsew signal output
rlabel locali 2055 649 2089 683 1 SUM
port 1 nsew signal output
rlabel locali 2055 427 2089 461 1 SUM
port 1 nsew signal output
rlabel locali 2055 945 2089 979 1 SUM
port 1 nsew signal output
rlabel locali 945 501 979 535 1 COUT
port 2 nsew signal output
rlabel locali 945 427 979 461 1 COUT
port 2 nsew signal output
rlabel locali 945 649 979 683 1 COUT
port 2 nsew signal output
rlabel locali 945 871 979 905 1 COUT
port 2 nsew signal output
rlabel locali 945 575 979 609 1 COUT
port 2 nsew signal output
rlabel locali 205 797 239 831 1 A
port 3 nsew signal input
rlabel locali 205 871 239 905 1 A
port 3 nsew signal input
rlabel locali 205 723 239 757 1 A
port 3 nsew signal input
rlabel locali 205 649 239 683 1 A
port 3 nsew signal input
rlabel locali 205 575 239 609 1 A
port 3 nsew signal input
rlabel locali 205 501 239 535 1 A
port 3 nsew signal input
rlabel locali 1241 871 1275 905 1 A
port 3 nsew signal input
rlabel locali 1241 797 1275 831 1 A
port 3 nsew signal input
rlabel locali 1241 649 1275 683 1 A
port 3 nsew signal input
rlabel locali 1241 575 1275 609 1 A
port 3 nsew signal input
rlabel locali 1241 501 1275 535 1 A
port 3 nsew signal input
rlabel locali 1759 871 1793 905 1 A
port 3 nsew signal input
rlabel locali 1759 797 1793 831 1 A
port 3 nsew signal input
rlabel locali 1759 649 1793 683 1 A
port 3 nsew signal input
rlabel locali 1759 575 1793 609 1 A
port 3 nsew signal input
rlabel locali 353 723 387 757 1 B
port 4 nsew signal input
rlabel locali 353 649 387 683 1 B
port 4 nsew signal input
rlabel locali 353 575 387 609 1 B
port 4 nsew signal input
rlabel locali 353 501 387 535 1 B
port 4 nsew signal input
rlabel locali 353 871 387 905 1 B
port 4 nsew signal input
rlabel locali 1907 723 1941 757 1 B
port 4 nsew signal input
rlabel locali 1907 797 1941 831 1 B
port 4 nsew signal input
rlabel locali 1907 871 1941 905 1 B
port 4 nsew signal input
rlabel locali 3165 723 3199 757 1 B
port 4 nsew signal input
rlabel locali 1981 575 2015 609 1 B
port 4 nsew signal input
rlabel locali 3165 575 3199 609 1 B
port 4 nsew signal input
rlabel locali 3165 649 3199 683 1 B
port 4 nsew signal input
rlabel locali 3165 501 3199 535 1 B
port 4 nsew signal input
rlabel locali 3165 797 3199 831 1 B
port 4 nsew signal input
rlabel locali 3165 871 3199 905 1 B
port 4 nsew signal input
rlabel locali 2425 871 2459 905 1 B
port 4 nsew signal input
rlabel metal1 -34 1446 3364 1514 1 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 -34 -34 3364 34 1 VGND
port 6 nsew ground bidirectional abutment
rlabel nwell 57 1463 91 1497 1 VPB
port 7 nsew power bidirectional
rlabel pwell 57 -17 91 17 1 VNB
port 8 nsew ground bidirectional
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
