VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DLATCH
  CLASS CORE ;
  FOREIGN DLATCH ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.980 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.027250 ;
    ANTENNADIFFAREA 0.963050 ;
    PORT
      LAYER li1 ;
        RECT 15.345 5.295 15.515 6.565 ;
        RECT 15.345 5.125 15.995 5.295 ;
        RECT 15.825 1.740 15.995 5.125 ;
        RECT 17.520 4.710 17.690 4.870 ;
        RECT 17.520 4.540 17.845 4.710 ;
        RECT 17.675 1.915 17.845 4.540 ;
        RECT 14.415 1.570 15.995 1.740 ;
        RECT 14.415 0.835 14.585 1.570 ;
        RECT 15.385 0.835 15.555 1.570 ;
      LAYER mcon ;
        RECT 15.825 3.245 15.995 3.415 ;
        RECT 17.675 3.245 17.845 3.415 ;
      LAYER met1 ;
        RECT 15.795 3.415 16.025 3.445 ;
        RECT 17.645 3.415 17.875 3.445 ;
        RECT 15.765 3.245 17.905 3.415 ;
        RECT 15.795 3.215 16.025 3.245 ;
        RECT 17.645 3.215 17.875 3.245 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.054500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.920 0.825 4.865 ;
        RECT 9.565 4.710 9.735 4.865 ;
        RECT 9.535 4.535 9.735 4.710 ;
        RECT 9.535 1.915 9.705 4.535 ;
      LAYER mcon ;
        RECT 0.655 3.985 0.825 4.155 ;
        RECT 9.535 3.985 9.705 4.155 ;
      LAYER met1 ;
        RECT 0.625 4.155 0.855 4.185 ;
        RECT 9.505 4.155 9.735 4.185 ;
        RECT 0.595 3.985 9.765 4.155 ;
        RECT 0.625 3.955 0.855 3.985 ;
        RECT 9.505 3.955 9.735 3.985 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 4.015 4.710 4.185 4.865 ;
        RECT 3.985 4.535 4.185 4.710 ;
        RECT 3.985 1.915 4.155 4.535 ;
        RECT 8.795 1.915 8.965 4.865 ;
      LAYER mcon ;
        RECT 3.985 2.875 4.155 3.045 ;
        RECT 8.795 2.875 8.965 3.045 ;
      LAYER met1 ;
        RECT 3.955 3.045 4.185 3.075 ;
        RECT 8.765 3.045 8.995 3.075 ;
        RECT 3.925 2.875 9.025 3.045 ;
        RECT 3.955 2.845 4.185 2.875 ;
        RECT 8.765 2.845 8.995 2.875 ;
    END
  END GATE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 20.415 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 20.150 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.590 5.185 0.760 7.230 ;
        RECT 1.470 5.185 1.640 7.230 ;
        RECT 2.050 4.110 2.390 7.230 ;
        RECT 2.925 5.135 3.095 7.230 ;
        RECT 3.805 5.555 3.975 7.230 ;
        RECT 4.685 5.555 4.855 7.230 ;
        RECT 5.380 4.110 5.720 7.230 ;
        RECT 6.140 5.185 6.310 7.230 ;
        RECT 7.020 5.185 7.190 7.230 ;
        RECT 7.600 4.110 7.940 7.230 ;
        RECT 8.475 5.135 8.645 7.230 ;
        RECT 9.355 5.555 9.525 7.230 ;
        RECT 10.235 5.555 10.405 7.230 ;
        RECT 10.930 4.110 11.270 7.230 ;
        RECT 11.690 5.185 11.860 7.230 ;
        RECT 12.570 5.185 12.740 7.230 ;
        RECT 13.150 4.110 13.490 7.230 ;
        RECT 14.465 5.555 14.635 7.230 ;
        RECT 16.480 4.110 16.820 7.230 ;
        RECT 17.795 5.555 17.965 7.230 ;
        RECT 19.810 4.110 20.150 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.245 7.315 3.415 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.575 7.315 6.745 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
        RECT 9.905 7.315 10.075 7.485 ;
        RECT 10.275 7.315 10.445 7.485 ;
        RECT 10.645 7.315 10.815 7.485 ;
        RECT 11.385 7.315 11.555 7.485 ;
        RECT 11.755 7.315 11.925 7.485 ;
        RECT 12.125 7.315 12.295 7.485 ;
        RECT 12.495 7.315 12.665 7.485 ;
        RECT 12.865 7.315 13.035 7.485 ;
        RECT 13.605 7.315 13.775 7.485 ;
        RECT 13.975 7.315 14.145 7.485 ;
        RECT 14.345 7.315 14.515 7.485 ;
        RECT 14.715 7.315 14.885 7.485 ;
        RECT 15.085 7.315 15.255 7.485 ;
        RECT 15.455 7.315 15.625 7.485 ;
        RECT 15.825 7.315 15.995 7.485 ;
        RECT 16.195 7.315 16.365 7.485 ;
        RECT 16.935 7.315 17.105 7.485 ;
        RECT 17.305 7.315 17.475 7.485 ;
        RECT 17.675 7.315 17.845 7.485 ;
        RECT 18.045 7.315 18.215 7.485 ;
        RECT 18.415 7.315 18.585 7.485 ;
        RECT 18.785 7.315 18.955 7.485 ;
        RECT 19.155 7.315 19.325 7.485 ;
        RECT 19.525 7.315 19.695 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 20.150 7.570 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 20.150 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.545 0.620 0.715 1.750 ;
        RECT 1.515 0.620 1.685 1.750 ;
        RECT 0.545 0.450 1.685 0.620 ;
        RECT 0.545 0.170 0.715 0.450 ;
        RECT 1.030 0.170 1.200 0.450 ;
        RECT 1.515 0.170 1.685 0.450 ;
        RECT 2.050 0.170 2.390 2.720 ;
        RECT 3.315 0.170 3.485 1.120 ;
        RECT 5.380 0.170 5.720 2.720 ;
        RECT 6.095 0.620 6.265 1.750 ;
        RECT 7.065 0.620 7.235 1.750 ;
        RECT 6.095 0.450 7.235 0.620 ;
        RECT 6.095 0.170 6.265 0.450 ;
        RECT 6.580 0.170 6.750 0.450 ;
        RECT 7.065 0.170 7.235 0.450 ;
        RECT 7.600 0.170 7.940 2.720 ;
        RECT 8.865 0.170 9.035 1.120 ;
        RECT 10.930 0.170 11.270 2.720 ;
        RECT 11.645 0.620 11.815 1.750 ;
        RECT 12.615 0.620 12.785 1.750 ;
        RECT 11.645 0.450 12.785 0.620 ;
        RECT 11.645 0.170 11.815 0.450 ;
        RECT 12.130 0.170 12.300 0.450 ;
        RECT 12.615 0.170 12.785 0.450 ;
        RECT 13.150 0.170 13.490 2.720 ;
        RECT 13.930 0.615 14.100 1.745 ;
        RECT 14.900 0.615 15.070 1.390 ;
        RECT 15.870 0.615 16.040 1.390 ;
        RECT 13.930 0.445 16.040 0.615 ;
        RECT 13.930 0.170 14.100 0.445 ;
        RECT 14.415 0.170 14.585 0.445 ;
        RECT 14.900 0.170 15.070 0.445 ;
        RECT 15.385 0.170 15.555 0.445 ;
        RECT 15.870 0.170 16.040 0.445 ;
        RECT 16.480 0.170 16.820 2.720 ;
        RECT 17.260 0.615 17.430 1.745 ;
        RECT 18.230 0.615 18.400 1.390 ;
        RECT 19.200 0.615 19.370 1.390 ;
        RECT 17.260 0.445 19.370 0.615 ;
        RECT 17.260 0.170 17.430 0.445 ;
        RECT 17.745 0.170 17.915 0.445 ;
        RECT 18.230 0.170 18.400 0.445 ;
        RECT 18.715 0.170 18.885 0.445 ;
        RECT 19.200 0.170 19.370 0.445 ;
        RECT 19.810 0.170 20.150 2.720 ;
        RECT -0.170 -0.170 20.150 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.245 -0.085 3.415 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
        RECT 9.905 -0.085 10.075 0.085 ;
        RECT 10.275 -0.085 10.445 0.085 ;
        RECT 10.645 -0.085 10.815 0.085 ;
        RECT 11.385 -0.085 11.555 0.085 ;
        RECT 11.755 -0.085 11.925 0.085 ;
        RECT 12.125 -0.085 12.295 0.085 ;
        RECT 12.495 -0.085 12.665 0.085 ;
        RECT 12.865 -0.085 13.035 0.085 ;
        RECT 13.605 -0.085 13.775 0.085 ;
        RECT 13.975 -0.085 14.145 0.085 ;
        RECT 14.345 -0.085 14.515 0.085 ;
        RECT 14.715 -0.085 14.885 0.085 ;
        RECT 15.085 -0.085 15.255 0.085 ;
        RECT 15.455 -0.085 15.625 0.085 ;
        RECT 15.825 -0.085 15.995 0.085 ;
        RECT 16.195 -0.085 16.365 0.085 ;
        RECT 16.935 -0.085 17.105 0.085 ;
        RECT 17.305 -0.085 17.475 0.085 ;
        RECT 17.675 -0.085 17.845 0.085 ;
        RECT 18.045 -0.085 18.215 0.085 ;
        RECT 18.415 -0.085 18.585 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.155 -0.085 19.325 0.085 ;
        RECT 19.525 -0.085 19.695 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 20.150 0.170 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 1.030 4.665 1.200 7.020 ;
        RECT 3.365 5.285 3.535 7.020 ;
        RECT 4.245 5.285 4.415 7.020 ;
        RECT 3.365 5.115 4.895 5.285 ;
        RECT 1.030 4.495 1.565 4.665 ;
        RECT 1.395 2.165 1.565 4.495 ;
        RECT 1.025 1.995 1.565 2.165 ;
        RECT 1.025 0.840 1.195 1.995 ;
        RECT 3.245 1.915 3.415 4.865 ;
        RECT 2.830 1.665 3.000 1.745 ;
        RECT 3.800 1.665 3.970 1.745 ;
        RECT 4.725 1.740 4.895 5.115 ;
        RECT 6.205 1.920 6.375 4.865 ;
        RECT 6.580 4.665 6.750 7.020 ;
        RECT 8.915 5.285 9.085 7.020 ;
        RECT 9.795 5.285 9.965 7.020 ;
        RECT 8.915 5.115 10.445 5.285 ;
        RECT 6.580 4.495 7.115 4.665 ;
        RECT 6.945 2.165 7.115 4.495 ;
        RECT 6.575 1.995 7.115 2.165 ;
        RECT 2.830 1.495 3.970 1.665 ;
        RECT 2.830 0.365 3.000 1.495 ;
        RECT 3.800 0.615 3.970 1.495 ;
        RECT 4.285 1.570 4.895 1.740 ;
        RECT 4.285 0.835 4.455 1.570 ;
        RECT 4.770 0.615 4.940 1.385 ;
        RECT 6.575 0.840 6.745 1.995 ;
        RECT 8.380 1.665 8.550 1.745 ;
        RECT 9.350 1.665 9.520 1.745 ;
        RECT 10.275 1.740 10.445 5.115 ;
        RECT 11.755 1.920 11.925 4.865 ;
        RECT 12.130 4.665 12.300 7.020 ;
        RECT 14.025 5.295 14.195 7.025 ;
        RECT 14.905 6.825 15.955 6.995 ;
        RECT 14.905 5.295 15.075 6.825 ;
        RECT 15.785 5.555 15.955 6.825 ;
        RECT 14.025 5.125 15.075 5.295 ;
        RECT 17.355 5.295 17.525 7.025 ;
        RECT 18.235 6.825 19.285 6.995 ;
        RECT 18.235 5.295 18.405 6.825 ;
        RECT 17.355 5.125 18.405 5.295 ;
        RECT 18.675 5.295 18.845 6.565 ;
        RECT 19.115 5.555 19.285 6.825 ;
        RECT 18.675 5.125 19.325 5.295 ;
        RECT 14.190 4.710 14.360 4.870 ;
        RECT 15.120 4.710 15.290 4.870 ;
        RECT 18.450 4.710 18.620 4.870 ;
        RECT 12.130 4.495 12.665 4.665 ;
        RECT 14.190 4.540 14.515 4.710 ;
        RECT 12.495 2.165 12.665 4.495 ;
        RECT 12.125 1.995 12.665 2.165 ;
        RECT 8.380 1.495 9.520 1.665 ;
        RECT 3.800 0.445 4.940 0.615 ;
        RECT 3.800 0.365 3.970 0.445 ;
        RECT 4.770 0.365 4.940 0.445 ;
        RECT 8.380 0.365 8.550 1.495 ;
        RECT 9.350 0.615 9.520 1.495 ;
        RECT 9.835 1.570 10.445 1.740 ;
        RECT 9.835 0.835 10.005 1.570 ;
        RECT 10.320 0.615 10.490 1.385 ;
        RECT 12.125 0.840 12.295 1.995 ;
        RECT 14.345 1.915 14.515 4.540 ;
        RECT 15.085 4.540 15.290 4.710 ;
        RECT 18.415 4.540 18.620 4.710 ;
        RECT 15.085 1.915 15.255 4.540 ;
        RECT 18.415 1.915 18.585 4.540 ;
        RECT 19.155 1.740 19.325 5.125 ;
        RECT 17.745 1.570 19.325 1.740 ;
        RECT 17.745 0.835 17.915 1.570 ;
        RECT 18.715 0.835 18.885 1.570 ;
        RECT 9.350 0.445 10.490 0.615 ;
        RECT 9.350 0.365 9.520 0.445 ;
        RECT 10.320 0.365 10.490 0.445 ;
      LAYER mcon ;
        RECT 1.395 3.615 1.565 3.785 ;
        RECT 3.245 3.615 3.415 3.785 ;
        RECT 4.725 3.245 4.895 3.415 ;
        RECT 6.205 3.245 6.375 3.415 ;
        RECT 6.945 3.615 7.115 3.785 ;
        RECT 10.275 3.245 10.445 3.415 ;
        RECT 11.755 3.245 11.925 3.415 ;
        RECT 12.495 3.985 12.665 4.155 ;
        RECT 14.345 3.615 14.515 3.785 ;
        RECT 15.085 3.615 15.255 3.785 ;
        RECT 18.415 3.985 18.585 4.155 ;
        RECT 19.155 3.615 19.325 3.785 ;
      LAYER met1 ;
        RECT 12.465 4.155 12.695 4.185 ;
        RECT 18.385 4.155 18.615 4.185 ;
        RECT 12.435 3.985 18.645 4.155 ;
        RECT 12.465 3.955 12.695 3.985 ;
        RECT 18.385 3.955 18.615 3.985 ;
        RECT 1.365 3.785 1.595 3.815 ;
        RECT 3.215 3.785 3.445 3.815 ;
        RECT 6.915 3.785 7.145 3.815 ;
        RECT 14.315 3.785 14.545 3.815 ;
        RECT 15.055 3.785 15.285 3.815 ;
        RECT 19.125 3.785 19.355 3.815 ;
        RECT 1.335 3.615 3.475 3.785 ;
        RECT 6.885 3.615 14.575 3.785 ;
        RECT 15.025 3.615 19.385 3.785 ;
        RECT 1.365 3.585 1.595 3.615 ;
        RECT 3.215 3.585 3.445 3.615 ;
        RECT 6.915 3.585 7.145 3.615 ;
        RECT 14.315 3.585 14.545 3.615 ;
        RECT 15.055 3.585 15.285 3.615 ;
        RECT 19.125 3.585 19.355 3.615 ;
        RECT 4.695 3.415 4.925 3.445 ;
        RECT 6.175 3.415 6.405 3.445 ;
        RECT 10.245 3.415 10.475 3.445 ;
        RECT 11.725 3.415 11.955 3.445 ;
        RECT 4.665 3.245 6.435 3.415 ;
        RECT 10.215 3.245 11.985 3.415 ;
        RECT 4.695 3.215 4.925 3.245 ;
        RECT 6.175 3.215 6.405 3.245 ;
        RECT 10.245 3.215 10.475 3.245 ;
        RECT 11.725 3.215 11.955 3.245 ;
  END
END DLATCH
END LIBRARY

