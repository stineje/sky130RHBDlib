* SPICE3 file created from TMRDFFQX1.ext - technology: sky130A

.subckt TMRDFFQX1 Q D CLK VDD GND
X0 GND dffx1_pcell_0/m1_2165_649# dffx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X1 dffx1_pcell_0/m1_258_797# CLK dffx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X2 VDD dffx1_pcell_0/m1_2165_649# dffx1_pcell_0/m1_258_797# VDD pshort w=2 l=0.15
X3 VDD CLK dffx1_pcell_0/m1_258_797# VDD pshort w=2 l=0.15
X4 GND dffx1_pcell_0/m1_833_723# dffx1_pcell_0/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X5 m1_3495_723# m1_3348_575# dffx1_pcell_0/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X6 VDD dffx1_pcell_0/m1_833_723# m1_3495_723# VDD pshort w=2 l=0.15
X7 VDD m1_3348_575# m1_3495_723# VDD pshort w=2 l=0.15
X8 GND m1_3495_723# dffx1_pcell_0/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X9 m1_3348_575# dffx1_pcell_0/m1_258_797# dffx1_pcell_0/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X10 VDD m1_3495_723# m1_3348_575# VDD pshort w=2 l=0.15
X11 VDD dffx1_pcell_0/m1_258_797# m1_3348_575# VDD pshort w=2 l=0.15
X12 GND dffx1_pcell_0/m1_258_797# dffx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X13 dffx1_pcell_0/m1_833_723# dffx1_pcell_0/m1_685_649# dffx1_pcell_0/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X14 dffx1_pcell_0/nand3x1_pcell_0/li_393_182# CLK dffx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X15 VDD dffx1_pcell_0/m1_258_797# dffx1_pcell_0/m1_833_723# VDD pshort w=2 l=0.15
X16 VDD CLK dffx1_pcell_0/m1_833_723# VDD pshort w=2 l=0.15
X17 VDD dffx1_pcell_0/m1_685_649# dffx1_pcell_0/m1_833_723# VDD pshort w=2 l=0.15
X18 GND dffx1_pcell_0/m1_833_723# dffx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X19 dffx1_pcell_0/m1_685_649# D dffx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X20 VDD dffx1_pcell_0/m1_833_723# dffx1_pcell_0/m1_685_649# VDD pshort w=2 l=0.15
X21 VDD D dffx1_pcell_0/m1_685_649# VDD pshort w=2 l=0.15
X22 GND dffx1_pcell_0/m1_685_649# dffx1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X23 dffx1_pcell_0/m1_2165_649# dffx1_pcell_0/m1_258_797# dffx1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X24 VDD dffx1_pcell_0/m1_685_649# dffx1_pcell_0/m1_2165_649# VDD pshort w=2 l=0.15
X25 VDD dffx1_pcell_0/m1_258_797# dffx1_pcell_0/m1_2165_649# VDD pshort w=2 l=0.15
X26 GND dffx1_pcell_1/m1_2165_649# dffx1_pcell_1/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X27 dffx1_pcell_1/m1_258_797# CLK dffx1_pcell_1/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X28 VDD dffx1_pcell_1/m1_2165_649# dffx1_pcell_1/m1_258_797# VDD pshort w=2 l=0.15
X29 VDD CLK dffx1_pcell_1/m1_258_797# VDD pshort w=2 l=0.15
X30 GND dffx1_pcell_1/m1_833_723# dffx1_pcell_1/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X31 m1_7741_723# m1_7639_427# dffx1_pcell_1/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X32 VDD dffx1_pcell_1/m1_833_723# m1_7741_723# VDD pshort w=2 l=0.15
X33 VDD m1_7639_427# m1_7741_723# VDD pshort w=2 l=0.15
X34 GND m1_7741_723# dffx1_pcell_1/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X35 m1_7639_427# dffx1_pcell_1/m1_258_797# dffx1_pcell_1/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X36 VDD m1_7741_723# m1_7639_427# VDD pshort w=2 l=0.15
X37 VDD dffx1_pcell_1/m1_258_797# m1_7639_427# VDD pshort w=2 l=0.15
X38 GND dffx1_pcell_1/m1_258_797# dffx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X39 dffx1_pcell_1/m1_833_723# dffx1_pcell_1/m1_685_649# dffx1_pcell_1/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X40 dffx1_pcell_1/nand3x1_pcell_0/li_393_182# CLK dffx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X41 VDD dffx1_pcell_1/m1_258_797# dffx1_pcell_1/m1_833_723# VDD pshort w=2 l=0.15
X42 VDD CLK dffx1_pcell_1/m1_833_723# VDD pshort w=2 l=0.15
X43 VDD dffx1_pcell_1/m1_685_649# dffx1_pcell_1/m1_833_723# VDD pshort w=2 l=0.15
X44 GND dffx1_pcell_1/m1_833_723# dffx1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X45 dffx1_pcell_1/m1_685_649# D dffx1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X46 VDD dffx1_pcell_1/m1_833_723# dffx1_pcell_1/m1_685_649# VDD pshort w=2 l=0.15
X47 VDD D dffx1_pcell_1/m1_685_649# VDD pshort w=2 l=0.15
X48 GND dffx1_pcell_1/m1_685_649# dffx1_pcell_1/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X49 dffx1_pcell_1/m1_2165_649# dffx1_pcell_1/m1_258_797# dffx1_pcell_1/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X50 VDD dffx1_pcell_1/m1_685_649# dffx1_pcell_1/m1_2165_649# VDD pshort w=2 l=0.15
X51 VDD dffx1_pcell_1/m1_258_797# dffx1_pcell_1/m1_2165_649# VDD pshort w=2 l=0.15
X52 GND dffx1_pcell_2/m1_2165_649# dffx1_pcell_2/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X53 dffx1_pcell_2/m1_258_797# CLK dffx1_pcell_2/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X54 VDD dffx1_pcell_2/m1_2165_649# dffx1_pcell_2/m1_258_797# VDD pshort w=2 l=0.15
X55 VDD CLK dffx1_pcell_2/m1_258_797# VDD pshort w=2 l=0.15
X56 GND dffx1_pcell_2/m1_833_723# dffx1_pcell_2/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X57 m1_12079_871# m1_11931_723# dffx1_pcell_2/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X58 VDD dffx1_pcell_2/m1_833_723# m1_12079_871# VDD pshort w=2 l=0.15
X59 VDD m1_11931_723# m1_12079_871# VDD pshort w=2 l=0.15
X60 GND m1_12079_871# dffx1_pcell_2/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X61 m1_11931_723# dffx1_pcell_2/m1_258_797# dffx1_pcell_2/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X62 VDD m1_12079_871# m1_11931_723# VDD pshort w=2 l=0.15
X63 VDD dffx1_pcell_2/m1_258_797# m1_11931_723# VDD pshort w=2 l=0.15
X64 GND dffx1_pcell_2/m1_258_797# dffx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X65 dffx1_pcell_2/m1_833_723# dffx1_pcell_2/m1_685_649# dffx1_pcell_2/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X66 dffx1_pcell_2/nand3x1_pcell_0/li_393_182# CLK dffx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X67 VDD dffx1_pcell_2/m1_258_797# dffx1_pcell_2/m1_833_723# VDD pshort w=2 l=0.15
X68 VDD CLK dffx1_pcell_2/m1_833_723# VDD pshort w=2 l=0.15
X69 VDD dffx1_pcell_2/m1_685_649# dffx1_pcell_2/m1_833_723# VDD pshort w=2 l=0.15
X70 GND dffx1_pcell_2/m1_833_723# dffx1_pcell_2/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X71 dffx1_pcell_2/m1_685_649# D dffx1_pcell_2/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X72 VDD dffx1_pcell_2/m1_833_723# dffx1_pcell_2/m1_685_649# VDD pshort w=2 l=0.15
X73 VDD D dffx1_pcell_2/m1_685_649# VDD pshort w=2 l=0.15
X74 GND dffx1_pcell_2/m1_685_649# dffx1_pcell_2/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X75 dffx1_pcell_2/m1_2165_649# dffx1_pcell_2/m1_258_797# dffx1_pcell_2/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X76 VDD dffx1_pcell_2/m1_685_649# dffx1_pcell_2/m1_2165_649# VDD pshort w=2 l=0.15
X77 VDD dffx1_pcell_2/m1_258_797# dffx1_pcell_2/m1_2165_649# VDD pshort w=2 l=0.15
X78 GND m1_11931_723# voter3x1_pcell_0/votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X79 GND m1_11931_723# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X80 GND m1_3348_575# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X81 voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# m1_11931_723# VDD VDD pshort w=2 l=0.15
X82 voter3x1_pcell_0/m1_1867_797# m1_3348_575# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X83 voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# m1_7639_427# VDD VDD pshort w=2 l=0.15
X84 voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# m1_3348_575# voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X85 voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# m1_11931_723# voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X86 voter3x1_pcell_0/m1_1867_797# m1_3348_575# voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X87 voter3x1_pcell_0/m1_1867_797# m1_7639_427# voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X88 voter3x1_pcell_0/m1_1867_797# m1_7639_427# voter3x1_pcell_0/votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X89 voter3x1_pcell_0/m1_1867_797# m1_7639_427# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X90 Q voter3x1_pcell_0/m1_1867_797# GND GND nshort w=3 l=0.15
X91 VDD voter3x1_pcell_0/m1_1867_797# Q VDD pshort w=2 l=0.15
C0 dffx1_pcell_1/m1_258_797# dffx1_pcell_1/m1_833_723# 3.00fF
C1 m1_7639_427# D 2.68fF
C2 dffx1_pcell_2/m1_258_797# CLK 3.24fF
C3 VDD m1_3348_575# 2.13fF
C4 dffx1_pcell_0/m1_258_797# CLK 4.48fF
C5 m1_7639_427# m1_3348_575# 2.76fF
C6 dffx1_pcell_1/m1_258_797# CLK 4.80fF
C7 VDD dffx1_pcell_2/m1_258_797# 2.53fF
C8 m1_7639_427# VDD 2.21fF
C9 dffx1_pcell_0/m1_258_797# dffx1_pcell_0/m1_833_723# 3.00fF
C10 dffx1_pcell_0/m1_258_797# VDD 2.51fF
C11 m1_3348_575# D 7.42fF
C12 dffx1_pcell_1/m1_258_797# VDD 2.49fF
C13 VDD voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# 2.08fF
C14 VDD CLK 4.72fF
C15 dffx1_pcell_2/m1_258_797# dffx1_pcell_2/m1_833_723# 3.01fF
.ends
