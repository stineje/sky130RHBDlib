* SPICE3 file created from DFFSNRNQX1.ext - technology: sky130A

.subckt DFFSNRNQX1 Q D CLK SN RN VDD GND
X0 VDD RN a_277_1004 VDD pshort w=2 l=0.15 M=2
X1 a_599_943 a_1561_943 VDD VDD pshort w=2 l=0.15 M=2
X2 VDD RN a_1561_943 VDD pshort w=2 l=0.15 M=2
X3 GND D a_91_75 GND nshort w=3 l=0.15
X4 VDD SN a_2201_1004 VDD pshort w=2 l=0.15 M=2
X5 a_4125_1004 a_599_943 VDD VDD pshort w=2 l=0.15 M=2
X6 a_4125_1004 Q VDD VDD pshort w=2 l=0.15 M=2
X7 a_1561_943 CLK VDD VDD pshort w=2 l=0.15 M=2
X8 VDD a_599_943 a_277_1004 VDD pshort w=2 l=0.15 M=2
X9 VDD a_1561_943 a_2201_1004 VDD pshort w=2 l=0.15 M=2
X10 a_4125_1004 RN VDD VDD pshort w=2 l=0.15 M=2
X11 a_1561_943 a_2201_1004 VDD VDD pshort w=2 l=0.15 M=2
X12 VDD a_4125_1004 Q VDD pshort w=2 l=0.15 M=2
X13 a_372_182 RN a_91_75 GND nshort w=3 l=0.15
X14 a_2201_1004 a_1561_943 a_2296_182 GND nshort w=3 l=0.15
X15 a_4125_1004 Q a_4220_182 GND nshort w=3 l=0.15
X16 a_277_1004 D VDD VDD pshort w=2 l=0.15 M=2
X17 VDD a_277_1004 a_599_943 VDD pshort w=2 l=0.15 M=2
X18 VDD SN Q VDD pshort w=2 l=0.15 M=2
X19 a_599_943 a_1561_943 a_1334_182 GND nshort w=3 l=0.15
X20 GND a_277_1004 a_2015_75 GND nshort w=3 l=0.15
X21 a_1561_943 RN a_3258_182 GND nshort w=3 l=0.15
X22 Q a_1561_943 a_5182_182 GND nshort w=3 l=0.15
X23 VDD CLK a_599_943 VDD pshort w=2 l=0.15 M=2
X24 GND a_2201_1004 a_2977_75 GND nshort w=3 l=0.15
X25 VDD a_1561_943 Q VDD pshort w=2 l=0.15 M=2
X26 GND a_277_1004 a_1053_75 GND nshort w=3 l=0.15
X27 a_4220_182 RN a_3939_75 GND nshort w=3 l=0.15
X28 a_2296_182 SN a_2015_75 GND nshort w=3 l=0.15
X29 GND a_599_943 a_3939_75 GND nshort w=3 l=0.15
X30 a_2201_1004 a_277_1004 VDD VDD pshort w=2 l=0.15 M=2
X31 a_1334_182 CLK a_1053_75 GND nshort w=3 l=0.15
X32 a_3258_182 CLK a_2977_75 GND nshort w=3 l=0.15
X33 a_5182_182 SN a_4901_75 GND nshort w=3 l=0.15
X34 GND a_4125_1004 a_4901_75 GND nshort w=3 l=0.15
X35 a_277_1004 a_599_943 a_372_182 GND nshort w=3 l=0.15
C0 RN a_1561_943 3.42fF
C1 VDD a_1561_943 3.40fF
C2 VDD a_2201_1004 2.07fF
C3 CLK a_599_943 2.41fF
C4 a_599_943 a_1561_943 3.20fF
C5 VDD a_277_1004 2.25fF
C6 VDD a_4125_1004 2.02fF
C7 VDD a_599_943 2.47fF
C8 VDD GND 13.96fF
.ends
