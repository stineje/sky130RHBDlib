* SPICE3 file created from FILL1.ext - technology: sky130A

.subckt FILL1 VPWR VGND VPB VNB
C0 VPWR VPB 0.08fF
C1 VPWR VNB 0.09fF
C2 VPB VNB 1.56fF
.ends
