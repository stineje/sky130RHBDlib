* SPICE3 file created from NOR2X1.ext - technology: sky130A

.subckt NOR2X1 Y A B VPB VNB
M1000 a_198_181.t2 a_343_383# a_131_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_131_1005.t1 a_164_908# VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_131_1005.t2 a_343_383# a_198_181.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t0 a_164_908# a_131_1005.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u



R0 a_131_1005.t0 a_131_1005.n0 101.66
R1 a_131_1005.n0 a_131_1005.t2 101.659
R2 a_131_1005.n0 a_131_1005.t3 14.294
R3 a_131_1005.n0 a_131_1005.t1 14.282
R4 a_198_181.n6 a_198_181.n1 321.065
R5 a_198_181.n6 a_198_181.n5 118.016
R6 a_198_181.n9 a_198_181.n0 55.263
R7 a_198_181.n8 a_198_181.n6 48.405
R8 a_198_181.n5 a_198_181.n4 30
R9 a_198_181.n8 a_198_181.n7 30
R10 a_198_181.n9 a_198_181.n8 25.263
R11 a_198_181.n3 a_198_181.n2 24.383
R12 a_198_181.n5 a_198_181.n3 23.684
R13 a_198_181.n1 a_198_181.t1 14.282
R14 a_198_181.n1 a_198_181.t2 14.282
R15 VNB VNB.n76 300.778
R16 VNB.n63 VNB.n62 76
R17 VNB.n58 VNB.n57 76
R18 VNB.n48 VNB.n47 62.533
R19 VNB.n37 VNB.n36 36.267
R20 VNB.n31 VNB.n28 20.452
R21 VNB.n64 VNB.n63 20.452
R22 VNB.n50 VNB.n43 19.735
R23 VNB.n54 VNB.n42 19.735
R24 VNB.n39 VNB.n10 19.735
R25 VNB.n32 VNB.n13 19.735
R26 VNB.n7 VNB.n6 19.735
R27 VNB.n5 VNB.t0 17.353
R28 VNB.n41 VNB.t1 13.654
R29 VNB.n35 VNB.n34 13.653
R30 VNB.n34 VNB.n33 13.653
R31 VNB.n38 VNB.n37 13.653
R32 VNB.n57 VNB.n56 13.653
R33 VNB.n56 VNB.n55 13.653
R34 VNB.n53 VNB.n52 13.653
R35 VNB.n52 VNB.n51 13.653
R36 VNB.n49 VNB.n48 13.653
R37 VNB.n46 VNB.n45 13.653
R38 VNB.n45 VNB.n44 13.653
R39 VNB.n63 VNB.n0 13.653
R40 VNB VNB.n0 13.653
R41 VNB.n31 VNB.n30 13.653
R42 VNB.n30 VNB.n29 13.653
R43 VNB.n71 VNB.n68 13.577
R44 VNB.n16 VNB.n14 13.276
R45 VNB.n28 VNB.n16 13.276
R46 VNB.n38 VNB.n35 13.276
R47 VNB.n49 VNB.n46 13.276
R48 VNB.n3 VNB.n1 13.276
R49 VNB.n64 VNB.n3 13.276
R50 VNB.n6 VNB.n5 12.837
R51 VNB.n32 VNB.n31 11.661
R52 VNB.n63 VNB.n7 11.661
R53 VNB.n13 VNB.n12 11.605
R54 VNB.n57 VNB.n39 10.764
R55 VNB.n53 VNB.n50 10.764
R56 VNB.n12 VNB.n11 9.809
R57 VNB.n5 VNB.n4 7.566
R58 VNB.n73 VNB.n72 7.5
R59 VNB.n65 VNB.n64 7.5
R60 VNB.n3 VNB.n2 7.5
R61 VNB.n70 VNB.n69 7.5
R62 VNB.n22 VNB.n21 7.5
R63 VNB.n18 VNB.n17 7.5
R64 VNB.n16 VNB.n15 7.5
R65 VNB.n28 VNB.n27 7.5
R66 VNB.t1 VNB.n40 7.04
R67 VNB.n75 VNB.n73 7.011
R68 VNB.n24 VNB.n22 7.011
R69 VNB.n20 VNB.n18 7.011
R70 VNB.n27 VNB.n26 7.01
R71 VNB.n20 VNB.n19 7.01
R72 VNB.n24 VNB.n23 7.01
R73 VNB.n75 VNB.n74 7.01
R74 VNB.n71 VNB.n70 6.788
R75 VNB.n66 VNB.n65 6.788
R76 VNB.n57 VNB.n54 6.638
R77 VNB.n54 VNB.n53 6.638
R78 VNB.n42 VNB.n41 5.774
R79 VNB.n39 VNB.n38 2.511
R80 VNB.n50 VNB.n49 2.511
R81 VNB.n35 VNB.n32 1.614
R82 VNB.n46 VNB.n7 1.614
R83 VNB.n76 VNB.n67 0.921
R84 VNB.n76 VNB.n71 0.476
R85 VNB.n76 VNB.n66 0.475
R86 VNB.n25 VNB.n20 0.246
R87 VNB.n26 VNB.n25 0.246
R88 VNB.n25 VNB.n24 0.246
R89 VNB.n76 VNB.n75 0.246
R90 VNB.n62 VNB 0.198
R91 VNB.n9 VNB.n8 0.136
R92 VNB.n58 VNB.n9 0.136
R93 VNB.n60 VNB.n59 0.136
R94 VNB.n61 VNB.n60 0.136
R95 VNB.n62 VNB.n61 0.136
R96 VNB VNB.n58 0.068
R97 VNB.n59 VNB 0.068
R98 VPB VPB.n74 126.832
R99 VPB.n67 VPB.n66 76
R100 VPB.n43 VPB.n42 44.502
R101 VPB.n46 VPB.n41 41.183
R102 VPB.n61 VPB.n60 35.118
R103 VPB.n71 VPB.n67 20.452
R104 VPB.n40 VPB.n37 20.452
R105 VPB.n41 VPB.t1 14.282
R106 VPB.n41 VPB.t0 14.282
R107 VPB.n40 VPB.n39 13.653
R108 VPB.n39 VPB.n38 13.653
R109 VPB.n59 VPB.n58 13.653
R110 VPB.n58 VPB.n57 13.653
R111 VPB.n56 VPB.n55 13.653
R112 VPB.n55 VPB.n54 13.653
R113 VPB.n53 VPB.n52 13.653
R114 VPB.n52 VPB.n51 13.653
R115 VPB.n50 VPB.n49 13.653
R116 VPB.n49 VPB.n48 13.653
R117 VPB.n45 VPB.n44 13.653
R118 VPB.n44 VPB.n43 13.653
R119 VPB.n16 VPB.n15 13.653
R120 VPB.n15 VPB.n14 13.653
R121 VPB.n67 VPB.n0 13.653
R122 VPB VPB.n0 13.653
R123 VPB.n48 VPB.n47 13.35
R124 VPB.n71 VPB.n70 13.276
R125 VPB.n70 VPB.n68 13.276
R126 VPB.n59 VPB.n56 13.276
R127 VPB.n56 VPB.n53 13.276
R128 VPB.n53 VPB.n50 13.276
R129 VPB.n45 VPB.n16 13.276
R130 VPB.n67 VPB.n16 13.276
R131 VPB.n37 VPB.n19 13.276
R132 VPB.n19 VPB.n17 13.276
R133 VPB.n24 VPB.n22 12.796
R134 VPB.n24 VPB.n23 12.564
R135 VPB.n33 VPB.n32 12.198
R136 VPB.n30 VPB.n29 12.198
R137 VPB.n30 VPB.n27 12.198
R138 VPB.n50 VPB.n46 8.97
R139 VPB.n37 VPB.n36 7.5
R140 VPB.n22 VPB.n21 7.5
R141 VPB.n29 VPB.n28 7.5
R142 VPB.n27 VPB.n26 7.5
R143 VPB.n19 VPB.n18 7.5
R144 VPB.n34 VPB.n20 7.5
R145 VPB.n70 VPB.n69 7.5
R146 VPB.n12 VPB.n11 7.5
R147 VPB.n6 VPB.n5 7.5
R148 VPB.n8 VPB.n7 7.5
R149 VPB.n2 VPB.n1 7.5
R150 VPB.n72 VPB.n71 7.5
R151 VPB.n13 VPB.n10 6.729
R152 VPB.n9 VPB.n6 6.729
R153 VPB.n4 VPB.n2 6.729
R154 VPB.n4 VPB.n3 6.728
R155 VPB.n9 VPB.n8 6.728
R156 VPB.n13 VPB.n12 6.728
R157 VPB.n73 VPB.n72 6.728
R158 VPB.n36 VPB.n35 6.398
R159 VPB.n60 VPB.n40 6.112
R160 VPB.n60 VPB.n59 6.101
R161 VPB.n46 VPB.n45 4.305
R162 VPB.n34 VPB.n25 1.402
R163 VPB.n34 VPB.n30 1.402
R164 VPB.n34 VPB.n31 1.402
R165 VPB.n34 VPB.n33 1.402
R166 VPB.n35 VPB.n34 0.735
R167 VPB.n34 VPB.n24 0.735
R168 VPB.n74 VPB.n13 0.387
R169 VPB.n74 VPB.n9 0.387
R170 VPB.n74 VPB.n4 0.387
R171 VPB.n74 VPB.n73 0.387
R172 VPB.n66 VPB 0.198
R173 VPB.n62 VPB.n61 0.136
R174 VPB.n64 VPB.n63 0.136
R175 VPB.n65 VPB.n64 0.136
R176 VPB.n66 VPB.n65 0.136
R177 VPB VPB.n62 0.068
R178 VPB.n63 VPB 0.068














































































.ends
