* SPICE3 file created from FA.ext - technology: sky130A

.subckt FA SUM COUT A B CIN VDD GND
X0 a_836_182 a_807_943 a_575_1004 VDD pshort w=2 l=0.15 M=2
X1 a_1241_1004 a_185_182 a_836_182 VDD pshort w=2 l=0.15 M=2
X2 VDD a_5767_1004 a_6401_182 VDD pshort w=2 l=0.15 M=2
X3 a_2405_182 a_836_182 VDD VDD pshort w=2 l=0.15 M=2
X4 GND A a_556_74 GND nshort w=3 l=0.15
X5 VDD B a_807_943 VDD pshort w=2 l=0.15 M=2
X6 COUT a_6858_181 VDD VDD pshort w=2 l=0.15 M=2
X7 a_185_182 A GND GND nshort w=3 l=0.15
X8 VDD a_836_182 a_4657_1004 VDD pshort w=2 l=0.15 M=2
X9 VDD B a_5767_1004 VDD pshort w=2 l=0.15 M=2
X10 VDD A a_575_1004 VDD pshort w=2 l=0.15 M=2
X11 a_6401_182 a_5767_1004 GND GND nshort w=3 l=0.15
X12 a_4657_1004 CIN VDD VDD pshort w=2 l=0.15 M=2
X13 SUM a_2405_182 a_3461_1004 VDD pshort w=2 l=0.15 M=2
X14 a_3027_943 CIN VDD VDD pshort w=2 l=0.15 M=2
X15 VDD a_5291_182 a_6791_1005 VDD pshort w=2 l=0.15 M=2
X16 a_836_182 a_185_182 a_1222_74 GND nshort w=3 l=0.15
X17 VDD A a_185_182 VDD pshort w=2 l=0.15 M=2
X18 a_807_943 B GND GND nshort w=3 l=0.15
X19 a_2795_1004 a_3027_943 SUM VDD pshort w=2 l=0.15 M=2
X20 a_6791_1005 a_6401_182 a_6858_181 VDD pshort w=2 l=0.15 M=2
X21 GND a_3027_943 a_3442_74 GND nshort w=3 l=0.15
X22 VDD B a_1241_1004 VDD pshort w=2 l=0.15 M=2
X23 COUT a_6858_181 GND GND nshort w=3 l=0.15
X24 a_3461_1004 CIN VDD VDD pshort w=2 l=0.15 M=2
X25 a_5291_182 a_4657_1004 VDD VDD pshort w=2 l=0.15 M=2
X26 GND CIN a_4552_73 GND nshort w=3 l=0.15
X27 a_3027_943 CIN GND GND nshort w=3 l=0.15
X28 a_836_182 B a_556_74 GND nshort w=3 l=0.15
X29 VDD a_836_182 a_2795_1004 VDD pshort w=2 l=0.15 M=2
X30 VDD A a_5767_1004 VDD pshort w=2 l=0.15 M=2
X31 GND B a_5662_73 GND nshort w=3 l=0.15
X32 SUM a_2405_182 a_3442_74 GND nshort w=3 l=0.15
X33 a_4657_1004 a_836_182 a_4552_73 GND nshort w=3 l=0.15
X34 GND a_836_182 a_2776_74 GND nshort w=3 l=0.15
X35 a_2405_182 a_836_182 GND GND nshort w=3 l=0.15
X36 a_6858_181 a_5291_182 GND GND nshort w=3 l=0.15
X37 GND a_807_943 a_1222_74 GND nshort w=3 l=0.15
X38 a_6858_181 a_6401_182 GND GND nshort w=3 l=0.15
X39 SUM CIN a_2776_74 GND nshort w=3 l=0.15
X40 a_5291_182 a_4657_1004 GND GND nshort w=3 l=0.15
X41 a_5767_1004 A a_5662_73 GND nshort w=3 l=0.15
C0 a_836_182 a_807_943 2.38fF
C1 CIN a_3027_943 2.29fF
C2 A a_836_182 3.22fF
C3 B a_807_943 2.27fF
C4 VDD B 2.32fF
C5 VDD GND 18.70fF
C6 a_836_182 GND 2.30fF **FLOATING
.ends
