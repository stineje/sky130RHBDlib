* SPICE3 file created from DFFRNX1.ext - technology: sky130A

.subckt DFFRNX1 Q QN D CLK RN VDD GND
M1000 VDD.t22 RN.t0 a_147_187.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VDD.t1 a_147_187.t8 Q.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t6 a_147_187.t9 a_277_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 GND a_147_187.t10 a_91_103.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1004 QN Q.t6 a_3924_210.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1005 a_599_989.t1 D.t0 VDD.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VDD.t11 CLK.t0 a_277_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VDD.t8 a_599_989.t8 a_2141_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VDD.t15 a_277_1050.t7 QN.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_599_989.t6 RN.t2 VDD.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_147_187.t5 CLK.t1 VDD.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 QN.t2 Q.t5 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 GND a_277_1050.t8 a_3643_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1013 Q.t3 QN.t7 VDD.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t3 a_147_187.t11 a_2141_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VDD.t16 a_599_989.t9 a_277_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 VDD.t10 a_2141_1050.t5 a_147_187.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 GND QN.t8 a_4626_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1018 GND a_599_989.t10 a_2036_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1019 GND a_2141_1050.t6 a_2681_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_147_187.t2 RN.t3 VDD.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 Q.t1 a_147_187.t12 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_277_1050.t0 a_147_187.t13 VDD.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VDD.t31 a_277_1050.t9 a_599_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 GND a_277_1050.t11 a_1053_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1025 VDD.t24 RN.t5 a_599_989.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VDD.t13 Q.t7 QN.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_277_1050.t6 CLK.t3 VDD.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_2141_1050.t4 a_599_989.t11 VDD.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 QN.t3 a_277_1050.t10 VDD.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 VDD.t14 D.t1 a_599_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 VDD.t25 RN.t7 QN.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_599_989.t2 a_277_1050.t12 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 Q a_147_187.t15 a_4626_101.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1034 a_277_1050.t5 a_599_989.t12 VDD.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_2141_1050.t2 a_147_187.t14 VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_147_187.t4 a_2141_1050.t7 VDD.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 QN.t5 RN.t8 VDD.t26 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 VDD.t12 CLK.t5 a_147_187.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 VDD.t29 QN.t9 Q.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VDD QN 1.85fF
C1 VDD CLK 0.38fF
C2 RN Q 0.18fF
C3 D VDD 0.05fF
C4 RN QN 0.12fF
C5 RN VDD 0.17fF
C6 D CLK 0.07fF
C7 RN CLK 0.28fF
C8 D RN 0.18fF
C9 Q QN 0.93fF
C10 VDD Q 1.39fF
R0 a_147_187.n10 a_147_187.t9 512.525
R1 a_147_187.n8 a_147_187.t11 472.359
R2 a_147_187.n6 a_147_187.t8 472.359
R3 a_147_187.n8 a_147_187.t14 384.527
R4 a_147_187.n6 a_147_187.t12 384.527
R5 a_147_187.n10 a_147_187.t13 371.139
R6 a_147_187.n11 a_147_187.t10 340.774
R7 a_147_187.n9 a_147_187.t7 294.278
R8 a_147_187.n7 a_147_187.t15 294.278
R9 a_147_187.n16 a_147_187.n14 266.21
R10 a_147_187.n14 a_147_187.n5 117.693
R11 a_147_187.n11 a_147_187.n10 109.607
R12 a_147_187.n12 a_147_187.n11 83.572
R13 a_147_187.n13 a_147_187.n7 81.396
R14 a_147_187.n4 a_147_187.n3 79.232
R15 a_147_187.n12 a_147_187.n9 76
R16 a_147_187.n14 a_147_187.n13 76
R17 a_147_187.n5 a_147_187.n4 63.152
R18 a_147_187.n9 a_147_187.n8 56.954
R19 a_147_187.n7 a_147_187.n6 56.954
R20 a_147_187.n17 a_147_187.n0 55.263
R21 a_147_187.n16 a_147_187.n15 30
R22 a_147_187.n17 a_147_187.n16 23.684
R23 a_147_187.n5 a_147_187.n1 16.08
R24 a_147_187.n4 a_147_187.n2 16.08
R25 a_147_187.n1 a_147_187.t0 14.282
R26 a_147_187.n1 a_147_187.t2 14.282
R27 a_147_187.n2 a_147_187.t1 14.282
R28 a_147_187.n2 a_147_187.t5 14.282
R29 a_147_187.n3 a_147_187.t6 14.282
R30 a_147_187.n3 a_147_187.t4 14.282
R31 a_147_187.n13 a_147_187.n12 4.035
R32 a_2036_101.t0 a_2036_101.n1 34.62
R33 a_2036_101.t0 a_2036_101.n0 8.137
R34 a_2036_101.t0 a_2036_101.n2 4.69
R35 a_2141_1050.n3 a_2141_1050.t5 512.525
R36 a_2141_1050.n3 a_2141_1050.t7 371.139
R37 a_2141_1050.n4 a_2141_1050.t6 287.668
R38 a_2141_1050.n7 a_2141_1050.n5 217.114
R39 a_2141_1050.n4 a_2141_1050.n3 162.713
R40 a_2141_1050.n5 a_2141_1050.n4 153.315
R41 a_2141_1050.n5 a_2141_1050.n2 152.499
R42 a_2141_1050.n2 a_2141_1050.n1 76.002
R43 a_2141_1050.n7 a_2141_1050.n6 15.218
R44 a_2141_1050.n0 a_2141_1050.t0 14.282
R45 a_2141_1050.n0 a_2141_1050.t2 14.282
R46 a_2141_1050.n1 a_2141_1050.t3 14.282
R47 a_2141_1050.n1 a_2141_1050.t4 14.282
R48 a_2141_1050.n2 a_2141_1050.n0 12.85
R49 a_2141_1050.n8 a_2141_1050.n7 12.014
R50 RN.n0 RN.t7 479.223
R51 RN.n5 RN.t2 454.685
R52 RN.n2 RN.t3 454.685
R53 RN.n5 RN.t5 428.979
R54 RN.n2 RN.t0 428.979
R55 RN.n0 RN.t8 375.52
R56 RN.n6 RN.n5 178.106
R57 RN.n3 RN.n2 178.106
R58 RN.n1 RN.n0 175.429
R59 RN.n1 RN.t6 162.048
R60 RN.n6 RN.t4 158.3
R61 RN.n3 RN.t1 158.3
R62 RN.n4 RN.n1 78.675
R63 RN.n4 RN.n3 76
R64 RN.n7 RN.n6 76
R65 RN.n7 RN.n4 5.94
R66 RN.n7 RN 0.046
R67 VDD.n345 VDD.n343 144.705
R68 VDD.n462 VDD.n460 144.705
R69 VDD.n426 VDD.n424 144.705
R70 VDD.n164 VDD.n162 144.705
R71 VDD.n83 VDD.n81 144.705
R72 VDD.n44 VDD.n43 76
R73 VDD.n49 VDD.n48 76
R74 VDD.n54 VDD.n53 76
R75 VDD.n58 VDD.n57 76
R76 VDD.n85 VDD.n84 76
R77 VDD.n89 VDD.n88 76
R78 VDD.n93 VDD.n92 76
R79 VDD.n98 VDD.n97 76
R80 VDD.n105 VDD.n104 76
R81 VDD.n110 VDD.n109 76
R82 VDD.n115 VDD.n114 76
R83 VDD.n122 VDD.n121 76
R84 VDD.n127 VDD.n126 76
R85 VDD.n132 VDD.n131 76
R86 VDD.n136 VDD.n135 76
R87 VDD.n140 VDD.n139 76
R88 VDD.n166 VDD.n165 76
R89 VDD.n170 VDD.n169 76
R90 VDD.n174 VDD.n173 76
R91 VDD.n179 VDD.n178 76
R92 VDD.n186 VDD.n185 76
R93 VDD.n191 VDD.n190 76
R94 VDD.n196 VDD.n195 76
R95 VDD.n203 VDD.n202 76
R96 VDD.n208 VDD.n207 76
R97 VDD.n213 VDD.n212 76
R98 VDD.n217 VDD.n216 76
R99 VDD.n242 VDD.n241 76
R100 VDD.n464 VDD.n463 76
R101 VDD.n459 VDD.n458 76
R102 VDD.n454 VDD.n453 76
R103 VDD.n449 VDD.n448 76
R104 VDD.n443 VDD.n442 76
R105 VDD.n438 VDD.n437 76
R106 VDD.n433 VDD.n432 76
R107 VDD.n428 VDD.n427 76
R108 VDD.n402 VDD.n401 76
R109 VDD.n398 VDD.n397 76
R110 VDD.n394 VDD.n393 76
R111 VDD.n390 VDD.n389 76
R112 VDD.n385 VDD.n384 76
R113 VDD.n378 VDD.n377 76
R114 VDD.n373 VDD.n372 76
R115 VDD.n368 VDD.n367 76
R116 VDD.n361 VDD.n360 76
R117 VDD.n356 VDD.n355 76
R118 VDD.n351 VDD.n350 76
R119 VDD.n347 VDD.n346 76
R120 VDD.n320 VDD.n319 76
R121 VDD.n316 VDD.n315 76
R122 VDD.n312 VDD.n311 76
R123 VDD.n308 VDD.n307 76
R124 VDD.n303 VDD.n302 76
R125 VDD.n296 VDD.n295 76
R126 VDD.n291 VDD.n290 76
R127 VDD.n286 VDD.n285 76
R128 VDD.n279 VDD.n278 76
R129 VDD.n274 VDD.n273 76
R130 VDD.n269 VDD.n268 76
R131 VDD.n265 VDD.n264 76
R132 VDD.n95 VDD.n94 64.064
R133 VDD.n176 VDD.n175 64.064
R134 VDD.n387 VDD.n386 64.064
R135 VDD.n305 VDD.n304 64.064
R136 VDD.n124 VDD.n123 59.488
R137 VDD.n205 VDD.n204 59.488
R138 VDD.n358 VDD.n357 59.488
R139 VDD.n276 VDD.n275 59.488
R140 VDD.n270 VDD.t4 55.106
R141 VDD.n352 VDD.t0 55.106
R142 VDD.n429 VDD.t20 55.106
R143 VDD.n209 VDD.t9 55.106
R144 VDD.n128 VDD.t19 55.106
R145 VDD.n50 VDD.t7 55.106
R146 VDD.n311 VDD.t16 55.106
R147 VDD.n393 VDD.t24 55.106
R148 VDD.n173 VDD.t22 55.106
R149 VDD.n92 VDD.t13 55.106
R150 VDD.n455 VDD.t3 55.106
R151 VDD.n33 VDD.t1 55.106
R152 VDD.n281 VDD.n280 40.824
R153 VDD.n301 VDD.n300 40.824
R154 VDD.n363 VDD.n362 40.824
R155 VDD.n383 VDD.n382 40.824
R156 VDD.n445 VDD.n444 40.824
R157 VDD.n198 VDD.n197 40.824
R158 VDD.n184 VDD.n183 40.824
R159 VDD.n117 VDD.n116 40.824
R160 VDD.n103 VDD.n102 40.824
R161 VDD.n28 VDD.n27 40.824
R162 VDD.n407 VDD.n406 36.774
R163 VDD.n222 VDD.n221 36.774
R164 VDD.n145 VDD.n144 36.774
R165 VDD.n63 VDD.n62 36.774
R166 VDD.n336 VDD.n335 36.774
R167 VDD.n25 VDD.n24 36.608
R168 VDD.n451 VDD.n450 36.608
R169 VDD.n38 VDD.n37 34.942
R170 VDD.n46 VDD.n45 32.032
R171 VDD.n435 VDD.n434 32.032
R172 VDD.n100 VDD.n99 27.456
R173 VDD.n181 VDD.n180 27.456
R174 VDD.n380 VDD.n379 27.456
R175 VDD.n298 VDD.n297 27.456
R176 VDD.n119 VDD.n118 22.88
R177 VDD.n200 VDD.n199 22.88
R178 VDD.n365 VDD.n364 22.88
R179 VDD.n283 VDD.n282 22.88
R180 VDD.n264 VDD.n261 21.841
R181 VDD.n23 VDD.n20 21.841
R182 VDD.n280 VDD.t30 14.282
R183 VDD.n280 VDD.t6 14.282
R184 VDD.n300 VDD.t27 14.282
R185 VDD.n300 VDD.t11 14.282
R186 VDD.n362 VDD.t17 14.282
R187 VDD.n362 VDD.t31 14.282
R188 VDD.n382 VDD.t23 14.282
R189 VDD.n382 VDD.t14 14.282
R190 VDD.n444 VDD.t2 14.282
R191 VDD.n444 VDD.t8 14.282
R192 VDD.n197 VDD.t28 14.282
R193 VDD.n197 VDD.t10 14.282
R194 VDD.n183 VDD.t21 14.282
R195 VDD.n183 VDD.t12 14.282
R196 VDD.n116 VDD.t26 14.282
R197 VDD.n116 VDD.t15 14.282
R198 VDD.n102 VDD.t18 14.282
R199 VDD.n102 VDD.t25 14.282
R200 VDD.n27 VDD.t5 14.282
R201 VDD.n27 VDD.t29 14.282
R202 VDD.n261 VDD.n244 14.167
R203 VDD.n244 VDD.n243 14.167
R204 VDD.n422 VDD.n404 14.167
R205 VDD.n404 VDD.n403 14.167
R206 VDD.n237 VDD.n219 14.167
R207 VDD.n219 VDD.n218 14.167
R208 VDD.n160 VDD.n142 14.167
R209 VDD.n142 VDD.n141 14.167
R210 VDD.n79 VDD.n60 14.167
R211 VDD.n60 VDD.n59 14.167
R212 VDD.n341 VDD.n322 14.167
R213 VDD.n322 VDD.n321 14.167
R214 VDD.n20 VDD.n19 14.167
R215 VDD.n19 VDD.n17 14.167
R216 VDD.n32 VDD.n31 14.167
R217 VDD.n84 VDD.n80 14.167
R218 VDD.n165 VDD.n161 14.167
R219 VDD.n241 VDD.n238 14.167
R220 VDD.n427 VDD.n423 14.167
R221 VDD.n346 VDD.n342 14.167
R222 VDD.n112 VDD.n111 13.728
R223 VDD.n193 VDD.n192 13.728
R224 VDD.n370 VDD.n369 13.728
R225 VDD.n288 VDD.n287 13.728
R226 VDD.n23 VDD.n22 13.653
R227 VDD.n22 VDD.n21 13.653
R228 VDD.n36 VDD.n35 13.653
R229 VDD.n35 VDD.n34 13.653
R230 VDD.n32 VDD.n26 13.653
R231 VDD.n26 VDD.n25 13.653
R232 VDD.n31 VDD.n30 13.653
R233 VDD.n30 VDD.n29 13.653
R234 VDD.n43 VDD.n42 13.653
R235 VDD.n42 VDD.n41 13.653
R236 VDD.n48 VDD.n47 13.653
R237 VDD.n47 VDD.n46 13.653
R238 VDD.n53 VDD.n52 13.653
R239 VDD.n52 VDD.n51 13.653
R240 VDD.n57 VDD.n56 13.653
R241 VDD.n56 VDD.n55 13.653
R242 VDD.n84 VDD.n83 13.653
R243 VDD.n83 VDD.n82 13.653
R244 VDD.n88 VDD.n87 13.653
R245 VDD.n87 VDD.n86 13.653
R246 VDD.n92 VDD.n91 13.653
R247 VDD.n91 VDD.n90 13.653
R248 VDD.n97 VDD.n96 13.653
R249 VDD.n96 VDD.n95 13.653
R250 VDD.n104 VDD.n101 13.653
R251 VDD.n101 VDD.n100 13.653
R252 VDD.n109 VDD.n108 13.653
R253 VDD.n108 VDD.n107 13.653
R254 VDD.n114 VDD.n113 13.653
R255 VDD.n113 VDD.n112 13.653
R256 VDD.n121 VDD.n120 13.653
R257 VDD.n120 VDD.n119 13.653
R258 VDD.n126 VDD.n125 13.653
R259 VDD.n125 VDD.n124 13.653
R260 VDD.n131 VDD.n130 13.653
R261 VDD.n130 VDD.n129 13.653
R262 VDD.n135 VDD.n134 13.653
R263 VDD.n134 VDD.n133 13.653
R264 VDD.n139 VDD.n138 13.653
R265 VDD.n138 VDD.n137 13.653
R266 VDD.n165 VDD.n164 13.653
R267 VDD.n164 VDD.n163 13.653
R268 VDD.n169 VDD.n168 13.653
R269 VDD.n168 VDD.n167 13.653
R270 VDD.n173 VDD.n172 13.653
R271 VDD.n172 VDD.n171 13.653
R272 VDD.n178 VDD.n177 13.653
R273 VDD.n177 VDD.n176 13.653
R274 VDD.n185 VDD.n182 13.653
R275 VDD.n182 VDD.n181 13.653
R276 VDD.n190 VDD.n189 13.653
R277 VDD.n189 VDD.n188 13.653
R278 VDD.n195 VDD.n194 13.653
R279 VDD.n194 VDD.n193 13.653
R280 VDD.n202 VDD.n201 13.653
R281 VDD.n201 VDD.n200 13.653
R282 VDD.n207 VDD.n206 13.653
R283 VDD.n206 VDD.n205 13.653
R284 VDD.n212 VDD.n211 13.653
R285 VDD.n211 VDD.n210 13.653
R286 VDD.n216 VDD.n215 13.653
R287 VDD.n215 VDD.n214 13.653
R288 VDD.n241 VDD.n240 13.653
R289 VDD.n240 VDD.n239 13.653
R290 VDD.n463 VDD.n462 13.653
R291 VDD.n462 VDD.n461 13.653
R292 VDD.n458 VDD.n457 13.653
R293 VDD.n457 VDD.n456 13.653
R294 VDD.n453 VDD.n452 13.653
R295 VDD.n452 VDD.n451 13.653
R296 VDD.n448 VDD.n447 13.653
R297 VDD.n447 VDD.n446 13.653
R298 VDD.n442 VDD.n441 13.653
R299 VDD.n441 VDD.n440 13.653
R300 VDD.n437 VDD.n436 13.653
R301 VDD.n436 VDD.n435 13.653
R302 VDD.n432 VDD.n431 13.653
R303 VDD.n431 VDD.n430 13.653
R304 VDD.n427 VDD.n426 13.653
R305 VDD.n426 VDD.n425 13.653
R306 VDD.n401 VDD.n400 13.653
R307 VDD.n400 VDD.n399 13.653
R308 VDD.n397 VDD.n396 13.653
R309 VDD.n396 VDD.n395 13.653
R310 VDD.n393 VDD.n392 13.653
R311 VDD.n392 VDD.n391 13.653
R312 VDD.n389 VDD.n388 13.653
R313 VDD.n388 VDD.n387 13.653
R314 VDD.n384 VDD.n381 13.653
R315 VDD.n381 VDD.n380 13.653
R316 VDD.n377 VDD.n376 13.653
R317 VDD.n376 VDD.n375 13.653
R318 VDD.n372 VDD.n371 13.653
R319 VDD.n371 VDD.n370 13.653
R320 VDD.n367 VDD.n366 13.653
R321 VDD.n366 VDD.n365 13.653
R322 VDD.n360 VDD.n359 13.653
R323 VDD.n359 VDD.n358 13.653
R324 VDD.n355 VDD.n354 13.653
R325 VDD.n354 VDD.n353 13.653
R326 VDD.n350 VDD.n349 13.653
R327 VDD.n349 VDD.n348 13.653
R328 VDD.n346 VDD.n345 13.653
R329 VDD.n345 VDD.n344 13.653
R330 VDD.n319 VDD.n318 13.653
R331 VDD.n318 VDD.n317 13.653
R332 VDD.n315 VDD.n314 13.653
R333 VDD.n314 VDD.n313 13.653
R334 VDD.n311 VDD.n310 13.653
R335 VDD.n310 VDD.n309 13.653
R336 VDD.n307 VDD.n306 13.653
R337 VDD.n306 VDD.n305 13.653
R338 VDD.n302 VDD.n299 13.653
R339 VDD.n299 VDD.n298 13.653
R340 VDD.n295 VDD.n294 13.653
R341 VDD.n294 VDD.n293 13.653
R342 VDD.n290 VDD.n289 13.653
R343 VDD.n289 VDD.n288 13.653
R344 VDD.n285 VDD.n284 13.653
R345 VDD.n284 VDD.n283 13.653
R346 VDD.n278 VDD.n277 13.653
R347 VDD.n277 VDD.n276 13.653
R348 VDD.n273 VDD.n272 13.653
R349 VDD.n272 VDD.n271 13.653
R350 VDD.n268 VDD.n267 13.653
R351 VDD.n267 VDD.n266 13.653
R352 VDD.n264 VDD.n263 13.653
R353 VDD.n263 VDD.n262 13.653
R354 VDD.n4 VDD.n2 12.915
R355 VDD.n4 VDD.n3 12.66
R356 VDD.n10 VDD.n9 12.343
R357 VDD.n12 VDD.n11 12.343
R358 VDD.n10 VDD.n7 12.343
R359 VDD.n33 VDD.n32 11.806
R360 VDD.n107 VDD.n106 9.152
R361 VDD.n188 VDD.n187 9.152
R362 VDD.n375 VDD.n374 9.152
R363 VDD.n293 VDD.n292 9.152
R364 VDD.n31 VDD.n28 8.658
R365 VDD.n448 VDD.n445 8.658
R366 VDD.n423 VDD.n422 7.674
R367 VDD.n238 VDD.n237 7.674
R368 VDD.n161 VDD.n160 7.674
R369 VDD.n80 VDD.n79 7.674
R370 VDD.n342 VDD.n341 7.674
R371 VDD.n74 VDD.n73 7.5
R372 VDD.n68 VDD.n67 7.5
R373 VDD.n70 VDD.n69 7.5
R374 VDD.n65 VDD.n64 7.5
R375 VDD.n79 VDD.n78 7.5
R376 VDD.n155 VDD.n154 7.5
R377 VDD.n149 VDD.n148 7.5
R378 VDD.n151 VDD.n150 7.5
R379 VDD.n157 VDD.n147 7.5
R380 VDD.n157 VDD.n145 7.5
R381 VDD.n160 VDD.n159 7.5
R382 VDD.n232 VDD.n231 7.5
R383 VDD.n226 VDD.n225 7.5
R384 VDD.n228 VDD.n227 7.5
R385 VDD.n234 VDD.n224 7.5
R386 VDD.n234 VDD.n222 7.5
R387 VDD.n237 VDD.n236 7.5
R388 VDD.n417 VDD.n416 7.5
R389 VDD.n411 VDD.n410 7.5
R390 VDD.n413 VDD.n412 7.5
R391 VDD.n419 VDD.n409 7.5
R392 VDD.n419 VDD.n407 7.5
R393 VDD.n422 VDD.n421 7.5
R394 VDD.n326 VDD.n325 7.5
R395 VDD.n329 VDD.n328 7.5
R396 VDD.n331 VDD.n330 7.5
R397 VDD.n334 VDD.n333 7.5
R398 VDD.n341 VDD.n340 7.5
R399 VDD.n256 VDD.n255 7.5
R400 VDD.n250 VDD.n249 7.5
R401 VDD.n252 VDD.n251 7.5
R402 VDD.n258 VDD.n248 7.5
R403 VDD.n258 VDD.n246 7.5
R404 VDD.n261 VDD.n260 7.5
R405 VDD.n20 VDD.n16 7.5
R406 VDD.n2 VDD.n1 7.5
R407 VDD.n9 VDD.n8 7.5
R408 VDD.n7 VDD.n6 7.5
R409 VDD.n19 VDD.n18 7.5
R410 VDD.n14 VDD.n0 7.5
R411 VDD.n66 VDD.n63 6.772
R412 VDD.n77 VDD.n61 6.772
R413 VDD.n75 VDD.n72 6.772
R414 VDD.n71 VDD.n68 6.772
R415 VDD.n158 VDD.n143 6.772
R416 VDD.n156 VDD.n153 6.772
R417 VDD.n152 VDD.n149 6.772
R418 VDD.n235 VDD.n220 6.772
R419 VDD.n233 VDD.n230 6.772
R420 VDD.n229 VDD.n226 6.772
R421 VDD.n420 VDD.n405 6.772
R422 VDD.n418 VDD.n415 6.772
R423 VDD.n414 VDD.n411 6.772
R424 VDD.n259 VDD.n245 6.772
R425 VDD.n257 VDD.n254 6.772
R426 VDD.n253 VDD.n250 6.772
R427 VDD.n66 VDD.n65 6.772
R428 VDD.n71 VDD.n70 6.772
R429 VDD.n75 VDD.n74 6.772
R430 VDD.n78 VDD.n77 6.772
R431 VDD.n152 VDD.n151 6.772
R432 VDD.n156 VDD.n155 6.772
R433 VDD.n159 VDD.n158 6.772
R434 VDD.n229 VDD.n228 6.772
R435 VDD.n233 VDD.n232 6.772
R436 VDD.n236 VDD.n235 6.772
R437 VDD.n414 VDD.n413 6.772
R438 VDD.n418 VDD.n417 6.772
R439 VDD.n421 VDD.n420 6.772
R440 VDD.n253 VDD.n252 6.772
R441 VDD.n257 VDD.n256 6.772
R442 VDD.n260 VDD.n259 6.772
R443 VDD.n340 VDD.n339 6.772
R444 VDD.n327 VDD.n324 6.772
R445 VDD.n332 VDD.n329 6.772
R446 VDD.n337 VDD.n334 6.772
R447 VDD.n337 VDD.n336 6.772
R448 VDD.n332 VDD.n331 6.772
R449 VDD.n327 VDD.n326 6.772
R450 VDD.n339 VDD.n323 6.772
R451 VDD.n121 VDD.n117 6.69
R452 VDD.n202 VDD.n198 6.69
R453 VDD.n367 VDD.n363 6.69
R454 VDD.n285 VDD.n281 6.69
R455 VDD.n37 VDD.n23 6.487
R456 VDD.n37 VDD.n36 6.475
R457 VDD.n16 VDD.n15 6.458
R458 VDD.n104 VDD.n103 6.296
R459 VDD.n185 VDD.n184 6.296
R460 VDD.n384 VDD.n383 6.296
R461 VDD.n302 VDD.n301 6.296
R462 VDD.n147 VDD.n146 6.202
R463 VDD.n224 VDD.n223 6.202
R464 VDD.n409 VDD.n408 6.202
R465 VDD.n248 VDD.n247 6.202
R466 VDD.n41 VDD.n40 4.576
R467 VDD.n440 VDD.n439 4.576
R468 VDD.n53 VDD.n50 2.754
R469 VDD.n432 VDD.n429 2.754
R470 VDD.n36 VDD.n33 2.361
R471 VDD.n458 VDD.n455 2.361
R472 VDD.n14 VDD.n5 1.329
R473 VDD.n14 VDD.n10 1.329
R474 VDD.n14 VDD.n12 1.329
R475 VDD.n14 VDD.n13 1.329
R476 VDD.n15 VDD.n14 0.696
R477 VDD.n14 VDD.n4 0.696
R478 VDD.n131 VDD.n128 0.393
R479 VDD.n212 VDD.n209 0.393
R480 VDD.n355 VDD.n352 0.393
R481 VDD.n273 VDD.n270 0.393
R482 VDD.n76 VDD.n75 0.365
R483 VDD.n76 VDD.n71 0.365
R484 VDD.n76 VDD.n66 0.365
R485 VDD.n77 VDD.n76 0.365
R486 VDD.n157 VDD.n156 0.365
R487 VDD.n157 VDD.n152 0.365
R488 VDD.n158 VDD.n157 0.365
R489 VDD.n234 VDD.n233 0.365
R490 VDD.n234 VDD.n229 0.365
R491 VDD.n235 VDD.n234 0.365
R492 VDD.n419 VDD.n418 0.365
R493 VDD.n419 VDD.n414 0.365
R494 VDD.n420 VDD.n419 0.365
R495 VDD.n258 VDD.n257 0.365
R496 VDD.n258 VDD.n253 0.365
R497 VDD.n259 VDD.n258 0.365
R498 VDD.n338 VDD.n337 0.365
R499 VDD.n338 VDD.n332 0.365
R500 VDD.n338 VDD.n327 0.365
R501 VDD.n339 VDD.n338 0.365
R502 VDD.n85 VDD.n58 0.29
R503 VDD.n166 VDD.n140 0.29
R504 VDD.n428 VDD.n402 0.29
R505 VDD.n347 VDD.n320 0.29
R506 VDD.n265 VDD 0.207
R507 VDD.n115 VDD.n110 0.197
R508 VDD.n196 VDD.n191 0.197
R509 VDD.n378 VDD.n373 0.197
R510 VDD.n296 VDD.n291 0.197
R511 VDD.n44 VDD.n39 0.181
R512 VDD.n449 VDD.n443 0.181
R513 VDD.n39 VDD.n38 0.145
R514 VDD.n49 VDD.n44 0.145
R515 VDD.n54 VDD.n49 0.145
R516 VDD.n58 VDD.n54 0.145
R517 VDD.n89 VDD.n85 0.145
R518 VDD.n93 VDD.n89 0.145
R519 VDD.n98 VDD.n93 0.145
R520 VDD.n105 VDD.n98 0.145
R521 VDD.n110 VDD.n105 0.145
R522 VDD.n122 VDD.n115 0.145
R523 VDD.n127 VDD.n122 0.145
R524 VDD.n132 VDD.n127 0.145
R525 VDD.n136 VDD.n132 0.145
R526 VDD.n140 VDD.n136 0.145
R527 VDD.n170 VDD.n166 0.145
R528 VDD.n174 VDD.n170 0.145
R529 VDD.n179 VDD.n174 0.145
R530 VDD.n186 VDD.n179 0.145
R531 VDD.n191 VDD.n186 0.145
R532 VDD.n203 VDD.n196 0.145
R533 VDD.n208 VDD.n203 0.145
R534 VDD.n213 VDD.n208 0.145
R535 VDD.n217 VDD.n213 0.145
R536 VDD.n242 VDD.n217 0.145
R537 VDD VDD.n242 0.145
R538 VDD VDD.n464 0.145
R539 VDD.n464 VDD.n459 0.145
R540 VDD.n459 VDD.n454 0.145
R541 VDD.n454 VDD.n449 0.145
R542 VDD.n443 VDD.n438 0.145
R543 VDD.n438 VDD.n433 0.145
R544 VDD.n433 VDD.n428 0.145
R545 VDD.n402 VDD.n398 0.145
R546 VDD.n398 VDD.n394 0.145
R547 VDD.n394 VDD.n390 0.145
R548 VDD.n390 VDD.n385 0.145
R549 VDD.n385 VDD.n378 0.145
R550 VDD.n373 VDD.n368 0.145
R551 VDD.n368 VDD.n361 0.145
R552 VDD.n361 VDD.n356 0.145
R553 VDD.n356 VDD.n351 0.145
R554 VDD.n351 VDD.n347 0.145
R555 VDD.n320 VDD.n316 0.145
R556 VDD.n316 VDD.n312 0.145
R557 VDD.n312 VDD.n308 0.145
R558 VDD.n308 VDD.n303 0.145
R559 VDD.n303 VDD.n296 0.145
R560 VDD.n291 VDD.n286 0.145
R561 VDD.n286 VDD.n279 0.145
R562 VDD.n279 VDD.n274 0.145
R563 VDD.n274 VDD.n269 0.145
R564 VDD.n269 VDD.n265 0.145
R565 Q.n8 Q.t5 454.685
R566 Q.n8 Q.t7 428.979
R567 Q.n9 Q.t6 264.512
R568 Q.n7 Q.n6 237.145
R569 Q.n7 Q.n2 125.947
R570 Q Q.n9 78.901
R571 Q.n2 Q.n1 76.002
R572 Q.n10 Q.n7 76
R573 Q.n9 Q.n8 71.894
R574 Q.n6 Q.n5 30
R575 Q.n4 Q.n3 24.383
R576 Q.n6 Q.n4 23.684
R577 Q.n0 Q.t2 14.282
R578 Q.n0 Q.t1 14.282
R579 Q.n1 Q.t4 14.282
R580 Q.n1 Q.t3 14.282
R581 Q.n2 Q.n0 12.85
R582 Q.n10 Q 0.046
R583 a_277_1050.n4 a_277_1050.t9 512.525
R584 a_277_1050.n2 a_277_1050.t7 512.525
R585 a_277_1050.n4 a_277_1050.t12 371.139
R586 a_277_1050.n2 a_277_1050.t10 371.139
R587 a_277_1050.n5 a_277_1050.t11 314.221
R588 a_277_1050.n3 a_277_1050.t8 314.221
R589 a_277_1050.n8 a_277_1050.n7 261.396
R590 a_277_1050.n9 a_277_1050.n8 144.246
R591 a_277_1050.n5 a_277_1050.n4 136.16
R592 a_277_1050.n3 a_277_1050.n2 136.16
R593 a_277_1050.n6 a_277_1050.n3 85.476
R594 a_277_1050.n11 a_277_1050.n10 79.231
R595 a_277_1050.n8 a_277_1050.n6 77.315
R596 a_277_1050.n6 a_277_1050.n5 76
R597 a_277_1050.n10 a_277_1050.n9 63.152
R598 a_277_1050.n9 a_277_1050.n1 16.08
R599 a_277_1050.n10 a_277_1050.n0 16.08
R600 a_277_1050.n1 a_277_1050.t3 14.282
R601 a_277_1050.n1 a_277_1050.t5 14.282
R602 a_277_1050.n0 a_277_1050.t2 14.282
R603 a_277_1050.n0 a_277_1050.t6 14.282
R604 a_277_1050.t1 a_277_1050.n11 14.282
R605 a_277_1050.n11 a_277_1050.t0 14.282
R606 a_599_989.n2 a_599_989.t8 480.392
R607 a_599_989.n4 a_599_989.t12 454.685
R608 a_599_989.n4 a_599_989.t9 428.979
R609 a_599_989.n2 a_599_989.t11 403.272
R610 a_599_989.n3 a_599_989.t10 283.48
R611 a_599_989.n5 a_599_989.t7 237.959
R612 a_599_989.n11 a_599_989.n10 213.104
R613 a_599_989.n12 a_599_989.n11 170.799
R614 a_599_989.n5 a_599_989.n4 98.447
R615 a_599_989.n3 a_599_989.n2 98.447
R616 a_599_989.n6 a_599_989.n5 80.035
R617 a_599_989.n14 a_599_989.n13 79.231
R618 a_599_989.n6 a_599_989.n3 77.315
R619 a_599_989.n11 a_599_989.n6 76
R620 a_599_989.n13 a_599_989.n12 63.152
R621 a_599_989.n10 a_599_989.n9 30
R622 a_599_989.n8 a_599_989.n7 24.383
R623 a_599_989.n10 a_599_989.n8 23.684
R624 a_599_989.n12 a_599_989.n1 16.08
R625 a_599_989.n13 a_599_989.n0 16.08
R626 a_599_989.n1 a_599_989.t5 14.282
R627 a_599_989.n1 a_599_989.t6 14.282
R628 a_599_989.n0 a_599_989.t0 14.282
R629 a_599_989.n0 a_599_989.t1 14.282
R630 a_599_989.t3 a_599_989.n14 14.282
R631 a_599_989.n14 a_599_989.t2 14.282
R632 a_372_210.n8 a_372_210.n6 96.467
R633 a_372_210.n3 a_372_210.n1 44.628
R634 a_372_210.t0 a_372_210.n8 32.417
R635 a_372_210.n3 a_372_210.n2 23.284
R636 a_372_210.n6 a_372_210.n5 22.349
R637 a_372_210.t0 a_372_210.n10 20.241
R638 a_372_210.n10 a_372_210.n9 13.494
R639 a_372_210.n6 a_372_210.n4 8.443
R640 a_372_210.t0 a_372_210.n0 8.137
R641 a_372_210.t0 a_372_210.n3 5.727
R642 a_372_210.n8 a_372_210.n7 1.435
R643 D.n0 D.t1 479.223
R644 D.n0 D.t0 375.52
R645 D.n1 D.t2 215.154
R646 D.n1 D.n0 122.323
R647 D.n2 D.n1 76
R648 D.n2 D 0.046
R649 a_2962_210.n10 a_2962_210.n8 82.852
R650 a_2962_210.n11 a_2962_210.n0 49.6
R651 a_2962_210.n7 a_2962_210.n6 32.833
R652 a_2962_210.n8 a_2962_210.t1 32.416
R653 a_2962_210.n10 a_2962_210.n9 27.2
R654 a_2962_210.n3 a_2962_210.n2 23.284
R655 a_2962_210.n11 a_2962_210.n10 22.4
R656 a_2962_210.n7 a_2962_210.n4 19.017
R657 a_2962_210.n6 a_2962_210.n5 13.494
R658 a_2962_210.t1 a_2962_210.n1 7.04
R659 a_2962_210.t1 a_2962_210.n3 5.727
R660 a_2962_210.n8 a_2962_210.n7 1.435
R661 CLK.n2 CLK.t0 459.505
R662 CLK.n0 CLK.t5 459.505
R663 CLK.n2 CLK.t3 384.527
R664 CLK.n0 CLK.t1 384.527
R665 CLK.n3 CLK.t2 322.152
R666 CLK.n1 CLK.t4 322.151
R667 CLK.n4 CLK.n1 58.818
R668 CLK.n4 CLK.n3 49.342
R669 CLK.n3 CLK.n2 27.599
R670 CLK.n1 CLK.n0 27.599
R671 CLK.n4 CLK 0.046
R672 QN.n0 QN.t9 480.392
R673 QN.n0 QN.t7 403.272
R674 QN.n1 QN.t8 283.48
R675 QN.n11 QN.n10 213.104
R676 QN.n11 QN.n6 170.799
R677 QN.n1 QN.n0 98.447
R678 QN.n5 QN.n4 79.232
R679 QN.n12 QN.n1 77.315
R680 QN.n12 QN.n11 76
R681 QN.n6 QN.n5 63.152
R682 QN.n10 QN.n9 30
R683 QN.n8 QN.n7 24.383
R684 QN.n10 QN.n8 23.684
R685 QN.n6 QN.n2 16.08
R686 QN.n5 QN.n3 16.08
R687 QN.n2 QN.t1 14.282
R688 QN.n2 QN.t2 14.282
R689 QN.n3 QN.t6 14.282
R690 QN.n3 QN.t5 14.282
R691 QN.n4 QN.t4 14.282
R692 QN.n4 QN.t3 14.282
R693 QN.n12 QN 0.046
R694 a_91_103.t0 a_91_103.n3 117.777
R695 a_91_103.n6 a_91_103.n5 45.444
R696 a_91_103.t0 a_91_103.n6 21.213
R697 a_91_103.t0 a_91_103.n4 11.595
R698 a_91_103.n2 a_91_103.n1 2.455
R699 a_91_103.n2 a_91_103.n0 1.32
R700 a_91_103.t0 a_91_103.n2 0.246
R701 GND.n29 GND.n27 219.745
R702 GND.n158 GND.n157 219.745
R703 GND.n203 GND.n201 219.745
R704 GND.n229 GND.n227 219.745
R705 GND.n74 GND.n73 219.745
R706 GND.n125 GND.n124 85.559
R707 GND.n29 GND.n28 85.529
R708 GND.n158 GND.n156 85.529
R709 GND.n203 GND.n202 85.529
R710 GND.n229 GND.n228 85.529
R711 GND.n74 GND.n72 85.529
R712 GND.n211 GND.n210 84.842
R713 GND.n119 GND.n118 76
R714 GND.n12 GND.n11 76
R715 GND.n20 GND.n19 76
R716 GND.n23 GND.n22 76
R717 GND.n26 GND.n25 76
R718 GND.n33 GND.n32 76
R719 GND.n36 GND.n35 76
R720 GND.n39 GND.n38 76
R721 GND.n42 GND.n41 76
R722 GND.n45 GND.n44 76
R723 GND.n48 GND.n47 76
R724 GND.n51 GND.n50 76
R725 GND.n54 GND.n53 76
R726 GND.n57 GND.n56 76
R727 GND.n65 GND.n64 76
R728 GND.n68 GND.n67 76
R729 GND.n71 GND.n70 76
R730 GND.n78 GND.n77 76
R731 GND.n81 GND.n80 76
R732 GND.n84 GND.n83 76
R733 GND.n87 GND.n86 76
R734 GND.n90 GND.n89 76
R735 GND.n93 GND.n92 76
R736 GND.n96 GND.n95 76
R737 GND.n99 GND.n98 76
R738 GND.n102 GND.n101 76
R739 GND.n110 GND.n109 76
R740 GND.n113 GND.n112 76
R741 GND.n116 GND.n115 76
R742 GND.n233 GND.n232 76
R743 GND.n226 GND.n225 76
R744 GND.n223 GND.n222 76
R745 GND.n220 GND.n219 76
R746 GND.n217 GND.n216 76
R747 GND.n214 GND.n213 76
R748 GND.n209 GND.n208 76
R749 GND.n206 GND.n205 76
R750 GND.n199 GND.n198 76
R751 GND.n196 GND.n195 76
R752 GND.n193 GND.n192 76
R753 GND.n190 GND.n189 76
R754 GND.n187 GND.n186 76
R755 GND.n184 GND.n183 76
R756 GND.n181 GND.n180 76
R757 GND.n178 GND.n177 76
R758 GND.n175 GND.n174 76
R759 GND.n172 GND.n171 76
R760 GND.n164 GND.n163 76
R761 GND.n161 GND.n160 76
R762 GND.n154 GND.n153 76
R763 GND.n151 GND.n150 76
R764 GND.n148 GND.n147 76
R765 GND.n145 GND.n144 76
R766 GND.n142 GND.n141 76
R767 GND.n139 GND.n138 76
R768 GND.n136 GND.n135 76
R769 GND.n133 GND.n132 76
R770 GND.n130 GND.n129 76
R771 GND.n127 GND.n126 76
R772 GND.n122 GND.n121 76
R773 GND.n63 GND.n62 64.552
R774 GND.n108 GND.n107 64.552
R775 GND.n170 GND.n169 64.552
R776 GND.n17 GND.n16 63.835
R777 GND.n8 GND.n7 34.942
R778 GND.n16 GND.n15 28.421
R779 GND.n62 GND.n61 28.421
R780 GND.n107 GND.n106 28.421
R781 GND.n169 GND.n168 28.421
R782 GND.n16 GND.n14 25.263
R783 GND.n62 GND.n60 25.263
R784 GND.n107 GND.n105 25.263
R785 GND.n169 GND.n167 25.263
R786 GND.n14 GND.n13 24.383
R787 GND.n60 GND.n59 24.383
R788 GND.n105 GND.n104 24.383
R789 GND.n167 GND.n166 24.383
R790 GND.n6 GND.n5 14.167
R791 GND.n5 GND.n4 14.167
R792 GND.n32 GND.n30 14.167
R793 GND.n77 GND.n75 14.167
R794 GND.n232 GND.n230 14.167
R795 GND.n205 GND.n204 14.167
R796 GND.n160 GND.n159 14.167
R797 GND.n121 GND.n120 13.653
R798 GND.n126 GND.n123 13.653
R799 GND.n129 GND.n128 13.653
R800 GND.n132 GND.n131 13.653
R801 GND.n135 GND.n134 13.653
R802 GND.n138 GND.n137 13.653
R803 GND.n141 GND.n140 13.653
R804 GND.n144 GND.n143 13.653
R805 GND.n147 GND.n146 13.653
R806 GND.n150 GND.n149 13.653
R807 GND.n153 GND.n152 13.653
R808 GND.n160 GND.n155 13.653
R809 GND.n163 GND.n162 13.653
R810 GND.n171 GND.n165 13.653
R811 GND.n174 GND.n173 13.653
R812 GND.n177 GND.n176 13.653
R813 GND.n180 GND.n179 13.653
R814 GND.n183 GND.n182 13.653
R815 GND.n186 GND.n185 13.653
R816 GND.n189 GND.n188 13.653
R817 GND.n192 GND.n191 13.653
R818 GND.n195 GND.n194 13.653
R819 GND.n198 GND.n197 13.653
R820 GND.n205 GND.n200 13.653
R821 GND.n208 GND.n207 13.653
R822 GND.n213 GND.n212 13.653
R823 GND.n216 GND.n215 13.653
R824 GND.n219 GND.n218 13.653
R825 GND.n222 GND.n221 13.653
R826 GND.n225 GND.n224 13.653
R827 GND.n232 GND.n231 13.653
R828 GND.n115 GND.n114 13.653
R829 GND.n112 GND.n111 13.653
R830 GND.n109 GND.n103 13.653
R831 GND.n101 GND.n100 13.653
R832 GND.n98 GND.n97 13.653
R833 GND.n95 GND.n94 13.653
R834 GND.n92 GND.n91 13.653
R835 GND.n89 GND.n88 13.653
R836 GND.n86 GND.n85 13.653
R837 GND.n83 GND.n82 13.653
R838 GND.n80 GND.n79 13.653
R839 GND.n77 GND.n76 13.653
R840 GND.n70 GND.n69 13.653
R841 GND.n67 GND.n66 13.653
R842 GND.n64 GND.n58 13.653
R843 GND.n56 GND.n55 13.653
R844 GND.n53 GND.n52 13.653
R845 GND.n50 GND.n49 13.653
R846 GND.n47 GND.n46 13.653
R847 GND.n44 GND.n43 13.653
R848 GND.n41 GND.n40 13.653
R849 GND.n38 GND.n37 13.653
R850 GND.n35 GND.n34 13.653
R851 GND.n32 GND.n31 13.653
R852 GND.n25 GND.n24 13.653
R853 GND.n22 GND.n21 13.653
R854 GND.n19 GND.n18 13.653
R855 GND.n11 GND.n10 13.653
R856 GND.n4 GND.n3 13.653
R857 GND.n5 GND.n2 13.653
R858 GND.n6 GND.n1 13.653
R859 GND.n30 GND.n29 7.312
R860 GND.n159 GND.n158 7.312
R861 GND.n204 GND.n203 7.312
R862 GND.n230 GND.n229 7.312
R863 GND.n75 GND.n74 7.312
R864 GND.n7 GND.n0 7.083
R865 GND.n7 GND.n6 6.474
R866 GND.n19 GND.n17 3.935
R867 GND.n213 GND.n211 3.935
R868 GND.n118 GND.n117 0.596
R869 GND.n33 GND.n26 0.29
R870 GND.n78 GND.n71 0.29
R871 GND.n206 GND.n199 0.29
R872 GND.n161 GND.n154 0.29
R873 GND.n119 GND 0.207
R874 GND.n51 GND.n48 0.197
R875 GND.n96 GND.n93 0.197
R876 GND.n184 GND.n181 0.197
R877 GND.n139 GND.n136 0.197
R878 GND.n64 GND.n63 0.196
R879 GND.n109 GND.n108 0.196
R880 GND.n171 GND.n170 0.196
R881 GND.n126 GND.n125 0.196
R882 GND.n12 GND.n9 0.181
R883 GND.n220 GND.n217 0.181
R884 GND.n9 GND.n8 0.145
R885 GND.n20 GND.n12 0.145
R886 GND.n23 GND.n20 0.145
R887 GND.n26 GND.n23 0.145
R888 GND.n36 GND.n33 0.145
R889 GND.n39 GND.n36 0.145
R890 GND.n42 GND.n39 0.145
R891 GND.n45 GND.n42 0.145
R892 GND.n48 GND.n45 0.145
R893 GND.n54 GND.n51 0.145
R894 GND.n57 GND.n54 0.145
R895 GND.n65 GND.n57 0.145
R896 GND.n68 GND.n65 0.145
R897 GND.n71 GND.n68 0.145
R898 GND.n81 GND.n78 0.145
R899 GND.n84 GND.n81 0.145
R900 GND.n87 GND.n84 0.145
R901 GND.n90 GND.n87 0.145
R902 GND.n93 GND.n90 0.145
R903 GND.n99 GND.n96 0.145
R904 GND.n102 GND.n99 0.145
R905 GND.n110 GND.n102 0.145
R906 GND.n113 GND.n110 0.145
R907 GND.n116 GND.n113 0.145
R908 GND GND.n116 0.145
R909 GND GND.n233 0.145
R910 GND.n233 GND.n226 0.145
R911 GND.n226 GND.n223 0.145
R912 GND.n223 GND.n220 0.145
R913 GND.n217 GND.n214 0.145
R914 GND.n214 GND.n209 0.145
R915 GND.n209 GND.n206 0.145
R916 GND.n199 GND.n196 0.145
R917 GND.n196 GND.n193 0.145
R918 GND.n193 GND.n190 0.145
R919 GND.n190 GND.n187 0.145
R920 GND.n187 GND.n184 0.145
R921 GND.n181 GND.n178 0.145
R922 GND.n178 GND.n175 0.145
R923 GND.n175 GND.n172 0.145
R924 GND.n172 GND.n164 0.145
R925 GND.n164 GND.n161 0.145
R926 GND.n154 GND.n151 0.145
R927 GND.n151 GND.n148 0.145
R928 GND.n148 GND.n145 0.145
R929 GND.n145 GND.n142 0.145
R930 GND.n142 GND.n139 0.145
R931 GND.n136 GND.n133 0.145
R932 GND.n133 GND.n130 0.145
R933 GND.n130 GND.n127 0.145
R934 GND.n127 GND.n122 0.145
R935 GND.n122 GND.n119 0.145
R936 a_3924_210.n9 a_3924_210.n7 82.852
R937 a_3924_210.n3 a_3924_210.n1 44.628
R938 a_3924_210.t0 a_3924_210.n9 32.417
R939 a_3924_210.n7 a_3924_210.n6 27.2
R940 a_3924_210.n5 a_3924_210.n4 23.498
R941 a_3924_210.n3 a_3924_210.n2 23.284
R942 a_3924_210.n7 a_3924_210.n5 22.4
R943 a_3924_210.t0 a_3924_210.n11 20.241
R944 a_3924_210.n11 a_3924_210.n10 13.494
R945 a_3924_210.t0 a_3924_210.n0 8.137
R946 a_3924_210.t0 a_3924_210.n3 5.727
R947 a_3924_210.n9 a_3924_210.n8 1.435
R948 a_3643_103.n5 a_3643_103.n4 19.724
R949 a_3643_103.t0 a_3643_103.n3 11.595
R950 a_3643_103.t0 a_3643_103.n5 9.207
R951 a_3643_103.n2 a_3643_103.n1 2.455
R952 a_3643_103.n2 a_3643_103.n0 1.32
R953 a_3643_103.t0 a_3643_103.n2 0.246
R954 a_4626_101.t0 a_4626_101.n1 34.62
R955 a_4626_101.t0 a_4626_101.n0 8.137
R956 a_4626_101.t0 a_4626_101.n2 4.69
R957 a_1334_210.n9 a_1334_210.n7 82.852
R958 a_1334_210.n3 a_1334_210.n1 44.628
R959 a_1334_210.t0 a_1334_210.n9 32.417
R960 a_1334_210.n7 a_1334_210.n6 27.2
R961 a_1334_210.n5 a_1334_210.n4 23.498
R962 a_1334_210.n3 a_1334_210.n2 23.284
R963 a_1334_210.n7 a_1334_210.n5 22.4
R964 a_1334_210.t0 a_1334_210.n11 20.241
R965 a_1334_210.n11 a_1334_210.n10 13.494
R966 a_1334_210.t0 a_1334_210.n0 8.137
R967 a_1334_210.t0 a_1334_210.n3 5.727
R968 a_1334_210.n9 a_1334_210.n8 1.435
R969 a_2681_103.n5 a_2681_103.n4 19.724
R970 a_2681_103.t0 a_2681_103.n3 11.595
R971 a_2681_103.t0 a_2681_103.n5 9.207
R972 a_2681_103.n2 a_2681_103.n1 2.455
R973 a_2681_103.n2 a_2681_103.n0 1.32
R974 a_2681_103.t0 a_2681_103.n2 0.246
R975 a_1053_103.n5 a_1053_103.n4 19.724
R976 a_1053_103.t0 a_1053_103.n3 11.595
R977 a_1053_103.t0 a_1053_103.n5 9.207
R978 a_1053_103.n2 a_1053_103.n1 2.455
R979 a_1053_103.n2 a_1053_103.n0 1.32
R980 a_1053_103.t0 a_1053_103.n2 0.246
C11 RN GND 2.65fF
C12 VDD GND 19.27fF
C13 a_1053_103.n0 GND 0.10fF
C14 a_1053_103.n1 GND 0.04fF
C15 a_1053_103.n2 GND 0.03fF
C16 a_1053_103.n3 GND 0.07fF
C17 a_1053_103.n4 GND 0.08fF
C18 a_1053_103.n5 GND 0.06fF
C19 a_2681_103.n0 GND 0.10fF
C20 a_2681_103.n1 GND 0.04fF
C21 a_2681_103.n2 GND 0.03fF
C22 a_2681_103.n3 GND 0.07fF
C23 a_2681_103.n4 GND 0.08fF
C24 a_2681_103.n5 GND 0.06fF
C25 a_1334_210.n0 GND 0.07fF
C26 a_1334_210.n1 GND 0.09fF
C27 a_1334_210.n2 GND 0.13fF
C28 a_1334_210.n3 GND 0.11fF
C29 a_1334_210.n4 GND 0.02fF
C30 a_1334_210.n5 GND 0.03fF
C31 a_1334_210.n6 GND 0.02fF
C32 a_1334_210.n7 GND 0.05fF
C33 a_1334_210.n8 GND 0.03fF
C34 a_1334_210.n9 GND 0.11fF
C35 a_1334_210.n10 GND 0.06fF
C36 a_1334_210.n11 GND 0.01fF
C37 a_1334_210.t0 GND 0.33fF
C38 a_4626_101.n0 GND 0.05fF
C39 a_4626_101.n1 GND 0.12fF
C40 a_4626_101.n2 GND 0.04fF
C41 a_3643_103.n0 GND 0.10fF
C42 a_3643_103.n1 GND 0.04fF
C43 a_3643_103.n2 GND 0.03fF
C44 a_3643_103.n3 GND 0.07fF
C45 a_3643_103.n4 GND 0.08fF
C46 a_3643_103.n5 GND 0.06fF
C47 a_3924_210.n0 GND 0.07fF
C48 a_3924_210.n1 GND 0.09fF
C49 a_3924_210.n2 GND 0.13fF
C50 a_3924_210.n3 GND 0.11fF
C51 a_3924_210.n4 GND 0.02fF
C52 a_3924_210.n5 GND 0.03fF
C53 a_3924_210.n6 GND 0.02fF
C54 a_3924_210.n7 GND 0.05fF
C55 a_3924_210.n8 GND 0.03fF
C56 a_3924_210.n9 GND 0.11fF
C57 a_3924_210.n10 GND 0.06fF
C58 a_3924_210.n11 GND 0.01fF
C59 a_91_103.n0 GND 0.10fF
C60 a_91_103.n1 GND 0.04fF
C61 a_91_103.n2 GND 0.03fF
C62 a_91_103.n3 GND 0.03fF
C63 a_91_103.n4 GND 0.05fF
C64 a_91_103.n5 GND 0.08fF
C65 a_91_103.n6 GND 0.07fF
C66 QN.n0 GND 0.32fF
C67 QN.n1 GND 0.34fF
C68 QN.n2 GND 0.46fF
C69 QN.n3 GND 0.46fF
C70 QN.n4 GND 0.54fF
C71 QN.n5 GND 0.17fF
C72 QN.n6 GND 0.26fF
C73 QN.n7 GND 0.03fF
C74 QN.n8 GND 0.05fF
C75 QN.n9 GND 0.03fF
C76 QN.n10 GND 0.26fF
C77 QN.n11 GND 0.38fF
C78 QN.n12 GND 0.29fF
C79 a_2962_210.n0 GND 0.02fF
C80 a_2962_210.n1 GND 0.09fF
C81 a_2962_210.n2 GND 0.13fF
C82 a_2962_210.n3 GND 0.11fF
C83 a_2962_210.t1 GND 0.30fF
C84 a_2962_210.n4 GND 0.09fF
C85 a_2962_210.n5 GND 0.06fF
C86 a_2962_210.n6 GND 0.01fF
C87 a_2962_210.n7 GND 0.03fF
C88 a_2962_210.n8 GND 0.11fF
C89 a_2962_210.n9 GND 0.02fF
C90 a_2962_210.n10 GND 0.05fF
C91 a_2962_210.n11 GND 0.02fF
C92 a_372_210.n0 GND 0.07fF
C93 a_372_210.n1 GND 0.09fF
C94 a_372_210.n2 GND 0.13fF
C95 a_372_210.n3 GND 0.11fF
C96 a_372_210.n4 GND 0.02fF
C97 a_372_210.n5 GND 0.03fF
C98 a_372_210.n6 GND 0.06fF
C99 a_372_210.n7 GND 0.03fF
C100 a_372_210.n8 GND 0.12fF
C101 a_372_210.n9 GND 0.06fF
C102 a_372_210.n10 GND 0.01fF
C103 a_372_210.t0 GND 0.33fF
C104 a_599_989.n0 GND 0.57fF
C105 a_599_989.n1 GND 0.57fF
C106 a_599_989.n2 GND 0.40fF
C107 a_599_989.n3 GND 0.42fF
C108 a_599_989.n4 GND 0.40fF
C109 a_599_989.t7 GND 0.57fF
C110 a_599_989.n5 GND 0.42fF
C111 a_599_989.n6 GND 1.32fF
C112 a_599_989.n7 GND 0.04fF
C113 a_599_989.n8 GND 0.06fF
C114 a_599_989.n9 GND 0.04fF
C115 a_599_989.n10 GND 0.32fF
C116 a_599_989.n11 GND 0.48fF
C117 a_599_989.n12 GND 0.32fF
C118 a_599_989.n13 GND 0.21fF
C119 a_599_989.n14 GND 0.67fF
C120 a_277_1050.n0 GND 0.74fF
C121 a_277_1050.n1 GND 0.74fF
C122 a_277_1050.n2 GND 0.42fF
C123 a_277_1050.n3 GND 0.83fF
C124 a_277_1050.n4 GND 0.42fF
C125 a_277_1050.n5 GND 0.66fF
C126 a_277_1050.n6 GND 3.24fF
C127 a_277_1050.n7 GND 0.59fF
C128 a_277_1050.n8 GND 0.66fF
C129 a_277_1050.n9 GND 0.38fF
C130 a_277_1050.n10 GND 0.27fF
C131 a_277_1050.n11 GND 0.87fF
C132 Q.n0 GND 0.54fF
C133 Q.n1 GND 0.64fF
C134 Q.n2 GND 0.28fF
C135 Q.n3 GND 0.04fF
C136 Q.n4 GND 0.05fF
C137 Q.n5 GND 0.03fF
C138 Q.n6 GND 0.34fF
C139 Q.n7 GND 0.43fF
C140 Q.n8 GND 0.35fF
C141 Q.n9 GND 0.39fF
C142 Q.n10 GND 0.03fF
C143 VDD.n0 GND 0.15fF
C144 VDD.n1 GND 0.02fF
C145 VDD.n2 GND 0.02fF
C146 VDD.n3 GND 0.04fF
C147 VDD.n4 GND 0.01fF
C148 VDD.n6 GND 0.02fF
C149 VDD.n7 GND 0.02fF
C150 VDD.n8 GND 0.02fF
C151 VDD.n9 GND 0.02fF
C152 VDD.n11 GND 0.02fF
C153 VDD.n14 GND 0.45fF
C154 VDD.n16 GND 0.03fF
C155 VDD.n17 GND 0.02fF
C156 VDD.n18 GND 0.02fF
C157 VDD.n19 GND 0.02fF
C158 VDD.n20 GND 0.04fF
C159 VDD.n21 GND 0.27fF
C160 VDD.n22 GND 0.02fF
C161 VDD.n23 GND 0.03fF
C162 VDD.n24 GND 0.14fF
C163 VDD.n25 GND 0.17fF
C164 VDD.n26 GND 0.01fF
C165 VDD.n27 GND 0.11fF
C166 VDD.n28 GND 0.03fF
C167 VDD.n29 GND 0.30fF
C168 VDD.n30 GND 0.01fF
C169 VDD.n31 GND 0.02fF
C170 VDD.n32 GND 0.02fF
C171 VDD.n33 GND 0.06fF
C172 VDD.n34 GND 0.24fF
C173 VDD.n35 GND 0.01fF
C174 VDD.n36 GND 0.01fF
C175 VDD.n37 GND 0.00fF
C176 VDD.n38 GND 0.09fF
C177 VDD.n39 GND 0.03fF
C178 VDD.n40 GND 0.17fF
C179 VDD.n41 GND 0.14fF
C180 VDD.n42 GND 0.01fF
C181 VDD.n43 GND 0.02fF
C182 VDD.n44 GND 0.03fF
C183 VDD.n45 GND 0.14fF
C184 VDD.n46 GND 0.16fF
C185 VDD.n47 GND 0.01fF
C186 VDD.n48 GND 0.02fF
C187 VDD.n49 GND 0.02fF
C188 VDD.n50 GND 0.06fF
C189 VDD.n51 GND 0.25fF
C190 VDD.n52 GND 0.01fF
C191 VDD.n53 GND 0.01fF
C192 VDD.n54 GND 0.02fF
C193 VDD.n55 GND 0.27fF
C194 VDD.n56 GND 0.01fF
C195 VDD.n57 GND 0.02fF
C196 VDD.n58 GND 0.03fF
C197 VDD.n59 GND 0.02fF
C198 VDD.n60 GND 0.02fF
C199 VDD.n61 GND 0.02fF
C200 VDD.n62 GND 0.26fF
C201 VDD.n63 GND 0.04fF
C202 VDD.n64 GND 0.04fF
C203 VDD.n65 GND 0.02fF
C204 VDD.n67 GND 0.02fF
C205 VDD.n68 GND 0.02fF
C206 VDD.n69 GND 0.02fF
C207 VDD.n70 GND 0.02fF
C208 VDD.n72 GND 0.02fF
C209 VDD.n73 GND 0.02fF
C210 VDD.n74 GND 0.02fF
C211 VDD.n76 GND 0.27fF
C212 VDD.n78 GND 0.02fF
C213 VDD.n79 GND 0.02fF
C214 VDD.n80 GND 0.03fF
C215 VDD.n81 GND 0.02fF
C216 VDD.n82 GND 0.27fF
C217 VDD.n83 GND 0.01fF
C218 VDD.n84 GND 0.02fF
C219 VDD.n85 GND 0.03fF
C220 VDD.n86 GND 0.27fF
C221 VDD.n87 GND 0.01fF
C222 VDD.n88 GND 0.02fF
C223 VDD.n89 GND 0.02fF
C224 VDD.n90 GND 0.22fF
C225 VDD.n91 GND 0.01fF
C226 VDD.n92 GND 0.07fF
C227 VDD.n93 GND 0.02fF
C228 VDD.n94 GND 0.14fF
C229 VDD.n95 GND 0.17fF
C230 VDD.n96 GND 0.01fF
C231 VDD.n97 GND 0.02fF
C232 VDD.n98 GND 0.02fF
C233 VDD.n99 GND 0.14fF
C234 VDD.n100 GND 0.16fF
C235 VDD.n101 GND 0.01fF
C236 VDD.n102 GND 0.11fF
C237 VDD.n103 GND 0.02fF
C238 VDD.n104 GND 0.02fF
C239 VDD.n105 GND 0.02fF
C240 VDD.n106 GND 0.17fF
C241 VDD.n107 GND 0.14fF
C242 VDD.n108 GND 0.01fF
C243 VDD.n109 GND 0.02fF
C244 VDD.n110 GND 0.03fF
C245 VDD.n111 GND 0.18fF
C246 VDD.n112 GND 0.15fF
C247 VDD.n113 GND 0.01fF
C248 VDD.n114 GND 0.02fF
C249 VDD.n115 GND 0.03fF
C250 VDD.n116 GND 0.11fF
C251 VDD.n117 GND 0.02fF
C252 VDD.n118 GND 0.14fF
C253 VDD.n119 GND 0.15fF
C254 VDD.n120 GND 0.01fF
C255 VDD.n121 GND 0.02fF
C256 VDD.n122 GND 0.02fF
C257 VDD.n123 GND 0.14fF
C258 VDD.n124 GND 0.17fF
C259 VDD.n125 GND 0.01fF
C260 VDD.n126 GND 0.02fF
C261 VDD.n127 GND 0.02fF
C262 VDD.n128 GND 0.06fF
C263 VDD.n129 GND 0.22fF
C264 VDD.n130 GND 0.01fF
C265 VDD.n131 GND 0.01fF
C266 VDD.n132 GND 0.02fF
C267 VDD.n133 GND 0.27fF
C268 VDD.n134 GND 0.01fF
C269 VDD.n135 GND 0.02fF
C270 VDD.n136 GND 0.02fF
C271 VDD.n137 GND 0.27fF
C272 VDD.n138 GND 0.01fF
C273 VDD.n139 GND 0.02fF
C274 VDD.n140 GND 0.03fF
C275 VDD.n141 GND 0.02fF
C276 VDD.n142 GND 0.02fF
C277 VDD.n143 GND 0.02fF
C278 VDD.n144 GND 0.31fF
C279 VDD.n145 GND 0.04fF
C280 VDD.n146 GND 0.03fF
C281 VDD.n147 GND 0.02fF
C282 VDD.n148 GND 0.02fF
C283 VDD.n149 GND 0.02fF
C284 VDD.n150 GND 0.02fF
C285 VDD.n151 GND 0.02fF
C286 VDD.n153 GND 0.02fF
C287 VDD.n154 GND 0.02fF
C288 VDD.n155 GND 0.02fF
C289 VDD.n157 GND 0.27fF
C290 VDD.n159 GND 0.02fF
C291 VDD.n160 GND 0.02fF
C292 VDD.n161 GND 0.03fF
C293 VDD.n162 GND 0.02fF
C294 VDD.n163 GND 0.27fF
C295 VDD.n164 GND 0.01fF
C296 VDD.n165 GND 0.02fF
C297 VDD.n166 GND 0.03fF
C298 VDD.n167 GND 0.27fF
C299 VDD.n168 GND 0.01fF
C300 VDD.n169 GND 0.02fF
C301 VDD.n170 GND 0.02fF
C302 VDD.n171 GND 0.22fF
C303 VDD.n172 GND 0.01fF
C304 VDD.n173 GND 0.07fF
C305 VDD.n174 GND 0.02fF
C306 VDD.n175 GND 0.14fF
C307 VDD.n176 GND 0.17fF
C308 VDD.n177 GND 0.01fF
C309 VDD.n178 GND 0.02fF
C310 VDD.n179 GND 0.02fF
C311 VDD.n180 GND 0.14fF
C312 VDD.n181 GND 0.16fF
C313 VDD.n182 GND 0.01fF
C314 VDD.n183 GND 0.11fF
C315 VDD.n184 GND 0.02fF
C316 VDD.n185 GND 0.02fF
C317 VDD.n186 GND 0.02fF
C318 VDD.n187 GND 0.17fF
C319 VDD.n188 GND 0.14fF
C320 VDD.n189 GND 0.01fF
C321 VDD.n190 GND 0.02fF
C322 VDD.n191 GND 0.03fF
C323 VDD.n192 GND 0.18fF
C324 VDD.n193 GND 0.15fF
C325 VDD.n194 GND 0.01fF
C326 VDD.n195 GND 0.02fF
C327 VDD.n196 GND 0.03fF
C328 VDD.n197 GND 0.11fF
C329 VDD.n198 GND 0.02fF
C330 VDD.n199 GND 0.14fF
C331 VDD.n200 GND 0.15fF
C332 VDD.n201 GND 0.01fF
C333 VDD.n202 GND 0.02fF
C334 VDD.n203 GND 0.02fF
C335 VDD.n204 GND 0.14fF
C336 VDD.n205 GND 0.17fF
C337 VDD.n206 GND 0.01fF
C338 VDD.n207 GND 0.02fF
C339 VDD.n208 GND 0.02fF
C340 VDD.n209 GND 0.06fF
C341 VDD.n210 GND 0.22fF
C342 VDD.n211 GND 0.01fF
C343 VDD.n212 GND 0.01fF
C344 VDD.n213 GND 0.02fF
C345 VDD.n214 GND 0.27fF
C346 VDD.n215 GND 0.01fF
C347 VDD.n216 GND 0.02fF
C348 VDD.n217 GND 0.02fF
C349 VDD.n218 GND 0.02fF
C350 VDD.n219 GND 0.02fF
C351 VDD.n220 GND 0.02fF
C352 VDD.n221 GND 0.26fF
C353 VDD.n222 GND 0.04fF
C354 VDD.n223 GND 0.03fF
C355 VDD.n224 GND 0.02fF
C356 VDD.n225 GND 0.02fF
C357 VDD.n226 GND 0.02fF
C358 VDD.n227 GND 0.02fF
C359 VDD.n228 GND 0.02fF
C360 VDD.n230 GND 0.02fF
C361 VDD.n231 GND 0.02fF
C362 VDD.n232 GND 0.02fF
C363 VDD.n234 GND 0.27fF
C364 VDD.n236 GND 0.02fF
C365 VDD.n237 GND 0.02fF
C366 VDD.n238 GND 0.03fF
C367 VDD.n239 GND 0.27fF
C368 VDD.n240 GND 0.01fF
C369 VDD.n241 GND 0.02fF
C370 VDD.n242 GND 0.02fF
C371 VDD.n243 GND 0.02fF
C372 VDD.n244 GND 0.02fF
C373 VDD.n245 GND 0.02fF
C374 VDD.n246 GND 0.20fF
C375 VDD.n247 GND 0.03fF
C376 VDD.n248 GND 0.02fF
C377 VDD.n249 GND 0.02fF
C378 VDD.n250 GND 0.02fF
C379 VDD.n251 GND 0.02fF
C380 VDD.n252 GND 0.02fF
C381 VDD.n254 GND 0.02fF
C382 VDD.n255 GND 0.02fF
C383 VDD.n256 GND 0.02fF
C384 VDD.n258 GND 0.45fF
C385 VDD.n260 GND 0.03fF
C386 VDD.n261 GND 0.04fF
C387 VDD.n262 GND 0.27fF
C388 VDD.n263 GND 0.02fF
C389 VDD.n264 GND 0.03fF
C390 VDD.n265 GND 0.03fF
C391 VDD.n266 GND 0.27fF
C392 VDD.n267 GND 0.01fF
C393 VDD.n268 GND 0.02fF
C394 VDD.n269 GND 0.02fF
C395 VDD.n270 GND 0.06fF
C396 VDD.n271 GND 0.22fF
C397 VDD.n272 GND 0.01fF
C398 VDD.n273 GND 0.01fF
C399 VDD.n274 GND 0.02fF
C400 VDD.n275 GND 0.14fF
C401 VDD.n276 GND 0.17fF
C402 VDD.n277 GND 0.01fF
C403 VDD.n278 GND 0.02fF
C404 VDD.n279 GND 0.02fF
C405 VDD.n280 GND 0.11fF
C406 VDD.n281 GND 0.02fF
C407 VDD.n282 GND 0.14fF
C408 VDD.n283 GND 0.15fF
C409 VDD.n284 GND 0.01fF
C410 VDD.n285 GND 0.02fF
C411 VDD.n286 GND 0.02fF
C412 VDD.n287 GND 0.18fF
C413 VDD.n288 GND 0.15fF
C414 VDD.n289 GND 0.01fF
C415 VDD.n290 GND 0.02fF
C416 VDD.n291 GND 0.03fF
C417 VDD.n292 GND 0.17fF
C418 VDD.n293 GND 0.14fF
C419 VDD.n294 GND 0.01fF
C420 VDD.n295 GND 0.02fF
C421 VDD.n296 GND 0.03fF
C422 VDD.n297 GND 0.14fF
C423 VDD.n298 GND 0.16fF
C424 VDD.n299 GND 0.01fF
C425 VDD.n300 GND 0.11fF
C426 VDD.n301 GND 0.02fF
C427 VDD.n302 GND 0.02fF
C428 VDD.n303 GND 0.02fF
C429 VDD.n304 GND 0.14fF
C430 VDD.n305 GND 0.17fF
C431 VDD.n306 GND 0.01fF
C432 VDD.n307 GND 0.02fF
C433 VDD.n308 GND 0.02fF
C434 VDD.n309 GND 0.22fF
C435 VDD.n310 GND 0.01fF
C436 VDD.n311 GND 0.07fF
C437 VDD.n312 GND 0.02fF
C438 VDD.n313 GND 0.27fF
C439 VDD.n314 GND 0.01fF
C440 VDD.n315 GND 0.02fF
C441 VDD.n316 GND 0.02fF
C442 VDD.n317 GND 0.27fF
C443 VDD.n318 GND 0.01fF
C444 VDD.n319 GND 0.02fF
C445 VDD.n320 GND 0.03fF
C446 VDD.n321 GND 0.02fF
C447 VDD.n322 GND 0.02fF
C448 VDD.n323 GND 0.02fF
C449 VDD.n324 GND 0.02fF
C450 VDD.n325 GND 0.02fF
C451 VDD.n326 GND 0.02fF
C452 VDD.n328 GND 0.02fF
C453 VDD.n329 GND 0.02fF
C454 VDD.n330 GND 0.02fF
C455 VDD.n331 GND 0.02fF
C456 VDD.n333 GND 0.04fF
C457 VDD.n334 GND 0.02fF
C458 VDD.n335 GND 0.31fF
C459 VDD.n336 GND 0.04fF
C460 VDD.n338 GND 0.27fF
C461 VDD.n340 GND 0.02fF
C462 VDD.n341 GND 0.02fF
C463 VDD.n342 GND 0.03fF
C464 VDD.n343 GND 0.02fF
C465 VDD.n344 GND 0.27fF
C466 VDD.n345 GND 0.01fF
C467 VDD.n346 GND 0.02fF
C468 VDD.n347 GND 0.03fF
C469 VDD.n348 GND 0.27fF
C470 VDD.n349 GND 0.01fF
C471 VDD.n350 GND 0.02fF
C472 VDD.n351 GND 0.02fF
C473 VDD.n352 GND 0.06fF
C474 VDD.n353 GND 0.22fF
C475 VDD.n354 GND 0.01fF
C476 VDD.n355 GND 0.01fF
C477 VDD.n356 GND 0.02fF
C478 VDD.n357 GND 0.14fF
C479 VDD.n358 GND 0.17fF
C480 VDD.n359 GND 0.01fF
C481 VDD.n360 GND 0.02fF
C482 VDD.n361 GND 0.02fF
C483 VDD.n362 GND 0.11fF
C484 VDD.n363 GND 0.02fF
C485 VDD.n364 GND 0.14fF
C486 VDD.n365 GND 0.15fF
C487 VDD.n366 GND 0.01fF
C488 VDD.n367 GND 0.02fF
C489 VDD.n368 GND 0.02fF
C490 VDD.n369 GND 0.18fF
C491 VDD.n370 GND 0.15fF
C492 VDD.n371 GND 0.01fF
C493 VDD.n372 GND 0.02fF
C494 VDD.n373 GND 0.03fF
C495 VDD.n374 GND 0.17fF
C496 VDD.n375 GND 0.14fF
C497 VDD.n376 GND 0.01fF
C498 VDD.n377 GND 0.02fF
C499 VDD.n378 GND 0.03fF
C500 VDD.n379 GND 0.14fF
C501 VDD.n380 GND 0.16fF
C502 VDD.n381 GND 0.01fF
C503 VDD.n382 GND 0.11fF
C504 VDD.n383 GND 0.02fF
C505 VDD.n384 GND 0.02fF
C506 VDD.n385 GND 0.02fF
C507 VDD.n386 GND 0.14fF
C508 VDD.n387 GND 0.17fF
C509 VDD.n388 GND 0.01fF
C510 VDD.n389 GND 0.02fF
C511 VDD.n390 GND 0.02fF
C512 VDD.n391 GND 0.22fF
C513 VDD.n392 GND 0.01fF
C514 VDD.n393 GND 0.07fF
C515 VDD.n394 GND 0.02fF
C516 VDD.n395 GND 0.27fF
C517 VDD.n396 GND 0.01fF
C518 VDD.n397 GND 0.02fF
C519 VDD.n398 GND 0.02fF
C520 VDD.n399 GND 0.27fF
C521 VDD.n400 GND 0.01fF
C522 VDD.n401 GND 0.02fF
C523 VDD.n402 GND 0.03fF
C524 VDD.n403 GND 0.02fF
C525 VDD.n404 GND 0.02fF
C526 VDD.n405 GND 0.02fF
C527 VDD.n406 GND 0.26fF
C528 VDD.n407 GND 0.04fF
C529 VDD.n408 GND 0.03fF
C530 VDD.n409 GND 0.02fF
C531 VDD.n410 GND 0.02fF
C532 VDD.n411 GND 0.02fF
C533 VDD.n412 GND 0.02fF
C534 VDD.n413 GND 0.02fF
C535 VDD.n415 GND 0.02fF
C536 VDD.n416 GND 0.02fF
C537 VDD.n417 GND 0.02fF
C538 VDD.n419 GND 0.27fF
C539 VDD.n421 GND 0.02fF
C540 VDD.n422 GND 0.02fF
C541 VDD.n423 GND 0.03fF
C542 VDD.n424 GND 0.02fF
C543 VDD.n425 GND 0.27fF
C544 VDD.n426 GND 0.01fF
C545 VDD.n427 GND 0.02fF
C546 VDD.n428 GND 0.03fF
C547 VDD.n429 GND 0.06fF
C548 VDD.n430 GND 0.25fF
C549 VDD.n431 GND 0.01fF
C550 VDD.n432 GND 0.01fF
C551 VDD.n433 GND 0.02fF
C552 VDD.n434 GND 0.14fF
C553 VDD.n435 GND 0.16fF
C554 VDD.n436 GND 0.01fF
C555 VDD.n437 GND 0.02fF
C556 VDD.n438 GND 0.02fF
C557 VDD.n439 GND 0.17fF
C558 VDD.n440 GND 0.14fF
C559 VDD.n441 GND 0.01fF
C560 VDD.n442 GND 0.02fF
C561 VDD.n443 GND 0.03fF
C562 VDD.n444 GND 0.11fF
C563 VDD.n445 GND 0.03fF
C564 VDD.n446 GND 0.30fF
C565 VDD.n447 GND 0.01fF
C566 VDD.n448 GND 0.02fF
C567 VDD.n449 GND 0.03fF
C568 VDD.n450 GND 0.14fF
C569 VDD.n451 GND 0.17fF
C570 VDD.n452 GND 0.01fF
C571 VDD.n453 GND 0.02fF
C572 VDD.n454 GND 0.02fF
C573 VDD.n455 GND 0.06fF
C574 VDD.n456 GND 0.24fF
C575 VDD.n457 GND 0.01fF
C576 VDD.n458 GND 0.01fF
C577 VDD.n459 GND 0.02fF
C578 VDD.n460 GND 0.02fF
C579 VDD.n461 GND 0.27fF
C580 VDD.n462 GND 0.01fF
C581 VDD.n463 GND 0.02fF
C582 VDD.n464 GND 0.02fF
C583 RN.n0 GND 0.39fF
C584 RN.t6 GND 0.35fF
C585 RN.n1 GND 0.30fF
C586 RN.n2 GND 0.38fF
C587 RN.t1 GND 0.36fF
C588 RN.n3 GND 0.29fF
C589 RN.n4 GND 1.05fF
C590 RN.n5 GND 0.38fF
C591 RN.t4 GND 0.37fF
C592 RN.n6 GND 0.29fF
C593 RN.n7 GND 0.55fF
C594 a_2141_1050.n0 GND 0.52fF
C595 a_2141_1050.n1 GND 0.61fF
C596 a_2141_1050.n2 GND 0.30fF
C597 a_2141_1050.n3 GND 0.33fF
C598 a_2141_1050.n4 GND 0.64fF
C599 a_2141_1050.n5 GND 0.60fF
C600 a_2141_1050.n6 GND 0.08fF
C601 a_2141_1050.n7 GND 0.28fF
C602 a_2141_1050.n8 GND 0.04fF
C603 a_2036_101.n0 GND 0.05fF
C604 a_2036_101.n1 GND 0.12fF
C605 a_2036_101.n2 GND 0.04fF
C606 a_147_187.n0 GND 0.06fF
C607 a_147_187.n1 GND 0.73fF
C608 a_147_187.n2 GND 0.73fF
C609 a_147_187.n3 GND 0.86fF
C610 a_147_187.n4 GND 0.27fF
C611 a_147_187.n5 GND 0.33fF
C612 a_147_187.n6 GND 0.38fF
C613 a_147_187.n7 GND 0.58fF
C614 a_147_187.n8 GND 0.38fF
C615 a_147_187.t7 GND 0.81fF
C616 a_147_187.n9 GND 0.52fF
C617 a_147_187.n10 GND 0.37fF
C618 a_147_187.n11 GND 0.77fF
C619 a_147_187.n12 GND 2.88fF
C620 a_147_187.n13 GND 2.27fF
C621 a_147_187.n14 GND 0.62fF
C622 a_147_187.n15 GND 0.06fF
C623 a_147_187.n16 GND 0.50fF
C624 a_147_187.n17 GND 0.06fF
.ends
