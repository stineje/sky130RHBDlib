magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 106 157 584 203
rect 1 21 735 157
rect 30 -17 64 21
<< locali >>
rect 17 215 97 264
rect 607 313 719 493
rect 646 128 719 313
rect 603 51 719 128
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 332 86 493
rect 120 366 185 527
rect 239 358 329 493
rect 17 298 201 332
rect 131 259 201 298
rect 131 205 221 259
rect 294 250 329 358
rect 363 333 413 493
rect 447 367 569 527
rect 363 299 553 333
rect 519 265 553 299
rect 294 215 484 250
rect 131 181 201 205
rect 17 147 201 181
rect 294 171 329 215
rect 519 198 610 265
rect 519 181 553 198
rect 17 51 82 147
rect 116 17 182 113
rect 235 51 329 171
rect 363 147 553 181
rect 363 51 413 147
rect 448 17 569 113
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 17 215 97 264 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 735 157 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 106 157 584 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 603 51 719 128 6 X
port 6 nsew signal output
rlabel locali s 646 128 719 313 6 X
port 6 nsew signal output
rlabel locali s 607 313 719 493 6 X
port 6 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3261692
string GDS_START 3255572
<< end >>
