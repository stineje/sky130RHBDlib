* SPICE3 file created from BUFX1.ext - technology: sky130A

.subckt BUFX1 Y A VPB VNB
M1000 VPB.t3 a_185_182.t3 a_629_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_629_182.t0 a_185_182.t4 VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPB.t1 a_121_384# a_185_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_185_182.t0 a_121_384# VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u

R0 a_185_182.n2 a_185_182.t3 512.525
R1 a_185_182.n2 a_185_182.t4 371.139
R2 a_185_182.n4 a_185_182.n1 220.249
R3 a_185_182.n3 a_185_182.n2 211.406
R4 a_185_182.n3 a_185_182.t5 167.157
R5 a_185_182.n4 a_185_182.n3 153.043
R6 a_185_182.n6 a_185_182.n4 135.599
R7 a_185_182.n6 a_185_182.n5 30
R8 a_185_182.n7 a_185_182.n0 24.383
R9 a_185_182.n7 a_185_182.n6 23.684
R10 a_185_182.n1 a_185_182.t1 14.282
R11 a_185_182.n1 a_185_182.t0 14.282
R12 a_629_182.n3 a_629_182.n1 355.848
R13 a_629_182.n3 a_629_182.n2 30
R14 a_629_182.n4 a_629_182.n0 24.383
R15 a_629_182.n4 a_629_182.n3 23.684
R16 a_629_182.n1 a_629_182.t1 14.282
R17 a_629_182.n1 a_629_182.t0 14.282
R18 VPB VPB.n109 126.832
R19 VPB.n90 VPB.n88 94.117
R20 VPB.n96 VPB.n95 76
R21 VPB.n102 VPB.n101 76
R22 VPB.n51 VPB.n50 68.979
R23 VPB.n77 VPB.n76 68.979
R24 VPB.n44 VPB.n43 64.528
R25 VPB.n84 VPB.n83 64.528
R26 VPB.n61 VPB.n60 61.764
R27 VPB.n14 VPB.t0 55.106
R28 VPB.n87 VPB.t1 55.106
R29 VPB.n54 VPB.t2 55.106
R30 VPB.n42 VPB.t3 55.106
R31 VPB.n106 VPB.n102 20.452
R32 VPB.n41 VPB.n38 20.452
R33 VPB.n41 VPB.n40 13.653
R34 VPB.n40 VPB.n39 13.653
R35 VPB.n46 VPB.n45 13.653
R36 VPB.n45 VPB.n44 13.653
R37 VPB.n49 VPB.n48 13.653
R38 VPB.n48 VPB.n47 13.653
R39 VPB.n53 VPB.n52 13.653
R40 VPB.n52 VPB.n51 13.653
R41 VPB.n95 VPB.n94 13.653
R42 VPB.n94 VPB.n93 13.653
R43 VPB.n91 VPB.n90 13.653
R44 VPB.n90 VPB.n89 13.653
R45 VPB.n86 VPB.n85 13.653
R46 VPB.n85 VPB.n84 13.653
R47 VPB.n82 VPB.n81 13.653
R48 VPB.n81 VPB.n80 13.653
R49 VPB.n79 VPB.n78 13.653
R50 VPB.n78 VPB.n77 13.653
R51 VPB.n102 VPB.n0 13.653
R52 VPB VPB.n0 13.653
R53 VPB.n106 VPB.n105 13.276
R54 VPB.n105 VPB.n103 13.276
R55 VPB.n75 VPB.n57 13.276
R56 VPB.n57 VPB.n55 13.276
R57 VPB.n49 VPB.n46 13.276
R58 VPB.n53 VPB.n49 13.276
R59 VPB.n95 VPB.n92 13.276
R60 VPB.n92 VPB.n91 13.276
R61 VPB.n86 VPB.n82 13.276
R62 VPB.n82 VPB.n79 13.276
R63 VPB.n38 VPB.n20 13.276
R64 VPB.n20 VPB.n18 13.276
R65 VPB.n25 VPB.n23 12.796
R66 VPB.n25 VPB.n24 12.564
R67 VPB.n34 VPB.n33 12.198
R68 VPB.n31 VPB.n30 12.198
R69 VPB.n28 VPB.n27 12.198
R70 VPB.n95 VPB.n54 10.944
R71 VPB.n102 VPB.n14 10.944
R72 VPB.n42 VPB.n41 10.585
R73 VPB.n91 VPB.n87 10.585
R74 VPB.n38 VPB.n37 7.5
R75 VPB.n23 VPB.n22 7.5
R76 VPB.n27 VPB.n26 7.5
R77 VPB.n30 VPB.n29 7.5
R78 VPB.n20 VPB.n19 7.5
R79 VPB.n35 VPB.n21 7.5
R80 VPB.n57 VPB.n56 7.5
R81 VPB.n70 VPB.n69 7.5
R82 VPB.n64 VPB.n63 7.5
R83 VPB.n66 VPB.n65 7.5
R84 VPB.n59 VPB.n58 7.5
R85 VPB.n75 VPB.n74 7.5
R86 VPB.n105 VPB.n104 7.5
R87 VPB.n12 VPB.n11 7.5
R88 VPB.n6 VPB.n5 7.5
R89 VPB.n8 VPB.n7 7.5
R90 VPB.n2 VPB.n1 7.5
R91 VPB.n107 VPB.n106 7.5
R92 VPB.n92 VPB.n75 7.176
R93 VPB.n71 VPB.n68 6.729
R94 VPB.n67 VPB.n64 6.729
R95 VPB.n62 VPB.n59 6.729
R96 VPB.n13 VPB.n10 6.729
R97 VPB.n9 VPB.n6 6.729
R98 VPB.n4 VPB.n2 6.729
R99 VPB.n62 VPB.n61 6.728
R100 VPB.n67 VPB.n66 6.728
R101 VPB.n71 VPB.n70 6.728
R102 VPB.n74 VPB.n73 6.728
R103 VPB.n4 VPB.n3 6.728
R104 VPB.n9 VPB.n8 6.728
R105 VPB.n13 VPB.n12 6.728
R106 VPB.n108 VPB.n107 6.728
R107 VPB.n37 VPB.n36 6.398
R108 VPB.n46 VPB.n42 2.691
R109 VPB.n87 VPB.n86 2.691
R110 VPB.n54 VPB.n53 2.332
R111 VPB.n79 VPB.n14 2.332
R112 VPB.n35 VPB.n28 1.402
R113 VPB.n35 VPB.n31 1.402
R114 VPB.n35 VPB.n32 1.402
R115 VPB.n35 VPB.n34 1.402
R116 VPB.n36 VPB.n35 0.735
R117 VPB.n35 VPB.n25 0.735
R118 VPB.n72 VPB.n71 0.387
R119 VPB.n72 VPB.n67 0.387
R120 VPB.n72 VPB.n62 0.387
R121 VPB.n73 VPB.n72 0.387
R122 VPB.n109 VPB.n13 0.387
R123 VPB.n109 VPB.n9 0.387
R124 VPB.n109 VPB.n4 0.387
R125 VPB.n109 VPB.n108 0.387
R126 VPB.n101 VPB 0.198
R127 VPB.n16 VPB.n15 0.136
R128 VPB.n17 VPB.n16 0.136
R129 VPB.n96 VPB.n17 0.136
R130 VPB VPB.n96 0.136
R131 VPB.n97 VPB 0.136
R132 VPB.n98 VPB.n97 0.136
R133 VPB.n99 VPB.n98 0.136
R134 VPB.n100 VPB.n99 0.136
R135 VPB.n101 VPB.n100 0.136
R136 VNB VNB.n114 300.778
R137 VNB.n65 VNB.n64 199.897
R138 VNB.n89 VNB.n87 154.509
R139 VNB.n101 VNB.n100 76
R140 VNB.n95 VNB.n94 76
R141 VNB.n49 VNB.n48 49.896
R142 VNB.n80 VNB.n79 49.896
R143 VNB.n24 VNB.n23 35.01
R144 VNB.n73 VNB.n72 35.01
R145 VNB.t1 VNB.n16 32.601
R146 VNB.t0 VNB.n6 32.601
R147 VNB.n42 VNB.n39 20.452
R148 VNB.n102 VNB.n101 20.452
R149 VNB.n43 VNB.n24 20.094
R150 VNB.n47 VNB.n21 20.094
R151 VNB.n54 VNB.n19 20.094
R152 VNB.n86 VNB.n73 20.094
R153 VNB.n82 VNB.n75 20.094
R154 VNB.n10 VNB.n9 20.094
R155 VNB.n24 VNB.n22 19.017
R156 VNB.n73 VNB.n71 19.017
R157 VNB.n18 VNB.t1 17.353
R158 VNB.n8 VNB.t0 17.353
R159 VNB.n46 VNB.n45 13.653
R160 VNB.n45 VNB.n44 13.653
R161 VNB.n50 VNB.n49 13.653
R162 VNB.n53 VNB.n52 13.653
R163 VNB.n52 VNB.n51 13.653
R164 VNB.n94 VNB.n93 13.653
R165 VNB.n93 VNB.n92 13.653
R166 VNB.n90 VNB.n89 13.653
R167 VNB.n89 VNB.n88 13.653
R168 VNB.n85 VNB.n84 13.653
R169 VNB.n84 VNB.n83 13.653
R170 VNB.n81 VNB.n80 13.653
R171 VNB.n78 VNB.n77 13.653
R172 VNB.n77 VNB.n76 13.653
R173 VNB.n101 VNB.n0 13.653
R174 VNB VNB.n0 13.653
R175 VNB.n42 VNB.n41 13.653
R176 VNB.n41 VNB.n40 13.653
R177 VNB.n109 VNB.n106 13.577
R178 VNB.n27 VNB.n25 13.276
R179 VNB.n39 VNB.n27 13.276
R180 VNB.n57 VNB.n55 13.276
R181 VNB.n70 VNB.n57 13.276
R182 VNB.n53 VNB.n50 13.276
R183 VNB.n94 VNB.n91 13.276
R184 VNB.n91 VNB.n90 13.276
R185 VNB.n81 VNB.n78 13.276
R186 VNB.n3 VNB.n1 13.276
R187 VNB.n102 VNB.n3 13.276
R188 VNB.n47 VNB.n46 13.097
R189 VNB.n85 VNB.n82 13.097
R190 VNB.n19 VNB.n18 12.837
R191 VNB.n9 VNB.n8 12.837
R192 VNB.n94 VNB.n54 9.329
R193 VNB.n101 VNB.n10 9.329
R194 VNB.n43 VNB.n42 8.97
R195 VNB.n90 VNB.n86 8.97
R196 VNB.n18 VNB.n17 7.566
R197 VNB.n8 VNB.n7 7.566
R198 VNB.n111 VNB.n110 7.5
R199 VNB.n63 VNB.n62 7.5
R200 VNB.n59 VNB.n58 7.5
R201 VNB.n57 VNB.n56 7.5
R202 VNB.n70 VNB.n69 7.5
R203 VNB.n103 VNB.n102 7.5
R204 VNB.n3 VNB.n2 7.5
R205 VNB.n108 VNB.n107 7.5
R206 VNB.n33 VNB.n32 7.5
R207 VNB.n29 VNB.n28 7.5
R208 VNB.n27 VNB.n26 7.5
R209 VNB.n39 VNB.n38 7.5
R210 VNB.n91 VNB.n70 7.176
R211 VNB.n113 VNB.n111 7.011
R212 VNB.n66 VNB.n63 7.011
R213 VNB.n61 VNB.n59 7.011
R214 VNB.n35 VNB.n33 7.011
R215 VNB.n31 VNB.n29 7.011
R216 VNB.n69 VNB.n68 7.01
R217 VNB.n61 VNB.n60 7.01
R218 VNB.n66 VNB.n65 7.01
R219 VNB.n38 VNB.n37 7.01
R220 VNB.n31 VNB.n30 7.01
R221 VNB.n35 VNB.n34 7.01
R222 VNB.n113 VNB.n112 7.01
R223 VNB.n109 VNB.n108 6.788
R224 VNB.n104 VNB.n103 6.788
R225 VNB.n15 VNB.n14 4.551
R226 VNB.n5 VNB.n4 4.551
R227 VNB.n46 VNB.n43 4.305
R228 VNB.n86 VNB.n85 4.305
R229 VNB.n54 VNB.n53 3.947
R230 VNB.n78 VNB.n10 3.947
R231 VNB.t1 VNB.n15 2.238
R232 VNB.t0 VNB.n5 2.238
R233 VNB.n114 VNB.n105 0.921
R234 VNB.n114 VNB.n109 0.476
R235 VNB.n114 VNB.n104 0.475
R236 VNB.n21 VNB.n20 0.358
R237 VNB.n75 VNB.n74 0.358
R238 VNB.n67 VNB.n61 0.246
R239 VNB.n68 VNB.n67 0.246
R240 VNB.n67 VNB.n66 0.246
R241 VNB.n36 VNB.n31 0.246
R242 VNB.n37 VNB.n36 0.246
R243 VNB.n36 VNB.n35 0.246
R244 VNB.n114 VNB.n113 0.246
R245 VNB.n100 VNB 0.198
R246 VNB.n50 VNB.n47 0.179
R247 VNB.n82 VNB.n81 0.179
R248 VNB.n12 VNB.n11 0.136
R249 VNB.n13 VNB.n12 0.136
R250 VNB.n95 VNB.n13 0.136
R251 VNB VNB.n95 0.136
R252 VNB.n96 VNB 0.136
R253 VNB.n97 VNB.n96 0.136
R254 VNB.n98 VNB.n97 0.136
R255 VNB.n99 VNB.n98 0.136
R256 VNB.n100 VNB.n99 0.136
















































































































.ends
