* SPICE3 file created from VOTER3X1.ext - technology: sky130A

.subckt VOTER3X1 Y A B C VDD GND
M1000 a_217_1051.t5 B.t0 a_881_1051.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_881_1051.t0 A.t0 a_392_209.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 GND B.t1 a_778_101.t0 nshort w=-1.605u l=1.765u
+  ad=1.6781p pd=12.81u as=0p ps=0u
M1003 a_217_1051.t3 A.t1 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_217_1051.t1 C.t0 a_881_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_392_209.t5 C.t1 a_881_1051.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 GND B.t2 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1007 GND C.t2 a_1444_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y.t2 a_392_209.t7 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_392_209.t9 GND.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1010 VDD.t5 B.t3 a_217_1051.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_392_209.t1 A.t3 a_881_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VDD.t1 a_392_209.t8 Y.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_881_1051.t3 C.t3 a_217_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t2 A.t5 a_217_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_881_1051.t4 C.t4 a_392_209.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_881_1051.t5 B.t4 a_217_1051.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_217_1051.t7 B.t5 VDD.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 A VDD 0.85fF
C1 A B 0.96fF
C2 C VDD 0.18fF
C3 B C 0.15fF
C4 Y VDD 0.76fF
C5 B VDD 0.28fF
C6 A C 0.26fF
R0 B.n2 B.t3 512.525
R1 B.n0 B.t0 477.179
R2 B.n0 B.t4 406.485
R3 B.n2 B.t5 371.139
R4 B.n1 B.t1 363.924
R5 B.n3 B.t2 357.498
R6 B.n3 B.n2 71.88
R7 B.n4 B.n1 52.017
R8 B.n4 B.n3 49.342
R9 B.n1 B.n0 15.776
R10 B.n4 B 0.046
R11 a_881_1051.n4 a_881_1051.n3 196.002
R12 a_881_1051.t0 a_881_1051.n5 89.556
R13 a_881_1051.n3 a_881_1051.n2 75.271
R14 a_881_1051.n5 a_881_1051.n4 75.214
R15 a_881_1051.n3 a_881_1051.n1 36.52
R16 a_881_1051.n4 a_881_1051.t7 14.338
R17 a_881_1051.n1 a_881_1051.t2 14.282
R18 a_881_1051.n1 a_881_1051.t3 14.282
R19 a_881_1051.n2 a_881_1051.t6 14.282
R20 a_881_1051.n2 a_881_1051.t5 14.282
R21 a_881_1051.n0 a_881_1051.t1 14.282
R22 a_881_1051.n0 a_881_1051.t4 14.282
R23 a_881_1051.n5 a_881_1051.n0 12.119
R24 a_217_1051.n3 a_217_1051.n2 195.987
R25 a_217_1051.n4 a_217_1051.t1 89.553
R26 a_217_1051.n2 a_217_1051.n1 75.271
R27 a_217_1051.n4 a_217_1051.n3 75.214
R28 a_217_1051.n2 a_217_1051.n0 36.519
R29 a_217_1051.n3 a_217_1051.t4 14.338
R30 a_217_1051.n0 a_217_1051.t0 14.282
R31 a_217_1051.n0 a_217_1051.t3 14.282
R32 a_217_1051.n1 a_217_1051.t6 14.282
R33 a_217_1051.n1 a_217_1051.t7 14.282
R34 a_217_1051.n5 a_217_1051.t2 14.282
R35 a_217_1051.t5 a_217_1051.n5 14.282
R36 a_217_1051.n5 a_217_1051.n4 12.122
R37 A.n0 A.t0 475.572
R38 A.n2 A.t5 469.145
R39 A.n2 A.t1 384.527
R40 A.n0 A.t3 384.527
R41 A.n3 A.t4 294.278
R42 A.n1 A.t2 294.278
R43 A.n4 A.n1 80.851
R44 A.n4 A.n3 76
R45 A.n1 A.n0 57.842
R46 A.n3 A.n2 56.833
R47 A.n4 A 0.046
R48 a_392_209.n0 a_392_209.t8 512.525
R49 a_392_209.n0 a_392_209.t7 371.139
R50 a_392_209.n1 a_392_209.t9 263.54
R51 a_392_209.n14 a_392_209.n13 216.728
R52 a_392_209.n14 a_392_209.n1 153.043
R53 a_392_209.n16 a_392_209.n14 126.664
R54 a_392_209.n1 a_392_209.n0 120.094
R55 a_392_209.n9 a_392_209.n4 111.94
R56 a_392_209.n9 a_392_209.n8 98.501
R57 a_392_209.n12 a_392_209.n10 80.526
R58 a_392_209.n13 a_392_209.n9 78.403
R59 a_392_209.n16 a_392_209.n15 75.271
R60 a_392_209.n8 a_392_209.n7 30
R61 a_392_209.n12 a_392_209.n11 30
R62 a_392_209.n6 a_392_209.n5 24.383
R63 a_392_209.n8 a_392_209.n6 23.684
R64 a_392_209.n4 a_392_209.n3 22.578
R65 a_392_209.n13 a_392_209.n12 20.417
R66 a_392_209.n15 a_392_209.t0 14.282
R67 a_392_209.n15 a_392_209.t5 14.282
R68 a_392_209.t2 a_392_209.n17 14.282
R69 a_392_209.n17 a_392_209.t1 14.282
R70 a_392_209.n17 a_392_209.n16 12.117
R71 a_392_209.n4 a_392_209.n2 8.58
R72 VDD.n122 VDD.n120 144.705
R73 VDD.n207 VDD.n205 144.705
R74 VDD.n68 VDD.n66 144.705
R75 VDD.n26 VDD.n25 77.792
R76 VDD.n35 VDD.n34 77.792
R77 VDD.n29 VDD.n23 76.145
R78 VDD.n29 VDD.n28 76
R79 VDD.n33 VDD.n32 76
R80 VDD.n39 VDD.n38 76
R81 VDD.n43 VDD.n42 76
R82 VDD.n70 VDD.n69 76
R83 VDD.n74 VDD.n73 76
R84 VDD.n78 VDD.n77 76
R85 VDD.n82 VDD.n81 76
R86 VDD.n86 VDD.n85 76
R87 VDD.n90 VDD.n89 76
R88 VDD.n94 VDD.n93 76
R89 VDD.n98 VDD.n97 76
R90 VDD.n124 VDD.n123 76
R91 VDD.n233 VDD.n232 76
R92 VDD.n229 VDD.n228 76
R93 VDD.n225 VDD.n224 76
R94 VDD.n221 VDD.n220 76
R95 VDD.n217 VDD.n216 76
R96 VDD.n213 VDD.n212 76
R97 VDD.n209 VDD.n208 76
R98 VDD.n182 VDD.n181 76
R99 VDD.n178 VDD.n177 76
R100 VDD.n173 VDD.n172 76
R101 VDD.n168 VDD.n167 76
R102 VDD.n162 VDD.n161 76
R103 VDD.n157 VDD.n156 76
R104 VDD.n152 VDD.n151 76
R105 VDD.n147 VDD.n146 76
R106 VDD.n148 VDD.t4 55.465
R107 VDD.n174 VDD.t2 55.465
R108 VDD.n37 VDD.t0 55.106
R109 VDD.n24 VDD.t1 55.106
R110 VDD.n164 VDD.n163 41.183
R111 VDD.n103 VDD.n102 36.774
R112 VDD.n48 VDD.n47 36.774
R113 VDD.n198 VDD.n197 36.774
R114 VDD.n170 VDD.n169 36.608
R115 VDD.n154 VDD.n153 32.032
R116 VDD.n146 VDD.n143 21.841
R117 VDD.n23 VDD.n20 21.841
R118 VDD.n163 VDD.t3 14.282
R119 VDD.n163 VDD.t5 14.282
R120 VDD.n143 VDD.n126 14.167
R121 VDD.n126 VDD.n125 14.167
R122 VDD.n118 VDD.n100 14.167
R123 VDD.n100 VDD.n99 14.167
R124 VDD.n64 VDD.n45 14.167
R125 VDD.n45 VDD.n44 14.167
R126 VDD.n203 VDD.n184 14.167
R127 VDD.n184 VDD.n183 14.167
R128 VDD.n20 VDD.n19 14.167
R129 VDD.n19 VDD.n17 14.167
R130 VDD.n69 VDD.n65 14.167
R131 VDD.n123 VDD.n119 14.167
R132 VDD.n208 VDD.n204 14.167
R133 VDD.n23 VDD.n22 13.653
R134 VDD.n22 VDD.n21 13.653
R135 VDD.n28 VDD.n27 13.653
R136 VDD.n27 VDD.n26 13.653
R137 VDD.n32 VDD.n31 13.653
R138 VDD.n31 VDD.n30 13.653
R139 VDD.n38 VDD.n36 13.653
R140 VDD.n36 VDD.n35 13.653
R141 VDD.n42 VDD.n41 13.653
R142 VDD.n41 VDD.n40 13.653
R143 VDD.n69 VDD.n68 13.653
R144 VDD.n68 VDD.n67 13.653
R145 VDD.n73 VDD.n72 13.653
R146 VDD.n72 VDD.n71 13.653
R147 VDD.n77 VDD.n76 13.653
R148 VDD.n76 VDD.n75 13.653
R149 VDD.n81 VDD.n80 13.653
R150 VDD.n80 VDD.n79 13.653
R151 VDD.n85 VDD.n84 13.653
R152 VDD.n84 VDD.n83 13.653
R153 VDD.n89 VDD.n88 13.653
R154 VDD.n88 VDD.n87 13.653
R155 VDD.n93 VDD.n92 13.653
R156 VDD.n92 VDD.n91 13.653
R157 VDD.n97 VDD.n96 13.653
R158 VDD.n96 VDD.n95 13.653
R159 VDD.n123 VDD.n122 13.653
R160 VDD.n122 VDD.n121 13.653
R161 VDD.n232 VDD.n231 13.653
R162 VDD.n231 VDD.n230 13.653
R163 VDD.n228 VDD.n227 13.653
R164 VDD.n227 VDD.n226 13.653
R165 VDD.n224 VDD.n223 13.653
R166 VDD.n223 VDD.n222 13.653
R167 VDD.n220 VDD.n219 13.653
R168 VDD.n219 VDD.n218 13.653
R169 VDD.n216 VDD.n215 13.653
R170 VDD.n215 VDD.n214 13.653
R171 VDD.n212 VDD.n211 13.653
R172 VDD.n211 VDD.n210 13.653
R173 VDD.n208 VDD.n207 13.653
R174 VDD.n207 VDD.n206 13.653
R175 VDD.n181 VDD.n180 13.653
R176 VDD.n180 VDD.n179 13.653
R177 VDD.n177 VDD.n176 13.653
R178 VDD.n176 VDD.n175 13.653
R179 VDD.n172 VDD.n171 13.653
R180 VDD.n171 VDD.n170 13.653
R181 VDD.n167 VDD.n166 13.653
R182 VDD.n166 VDD.n165 13.653
R183 VDD.n161 VDD.n160 13.653
R184 VDD.n160 VDD.n159 13.653
R185 VDD.n156 VDD.n155 13.653
R186 VDD.n155 VDD.n154 13.653
R187 VDD.n151 VDD.n150 13.653
R188 VDD.n150 VDD.n149 13.653
R189 VDD.n146 VDD.n145 13.653
R190 VDD.n145 VDD.n144 13.653
R191 VDD.n4 VDD.n2 12.915
R192 VDD.n4 VDD.n3 12.66
R193 VDD.n13 VDD.n12 12.343
R194 VDD.n11 VDD.n10 12.343
R195 VDD.n7 VDD.n6 12.343
R196 VDD.n167 VDD.n164 8.658
R197 VDD.n119 VDD.n118 7.674
R198 VDD.n65 VDD.n64 7.674
R199 VDD.n204 VDD.n203 7.674
R200 VDD.n59 VDD.n58 7.5
R201 VDD.n53 VDD.n52 7.5
R202 VDD.n55 VDD.n54 7.5
R203 VDD.n50 VDD.n49 7.5
R204 VDD.n64 VDD.n63 7.5
R205 VDD.n113 VDD.n112 7.5
R206 VDD.n107 VDD.n106 7.5
R207 VDD.n109 VDD.n108 7.5
R208 VDD.n115 VDD.n105 7.5
R209 VDD.n115 VDD.n103 7.5
R210 VDD.n118 VDD.n117 7.5
R211 VDD.n188 VDD.n187 7.5
R212 VDD.n191 VDD.n190 7.5
R213 VDD.n193 VDD.n192 7.5
R214 VDD.n196 VDD.n195 7.5
R215 VDD.n203 VDD.n202 7.5
R216 VDD.n138 VDD.n137 7.5
R217 VDD.n132 VDD.n131 7.5
R218 VDD.n134 VDD.n133 7.5
R219 VDD.n140 VDD.n130 7.5
R220 VDD.n140 VDD.n128 7.5
R221 VDD.n143 VDD.n142 7.5
R222 VDD.n20 VDD.n16 7.5
R223 VDD.n2 VDD.n1 7.5
R224 VDD.n6 VDD.n5 7.5
R225 VDD.n10 VDD.n9 7.5
R226 VDD.n19 VDD.n18 7.5
R227 VDD.n14 VDD.n0 7.5
R228 VDD.n51 VDD.n48 6.772
R229 VDD.n62 VDD.n46 6.772
R230 VDD.n60 VDD.n57 6.772
R231 VDD.n56 VDD.n53 6.772
R232 VDD.n116 VDD.n101 6.772
R233 VDD.n114 VDD.n111 6.772
R234 VDD.n110 VDD.n107 6.772
R235 VDD.n141 VDD.n127 6.772
R236 VDD.n139 VDD.n136 6.772
R237 VDD.n135 VDD.n132 6.772
R238 VDD.n51 VDD.n50 6.772
R239 VDD.n56 VDD.n55 6.772
R240 VDD.n60 VDD.n59 6.772
R241 VDD.n63 VDD.n62 6.772
R242 VDD.n110 VDD.n109 6.772
R243 VDD.n114 VDD.n113 6.772
R244 VDD.n117 VDD.n116 6.772
R245 VDD.n135 VDD.n134 6.772
R246 VDD.n139 VDD.n138 6.772
R247 VDD.n142 VDD.n141 6.772
R248 VDD.n202 VDD.n201 6.772
R249 VDD.n189 VDD.n186 6.772
R250 VDD.n194 VDD.n191 6.772
R251 VDD.n199 VDD.n196 6.772
R252 VDD.n199 VDD.n198 6.772
R253 VDD.n194 VDD.n193 6.772
R254 VDD.n189 VDD.n188 6.772
R255 VDD.n201 VDD.n185 6.772
R256 VDD.n16 VDD.n15 6.458
R257 VDD.n105 VDD.n104 6.202
R258 VDD.n130 VDD.n129 6.202
R259 VDD.n159 VDD.n158 4.576
R260 VDD.n151 VDD.n148 2.754
R261 VDD.n177 VDD.n174 2.361
R262 VDD.n28 VDD.n24 1.967
R263 VDD.n38 VDD.n37 1.967
R264 VDD.n14 VDD.n7 1.329
R265 VDD.n14 VDD.n8 1.329
R266 VDD.n14 VDD.n11 1.329
R267 VDD.n14 VDD.n13 1.329
R268 VDD.n15 VDD.n14 0.696
R269 VDD.n14 VDD.n4 0.696
R270 VDD.n61 VDD.n60 0.365
R271 VDD.n61 VDD.n56 0.365
R272 VDD.n61 VDD.n51 0.365
R273 VDD.n62 VDD.n61 0.365
R274 VDD.n115 VDD.n114 0.365
R275 VDD.n115 VDD.n110 0.365
R276 VDD.n116 VDD.n115 0.365
R277 VDD.n140 VDD.n139 0.365
R278 VDD.n140 VDD.n135 0.365
R279 VDD.n141 VDD.n140 0.365
R280 VDD.n200 VDD.n199 0.365
R281 VDD.n200 VDD.n194 0.365
R282 VDD.n200 VDD.n189 0.365
R283 VDD.n201 VDD.n200 0.365
R284 VDD.n70 VDD.n43 0.29
R285 VDD.n124 VDD.n98 0.29
R286 VDD.n209 VDD.n182 0.29
R287 VDD.n147 VDD 0.207
R288 VDD.n86 VDD.n82 0.181
R289 VDD.n225 VDD.n221 0.181
R290 VDD.n168 VDD.n162 0.181
R291 VDD.n33 VDD.n29 0.157
R292 VDD.n39 VDD.n33 0.157
R293 VDD.n43 VDD.n39 0.145
R294 VDD.n74 VDD.n70 0.145
R295 VDD.n78 VDD.n74 0.145
R296 VDD.n82 VDD.n78 0.145
R297 VDD.n90 VDD.n86 0.145
R298 VDD.n94 VDD.n90 0.145
R299 VDD.n98 VDD.n94 0.145
R300 VDD.n233 VDD.n229 0.145
R301 VDD.n229 VDD.n225 0.145
R302 VDD.n221 VDD.n217 0.145
R303 VDD.n217 VDD.n213 0.145
R304 VDD.n213 VDD.n209 0.145
R305 VDD.n182 VDD.n178 0.145
R306 VDD.n178 VDD.n173 0.145
R307 VDD.n173 VDD.n168 0.145
R308 VDD.n162 VDD.n157 0.145
R309 VDD.n157 VDD.n152 0.145
R310 VDD.n152 VDD.n147 0.145
R311 VDD VDD.n124 0.078
R312 VDD VDD.n233 0.066
R313 C.n2 C.t3 512.525
R314 C.n0 C.t4 512.525
R315 C.n2 C.t0 371.139
R316 C.n0 C.t1 371.139
R317 C.n3 C.n2 265.439
R318 C.n1 C.n0 265.439
R319 C.n1 C.t2 176.995
R320 C.n3 C.t5 170.569
R321 C.n4 C.n1 77.043
R322 C.n4 C.n3 76
R323 C.n4 C 0.046
R324 Y.n5 Y.n4 232.48
R325 Y.n5 Y.n0 130.543
R326 Y.n6 Y.n5 76
R327 Y.n4 Y.n3 30
R328 Y.n2 Y.n1 24.383
R329 Y.n4 Y.n2 23.684
R330 Y.n0 Y.t1 14.282
R331 Y.n0 Y.t2 14.282
R332 Y.n6 Y 0.046
R333 a_778_101.t0 a_778_101.n0 93.333
R334 a_778_101.n3 a_778_101.n1 55.048
R335 a_778_101.n3 a_778_101.n2 2.097
R336 a_778_101.t0 a_778_101.n3 0.11
R337 GND.n30 GND.n29 219.745
R338 GND.n63 GND.n61 219.745
R339 GND.n100 GND.n99 219.745
R340 GND.n30 GND.n28 85.529
R341 GND.n63 GND.n62 85.529
R342 GND.n100 GND.n98 85.529
R343 GND.n108 GND.n107 84.842
R344 GND.n9 GND.n1 76.145
R345 GND.n70 GND.n69 76
R346 GND.n117 GND.n116 76
R347 GND.n114 GND.n113 76
R348 GND.n111 GND.n110 76
R349 GND.n106 GND.n105 76
R350 GND.n103 GND.n102 76
R351 GND.n96 GND.n95 76
R352 GND.n93 GND.n92 76
R353 GND.n90 GND.n89 76
R354 GND.n87 GND.n86 76
R355 GND.n84 GND.n83 76
R356 GND.n81 GND.n80 76
R357 GND.n73 GND.n72 76
R358 GND.n9 GND.n8 76
R359 GND.n17 GND.n16 76
R360 GND.n24 GND.n23 76
R361 GND.n27 GND.n26 76
R362 GND.n34 GND.n33 76
R363 GND.n37 GND.n36 76
R364 GND.n40 GND.n39 76
R365 GND.n43 GND.n42 76
R366 GND.n46 GND.n45 76
R367 GND.n54 GND.n53 76
R368 GND.n57 GND.n56 76
R369 GND.n60 GND.n59 76
R370 GND.n67 GND.n66 76
R371 GND.n123 GND.n122 76
R372 GND.n120 GND.n119 76
R373 GND.n78 GND.n77 63.835
R374 GND.n51 GND.n50 63.835
R375 GND.n5 GND.n4 35.01
R376 GND.n3 GND.n2 29.127
R377 GND.n77 GND.n76 28.421
R378 GND.n50 GND.n49 28.421
R379 GND.n77 GND.n75 25.263
R380 GND.n50 GND.n48 25.263
R381 GND.n75 GND.n74 24.383
R382 GND.n48 GND.n47 24.383
R383 GND.n12 GND.t0 20.794
R384 GND.n6 GND.n5 19.735
R385 GND.n14 GND.n13 19.735
R386 GND.n21 GND.n20 19.735
R387 GND.n5 GND.n3 19.017
R388 GND.n33 GND.n31 14.167
R389 GND.n66 GND.n64 14.167
R390 GND.n102 GND.n101 14.167
R391 GND.n72 GND.n71 13.653
R392 GND.n80 GND.n79 13.653
R393 GND.n83 GND.n82 13.653
R394 GND.n86 GND.n85 13.653
R395 GND.n89 GND.n88 13.653
R396 GND.n92 GND.n91 13.653
R397 GND.n95 GND.n94 13.653
R398 GND.n102 GND.n97 13.653
R399 GND.n105 GND.n104 13.653
R400 GND.n110 GND.n109 13.653
R401 GND.n113 GND.n112 13.653
R402 GND.n116 GND.n115 13.653
R403 GND.n8 GND.n7 13.653
R404 GND.n16 GND.n15 13.653
R405 GND.n23 GND.n22 13.653
R406 GND.n26 GND.n25 13.653
R407 GND.n33 GND.n32 13.653
R408 GND.n36 GND.n35 13.653
R409 GND.n39 GND.n38 13.653
R410 GND.n42 GND.n41 13.653
R411 GND.n45 GND.n44 13.653
R412 GND.n53 GND.n52 13.653
R413 GND.n56 GND.n55 13.653
R414 GND.n59 GND.n58 13.653
R415 GND.n66 GND.n65 13.653
R416 GND.n122 GND.n121 13.653
R417 GND.n119 GND.n118 13.653
R418 GND.n20 GND.n19 12.837
R419 GND.n19 GND.n18 7.566
R420 GND.n31 GND.n30 7.312
R421 GND.n64 GND.n63 7.312
R422 GND.n101 GND.n100 7.312
R423 GND.n11 GND.n10 4.551
R424 GND.n8 GND.n6 3.935
R425 GND.n53 GND.n51 3.935
R426 GND.n110 GND.n108 3.935
R427 GND.n80 GND.n78 3.935
R428 GND.n23 GND.n21 3.541
R429 GND.t0 GND.n11 2.238
R430 GND.n69 GND.n68 0.596
R431 GND.n1 GND.n0 0.596
R432 GND.n13 GND.n12 0.358
R433 GND.n34 GND.n27 0.29
R434 GND.n67 GND.n60 0.29
R435 GND.n103 GND.n96 0.29
R436 GND.n70 GND 0.207
R437 GND.n16 GND.n14 0.196
R438 GND.n46 GND.n43 0.181
R439 GND.n117 GND.n114 0.181
R440 GND.n87 GND.n84 0.181
R441 GND.n17 GND.n9 0.157
R442 GND.n24 GND.n17 0.157
R443 GND.n27 GND.n24 0.145
R444 GND.n37 GND.n34 0.145
R445 GND.n40 GND.n37 0.145
R446 GND.n43 GND.n40 0.145
R447 GND.n54 GND.n46 0.145
R448 GND.n57 GND.n54 0.145
R449 GND.n60 GND.n57 0.145
R450 GND.n123 GND.n120 0.145
R451 GND.n120 GND.n117 0.145
R452 GND.n114 GND.n111 0.145
R453 GND.n111 GND.n106 0.145
R454 GND.n106 GND.n103 0.145
R455 GND.n96 GND.n93 0.145
R456 GND.n93 GND.n90 0.145
R457 GND.n90 GND.n87 0.145
R458 GND.n84 GND.n81 0.145
R459 GND.n81 GND.n73 0.145
R460 GND.n73 GND.n70 0.145
R461 GND GND.n67 0.078
R462 GND GND.n123 0.066
R463 a_112_101.n1 a_112_101.n0 32.249
R464 a_112_101.t0 a_112_101.n5 7.911
R465 a_112_101.n4 a_112_101.n2 4.032
R466 a_112_101.n4 a_112_101.n3 3.644
R467 a_112_101.t0 a_112_101.n1 2.534
R468 a_112_101.t0 a_112_101.n4 1.099
R469 a_1444_101.t0 a_1444_101.n1 34.62
R470 a_1444_101.t0 a_1444_101.n0 8.137
R471 a_1444_101.t0 a_1444_101.n2 4.69
C7 VDD GND 9.83fF
C8 a_1444_101.n0 GND 0.06fF
C9 a_1444_101.n1 GND 0.14fF
C10 a_1444_101.n2 GND 0.04fF
C11 a_112_101.n0 GND 0.10fF
C12 a_112_101.n1 GND 0.09fF
C13 a_112_101.n2 GND 0.08fF
C14 a_112_101.n3 GND 0.02fF
C15 a_112_101.n4 GND 0.01fF
C16 a_112_101.n5 GND 0.06fF
C17 a_778_101.n0 GND 0.03fF
C18 a_778_101.n1 GND 0.13fF
C19 a_778_101.n2 GND 0.13fF
C20 a_778_101.n3 GND 0.15fF
C21 Y.n0 GND 0.75fF
C22 Y.n1 GND 0.04fF
C23 Y.n2 GND 0.06fF
C24 Y.n3 GND 0.04fF
C25 Y.n4 GND 0.35fF
C26 Y.n5 GND 0.48fF
C27 Y.n6 GND 0.01fF
C28 VDD.n0 GND 0.12fF
C29 VDD.n1 GND 0.02fF
C30 VDD.n2 GND 0.02fF
C31 VDD.n3 GND 0.04fF
C32 VDD.n4 GND 0.01fF
C33 VDD.n5 GND 0.02fF
C34 VDD.n6 GND 0.02fF
C35 VDD.n9 GND 0.02fF
C36 VDD.n10 GND 0.02fF
C37 VDD.n12 GND 0.02fF
C38 VDD.n14 GND 0.45fF
C39 VDD.n16 GND 0.03fF
C40 VDD.n17 GND 0.02fF
C41 VDD.n18 GND 0.02fF
C42 VDD.n19 GND 0.02fF
C43 VDD.n20 GND 0.03fF
C44 VDD.n21 GND 0.27fF
C45 VDD.n22 GND 0.02fF
C46 VDD.n23 GND 0.03fF
C47 VDD.n24 GND 0.06fF
C48 VDD.n25 GND 0.14fF
C49 VDD.n26 GND 0.20fF
C50 VDD.n27 GND 0.01fF
C51 VDD.n28 GND 0.01fF
C52 VDD.n29 GND 0.07fF
C53 VDD.n30 GND 0.16fF
C54 VDD.n31 GND 0.01fF
C55 VDD.n32 GND 0.02fF
C56 VDD.n33 GND 0.02fF
C57 VDD.n34 GND 0.14fF
C58 VDD.n35 GND 0.20fF
C59 VDD.n36 GND 0.01fF
C60 VDD.n37 GND 0.06fF
C61 VDD.n38 GND 0.01fF
C62 VDD.n39 GND 0.02fF
C63 VDD.n40 GND 0.27fF
C64 VDD.n41 GND 0.01fF
C65 VDD.n42 GND 0.02fF
C66 VDD.n43 GND 0.03fF
C67 VDD.n44 GND 0.02fF
C68 VDD.n45 GND 0.02fF
C69 VDD.n46 GND 0.02fF
C70 VDD.n47 GND 0.18fF
C71 VDD.n48 GND 0.04fF
C72 VDD.n49 GND 0.03fF
C73 VDD.n50 GND 0.02fF
C74 VDD.n52 GND 0.02fF
C75 VDD.n53 GND 0.02fF
C76 VDD.n54 GND 0.02fF
C77 VDD.n55 GND 0.02fF
C78 VDD.n57 GND 0.02fF
C79 VDD.n58 GND 0.02fF
C80 VDD.n59 GND 0.02fF
C81 VDD.n61 GND 0.27fF
C82 VDD.n63 GND 0.02fF
C83 VDD.n64 GND 0.02fF
C84 VDD.n65 GND 0.03fF
C85 VDD.n66 GND 0.02fF
C86 VDD.n67 GND 0.27fF
C87 VDD.n68 GND 0.01fF
C88 VDD.n69 GND 0.02fF
C89 VDD.n70 GND 0.03fF
C90 VDD.n71 GND 0.27fF
C91 VDD.n72 GND 0.01fF
C92 VDD.n73 GND 0.02fF
C93 VDD.n74 GND 0.02fF
C94 VDD.n75 GND 0.27fF
C95 VDD.n76 GND 0.01fF
C96 VDD.n77 GND 0.02fF
C97 VDD.n78 GND 0.02fF
C98 VDD.n79 GND 0.30fF
C99 VDD.n80 GND 0.01fF
C100 VDD.n81 GND 0.03fF
C101 VDD.n82 GND 0.03fF
C102 VDD.n83 GND 0.30fF
C103 VDD.n84 GND 0.01fF
C104 VDD.n85 GND 0.03fF
C105 VDD.n86 GND 0.03fF
C106 VDD.n87 GND 0.27fF
C107 VDD.n88 GND 0.01fF
C108 VDD.n89 GND 0.02fF
C109 VDD.n90 GND 0.02fF
C110 VDD.n91 GND 0.27fF
C111 VDD.n92 GND 0.01fF
C112 VDD.n93 GND 0.02fF
C113 VDD.n94 GND 0.02fF
C114 VDD.n95 GND 0.27fF
C115 VDD.n96 GND 0.01fF
C116 VDD.n97 GND 0.02fF
C117 VDD.n98 GND 0.03fF
C118 VDD.n99 GND 0.02fF
C119 VDD.n100 GND 0.02fF
C120 VDD.n101 GND 0.02fF
C121 VDD.n102 GND 0.21fF
C122 VDD.n103 GND 0.04fF
C123 VDD.n104 GND 0.03fF
C124 VDD.n105 GND 0.02fF
C125 VDD.n106 GND 0.02fF
C126 VDD.n107 GND 0.02fF
C127 VDD.n108 GND 0.02fF
C128 VDD.n109 GND 0.02fF
C129 VDD.n111 GND 0.02fF
C130 VDD.n112 GND 0.02fF
C131 VDD.n113 GND 0.02fF
C132 VDD.n115 GND 0.27fF
C133 VDD.n117 GND 0.02fF
C134 VDD.n118 GND 0.02fF
C135 VDD.n119 GND 0.03fF
C136 VDD.n120 GND 0.02fF
C137 VDD.n121 GND 0.27fF
C138 VDD.n122 GND 0.01fF
C139 VDD.n123 GND 0.02fF
C140 VDD.n124 GND 0.03fF
C141 VDD.n125 GND 0.02fF
C142 VDD.n126 GND 0.02fF
C143 VDD.n127 GND 0.02fF
C144 VDD.n128 GND 0.15fF
C145 VDD.n129 GND 0.03fF
C146 VDD.n130 GND 0.02fF
C147 VDD.n131 GND 0.02fF
C148 VDD.n132 GND 0.02fF
C149 VDD.n133 GND 0.02fF
C150 VDD.n134 GND 0.02fF
C151 VDD.n136 GND 0.02fF
C152 VDD.n137 GND 0.02fF
C153 VDD.n138 GND 0.02fF
C154 VDD.n140 GND 0.45fF
C155 VDD.n142 GND 0.03fF
C156 VDD.n143 GND 0.03fF
C157 VDD.n144 GND 0.27fF
C158 VDD.n145 GND 0.02fF
C159 VDD.n146 GND 0.03fF
C160 VDD.n147 GND 0.03fF
C161 VDD.n148 GND 0.06fF
C162 VDD.n149 GND 0.24fF
C163 VDD.n150 GND 0.01fF
C164 VDD.n151 GND 0.01fF
C165 VDD.n152 GND 0.02fF
C166 VDD.n153 GND 0.13fF
C167 VDD.n154 GND 0.16fF
C168 VDD.n155 GND 0.01fF
C169 VDD.n156 GND 0.02fF
C170 VDD.n157 GND 0.02fF
C171 VDD.n158 GND 0.17fF
C172 VDD.n159 GND 0.14fF
C173 VDD.n160 GND 0.01fF
C174 VDD.n161 GND 0.02fF
C175 VDD.n162 GND 0.03fF
C176 VDD.n163 GND 0.10fF
C177 VDD.n164 GND 0.02fF
C178 VDD.n165 GND 0.30fF
C179 VDD.n166 GND 0.01fF
C180 VDD.n167 GND 0.02fF
C181 VDD.n168 GND 0.03fF
C182 VDD.n169 GND 0.13fF
C183 VDD.n170 GND 0.16fF
C184 VDD.n171 GND 0.01fF
C185 VDD.n172 GND 0.02fF
C186 VDD.n173 GND 0.02fF
C187 VDD.n174 GND 0.06fF
C188 VDD.n175 GND 0.24fF
C189 VDD.n176 GND 0.01fF
C190 VDD.n177 GND 0.01fF
C191 VDD.n178 GND 0.02fF
C192 VDD.n179 GND 0.27fF
C193 VDD.n180 GND 0.01fF
C194 VDD.n181 GND 0.02fF
C195 VDD.n182 GND 0.03fF
C196 VDD.n183 GND 0.02fF
C197 VDD.n184 GND 0.02fF
C198 VDD.n185 GND 0.02fF
C199 VDD.n186 GND 0.02fF
C200 VDD.n187 GND 0.02fF
C201 VDD.n188 GND 0.02fF
C202 VDD.n190 GND 0.02fF
C203 VDD.n191 GND 0.02fF
C204 VDD.n192 GND 0.02fF
C205 VDD.n193 GND 0.02fF
C206 VDD.n195 GND 0.03fF
C207 VDD.n196 GND 0.02fF
C208 VDD.n197 GND 0.21fF
C209 VDD.n198 GND 0.04fF
C210 VDD.n200 GND 0.27fF
C211 VDD.n202 GND 0.02fF
C212 VDD.n203 GND 0.02fF
C213 VDD.n204 GND 0.03fF
C214 VDD.n205 GND 0.02fF
C215 VDD.n206 GND 0.27fF
C216 VDD.n207 GND 0.01fF
C217 VDD.n208 GND 0.02fF
C218 VDD.n209 GND 0.03fF
C219 VDD.n210 GND 0.27fF
C220 VDD.n211 GND 0.01fF
C221 VDD.n212 GND 0.02fF
C222 VDD.n213 GND 0.02fF
C223 VDD.n214 GND 0.27fF
C224 VDD.n215 GND 0.01fF
C225 VDD.n216 GND 0.02fF
C226 VDD.n217 GND 0.02fF
C227 VDD.n218 GND 0.30fF
C228 VDD.n219 GND 0.01fF
C229 VDD.n220 GND 0.03fF
C230 VDD.n221 GND 0.03fF
C231 VDD.n222 GND 0.30fF
C232 VDD.n223 GND 0.01fF
C233 VDD.n224 GND 0.03fF
C234 VDD.n225 GND 0.03fF
C235 VDD.n226 GND 0.27fF
C236 VDD.n227 GND 0.01fF
C237 VDD.n228 GND 0.02fF
C238 VDD.n229 GND 0.02fF
C239 VDD.n230 GND 0.27fF
C240 VDD.n231 GND 0.01fF
C241 VDD.n232 GND 0.02fF
C242 VDD.n233 GND 0.02fF
C243 a_392_209.n0 GND 0.25fF
C244 a_392_209.n1 GND 0.47fF
C245 a_392_209.n2 GND 0.03fF
C246 a_392_209.n3 GND 0.04fF
C247 a_392_209.n4 GND 0.09fF
C248 a_392_209.n5 GND 0.03fF
C249 a_392_209.n6 GND 0.04fF
C250 a_392_209.n7 GND 0.03fF
C251 a_392_209.n8 GND 0.09fF
C252 a_392_209.n9 GND 0.95fF
C253 a_392_209.n10 GND 0.05fF
C254 a_392_209.n11 GND 0.03fF
C255 a_392_209.n12 GND 0.07fF
C256 a_392_209.n13 GND 0.25fF
C257 a_392_209.n14 GND 0.44fF
C258 a_392_209.n15 GND 0.45fF
C259 a_392_209.n16 GND 0.22fF
C260 a_392_209.n17 GND 0.37fF
C261 a_217_1051.n0 GND 0.36fF
C262 a_217_1051.n1 GND 0.40fF
C263 a_217_1051.n2 GND 0.28fF
C264 a_217_1051.n3 GND 0.62fF
C265 a_217_1051.n4 GND 0.23fF
C266 a_217_1051.n5 GND 0.32fF
C267 a_881_1051.n0 GND 0.29fF
C268 a_881_1051.n1 GND 0.28fF
C269 a_881_1051.n2 GND 0.35fF
C270 a_881_1051.n3 GND 0.25fF
C271 a_881_1051.n4 GND 0.57fF
C272 a_881_1051.n5 GND 0.20fF
.ends
