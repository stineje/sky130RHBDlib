* SPICE3 file created from TIEHI.ext - technology: sky130A

.subckt TIEHI Y VPB VNB
X0 VPB a_121_383# a_193_1004# VPB sky130_fd_pr__pfet_01v8 ad=1.1e+12p pd=9.1e+06u as=0p ps=0u w=2e+06u l=150000u M=2
X1 a_121_383# a_121_383# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.1408e+12p ps=8.1e+06u w=3e+06u l=150000u
.ends
