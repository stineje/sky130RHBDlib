magic
tech sky130A
magscale 1 2
timestamp 1652326224
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 797 945 831 979
rect 205 871 239 905
rect 427 871 461 905
rect 649 871 683 905
rect 797 871 831 905
rect 205 797 239 831
rect 427 797 461 831
rect 649 797 683 831
rect 797 797 831 831
rect 205 723 239 757
rect 427 723 461 757
rect 649 723 683 757
rect 797 723 831 757
rect 205 649 239 683
rect 427 649 461 683
rect 649 649 683 683
rect 797 649 831 683
rect 205 575 239 609
rect 427 575 461 609
rect 649 575 683 609
rect 797 575 831 609
rect 205 501 239 535
rect 427 501 461 535
rect 649 501 683 535
rect 797 501 831 535
rect 205 427 239 461
rect 427 427 461 461
rect 649 427 683 461
rect 797 427 831 461
<< metal1 >>
rect -34 1446 996 1514
rect -34 -34 996 34
use nand3x1_pcell  nand3x1_pcell_0 pcells
timestamp 1652319931
transform 1 0 0 0 1 0
box -87 -34 1049 1550
<< labels >>
rlabel locali 797 427 831 461 1 Y
port 1 nsew signal output
rlabel locali 797 501 831 535 1 Y
port 1 nsew signal output
rlabel locali 797 575 831 609 1 Y
port 1 nsew signal output
rlabel locali 797 649 831 683 1 Y
port 1 nsew signal output
rlabel locali 797 723 831 757 1 Y
port 1 nsew signal output
rlabel locali 797 871 831 905 1 Y
port 1 nsew signal output
rlabel locali 797 945 831 979 1 Y
port 1 nsew signal output
rlabel locali 797 797 831 831 1 Y
port 1 nsew signal output
rlabel locali 205 575 239 609 1 A
port 2 nsew signal input
rlabel locali 205 501 239 535 1 A
port 2 nsew signal input
rlabel locali 205 427 239 461 1 A
port 2 nsew signal input
rlabel locali 205 649 239 683 1 A
port 2 nsew signal input
rlabel locali 205 723 239 757 1 A
port 2 nsew signal input
rlabel locali 205 797 239 831 1 A
port 2 nsew signal input
rlabel locali 205 871 239 905 1 A
port 2 nsew signal input
rlabel locali 427 649 461 683 1 B
port 3 nsew signal input
rlabel locali 427 723 461 757 1 B
port 3 nsew signal input
rlabel locali 427 797 461 831 1 B
port 3 nsew signal input
rlabel locali 427 871 461 905 1 B
port 3 nsew signal input
rlabel locali 427 575 461 609 1 B
port 3 nsew signal input
rlabel locali 427 501 461 535 1 B
port 3 nsew signal input
rlabel locali 427 427 461 461 1 B
port 3 nsew signal input
rlabel locali 649 575 683 609 1 C
port 4 nsew signal input
rlabel locali 649 501 683 535 1 C
port 4 nsew signal input
rlabel locali 649 427 683 461 1 C
port 4 nsew signal input
rlabel locali 649 649 683 683 1 C
port 4 nsew signal input
rlabel locali 649 723 683 757 1 C
port 4 nsew signal input
rlabel locali 649 797 683 831 1 C
port 4 nsew signal input
rlabel locali 649 871 683 905 1 C
port 4 nsew signal input
rlabel metal1 -34 1446 996 1514 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 -34 -34 996 34 1 VGND
port 6 nsew ground bidirectional abutment
rlabel nwell 57 1463 91 1497 1 VPB
port 6 nsew power bidirectional
rlabel pwell 57 -17 91 17 1 VNB
port 6 nsew ground bidirectional
<< properties >>                                                                
string LEFsite unithd                                                           
string LEFclass CORE
string LEFsymmetry X Y R90
<< end >>
