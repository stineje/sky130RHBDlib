VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOR2X1
  CLASS CORE ;
  FOREIGN NOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.330 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.963050 ;
    PORT
      LAYER li1 ;
        RECT 2.025 5.295 2.195 6.565 ;
        RECT 2.025 5.125 2.675 5.295 ;
        RECT 2.505 1.740 2.675 5.125 ;
        RECT 1.095 1.570 2.675 1.740 ;
        RECT 1.095 0.835 1.265 1.570 ;
        RECT 2.065 0.835 2.235 1.570 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 0.870 4.710 1.040 4.870 ;
        RECT 0.870 4.540 1.195 4.710 ;
        RECT 1.025 1.915 1.195 4.540 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.026450 ;
    PORT
      LAYER li1 ;
        RECT 1.800 4.710 1.970 4.870 ;
        RECT 1.765 4.540 1.970 4.710 ;
        RECT 1.765 1.915 1.935 4.540 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 3.765 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 3.500 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 1.145 5.555 1.315 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 3.500 7.570 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 3.500 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 0.610 0.615 0.780 1.745 ;
        RECT 1.580 0.615 1.750 1.390 ;
        RECT 2.550 0.615 2.720 1.390 ;
        RECT 0.610 0.445 2.720 0.615 ;
        RECT 0.610 0.170 0.780 0.445 ;
        RECT 1.095 0.170 1.265 0.445 ;
        RECT 1.580 0.170 1.750 0.445 ;
        RECT 2.065 0.170 2.235 0.445 ;
        RECT 2.550 0.170 2.720 0.445 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT -0.170 -0.170 3.500 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 3.500 0.170 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 0.705 5.295 0.875 7.025 ;
        RECT 1.585 6.825 2.635 6.995 ;
        RECT 1.585 5.295 1.755 6.825 ;
        RECT 2.465 5.555 2.635 6.825 ;
        RECT 0.705 5.125 1.755 5.295 ;
  END
END NOR2X1
END LIBRARY

