* SPICE3 file created from tmp.ext - technology: sky130A

.subckt tmp Y A B VDD VSS
X0 Y or2x1_pcell_0/m1_547_649 VSS VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=3.07743p ps=2.1045u w=3u l=0.15u
X1 VDD or2x1_pcell_0/m1_547_649 Y VDD sky130_fd_pr__pfet_01v8 ad=5.4545p pd=1.369u as=-4.325p ps=4.585u w=2u l=0.15u M=2
X2 VDD A or2x1_pcell_0/nor2x1_pcell_0/a_317_1377 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X3 or2x1_pcell_0/m1_547_649 B or2x1_pcell_0/nor2x1_pcell_0/a_317_1377 VDD sky130_fd_pr__pfet_01v8 ad=-0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X4 or2x1_pcell_0/m1_547_649 A VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X5 or2x1_pcell_0/m1_547_649 B VSS VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
C0 VDD VSS 2.58fF
.ends
