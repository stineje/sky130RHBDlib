magic
tech sky130A
magscale 1 2
timestamp 1652453496
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 131 871 165 905
rect 575 871 609 905
rect 2351 871 2385 905
rect 3609 871 3643 905
rect 3979 871 4013 905
rect 131 797 165 831
rect 575 797 609 831
rect 2351 797 2385 831
rect 131 723 165 757
rect 575 723 609 757
rect 131 649 165 683
rect 575 649 609 683
rect 2351 649 2385 683
rect 3609 649 3643 683
rect 3979 649 4013 683
rect 131 575 165 609
rect 2351 575 2385 609
rect 3609 575 3643 609
rect 3979 575 4013 609
rect 131 501 165 535
rect 575 501 609 535
rect 2351 501 2385 535
rect 3609 501 3643 535
rect 3979 501 4013 535
rect 3609 427 3643 461
rect 3979 427 4013 461
<< metal1 >>
rect -34 1446 4474 1514
rect 645 797 2315 831
rect 3013 797 4091 831
rect 793 723 1057 757
rect 1903 723 3277 757
rect 3531 723 4239 757
rect 3679 649 3943 683
rect 349 575 2167 609
rect -34 -34 4474 34
use li1_M1_contact  li1_M1_contact_14 pcells
timestamp 1648061256
transform -1 0 296 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform -1 0 592 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 740 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform -1 0 1850 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform 1 0 1110 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 1258 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform -1 0 2960 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 3330 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 2220 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform 1 0 2368 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform 1 0 3996 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform -1 0 3478 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform -1 0 3626 0 -1 666
box -53 -33 29 33
use invx1_pcell  invx1_pcell_1 pcells
timestamp 1652329846
transform 1 0 0 0 1 0
box -87 -34 531 1550
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform 1 0 4292 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 4144 0 1 814
box -53 -33 29 33
use nor2x1_pcell  nor2x1_pcell_0 pcells
timestamp 1652323563
transform 1 0 3108 0 1 0
box -87 -34 753 1550
use nor2x1_pcell  nor2x1_pcell_1
timestamp 1652323563
transform 1 0 3774 0 1 0
box -87 -34 753 1550
use and2x1_pcell  and2x1_pcell_1 pcells
timestamp 1652453496
transform 1 0 1998 0 1 0
box -87 -34 1197 1550
use invx1_pcell  invx1_pcell_0
timestamp 1652329846
transform 1 0 444 0 1 0
box -87 -34 531 1550
use and2x1_pcell  and2x1_pcell_0
timestamp 1652453496
transform 1 0 888 0 1 0
box -87 -34 1197 1550
<< labels >>
rlabel locali 3609 649 3643 683 1 Q
port 1 nsew signal output
rlabel locali 3609 575 3643 609 1 Q
port 1 nsew signal output
rlabel locali 3609 501 3643 535 1 Q
port 1 nsew signal output
rlabel locali 3609 427 3643 461 1 Q
port 1 nsew signal output
rlabel locali 3609 871 3643 905 1 Q
port 1 nsew signal output
rlabel locali 3979 427 4013 461 1 Q
port 1 nsew signal output
rlabel locali 3979 501 4013 535 1 Q
port 1 nsew signal output
rlabel locali 3979 575 4013 609 1 Q
port 1 nsew signal output
rlabel locali 3979 649 4013 683 1 Q
port 1 nsew signal output
rlabel locali 3979 871 4013 905 1 Q
port 1 nsew signal output
rlabel locali 575 797 609 831 1 D
port 2 nsew signal input
rlabel locali 575 871 609 905 1 D
port 2 nsew signal input
rlabel locali 575 723 609 757 1 D
port 2 nsew signal input
rlabel locali 575 649 609 683 1 D
port 2 nsew signal input
rlabel locali 575 501 609 535 1 D
port 2 nsew signal input
rlabel locali 2351 649 2385 683 1 D
port 2 nsew signal input
rlabel locali 2351 797 2385 831 1 D
port 2 nsew signal input
rlabel locali 2351 871 2385 905 1 D
port 2 nsew signal input
rlabel locali 2351 575 2385 609 1 D
port 2 nsew signal input
rlabel locali 2351 501 2385 535 1 D
port 2 nsew signal input
rlabel locali 131 575 165 609 1 GATE_N
port 3 nsew signal input
rlabel locali 131 501 165 535 1 GATE_N
port 3 nsew signal input
rlabel locali 131 649 165 683 1 GATE_N
port 3 nsew signal input
rlabel locali 131 723 165 757 1 GATE_N
port 3 nsew signal input
rlabel locali 131 797 165 831 1 GATE_N
port 3 nsew signal input
rlabel locali 131 871 165 905 1 GATE_N
port 3 nsew signal input
rlabel metal1 -34 1446 4474 1514 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 -34 -34 4474 34 1 GND
port 5 nsew ground bidirectional abutment


<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 4440 1480
string LEFsymmetry X Y R90
<< end >>
