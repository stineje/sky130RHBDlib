// File: nand2x1_pcell.spi.pex
// Created: Tue Oct 15 15:57:39 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_NAND2X1_PCELL\%noxref_2 ( 7 19 27 42 45 46 47 48 )
c35 ( 48 0 ) capacitor c=0.0383753f //x=2.405 //y=5.02
c36 ( 47 0 ) capacitor c=0.0243052f //x=1.525 //y=5.02
c37 ( 46 0 ) capacitor c=0.053196f //x=0.655 //y=5.02
c38 ( 45 0 ) capacitor c=0.243792f //x=2.59 //y=7.4
c39 ( 43 0 ) capacitor c=0.00591168f //x=1.67 //y=7.4
c40 ( 42 0 ) capacitor c=0.24846f //x=0.74 //y=7.4
c41 ( 27 0 ) capacitor c=0.0285035f //x=2.465 //y=7.4
c42 ( 19 0 ) capacitor c=0.0286367f //x=1.585 //y=7.4
c43 ( 7 0 ) capacitor c=0.153489f //x=2.59 //y=7.4
r44 (  31 45 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.55 //y=7.23 //x2=2.55 //y2=7.4
r45 (  31 48 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=6.745
r46 (  28 43 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.67 //y2=7.4
r47 (  28 30 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.85 //y2=7.4
r48 (  27 45 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=2.55 //y2=7.4
r49 (  27 30 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=1.85 //y2=7.4
r50 (  21 43 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.67 //y=7.23 //x2=1.67 //y2=7.4
r51 (  21 47 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=6.745
r52 (  20 42 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.875 //y=7.4 //x2=0.79 //y2=7.4
r53 (  19 43 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=1.67 //y2=7.4
r54 (  19 20 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=0.875 //y2=7.4
r55 (  13 42 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=0.79 //y=7.23 //x2=0.79 //y2=7.4
r56 (  13 46 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=6.405
r57 (  7 45 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=2.59 //y=7.4 //x2=2.59 //y2=7.4
r58 (  5 30 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=1.85 \
 //y=7.4 //x2=1.85 //y2=7.4
r59 (  5 7 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.59 //y2=7.4
r60 (  2 42 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=0.74 \
 //y=7.4 //x2=0.74 //y2=7.4
r61 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_NAND2X1_PCELL\%noxref_2

subckt PM_NAND2X1_PCELL\%noxref_3 ( 2 7 8 9 10 11 12 13 17 19 22 23 33 )
c53 ( 33 0 ) capacitor c=0.0667949f //x=1.11 //y=4.7
c54 ( 23 0 ) capacitor c=0.0318948f //x=1.445 //y=1.21
c55 ( 22 0 ) capacitor c=0.0187384f //x=1.445 //y=0.865
c56 ( 19 0 ) capacitor c=0.0141798f //x=1.29 //y=1.365
c57 ( 17 0 ) capacitor c=0.0149844f //x=1.29 //y=0.71
c58 ( 13 0 ) capacitor c=0.0860049f //x=0.915 //y=1.915
c59 ( 12 0 ) capacitor c=0.0229722f //x=0.915 //y=1.52
c60 ( 11 0 ) capacitor c=0.0234352f //x=0.915 //y=1.21
c61 ( 10 0 ) capacitor c=0.0199343f //x=0.915 //y=0.865
c62 ( 9 0 ) capacitor c=0.110275f //x=1.45 //y=6.02
c63 ( 8 0 ) capacitor c=0.154305f //x=1.01 //y=6.02
c64 ( 2 0 ) capacitor c=0.116968f //x=1.11 //y=2.08
r65 (  31 33 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.7 //x2=1.11 //y2=4.7
r66 (  24 33 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=1.45 //y=4.865 //x2=1.11 //y2=4.7
r67 (  23 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.21 //x2=1.405 //y2=1.365
r68 (  22 34 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.405 //y2=0.71
r69 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.445 //y2=1.21
r70 (  20 30 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.365 //x2=0.955 //y2=1.365
r71 (  19 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.365 //x2=1.405 //y2=1.365
r72 (  18 29 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.71 //x2=0.955 //y2=0.71
r73 (  17 34 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.405 //y2=0.71
r74 (  17 18 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.07 //y2=0.71
r75 (  14 31 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.865 //x2=1.01 //y2=4.7
r76 (  13 28 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r77 (  12 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.955 //y2=1.365
r78 (  12 13 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.915 //y2=1.915
r79 (  11 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.21 //x2=0.955 //y2=1.365
r80 (  10 29 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.955 //y2=0.71
r81 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.915 //y2=1.21
r82 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.02 //x2=1.45 //y2=4.865
r83 (  8 14 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.02 //x2=1.01 //y2=4.865
r84 (  7 19 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.29 //y2=1.365
r85 (  7 20 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.07 //y2=1.365
r86 (  5 33 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r87 (  2 28 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r88 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=4.7
ends PM_NAND2X1_PCELL\%noxref_3

subckt PM_NAND2X1_PCELL\%noxref_4 ( 1 3 7 8 9 10 11 12 17 19 21 27 28 30 31 34 )
c61 ( 34 0 ) capacitor c=0.034715f //x=1.88 //y=4.7
c62 ( 31 0 ) capacitor c=0.0279499f //x=1.85 //y=1.915
c63 ( 30 0 ) capacitor c=0.0437302f //x=1.85 //y=2.08
c64 ( 28 0 ) capacitor c=0.0429696f //x=2.415 //y=1.25
c65 ( 27 0 ) capacitor c=0.0192208f //x=2.415 //y=0.905
c66 ( 21 0 ) capacitor c=0.0158629f //x=2.26 //y=1.405
c67 ( 19 0 ) capacitor c=0.0157803f //x=2.26 //y=0.75
c68 ( 17 0 ) capacitor c=0.0366192f //x=2.255 //y=4.79
c69 ( 12 0 ) capacitor c=0.0205163f //x=1.885 //y=1.56
c70 ( 11 0 ) capacitor c=0.0168481f //x=1.885 //y=1.25
c71 ( 10 0 ) capacitor c=0.0174783f //x=1.885 //y=0.905
c72 ( 9 0 ) capacitor c=0.15358f //x=2.33 //y=6.02
c73 ( 8 0 ) capacitor c=0.110281f //x=1.89 //y=6.02
c74 ( 3 0 ) capacitor c=0.0822126f //x=1.85 //y=2.08
c75 ( 1 0 ) capacitor c=0.00453889f //x=1.85 //y=4.535
r76 (  36 37 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.79 //x2=1.88 //y2=4.865
r77 (  34 36 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.7 //x2=1.88 //y2=4.79
r78 (  30 31 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r79 (  28 41 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.25 //x2=2.375 //y2=1.405
r80 (  27 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r81 (  27 28 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.25
r82 (  22 39 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r83 (  21 41 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.375 //y2=1.405
r84 (  20 38 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r85 (  19 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r86 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r87 (  18 36 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.015 //y=4.79 //x2=1.88 //y2=4.79
r88 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.33 //y2=4.865
r89 (  17 18 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.015 //y2=4.79
r90 (  12 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r91 (  12 31 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r92 (  11 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.25 //x2=1.925 //y2=1.405
r93 (  10 38 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r94 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.25
r95 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.02 //x2=2.33 //y2=4.865
r96 (  8 37 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.02 //x2=1.89 //y2=4.865
r97 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r98 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r99 (  6 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.88 //y=4.7 //x2=1.88 //y2=4.7
r100 (  3 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r101 (  1 6 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.865 //y2=4.7
r102 (  1 3 ) resistor r=168.043 //w=0.187 //l=2.455 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.85 //y2=2.08
ends PM_NAND2X1_PCELL\%noxref_4

subckt PM_NAND2X1_PCELL\%noxref_5 ( 7 8 19 21 22 24 25 26 28 29 )
c57 ( 29 0 ) capacitor c=0.0220291f //x=1.965 //y=5.02
c58 ( 28 0 ) capacitor c=0.0217503f //x=1.085 //y=5.02
c59 ( 26 0 ) capacitor c=0.0084702f //x=1.96 //y=0.905
c60 ( 25 0 ) capacitor c=0.00427536f //x=2.11 //y=5.2
c61 ( 24 0 ) capacitor c=0.133595f //x=2.59 //y=5.115
c62 ( 22 0 ) capacitor c=0.00781917f //x=2.235 //y=1.655
c63 ( 21 0 ) capacitor c=0.0167625f //x=2.505 //y=1.655
c64 ( 19 0 ) capacitor c=0.017841f //x=2.505 //y=5.2
c65 ( 8 0 ) capacitor c=0.00387264f //x=1.315 //y=5.2
c66 ( 7 0 ) capacitor c=0.0222171f //x=2.025 //y=5.2
r67 (  23 24 ) resistor r=231.016 //w=0.187 //l=3.375 //layer=li \
 //thickness=0.1 //x=2.59 //y=1.74 //x2=2.59 //y2=5.115
r68 (  21 23 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.59 //y2=1.74
r69 (  21 22 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.235 //y2=1.655
r70 (  20 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.195 //y=5.2 //x2=2.11 //y2=5.2
r71 (  19 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.59 //y2=5.115
r72 (  19 20 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.195 //y2=5.2
r73 (  15 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.235 //y2=1.655
r74 (  15 26 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r75 (  9 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.11 //y=5.285 //x2=2.11 //y2=5.2
r76 (  9 29 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li //thickness=0.1 \
 //x=2.11 //y=5.285 //x2=2.11 //y2=5.725
r77 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.025 //y=5.2 //x2=2.11 //y2=5.2
r78 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=2.025 //y=5.2 //x2=1.315 //y2=5.2
r79 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.315 //y2=5.2
r80 (  1 28 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li //thickness=0.1 \
 //x=1.23 //y=5.285 //x2=1.23 //y2=5.725
ends PM_NAND2X1_PCELL\%noxref_5

subckt PM_NAND2X1_PCELL\%noxref_6 ( 1 5 9 10 13 17 29 )
c31 ( 29 0 ) capacitor c=0.0642544f //x=0.56 //y=0.365
c32 ( 17 0 ) capacitor c=0.00722223f //x=2.635 //y=0.615
c33 ( 13 0 ) capacitor c=0.0154622f //x=2.55 //y=0.53
c34 ( 10 0 ) capacitor c=0.0092508f //x=1.665 //y=1.495
c35 ( 9 0 ) capacitor c=0.006761f //x=1.665 //y=0.615
c36 ( 5 0 ) capacitor c=0.0255599f //x=1.58 //y=1.58
c37 ( 1 0 ) capacitor c=0.0113547f //x=0.695 //y=1.495
r38 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.49
r39 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r40 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.75 //y=0.53 //x2=1.665 //y2=0.49
r41 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=2.15 //y2=0.53
r42 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.49
r43 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.55 //y=0.53 //x2=2.15 //y2=0.53
r44 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=1.62
r45 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=0.88
r46 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.49
r47 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r48 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.78 //y=1.58 //x2=0.695 //y2=1.62
r49 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.78 //y=1.58 //x2=1.18 //y2=1.58
r50 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.58 //y=1.58 //x2=1.665 //y2=1.62
r51 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.58 //y=1.58 //x2=1.18 //y2=1.58
r52 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.695 //y=1.495 //x2=0.695 //y2=1.62
r53 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.695 //y=1.495 //x2=0.695 //y2=0.88
ends PM_NAND2X1_PCELL\%noxref_6

