* SPICE3 file created from NAND3X1.ext - technology: sky130A

.subckt NAND3X1 Y A B C VPB VNB
X0 VPB a_342_166# a_277_1004# VPB sky130_fd_pr__pfet_01v8 ad=2.26e+12p pd=1.826e+07u as=0p ps=0u w=2e+06u l=150000u M=2
X1 VNB a_147_159# a_91_75# VNB sky130_fd_pr__nfet_01v8 ad=1.791e+11p pd=1.57e+06u as=0p ps=0u w=3e+06u l=150000u
X2 VPB a_599_943# a_277_1004# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X3 a_372_182# a_342_166# a_91_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X4 a_277_1004# a_147_159# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X5 a_277_1004# a_599_943# a_372_182# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
.ends
