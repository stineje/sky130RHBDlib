* SPICE3 file created from DFFSNQNX1.ext - technology: sky130A

.subckt DFFSNQNX1 QN D CLK SN VDD GND
M1000 a_3599_411.t4 QN.t5 VDD.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_343_411.t4 a_1265_989.t5 VDD.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t3 SN.t1 a_1905_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_1265_989.t4 CLK.t0 VDD.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VDD.t19 a_343_411.t7 QN.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_3599_411.t2 SN.t2 VDD.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 GND a_217_1050.t6 a_757_103.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1007 GND D.t1 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1008 GND a_343_411.t8 a_3368_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1009 VDD.t11 D.t0 a_217_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VDD.t0 a_1265_989.t7 a_1905_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_3599_411.t0 a_1265_989.t8 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1905_1050.t4 a_217_1050.t5 VDD.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VDD.t13 a_343_411.t9 a_217_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t2 a_217_1050.t7 a_343_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 GND a_217_1050.t8 a_1719_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1016 QN.t4 a_3599_411.t7 VDD.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VDD.t29 CLK.t1 a_343_411.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 GND a_1905_1050.t8 a_2702_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1019 VDD.t4 a_1905_1050.t7 a_1265_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 QN.t1 a_343_411.t10 VDD.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VDD.t23 QN.t6 a_3599_411.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VDD.t26 a_1265_989.t10 a_3599_411.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 QN a_3599_411.t8 a_3368_101.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1024 a_217_1050.t3 D.t2 VDD.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 VDD.t9 a_1265_989.t11 a_343_411.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1905_1050.t2 a_1265_989.t12 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 GND QN.t7 a_4013_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1028 VDD.t16 SN.t3 a_3599_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1905_1050.t5 SN.t5 VDD.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_217_1050.t1 a_343_411.t12 VDD.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_343_411.t0 a_217_1050.t9 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 VDD.t7 a_217_1050.t10 a_1905_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_343_411.t5 CLK.t3 VDD.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1265_989.t1 a_1905_1050.t9 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 VDD.t17 a_3599_411.t9 QN.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 VDD.t20 CLK.t4 a_1265_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VDD D 0.08fF
C1 VDD CLK 0.31fF
C2 VDD SN 0.10fF
C3 SN CLK 0.09fF
C4 VDD QN 1.44fF
C5 SN QN 0.42fF
R0 QN.n0 QN.t6 512.525
R1 QN.n0 QN.t5 371.139
R2 QN.n1 QN.t7 261.115
R3 QN.n6 QN.n5 205.778
R4 QN.n1 QN.n0 189.266
R5 QN.n6 QN.n4 179.052
R6 QN QN.n6 77.269
R7 QN.n4 QN.n3 76.002
R8 QN.n7 QN.n1 76
R9 QN.n2 QN.t2 14.282
R10 QN.n2 QN.t4 14.282
R11 QN.n3 QN.t3 14.282
R12 QN.n3 QN.t1 14.282
R13 QN.n4 QN.n2 12.85
R14 QN.n7 QN 0.046
R15 VDD.n314 VDD.n312 144.705
R16 VDD.n225 VDD.n223 144.705
R17 VDD.n395 VDD.n393 144.705
R18 VDD.n164 VDD.n162 144.705
R19 VDD.n103 VDD.n101 144.705
R20 VDD.n43 VDD.n42 76
R21 VDD.n48 VDD.n47 76
R22 VDD.n53 VDD.n52 76
R23 VDD.n60 VDD.n59 76
R24 VDD.n65 VDD.n64 76
R25 VDD.n70 VDD.n69 76
R26 VDD.n74 VDD.n73 76
R27 VDD.n78 VDD.n77 76
R28 VDD.n105 VDD.n104 76
R29 VDD.n110 VDD.n109 76
R30 VDD.n115 VDD.n114 76
R31 VDD.n121 VDD.n120 76
R32 VDD.n126 VDD.n125 76
R33 VDD.n131 VDD.n130 76
R34 VDD.n136 VDD.n135 76
R35 VDD.n140 VDD.n139 76
R36 VDD.n166 VDD.n165 76
R37 VDD.n171 VDD.n170 76
R38 VDD.n176 VDD.n175 76
R39 VDD.n182 VDD.n181 76
R40 VDD.n187 VDD.n186 76
R41 VDD.n192 VDD.n191 76
R42 VDD.n197 VDD.n196 76
R43 VDD.n201 VDD.n200 76
R44 VDD.n227 VDD.n226 76
R45 VDD.n231 VDD.n230 76
R46 VDD.n444 VDD.n443 76
R47 VDD.n440 VDD.n439 76
R48 VDD.n435 VDD.n434 76
R49 VDD.n428 VDD.n427 76
R50 VDD.n423 VDD.n422 76
R51 VDD.n418 VDD.n417 76
R52 VDD.n411 VDD.n410 76
R53 VDD.n406 VDD.n405 76
R54 VDD.n401 VDD.n400 76
R55 VDD.n397 VDD.n396 76
R56 VDD.n371 VDD.n370 76
R57 VDD.n367 VDD.n366 76
R58 VDD.n363 VDD.n362 76
R59 VDD.n359 VDD.n358 76
R60 VDD.n354 VDD.n353 76
R61 VDD.n347 VDD.n346 76
R62 VDD.n342 VDD.n341 76
R63 VDD.n337 VDD.n336 76
R64 VDD.n330 VDD.n329 76
R65 VDD.n325 VDD.n324 76
R66 VDD.n320 VDD.n319 76
R67 VDD.n316 VDD.n315 76
R68 VDD.n289 VDD.n288 76
R69 VDD.n285 VDD.n284 76
R70 VDD.n280 VDD.n279 76
R71 VDD.n275 VDD.n274 76
R72 VDD.n269 VDD.n268 76
R73 VDD.n264 VDD.n263 76
R74 VDD.n259 VDD.n258 76
R75 VDD.n254 VDD.n253 76
R76 VDD.n27 VDD.n26 64.064
R77 VDD.n437 VDD.n436 64.064
R78 VDD.n356 VDD.n355 64.064
R79 VDD.n62 VDD.n61 59.488
R80 VDD.n408 VDD.n407 59.488
R81 VDD.n327 VDD.n326 59.488
R82 VDD.n255 VDD.t12 55.106
R83 VDD.n321 VDD.t1 55.106
R84 VDD.n402 VDD.t10 55.106
R85 VDD.n193 VDD.t8 55.106
R86 VDD.n132 VDD.t14 55.106
R87 VDD.n66 VDD.t24 55.106
R88 VDD.n362 VDD.t9 55.106
R89 VDD.n443 VDD.t0 55.106
R90 VDD.n30 VDD.t26 55.106
R91 VDD.n281 VDD.t13 55.106
R92 VDD.n167 VDD.t20 55.106
R93 VDD.n106 VDD.t17 55.106
R94 VDD.n271 VDD.n270 40.824
R95 VDD.n332 VDD.n331 40.824
R96 VDD.n352 VDD.n351 40.824
R97 VDD.n413 VDD.n412 40.824
R98 VDD.n433 VDD.n432 40.824
R99 VDD.n178 VDD.n177 40.824
R100 VDD.n117 VDD.n116 40.824
R101 VDD.n55 VDD.n54 40.824
R102 VDD.n41 VDD.n40 40.824
R103 VDD.n376 VDD.n375 36.774
R104 VDD.n206 VDD.n205 36.774
R105 VDD.n145 VDD.n144 36.774
R106 VDD.n83 VDD.n82 36.774
R107 VDD.n305 VDD.n304 36.774
R108 VDD.n112 VDD.n111 36.608
R109 VDD.n173 VDD.n172 36.608
R110 VDD.n277 VDD.n276 36.608
R111 VDD.n35 VDD.n34 34.942
R112 VDD.n128 VDD.n127 32.032
R113 VDD.n189 VDD.n188 32.032
R114 VDD.n261 VDD.n260 32.032
R115 VDD.n38 VDD.n37 27.456
R116 VDD.n430 VDD.n429 27.456
R117 VDD.n349 VDD.n348 27.456
R118 VDD.n57 VDD.n56 22.88
R119 VDD.n415 VDD.n414 22.88
R120 VDD.n334 VDD.n333 22.88
R121 VDD.n253 VDD.n250 21.841
R122 VDD.n23 VDD.n20 21.841
R123 VDD.n270 VDD.t15 14.282
R124 VDD.n270 VDD.t11 14.282
R125 VDD.n331 VDD.t27 14.282
R126 VDD.n331 VDD.t2 14.282
R127 VDD.n351 VDD.t6 14.282
R128 VDD.n351 VDD.t29 14.282
R129 VDD.n412 VDD.t28 14.282
R130 VDD.n412 VDD.t7 14.282
R131 VDD.n432 VDD.t18 14.282
R132 VDD.n432 VDD.t3 14.282
R133 VDD.n177 VDD.t22 14.282
R134 VDD.n177 VDD.t4 14.282
R135 VDD.n116 VDD.t25 14.282
R136 VDD.n116 VDD.t19 14.282
R137 VDD.n54 VDD.t21 14.282
R138 VDD.n54 VDD.t23 14.282
R139 VDD.n40 VDD.t5 14.282
R140 VDD.n40 VDD.t16 14.282
R141 VDD.n250 VDD.n233 14.167
R142 VDD.n233 VDD.n232 14.167
R143 VDD.n391 VDD.n373 14.167
R144 VDD.n373 VDD.n372 14.167
R145 VDD.n221 VDD.n203 14.167
R146 VDD.n203 VDD.n202 14.167
R147 VDD.n160 VDD.n142 14.167
R148 VDD.n142 VDD.n141 14.167
R149 VDD.n99 VDD.n80 14.167
R150 VDD.n80 VDD.n79 14.167
R151 VDD.n310 VDD.n291 14.167
R152 VDD.n291 VDD.n290 14.167
R153 VDD.n20 VDD.n19 14.167
R154 VDD.n19 VDD.n17 14.167
R155 VDD.n33 VDD.n30 14.167
R156 VDD.n30 VDD.n29 14.167
R157 VDD.n104 VDD.n100 14.167
R158 VDD.n165 VDD.n161 14.167
R159 VDD.n226 VDD.n222 14.167
R160 VDD.n396 VDD.n392 14.167
R161 VDD.n315 VDD.n311 14.167
R162 VDD.n50 VDD.n49 13.728
R163 VDD.n420 VDD.n419 13.728
R164 VDD.n339 VDD.n338 13.728
R165 VDD.n23 VDD.n22 13.653
R166 VDD.n22 VDD.n21 13.653
R167 VDD.n33 VDD.n32 13.653
R168 VDD.n32 VDD.n31 13.653
R169 VDD.n30 VDD.n25 13.653
R170 VDD.n25 VDD.n24 13.653
R171 VDD.n29 VDD.n28 13.653
R172 VDD.n28 VDD.n27 13.653
R173 VDD.n42 VDD.n39 13.653
R174 VDD.n39 VDD.n38 13.653
R175 VDD.n47 VDD.n46 13.653
R176 VDD.n46 VDD.n45 13.653
R177 VDD.n52 VDD.n51 13.653
R178 VDD.n51 VDD.n50 13.653
R179 VDD.n59 VDD.n58 13.653
R180 VDD.n58 VDD.n57 13.653
R181 VDD.n64 VDD.n63 13.653
R182 VDD.n63 VDD.n62 13.653
R183 VDD.n69 VDD.n68 13.653
R184 VDD.n68 VDD.n67 13.653
R185 VDD.n73 VDD.n72 13.653
R186 VDD.n72 VDD.n71 13.653
R187 VDD.n77 VDD.n76 13.653
R188 VDD.n76 VDD.n75 13.653
R189 VDD.n104 VDD.n103 13.653
R190 VDD.n103 VDD.n102 13.653
R191 VDD.n109 VDD.n108 13.653
R192 VDD.n108 VDD.n107 13.653
R193 VDD.n114 VDD.n113 13.653
R194 VDD.n113 VDD.n112 13.653
R195 VDD.n120 VDD.n119 13.653
R196 VDD.n119 VDD.n118 13.653
R197 VDD.n125 VDD.n124 13.653
R198 VDD.n124 VDD.n123 13.653
R199 VDD.n130 VDD.n129 13.653
R200 VDD.n129 VDD.n128 13.653
R201 VDD.n135 VDD.n134 13.653
R202 VDD.n134 VDD.n133 13.653
R203 VDD.n139 VDD.n138 13.653
R204 VDD.n138 VDD.n137 13.653
R205 VDD.n165 VDD.n164 13.653
R206 VDD.n164 VDD.n163 13.653
R207 VDD.n170 VDD.n169 13.653
R208 VDD.n169 VDD.n168 13.653
R209 VDD.n175 VDD.n174 13.653
R210 VDD.n174 VDD.n173 13.653
R211 VDD.n181 VDD.n180 13.653
R212 VDD.n180 VDD.n179 13.653
R213 VDD.n186 VDD.n185 13.653
R214 VDD.n185 VDD.n184 13.653
R215 VDD.n191 VDD.n190 13.653
R216 VDD.n190 VDD.n189 13.653
R217 VDD.n196 VDD.n195 13.653
R218 VDD.n195 VDD.n194 13.653
R219 VDD.n200 VDD.n199 13.653
R220 VDD.n199 VDD.n198 13.653
R221 VDD.n226 VDD.n225 13.653
R222 VDD.n225 VDD.n224 13.653
R223 VDD.n230 VDD.n229 13.653
R224 VDD.n229 VDD.n228 13.653
R225 VDD.n443 VDD.n442 13.653
R226 VDD.n442 VDD.n441 13.653
R227 VDD.n439 VDD.n438 13.653
R228 VDD.n438 VDD.n437 13.653
R229 VDD.n434 VDD.n431 13.653
R230 VDD.n431 VDD.n430 13.653
R231 VDD.n427 VDD.n426 13.653
R232 VDD.n426 VDD.n425 13.653
R233 VDD.n422 VDD.n421 13.653
R234 VDD.n421 VDD.n420 13.653
R235 VDD.n417 VDD.n416 13.653
R236 VDD.n416 VDD.n415 13.653
R237 VDD.n410 VDD.n409 13.653
R238 VDD.n409 VDD.n408 13.653
R239 VDD.n405 VDD.n404 13.653
R240 VDD.n404 VDD.n403 13.653
R241 VDD.n400 VDD.n399 13.653
R242 VDD.n399 VDD.n398 13.653
R243 VDD.n396 VDD.n395 13.653
R244 VDD.n395 VDD.n394 13.653
R245 VDD.n370 VDD.n369 13.653
R246 VDD.n369 VDD.n368 13.653
R247 VDD.n366 VDD.n365 13.653
R248 VDD.n365 VDD.n364 13.653
R249 VDD.n362 VDD.n361 13.653
R250 VDD.n361 VDD.n360 13.653
R251 VDD.n358 VDD.n357 13.653
R252 VDD.n357 VDD.n356 13.653
R253 VDD.n353 VDD.n350 13.653
R254 VDD.n350 VDD.n349 13.653
R255 VDD.n346 VDD.n345 13.653
R256 VDD.n345 VDD.n344 13.653
R257 VDD.n341 VDD.n340 13.653
R258 VDD.n340 VDD.n339 13.653
R259 VDD.n336 VDD.n335 13.653
R260 VDD.n335 VDD.n334 13.653
R261 VDD.n329 VDD.n328 13.653
R262 VDD.n328 VDD.n327 13.653
R263 VDD.n324 VDD.n323 13.653
R264 VDD.n323 VDD.n322 13.653
R265 VDD.n319 VDD.n318 13.653
R266 VDD.n318 VDD.n317 13.653
R267 VDD.n315 VDD.n314 13.653
R268 VDD.n314 VDD.n313 13.653
R269 VDD.n288 VDD.n287 13.653
R270 VDD.n287 VDD.n286 13.653
R271 VDD.n284 VDD.n283 13.653
R272 VDD.n283 VDD.n282 13.653
R273 VDD.n279 VDD.n278 13.653
R274 VDD.n278 VDD.n277 13.653
R275 VDD.n274 VDD.n273 13.653
R276 VDD.n273 VDD.n272 13.653
R277 VDD.n268 VDD.n267 13.653
R278 VDD.n267 VDD.n266 13.653
R279 VDD.n263 VDD.n262 13.653
R280 VDD.n262 VDD.n261 13.653
R281 VDD.n258 VDD.n257 13.653
R282 VDD.n257 VDD.n256 13.653
R283 VDD.n253 VDD.n252 13.653
R284 VDD.n252 VDD.n251 13.653
R285 VDD.n4 VDD.n2 12.915
R286 VDD.n4 VDD.n3 12.66
R287 VDD.n13 VDD.n12 12.343
R288 VDD.n10 VDD.n9 12.343
R289 VDD.n7 VDD.n6 12.343
R290 VDD.n45 VDD.n44 9.152
R291 VDD.n425 VDD.n424 9.152
R292 VDD.n344 VDD.n343 9.152
R293 VDD.n120 VDD.n117 8.658
R294 VDD.n181 VDD.n178 8.658
R295 VDD.n274 VDD.n271 8.658
R296 VDD.n392 VDD.n391 7.674
R297 VDD.n222 VDD.n221 7.674
R298 VDD.n161 VDD.n160 7.674
R299 VDD.n100 VDD.n99 7.674
R300 VDD.n311 VDD.n310 7.674
R301 VDD.n94 VDD.n93 7.5
R302 VDD.n88 VDD.n87 7.5
R303 VDD.n90 VDD.n89 7.5
R304 VDD.n85 VDD.n84 7.5
R305 VDD.n99 VDD.n98 7.5
R306 VDD.n155 VDD.n154 7.5
R307 VDD.n149 VDD.n148 7.5
R308 VDD.n151 VDD.n150 7.5
R309 VDD.n157 VDD.n147 7.5
R310 VDD.n157 VDD.n145 7.5
R311 VDD.n160 VDD.n159 7.5
R312 VDD.n216 VDD.n215 7.5
R313 VDD.n210 VDD.n209 7.5
R314 VDD.n212 VDD.n211 7.5
R315 VDD.n218 VDD.n208 7.5
R316 VDD.n218 VDD.n206 7.5
R317 VDD.n221 VDD.n220 7.5
R318 VDD.n386 VDD.n385 7.5
R319 VDD.n380 VDD.n379 7.5
R320 VDD.n382 VDD.n381 7.5
R321 VDD.n388 VDD.n378 7.5
R322 VDD.n388 VDD.n376 7.5
R323 VDD.n391 VDD.n390 7.5
R324 VDD.n295 VDD.n294 7.5
R325 VDD.n298 VDD.n297 7.5
R326 VDD.n300 VDD.n299 7.5
R327 VDD.n303 VDD.n302 7.5
R328 VDD.n310 VDD.n309 7.5
R329 VDD.n245 VDD.n244 7.5
R330 VDD.n239 VDD.n238 7.5
R331 VDD.n241 VDD.n240 7.5
R332 VDD.n247 VDD.n237 7.5
R333 VDD.n247 VDD.n235 7.5
R334 VDD.n250 VDD.n249 7.5
R335 VDD.n20 VDD.n16 7.5
R336 VDD.n2 VDD.n1 7.5
R337 VDD.n6 VDD.n5 7.5
R338 VDD.n9 VDD.n8 7.5
R339 VDD.n19 VDD.n18 7.5
R340 VDD.n14 VDD.n0 7.5
R341 VDD.n86 VDD.n83 6.772
R342 VDD.n97 VDD.n81 6.772
R343 VDD.n95 VDD.n92 6.772
R344 VDD.n91 VDD.n88 6.772
R345 VDD.n158 VDD.n143 6.772
R346 VDD.n156 VDD.n153 6.772
R347 VDD.n152 VDD.n149 6.772
R348 VDD.n219 VDD.n204 6.772
R349 VDD.n217 VDD.n214 6.772
R350 VDD.n213 VDD.n210 6.772
R351 VDD.n389 VDD.n374 6.772
R352 VDD.n387 VDD.n384 6.772
R353 VDD.n383 VDD.n380 6.772
R354 VDD.n248 VDD.n234 6.772
R355 VDD.n246 VDD.n243 6.772
R356 VDD.n242 VDD.n239 6.772
R357 VDD.n86 VDD.n85 6.772
R358 VDD.n91 VDD.n90 6.772
R359 VDD.n95 VDD.n94 6.772
R360 VDD.n98 VDD.n97 6.772
R361 VDD.n152 VDD.n151 6.772
R362 VDD.n156 VDD.n155 6.772
R363 VDD.n159 VDD.n158 6.772
R364 VDD.n213 VDD.n212 6.772
R365 VDD.n217 VDD.n216 6.772
R366 VDD.n220 VDD.n219 6.772
R367 VDD.n383 VDD.n382 6.772
R368 VDD.n387 VDD.n386 6.772
R369 VDD.n390 VDD.n389 6.772
R370 VDD.n242 VDD.n241 6.772
R371 VDD.n246 VDD.n245 6.772
R372 VDD.n249 VDD.n248 6.772
R373 VDD.n309 VDD.n308 6.772
R374 VDD.n296 VDD.n293 6.772
R375 VDD.n301 VDD.n298 6.772
R376 VDD.n306 VDD.n303 6.772
R377 VDD.n306 VDD.n305 6.772
R378 VDD.n301 VDD.n300 6.772
R379 VDD.n296 VDD.n295 6.772
R380 VDD.n308 VDD.n292 6.772
R381 VDD.n59 VDD.n55 6.69
R382 VDD.n417 VDD.n413 6.69
R383 VDD.n336 VDD.n332 6.69
R384 VDD.n34 VDD.n23 6.487
R385 VDD.n34 VDD.n33 6.475
R386 VDD.n16 VDD.n15 6.458
R387 VDD.n42 VDD.n41 6.296
R388 VDD.n434 VDD.n433 6.296
R389 VDD.n353 VDD.n352 6.296
R390 VDD.n147 VDD.n146 6.202
R391 VDD.n208 VDD.n207 6.202
R392 VDD.n378 VDD.n377 6.202
R393 VDD.n237 VDD.n236 6.202
R394 VDD.n123 VDD.n122 4.576
R395 VDD.n184 VDD.n183 4.576
R396 VDD.n266 VDD.n265 4.576
R397 VDD.n135 VDD.n132 2.754
R398 VDD.n196 VDD.n193 2.754
R399 VDD.n258 VDD.n255 2.754
R400 VDD.n109 VDD.n106 2.361
R401 VDD.n170 VDD.n167 2.361
R402 VDD.n284 VDD.n281 2.361
R403 VDD.n14 VDD.n7 1.329
R404 VDD.n14 VDD.n10 1.329
R405 VDD.n14 VDD.n11 1.329
R406 VDD.n14 VDD.n13 1.329
R407 VDD.n15 VDD.n14 0.696
R408 VDD.n14 VDD.n4 0.696
R409 VDD.n69 VDD.n66 0.393
R410 VDD.n405 VDD.n402 0.393
R411 VDD.n324 VDD.n321 0.393
R412 VDD.n96 VDD.n95 0.365
R413 VDD.n96 VDD.n91 0.365
R414 VDD.n96 VDD.n86 0.365
R415 VDD.n97 VDD.n96 0.365
R416 VDD.n157 VDD.n156 0.365
R417 VDD.n157 VDD.n152 0.365
R418 VDD.n158 VDD.n157 0.365
R419 VDD.n218 VDD.n217 0.365
R420 VDD.n218 VDD.n213 0.365
R421 VDD.n219 VDD.n218 0.365
R422 VDD.n388 VDD.n387 0.365
R423 VDD.n388 VDD.n383 0.365
R424 VDD.n389 VDD.n388 0.365
R425 VDD.n247 VDD.n246 0.365
R426 VDD.n247 VDD.n242 0.365
R427 VDD.n248 VDD.n247 0.365
R428 VDD.n307 VDD.n306 0.365
R429 VDD.n307 VDD.n301 0.365
R430 VDD.n307 VDD.n296 0.365
R431 VDD.n308 VDD.n307 0.365
R432 VDD.n105 VDD.n78 0.29
R433 VDD.n166 VDD.n140 0.29
R434 VDD.n227 VDD.n201 0.29
R435 VDD.n397 VDD.n371 0.29
R436 VDD.n316 VDD.n289 0.29
R437 VDD.n254 VDD 0.207
R438 VDD.n53 VDD.n48 0.197
R439 VDD.n428 VDD.n423 0.197
R440 VDD.n347 VDD.n342 0.197
R441 VDD.n126 VDD.n121 0.181
R442 VDD.n187 VDD.n182 0.181
R443 VDD.n275 VDD.n269 0.181
R444 VDD.n36 VDD.n35 0.145
R445 VDD.n43 VDD.n36 0.145
R446 VDD.n48 VDD.n43 0.145
R447 VDD.n60 VDD.n53 0.145
R448 VDD.n65 VDD.n60 0.145
R449 VDD.n70 VDD.n65 0.145
R450 VDD.n74 VDD.n70 0.145
R451 VDD.n78 VDD.n74 0.145
R452 VDD.n110 VDD.n105 0.145
R453 VDD.n115 VDD.n110 0.145
R454 VDD.n121 VDD.n115 0.145
R455 VDD.n131 VDD.n126 0.145
R456 VDD.n136 VDD.n131 0.145
R457 VDD.n140 VDD.n136 0.145
R458 VDD.n171 VDD.n166 0.145
R459 VDD.n176 VDD.n171 0.145
R460 VDD.n182 VDD.n176 0.145
R461 VDD.n192 VDD.n187 0.145
R462 VDD.n197 VDD.n192 0.145
R463 VDD.n201 VDD.n197 0.145
R464 VDD.n231 VDD.n227 0.145
R465 VDD.n444 VDD.n440 0.145
R466 VDD.n440 VDD.n435 0.145
R467 VDD.n435 VDD.n428 0.145
R468 VDD.n423 VDD.n418 0.145
R469 VDD.n418 VDD.n411 0.145
R470 VDD.n411 VDD.n406 0.145
R471 VDD.n406 VDD.n401 0.145
R472 VDD.n401 VDD.n397 0.145
R473 VDD.n371 VDD.n367 0.145
R474 VDD.n367 VDD.n363 0.145
R475 VDD.n363 VDD.n359 0.145
R476 VDD.n359 VDD.n354 0.145
R477 VDD.n354 VDD.n347 0.145
R478 VDD.n342 VDD.n337 0.145
R479 VDD.n337 VDD.n330 0.145
R480 VDD.n330 VDD.n325 0.145
R481 VDD.n325 VDD.n320 0.145
R482 VDD.n320 VDD.n316 0.145
R483 VDD.n289 VDD.n285 0.145
R484 VDD.n285 VDD.n280 0.145
R485 VDD.n280 VDD.n275 0.145
R486 VDD.n269 VDD.n264 0.145
R487 VDD.n264 VDD.n259 0.145
R488 VDD.n259 VDD.n254 0.145
R489 VDD VDD.n444 0.137
R490 VDD VDD.n231 0.008
R491 a_3599_411.n2 a_3599_411.t9 472.359
R492 a_3599_411.n2 a_3599_411.t7 384.527
R493 a_3599_411.n3 a_3599_411.t8 241.172
R494 a_3599_411.n8 a_3599_411.n7 213.104
R495 a_3599_411.n9 a_3599_411.n8 170.799
R496 a_3599_411.n8 a_3599_411.n3 156.035
R497 a_3599_411.n3 a_3599_411.n2 110.06
R498 a_3599_411.n11 a_3599_411.n10 79.231
R499 a_3599_411.n10 a_3599_411.n9 63.152
R500 a_3599_411.n7 a_3599_411.n6 30
R501 a_3599_411.n5 a_3599_411.n4 24.383
R502 a_3599_411.n7 a_3599_411.n5 23.684
R503 a_3599_411.n9 a_3599_411.n1 16.08
R504 a_3599_411.n10 a_3599_411.n0 16.08
R505 a_3599_411.n1 a_3599_411.t5 14.282
R506 a_3599_411.n1 a_3599_411.t0 14.282
R507 a_3599_411.n0 a_3599_411.t1 14.282
R508 a_3599_411.n0 a_3599_411.t2 14.282
R509 a_3599_411.n11 a_3599_411.t3 14.282
R510 a_3599_411.t4 a_3599_411.n11 14.282
R511 SN.n2 SN.t1 479.223
R512 SN.n0 SN.t3 479.223
R513 SN.n2 SN.t5 375.52
R514 SN.n0 SN.t2 375.52
R515 SN.n3 SN.n2 175.429
R516 SN.n1 SN.n0 175.429
R517 SN.n3 SN.t4 162.048
R518 SN.n1 SN.t0 162.048
R519 SN.n4 SN.n1 84.388
R520 SN.n4 SN.n3 76
R521 SN.n4 SN 0.046
R522 a_4013_103.t0 a_4013_103.n0 117.777
R523 a_4013_103.n2 a_4013_103.n1 55.228
R524 a_4013_103.n4 a_4013_103.n3 9.111
R525 a_4013_103.n8 a_4013_103.n6 7.859
R526 a_4013_103.t0 a_4013_103.n2 4.04
R527 a_4013_103.t0 a_4013_103.n8 3.034
R528 a_4013_103.n6 a_4013_103.n4 1.964
R529 a_4013_103.n6 a_4013_103.n5 1.964
R530 a_4013_103.n8 a_4013_103.n7 0.443
R531 a_4294_210.n10 a_4294_210.n8 82.852
R532 a_4294_210.n11 a_4294_210.n0 49.6
R533 a_4294_210.n7 a_4294_210.n6 32.833
R534 a_4294_210.n8 a_4294_210.t1 32.416
R535 a_4294_210.n10 a_4294_210.n9 27.2
R536 a_4294_210.n3 a_4294_210.n2 23.284
R537 a_4294_210.n11 a_4294_210.n10 22.4
R538 a_4294_210.n7 a_4294_210.n4 19.017
R539 a_4294_210.n6 a_4294_210.n5 13.494
R540 a_4294_210.t1 a_4294_210.n1 7.04
R541 a_4294_210.t1 a_4294_210.n3 5.727
R542 a_4294_210.n8 a_4294_210.n7 1.435
R543 a_1265_989.n6 a_1265_989.t12 454.685
R544 a_1265_989.n8 a_1265_989.t5 454.685
R545 a_1265_989.n4 a_1265_989.t8 454.685
R546 a_1265_989.n6 a_1265_989.t7 428.979
R547 a_1265_989.n8 a_1265_989.t11 428.979
R548 a_1265_989.n4 a_1265_989.t10 428.979
R549 a_1265_989.n7 a_1265_989.t6 264.512
R550 a_1265_989.n9 a_1265_989.t9 264.512
R551 a_1265_989.n5 a_1265_989.t13 264.512
R552 a_1265_989.n14 a_1265_989.n12 237.145
R553 a_1265_989.n12 a_1265_989.n3 125.947
R554 a_1265_989.n11 a_1265_989.n5 81.396
R555 a_1265_989.n10 a_1265_989.n9 79.491
R556 a_1265_989.n3 a_1265_989.n2 76.002
R557 a_1265_989.n10 a_1265_989.n7 76
R558 a_1265_989.n12 a_1265_989.n11 76
R559 a_1265_989.n7 a_1265_989.n6 71.894
R560 a_1265_989.n9 a_1265_989.n8 71.894
R561 a_1265_989.n5 a_1265_989.n4 71.894
R562 a_1265_989.n15 a_1265_989.n0 55.263
R563 a_1265_989.n14 a_1265_989.n13 30
R564 a_1265_989.n15 a_1265_989.n14 23.684
R565 a_1265_989.n1 a_1265_989.t2 14.282
R566 a_1265_989.n1 a_1265_989.t4 14.282
R567 a_1265_989.n2 a_1265_989.t0 14.282
R568 a_1265_989.n2 a_1265_989.t1 14.282
R569 a_1265_989.n3 a_1265_989.n1 12.85
R570 a_1265_989.n11 a_1265_989.n10 2.947
R571 a_343_411.n0 a_343_411.t7 480.392
R572 a_343_411.n2 a_343_411.t9 472.359
R573 a_343_411.n0 a_343_411.t10 403.272
R574 a_343_411.n2 a_343_411.t12 384.527
R575 a_343_411.n1 a_343_411.t8 336.586
R576 a_343_411.n3 a_343_411.t11 294.278
R577 a_343_411.n9 a_343_411.n8 265.87
R578 a_343_411.n13 a_343_411.n9 117.354
R579 a_343_411.n4 a_343_411.n1 83.304
R580 a_343_411.n4 a_343_411.n3 80.032
R581 a_343_411.n12 a_343_411.n11 79.232
R582 a_343_411.n9 a_343_411.n4 76
R583 a_343_411.n13 a_343_411.n12 63.152
R584 a_343_411.n3 a_343_411.n2 56.954
R585 a_343_411.n1 a_343_411.n0 45.341
R586 a_343_411.n8 a_343_411.n7 30
R587 a_343_411.n6 a_343_411.n5 24.383
R588 a_343_411.n8 a_343_411.n6 23.684
R589 a_343_411.n12 a_343_411.n10 16.08
R590 a_343_411.n14 a_343_411.n13 16.078
R591 a_343_411.n10 a_343_411.t6 14.282
R592 a_343_411.n10 a_343_411.t5 14.282
R593 a_343_411.n11 a_343_411.t1 14.282
R594 a_343_411.n11 a_343_411.t0 14.282
R595 a_343_411.n14 a_343_411.t3 14.282
R596 a_343_411.t4 a_343_411.n14 14.282
R597 a_1905_1050.n0 a_1905_1050.t7 480.392
R598 a_1905_1050.n0 a_1905_1050.t9 403.272
R599 a_1905_1050.n1 a_1905_1050.t8 230.374
R600 a_1905_1050.n10 a_1905_1050.n6 223.905
R601 a_1905_1050.n6 a_1905_1050.n5 159.998
R602 a_1905_1050.n6 a_1905_1050.n1 153.315
R603 a_1905_1050.n1 a_1905_1050.n0 151.553
R604 a_1905_1050.n9 a_1905_1050.n8 79.232
R605 a_1905_1050.n10 a_1905_1050.n9 63.152
R606 a_1905_1050.n5 a_1905_1050.n4 30
R607 a_1905_1050.n3 a_1905_1050.n2 24.383
R608 a_1905_1050.n5 a_1905_1050.n3 23.684
R609 a_1905_1050.n9 a_1905_1050.n7 16.08
R610 a_1905_1050.n11 a_1905_1050.n10 16.078
R611 a_1905_1050.n7 a_1905_1050.t6 14.282
R612 a_1905_1050.n7 a_1905_1050.t5 14.282
R613 a_1905_1050.n8 a_1905_1050.t0 14.282
R614 a_1905_1050.n8 a_1905_1050.t4 14.282
R615 a_1905_1050.t3 a_1905_1050.n11 14.282
R616 a_1905_1050.n11 a_1905_1050.t2 14.282
R617 CLK.n0 CLK.t4 472.359
R618 CLK.n2 CLK.t1 459.505
R619 CLK.n2 CLK.t3 384.527
R620 CLK.n0 CLK.t0 384.527
R621 CLK.n3 CLK.t2 322.152
R622 CLK.n1 CLK.t5 321.724
R623 CLK.n4 CLK.n3 49.342
R624 CLK.n4 CLK.n1 43.573
R625 CLK.n3 CLK.n2 27.599
R626 CLK.n1 CLK.n0 23.329
R627 CLK.n4 CLK 0.046
R628 a_2000_210.n9 a_2000_210.n7 82.852
R629 a_2000_210.n3 a_2000_210.n1 44.628
R630 a_2000_210.t0 a_2000_210.n9 32.417
R631 a_2000_210.n7 a_2000_210.n6 27.2
R632 a_2000_210.n5 a_2000_210.n4 23.498
R633 a_2000_210.n3 a_2000_210.n2 23.284
R634 a_2000_210.n7 a_2000_210.n5 22.4
R635 a_2000_210.t0 a_2000_210.n11 20.241
R636 a_2000_210.n11 a_2000_210.n10 13.494
R637 a_2000_210.t0 a_2000_210.n0 8.137
R638 a_2000_210.t0 a_2000_210.n3 5.727
R639 a_2000_210.n9 a_2000_210.n8 1.435
R640 D.n0 D.t0 480.392
R641 D.n0 D.t2 403.272
R642 D.n1 D.t1 310.033
R643 D.n2 D.n1 76
R644 D.n1 D.n0 71.894
R645 D.n2 D 0.046
R646 a_217_1050.n2 a_217_1050.t7 512.525
R647 a_217_1050.n0 a_217_1050.t10 512.525
R648 a_217_1050.n2 a_217_1050.t9 371.139
R649 a_217_1050.n0 a_217_1050.t5 371.139
R650 a_217_1050.n1 a_217_1050.t8 234.562
R651 a_217_1050.n3 a_217_1050.t6 234.204
R652 a_217_1050.n3 a_217_1050.n2 216.178
R653 a_217_1050.n1 a_217_1050.n0 215.819
R654 a_217_1050.n11 a_217_1050.n9 205.605
R655 a_217_1050.n9 a_217_1050.n8 157.486
R656 a_217_1050.n4 a_217_1050.n1 79.488
R657 a_217_1050.n9 a_217_1050.n4 77.314
R658 a_217_1050.n11 a_217_1050.n10 76.002
R659 a_217_1050.n4 a_217_1050.n3 76
R660 a_217_1050.n8 a_217_1050.n7 30
R661 a_217_1050.n6 a_217_1050.n5 24.383
R662 a_217_1050.n8 a_217_1050.n6 23.684
R663 a_217_1050.n10 a_217_1050.t4 14.282
R664 a_217_1050.n10 a_217_1050.t3 14.282
R665 a_217_1050.t2 a_217_1050.n12 14.282
R666 a_217_1050.n12 a_217_1050.t1 14.282
R667 a_217_1050.n12 a_217_1050.n11 12.848
R668 a_1038_210.n10 a_1038_210.n8 82.852
R669 a_1038_210.n7 a_1038_210.n6 32.833
R670 a_1038_210.n8 a_1038_210.t1 32.416
R671 a_1038_210.n10 a_1038_210.n9 27.2
R672 a_1038_210.n11 a_1038_210.n0 23.498
R673 a_1038_210.n3 a_1038_210.n2 23.284
R674 a_1038_210.n11 a_1038_210.n10 22.4
R675 a_1038_210.n7 a_1038_210.n4 19.017
R676 a_1038_210.n6 a_1038_210.n5 13.494
R677 a_1038_210.t1 a_1038_210.n1 7.04
R678 a_1038_210.t1 a_1038_210.n3 5.727
R679 a_1038_210.n8 a_1038_210.n7 1.435
R680 a_757_103.t0 a_757_103.n0 117.777
R681 a_757_103.n2 a_757_103.n1 55.228
R682 a_757_103.n4 a_757_103.n3 9.111
R683 a_757_103.t0 a_757_103.n2 4.04
R684 a_757_103.n8 a_757_103.n7 2.455
R685 a_757_103.n6 a_757_103.n4 1.964
R686 a_757_103.n6 a_757_103.n5 1.964
R687 a_757_103.n8 a_757_103.n6 0.636
R688 a_757_103.t0 a_757_103.n8 0.246
R689 GND.n38 GND.n36 219.745
R690 GND.n144 GND.n143 219.745
R691 GND.n186 GND.n184 219.745
R692 GND.n104 GND.n102 219.745
R693 GND.n71 GND.n70 219.745
R694 GND.n27 GND.n26 85.559
R695 GND.n153 GND.n152 85.559
R696 GND.n38 GND.n37 85.529
R697 GND.n144 GND.n142 85.529
R698 GND.n186 GND.n185 85.529
R699 GND.n104 GND.n103 85.529
R700 GND.n71 GND.n69 85.529
R701 GND.n114 GND.n113 76
R702 GND.n12 GND.n11 76
R703 GND.n15 GND.n14 76
R704 GND.n18 GND.n17 76
R705 GND.n21 GND.n20 76
R706 GND.n24 GND.n23 76
R707 GND.n29 GND.n28 76
R708 GND.n32 GND.n31 76
R709 GND.n35 GND.n34 76
R710 GND.n42 GND.n41 76
R711 GND.n45 GND.n44 76
R712 GND.n48 GND.n47 76
R713 GND.n51 GND.n50 76
R714 GND.n54 GND.n53 76
R715 GND.n62 GND.n61 76
R716 GND.n65 GND.n64 76
R717 GND.n68 GND.n67 76
R718 GND.n75 GND.n74 76
R719 GND.n78 GND.n77 76
R720 GND.n81 GND.n80 76
R721 GND.n84 GND.n83 76
R722 GND.n87 GND.n86 76
R723 GND.n95 GND.n94 76
R724 GND.n98 GND.n97 76
R725 GND.n101 GND.n100 76
R726 GND.n108 GND.n107 76
R727 GND.n111 GND.n110 76
R728 GND.n221 GND.n220 76
R729 GND.n218 GND.n217 76
R730 GND.n215 GND.n214 76
R731 GND.n212 GND.n211 76
R732 GND.n209 GND.n208 76
R733 GND.n206 GND.n205 76
R734 GND.n203 GND.n202 76
R735 GND.n200 GND.n199 76
R736 GND.n192 GND.n191 76
R737 GND.n189 GND.n188 76
R738 GND.n182 GND.n181 76
R739 GND.n179 GND.n178 76
R740 GND.n176 GND.n175 76
R741 GND.n173 GND.n172 76
R742 GND.n170 GND.n169 76
R743 GND.n167 GND.n166 76
R744 GND.n164 GND.n163 76
R745 GND.n161 GND.n160 76
R746 GND.n158 GND.n157 76
R747 GND.n155 GND.n154 76
R748 GND.n150 GND.n149 76
R749 GND.n147 GND.n146 76
R750 GND.n140 GND.n139 76
R751 GND.n137 GND.n136 76
R752 GND.n134 GND.n133 76
R753 GND.n131 GND.n130 76
R754 GND.n128 GND.n127 76
R755 GND.n125 GND.n124 76
R756 GND.n117 GND.n116 76
R757 GND.n198 GND.n197 64.552
R758 GND.n59 GND.n58 63.835
R759 GND.n92 GND.n91 63.835
R760 GND.n122 GND.n121 63.835
R761 GND.n8 GND.n7 34.942
R762 GND.n58 GND.n57 28.421
R763 GND.n91 GND.n90 28.421
R764 GND.n197 GND.n196 28.421
R765 GND.n121 GND.n120 28.421
R766 GND.n58 GND.n56 25.263
R767 GND.n91 GND.n89 25.263
R768 GND.n197 GND.n195 25.263
R769 GND.n121 GND.n119 25.263
R770 GND.n56 GND.n55 24.383
R771 GND.n89 GND.n88 24.383
R772 GND.n195 GND.n194 24.383
R773 GND.n119 GND.n118 24.383
R774 GND.n6 GND.n5 14.167
R775 GND.n5 GND.n4 14.167
R776 GND.n41 GND.n39 14.167
R777 GND.n74 GND.n72 14.167
R778 GND.n107 GND.n105 14.167
R779 GND.n188 GND.n187 14.167
R780 GND.n146 GND.n145 14.167
R781 GND.n116 GND.n115 13.653
R782 GND.n124 GND.n123 13.653
R783 GND.n127 GND.n126 13.653
R784 GND.n130 GND.n129 13.653
R785 GND.n133 GND.n132 13.653
R786 GND.n136 GND.n135 13.653
R787 GND.n139 GND.n138 13.653
R788 GND.n146 GND.n141 13.653
R789 GND.n149 GND.n148 13.653
R790 GND.n154 GND.n151 13.653
R791 GND.n157 GND.n156 13.653
R792 GND.n160 GND.n159 13.653
R793 GND.n163 GND.n162 13.653
R794 GND.n166 GND.n165 13.653
R795 GND.n169 GND.n168 13.653
R796 GND.n172 GND.n171 13.653
R797 GND.n175 GND.n174 13.653
R798 GND.n178 GND.n177 13.653
R799 GND.n181 GND.n180 13.653
R800 GND.n188 GND.n183 13.653
R801 GND.n191 GND.n190 13.653
R802 GND.n199 GND.n193 13.653
R803 GND.n202 GND.n201 13.653
R804 GND.n205 GND.n204 13.653
R805 GND.n208 GND.n207 13.653
R806 GND.n211 GND.n210 13.653
R807 GND.n214 GND.n213 13.653
R808 GND.n217 GND.n216 13.653
R809 GND.n220 GND.n219 13.653
R810 GND.n110 GND.n109 13.653
R811 GND.n107 GND.n106 13.653
R812 GND.n100 GND.n99 13.653
R813 GND.n97 GND.n96 13.653
R814 GND.n94 GND.n93 13.653
R815 GND.n86 GND.n85 13.653
R816 GND.n83 GND.n82 13.653
R817 GND.n80 GND.n79 13.653
R818 GND.n77 GND.n76 13.653
R819 GND.n74 GND.n73 13.653
R820 GND.n67 GND.n66 13.653
R821 GND.n64 GND.n63 13.653
R822 GND.n61 GND.n60 13.653
R823 GND.n53 GND.n52 13.653
R824 GND.n50 GND.n49 13.653
R825 GND.n47 GND.n46 13.653
R826 GND.n44 GND.n43 13.653
R827 GND.n41 GND.n40 13.653
R828 GND.n34 GND.n33 13.653
R829 GND.n31 GND.n30 13.653
R830 GND.n28 GND.n25 13.653
R831 GND.n23 GND.n22 13.653
R832 GND.n20 GND.n19 13.653
R833 GND.n17 GND.n16 13.653
R834 GND.n14 GND.n13 13.653
R835 GND.n11 GND.n10 13.653
R836 GND.n4 GND.n3 13.653
R837 GND.n5 GND.n2 13.653
R838 GND.n6 GND.n1 13.653
R839 GND.n39 GND.n38 7.312
R840 GND.n145 GND.n144 7.312
R841 GND.n187 GND.n186 7.312
R842 GND.n105 GND.n104 7.312
R843 GND.n72 GND.n71 7.312
R844 GND.n7 GND.n0 7.083
R845 GND.n7 GND.n6 6.474
R846 GND.n61 GND.n59 3.935
R847 GND.n94 GND.n92 3.935
R848 GND.n124 GND.n122 3.935
R849 GND.n113 GND.n112 0.596
R850 GND.n42 GND.n35 0.29
R851 GND.n75 GND.n68 0.29
R852 GND.n108 GND.n101 0.29
R853 GND.n189 GND.n182 0.29
R854 GND.n147 GND.n140 0.29
R855 GND.n114 GND 0.207
R856 GND.n18 GND.n15 0.197
R857 GND.n212 GND.n209 0.197
R858 GND.n167 GND.n164 0.197
R859 GND.n28 GND.n27 0.196
R860 GND.n199 GND.n198 0.196
R861 GND.n154 GND.n153 0.196
R862 GND.n54 GND.n51 0.181
R863 GND.n87 GND.n84 0.181
R864 GND.n131 GND.n128 0.181
R865 GND.n9 GND.n8 0.145
R866 GND.n12 GND.n9 0.145
R867 GND.n15 GND.n12 0.145
R868 GND.n21 GND.n18 0.145
R869 GND.n24 GND.n21 0.145
R870 GND.n29 GND.n24 0.145
R871 GND.n32 GND.n29 0.145
R872 GND.n35 GND.n32 0.145
R873 GND.n45 GND.n42 0.145
R874 GND.n48 GND.n45 0.145
R875 GND.n51 GND.n48 0.145
R876 GND.n62 GND.n54 0.145
R877 GND.n65 GND.n62 0.145
R878 GND.n68 GND.n65 0.145
R879 GND.n78 GND.n75 0.145
R880 GND.n81 GND.n78 0.145
R881 GND.n84 GND.n81 0.145
R882 GND.n95 GND.n87 0.145
R883 GND.n98 GND.n95 0.145
R884 GND.n101 GND.n98 0.145
R885 GND.n111 GND.n108 0.145
R886 GND.n221 GND.n218 0.145
R887 GND.n218 GND.n215 0.145
R888 GND.n215 GND.n212 0.145
R889 GND.n209 GND.n206 0.145
R890 GND.n206 GND.n203 0.145
R891 GND.n203 GND.n200 0.145
R892 GND.n200 GND.n192 0.145
R893 GND.n192 GND.n189 0.145
R894 GND.n182 GND.n179 0.145
R895 GND.n179 GND.n176 0.145
R896 GND.n176 GND.n173 0.145
R897 GND.n173 GND.n170 0.145
R898 GND.n170 GND.n167 0.145
R899 GND.n164 GND.n161 0.145
R900 GND.n161 GND.n158 0.145
R901 GND.n158 GND.n155 0.145
R902 GND.n155 GND.n150 0.145
R903 GND.n150 GND.n147 0.145
R904 GND.n140 GND.n137 0.145
R905 GND.n137 GND.n134 0.145
R906 GND.n134 GND.n131 0.145
R907 GND.n128 GND.n125 0.145
R908 GND.n125 GND.n117 0.145
R909 GND.n117 GND.n114 0.145
R910 GND GND.n221 0.137
R911 GND GND.n111 0.008
R912 a_112_101.t0 a_112_101.n1 34.62
R913 a_112_101.t0 a_112_101.n0 8.137
R914 a_112_101.t0 a_112_101.n2 4.69
R915 a_3368_101.t0 a_3368_101.n1 34.62
R916 a_3368_101.t0 a_3368_101.n0 8.137
R917 a_3368_101.t0 a_3368_101.n2 4.69
R918 a_1719_103.n1 a_1719_103.n0 25.576
R919 a_1719_103.n3 a_1719_103.n2 9.111
R920 a_1719_103.n7 a_1719_103.n6 2.455
R921 a_1719_103.n5 a_1719_103.n3 1.964
R922 a_1719_103.n5 a_1719_103.n4 1.964
R923 a_1719_103.t0 a_1719_103.n1 1.871
R924 a_1719_103.n7 a_1719_103.n5 0.636
R925 a_1719_103.t0 a_1719_103.n7 0.246
R926 a_2702_101.t0 a_2702_101.n1 34.62
R927 a_2702_101.t0 a_2702_101.n0 8.137
R928 a_2702_101.t0 a_2702_101.n2 4.69
C6 SN GND 2.06fF
C7 VDD GND 18.31fF
C8 a_2702_101.n0 GND 0.05fF
C9 a_2702_101.n1 GND 0.12fF
C10 a_2702_101.n2 GND 0.04fF
C11 a_1719_103.n0 GND 0.09fF
C12 a_1719_103.n1 GND 0.10fF
C13 a_1719_103.n2 GND 0.05fF
C14 a_1719_103.n3 GND 0.03fF
C15 a_1719_103.n4 GND 0.04fF
C16 a_1719_103.n5 GND 0.03fF
C17 a_1719_103.n6 GND 0.04fF
C18 a_3368_101.n0 GND 0.05fF
C19 a_3368_101.n1 GND 0.12fF
C20 a_3368_101.n2 GND 0.04fF
C21 a_112_101.n0 GND 0.05fF
C22 a_112_101.n1 GND 0.12fF
C23 a_112_101.n2 GND 0.04fF
C24 a_757_103.n0 GND 0.03fF
C25 a_757_103.n1 GND 0.10fF
C26 a_757_103.n2 GND 0.10fF
C27 a_757_103.n3 GND 0.05fF
C28 a_757_103.n4 GND 0.03fF
C29 a_757_103.n5 GND 0.04fF
C30 a_757_103.n6 GND 0.03fF
C31 a_757_103.n7 GND 0.04fF
C32 a_1038_210.n0 GND 0.02fF
C33 a_1038_210.n1 GND 0.09fF
C34 a_1038_210.n2 GND 0.13fF
C35 a_1038_210.n3 GND 0.11fF
C36 a_1038_210.t1 GND 0.30fF
C37 a_1038_210.n4 GND 0.09fF
C38 a_1038_210.n5 GND 0.06fF
C39 a_1038_210.n6 GND 0.01fF
C40 a_1038_210.n7 GND 0.03fF
C41 a_1038_210.n8 GND 0.11fF
C42 a_1038_210.n9 GND 0.02fF
C43 a_1038_210.n10 GND 0.05fF
C44 a_1038_210.n11 GND 0.03fF
C45 a_217_1050.n0 GND 0.31fF
C46 a_217_1050.n1 GND 0.38fF
C47 a_217_1050.n2 GND 0.31fF
C48 a_217_1050.n3 GND 0.36fF
C49 a_217_1050.n4 GND 0.88fF
C50 a_217_1050.n5 GND 0.03fF
C51 a_217_1050.n6 GND 0.04fF
C52 a_217_1050.n7 GND 0.03fF
C53 a_217_1050.n8 GND 0.18fF
C54 a_217_1050.n9 GND 0.33fF
C55 a_217_1050.n10 GND 0.49fF
C56 a_217_1050.n11 GND 0.28fF
C57 a_217_1050.n12 GND 0.41fF
C58 a_2000_210.n0 GND 0.07fF
C59 a_2000_210.n1 GND 0.09fF
C60 a_2000_210.n2 GND 0.13fF
C61 a_2000_210.n3 GND 0.11fF
C62 a_2000_210.n4 GND 0.02fF
C63 a_2000_210.n5 GND 0.03fF
C64 a_2000_210.n6 GND 0.02fF
C65 a_2000_210.n7 GND 0.05fF
C66 a_2000_210.n8 GND 0.03fF
C67 a_2000_210.n9 GND 0.11fF
C68 a_2000_210.n10 GND 0.06fF
C69 a_2000_210.n11 GND 0.01fF
C70 a_2000_210.t0 GND 0.33fF
C71 a_1905_1050.n0 GND 0.39fF
C72 a_1905_1050.n1 GND 0.50fF
C73 a_1905_1050.n2 GND 0.04fF
C74 a_1905_1050.n3 GND 0.05fF
C75 a_1905_1050.n4 GND 0.03fF
C76 a_1905_1050.n5 GND 0.21fF
C77 a_1905_1050.n6 GND 0.56fF
C78 a_1905_1050.n7 GND 0.48fF
C79 a_1905_1050.n8 GND 0.56fF
C80 a_1905_1050.n9 GND 0.18fF
C81 a_1905_1050.n10 GND 0.33fF
C82 a_1905_1050.n11 GND 0.48fF
C83 a_343_411.n0 GND 0.39fF
C84 a_343_411.n1 GND 0.60fF
C85 a_343_411.n2 GND 0.35fF
C86 a_343_411.t11 GND 0.74fF
C87 a_343_411.n3 GND 0.51fF
C88 a_343_411.n4 GND 3.15fF
C89 a_343_411.n5 GND 0.05fF
C90 a_343_411.n6 GND 0.07fF
C91 a_343_411.n7 GND 0.04fF
C92 a_343_411.n8 GND 0.46fF
C93 a_343_411.n9 GND 0.57fF
C94 a_343_411.n10 GND 0.68fF
C95 a_343_411.n11 GND 0.79fF
C96 a_343_411.n12 GND 0.25fF
C97 a_343_411.n13 GND 0.31fF
C98 a_343_411.n14 GND 0.68fF
C99 a_1265_989.n0 GND 0.07fF
C100 a_1265_989.n1 GND 0.64fF
C101 a_1265_989.n2 GND 0.76fF
C102 a_1265_989.n3 GND 0.33fF
C103 a_1265_989.n4 GND 0.42fF
C104 a_1265_989.t13 GND 0.68fF
C105 a_1265_989.n5 GND 0.50fF
C106 a_1265_989.n6 GND 0.42fF
C107 a_1265_989.t6 GND 0.68fF
C108 a_1265_989.n7 GND 0.45fF
C109 a_1265_989.n8 GND 0.42fF
C110 a_1265_989.t9 GND 0.68fF
C111 a_1265_989.n9 GND 0.47fF
C112 a_1265_989.n10 GND 1.37fF
C113 a_1265_989.n11 GND 1.85fF
C114 a_1265_989.n12 GND 0.51fF
C115 a_1265_989.n13 GND 0.03fF
C116 a_1265_989.n14 GND 0.40fF
C117 a_1265_989.n15 GND 0.05fF
C118 a_4294_210.n0 GND 0.02fF
C119 a_4294_210.n1 GND 0.09fF
C120 a_4294_210.n2 GND 0.13fF
C121 a_4294_210.n3 GND 0.11fF
C122 a_4294_210.t1 GND 0.29fF
C123 a_4294_210.n4 GND 0.09fF
C124 a_4294_210.n5 GND 0.05fF
C125 a_4294_210.n6 GND 0.01fF
C126 a_4294_210.n7 GND 0.03fF
C127 a_4294_210.n8 GND 0.11fF
C128 a_4294_210.n9 GND 0.02fF
C129 a_4294_210.n10 GND 0.05fF
C130 a_4294_210.n11 GND 0.02fF
C131 a_4013_103.n0 GND 0.03fF
C132 a_4013_103.n1 GND 0.10fF
C133 a_4013_103.n2 GND 0.10fF
C134 a_4013_103.n3 GND 0.05fF
C135 a_4013_103.n4 GND 0.03fF
C136 a_4013_103.n5 GND 0.04fF
C137 a_4013_103.n6 GND 0.11fF
C138 a_4013_103.n7 GND 0.04fF
C139 SN.n0 GND 0.47fF
C140 SN.t0 GND 0.43fF
C141 SN.n1 GND 0.45fF
C142 SN.n2 GND 0.47fF
C143 SN.t4 GND 0.43fF
C144 SN.n3 GND 0.35fF
C145 SN.n4 GND 1.78fF
C146 a_3599_411.n0 GND 0.55fF
C147 a_3599_411.n1 GND 0.55fF
C148 a_3599_411.n2 GND 0.34fF
C149 a_3599_411.n3 GND 0.88fF
C150 a_3599_411.n4 GND 0.04fF
C151 a_3599_411.n5 GND 0.06fF
C152 a_3599_411.n6 GND 0.03fF
C153 a_3599_411.n7 GND 0.31fF
C154 a_3599_411.n8 GND 0.95fF
C155 a_3599_411.n9 GND 0.31fF
C156 a_3599_411.n10 GND 0.20fF
C157 a_3599_411.n11 GND 0.65fF
C158 VDD.n0 GND 0.20fF
C159 VDD.n1 GND 0.02fF
C160 VDD.n2 GND 0.02fF
C161 VDD.n3 GND 0.04fF
C162 VDD.n4 GND 0.01fF
C163 VDD.n5 GND 0.02fF
C164 VDD.n6 GND 0.02fF
C165 VDD.n8 GND 0.02fF
C166 VDD.n9 GND 0.02fF
C167 VDD.n12 GND 0.02fF
C168 VDD.n14 GND 0.45fF
C169 VDD.n16 GND 0.03fF
C170 VDD.n17 GND 0.02fF
C171 VDD.n18 GND 0.02fF
C172 VDD.n19 GND 0.02fF
C173 VDD.n20 GND 0.03fF
C174 VDD.n21 GND 0.27fF
C175 VDD.n22 GND 0.02fF
C176 VDD.n23 GND 0.03fF
C177 VDD.n24 GND 0.22fF
C178 VDD.n25 GND 0.01fF
C179 VDD.n26 GND 0.13fF
C180 VDD.n27 GND 0.16fF
C181 VDD.n28 GND 0.01fF
C182 VDD.n29 GND 0.02fF
C183 VDD.n30 GND 0.07fF
C184 VDD.n31 GND 0.27fF
C185 VDD.n32 GND 0.01fF
C186 VDD.n33 GND 0.02fF
C187 VDD.n34 GND 0.00fF
C188 VDD.n35 GND 0.09fF
C189 VDD.n36 GND 0.02fF
C190 VDD.n37 GND 0.13fF
C191 VDD.n38 GND 0.16fF
C192 VDD.n39 GND 0.01fF
C193 VDD.n40 GND 0.10fF
C194 VDD.n41 GND 0.02fF
C195 VDD.n42 GND 0.02fF
C196 VDD.n43 GND 0.02fF
C197 VDD.n44 GND 0.17fF
C198 VDD.n45 GND 0.14fF
C199 VDD.n46 GND 0.01fF
C200 VDD.n47 GND 0.02fF
C201 VDD.n48 GND 0.03fF
C202 VDD.n49 GND 0.17fF
C203 VDD.n50 GND 0.14fF
C204 VDD.n51 GND 0.01fF
C205 VDD.n52 GND 0.02fF
C206 VDD.n53 GND 0.03fF
C207 VDD.n54 GND 0.10fF
C208 VDD.n55 GND 0.02fF
C209 VDD.n56 GND 0.13fF
C210 VDD.n57 GND 0.15fF
C211 VDD.n58 GND 0.01fF
C212 VDD.n59 GND 0.02fF
C213 VDD.n60 GND 0.02fF
C214 VDD.n61 GND 0.13fF
C215 VDD.n62 GND 0.16fF
C216 VDD.n63 GND 0.01fF
C217 VDD.n64 GND 0.02fF
C218 VDD.n65 GND 0.02fF
C219 VDD.n66 GND 0.06fF
C220 VDD.n67 GND 0.22fF
C221 VDD.n68 GND 0.01fF
C222 VDD.n69 GND 0.01fF
C223 VDD.n70 GND 0.02fF
C224 VDD.n71 GND 0.27fF
C225 VDD.n72 GND 0.01fF
C226 VDD.n73 GND 0.02fF
C227 VDD.n74 GND 0.02fF
C228 VDD.n75 GND 0.27fF
C229 VDD.n76 GND 0.01fF
C230 VDD.n77 GND 0.02fF
C231 VDD.n78 GND 0.03fF
C232 VDD.n79 GND 0.02fF
C233 VDD.n80 GND 0.02fF
C234 VDD.n81 GND 0.02fF
C235 VDD.n82 GND 0.26fF
C236 VDD.n83 GND 0.04fF
C237 VDD.n84 GND 0.03fF
C238 VDD.n85 GND 0.02fF
C239 VDD.n87 GND 0.02fF
C240 VDD.n88 GND 0.02fF
C241 VDD.n89 GND 0.02fF
C242 VDD.n90 GND 0.02fF
C243 VDD.n92 GND 0.02fF
C244 VDD.n93 GND 0.02fF
C245 VDD.n94 GND 0.02fF
C246 VDD.n96 GND 0.27fF
C247 VDD.n98 GND 0.02fF
C248 VDD.n99 GND 0.02fF
C249 VDD.n100 GND 0.03fF
C250 VDD.n101 GND 0.02fF
C251 VDD.n102 GND 0.27fF
C252 VDD.n103 GND 0.01fF
C253 VDD.n104 GND 0.02fF
C254 VDD.n105 GND 0.03fF
C255 VDD.n106 GND 0.05fF
C256 VDD.n107 GND 0.24fF
C257 VDD.n108 GND 0.01fF
C258 VDD.n109 GND 0.01fF
C259 VDD.n110 GND 0.02fF
C260 VDD.n111 GND 0.13fF
C261 VDD.n112 GND 0.16fF
C262 VDD.n113 GND 0.01fF
C263 VDD.n114 GND 0.02fF
C264 VDD.n115 GND 0.02fF
C265 VDD.n116 GND 0.10fF
C266 VDD.n117 GND 0.02fF
C267 VDD.n118 GND 0.30fF
C268 VDD.n119 GND 0.01fF
C269 VDD.n120 GND 0.02fF
C270 VDD.n121 GND 0.03fF
C271 VDD.n122 GND 0.17fF
C272 VDD.n123 GND 0.14fF
C273 VDD.n124 GND 0.01fF
C274 VDD.n125 GND 0.02fF
C275 VDD.n126 GND 0.03fF
C276 VDD.n127 GND 0.13fF
C277 VDD.n128 GND 0.16fF
C278 VDD.n129 GND 0.01fF
C279 VDD.n130 GND 0.02fF
C280 VDD.n131 GND 0.02fF
C281 VDD.n132 GND 0.06fF
C282 VDD.n133 GND 0.24fF
C283 VDD.n134 GND 0.01fF
C284 VDD.n135 GND 0.01fF
C285 VDD.n136 GND 0.02fF
C286 VDD.n137 GND 0.27fF
C287 VDD.n138 GND 0.01fF
C288 VDD.n139 GND 0.02fF
C289 VDD.n140 GND 0.03fF
C290 VDD.n141 GND 0.02fF
C291 VDD.n142 GND 0.02fF
C292 VDD.n143 GND 0.02fF
C293 VDD.n144 GND 0.21fF
C294 VDD.n145 GND 0.04fF
C295 VDD.n146 GND 0.03fF
C296 VDD.n147 GND 0.02fF
C297 VDD.n148 GND 0.02fF
C298 VDD.n149 GND 0.02fF
C299 VDD.n150 GND 0.02fF
C300 VDD.n151 GND 0.02fF
C301 VDD.n153 GND 0.02fF
C302 VDD.n154 GND 0.02fF
C303 VDD.n155 GND 0.02fF
C304 VDD.n157 GND 0.27fF
C305 VDD.n159 GND 0.02fF
C306 VDD.n160 GND 0.02fF
C307 VDD.n161 GND 0.03fF
C308 VDD.n162 GND 0.02fF
C309 VDD.n163 GND 0.27fF
C310 VDD.n164 GND 0.01fF
C311 VDD.n165 GND 0.02fF
C312 VDD.n166 GND 0.03fF
C313 VDD.n167 GND 0.05fF
C314 VDD.n168 GND 0.24fF
C315 VDD.n169 GND 0.01fF
C316 VDD.n170 GND 0.01fF
C317 VDD.n171 GND 0.02fF
C318 VDD.n172 GND 0.13fF
C319 VDD.n173 GND 0.16fF
C320 VDD.n174 GND 0.01fF
C321 VDD.n175 GND 0.02fF
C322 VDD.n176 GND 0.02fF
C323 VDD.n177 GND 0.10fF
C324 VDD.n178 GND 0.02fF
C325 VDD.n179 GND 0.30fF
C326 VDD.n180 GND 0.01fF
C327 VDD.n181 GND 0.02fF
C328 VDD.n182 GND 0.03fF
C329 VDD.n183 GND 0.17fF
C330 VDD.n184 GND 0.14fF
C331 VDD.n185 GND 0.01fF
C332 VDD.n186 GND 0.02fF
C333 VDD.n187 GND 0.03fF
C334 VDD.n188 GND 0.13fF
C335 VDD.n189 GND 0.16fF
C336 VDD.n190 GND 0.01fF
C337 VDD.n191 GND 0.02fF
C338 VDD.n192 GND 0.02fF
C339 VDD.n193 GND 0.06fF
C340 VDD.n194 GND 0.24fF
C341 VDD.n195 GND 0.01fF
C342 VDD.n196 GND 0.01fF
C343 VDD.n197 GND 0.02fF
C344 VDD.n198 GND 0.27fF
C345 VDD.n199 GND 0.01fF
C346 VDD.n200 GND 0.02fF
C347 VDD.n201 GND 0.03fF
C348 VDD.n202 GND 0.02fF
C349 VDD.n203 GND 0.02fF
C350 VDD.n204 GND 0.02fF
C351 VDD.n205 GND 0.26fF
C352 VDD.n206 GND 0.04fF
C353 VDD.n207 GND 0.03fF
C354 VDD.n208 GND 0.02fF
C355 VDD.n209 GND 0.02fF
C356 VDD.n210 GND 0.02fF
C357 VDD.n211 GND 0.02fF
C358 VDD.n212 GND 0.02fF
C359 VDD.n214 GND 0.02fF
C360 VDD.n215 GND 0.02fF
C361 VDD.n216 GND 0.02fF
C362 VDD.n218 GND 0.27fF
C363 VDD.n220 GND 0.02fF
C364 VDD.n221 GND 0.02fF
C365 VDD.n222 GND 0.03fF
C366 VDD.n223 GND 0.02fF
C367 VDD.n224 GND 0.27fF
C368 VDD.n225 GND 0.01fF
C369 VDD.n226 GND 0.02fF
C370 VDD.n227 GND 0.03fF
C371 VDD.n228 GND 0.27fF
C372 VDD.n229 GND 0.01fF
C373 VDD.n230 GND 0.02fF
C374 VDD.n231 GND 0.01fF
C375 VDD.n232 GND 0.02fF
C376 VDD.n233 GND 0.02fF
C377 VDD.n234 GND 0.02fF
C378 VDD.n235 GND 0.15fF
C379 VDD.n236 GND 0.03fF
C380 VDD.n237 GND 0.02fF
C381 VDD.n238 GND 0.02fF
C382 VDD.n239 GND 0.02fF
C383 VDD.n240 GND 0.02fF
C384 VDD.n241 GND 0.02fF
C385 VDD.n243 GND 0.02fF
C386 VDD.n244 GND 0.02fF
C387 VDD.n245 GND 0.02fF
C388 VDD.n247 GND 0.45fF
C389 VDD.n249 GND 0.03fF
C390 VDD.n250 GND 0.03fF
C391 VDD.n251 GND 0.27fF
C392 VDD.n252 GND 0.02fF
C393 VDD.n253 GND 0.03fF
C394 VDD.n254 GND 0.03fF
C395 VDD.n255 GND 0.06fF
C396 VDD.n256 GND 0.24fF
C397 VDD.n257 GND 0.01fF
C398 VDD.n258 GND 0.01fF
C399 VDD.n259 GND 0.02fF
C400 VDD.n260 GND 0.13fF
C401 VDD.n261 GND 0.16fF
C402 VDD.n262 GND 0.01fF
C403 VDD.n263 GND 0.02fF
C404 VDD.n264 GND 0.02fF
C405 VDD.n265 GND 0.17fF
C406 VDD.n266 GND 0.14fF
C407 VDD.n267 GND 0.01fF
C408 VDD.n268 GND 0.02fF
C409 VDD.n269 GND 0.03fF
C410 VDD.n270 GND 0.10fF
C411 VDD.n271 GND 0.02fF
C412 VDD.n272 GND 0.30fF
C413 VDD.n273 GND 0.01fF
C414 VDD.n274 GND 0.02fF
C415 VDD.n275 GND 0.03fF
C416 VDD.n276 GND 0.13fF
C417 VDD.n277 GND 0.16fF
C418 VDD.n278 GND 0.01fF
C419 VDD.n279 GND 0.02fF
C420 VDD.n280 GND 0.02fF
C421 VDD.n281 GND 0.05fF
C422 VDD.n282 GND 0.24fF
C423 VDD.n283 GND 0.01fF
C424 VDD.n284 GND 0.01fF
C425 VDD.n285 GND 0.02fF
C426 VDD.n286 GND 0.27fF
C427 VDD.n287 GND 0.01fF
C428 VDD.n288 GND 0.02fF
C429 VDD.n289 GND 0.03fF
C430 VDD.n290 GND 0.02fF
C431 VDD.n291 GND 0.02fF
C432 VDD.n292 GND 0.02fF
C433 VDD.n293 GND 0.02fF
C434 VDD.n294 GND 0.02fF
C435 VDD.n295 GND 0.02fF
C436 VDD.n297 GND 0.02fF
C437 VDD.n298 GND 0.02fF
C438 VDD.n299 GND 0.02fF
C439 VDD.n300 GND 0.02fF
C440 VDD.n302 GND 0.03fF
C441 VDD.n303 GND 0.02fF
C442 VDD.n304 GND 0.26fF
C443 VDD.n305 GND 0.04fF
C444 VDD.n307 GND 0.27fF
C445 VDD.n309 GND 0.02fF
C446 VDD.n310 GND 0.02fF
C447 VDD.n311 GND 0.03fF
C448 VDD.n312 GND 0.02fF
C449 VDD.n313 GND 0.27fF
C450 VDD.n314 GND 0.01fF
C451 VDD.n315 GND 0.02fF
C452 VDD.n316 GND 0.03fF
C453 VDD.n317 GND 0.27fF
C454 VDD.n318 GND 0.01fF
C455 VDD.n319 GND 0.02fF
C456 VDD.n320 GND 0.02fF
C457 VDD.n321 GND 0.06fF
C458 VDD.n322 GND 0.22fF
C459 VDD.n323 GND 0.01fF
C460 VDD.n324 GND 0.01fF
C461 VDD.n325 GND 0.02fF
C462 VDD.n326 GND 0.13fF
C463 VDD.n327 GND 0.16fF
C464 VDD.n328 GND 0.01fF
C465 VDD.n329 GND 0.02fF
C466 VDD.n330 GND 0.02fF
C467 VDD.n331 GND 0.10fF
C468 VDD.n332 GND 0.02fF
C469 VDD.n333 GND 0.13fF
C470 VDD.n334 GND 0.15fF
C471 VDD.n335 GND 0.01fF
C472 VDD.n336 GND 0.02fF
C473 VDD.n337 GND 0.02fF
C474 VDD.n338 GND 0.17fF
C475 VDD.n339 GND 0.14fF
C476 VDD.n340 GND 0.01fF
C477 VDD.n341 GND 0.02fF
C478 VDD.n342 GND 0.03fF
C479 VDD.n343 GND 0.17fF
C480 VDD.n344 GND 0.14fF
C481 VDD.n345 GND 0.01fF
C482 VDD.n346 GND 0.02fF
C483 VDD.n347 GND 0.03fF
C484 VDD.n348 GND 0.13fF
C485 VDD.n349 GND 0.16fF
C486 VDD.n350 GND 0.01fF
C487 VDD.n351 GND 0.10fF
C488 VDD.n352 GND 0.02fF
C489 VDD.n353 GND 0.02fF
C490 VDD.n354 GND 0.02fF
C491 VDD.n355 GND 0.13fF
C492 VDD.n356 GND 0.16fF
C493 VDD.n357 GND 0.01fF
C494 VDD.n358 GND 0.02fF
C495 VDD.n359 GND 0.02fF
C496 VDD.n360 GND 0.22fF
C497 VDD.n361 GND 0.01fF
C498 VDD.n362 GND 0.07fF
C499 VDD.n363 GND 0.02fF
C500 VDD.n364 GND 0.27fF
C501 VDD.n365 GND 0.01fF
C502 VDD.n366 GND 0.02fF
C503 VDD.n367 GND 0.02fF
C504 VDD.n368 GND 0.27fF
C505 VDD.n369 GND 0.01fF
C506 VDD.n370 GND 0.02fF
C507 VDD.n371 GND 0.03fF
C508 VDD.n372 GND 0.02fF
C509 VDD.n373 GND 0.02fF
C510 VDD.n374 GND 0.02fF
C511 VDD.n375 GND 0.30fF
C512 VDD.n376 GND 0.04fF
C513 VDD.n377 GND 0.03fF
C514 VDD.n378 GND 0.02fF
C515 VDD.n379 GND 0.02fF
C516 VDD.n380 GND 0.02fF
C517 VDD.n381 GND 0.02fF
C518 VDD.n382 GND 0.02fF
C519 VDD.n384 GND 0.02fF
C520 VDD.n385 GND 0.02fF
C521 VDD.n386 GND 0.02fF
C522 VDD.n388 GND 0.27fF
C523 VDD.n390 GND 0.02fF
C524 VDD.n391 GND 0.02fF
C525 VDD.n392 GND 0.03fF
C526 VDD.n393 GND 0.02fF
C527 VDD.n394 GND 0.27fF
C528 VDD.n395 GND 0.01fF
C529 VDD.n396 GND 0.02fF
C530 VDD.n397 GND 0.03fF
C531 VDD.n398 GND 0.27fF
C532 VDD.n399 GND 0.01fF
C533 VDD.n400 GND 0.02fF
C534 VDD.n401 GND 0.02fF
C535 VDD.n402 GND 0.06fF
C536 VDD.n403 GND 0.22fF
C537 VDD.n404 GND 0.01fF
C538 VDD.n405 GND 0.01fF
C539 VDD.n406 GND 0.02fF
C540 VDD.n407 GND 0.13fF
C541 VDD.n408 GND 0.16fF
C542 VDD.n409 GND 0.01fF
C543 VDD.n410 GND 0.02fF
C544 VDD.n411 GND 0.02fF
C545 VDD.n412 GND 0.10fF
C546 VDD.n413 GND 0.02fF
C547 VDD.n414 GND 0.13fF
C548 VDD.n415 GND 0.15fF
C549 VDD.n416 GND 0.01fF
C550 VDD.n417 GND 0.02fF
C551 VDD.n418 GND 0.02fF
C552 VDD.n419 GND 0.17fF
C553 VDD.n420 GND 0.14fF
C554 VDD.n421 GND 0.01fF
C555 VDD.n422 GND 0.02fF
C556 VDD.n423 GND 0.03fF
C557 VDD.n424 GND 0.17fF
C558 VDD.n425 GND 0.14fF
C559 VDD.n426 GND 0.01fF
C560 VDD.n427 GND 0.02fF
C561 VDD.n428 GND 0.03fF
C562 VDD.n429 GND 0.13fF
C563 VDD.n430 GND 0.16fF
C564 VDD.n431 GND 0.01fF
C565 VDD.n432 GND 0.10fF
C566 VDD.n433 GND 0.02fF
C567 VDD.n434 GND 0.02fF
C568 VDD.n435 GND 0.02fF
C569 VDD.n436 GND 0.13fF
C570 VDD.n437 GND 0.16fF
C571 VDD.n438 GND 0.01fF
C572 VDD.n439 GND 0.02fF
C573 VDD.n440 GND 0.02fF
C574 VDD.n441 GND 0.22fF
C575 VDD.n442 GND 0.01fF
C576 VDD.n443 GND 0.07fF
C577 VDD.n444 GND 0.02fF
C578 QN.n0 GND 0.35fF
C579 QN.n1 GND 0.45fF
C580 QN.n2 GND 0.51fF
C581 QN.n3 GND 0.60fF
C582 QN.n4 GND 0.32fF
C583 QN.n5 GND 0.35fF
C584 QN.n6 GND 0.44fF
C585 QN.n7 GND 0.03fF
.ends
