* SPICE3 file created from TMRDFFQX1.ext - technology: sky130A

.subckt TMRDFFQX1 Q D CLK VPB
M1000 a_13093_1005.t5 a_11887_383.t5 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=96.4069p ps=682.92u
M1001 VPB a_147_159.t5 a_1845_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_6137_1004.t4 a_4891_943.t5 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB a_4569_1004.t7 a_4891_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_13093_1005.t3 a_11887_383.t6 a_13757_1005.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPB a_4439_159.t6 a_7595_383.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPB a_147_159.t6 a_277_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPB a_6137_1004.t5 a_4439_159.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPB a_8861_1004.t11 a_11656_73.t0 nshort w=-1.605u l=1.765u
+  ad=71.008p pd=467.45u as=0p ps=0u
M1009 VPB a_8731_159.t5 a_8861_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_3177_1004.t3 a_277_1004.t7 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_15059_182.t2 a_13268_181.t7 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB a_1845_1004.t5 a_147_159.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_11887_383.t4 a_11761_1004.t5 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPB D a_9183_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPB a_10429_1004.t5 a_10990_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPB a_8731_159.t9 a_8675_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPB D a_4891_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPB a_7469_1004.t5 a_7595_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPB CLK a_277_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPB a_4569_1004.t8 a_5366_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPB a_599_943.t5 a_1740_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_13757_1005.t0 a_7595_383.t5 a_13268_181.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPB a_11887_383.t7 a_13654_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_3177_1004.t0 a_3303_383.t5 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPB CLK a_147_159.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_11887_383.t1 a_8731_159.t6 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPB a_11887_383.t9 a_11761_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPB a_11887_383.t8 a_12988_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPB CLK a_4439_159.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_9183_943.t2 D VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_3303_383.t1 a_3177_1004.t6 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPB a_599_943.t6 a_277_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPB a_147_159.t13 a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPB a_277_1004.t8 a_599_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_8731_159.t1 a_10429_1004.t6 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_4569_1004.t4 a_4891_943.t6 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_13757_1005.t2 a_3303_383.t6 a_13268_181.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPB a_9183_943.t7 a_10429_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPB a_147_159.t7 a_3303_383.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_7595_383.t4 a_7469_1004.t6 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPB a_4569_1004.t9 a_7364_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPB a_3177_1004.t5 a_3738_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1043 VPB a_4569_1004.t10 a_7469_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPB a_9183_943.t5 a_10324_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_4439_159.t2 CLK VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_1845_1004.t3 a_147_159.t8 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_8861_1004.t1 a_9183_943.t8 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 VPB a_4439_159.t8 a_4569_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_6137_1004.t1 a_4439_159.t9 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_9183_943.t1 a_8861_1004.t7 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1051 VPB a_4439_159.t5 a_4383_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1052 a_13093_1005.t2 a_3303_383.t7 a_13757_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 a_11761_1004.t3 a_11887_383.t11 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_3303_383.t3 a_147_159.t10 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 VPB a_7595_383.t6 a_13093_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 VPB a_277_1004.t9 a_1074_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1057 VPB D a_599_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_13757_1005.t5 a_11887_383.t12 a_13093_1005.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1059 a_8731_159.t4 CLK VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1060 VPB a_8731_159.t7 a_10429_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 a_277_1004.t3 a_147_159.t11 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 a_4439_159.t0 a_6137_1004.t6 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 VPB a_7595_383.t7 a_7469_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1064 VPB CLK a_4569_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 VPB a_599_943.t7 a_1845_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 a_11761_1004.t1 a_8861_1004.t8 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1067 VPB a_11761_1004.t6 a_12322_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1068 VPB a_11887_383.t13 a_13093_1005.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 a_4891_943.t2 D VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 a_13757_1005.t7 a_3303_383.t10 a_13093_1005.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 a_277_1004.t5 CLK VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1072 VPB a_6137_1004.t7 a_6698_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1073 VPB a_277_1004.t10 a_3072_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1074 VPB a_4891_943.t8 a_4569_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 VPB a_277_1004.t11 a_3177_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1076 a_147_159.t3 CLK VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 VPB a_13268_181.t9 a_15059_182.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1078 VPB a_11761_1004.t7 a_11887_383.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 VPB a_4891_943.t7 a_6032_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1080 VPB a_3303_383.t9 a_14320_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1081 a_4891_943.t0 a_4569_1004.t11 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1082 a_7595_383.t1 a_4439_159.t10 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_277_1004.t1 a_599_943.t8 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 a_599_943.t0 a_277_1004.t12 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 a_8861_1004.t3 a_8731_159.t10 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_13268_181.t5 a_3303_383.t11 a_13757_1005.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 VPB CLK a_8731_159.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 a_10429_1004.t1 a_9183_943.t9 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 a_147_159.t0 a_1845_1004.t6 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 a_7469_1004.t0 a_4569_1004.t12 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 VPB a_3303_383.t12 a_3177_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1092 VPB a_8731_159.t12 a_11887_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1093 VPB CLK a_8861_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 a_4569_1004.t0 a_4439_159.t11 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1095 VPB a_4891_943.t9 a_6137_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1096 VPB a_7469_1004.t7 a_8030_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1097 VPB a_8861_1004.t10 a_11761_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 VPB a_3177_1004.t7 a_3303_383.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1099 a_13093_1005.t0 a_7595_383.t10 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 a_599_943.t3 D VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1101 VPB a_10429_1004.t7 a_8731_159.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 VPB a_1845_1004.t7 a_2406_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_13268_181.t3 a_7595_383.t11 a_13757_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 a_10429_1004.t2 a_8731_159.t13 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 a_7469_1004.t3 a_7595_383.t12 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 VPB a_8861_1004.t9 a_9658_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1107 VPB a_9183_943.t10 a_8861_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 a_4569_1004.t5 CLK VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 VPB a_4439_159.t13 a_6137_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 VPB a_8861_1004.t12 a_9183_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 a_1845_1004.t0 a_599_943.t10 VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1112 a_8861_1004.t5 CLK VPB pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u

R0 a_10429_1004.n3 a_10429_1004.t7 480.392
R1 a_10429_1004.n3 a_10429_1004.t6 403.272
R2 a_10429_1004.n4 a_10429_1004.t5 266.974
R3 a_10429_1004.n7 a_10429_1004.n5 200.608
R4 a_10429_1004.n5 a_10429_1004.n2 162.547
R5 a_10429_1004.n5 a_10429_1004.n4 153.315
R6 a_10429_1004.n4 a_10429_1004.n3 108.494
R7 a_10429_1004.n2 a_10429_1004.n1 76.002
R8 a_10429_1004.n7 a_10429_1004.n6 15.218
R9 a_10429_1004.n0 a_10429_1004.t3 14.282
R10 a_10429_1004.n0 a_10429_1004.t2 14.282
R11 a_10429_1004.n1 a_10429_1004.t4 14.282
R12 a_10429_1004.n1 a_10429_1004.t1 14.282
R13 a_10429_1004.n2 a_10429_1004.n0 12.85
R14 a_10429_1004.n8 a_10429_1004.n7 12.014
R15 a_10990_73.n5 a_10990_73.n4 24.877
R16 a_10990_73.t0 a_10990_73.n5 12.677
R17 a_10990_73.t0 a_10990_73.n3 11.595
R18 a_10990_73.t0 a_10990_73.n6 8.137
R19 a_10990_73.n2 a_10990_73.n0 4.031
R20 a_10990_73.n2 a_10990_73.n1 3.644
R21 a_10990_73.t0 a_10990_73.n2 1.093
R22 a_4439_159.n8 a_4439_159.t8 512.525
R23 a_4439_159.n6 a_4439_159.t13 472.359
R24 a_4439_159.n4 a_4439_159.t6 472.359
R25 a_4439_159.n6 a_4439_159.t9 384.527
R26 a_4439_159.n4 a_4439_159.t10 384.527
R27 a_4439_159.n8 a_4439_159.t11 371.139
R28 a_4439_159.n9 a_4439_159.t5 324.268
R29 a_4439_159.n7 a_4439_159.t12 277.772
R30 a_4439_159.n5 a_4439_159.t7 277.772
R31 a_4439_159.n14 a_4439_159.n12 247.192
R32 a_4439_159.n9 a_4439_159.n8 119.654
R33 a_4439_159.n12 a_4439_159.n3 109.441
R34 a_4439_159.n10 a_4439_159.n9 82.484
R35 a_4439_159.n11 a_4439_159.n5 80.307
R36 a_4439_159.n3 a_4439_159.n2 76.002
R37 a_4439_159.n10 a_4439_159.n7 76
R38 a_4439_159.n12 a_4439_159.n11 76
R39 a_4439_159.n7 a_4439_159.n6 67.001
R40 a_4439_159.n5 a_4439_159.n4 67.001
R41 a_4439_159.n14 a_4439_159.n13 30
R42 a_4439_159.n15 a_4439_159.n0 24.383
R43 a_4439_159.n15 a_4439_159.n14 23.684
R44 a_4439_159.n1 a_4439_159.t3 14.282
R45 a_4439_159.n1 a_4439_159.t2 14.282
R46 a_4439_159.n2 a_4439_159.t1 14.282
R47 a_4439_159.n2 a_4439_159.t0 14.282
R48 a_4439_159.n3 a_4439_159.n1 12.85
R49 a_4439_159.n11 a_4439_159.n10 2.947
R50 a_4383_75.n4 a_4383_75.n3 19.724
R51 a_4383_75.t0 a_4383_75.n5 11.595
R52 a_4383_75.t0 a_4383_75.n4 9.207
R53 a_4383_75.n2 a_4383_75.n0 8.543
R54 a_4383_75.t0 a_4383_75.n2 3.034
R55 a_4383_75.n2 a_4383_75.n1 0.443
R56 a_11887_383.n3 a_11887_383.t13 512.525
R57 a_11887_383.n4 a_11887_383.t6 477.179
R58 a_11887_383.n8 a_11887_383.t9 472.359
R59 a_11887_383.n4 a_11887_383.t12 406.485
R60 a_11887_383.n8 a_11887_383.t11 384.527
R61 a_11887_383.n3 a_11887_383.t5 371.139
R62 a_11887_383.n5 a_11887_383.t7 346.633
R63 a_11887_383.n7 a_11887_383.t8 287.1
R64 a_11887_383.n9 a_11887_383.t10 251.219
R65 a_11887_383.n13 a_11887_383.n11 227.161
R66 a_11887_383.n6 a_11887_383.n5 154.675
R67 a_11887_383.n11 a_11887_383.n2 135.994
R68 a_11887_383.n9 a_11887_383.n8 93.554
R69 a_11887_383.n6 a_11887_383.n3 89.615
R70 a_11887_383.n10 a_11887_383.n9 78.947
R71 a_11887_383.n10 a_11887_383.n7 77.043
R72 a_11887_383.n2 a_11887_383.n1 76.002
R73 a_11887_383.n11 a_11887_383.n10 76
R74 a_11887_383.n7 a_11887_383.n6 53.105
R75 a_11887_383.n5 a_11887_383.n4 29.194
R76 a_11887_383.n13 a_11887_383.n12 15.218
R77 a_11887_383.n0 a_11887_383.t3 14.282
R78 a_11887_383.n0 a_11887_383.t1 14.282
R79 a_11887_383.n1 a_11887_383.t2 14.282
R80 a_11887_383.n1 a_11887_383.t4 14.282
R81 a_11887_383.n2 a_11887_383.n0 12.85
R82 a_11887_383.n14 a_11887_383.n13 12.014
R83 a_13093_1005.n4 a_13093_1005.n3 195.987
R84 a_13093_1005.n2 a_13093_1005.t2 89.553
R85 a_13093_1005.n5 a_13093_1005.n4 75.27
R86 a_13093_1005.n3 a_13093_1005.n2 75.214
R87 a_13093_1005.n4 a_13093_1005.n0 36.519
R88 a_13093_1005.n3 a_13093_1005.t6 14.338
R89 a_13093_1005.n0 a_13093_1005.t1 14.282
R90 a_13093_1005.n0 a_13093_1005.t0 14.282
R91 a_13093_1005.n1 a_13093_1005.t7 14.282
R92 a_13093_1005.n1 a_13093_1005.t3 14.282
R93 a_13093_1005.n5 a_13093_1005.t4 14.282
R94 a_13093_1005.t5 a_13093_1005.n5 14.282
R95 a_13093_1005.n2 a_13093_1005.n1 12.119
R96 a_147_159.n8 a_147_159.t6 512.525
R97 a_147_159.n6 a_147_159.t5 472.359
R98 a_147_159.n4 a_147_159.t7 472.359
R99 a_147_159.n6 a_147_159.t8 384.527
R100 a_147_159.n4 a_147_159.t10 384.527
R101 a_147_159.n8 a_147_159.t11 371.139
R102 a_147_159.n9 a_147_159.t13 324.268
R103 a_147_159.n7 a_147_159.t9 277.772
R104 a_147_159.n5 a_147_159.t12 277.772
R105 a_147_159.n14 a_147_159.n12 247.192
R106 a_147_159.n9 a_147_159.n8 119.654
R107 a_147_159.n12 a_147_159.n3 109.441
R108 a_147_159.n10 a_147_159.n9 82.484
R109 a_147_159.n11 a_147_159.n5 80.307
R110 a_147_159.n3 a_147_159.n2 76.002
R111 a_147_159.n10 a_147_159.n7 76
R112 a_147_159.n12 a_147_159.n11 76
R113 a_147_159.n7 a_147_159.n6 67.001
R114 a_147_159.n5 a_147_159.n4 67.001
R115 a_147_159.n14 a_147_159.n13 30
R116 a_147_159.n15 a_147_159.n0 24.383
R117 a_147_159.n15 a_147_159.n14 23.684
R118 a_147_159.n1 a_147_159.t4 14.282
R119 a_147_159.n1 a_147_159.t3 14.282
R120 a_147_159.n2 a_147_159.t1 14.282
R121 a_147_159.n2 a_147_159.t0 14.282
R122 a_147_159.n3 a_147_159.n1 12.85
R123 a_147_159.n11 a_147_159.n10 2.947
R124 a_1845_1004.n4 a_1845_1004.t5 480.392
R125 a_1845_1004.n4 a_1845_1004.t6 403.272
R126 a_1845_1004.n5 a_1845_1004.t7 266.974
R127 a_1845_1004.n8 a_1845_1004.n6 194.086
R128 a_1845_1004.n6 a_1845_1004.n3 162.547
R129 a_1845_1004.n6 a_1845_1004.n5 153.315
R130 a_1845_1004.n5 a_1845_1004.n4 108.494
R131 a_1845_1004.n3 a_1845_1004.n2 76.002
R132 a_1845_1004.n8 a_1845_1004.n7 30
R133 a_1845_1004.n9 a_1845_1004.n0 24.383
R134 a_1845_1004.n9 a_1845_1004.n8 23.684
R135 a_1845_1004.n1 a_1845_1004.t4 14.282
R136 a_1845_1004.n1 a_1845_1004.t3 14.282
R137 a_1845_1004.n2 a_1845_1004.t1 14.282
R138 a_1845_1004.n2 a_1845_1004.t0 14.282
R139 a_1845_1004.n3 a_1845_1004.n1 12.85
R140 a_4891_943.n4 a_4891_943.t9 480.392
R141 a_4891_943.n6 a_4891_943.t6 454.685
R142 a_4891_943.n6 a_4891_943.t8 428.979
R143 a_4891_943.n4 a_4891_943.t5 403.272
R144 a_4891_943.n5 a_4891_943.t7 266.974
R145 a_4891_943.n7 a_4891_943.t10 221.453
R146 a_4891_943.n11 a_4891_943.n9 194.086
R147 a_4891_943.n9 a_4891_943.n3 162.547
R148 a_4891_943.n7 a_4891_943.n6 108.494
R149 a_4891_943.n5 a_4891_943.n4 108.494
R150 a_4891_943.n8 a_4891_943.n7 78.947
R151 a_4891_943.n8 a_4891_943.n5 77.315
R152 a_4891_943.n3 a_4891_943.n2 76.002
R153 a_4891_943.n9 a_4891_943.n8 76
R154 a_4891_943.n11 a_4891_943.n10 30
R155 a_4891_943.n12 a_4891_943.n0 24.383
R156 a_4891_943.n12 a_4891_943.n11 23.684
R157 a_4891_943.n1 a_4891_943.t3 14.282
R158 a_4891_943.n1 a_4891_943.t2 14.282
R159 a_4891_943.n2 a_4891_943.t1 14.282
R160 a_4891_943.n2 a_4891_943.t0 14.282
R161 a_4891_943.n3 a_4891_943.n1 12.85
R162 a_6137_1004.n4 a_6137_1004.t5 480.392
R163 a_6137_1004.n4 a_6137_1004.t6 403.272
R164 a_6137_1004.n5 a_6137_1004.t7 266.974
R165 a_6137_1004.n8 a_6137_1004.n6 194.086
R166 a_6137_1004.n6 a_6137_1004.n3 162.547
R167 a_6137_1004.n6 a_6137_1004.n5 153.315
R168 a_6137_1004.n5 a_6137_1004.n4 108.494
R169 a_6137_1004.n3 a_6137_1004.n2 76.002
R170 a_6137_1004.n8 a_6137_1004.n7 30
R171 a_6137_1004.n9 a_6137_1004.n0 24.383
R172 a_6137_1004.n9 a_6137_1004.n8 23.684
R173 a_6137_1004.n1 a_6137_1004.t0 14.282
R174 a_6137_1004.n1 a_6137_1004.t1 14.282
R175 a_6137_1004.n2 a_6137_1004.t3 14.282
R176 a_6137_1004.n2 a_6137_1004.t4 14.282
R177 a_6137_1004.n3 a_6137_1004.n1 12.85
R178 a_4569_1004.n8 a_4569_1004.t7 480.392
R179 a_4569_1004.n6 a_4569_1004.t10 480.392
R180 a_4569_1004.n8 a_4569_1004.t11 403.272
R181 a_4569_1004.n6 a_4569_1004.t12 403.272
R182 a_4569_1004.n9 a_4569_1004.t8 293.527
R183 a_4569_1004.n7 a_4569_1004.t9 293.527
R184 a_4569_1004.n13 a_4569_1004.n11 223.151
R185 a_4569_1004.n11 a_4569_1004.n5 154.293
R186 a_4569_1004.n10 a_4569_1004.n7 83.3
R187 a_4569_1004.n9 a_4569_1004.n8 81.941
R188 a_4569_1004.n7 a_4569_1004.n6 81.941
R189 a_4569_1004.n4 a_4569_1004.n3 79.232
R190 a_4569_1004.n11 a_4569_1004.n10 77.315
R191 a_4569_1004.n10 a_4569_1004.n9 76
R192 a_4569_1004.n5 a_4569_1004.n4 63.152
R193 a_4569_1004.n13 a_4569_1004.n12 30
R194 a_4569_1004.n14 a_4569_1004.n0 24.383
R195 a_4569_1004.n14 a_4569_1004.n13 23.684
R196 a_4569_1004.n5 a_4569_1004.n1 16.08
R197 a_4569_1004.n4 a_4569_1004.n2 16.08
R198 a_4569_1004.n1 a_4569_1004.t3 14.282
R199 a_4569_1004.n1 a_4569_1004.t4 14.282
R200 a_4569_1004.n2 a_4569_1004.t6 14.282
R201 a_4569_1004.n2 a_4569_1004.t5 14.282
R202 a_4569_1004.n3 a_4569_1004.t1 14.282
R203 a_4569_1004.n3 a_4569_1004.t0 14.282
R204 a_13757_1005.n4 a_13757_1005.n3 196.002
R205 a_13757_1005.n2 a_13757_1005.t0 89.553
R206 a_13757_1005.n5 a_13757_1005.n4 75.27
R207 a_13757_1005.n3 a_13757_1005.n2 75.214
R208 a_13757_1005.n4 a_13757_1005.n0 36.52
R209 a_13757_1005.n3 a_13757_1005.t4 14.338
R210 a_13757_1005.n0 a_13757_1005.t3 14.282
R211 a_13757_1005.n0 a_13757_1005.t7 14.282
R212 a_13757_1005.n1 a_13757_1005.t1 14.282
R213 a_13757_1005.n1 a_13757_1005.t2 14.282
R214 a_13757_1005.t6 a_13757_1005.n5 14.282
R215 a_13757_1005.n5 a_13757_1005.t5 14.282
R216 a_13757_1005.n2 a_13757_1005.n1 12.119
R217 a_7595_383.n5 a_7595_383.t5 475.572
R218 a_7595_383.n9 a_7595_383.t7 472.359
R219 a_7595_383.n4 a_7595_383.t6 469.145
R220 a_7595_383.n9 a_7595_383.t12 384.527
R221 a_7595_383.n5 a_7595_383.t11 384.527
R222 a_7595_383.n4 a_7595_383.t10 384.527
R223 a_7595_383.n6 a_7595_383.t13 277.772
R224 a_7595_383.n12 a_7595_383.n3 242.205
R225 a_7595_383.n10 a_7595_383.n9 201.031
R226 a_7595_383.n7 a_7595_383.n6 156.851
R227 a_7595_383.n10 a_7595_383.t9 141.018
R228 a_7595_383.n8 a_7595_383.t8 141.018
R229 a_7595_383.n8 a_7595_383.n7 134.03
R230 a_7595_383.n14 a_7595_383.n12 114.428
R231 a_7595_383.n3 a_7595_383.n2 76.002
R232 a_7595_383.n12 a_7595_383.n11 76
R233 a_7595_383.n6 a_7595_383.n5 67.889
R234 a_7595_383.n11 a_7595_383.n8 66.982
R235 a_7595_383.n7 a_7595_383.n4 66.88
R236 a_7595_383.n11 a_7595_383.n10 52.291
R237 a_7595_383.n14 a_7595_383.n13 30
R238 a_7595_383.n15 a_7595_383.n0 24.383
R239 a_7595_383.n15 a_7595_383.n14 23.684
R240 a_7595_383.n1 a_7595_383.t2 14.282
R241 a_7595_383.n1 a_7595_383.t1 14.282
R242 a_7595_383.n2 a_7595_383.t3 14.282
R243 a_7595_383.n2 a_7595_383.t4 14.282
R244 a_7595_383.n3 a_7595_383.n1 12.85
R245 a_277_1004.n7 a_277_1004.t8 480.392
R246 a_277_1004.n5 a_277_1004.t11 480.392
R247 a_277_1004.n7 a_277_1004.t12 403.272
R248 a_277_1004.n5 a_277_1004.t7 403.272
R249 a_277_1004.n8 a_277_1004.t9 293.527
R250 a_277_1004.n6 a_277_1004.t10 293.527
R251 a_277_1004.n12 a_277_1004.n10 229.673
R252 a_277_1004.n10 a_277_1004.n4 154.293
R253 a_277_1004.n9 a_277_1004.n6 83.3
R254 a_277_1004.n8 a_277_1004.n7 81.941
R255 a_277_1004.n6 a_277_1004.n5 81.941
R256 a_277_1004.n3 a_277_1004.n2 79.232
R257 a_277_1004.n10 a_277_1004.n9 77.315
R258 a_277_1004.n9 a_277_1004.n8 76
R259 a_277_1004.n4 a_277_1004.n3 63.152
R260 a_277_1004.n4 a_277_1004.n0 16.08
R261 a_277_1004.n3 a_277_1004.n1 16.08
R262 a_277_1004.n12 a_277_1004.n11 15.218
R263 a_277_1004.n0 a_277_1004.t0 14.282
R264 a_277_1004.n0 a_277_1004.t1 14.282
R265 a_277_1004.n1 a_277_1004.t6 14.282
R266 a_277_1004.n1 a_277_1004.t5 14.282
R267 a_277_1004.n2 a_277_1004.t4 14.282
R268 a_277_1004.n2 a_277_1004.t3 14.282
R269 a_277_1004.n13 a_277_1004.n12 12.014
R270 a_8030_73.t0 a_8030_73.n1 34.62
R271 a_8030_73.t0 a_8030_73.n0 8.137
R272 a_8030_73.t0 a_8030_73.n2 4.69
R273 a_8731_159.n7 a_8731_159.t5 512.525
R274 a_8731_159.n5 a_8731_159.t7 472.359
R275 a_8731_159.n3 a_8731_159.t12 472.359
R276 a_8731_159.n5 a_8731_159.t13 384.527
R277 a_8731_159.n3 a_8731_159.t6 384.527
R278 a_8731_159.n7 a_8731_159.t10 371.139
R279 a_8731_159.n8 a_8731_159.t9 324.268
R280 a_8731_159.n6 a_8731_159.t8 277.772
R281 a_8731_159.n4 a_8731_159.t11 277.772
R282 a_8731_159.n13 a_8731_159.n11 253.714
R283 a_8731_159.n8 a_8731_159.n7 119.654
R284 a_8731_159.n11 a_8731_159.n2 109.441
R285 a_8731_159.n9 a_8731_159.n8 82.484
R286 a_8731_159.n10 a_8731_159.n4 80.307
R287 a_8731_159.n2 a_8731_159.n1 76.002
R288 a_8731_159.n9 a_8731_159.n6 76
R289 a_8731_159.n11 a_8731_159.n10 76
R290 a_8731_159.n6 a_8731_159.n5 67.001
R291 a_8731_159.n4 a_8731_159.n3 67.001
R292 a_8731_159.n13 a_8731_159.n12 15.218
R293 a_8731_159.n0 a_8731_159.t3 14.282
R294 a_8731_159.n0 a_8731_159.t4 14.282
R295 a_8731_159.n1 a_8731_159.t0 14.282
R296 a_8731_159.n1 a_8731_159.t1 14.282
R297 a_8731_159.n2 a_8731_159.n0 12.85
R298 a_8731_159.n14 a_8731_159.n13 12.014
R299 a_8731_159.n10 a_8731_159.n9 2.947
R300 a_8861_1004.n7 a_8861_1004.t12 480.392
R301 a_8861_1004.n5 a_8861_1004.t10 480.392
R302 a_8861_1004.n7 a_8861_1004.t7 403.272
R303 a_8861_1004.n5 a_8861_1004.t8 403.272
R304 a_8861_1004.n8 a_8861_1004.t9 293.527
R305 a_8861_1004.n6 a_8861_1004.t11 293.527
R306 a_8861_1004.n12 a_8861_1004.n10 229.673
R307 a_8861_1004.n10 a_8861_1004.n4 154.293
R308 a_8861_1004.n9 a_8861_1004.n6 83.3
R309 a_8861_1004.n8 a_8861_1004.n7 81.941
R310 a_8861_1004.n6 a_8861_1004.n5 81.941
R311 a_8861_1004.n3 a_8861_1004.n2 79.232
R312 a_8861_1004.n10 a_8861_1004.n9 77.315
R313 a_8861_1004.n9 a_8861_1004.n8 76
R314 a_8861_1004.n4 a_8861_1004.n3 63.152
R315 a_8861_1004.n4 a_8861_1004.n0 16.08
R316 a_8861_1004.n3 a_8861_1004.n1 16.08
R317 a_8861_1004.n12 a_8861_1004.n11 15.218
R318 a_8861_1004.n0 a_8861_1004.t2 14.282
R319 a_8861_1004.n0 a_8861_1004.t1 14.282
R320 a_8861_1004.n1 a_8861_1004.t6 14.282
R321 a_8861_1004.n1 a_8861_1004.t5 14.282
R322 a_8861_1004.n2 a_8861_1004.t4 14.282
R323 a_8861_1004.n2 a_8861_1004.t3 14.282
R324 a_8861_1004.n13 a_8861_1004.n12 12.014
R325 a_5366_73.n12 a_5366_73.n11 26.811
R326 a_5366_73.n6 a_5366_73.n5 24.977
R327 a_5366_73.n2 a_5366_73.n1 24.877
R328 a_5366_73.t0 a_5366_73.n2 12.677
R329 a_5366_73.t0 a_5366_73.n3 11.595
R330 a_5366_73.t1 a_5366_73.n8 8.137
R331 a_5366_73.t0 a_5366_73.n4 7.273
R332 a_5366_73.t0 a_5366_73.n0 6.109
R333 a_5366_73.t1 a_5366_73.n7 4.864
R334 a_5366_73.t0 a_5366_73.n12 2.074
R335 a_5366_73.n7 a_5366_73.n6 1.13
R336 a_5366_73.n12 a_5366_73.t1 0.937
R337 a_5366_73.t1 a_5366_73.n10 0.804
R338 a_5366_73.n10 a_5366_73.n9 0.136
R339 a_599_943.n4 a_599_943.t7 480.392
R340 a_599_943.n6 a_599_943.t8 454.685
R341 a_599_943.n6 a_599_943.t6 428.979
R342 a_599_943.n4 a_599_943.t10 403.272
R343 a_599_943.n5 a_599_943.t5 266.974
R344 a_599_943.n7 a_599_943.t9 221.453
R345 a_599_943.n11 a_599_943.n9 194.086
R346 a_599_943.n9 a_599_943.n3 162.547
R347 a_599_943.n7 a_599_943.n6 108.494
R348 a_599_943.n5 a_599_943.n4 108.494
R349 a_599_943.n8 a_599_943.n7 78.947
R350 a_599_943.n8 a_599_943.n5 77.315
R351 a_599_943.n3 a_599_943.n2 76.002
R352 a_599_943.n9 a_599_943.n8 76
R353 a_599_943.n11 a_599_943.n10 30
R354 a_599_943.n12 a_599_943.n0 24.383
R355 a_599_943.n12 a_599_943.n11 23.684
R356 a_599_943.n1 a_599_943.t4 14.282
R357 a_599_943.n1 a_599_943.t3 14.282
R358 a_599_943.n2 a_599_943.t1 14.282
R359 a_599_943.n2 a_599_943.t0 14.282
R360 a_599_943.n3 a_599_943.n1 12.85
R361 a_1740_73.n12 a_1740_73.n11 26.811
R362 a_1740_73.n6 a_1740_73.n5 24.977
R363 a_1740_73.n2 a_1740_73.n1 24.877
R364 a_1740_73.t0 a_1740_73.n2 12.677
R365 a_1740_73.t0 a_1740_73.n3 11.595
R366 a_1740_73.t1 a_1740_73.n8 8.137
R367 a_1740_73.t0 a_1740_73.n4 7.273
R368 a_1740_73.t0 a_1740_73.n0 6.109
R369 a_1740_73.t1 a_1740_73.n7 4.864
R370 a_1740_73.t0 a_1740_73.n12 2.074
R371 a_1740_73.n7 a_1740_73.n6 1.13
R372 a_1740_73.n12 a_1740_73.t1 0.937
R373 a_1740_73.t1 a_1740_73.n10 0.804
R374 a_1740_73.n10 a_1740_73.n9 0.136
R375 a_3177_1004.n3 a_3177_1004.t7 480.392
R376 a_3177_1004.n3 a_3177_1004.t6 403.272
R377 a_3177_1004.n4 a_3177_1004.t5 293.527
R378 a_3177_1004.n7 a_3177_1004.n5 227.161
R379 a_3177_1004.n5 a_3177_1004.n4 153.315
R380 a_3177_1004.n5 a_3177_1004.n2 135.994
R381 a_3177_1004.n4 a_3177_1004.n3 81.941
R382 a_3177_1004.n2 a_3177_1004.n1 76.002
R383 a_3177_1004.n7 a_3177_1004.n6 15.218
R384 a_3177_1004.n0 a_3177_1004.t1 14.282
R385 a_3177_1004.n0 a_3177_1004.t0 14.282
R386 a_3177_1004.n1 a_3177_1004.t2 14.282
R387 a_3177_1004.n1 a_3177_1004.t3 14.282
R388 a_3177_1004.n2 a_3177_1004.n0 12.85
R389 a_3177_1004.n8 a_3177_1004.n7 12.014
R390 a_13268_181.n4 a_13268_181.t9 512.525
R391 a_13268_181.n4 a_13268_181.t7 371.139
R392 a_13268_181.n5 a_13268_181.t8 273.368
R393 a_13268_181.n16 a_13268_181.n6 226.775
R394 a_13268_181.n6 a_13268_181.n5 153.043
R395 a_13268_181.n6 a_13268_181.n3 110.158
R396 a_13268_181.n5 a_13268_181.n4 105.194
R397 a_13268_181.n15 a_13268_181.n14 98.501
R398 a_13268_181.n15 a_13268_181.n10 96.417
R399 a_13268_181.n16 a_13268_181.n15 78.403
R400 a_13268_181.n3 a_13268_181.n2 75.271
R401 a_13268_181.n19 a_13268_181.n0 55.263
R402 a_13268_181.n10 a_13268_181.n9 30
R403 a_13268_181.n14 a_13268_181.n13 30
R404 a_13268_181.n18 a_13268_181.n17 30
R405 a_13268_181.n19 a_13268_181.n18 25.263
R406 a_13268_181.n8 a_13268_181.n7 24.383
R407 a_13268_181.n12 a_13268_181.n11 24.383
R408 a_13268_181.n10 a_13268_181.n8 23.684
R409 a_13268_181.n14 a_13268_181.n12 23.684
R410 a_13268_181.n18 a_13268_181.n16 20.417
R411 a_13268_181.n1 a_13268_181.t4 14.282
R412 a_13268_181.n1 a_13268_181.t3 14.282
R413 a_13268_181.n2 a_13268_181.t0 14.282
R414 a_13268_181.n2 a_13268_181.t5 14.282
R415 a_13268_181.n3 a_13268_181.n1 12.119
R416 a_15059_182.n2 a_15059_182.n0 362.371
R417 a_15059_182.n2 a_15059_182.n1 15.218
R418 a_15059_182.n0 a_15059_182.t0 14.282
R419 a_15059_182.n0 a_15059_182.t2 14.282
R420 a_15059_182.n3 a_15059_182.n2 12.014
R421 a_11761_1004.n4 a_11761_1004.t7 480.392
R422 a_11761_1004.n4 a_11761_1004.t5 403.272
R423 a_11761_1004.n5 a_11761_1004.t6 346.633
R424 a_11761_1004.n8 a_11761_1004.n6 273.745
R425 a_11761_1004.n6 a_11761_1004.n5 153.315
R426 a_11761_1004.n6 a_11761_1004.n3 82.888
R427 a_11761_1004.n3 a_11761_1004.n2 76.002
R428 a_11761_1004.n8 a_11761_1004.n7 30
R429 a_11761_1004.n5 a_11761_1004.n4 28.835
R430 a_11761_1004.n9 a_11761_1004.n0 24.383
R431 a_11761_1004.n9 a_11761_1004.n8 23.684
R432 a_11761_1004.n1 a_11761_1004.t4 14.282
R433 a_11761_1004.n1 a_11761_1004.t3 14.282
R434 a_11761_1004.n2 a_11761_1004.t0 14.282
R435 a_11761_1004.n2 a_11761_1004.t1 14.282
R436 a_11761_1004.n3 a_11761_1004.n1 12.85
R437 a_9183_943.n4 a_9183_943.t7 480.392
R438 a_9183_943.n6 a_9183_943.t8 454.685
R439 a_9183_943.n6 a_9183_943.t10 428.979
R440 a_9183_943.n4 a_9183_943.t9 403.272
R441 a_9183_943.n5 a_9183_943.t5 266.974
R442 a_9183_943.n7 a_9183_943.t6 221.453
R443 a_9183_943.n11 a_9183_943.n9 194.086
R444 a_9183_943.n9 a_9183_943.n3 162.547
R445 a_9183_943.n7 a_9183_943.n6 108.494
R446 a_9183_943.n5 a_9183_943.n4 108.494
R447 a_9183_943.n8 a_9183_943.n7 78.947
R448 a_9183_943.n8 a_9183_943.n5 77.315
R449 a_9183_943.n3 a_9183_943.n2 76.002
R450 a_9183_943.n9 a_9183_943.n8 76
R451 a_9183_943.n11 a_9183_943.n10 30
R452 a_9183_943.n12 a_9183_943.n0 24.383
R453 a_9183_943.n12 a_9183_943.n11 23.684
R454 a_9183_943.n1 a_9183_943.t3 14.282
R455 a_9183_943.n1 a_9183_943.t2 14.282
R456 a_9183_943.n2 a_9183_943.t0 14.282
R457 a_9183_943.n2 a_9183_943.t1 14.282
R458 a_9183_943.n3 a_9183_943.n1 12.85
R459 a_91_75.n4 a_91_75.n3 19.724
R460 a_91_75.t0 a_91_75.n5 11.595
R461 a_91_75.t0 a_91_75.n4 9.207
R462 a_91_75.n2 a_91_75.n0 8.543
R463 a_91_75.t0 a_91_75.n2 3.034
R464 a_91_75.n2 a_91_75.n1 0.443
R465 a_372_182.n8 a_372_182.n6 96.467
R466 a_372_182.n3 a_372_182.n1 44.628
R467 a_372_182.t0 a_372_182.n8 32.417
R468 a_372_182.n3 a_372_182.n2 23.284
R469 a_372_182.n6 a_372_182.n5 22.349
R470 a_372_182.t0 a_372_182.n10 20.241
R471 a_372_182.n10 a_372_182.n9 13.494
R472 a_372_182.n6 a_372_182.n4 8.443
R473 a_372_182.t0 a_372_182.n0 8.137
R474 a_372_182.t0 a_372_182.n3 5.727
R475 a_372_182.n8 a_372_182.n7 1.435
R476 a_13654_73.n2 a_13654_73.n0 34.602
R477 a_13654_73.n2 a_13654_73.n1 2.138
R478 a_13654_73.t0 a_13654_73.n2 0.069
R479 a_12988_73.n1 a_12988_73.n0 32.249
R480 a_12988_73.t0 a_12988_73.n5 7.911
R481 a_12988_73.n4 a_12988_73.n2 4.032
R482 a_12988_73.n4 a_12988_73.n3 3.644
R483 a_12988_73.t0 a_12988_73.n1 2.534
R484 a_12988_73.t0 a_12988_73.n4 1.099
R485 a_7469_1004.n4 a_7469_1004.t5 480.392
R486 a_7469_1004.n4 a_7469_1004.t6 403.272
R487 a_7469_1004.n5 a_7469_1004.t7 293.527
R488 a_7469_1004.n8 a_7469_1004.n6 220.639
R489 a_7469_1004.n6 a_7469_1004.n5 153.315
R490 a_7469_1004.n6 a_7469_1004.n3 135.994
R491 a_7469_1004.n5 a_7469_1004.n4 81.941
R492 a_7469_1004.n3 a_7469_1004.n2 76.002
R493 a_7469_1004.n8 a_7469_1004.n7 30
R494 a_7469_1004.n9 a_7469_1004.n0 24.383
R495 a_7469_1004.n9 a_7469_1004.n8 23.684
R496 a_7469_1004.n1 a_7469_1004.t4 14.282
R497 a_7469_1004.n1 a_7469_1004.t3 14.282
R498 a_7469_1004.n2 a_7469_1004.t1 14.282
R499 a_7469_1004.n2 a_7469_1004.t0 14.282
R500 a_7469_1004.n3 a_7469_1004.n1 12.85
R501 a_2406_73.n12 a_2406_73.n11 26.811
R502 a_2406_73.n6 a_2406_73.n5 24.977
R503 a_2406_73.n2 a_2406_73.n1 24.877
R504 a_2406_73.t0 a_2406_73.n2 12.677
R505 a_2406_73.t0 a_2406_73.n3 11.595
R506 a_2406_73.t1 a_2406_73.n8 8.137
R507 a_2406_73.t0 a_2406_73.n4 7.273
R508 a_2406_73.t0 a_2406_73.n0 6.109
R509 a_2406_73.t1 a_2406_73.n7 4.864
R510 a_2406_73.t0 a_2406_73.n12 2.074
R511 a_2406_73.n7 a_2406_73.n6 1.13
R512 a_2406_73.n12 a_2406_73.t1 0.937
R513 a_2406_73.t1 a_2406_73.n10 0.804
R514 a_2406_73.n10 a_2406_73.n9 0.136
R515 a_4664_182.n8 a_4664_182.n6 96.467
R516 a_4664_182.n3 a_4664_182.n1 44.628
R517 a_4664_182.t0 a_4664_182.n8 32.417
R518 a_4664_182.n3 a_4664_182.n2 23.284
R519 a_4664_182.n6 a_4664_182.n5 22.349
R520 a_4664_182.t0 a_4664_182.n10 20.241
R521 a_4664_182.n10 a_4664_182.n9 13.494
R522 a_4664_182.n6 a_4664_182.n4 8.443
R523 a_4664_182.t0 a_4664_182.n0 8.137
R524 a_4664_182.t0 a_4664_182.n3 5.727
R525 a_4664_182.n8 a_4664_182.n7 1.435
R526 a_9658_73.n12 a_9658_73.n11 26.811
R527 a_9658_73.n6 a_9658_73.n5 24.977
R528 a_9658_73.n2 a_9658_73.n1 24.877
R529 a_9658_73.t0 a_9658_73.n2 12.677
R530 a_9658_73.t0 a_9658_73.n3 11.595
R531 a_9658_73.t1 a_9658_73.n8 8.137
R532 a_9658_73.t0 a_9658_73.n4 7.273
R533 a_9658_73.t0 a_9658_73.n0 6.109
R534 a_9658_73.t1 a_9658_73.n7 4.864
R535 a_9658_73.t0 a_9658_73.n12 2.074
R536 a_9658_73.n7 a_9658_73.n6 1.13
R537 a_9658_73.n12 a_9658_73.t1 0.937
R538 a_9658_73.t1 a_9658_73.n10 0.804
R539 a_9658_73.n10 a_9658_73.n9 0.136
R540 a_3303_383.n5 a_3303_383.t6 512.525
R541 a_3303_383.n4 a_3303_383.t10 512.525
R542 a_3303_383.n9 a_3303_383.t12 472.359
R543 a_3303_383.n9 a_3303_383.t5 384.527
R544 a_3303_383.n5 a_3303_383.t11 371.139
R545 a_3303_383.n4 a_3303_383.t7 371.139
R546 a_3303_383.n6 a_3303_383.n5 258.98
R547 a_3303_383.n10 a_3303_383.t13 198.113
R548 a_3303_383.n8 a_3303_383.n4 195.827
R549 a_3303_383.n12 a_3303_383.n3 189.099
R550 a_3303_383.n6 a_3303_383.t9 176.995
R551 a_3303_383.n7 a_3303_383.t8 170.569
R552 a_3303_383.n14 a_3303_383.n12 167.533
R553 a_3303_383.n7 a_3303_383.n6 153.043
R554 a_3303_383.n10 a_3303_383.n9 146.66
R555 a_3303_383.n11 a_3303_383.n8 112.41
R556 a_3303_383.n11 a_3303_383.n10 78.947
R557 a_3303_383.n3 a_3303_383.n2 76.002
R558 a_3303_383.n12 a_3303_383.n11 76
R559 a_3303_383.n8 a_3303_383.n7 63.152
R560 a_3303_383.n14 a_3303_383.n13 30
R561 a_3303_383.n15 a_3303_383.n0 24.383
R562 a_3303_383.n15 a_3303_383.n14 23.684
R563 a_3303_383.n1 a_3303_383.t4 14.282
R564 a_3303_383.n1 a_3303_383.t3 14.282
R565 a_3303_383.n2 a_3303_383.t0 14.282
R566 a_3303_383.n2 a_3303_383.t1 14.282
R567 a_3303_383.n3 a_3303_383.n1 12.85
R568 a_7364_73.n12 a_7364_73.n11 26.811
R569 a_7364_73.n6 a_7364_73.n5 24.977
R570 a_7364_73.n2 a_7364_73.n1 24.877
R571 a_7364_73.t0 a_7364_73.n2 12.677
R572 a_7364_73.t0 a_7364_73.n3 11.595
R573 a_7364_73.t1 a_7364_73.n8 8.137
R574 a_7364_73.t0 a_7364_73.n4 7.273
R575 a_7364_73.t0 a_7364_73.n0 6.109
R576 a_7364_73.t1 a_7364_73.n7 4.864
R577 a_7364_73.t0 a_7364_73.n12 2.074
R578 a_7364_73.n7 a_7364_73.n6 1.13
R579 a_7364_73.n12 a_7364_73.t1 0.937
R580 a_7364_73.t1 a_7364_73.n10 0.804
R581 a_7364_73.n10 a_7364_73.n9 0.136
R582 a_3738_73.n12 a_3738_73.n11 26.811
R583 a_3738_73.n6 a_3738_73.n5 24.977
R584 a_3738_73.n2 a_3738_73.n1 24.877
R585 a_3738_73.t0 a_3738_73.n2 12.677
R586 a_3738_73.t0 a_3738_73.n3 11.595
R587 a_3738_73.t1 a_3738_73.n8 8.137
R588 a_3738_73.t0 a_3738_73.n4 7.273
R589 a_3738_73.t0 a_3738_73.n0 6.109
R590 a_3738_73.t1 a_3738_73.n7 4.864
R591 a_3738_73.t0 a_3738_73.n12 2.074
R592 a_3738_73.n7 a_3738_73.n6 1.13
R593 a_3738_73.n12 a_3738_73.t1 0.937
R594 a_3738_73.t1 a_3738_73.n10 0.804
R595 a_3738_73.n10 a_3738_73.n9 0.136
R596 a_10324_73.t0 a_10324_73.n1 34.62
R597 a_10324_73.t0 a_10324_73.n0 8.137
R598 a_10324_73.t0 a_10324_73.n2 4.69
R599 a_8956_182.n10 a_8956_182.n8 82.852
R600 a_8956_182.n7 a_8956_182.n6 32.833
R601 a_8956_182.n8 a_8956_182.t1 32.416
R602 a_8956_182.n10 a_8956_182.n9 27.2
R603 a_8956_182.n11 a_8956_182.n0 23.498
R604 a_8956_182.n3 a_8956_182.n2 23.284
R605 a_8956_182.n11 a_8956_182.n10 22.4
R606 a_8956_182.n7 a_8956_182.n4 19.017
R607 a_8956_182.n6 a_8956_182.n5 13.494
R608 a_8956_182.t1 a_8956_182.n1 7.04
R609 a_8956_182.t1 a_8956_182.n3 5.727
R610 a_8956_182.n8 a_8956_182.n7 1.435
R611 a_11656_73.n12 a_11656_73.n11 26.811
R612 a_11656_73.n6 a_11656_73.n5 24.977
R613 a_11656_73.n2 a_11656_73.n1 24.877
R614 a_11656_73.t0 a_11656_73.n2 12.677
R615 a_11656_73.t0 a_11656_73.n3 11.595
R616 a_11656_73.t1 a_11656_73.n8 8.137
R617 a_11656_73.t0 a_11656_73.n4 7.273
R618 a_11656_73.t0 a_11656_73.n0 6.109
R619 a_11656_73.t1 a_11656_73.n7 4.864
R620 a_11656_73.t0 a_11656_73.n12 2.074
R621 a_11656_73.n7 a_11656_73.n6 1.13
R622 a_11656_73.n12 a_11656_73.t1 0.937
R623 a_11656_73.t1 a_11656_73.n10 0.804
R624 a_11656_73.n10 a_11656_73.n9 0.136
R625 a_1074_73.n12 a_1074_73.n11 26.811
R626 a_1074_73.n6 a_1074_73.n5 24.977
R627 a_1074_73.n2 a_1074_73.n1 24.877
R628 a_1074_73.t0 a_1074_73.n2 12.677
R629 a_1074_73.t0 a_1074_73.n3 11.595
R630 a_1074_73.t1 a_1074_73.n8 8.137
R631 a_1074_73.t0 a_1074_73.n4 7.273
R632 a_1074_73.t0 a_1074_73.n0 6.109
R633 a_1074_73.t1 a_1074_73.n7 4.864
R634 a_1074_73.t0 a_1074_73.n12 2.074
R635 a_1074_73.n7 a_1074_73.n6 1.13
R636 a_1074_73.n12 a_1074_73.t1 0.937
R637 a_1074_73.t1 a_1074_73.n10 0.804
R638 a_1074_73.n10 a_1074_73.n9 0.136
R639 a_12322_73.n12 a_12322_73.n11 26.811
R640 a_12322_73.n6 a_12322_73.n5 24.977
R641 a_12322_73.n2 a_12322_73.n1 24.877
R642 a_12322_73.t0 a_12322_73.n2 12.677
R643 a_12322_73.t0 a_12322_73.n3 11.595
R644 a_12322_73.t1 a_12322_73.n8 8.137
R645 a_12322_73.t0 a_12322_73.n4 7.273
R646 a_12322_73.t0 a_12322_73.n0 6.109
R647 a_12322_73.t1 a_12322_73.n7 4.864
R648 a_12322_73.t0 a_12322_73.n12 2.074
R649 a_12322_73.n7 a_12322_73.n6 1.13
R650 a_12322_73.n12 a_12322_73.t1 0.937
R651 a_12322_73.t1 a_12322_73.n10 0.804
R652 a_12322_73.n10 a_12322_73.n9 0.136
R653 a_6698_73.n12 a_6698_73.n11 26.811
R654 a_6698_73.n6 a_6698_73.n5 24.977
R655 a_6698_73.n2 a_6698_73.n1 24.877
R656 a_6698_73.t0 a_6698_73.n2 12.677
R657 a_6698_73.t0 a_6698_73.n3 11.595
R658 a_6698_73.t1 a_6698_73.n8 8.137
R659 a_6698_73.t0 a_6698_73.n4 7.273
R660 a_6698_73.t0 a_6698_73.n0 6.109
R661 a_6698_73.t1 a_6698_73.n7 4.864
R662 a_6698_73.t0 a_6698_73.n12 2.074
R663 a_6698_73.n7 a_6698_73.n6 1.13
R664 a_6698_73.n12 a_6698_73.t1 0.937
R665 a_6698_73.t1 a_6698_73.n10 0.804
R666 a_6698_73.n10 a_6698_73.n9 0.136
R667 a_3072_73.n12 a_3072_73.n11 26.811
R668 a_3072_73.n6 a_3072_73.n5 24.977
R669 a_3072_73.n2 a_3072_73.n1 24.877
R670 a_3072_73.t0 a_3072_73.n2 12.677
R671 a_3072_73.t0 a_3072_73.n3 11.595
R672 a_3072_73.t1 a_3072_73.n8 8.137
R673 a_3072_73.t0 a_3072_73.n4 7.273
R674 a_3072_73.t0 a_3072_73.n0 6.109
R675 a_3072_73.t1 a_3072_73.n7 4.864
R676 a_3072_73.t0 a_3072_73.n12 2.074
R677 a_3072_73.n7 a_3072_73.n6 1.13
R678 a_3072_73.n12 a_3072_73.t1 0.937
R679 a_3072_73.t1 a_3072_73.n10 0.804
R680 a_3072_73.n10 a_3072_73.n9 0.136
R681 a_6032_73.t0 a_6032_73.n1 34.62
R682 a_6032_73.t0 a_6032_73.n0 8.137
R683 a_6032_73.t0 a_6032_73.n2 4.69
R684 a_14320_73.t0 a_14320_73.n1 34.62
R685 a_14320_73.t0 a_14320_73.n0 8.137
R686 a_14320_73.t0 a_14320_73.n2 4.69
R687 a_8675_75.n5 a_8675_75.n4 19.724
R688 a_8675_75.t0 a_8675_75.n3 11.595
R689 a_8675_75.t0 a_8675_75.n5 9.207
R690 a_8675_75.n2 a_8675_75.n1 2.455
R691 a_8675_75.n2 a_8675_75.n0 1.32
R692 a_8675_75.t0 a_8675_75.n2 0.246











































































































































































































































































































































































































































































































































.ends
