magic
tech sky130A
magscale 1 2
timestamp 1652468990
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 2055 945 2089 979
rect 5755 945 5789 979
rect 131 871 165 905
rect 649 871 683 905
rect 1315 871 1349 905
rect 2055 871 2089 905
rect 3165 871 3199 905
rect 3535 871 3569 905
rect 4275 871 4309 905
rect 4645 871 4679 905
rect 5755 871 5789 905
rect 5903 871 5937 905
rect 7605 871 7639 905
rect 131 797 165 831
rect 649 797 683 831
rect 2055 797 2089 831
rect 4275 797 4309 831
rect 4645 797 4679 831
rect 5755 797 5789 831
rect 5903 797 5937 831
rect 7605 797 7639 831
rect 131 723 165 757
rect 649 723 683 757
rect 3165 723 3199 757
rect 3831 723 3865 757
rect 4275 723 4309 757
rect 4645 723 4679 757
rect 5755 723 5789 757
rect 5903 723 5937 757
rect 7605 723 7639 757
rect 131 649 165 683
rect 649 649 683 683
rect 2055 649 2089 683
rect 3165 649 3199 683
rect 4275 649 4309 683
rect 4645 649 4679 683
rect 5755 649 5789 683
rect 5903 649 5937 683
rect 7605 649 7639 683
rect 131 575 165 609
rect 649 575 683 609
rect 871 575 905 609
rect 2055 575 2089 609
rect 3091 575 3125 609
rect 4275 575 4309 609
rect 4645 575 4679 609
rect 7605 575 7639 609
rect 131 501 165 535
rect 2055 501 2089 535
rect 3831 501 3865 535
rect 4275 501 4309 535
rect 4645 501 4679 535
rect 5755 501 5789 535
rect 5903 501 5937 535
rect 7605 501 7639 535
rect 649 427 683 461
rect 871 427 905 461
rect 5903 427 5937 461
rect 7605 427 7639 461
<< metal1 >>
rect -34 1446 7804 1514
rect 2125 945 5755 979
rect 4321 871 4609 905
rect 1657 723 2349 757
rect 6565 649 6977 683
rect 5455 575 6829 609
rect 2421 427 4757 461
rect 649 387 683 391
rect 5903 387 5937 391
rect 649 353 5937 387
rect -34 -34 7804 34
use li1_M1_contact  li1_M1_contact_3 pcells
timestamp 1648061256
transform 0 -1 666 1 0 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 2072 0 -1 962
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform 1 0 2368 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform -1 0 2368 0 -1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform 1 0 4662 0 1 888
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 0 1 5772 -1 0 926
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 4810 0 1 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 5402 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform 0 -1 5920 1 0 444
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform -1 0 6512 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform 1 0 6882 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 7030 0 1 666
box -53 -33 29 33
use xor2X1_pcell  xor2X1_pcell_0 pcells
timestamp 1652468990
transform 1 0 0 0 1 0
box -87 -34 2307 1550
use xor2X1_pcell  xor2X1_pcell_1
timestamp 1652468990
transform 1 0 2220 0 1 0
box -87 -34 2307 1550
use and2x1_pcell  and2x1_pcell_0 pcells
timestamp 1652468990
transform 1 0 4440 0 1 0
box -87 -34 1197 1550
use and2x1_pcell  and2x1_pcell_1
timestamp 1652468990
transform 1 0 5550 0 1 0
box -87 -34 1197 1550
use or2x1_pcell  or2x1_pcell_0 pcells
timestamp 1652468990
transform 1 0 6660 0 1 0
box -87 -34 1197 1550
<< labels >>
rlabel locali 3831 723 3865 757 1 SUM
port 1 nsew signal output
rlabel locali 3831 501 3865 535 1 SUM
port 1 nsew signal output
rlabel locali 3165 723 3199 757 1 SUM
port 1 nsew signal output
rlabel locali 3165 649 3199 683 1 SUM
port 1 nsew signal output
rlabel locali 3165 871 3199 905 1 SUM
port 1 nsew signal output
rlabel locali 7605 649 7639 683 1 COUT
port 2 nsew signal output
rlabel locali 7605 723 7639 757 1 COUT
port 2 nsew signal output
rlabel locali 7605 797 7639 831 1 COUT
port 2 nsew signal output
rlabel locali 7605 871 7639 905 1 COUT
port 2 nsew signal output
rlabel locali 7605 575 7639 609 1 COUT
port 2 nsew signal output
rlabel locali 7605 501 7639 535 1 COUT
port 2 nsew signal output
rlabel locali 7605 427 7639 461 1 COUT
port 2 nsew signal output
rlabel locali 131 871 165 905 1 A
port 3 nsew signal input
rlabel locali 131 723 165 757 1 A
port 3 nsew signal input
rlabel locali 131 649 165 683 1 A
port 3 nsew signal input
rlabel locali 131 575 165 609 1 A
port 3 nsew signal input
rlabel locali 131 501 165 535 1 A
port 3 nsew signal input
rlabel locali 649 871 683 905 1 A
port 3 nsew signal input
rlabel locali 649 797 683 831 1 A
port 3 nsew signal input
rlabel locali 649 723 683 757 1 A
port 3 nsew signal input
rlabel locali 649 649 683 683 1 A
port 3 nsew signal input
rlabel locali 649 575 683 609 1 A
port 3 nsew signal input
rlabel locali 649 427 683 461 1 A
port 3 nsew signal input
rlabel locali 5903 871 5937 905 1 A
port 3 nsew signal input
rlabel locali 5903 797 5937 831 1 A
port 3 nsew signal input
rlabel locali 5903 723 5937 757 1 A
port 3 nsew signal input
rlabel locali 5903 649 5937 683 1 A
port 3 nsew signal input
rlabel locali 5903 501 5937 535 1 A
port 3 nsew signal input
rlabel locali 5903 427 5937 461 1 A
port 3 nsew signal input
rlabel locali 131 797 165 831 1 A
port 3 nsew signal input
rlabel locali 1315 871 1349 905 1 B
port 4 nsew signal input
rlabel locali 2055 871 2089 905 1 B
port 4 nsew signal input
rlabel locali 2055 945 2089 979 1 B
port 4 nsew signal input
rlabel locali 2055 797 2089 831 1 B
port 4 nsew signal input
rlabel locali 2055 649 2089 683 1 B
port 4 nsew signal input
rlabel locali 2055 501 2089 535 1 B
port 4 nsew signal input
rlabel locali 2055 575 2089 609 1 B
port 4 nsew signal input
rlabel locali 871 575 905 609 1 B
port 4 nsew signal input
rlabel locali 871 427 905 461 1 B
port 4 nsew signal input
rlabel locali 5755 649 5789 683 1 B
port 4 nsew signal input
rlabel locali 5755 723 5789 757 1 B
port 4 nsew signal input
rlabel locali 5755 797 5789 831 1 B
port 4 nsew signal input
rlabel locali 5755 871 5789 905 1 B
port 4 nsew signal input
rlabel locali 5755 945 5789 979 1 B
port 4 nsew signal input
rlabel locali 5755 501 5789 535 1 B
port 4 nsew signal input
rlabel locali 4645 871 4679 905 1 CIN
port 5 nsew signal input
rlabel locali 4645 797 4679 831 1 CIN
port 5 nsew signal input
rlabel locali 4645 723 4679 757 1 CIN
port 5 nsew signal input
rlabel locali 4645 649 4679 683 1 CIN
port 5 nsew signal input
rlabel locali 4645 575 4679 609 1 CIN
port 5 nsew signal input
rlabel locali 4645 501 4679 535 1 CIN
port 5 nsew signal input
rlabel locali 4275 871 4309 905 1 CIN
port 5 nsew signal input
rlabel locali 4275 575 4309 609 1 CIN
port 5 nsew signal input
rlabel locali 4275 649 4309 683 1 CIN
port 5 nsew signal input
rlabel locali 4275 723 4309 757 1 CIN
port 5 nsew signal input
rlabel locali 4275 797 4309 831 1 CIN
port 5 nsew signal input
rlabel locali 4275 501 4309 535 1 CIN
port 5 nsew signal input
rlabel locali 3535 871 3569 905 1 CIN
port 5 nsew signal input
rlabel locali 3091 575 3125 609 1 CIN
port 5 nsew signal input
rlabel metal1 -34 1446 7804 1514 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 -34 -34 7804 34 1 VGND
port 7 nsew ground bidirectional abutment
rlabel nwell 57 1463 91 1497 1 VPB
port 8 nsew power bidirectional
rlabel pwell 57 -17 91 17 1 VNB
port 9 nsew ground bidirectional
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
