* SPICE3 file created from DLATCHN.ext - technology: sky130A

.subckt DLATCHN Q D GATE_N VDD GND
X0 m1_793_723# D invx1_pcell_0/pmos2_0/VSUBS invx1_pcell_0/pmos2_0/VSUBS nshort w=3 l=0.15
X1 VDD D m1_793_723# VDD pshort w=2 l=0.15
X2 m1_349_575# GATE_N GND GND nshort w=3 l=0.15
X3 VDD GATE_N m1_349_575# VDD pshort w=2 l=0.15
X4 m1_1903_723# and2x1_pcell_0/m1_547_649# GND GND nshort w=3 l=0.15
X5 VDD and2x1_pcell_0/m1_547_649# m1_1903_723# VDD pshort w=2 l=0.15
X6 GND m1_793_723# and2x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X7 and2x1_pcell_0/m1_547_649# m1_349_575# and2x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X8 VDD m1_793_723# and2x1_pcell_0/m1_547_649# VDD pshort w=2 l=0.15
X9 VDD m1_349_575# and2x1_pcell_0/m1_547_649# VDD pshort w=2 l=0.15
X10 m1_3013_797# and2x1_pcell_1/m1_547_649# and2x1_pcell_1/VSUBS and2x1_pcell_1/VSUBS nshort w=3 l=0.15
X11 VDD and2x1_pcell_1/m1_547_649# m1_3013_797# VDD pshort w=2 l=0.15
X12 and2x1_pcell_1/VSUBS m1_349_575# and2x1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# and2x1_pcell_1/VSUBS nshort w=3 l=0.15
X13 and2x1_pcell_1/m1_547_649# D and2x1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# and2x1_pcell_1/VSUBS nshort w=3 l=0.15
X14 VDD m1_349_575# and2x1_pcell_1/m1_547_649# VDD pshort w=2 l=0.15
X15 VDD D and2x1_pcell_1/m1_547_649# VDD pshort w=2 l=0.15
X16 VDD m1_1903_723# nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X17 Q m1_3531_723# nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X18 Q m1_1903_723# nor2x1_pcell_0/pmos2_1_1/VSUBS nor2x1_pcell_0/pmos2_1_1/VSUBS nshort w=3 l=0.15
X19 Q m1_3531_723# nor2x1_pcell_0/pmos2_1_1/VSUBS nor2x1_pcell_0/pmos2_1_1/VSUBS nshort w=3 l=0.15
X20 VDD Q nor2x1_pcell_1/a_317_1331# VDD pshort w=2 l=0.15
X21 m1_3531_723# m1_3013_797# nor2x1_pcell_1/a_317_1331# VDD pshort w=2 l=0.15
X22 m1_3531_723# Q li1_M1_contact_12/VSUBS li1_M1_contact_12/VSUBS nshort w=3 l=0.15
X23 m1_3531_723# m1_3013_797# li1_M1_contact_12/VSUBS li1_M1_contact_12/VSUBS nshort w=3 l=0.15
.ends
