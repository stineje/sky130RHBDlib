magic
tech sky130A
magscale 1 2
timestamp 1652394001
<< nwell >>
rect 55 1463 89 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 131 871 165 905
rect 871 871 905 905
rect 1167 871 1201 905
rect 1463 871 1497 905
rect 1685 871 1719 905
rect 2277 872 2311 906
rect 131 797 165 831
rect 353 797 387 831
rect 1685 797 1719 831
rect 2277 798 2311 832
rect 131 723 165 757
rect 353 723 387 757
rect 871 723 905 757
rect 1167 723 1201 757
rect 1463 723 1497 757
rect 1685 723 1719 757
rect 2277 724 2311 758
rect 131 649 165 683
rect 353 649 387 683
rect 871 649 905 683
rect 1167 649 1201 683
rect 1463 649 1497 683
rect 1685 649 1719 683
rect 2277 650 2311 684
rect 131 575 165 609
rect 353 575 387 609
rect 871 575 905 609
rect 1167 575 1201 609
rect 1463 575 1497 609
rect 1685 575 1719 609
rect 2277 576 2311 610
rect 131 501 165 535
rect 353 501 387 535
rect 871 501 905 535
rect 1167 501 1201 535
rect 1463 501 1497 535
rect 1685 501 1719 535
rect 2277 502 2311 536
rect 2277 428 2311 462
<< metal1 >>
rect -34 1446 2476 1514
rect -34 -34 2476 34
use voter3x1_pcell  voter3x1_pcell_0 pcells
timestamp 1652393968
transform 1 0 0 0 1 0
box -87 -34 2529 1550
<< labels >>
rlabel locali 2277 798 2311 832 1 Y
port 1 nsew signal output
rlabel locali 2277 724 2311 758 1 Y
port 1 nsew signal output
rlabel locali 2277 872 2311 906 1 Y
port 1 nsew signal output
rlabel locali 2277 650 2311 684 1 Y
port 1 nsew signal output
rlabel locali 2277 576 2311 610 1 Y
port 1 nsew signal output
rlabel locali 2277 502 2311 536 1 Y
port 1 nsew signal output
rlabel locali 2277 428 2311 462 1 Y
port 1 nsew signal output
rlabel locali 1685 871 1719 905 1 A
port 2 nsew signal input
rlabel locali 353 797 387 831 1 A
port 2 nsew signal input
rlabel locali 353 723 387 757 1 A
port 2 nsew signal input
rlabel locali 353 649 387 683 1 A
port 2 nsew signal input
rlabel locali 353 575 387 609 1 A
port 2 nsew signal input
rlabel locali 353 501 387 535 1 A
port 2 nsew signal input
rlabel locali 1685 501 1719 535 1 A
port 2 nsew signal input
rlabel locali 1685 575 1719 609 1 A
port 2 nsew signal input
rlabel locali 1685 649 1719 683 1 A
port 2 nsew signal input
rlabel locali 1685 723 1719 757 1 A
port 2 nsew signal input
rlabel locali 1685 797 1719 831 1 A
port 2 nsew signal input
rlabel locali 131 871 165 905 1 B
port 3 nsew signal input
rlabel locali 131 797 165 831 1 B
port 3 nsew signal input
rlabel locali 131 723 165 757 1 B
port 3 nsew signal input
rlabel locali 131 649 165 683 1 B
port 3 nsew signal input
rlabel locali 131 575 165 609 1 B
port 3 nsew signal input
rlabel locali 131 501 165 535 1 B
port 3 nsew signal input
rlabel locali 871 501 905 535 1 B
port 3 nsew signal input
rlabel locali 871 575 905 609 1 B
port 3 nsew signal input
rlabel locali 871 649 905 683 1 B
port 3 nsew signal input
rlabel locali 871 723 905 757 1 B
port 3 nsew signal input
rlabel locali 871 871 905 905 1 B
port 3 nsew signal input
rlabel locali 1167 501 1201 535 1 C
port 4 nsew signal input
rlabel locali 1167 575 1201 609 1 C
port 4 nsew signal input
rlabel locali 1167 649 1201 683 1 C
port 4 nsew signal input
rlabel locali 1167 723 1201 757 1 C
port 4 nsew signal input
rlabel locali 1167 871 1201 905 1 C
port 4 nsew signal input
rlabel locali 1463 501 1497 535 1 C
port 4 nsew signal input
rlabel locali 1463 575 1497 609 1 C
port 4 nsew signal input
rlabel locali 1463 649 1497 683 1 C
port 4 nsew signal input
rlabel locali 1463 723 1497 757 1 C
port 4 nsew signal input
rlabel locali 1463 871 1497 905 1 C
port 4 nsew signal input
rlabel metal1 -34 1446 2476 1514 1 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 -34 -34 2476 34 1 VGND
port 6 nsew ground bidirectional abutment
rlabel nwell 55 1463 89 1497 1 VPB
rlabel pwell 57 -17 91 17 1 VNB
<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 2442 1480
string LEFsymmetry X Y R90
<< end >>
