* SPICE3 file created from AO3X1.ext - technology: sky130A

.subckt AO3X1 Y A B C VDD GND
X0 a_864_181 a_217_1004 GND GND nshort w=3 l=0.15
X1 VDD B a_217_1004 VDD pshort w=2 l=0.15 M=2
X2 GND A a_112_73 GND nshort w=3 l=0.15
X3 Y a_864_181 VDD VDD pshort w=2 l=0.15 M=2
X4 a_797_1005 C a_864_181 VDD pshort w=2 l=0.15 M=2
X5 a_217_1004 A VDD VDD pshort w=2 l=0.15 M=2
X6 a_217_1004 B a_112_73 GND nshort w=3 l=0.15
X7 a_864_181 C GND GND nshort w=3 l=0.15
X8 a_797_1005 a_217_1004 VDD VDD pshort w=2 l=0.15 M=2
X9 Y a_864_181 GND GND nshort w=3 l=0.15
C0 VDD GND 4.59fF
.ends
