* SPICE3 file created from AND2X1.ext - technology: sky130A

.subckt AND2X1 Y A B VPB VNB
M1000 VNB a_168_157# a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=1.3199p pd=9.67u as=0p ps=0u
M1001 VPB.t1 a_168_157# a_217_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_851_182.t1 a_217_1004.t5 VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t3 a_343_383# a_217_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPB.t5 a_217_1004.t6 a_851_182.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_217_1004.t1 a_168_157# VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_217_1004.t3 a_343_383# VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 a_343_383# VPB 0.07fF
C1 a_343_383# a_168_157# 0.26fF
C2 VPB a_168_157# 0.08fF
R0 a_217_1004.n4 a_217_1004.t6 512.525
R1 a_217_1004.n4 a_217_1004.t5 371.139
R2 a_217_1004.n5 a_217_1004.t7 220.263
R3 a_217_1004.n8 a_217_1004.n6 194.086
R4 a_217_1004.n6 a_217_1004.n3 162.547
R5 a_217_1004.n5 a_217_1004.n4 158.3
R6 a_217_1004.n6 a_217_1004.n5 153.043
R7 a_217_1004.n3 a_217_1004.n2 76.002
R8 a_217_1004.n8 a_217_1004.n7 30
R9 a_217_1004.n9 a_217_1004.n0 24.383
R10 a_217_1004.n9 a_217_1004.n8 23.684
R11 a_217_1004.n1 a_217_1004.t4 14.282
R12 a_217_1004.n1 a_217_1004.t3 14.282
R13 a_217_1004.n2 a_217_1004.t0 14.282
R14 a_217_1004.n2 a_217_1004.t1 14.282
R15 a_217_1004.n3 a_217_1004.n1 12.85
R16 VPB VPB.n125 126.832
R17 VPB.n108 VPB.n106 94.117
R18 VPB.n110 VPB.n109 76
R19 VPB.n118 VPB.n117 76
R20 VPB.n75 VPB.n74 68.979
R21 VPB.n68 VPB.n67 64.528
R22 VPB.n27 VPB.n26 61.764
R23 VPB.n84 VPB.t0 55.106
R24 VPB.n78 VPB.t4 55.106
R25 VPB.n66 VPB.t5 55.106
R26 VPB.n102 VPB.t3 55.106
R27 VPB.n99 VPB.n98 48.952
R28 VPB.n86 VPB.n85 44.502
R29 VPB.n93 VPB.n83 40.824
R30 VPB.n122 VPB.n118 20.452
R31 VPB.n65 VPB.n62 20.452
R32 VPB.n95 VPB.n94 17.801
R33 VPB.n83 VPB.t2 14.282
R34 VPB.n83 VPB.t1 14.282
R35 VPB.n65 VPB.n64 13.653
R36 VPB.n64 VPB.n63 13.653
R37 VPB.n70 VPB.n69 13.653
R38 VPB.n69 VPB.n68 13.653
R39 VPB.n73 VPB.n72 13.653
R40 VPB.n72 VPB.n71 13.653
R41 VPB.n77 VPB.n76 13.653
R42 VPB.n76 VPB.n75 13.653
R43 VPB.n81 VPB.n80 13.653
R44 VPB.n80 VPB.n79 13.653
R45 VPB.n109 VPB.n108 13.653
R46 VPB.n108 VPB.n107 13.653
R47 VPB.n105 VPB.n104 13.653
R48 VPB.n104 VPB.n103 13.653
R49 VPB.n101 VPB.n100 13.653
R50 VPB.n100 VPB.n99 13.653
R51 VPB.n97 VPB.n96 13.653
R52 VPB.n96 VPB.n95 13.653
R53 VPB.n92 VPB.n91 13.653
R54 VPB.n91 VPB.n90 13.653
R55 VPB.n88 VPB.n87 13.653
R56 VPB.n87 VPB.n86 13.653
R57 VPB.n16 VPB.n15 13.653
R58 VPB.n15 VPB.n14 13.653
R59 VPB.n118 VPB.n0 13.653
R60 VPB VPB.n0 13.653
R61 VPB.n90 VPB.n89 13.35
R62 VPB.n122 VPB.n121 13.276
R63 VPB.n121 VPB.n119 13.276
R64 VPB.n41 VPB.n23 13.276
R65 VPB.n23 VPB.n21 13.276
R66 VPB.n73 VPB.n70 13.276
R67 VPB.n77 VPB.n73 13.276
R68 VPB.n82 VPB.n81 13.276
R69 VPB.n109 VPB.n82 13.276
R70 VPB.n109 VPB.n105 13.276
R71 VPB.n101 VPB.n97 13.276
R72 VPB.n92 VPB.n88 13.276
R73 VPB.n118 VPB.n16 13.276
R74 VPB.n62 VPB.n44 13.276
R75 VPB.n44 VPB.n42 13.276
R76 VPB.n49 VPB.n47 12.796
R77 VPB.n49 VPB.n48 12.564
R78 VPB.n55 VPB.n54 12.198
R79 VPB.n57 VPB.n56 12.198
R80 VPB.n55 VPB.n52 12.198
R81 VPB.n102 VPB.n101 11.841
R82 VPB.n88 VPB.n84 11.482
R83 VPB.n81 VPB.n78 10.944
R84 VPB.n66 VPB.n65 10.585
R85 VPB.n62 VPB.n61 7.5
R86 VPB.n47 VPB.n46 7.5
R87 VPB.n54 VPB.n53 7.5
R88 VPB.n52 VPB.n51 7.5
R89 VPB.n44 VPB.n43 7.5
R90 VPB.n59 VPB.n45 7.5
R91 VPB.n23 VPB.n22 7.5
R92 VPB.n36 VPB.n35 7.5
R93 VPB.n30 VPB.n29 7.5
R94 VPB.n32 VPB.n31 7.5
R95 VPB.n25 VPB.n24 7.5
R96 VPB.n41 VPB.n40 7.5
R97 VPB.n121 VPB.n120 7.5
R98 VPB.n12 VPB.n11 7.5
R99 VPB.n6 VPB.n5 7.5
R100 VPB.n8 VPB.n7 7.5
R101 VPB.n2 VPB.n1 7.5
R102 VPB.n123 VPB.n122 7.5
R103 VPB.n82 VPB.n41 7.176
R104 VPB.n93 VPB.n92 6.817
R105 VPB.n37 VPB.n34 6.729
R106 VPB.n33 VPB.n30 6.729
R107 VPB.n28 VPB.n25 6.729
R108 VPB.n13 VPB.n10 6.729
R109 VPB.n9 VPB.n6 6.729
R110 VPB.n4 VPB.n2 6.729
R111 VPB.n28 VPB.n27 6.728
R112 VPB.n33 VPB.n32 6.728
R113 VPB.n37 VPB.n36 6.728
R114 VPB.n40 VPB.n39 6.728
R115 VPB.n4 VPB.n3 6.728
R116 VPB.n9 VPB.n8 6.728
R117 VPB.n13 VPB.n12 6.728
R118 VPB.n124 VPB.n123 6.728
R119 VPB.n97 VPB.n93 6.458
R120 VPB.n61 VPB.n60 6.398
R121 VPB.n70 VPB.n66 2.691
R122 VPB.n78 VPB.n77 2.332
R123 VPB.n84 VPB.n16 1.794
R124 VPB.n105 VPB.n102 1.435
R125 VPB.n59 VPB.n50 1.402
R126 VPB.n59 VPB.n55 1.402
R127 VPB.n59 VPB.n57 1.402
R128 VPB.n59 VPB.n58 1.402
R129 VPB.n60 VPB.n59 0.735
R130 VPB.n59 VPB.n49 0.735
R131 VPB.n38 VPB.n37 0.387
R132 VPB.n38 VPB.n33 0.387
R133 VPB.n38 VPB.n28 0.387
R134 VPB.n39 VPB.n38 0.387
R135 VPB.n125 VPB.n13 0.387
R136 VPB.n125 VPB.n9 0.387
R137 VPB.n125 VPB.n4 0.387
R138 VPB.n125 VPB.n124 0.387
R139 VPB.n110 VPB.n20 0.272
R140 VPB.n117 VPB 0.198
R141 VPB.n18 VPB.n17 0.136
R142 VPB.n19 VPB.n18 0.136
R143 VPB.n20 VPB.n19 0.136
R144 VPB.n112 VPB.n111 0.136
R145 VPB.n113 VPB.n112 0.136
R146 VPB.n114 VPB.n113 0.136
R147 VPB.n115 VPB.n114 0.136
R148 VPB.n116 VPB.n115 0.136
R149 VPB.n117 VPB.n116 0.136
R150 VPB VPB.n110 0.068
R151 VPB.n111 VPB 0.068
R152 a_851_182.n3 a_851_182.n1 355.848
R153 a_851_182.n3 a_851_182.n2 30
R154 a_851_182.n4 a_851_182.n0 24.383
R155 a_851_182.n4 a_851_182.n3 23.684
R156 a_851_182.n1 a_851_182.t0 14.282
R157 a_851_182.n1 a_851_182.t1 14.282
R158 a_112_73.n10 a_112_73.n9 93.333
R159 a_112_73.n2 a_112_73.n1 41.622
R160 a_112_73.n13 a_112_73.n12 26.667
R161 a_112_73.n6 a_112_73.n5 24.977
R162 a_112_73.t0 a_112_73.n2 21.209
R163 a_112_73.t0 a_112_73.n3 11.595
R164 a_112_73.t1 a_112_73.n8 8.137
R165 a_112_73.t0 a_112_73.n0 6.109
R166 a_112_73.t1 a_112_73.n7 4.864
R167 a_112_73.t0 a_112_73.n4 3.871
R168 a_112_73.t0 a_112_73.n13 2.535
R169 a_112_73.n13 a_112_73.t1 1.145
R170 a_112_73.n7 a_112_73.n6 1.13
R171 a_112_73.t1 a_112_73.n11 0.804
R172 a_112_73.n11 a_112_73.n10 0.136
R173 VNB VNB.n114 300.778
R174 VNB.n21 VNB.n20 199.897
R175 VNB.n91 VNB.n89 154.509
R176 VNB.n76 VNB.n72 84.842
R177 VNB.n101 VNB.n100 76
R178 VNB.n93 VNB.n92 76
R179 VNB.n62 VNB.n61 49.896
R180 VNB.n74 VNB.n73 36.678
R181 VNB.n37 VNB.n36 35.01
R182 VNB.t1 VNB.n29 32.601
R183 VNB.n55 VNB.n52 20.452
R184 VNB.n102 VNB.n101 20.452
R185 VNB.n56 VNB.n37 20.094
R186 VNB.n60 VNB.n34 20.094
R187 VNB.n67 VNB.n32 20.094
R188 VNB.n37 VNB.n35 19.017
R189 VNB.n31 VNB.t1 17.353
R190 VNB.n59 VNB.n58 13.653
R191 VNB.n58 VNB.n57 13.653
R192 VNB.n63 VNB.n62 13.653
R193 VNB.n66 VNB.n65 13.653
R194 VNB.n65 VNB.n64 13.653
R195 VNB.n70 VNB.n69 13.653
R196 VNB.n69 VNB.n68 13.653
R197 VNB.n92 VNB.n91 13.653
R198 VNB.n91 VNB.n90 13.653
R199 VNB.n88 VNB.n87 13.653
R200 VNB.n87 VNB.n86 13.653
R201 VNB.n85 VNB.n84 13.653
R202 VNB.n84 VNB.n83 13.653
R203 VNB.n82 VNB.n81 13.653
R204 VNB.n81 VNB.n80 13.653
R205 VNB.n79 VNB.n78 13.653
R206 VNB.n78 VNB.n77 13.653
R207 VNB.n75 VNB.n74 13.653
R208 VNB.n6 VNB.n5 13.653
R209 VNB.n5 VNB.n4 13.653
R210 VNB.n101 VNB.n0 13.653
R211 VNB VNB.n0 13.653
R212 VNB.n55 VNB.n54 13.653
R213 VNB.n54 VNB.n53 13.653
R214 VNB.n109 VNB.n106 13.577
R215 VNB.n40 VNB.n38 13.276
R216 VNB.n52 VNB.n40 13.276
R217 VNB.n13 VNB.n11 13.276
R218 VNB.n26 VNB.n13 13.276
R219 VNB.n66 VNB.n63 13.276
R220 VNB.n71 VNB.n70 13.276
R221 VNB.n92 VNB.n71 13.276
R222 VNB.n92 VNB.n88 13.276
R223 VNB.n88 VNB.n85 13.276
R224 VNB.n85 VNB.n82 13.276
R225 VNB.n82 VNB.n79 13.276
R226 VNB.n75 VNB.n6 13.276
R227 VNB.n101 VNB.n6 13.276
R228 VNB.n3 VNB.n1 13.276
R229 VNB.n102 VNB.n3 13.276
R230 VNB.n60 VNB.n59 13.097
R231 VNB.n32 VNB.n31 12.837
R232 VNB.n79 VNB.n76 10.764
R233 VNB.n70 VNB.n67 9.329
R234 VNB.n56 VNB.n55 8.97
R235 VNB.n31 VNB.n30 7.566
R236 VNB.n111 VNB.n110 7.5
R237 VNB.n19 VNB.n18 7.5
R238 VNB.n15 VNB.n14 7.5
R239 VNB.n13 VNB.n12 7.5
R240 VNB.n26 VNB.n25 7.5
R241 VNB.n103 VNB.n102 7.5
R242 VNB.n3 VNB.n2 7.5
R243 VNB.n108 VNB.n107 7.5
R244 VNB.n46 VNB.n45 7.5
R245 VNB.n42 VNB.n41 7.5
R246 VNB.n40 VNB.n39 7.5
R247 VNB.n52 VNB.n51 7.5
R248 VNB.n71 VNB.n26 7.176
R249 VNB.n113 VNB.n111 7.011
R250 VNB.n22 VNB.n19 7.011
R251 VNB.n17 VNB.n15 7.011
R252 VNB.n48 VNB.n46 7.011
R253 VNB.n44 VNB.n42 7.011
R254 VNB.n25 VNB.n24 7.01
R255 VNB.n17 VNB.n16 7.01
R256 VNB.n22 VNB.n21 7.01
R257 VNB.n51 VNB.n50 7.01
R258 VNB.n44 VNB.n43 7.01
R259 VNB.n48 VNB.n47 7.01
R260 VNB.n113 VNB.n112 7.01
R261 VNB.n109 VNB.n108 6.788
R262 VNB.n104 VNB.n103 6.788
R263 VNB.n28 VNB.n27 4.551
R264 VNB.n59 VNB.n56 4.305
R265 VNB.n67 VNB.n66 3.947
R266 VNB.n76 VNB.n75 2.511
R267 VNB.t1 VNB.n28 2.238
R268 VNB.n114 VNB.n105 0.921
R269 VNB.n114 VNB.n109 0.476
R270 VNB.n114 VNB.n104 0.475
R271 VNB.n34 VNB.n33 0.358
R272 VNB.n93 VNB.n10 0.272
R273 VNB.n23 VNB.n17 0.246
R274 VNB.n24 VNB.n23 0.246
R275 VNB.n23 VNB.n22 0.246
R276 VNB.n49 VNB.n44 0.246
R277 VNB.n50 VNB.n49 0.246
R278 VNB.n49 VNB.n48 0.246
R279 VNB.n114 VNB.n113 0.246
R280 VNB.n100 VNB 0.198
R281 VNB.n63 VNB.n60 0.179
R282 VNB.n8 VNB.n7 0.136
R283 VNB.n9 VNB.n8 0.136
R284 VNB.n10 VNB.n9 0.136
R285 VNB.n95 VNB.n94 0.136
R286 VNB.n96 VNB.n95 0.136
R287 VNB.n97 VNB.n96 0.136
R288 VNB.n98 VNB.n97 0.136
R289 VNB.n99 VNB.n98 0.136
R290 VNB.n100 VNB.n99 0.136
R291 VNB VNB.n93 0.068
R292 VNB.n94 VNB 0.068
C3 VPB VNB 5.42fF
C4 a_112_73.n0 VNB 0.02fF
C5 a_112_73.n1 VNB 0.10fF
C6 a_112_73.n2 VNB 0.07fF
C7 a_112_73.n3 VNB 0.05fF
C8 a_112_73.n4 VNB 0.00fF
C9 a_112_73.n5 VNB 0.04fF
C10 a_112_73.n6 VNB 0.05fF
C11 a_112_73.n7 VNB 0.02fF
C12 a_112_73.n8 VNB 0.05fF
C13 a_112_73.n9 VNB 0.02fF
C14 a_112_73.n10 VNB 0.07fF
C15 a_112_73.n11 VNB 0.17fF
C16 a_112_73.t1 VNB 0.22fF
C17 a_112_73.n12 VNB 0.09fF
C18 a_112_73.n13 VNB 0.00fF
C19 a_851_182.n0 VNB 0.04fF
C20 a_851_182.n1 VNB 1.02fF
C21 a_851_182.n2 VNB 0.04fF
C22 a_851_182.n3 VNB 0.50fF
C23 a_851_182.n4 VNB 0.06fF
C24 VPB.n0 VNB 0.03fF
C25 VPB.n1 VNB 0.03fF
C26 VPB.n2 VNB 0.02fF
C27 VPB.n3 VNB 0.13fF
C28 VPB.n5 VNB 0.02fF
C29 VPB.n6 VNB 0.02fF
C30 VPB.n7 VNB 0.02fF
C31 VPB.n8 VNB 0.02fF
C32 VPB.n10 VNB 0.02fF
C33 VPB.n11 VNB 0.02fF
C34 VPB.n12 VNB 0.02fF
C35 VPB.n14 VNB 0.22fF
C36 VPB.n15 VNB 0.02fF
C37 VPB.n16 VNB 0.01fF
C38 VPB.n17 VNB 0.07fF
C39 VPB.n18 VNB 0.02fF
C40 VPB.n19 VNB 0.02fF
C41 VPB.n20 VNB 0.03fF
C42 VPB.n21 VNB 0.02fF
C43 VPB.n22 VNB 0.02fF
C44 VPB.n23 VNB 0.02fF
C45 VPB.n24 VNB 0.03fF
C46 VPB.n25 VNB 0.02fF
C47 VPB.n26 VNB 0.16fF
C48 VPB.n27 VNB 0.04fF
C49 VPB.n29 VNB 0.02fF
C50 VPB.n30 VNB 0.02fF
C51 VPB.n31 VNB 0.02fF
C52 VPB.n32 VNB 0.02fF
C53 VPB.n34 VNB 0.02fF
C54 VPB.n35 VNB 0.02fF
C55 VPB.n36 VNB 0.02fF
C56 VPB.n38 VNB 0.25fF
C57 VPB.n40 VNB 0.02fF
C58 VPB.n41 VNB 0.02fF
C59 VPB.n42 VNB 0.02fF
C60 VPB.n43 VNB 0.02fF
C61 VPB.n44 VNB 0.02fF
C62 VPB.n45 VNB 0.10fF
C63 VPB.n46 VNB 0.02fF
C64 VPB.n47 VNB 0.02fF
C65 VPB.n48 VNB 0.04fF
C66 VPB.n49 VNB 0.01fF
C67 VPB.n51 VNB 0.02fF
C68 VPB.n52 VNB 0.02fF
C69 VPB.n53 VNB 0.02fF
C70 VPB.n54 VNB 0.02fF
C71 VPB.n56 VNB 0.02fF
C72 VPB.n59 VNB 0.42fF
C73 VPB.n61 VNB 0.03fF
C74 VPB.n62 VNB 0.04fF
C75 VPB.n63 VNB 0.25fF
C76 VPB.n64 VNB 0.03fF
C77 VPB.n65 VNB 0.03fF
C78 VPB.n66 VNB 0.05fF
C79 VPB.n67 VNB 0.13fF
C80 VPB.n68 VNB 0.18fF
C81 VPB.n69 VNB 0.02fF
C82 VPB.n70 VNB 0.01fF
C83 VPB.n71 VNB 0.15fF
C84 VPB.n72 VNB 0.02fF
C85 VPB.n73 VNB 0.02fF
C86 VPB.n74 VNB 0.13fF
C87 VPB.n75 VNB 0.18fF
C88 VPB.n76 VNB 0.02fF
C89 VPB.n77 VNB 0.01fF
C90 VPB.n78 VNB 0.05fF
C91 VPB.n79 VNB 0.25fF
C92 VPB.n80 VNB 0.01fF
C93 VPB.n81 VNB 0.02fF
C94 VPB.n82 VNB 0.03fF
C95 VPB.n83 VNB 0.09fF
C96 VPB.n84 VNB 0.05fF
C97 VPB.n85 VNB 0.13fF
C98 VPB.n86 VNB 0.15fF
C99 VPB.n87 VNB 0.02fF
C100 VPB.n88 VNB 0.02fF
C101 VPB.n89 VNB 0.13fF
C102 VPB.n90 VNB 0.14fF
C103 VPB.n91 VNB 0.02fF
C104 VPB.n92 VNB 0.02fF
C105 VPB.n93 VNB 0.02fF
C106 VPB.n94 VNB 0.13fF
C107 VPB.n95 VNB 0.14fF
C108 VPB.n96 VNB 0.02fF
C109 VPB.n97 VNB 0.02fF
C110 VPB.n98 VNB 0.13fF
C111 VPB.n99 VNB 0.15fF
C112 VPB.n100 VNB 0.02fF
C113 VPB.n101 VNB 0.02fF
C114 VPB.n102 VNB 0.05fF
C115 VPB.n103 VNB 0.21fF
C116 VPB.n104 VNB 0.02fF
C117 VPB.n105 VNB 0.01fF
C118 VPB.n106 VNB 0.03fF
C119 VPB.n107 VNB 0.25fF
C120 VPB.n108 VNB 0.01fF
C121 VPB.n109 VNB 0.02fF
C122 VPB.n110 VNB 0.03fF
C123 VPB.n111 VNB 0.02fF
C124 VPB.n112 VNB 0.02fF
C125 VPB.n113 VNB 0.02fF
C126 VPB.n114 VNB 0.02fF
C127 VPB.n115 VNB 0.02fF
C128 VPB.n116 VNB 0.02fF
C129 VPB.n117 VNB 0.03fF
C130 VPB.n118 VNB 0.03fF
C131 VPB.n119 VNB 0.02fF
C132 VPB.n120 VNB 0.02fF
C133 VPB.n121 VNB 0.02fF
C134 VPB.n122 VNB 0.04fF
C135 VPB.n123 VNB 0.03fF
C136 VPB.n125 VNB 0.39fF
C137 a_217_1004.n0 VNB 0.03fF
C138 a_217_1004.n1 VNB 0.42fF
C139 a_217_1004.n2 VNB 0.49fF
C140 a_217_1004.n3 VNB 0.25fF
C141 a_217_1004.n4 VNB 0.28fF
C142 a_217_1004.t7 VNB 0.41fF
C143 a_217_1004.n5 VNB 0.45fF
C144 a_217_1004.n6 VNB 0.44fF
C145 a_217_1004.n7 VNB 0.03fF
C146 a_217_1004.n8 VNB 0.22fF
C147 a_217_1004.n9 VNB 0.04fF
.ends
