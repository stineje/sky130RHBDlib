* SPICE3 file created from AOAI4X1.ext - technology: sky130A

.subckt AOAI4X1 YN A B C D VPB VNB
M1000 VNB a_168_157# a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=2.2948p pd=16.08u as=0p ps=0u
M1001 VNB a_864_181.t6 a_1444_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_1549_1004.t1 a_1675_383# VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t2 a_168_157# a_217_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPB.t8 a_217_1004.t5 a_797_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPB.t5 a_343_383# a_217_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPB.t7 a_864_181.t4 a_1549_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_797_1005.t3 a_1009_383# a_864_181.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_217_1004.t0 a_168_157# VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPB.t0 a_1675_383# a_1549_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_217_1004.t2 a_343_383# VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_797_1005.t0 a_217_1004.t6 VPB.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1549_1004.t3 a_864_181.t5 VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_864_181.t1 a_1009_383# a_797_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 a_343_383# a_168_157# 0.26fF
C1 VPB a_1675_383# 0.07fF
C2 VPB a_168_157# 0.08fF
C3 VPB a_343_383# 0.07fF
C4 VPB a_1009_383# 0.07fF
R0 a_1444_73.t0 a_1444_73.n1 34.62
R1 a_1444_73.t0 a_1444_73.n0 8.137
R2 a_1444_73.t0 a_1444_73.n2 4.69
R3 a_1549_1004.n4 a_1549_1004.n2 363.155
R4 a_1549_1004.n2 a_1549_1004.n1 76.002
R5 a_1549_1004.n4 a_1549_1004.n3 15.218
R6 a_1549_1004.n0 a_1549_1004.t0 14.282
R7 a_1549_1004.n0 a_1549_1004.t1 14.282
R8 a_1549_1004.n1 a_1549_1004.t4 14.282
R9 a_1549_1004.n1 a_1549_1004.t3 14.282
R10 a_1549_1004.n2 a_1549_1004.n0 12.85
R11 a_1549_1004.n5 a_1549_1004.n4 12.014
R12 VPB VPB.n200 126.832
R13 VPB.n51 VPB.n49 94.117
R14 VPB.n123 VPB.n121 94.117
R15 VPB.n176 VPB.n173 76
R16 VPB.n181 VPB.n180 76
R17 VPB.n193 VPB.n192 76
R18 VPB.n21 VPB.n20 61.764
R19 VPB.n84 VPB.n83 61.764
R20 VPB.n74 VPB.t3 55.106
R21 VPB.n113 VPB.t6 55.106
R22 VPB.n56 VPB.t5 55.106
R23 VPB.n159 VPB.t0 55.106
R24 VPB.n156 VPB.n155 48.952
R25 VPB.n58 VPB.n57 48.952
R26 VPB.n110 VPB.n109 44.502
R27 VPB.n39 VPB.n38 44.502
R28 VPB.n71 VPB.n70 44.502
R29 VPB.n37 VPB.n36 41.183
R30 VPB.n65 VPB.n14 40.824
R31 VPB.n104 VPB.n99 40.824
R32 VPB.n164 VPB.n163 35.118
R33 VPB.n197 VPB.n193 20.452
R34 VPB.n154 VPB.n151 20.452
R35 VPB.n101 VPB.n100 17.801
R36 VPB.n62 VPB.n61 17.801
R37 VPB.n14 VPB.t4 14.282
R38 VPB.n14 VPB.t2 14.282
R39 VPB.n36 VPB.t9 14.282
R40 VPB.n36 VPB.t8 14.282
R41 VPB.n99 VPB.t1 14.282
R42 VPB.n99 VPB.t7 14.282
R43 VPB.n154 VPB.n153 13.653
R44 VPB.n153 VPB.n152 13.653
R45 VPB.n162 VPB.n161 13.653
R46 VPB.n161 VPB.n160 13.653
R47 VPB.n158 VPB.n157 13.653
R48 VPB.n157 VPB.n156 13.653
R49 VPB.n103 VPB.n102 13.653
R50 VPB.n102 VPB.n101 13.653
R51 VPB.n108 VPB.n107 13.653
R52 VPB.n107 VPB.n106 13.653
R53 VPB.n112 VPB.n111 13.653
R54 VPB.n111 VPB.n110 13.653
R55 VPB.n116 VPB.n115 13.653
R56 VPB.n115 VPB.n114 13.653
R57 VPB.n119 VPB.n118 13.653
R58 VPB.n118 VPB.n117 13.653
R59 VPB.n124 VPB.n123 13.653
R60 VPB.n123 VPB.n122 13.653
R61 VPB.n127 VPB.n126 13.653
R62 VPB.n126 VPB.n125 13.653
R63 VPB.n130 VPB.n129 13.653
R64 VPB.n129 VPB.n128 13.653
R65 VPB.n176 VPB.n175 13.653
R66 VPB.n175 VPB.n174 13.653
R67 VPB.n180 VPB.n179 13.653
R68 VPB.n179 VPB.n178 13.653
R69 VPB.n41 VPB.n40 13.653
R70 VPB.n40 VPB.n39 13.653
R71 VPB.n44 VPB.n43 13.653
R72 VPB.n43 VPB.n42 13.653
R73 VPB.n47 VPB.n46 13.653
R74 VPB.n46 VPB.n45 13.653
R75 VPB.n52 VPB.n51 13.653
R76 VPB.n51 VPB.n50 13.653
R77 VPB.n55 VPB.n54 13.653
R78 VPB.n54 VPB.n53 13.653
R79 VPB.n60 VPB.n59 13.653
R80 VPB.n59 VPB.n58 13.653
R81 VPB.n64 VPB.n63 13.653
R82 VPB.n63 VPB.n62 13.653
R83 VPB.n69 VPB.n68 13.653
R84 VPB.n68 VPB.n67 13.653
R85 VPB.n73 VPB.n72 13.653
R86 VPB.n72 VPB.n71 13.653
R87 VPB.n77 VPB.n76 13.653
R88 VPB.n76 VPB.n75 13.653
R89 VPB.n193 VPB.n0 13.653
R90 VPB VPB.n0 13.653
R91 VPB.n106 VPB.n105 13.35
R92 VPB.n178 VPB.n177 13.35
R93 VPB.n67 VPB.n66 13.35
R94 VPB.n197 VPB.n196 13.276
R95 VPB.n196 VPB.n194 13.276
R96 VPB.n35 VPB.n17 13.276
R97 VPB.n17 VPB.n15 13.276
R98 VPB.n98 VPB.n80 13.276
R99 VPB.n80 VPB.n78 13.276
R100 VPB.n112 VPB.n108 13.276
R101 VPB.n119 VPB.n116 13.276
R102 VPB.n120 VPB.n119 13.276
R103 VPB.n124 VPB.n120 13.276
R104 VPB.n127 VPB.n124 13.276
R105 VPB.n130 VPB.n127 13.276
R106 VPB.n176 VPB.n130 13.276
R107 VPB.n180 VPB.n176 13.276
R108 VPB.n44 VPB.n41 13.276
R109 VPB.n47 VPB.n44 13.276
R110 VPB.n48 VPB.n47 13.276
R111 VPB.n52 VPB.n48 13.276
R112 VPB.n55 VPB.n52 13.276
R113 VPB.n64 VPB.n60 13.276
R114 VPB.n73 VPB.n69 13.276
R115 VPB.n193 VPB.n77 13.276
R116 VPB.n151 VPB.n133 13.276
R117 VPB.n133 VPB.n131 13.276
R118 VPB.n138 VPB.n136 12.796
R119 VPB.n138 VPB.n137 12.564
R120 VPB.n144 VPB.n143 12.198
R121 VPB.n146 VPB.n145 12.198
R122 VPB.n144 VPB.n141 12.198
R123 VPB.n159 VPB.n158 11.841
R124 VPB.n60 VPB.n56 11.841
R125 VPB.n113 VPB.n112 11.482
R126 VPB.n74 VPB.n73 11.482
R127 VPB.n151 VPB.n150 7.5
R128 VPB.n136 VPB.n135 7.5
R129 VPB.n143 VPB.n142 7.5
R130 VPB.n141 VPB.n140 7.5
R131 VPB.n133 VPB.n132 7.5
R132 VPB.n148 VPB.n134 7.5
R133 VPB.n80 VPB.n79 7.5
R134 VPB.n93 VPB.n92 7.5
R135 VPB.n87 VPB.n86 7.5
R136 VPB.n89 VPB.n88 7.5
R137 VPB.n82 VPB.n81 7.5
R138 VPB.n98 VPB.n97 7.5
R139 VPB.n17 VPB.n16 7.5
R140 VPB.n30 VPB.n29 7.5
R141 VPB.n24 VPB.n23 7.5
R142 VPB.n26 VPB.n25 7.5
R143 VPB.n19 VPB.n18 7.5
R144 VPB.n35 VPB.n34 7.5
R145 VPB.n196 VPB.n195 7.5
R146 VPB.n12 VPB.n11 7.5
R147 VPB.n6 VPB.n5 7.5
R148 VPB.n8 VPB.n7 7.5
R149 VPB.n2 VPB.n1 7.5
R150 VPB.n198 VPB.n197 7.5
R151 VPB.n48 VPB.n35 7.176
R152 VPB.n120 VPB.n98 7.176
R153 VPB.n108 VPB.n104 6.817
R154 VPB.n69 VPB.n65 6.817
R155 VPB.n94 VPB.n91 6.729
R156 VPB.n90 VPB.n87 6.729
R157 VPB.n85 VPB.n82 6.729
R158 VPB.n31 VPB.n28 6.729
R159 VPB.n27 VPB.n24 6.729
R160 VPB.n22 VPB.n19 6.729
R161 VPB.n13 VPB.n10 6.729
R162 VPB.n9 VPB.n6 6.729
R163 VPB.n4 VPB.n2 6.729
R164 VPB.n85 VPB.n84 6.728
R165 VPB.n90 VPB.n89 6.728
R166 VPB.n94 VPB.n93 6.728
R167 VPB.n97 VPB.n96 6.728
R168 VPB.n22 VPB.n21 6.728
R169 VPB.n27 VPB.n26 6.728
R170 VPB.n31 VPB.n30 6.728
R171 VPB.n34 VPB.n33 6.728
R172 VPB.n4 VPB.n3 6.728
R173 VPB.n9 VPB.n8 6.728
R174 VPB.n13 VPB.n12 6.728
R175 VPB.n199 VPB.n198 6.728
R176 VPB.n104 VPB.n103 6.458
R177 VPB.n65 VPB.n64 6.458
R178 VPB.n150 VPB.n149 6.398
R179 VPB.n163 VPB.n154 6.112
R180 VPB.n163 VPB.n162 6.101
R181 VPB.n41 VPB.n37 4.305
R182 VPB.n116 VPB.n113 1.794
R183 VPB.n77 VPB.n74 1.794
R184 VPB.n162 VPB.n159 1.435
R185 VPB.n56 VPB.n55 1.435
R186 VPB.n148 VPB.n139 1.402
R187 VPB.n148 VPB.n144 1.402
R188 VPB.n148 VPB.n146 1.402
R189 VPB.n148 VPB.n147 1.402
R190 VPB.n149 VPB.n148 0.735
R191 VPB.n148 VPB.n138 0.735
R192 VPB.n95 VPB.n94 0.387
R193 VPB.n95 VPB.n90 0.387
R194 VPB.n95 VPB.n85 0.387
R195 VPB.n96 VPB.n95 0.387
R196 VPB.n32 VPB.n31 0.387
R197 VPB.n32 VPB.n27 0.387
R198 VPB.n32 VPB.n22 0.387
R199 VPB.n33 VPB.n32 0.387
R200 VPB.n200 VPB.n13 0.387
R201 VPB.n200 VPB.n9 0.387
R202 VPB.n200 VPB.n4 0.387
R203 VPB.n200 VPB.n199 0.387
R204 VPB.n170 VPB.n169 0.272
R205 VPB.n185 VPB.n184 0.272
R206 VPB.n192 VPB 0.198
R207 VPB.n165 VPB.n164 0.136
R208 VPB.n166 VPB.n165 0.136
R209 VPB.n167 VPB.n166 0.136
R210 VPB.n168 VPB.n167 0.136
R211 VPB.n169 VPB.n168 0.136
R212 VPB.n171 VPB.n170 0.136
R213 VPB.n172 VPB.n171 0.136
R214 VPB.n173 VPB.n172 0.136
R215 VPB.n182 VPB.n181 0.136
R216 VPB.n183 VPB.n182 0.136
R217 VPB.n184 VPB.n183 0.136
R218 VPB.n186 VPB.n185 0.136
R219 VPB.n187 VPB.n186 0.136
R220 VPB.n188 VPB.n187 0.136
R221 VPB.n189 VPB.n188 0.136
R222 VPB.n190 VPB.n189 0.136
R223 VPB.n191 VPB.n190 0.136
R224 VPB.n192 VPB.n191 0.136
R225 VPB.n173 VPB 0.068
R226 VPB.n181 VPB 0.068
R227 a_217_1004.n4 a_217_1004.t6 486.819
R228 a_217_1004.n4 a_217_1004.t5 384.527
R229 a_217_1004.n6 a_217_1004.n3 215.652
R230 a_217_1004.n5 a_217_1004.t7 207.443
R231 a_217_1004.n5 a_217_1004.n4 169.7
R232 a_217_1004.n6 a_217_1004.n5 153.315
R233 a_217_1004.n8 a_217_1004.n6 140.981
R234 a_217_1004.n3 a_217_1004.n2 76.002
R235 a_217_1004.n8 a_217_1004.n7 30
R236 a_217_1004.n9 a_217_1004.n0 24.383
R237 a_217_1004.n9 a_217_1004.n8 23.684
R238 a_217_1004.n1 a_217_1004.t3 14.282
R239 a_217_1004.n1 a_217_1004.t2 14.282
R240 a_217_1004.n2 a_217_1004.t1 14.282
R241 a_217_1004.n2 a_217_1004.t0 14.282
R242 a_217_1004.n3 a_217_1004.n1 12.85
R243 a_797_1005.t1 a_797_1005.n0 101.66
R244 a_797_1005.n0 a_797_1005.t3 101.659
R245 a_797_1005.n0 a_797_1005.t2 14.294
R246 a_797_1005.n0 a_797_1005.t0 14.282
R247 a_864_181.n2 a_864_181.t4 480.392
R248 a_864_181.n2 a_864_181.t5 403.272
R249 a_864_181.n4 a_864_181.n1 228.489
R250 a_864_181.n3 a_864_181.t6 213.869
R251 a_864_181.n3 a_864_181.n2 161.6
R252 a_864_181.n4 a_864_181.n3 153.315
R253 a_864_181.n9 a_864_181.n8 118.016
R254 a_864_181.n9 a_864_181.n4 92.576
R255 a_864_181.n12 a_864_181.n0 55.263
R256 a_864_181.n11 a_864_181.n9 48.405
R257 a_864_181.n8 a_864_181.n7 30
R258 a_864_181.n11 a_864_181.n10 30
R259 a_864_181.n12 a_864_181.n11 25.263
R260 a_864_181.n6 a_864_181.n5 24.383
R261 a_864_181.n8 a_864_181.n6 23.684
R262 a_864_181.n1 a_864_181.t2 14.282
R263 a_864_181.n1 a_864_181.t1 14.282
R264 a_112_73.n10 a_112_73.n9 93.333
R265 a_112_73.n2 a_112_73.n1 41.622
R266 a_112_73.n13 a_112_73.n12 26.667
R267 a_112_73.n6 a_112_73.n5 24.977
R268 a_112_73.t0 a_112_73.n2 21.209
R269 a_112_73.t0 a_112_73.n3 11.595
R270 a_112_73.t1 a_112_73.n8 8.137
R271 a_112_73.t0 a_112_73.n0 6.109
R272 a_112_73.t1 a_112_73.n7 4.864
R273 a_112_73.t0 a_112_73.n4 3.871
R274 a_112_73.t0 a_112_73.n13 2.535
R275 a_112_73.n13 a_112_73.t1 1.145
R276 a_112_73.n7 a_112_73.n6 1.13
R277 a_112_73.t1 a_112_73.n11 0.804
R278 a_112_73.n11 a_112_73.n10 0.136
R279 VNB VNB.n180 300.778
R280 VNB.n76 VNB.n75 199.897
R281 VNB.n15 VNB.n14 199.897
R282 VNB.n102 VNB.n100 154.509
R283 VNB.n38 VNB.n36 154.509
R284 VNB.n89 VNB.n82 84.842
R285 VNB.n52 VNB.n4 84.842
R286 VNB.n167 VNB.n166 76
R287 VNB.n155 VNB.n154 76
R288 VNB.n149 VNB.n146 76
R289 VNB.n152 VNB.n151 36.937
R290 VNB.n91 VNB.n90 36.678
R291 VNB.n54 VNB.n53 36.678
R292 VNB.n109 VNB.n108 36.267
R293 VNB.n137 VNB.n136 35.118
R294 VNB.n129 VNB.n126 20.452
R295 VNB.n168 VNB.n167 20.452
R296 VNB.n25 VNB.n24 19.735
R297 VNB.n150 VNB.n61 19.735
R298 VNB.n111 VNB.n62 19.735
R299 VNB.n104 VNB.n65 19.735
R300 VNB.n31 VNB.n23 19.735
R301 VNB.n22 VNB.t0 17.353
R302 VNB.n60 VNB.t1 13.654
R303 VNB.n135 VNB.n134 13.653
R304 VNB.n134 VNB.n133 13.653
R305 VNB.n132 VNB.n131 13.653
R306 VNB.n131 VNB.n130 13.653
R307 VNB.n85 VNB.n84 13.653
R308 VNB.n84 VNB.n83 13.653
R309 VNB.n88 VNB.n87 13.653
R310 VNB.n87 VNB.n86 13.653
R311 VNB.n92 VNB.n91 13.653
R312 VNB.n95 VNB.n94 13.653
R313 VNB.n94 VNB.n93 13.653
R314 VNB.n98 VNB.n97 13.653
R315 VNB.n97 VNB.n96 13.653
R316 VNB.n103 VNB.n102 13.653
R317 VNB.n102 VNB.n101 13.653
R318 VNB.n107 VNB.n106 13.653
R319 VNB.n106 VNB.n105 13.653
R320 VNB.n110 VNB.n109 13.653
R321 VNB.n149 VNB.n148 13.653
R322 VNB.n148 VNB.n147 13.653
R323 VNB.n154 VNB.n153 13.653
R324 VNB.n153 VNB.n152 13.653
R325 VNB.n27 VNB.n26 13.653
R326 VNB.n30 VNB.n29 13.653
R327 VNB.n29 VNB.n28 13.653
R328 VNB.n34 VNB.n33 13.653
R329 VNB.n33 VNB.n32 13.653
R330 VNB.n39 VNB.n38 13.653
R331 VNB.n38 VNB.n37 13.653
R332 VNB.n42 VNB.n41 13.653
R333 VNB.n41 VNB.n40 13.653
R334 VNB.n45 VNB.n44 13.653
R335 VNB.n44 VNB.n43 13.653
R336 VNB.n48 VNB.n47 13.653
R337 VNB.n47 VNB.n46 13.653
R338 VNB.n51 VNB.n50 13.653
R339 VNB.n50 VNB.n49 13.653
R340 VNB.n55 VNB.n54 13.653
R341 VNB.n58 VNB.n57 13.653
R342 VNB.n57 VNB.n56 13.653
R343 VNB.n167 VNB.n0 13.653
R344 VNB VNB.n0 13.653
R345 VNB.n129 VNB.n128 13.653
R346 VNB.n128 VNB.n127 13.653
R347 VNB.n175 VNB.n172 13.577
R348 VNB.n114 VNB.n112 13.276
R349 VNB.n126 VNB.n114 13.276
R350 VNB.n68 VNB.n66 13.276
R351 VNB.n81 VNB.n68 13.276
R352 VNB.n7 VNB.n5 13.276
R353 VNB.n20 VNB.n7 13.276
R354 VNB.n135 VNB.n132 13.276
R355 VNB.n88 VNB.n85 13.276
R356 VNB.n95 VNB.n92 13.276
R357 VNB.n98 VNB.n95 13.276
R358 VNB.n99 VNB.n98 13.276
R359 VNB.n103 VNB.n99 13.276
R360 VNB.n110 VNB.n107 13.276
R361 VNB.n30 VNB.n27 13.276
R362 VNB.n35 VNB.n34 13.276
R363 VNB.n39 VNB.n35 13.276
R364 VNB.n42 VNB.n39 13.276
R365 VNB.n45 VNB.n42 13.276
R366 VNB.n48 VNB.n45 13.276
R367 VNB.n51 VNB.n48 13.276
R368 VNB.n58 VNB.n55 13.276
R369 VNB.n167 VNB.n58 13.276
R370 VNB.n3 VNB.n1 13.276
R371 VNB.n168 VNB.n3 13.276
R372 VNB.n23 VNB.n22 12.837
R373 VNB.n104 VNB.n103 11.661
R374 VNB.n34 VNB.n31 11.661
R375 VNB.n65 VNB.n64 11.605
R376 VNB.n89 VNB.n88 10.764
R377 VNB.n149 VNB.n111 10.764
R378 VNB.n52 VNB.n51 10.764
R379 VNB.n64 VNB.n63 9.809
R380 VNB.n22 VNB.n21 7.566
R381 VNB.n177 VNB.n176 7.5
R382 VNB.n74 VNB.n73 7.5
R383 VNB.n70 VNB.n69 7.5
R384 VNB.n68 VNB.n67 7.5
R385 VNB.n81 VNB.n80 7.5
R386 VNB.n13 VNB.n12 7.5
R387 VNB.n9 VNB.n8 7.5
R388 VNB.n7 VNB.n6 7.5
R389 VNB.n20 VNB.n19 7.5
R390 VNB.n169 VNB.n168 7.5
R391 VNB.n3 VNB.n2 7.5
R392 VNB.n174 VNB.n173 7.5
R393 VNB.n120 VNB.n119 7.5
R394 VNB.n116 VNB.n115 7.5
R395 VNB.n114 VNB.n113 7.5
R396 VNB.n126 VNB.n125 7.5
R397 VNB.n99 VNB.n81 7.176
R398 VNB.n35 VNB.n20 7.176
R399 VNB.t1 VNB.n59 7.04
R400 VNB.n179 VNB.n177 7.011
R401 VNB.n77 VNB.n74 7.011
R402 VNB.n72 VNB.n70 7.011
R403 VNB.n16 VNB.n13 7.011
R404 VNB.n11 VNB.n9 7.011
R405 VNB.n122 VNB.n120 7.011
R406 VNB.n118 VNB.n116 7.011
R407 VNB.n80 VNB.n79 7.01
R408 VNB.n72 VNB.n71 7.01
R409 VNB.n77 VNB.n76 7.01
R410 VNB.n19 VNB.n18 7.01
R411 VNB.n11 VNB.n10 7.01
R412 VNB.n16 VNB.n15 7.01
R413 VNB.n125 VNB.n124 7.01
R414 VNB.n118 VNB.n117 7.01
R415 VNB.n122 VNB.n121 7.01
R416 VNB.n179 VNB.n178 7.01
R417 VNB.n175 VNB.n174 6.788
R418 VNB.n170 VNB.n169 6.788
R419 VNB.n150 VNB.n149 6.638
R420 VNB.n154 VNB.n150 6.638
R421 VNB.n136 VNB.n129 6.111
R422 VNB.n136 VNB.n135 6.1
R423 VNB.n61 VNB.n60 5.774
R424 VNB.n92 VNB.n89 2.511
R425 VNB.n111 VNB.n110 2.511
R426 VNB.n27 VNB.n25 2.511
R427 VNB.n55 VNB.n52 2.511
R428 VNB.n107 VNB.n104 1.614
R429 VNB.n31 VNB.n30 1.614
R430 VNB.n180 VNB.n171 0.921
R431 VNB.n180 VNB.n175 0.476
R432 VNB.n180 VNB.n170 0.475
R433 VNB.n143 VNB.n142 0.272
R434 VNB.n159 VNB.n158 0.272
R435 VNB.n78 VNB.n72 0.246
R436 VNB.n79 VNB.n78 0.246
R437 VNB.n78 VNB.n77 0.246
R438 VNB.n17 VNB.n11 0.246
R439 VNB.n18 VNB.n17 0.246
R440 VNB.n17 VNB.n16 0.246
R441 VNB.n123 VNB.n118 0.246
R442 VNB.n124 VNB.n123 0.246
R443 VNB.n123 VNB.n122 0.246
R444 VNB.n180 VNB.n179 0.246
R445 VNB.n166 VNB 0.198
R446 VNB.n138 VNB.n137 0.136
R447 VNB.n139 VNB.n138 0.136
R448 VNB.n140 VNB.n139 0.136
R449 VNB.n141 VNB.n140 0.136
R450 VNB.n142 VNB.n141 0.136
R451 VNB.n144 VNB.n143 0.136
R452 VNB.n145 VNB.n144 0.136
R453 VNB.n146 VNB.n145 0.136
R454 VNB.n156 VNB.n155 0.136
R455 VNB.n157 VNB.n156 0.136
R456 VNB.n158 VNB.n157 0.136
R457 VNB.n160 VNB.n159 0.136
R458 VNB.n161 VNB.n160 0.136
R459 VNB.n162 VNB.n161 0.136
R460 VNB.n163 VNB.n162 0.136
R461 VNB.n164 VNB.n163 0.136
R462 VNB.n165 VNB.n164 0.136
R463 VNB.n166 VNB.n165 0.136
R464 VNB.n146 VNB 0.068
R465 VNB.n155 VNB 0.068
C5 VPB VNB 8.64fF
C6 a_112_73.n0 VNB 0.02fF
C7 a_112_73.n1 VNB 0.10fF
C8 a_112_73.n2 VNB 0.07fF
C9 a_112_73.n3 VNB 0.05fF
C10 a_112_73.n4 VNB 0.00fF
C11 a_112_73.n5 VNB 0.04fF
C12 a_112_73.n6 VNB 0.05fF
C13 a_112_73.n7 VNB 0.02fF
C14 a_112_73.n8 VNB 0.05fF
C15 a_112_73.n9 VNB 0.02fF
C16 a_112_73.n10 VNB 0.07fF
C17 a_112_73.n11 VNB 0.17fF
C18 a_112_73.t1 VNB 0.22fF
C19 a_112_73.n12 VNB 0.09fF
C20 a_112_73.n13 VNB 0.00fF
C21 a_864_181.n0 VNB 0.04fF
C22 a_864_181.n1 VNB 0.62fF
C23 a_864_181.n2 VNB 0.38fF
C24 a_864_181.n3 VNB 0.46fF
C25 a_864_181.n4 VNB 0.46fF
C26 a_864_181.n5 VNB 0.03fF
C27 a_864_181.n6 VNB 0.05fF
C28 a_864_181.n7 VNB 0.03fF
C29 a_864_181.n8 VNB 0.15fF
C30 a_864_181.n9 VNB 0.26fF
C31 a_864_181.n10 VNB 0.03fF
C32 a_864_181.n11 VNB 0.08fF
C33 a_864_181.n12 VNB 0.04fF
C34 a_797_1005.n0 VNB 0.55fF
C35 a_217_1004.n0 VNB 0.03fF
C36 a_217_1004.n1 VNB 0.43fF
C37 a_217_1004.n2 VNB 0.51fF
C38 a_217_1004.n3 VNB 0.31fF
C39 a_217_1004.n4 VNB 0.35fF
C40 a_217_1004.t7 VNB 0.38fF
C41 a_217_1004.n5 VNB 0.45fF
C42 a_217_1004.n6 VNB 0.49fF
C43 a_217_1004.n7 VNB 0.03fF
C44 a_217_1004.n8 VNB 0.17fF
C45 a_217_1004.n9 VNB 0.04fF
C46 VPB.n0 VNB 0.03fF
C47 VPB.n1 VNB 0.04fF
C48 VPB.n2 VNB 0.02fF
C49 VPB.n3 VNB 0.13fF
C50 VPB.n5 VNB 0.02fF
C51 VPB.n6 VNB 0.02fF
C52 VPB.n7 VNB 0.02fF
C53 VPB.n8 VNB 0.02fF
C54 VPB.n10 VNB 0.02fF
C55 VPB.n11 VNB 0.02fF
C56 VPB.n12 VNB 0.02fF
C57 VPB.n14 VNB 0.10fF
C58 VPB.n15 VNB 0.02fF
C59 VPB.n16 VNB 0.02fF
C60 VPB.n17 VNB 0.02fF
C61 VPB.n18 VNB 0.04fF
C62 VPB.n19 VNB 0.02fF
C63 VPB.n20 VNB 0.19fF
C64 VPB.n21 VNB 0.04fF
C65 VPB.n23 VNB 0.02fF
C66 VPB.n24 VNB 0.02fF
C67 VPB.n25 VNB 0.02fF
C68 VPB.n26 VNB 0.02fF
C69 VPB.n28 VNB 0.02fF
C70 VPB.n29 VNB 0.02fF
C71 VPB.n30 VNB 0.02fF
C72 VPB.n32 VNB 0.26fF
C73 VPB.n34 VNB 0.02fF
C74 VPB.n35 VNB 0.02fF
C75 VPB.n36 VNB 0.10fF
C76 VPB.n37 VNB 0.02fF
C77 VPB.n38 VNB 0.13fF
C78 VPB.n39 VNB 0.16fF
C79 VPB.n40 VNB 0.02fF
C80 VPB.n41 VNB 0.02fF
C81 VPB.n42 VNB 0.23fF
C82 VPB.n43 VNB 0.02fF
C83 VPB.n44 VNB 0.02fF
C84 VPB.n45 VNB 0.26fF
C85 VPB.n46 VNB 0.01fF
C86 VPB.n47 VNB 0.02fF
C87 VPB.n48 VNB 0.03fF
C88 VPB.n49 VNB 0.03fF
C89 VPB.n50 VNB 0.26fF
C90 VPB.n51 VNB 0.01fF
C91 VPB.n52 VNB 0.02fF
C92 VPB.n53 VNB 0.22fF
C93 VPB.n54 VNB 0.02fF
C94 VPB.n55 VNB 0.01fF
C95 VPB.n56 VNB 0.05fF
C96 VPB.n57 VNB 0.13fF
C97 VPB.n58 VNB 0.16fF
C98 VPB.n59 VNB 0.02fF
C99 VPB.n60 VNB 0.02fF
C100 VPB.n61 VNB 0.13fF
C101 VPB.n62 VNB 0.15fF
C102 VPB.n63 VNB 0.02fF
C103 VPB.n64 VNB 0.02fF
C104 VPB.n65 VNB 0.02fF
C105 VPB.n66 VNB 0.13fF
C106 VPB.n67 VNB 0.14fF
C107 VPB.n68 VNB 0.02fF
C108 VPB.n69 VNB 0.02fF
C109 VPB.n70 VNB 0.13fF
C110 VPB.n71 VNB 0.16fF
C111 VPB.n72 VNB 0.02fF
C112 VPB.n73 VNB 0.02fF
C113 VPB.n74 VNB 0.06fF
C114 VPB.n75 VNB 0.23fF
C115 VPB.n76 VNB 0.02fF
C116 VPB.n77 VNB 0.01fF
C117 VPB.n78 VNB 0.02fF
C118 VPB.n79 VNB 0.02fF
C119 VPB.n80 VNB 0.02fF
C120 VPB.n81 VNB 0.04fF
C121 VPB.n82 VNB 0.02fF
C122 VPB.n83 VNB 0.19fF
C123 VPB.n84 VNB 0.04fF
C124 VPB.n86 VNB 0.02fF
C125 VPB.n87 VNB 0.02fF
C126 VPB.n88 VNB 0.02fF
C127 VPB.n89 VNB 0.02fF
C128 VPB.n91 VNB 0.02fF
C129 VPB.n92 VNB 0.02fF
C130 VPB.n93 VNB 0.02fF
C131 VPB.n95 VNB 0.26fF
C132 VPB.n97 VNB 0.02fF
C133 VPB.n98 VNB 0.02fF
C134 VPB.n99 VNB 0.10fF
C135 VPB.n100 VNB 0.13fF
C136 VPB.n101 VNB 0.15fF
C137 VPB.n102 VNB 0.02fF
C138 VPB.n103 VNB 0.02fF
C139 VPB.n104 VNB 0.02fF
C140 VPB.n105 VNB 0.13fF
C141 VPB.n106 VNB 0.14fF
C142 VPB.n107 VNB 0.02fF
C143 VPB.n108 VNB 0.02fF
C144 VPB.n109 VNB 0.13fF
C145 VPB.n110 VNB 0.16fF
C146 VPB.n111 VNB 0.02fF
C147 VPB.n112 VNB 0.02fF
C148 VPB.n113 VNB 0.06fF
C149 VPB.n114 VNB 0.23fF
C150 VPB.n115 VNB 0.02fF
C151 VPB.n116 VNB 0.01fF
C152 VPB.n117 VNB 0.26fF
C153 VPB.n118 VNB 0.01fF
C154 VPB.n119 VNB 0.02fF
C155 VPB.n120 VNB 0.03fF
C156 VPB.n121 VNB 0.03fF
C157 VPB.n122 VNB 0.26fF
C158 VPB.n123 VNB 0.01fF
C159 VPB.n124 VNB 0.02fF
C160 VPB.n125 VNB 0.26fF
C161 VPB.n126 VNB 0.02fF
C162 VPB.n127 VNB 0.02fF
C163 VPB.n128 VNB 0.26fF
C164 VPB.n129 VNB 0.02fF
C165 VPB.n130 VNB 0.02fF
C166 VPB.n131 VNB 0.02fF
C167 VPB.n132 VNB 0.02fF
C168 VPB.n133 VNB 0.02fF
C169 VPB.n134 VNB 0.13fF
C170 VPB.n135 VNB 0.03fF
C171 VPB.n136 VNB 0.02fF
C172 VPB.n137 VNB 0.04fF
C173 VPB.n138 VNB 0.01fF
C174 VPB.n140 VNB 0.02fF
C175 VPB.n141 VNB 0.02fF
C176 VPB.n142 VNB 0.02fF
C177 VPB.n143 VNB 0.02fF
C178 VPB.n145 VNB 0.02fF
C179 VPB.n148 VNB 0.44fF
C180 VPB.n150 VNB 0.03fF
C181 VPB.n151 VNB 0.04fF
C182 VPB.n152 VNB 0.26fF
C183 VPB.n153 VNB 0.03fF
C184 VPB.n154 VNB 0.03fF
C185 VPB.n155 VNB 0.13fF
C186 VPB.n156 VNB 0.16fF
C187 VPB.n157 VNB 0.02fF
C188 VPB.n158 VNB 0.02fF
C189 VPB.n159 VNB 0.05fF
C190 VPB.n160 VNB 0.22fF
C191 VPB.n161 VNB 0.02fF
C192 VPB.n162 VNB 0.01fF
C193 VPB.n163 VNB 0.00fF
C194 VPB.n164 VNB 0.09fF
C195 VPB.n165 VNB 0.02fF
C196 VPB.n166 VNB 0.02fF
C197 VPB.n167 VNB 0.02fF
C198 VPB.n168 VNB 0.02fF
C199 VPB.n169 VNB 0.03fF
C200 VPB.n170 VNB 0.03fF
C201 VPB.n171 VNB 0.02fF
C202 VPB.n172 VNB 0.02fF
C203 VPB.n173 VNB 0.02fF
C204 VPB.n174 VNB 0.26fF
C205 VPB.n175 VNB 0.02fF
C206 VPB.n176 VNB 0.02fF
C207 VPB.n177 VNB 0.13fF
C208 VPB.n178 VNB 0.14fF
C209 VPB.n179 VNB 0.02fF
C210 VPB.n180 VNB 0.02fF
C211 VPB.n181 VNB 0.02fF
C212 VPB.n182 VNB 0.02fF
C213 VPB.n183 VNB 0.02fF
C214 VPB.n184 VNB 0.03fF
C215 VPB.n185 VNB 0.03fF
C216 VPB.n186 VNB 0.02fF
C217 VPB.n187 VNB 0.02fF
C218 VPB.n188 VNB 0.02fF
C219 VPB.n189 VNB 0.02fF
C220 VPB.n190 VNB 0.02fF
C221 VPB.n191 VNB 0.02fF
C222 VPB.n192 VNB 0.03fF
C223 VPB.n193 VNB 0.03fF
C224 VPB.n194 VNB 0.02fF
C225 VPB.n195 VNB 0.02fF
C226 VPB.n196 VNB 0.02fF
C227 VPB.n197 VNB 0.04fF
C228 VPB.n198 VNB 0.03fF
C229 VPB.n200 VNB 0.41fF
C230 a_1549_1004.n0 VNB 0.47fF
C231 a_1549_1004.n1 VNB 0.56fF
C232 a_1549_1004.n2 VNB 0.49fF
C233 a_1549_1004.n3 VNB 0.07fF
C234 a_1549_1004.n4 VNB 0.41fF
C235 a_1549_1004.n5 VNB 0.04fF
C236 a_1444_73.n0 VNB 0.05fF
C237 a_1444_73.n1 VNB 0.12fF
C238 a_1444_73.n2 VNB 0.04fF
.ends
