magic
tech sky130A
magscale 1 2
timestamp 1648062456
<< nmos >>
tri 146 215 162 231 se
rect 162 215 192 276
tri 56 185 86 215 se
rect 86 185 192 215
rect 56 84 86 185
tri 86 169 102 185 nw
tri 146 169 162 185 ne
tri 86 84 102 100 sw
tri 146 84 162 100 se
rect 162 84 192 185
tri 56 54 86 84 ne
rect 86 54 162 84
tri 162 54 192 84 nw
<< ndiff >>
rect 0 260 162 276
rect 0 226 10 260
rect 44 226 107 260
rect 141 231 162 260
rect 141 226 146 231
rect 0 215 146 226
tri 146 215 162 231 nw
rect 192 260 248 276
rect 192 226 204 260
rect 238 226 248 260
rect 0 188 56 215
rect 0 154 10 188
rect 44 154 56 188
tri 56 185 86 215 nw
rect 192 188 248 226
rect 0 120 56 154
rect 0 86 10 120
rect 44 86 56 120
rect 0 54 56 86
tri 86 169 102 185 se
rect 102 169 146 185
tri 146 169 162 185 sw
rect 86 135 162 169
rect 86 101 107 135
rect 141 101 162 135
rect 86 100 162 101
tri 86 84 102 100 ne
rect 102 84 146 100
tri 146 84 162 100 nw
rect 192 154 204 188
rect 238 154 248 188
rect 192 120 248 154
rect 192 86 204 120
rect 238 86 248 120
tri 56 54 86 84 sw
tri 162 54 192 84 se
rect 192 54 248 86
rect 0 50 248 54
rect 0 16 10 50
rect 44 16 204 50
rect 238 16 248 50
rect 0 0 248 16
<< ndiffc >>
rect 10 226 44 260
rect 107 226 141 260
rect 204 226 238 260
rect 10 154 44 188
rect 10 86 44 120
rect 107 101 141 135
rect 204 154 238 188
rect 204 86 238 120
rect 10 16 44 50
rect 204 16 238 50
<< poly >>
rect 162 276 192 302
<< locali >>
rect 10 260 44 276
rect 204 260 238 276
rect 44 226 107 260
rect 141 226 204 260
rect 10 188 44 226
rect 10 120 44 154
rect 204 188 238 226
rect 10 50 44 86
rect 107 135 141 151
rect 107 85 141 101
rect 204 120 238 154
rect 10 0 44 16
rect 204 50 238 86
rect 204 0 238 16
<< end >>
