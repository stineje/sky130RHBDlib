magic
tech sky130A
magscale 1 2
timestamp 1654964768
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 131 871 165 905
rect 279 871 313 905
rect 131 797 165 831
rect 279 797 313 831
rect 131 723 165 757
rect 279 723 313 757
rect 131 649 165 683
rect 279 649 313 683
rect 131 575 165 609
rect 279 575 313 609
rect 131 501 165 535
rect 279 501 313 535
rect 131 427 165 461
rect 279 427 313 461
<< metal1 >>
rect -34 1446 478 1514
rect -34 -34 478 34
use invx1_pcell  invx1_pcell_0 pcells
timestamp 1652329846
transform 1 0 0 0 1 0
box -87 -34 531 1550
<< labels >>
rlabel locali 279 649 313 683 1 Y
port 1 nsew signal output
rlabel locali 279 723 313 757 1 Y
port 1 nsew signal output
rlabel locali 279 797 313 831 1 Y
port 1 nsew signal output
rlabel locali 279 575 313 609 1 Y
port 1 nsew signal output
rlabel locali 279 871 313 905 1 Y
port 1 nsew signal output
rlabel locali 279 501 313 535 1 Y
port 1 nsew signal output
rlabel locali 279 427 313 461 1 Y
port 1 nsew signal output
rlabel locali 131 649 165 683 1 A
port 2 nsew signal input
rlabel locali 131 723 165 757 1 A
port 2 nsew signal input
rlabel locali 131 797 165 831 1 A
port 2 nsew signal input
rlabel locali 131 575 165 609 1 A
port 2 nsew signal input
rlabel locali 131 871 165 905 1 A
port 2 nsew signal input
rlabel locali 131 501 165 535 1 A
port 2 nsew signal input
rlabel locali 131 427 165 461 1 A
port 2 nsew signal input
rlabel metal1 -34 1446 478 1514 1 VPWR
port 3 nsew power bidirectional abutment
rlabel metal1 -34 -34 478 34 1 VGND
port 4 nsew ground bidirectional abutment
rlabel nwell 57 1463 91 1497 1 VPB
rlabel pwell 57 -17 91 17 1 VNB
<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 444 1480
string LEFsymmetry X Y R90
<< end >>
