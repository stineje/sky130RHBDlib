* SPICE3 file created from DFFSNRNQNX1.ext - technology: sky130A

.subckt DFFSNRNQNX1 QN D CLK RN SN VPB VNB
M1000 a_4447_943.t1 SN.t0 VPB.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VNB QN a_4901_75.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1002 VPB.t35 a_147_159# a_277_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_599_943.t6 CLK VPB.t32 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPB.t33 CLK a_1561_943.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPB.t24 a_277_1004.t7 a_2201_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPB.t3 RN a_277_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 QN a_4447_943.t7 a_4220_182.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1008 a_599_943.t4 a_1561_943.t8 VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPB.t14 SN.t1 a_2201_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t4 RN a_1561_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 QN a_599_943.t7 VPB.t13 pshort w=2u l=0.15u
+  ad=1.74p pd=13.74u as=0p ps=0u
M1012 a_1561_943.t5 CLK VPB.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 QN a_4447_943.t8 VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VNB a_147_159# a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPB.t20 a_599_943.t8 a_277_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 QN RN VPB.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPB.t11 a_1561_943.t11 a_2201_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1561_943.t3 a_2201_1004.t8 VPB.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPB.t26 QN a_4447_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_277_1004.t5 a_147_159# VPB.t34 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPB.t23 a_277_1004.t10 a_599_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t9 a_1561_943.t12 a_599_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPB.t16 SN.t3 a_4447_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VNB a_277_1004.t8 a_2015_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_277_1004.t0 RN VPB.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPB.t31 CLK a_599_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_2201_1004.t2 SN.t5 VPB.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1561_943.t1 RN VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPB.t6 RN QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPB.t27 a_1561_943.t13 a_4447_943.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_599_943.t0 a_277_1004.t11 VPB.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_277_1004.t2 a_599_943.t10 VPB.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 VNB a_2201_1004.t7 a_2977_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1034 VNB a_277_1004.t9 a_1053_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_2201_1004.t0 a_277_1004.t12 VPB.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_2201_1004.t4 a_1561_943.t14 VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPB.t19 a_599_943.t12 QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPB.t18 a_4447_943.t9 QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_4447_943.t2 QN VPB.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_4447_943.t6 a_1561_943.t15 VPB.t29 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 VNB a_599_943.t9 a_3939_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPB.t28 a_2201_1004.t9 a_1561_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u











R0 SN.n2 SN.t1 479.223
R1 SN.n0 SN.t3 479.223
R2 SN.n2 SN.t5 375.52
R3 SN.n0 SN.t0 375.52
R4 SN.n3 SN.t2 172.454
R5 SN.n1 SN.t4 172.096
R6 SN.n1 SN.n0 158.923
R7 SN.n3 SN.n2 158.564
R8 SN.n4 SN.n1 86.564
R9 SN.n4 SN.n3 76
R10 SN.n4 SN 0.046
R11 VPB VPB.n513 126.832
R12 VPB.n40 VPB.n38 94.117
R13 VPB.n435 VPB.n433 94.117
R14 VPB.n352 VPB.n350 94.117
R15 VPB.n129 VPB.n127 94.117
R16 VPB.n275 VPB.n273 94.117
R17 VPB.n199 VPB.n198 84.554
R18 VPB.n288 VPB.n287 80.104
R19 VPB.n139 VPB.n138 80.104
R20 VPB.n365 VPB.n364 80.104
R21 VPB.n448 VPB.n447 80.104
R22 VPB.n50 VPB.n49 80.104
R23 VPB.n215 VPB.n214 76
R24 VPB.n220 VPB.n219 76
R25 VPB.n225 VPB.n224 76
R26 VPB.n232 VPB.n231 76
R27 VPB.n237 VPB.n236 76
R28 VPB.n242 VPB.n241 76
R29 VPB.n246 VPB.n245 76
R30 VPB.n250 VPB.n249 76
R31 VPB.n277 VPB.n276 76
R32 VPB.n281 VPB.n280 76
R33 VPB.n286 VPB.n285 76
R34 VPB.n291 VPB.n290 76
R35 VPB.n298 VPB.n297 76
R36 VPB.n303 VPB.n302 76
R37 VPB.n308 VPB.n307 76
R38 VPB.n315 VPB.n314 76
R39 VPB.n320 VPB.n319 76
R40 VPB.n325 VPB.n324 76
R41 VPB.n329 VPB.n328 76
R42 VPB.n333 VPB.n332 76
R43 VPB.n348 VPB.n345 76
R44 VPB.n354 VPB.n353 76
R45 VPB.n358 VPB.n357 76
R46 VPB.n363 VPB.n362 76
R47 VPB.n368 VPB.n367 76
R48 VPB.n375 VPB.n374 76
R49 VPB.n380 VPB.n379 76
R50 VPB.n385 VPB.n384 76
R51 VPB.n392 VPB.n391 76
R52 VPB.n397 VPB.n396 76
R53 VPB.n402 VPB.n401 76
R54 VPB.n406 VPB.n405 76
R55 VPB.n410 VPB.n409 76
R56 VPB.n437 VPB.n436 76
R57 VPB.n441 VPB.n440 76
R58 VPB.n446 VPB.n445 76
R59 VPB.n451 VPB.n450 76
R60 VPB.n458 VPB.n457 76
R61 VPB.n463 VPB.n462 76
R62 VPB.n468 VPB.n467 76
R63 VPB.n475 VPB.n474 76
R64 VPB.n480 VPB.n479 76
R65 VPB.n485 VPB.n484 76
R66 VPB.n489 VPB.n488 76
R67 VPB.n493 VPB.n492 76
R68 VPB.n506 VPB.n505 76
R69 VPB.n234 VPB.n233 75.654
R70 VPB.n317 VPB.n316 75.654
R71 VPB.n161 VPB.n160 75.654
R72 VPB.n394 VPB.n393 75.654
R73 VPB.n477 VPB.n476 75.654
R74 VPB.n72 VPB.n71 75.654
R75 VPB.n22 VPB.n21 61.764
R76 VPB.n417 VPB.n416 61.764
R77 VPB.n88 VPB.n87 61.764
R78 VPB.n111 VPB.n110 61.764
R79 VPB.n257 VPB.n256 61.764
R80 VPB.n78 VPB.t34 55.106
R81 VPB.n481 VPB.t10 55.106
R82 VPB.n398 VPB.t21 55.106
R83 VPB.n167 VPB.t22 55.106
R84 VPB.n321 VPB.t13 55.106
R85 VPB.n238 VPB.t25 55.106
R86 VPB.n45 VPB.t20 55.106
R87 VPB.n442 VPB.t9 55.106
R88 VPB.n359 VPB.t11 55.106
R89 VPB.n134 VPB.t4 55.106
R90 VPB.n282 VPB.t18 55.106
R91 VPB.n202 VPB.t27 55.106
R92 VPB.n212 VPB.n211 48.952
R93 VPB.n295 VPB.n294 48.952
R94 VPB.n143 VPB.n142 48.952
R95 VPB.n372 VPB.n371 48.952
R96 VPB.n455 VPB.n454 48.952
R97 VPB.n54 VPB.n53 48.952
R98 VPB.n229 VPB.n228 44.502
R99 VPB.n312 VPB.n311 44.502
R100 VPB.n157 VPB.n156 44.502
R101 VPB.n389 VPB.n388 44.502
R102 VPB.n472 VPB.n471 44.502
R103 VPB.n68 VPB.n67 44.502
R104 VPB.n66 VPB.n14 40.824
R105 VPB.n57 VPB.n15 40.824
R106 VPB.n470 VPB.n469 40.824
R107 VPB.n453 VPB.n452 40.824
R108 VPB.n387 VPB.n386 40.824
R109 VPB.n370 VPB.n369 40.824
R110 VPB.n155 VPB.n103 40.824
R111 VPB.n146 VPB.n104 40.824
R112 VPB.n310 VPB.n309 40.824
R113 VPB.n293 VPB.n292 40.824
R114 VPB.n227 VPB.n226 40.824
R115 VPB.n210 VPB.n209 40.824
R116 VPB.n207 VPB.n206 35.118
R117 VPB.n510 VPB.n506 20.452
R118 VPB.n194 VPB.n191 20.452
R119 VPB.n217 VPB.n216 17.801
R120 VPB.n300 VPB.n299 17.801
R121 VPB.n148 VPB.n147 17.801
R122 VPB.n377 VPB.n376 17.801
R123 VPB.n460 VPB.n459 17.801
R124 VPB.n59 VPB.n58 17.801
R125 VPB.n14 VPB.t5 14.282
R126 VPB.n14 VPB.t35 14.282
R127 VPB.n15 VPB.t8 14.282
R128 VPB.n15 VPB.t3 14.282
R129 VPB.n469 VPB.t32 14.282
R130 VPB.n469 VPB.t23 14.282
R131 VPB.n452 VPB.t12 14.282
R132 VPB.n452 VPB.t31 14.282
R133 VPB.n386 VPB.t15 14.282
R134 VPB.n386 VPB.t24 14.282
R135 VPB.n369 VPB.t1 14.282
R136 VPB.n369 VPB.t14 14.282
R137 VPB.n103 VPB.t30 14.282
R138 VPB.n103 VPB.t28 14.282
R139 VPB.n104 VPB.t2 14.282
R140 VPB.n104 VPB.t33 14.282
R141 VPB.n309 VPB.t7 14.282
R142 VPB.n309 VPB.t19 14.282
R143 VPB.n292 VPB.t0 14.282
R144 VPB.n292 VPB.t6 14.282
R145 VPB.n226 VPB.t17 14.282
R146 VPB.n226 VPB.t26 14.282
R147 VPB.n209 VPB.t29 14.282
R148 VPB.n209 VPB.t16 14.282
R149 VPB.n194 VPB.n193 13.653
R150 VPB.n193 VPB.n192 13.653
R151 VPB.n205 VPB.n204 13.653
R152 VPB.n204 VPB.n203 13.653
R153 VPB.n201 VPB.n200 13.653
R154 VPB.n200 VPB.n199 13.653
R155 VPB.n197 VPB.n196 13.653
R156 VPB.n196 VPB.n195 13.653
R157 VPB.n214 VPB.n213 13.653
R158 VPB.n213 VPB.n212 13.653
R159 VPB.n219 VPB.n218 13.653
R160 VPB.n218 VPB.n217 13.653
R161 VPB.n224 VPB.n223 13.653
R162 VPB.n223 VPB.n222 13.653
R163 VPB.n231 VPB.n230 13.653
R164 VPB.n230 VPB.n229 13.653
R165 VPB.n236 VPB.n235 13.653
R166 VPB.n235 VPB.n234 13.653
R167 VPB.n241 VPB.n240 13.653
R168 VPB.n240 VPB.n239 13.653
R169 VPB.n245 VPB.n244 13.653
R170 VPB.n244 VPB.n243 13.653
R171 VPB.n249 VPB.n248 13.653
R172 VPB.n248 VPB.n247 13.653
R173 VPB.n276 VPB.n275 13.653
R174 VPB.n275 VPB.n274 13.653
R175 VPB.n280 VPB.n279 13.653
R176 VPB.n279 VPB.n278 13.653
R177 VPB.n285 VPB.n284 13.653
R178 VPB.n284 VPB.n283 13.653
R179 VPB.n290 VPB.n289 13.653
R180 VPB.n289 VPB.n288 13.653
R181 VPB.n297 VPB.n296 13.653
R182 VPB.n296 VPB.n295 13.653
R183 VPB.n302 VPB.n301 13.653
R184 VPB.n301 VPB.n300 13.653
R185 VPB.n307 VPB.n306 13.653
R186 VPB.n306 VPB.n305 13.653
R187 VPB.n314 VPB.n313 13.653
R188 VPB.n313 VPB.n312 13.653
R189 VPB.n319 VPB.n318 13.653
R190 VPB.n318 VPB.n317 13.653
R191 VPB.n324 VPB.n323 13.653
R192 VPB.n323 VPB.n322 13.653
R193 VPB.n328 VPB.n327 13.653
R194 VPB.n327 VPB.n326 13.653
R195 VPB.n332 VPB.n331 13.653
R196 VPB.n331 VPB.n330 13.653
R197 VPB.n130 VPB.n129 13.653
R198 VPB.n129 VPB.n128 13.653
R199 VPB.n133 VPB.n132 13.653
R200 VPB.n132 VPB.n131 13.653
R201 VPB.n137 VPB.n136 13.653
R202 VPB.n136 VPB.n135 13.653
R203 VPB.n141 VPB.n140 13.653
R204 VPB.n140 VPB.n139 13.653
R205 VPB.n145 VPB.n144 13.653
R206 VPB.n144 VPB.n143 13.653
R207 VPB.n150 VPB.n149 13.653
R208 VPB.n149 VPB.n148 13.653
R209 VPB.n154 VPB.n153 13.653
R210 VPB.n153 VPB.n152 13.653
R211 VPB.n159 VPB.n158 13.653
R212 VPB.n158 VPB.n157 13.653
R213 VPB.n163 VPB.n162 13.653
R214 VPB.n162 VPB.n161 13.653
R215 VPB.n166 VPB.n165 13.653
R216 VPB.n165 VPB.n164 13.653
R217 VPB.n170 VPB.n169 13.653
R218 VPB.n169 VPB.n168 13.653
R219 VPB.n348 VPB.n347 13.653
R220 VPB.n347 VPB.n346 13.653
R221 VPB.n353 VPB.n352 13.653
R222 VPB.n352 VPB.n351 13.653
R223 VPB.n357 VPB.n356 13.653
R224 VPB.n356 VPB.n355 13.653
R225 VPB.n362 VPB.n361 13.653
R226 VPB.n361 VPB.n360 13.653
R227 VPB.n367 VPB.n366 13.653
R228 VPB.n366 VPB.n365 13.653
R229 VPB.n374 VPB.n373 13.653
R230 VPB.n373 VPB.n372 13.653
R231 VPB.n379 VPB.n378 13.653
R232 VPB.n378 VPB.n377 13.653
R233 VPB.n384 VPB.n383 13.653
R234 VPB.n383 VPB.n382 13.653
R235 VPB.n391 VPB.n390 13.653
R236 VPB.n390 VPB.n389 13.653
R237 VPB.n396 VPB.n395 13.653
R238 VPB.n395 VPB.n394 13.653
R239 VPB.n401 VPB.n400 13.653
R240 VPB.n400 VPB.n399 13.653
R241 VPB.n405 VPB.n404 13.653
R242 VPB.n404 VPB.n403 13.653
R243 VPB.n409 VPB.n408 13.653
R244 VPB.n408 VPB.n407 13.653
R245 VPB.n436 VPB.n435 13.653
R246 VPB.n435 VPB.n434 13.653
R247 VPB.n440 VPB.n439 13.653
R248 VPB.n439 VPB.n438 13.653
R249 VPB.n445 VPB.n444 13.653
R250 VPB.n444 VPB.n443 13.653
R251 VPB.n450 VPB.n449 13.653
R252 VPB.n449 VPB.n448 13.653
R253 VPB.n457 VPB.n456 13.653
R254 VPB.n456 VPB.n455 13.653
R255 VPB.n462 VPB.n461 13.653
R256 VPB.n461 VPB.n460 13.653
R257 VPB.n467 VPB.n466 13.653
R258 VPB.n466 VPB.n465 13.653
R259 VPB.n474 VPB.n473 13.653
R260 VPB.n473 VPB.n472 13.653
R261 VPB.n479 VPB.n478 13.653
R262 VPB.n478 VPB.n477 13.653
R263 VPB.n484 VPB.n483 13.653
R264 VPB.n483 VPB.n482 13.653
R265 VPB.n488 VPB.n487 13.653
R266 VPB.n487 VPB.n486 13.653
R267 VPB.n492 VPB.n491 13.653
R268 VPB.n491 VPB.n490 13.653
R269 VPB.n41 VPB.n40 13.653
R270 VPB.n40 VPB.n39 13.653
R271 VPB.n44 VPB.n43 13.653
R272 VPB.n43 VPB.n42 13.653
R273 VPB.n48 VPB.n47 13.653
R274 VPB.n47 VPB.n46 13.653
R275 VPB.n52 VPB.n51 13.653
R276 VPB.n51 VPB.n50 13.653
R277 VPB.n56 VPB.n55 13.653
R278 VPB.n55 VPB.n54 13.653
R279 VPB.n61 VPB.n60 13.653
R280 VPB.n60 VPB.n59 13.653
R281 VPB.n65 VPB.n64 13.653
R282 VPB.n64 VPB.n63 13.653
R283 VPB.n70 VPB.n69 13.653
R284 VPB.n69 VPB.n68 13.653
R285 VPB.n74 VPB.n73 13.653
R286 VPB.n73 VPB.n72 13.653
R287 VPB.n77 VPB.n76 13.653
R288 VPB.n76 VPB.n75 13.653
R289 VPB.n81 VPB.n80 13.653
R290 VPB.n80 VPB.n79 13.653
R291 VPB.n506 VPB.n0 13.653
R292 VPB VPB.n0 13.653
R293 VPB.n222 VPB.n221 13.35
R294 VPB.n305 VPB.n304 13.35
R295 VPB.n152 VPB.n151 13.35
R296 VPB.n382 VPB.n381 13.35
R297 VPB.n465 VPB.n464 13.35
R298 VPB.n63 VPB.n62 13.35
R299 VPB.n510 VPB.n509 13.276
R300 VPB.n509 VPB.n507 13.276
R301 VPB.n36 VPB.n18 13.276
R302 VPB.n18 VPB.n16 13.276
R303 VPB.n431 VPB.n413 13.276
R304 VPB.n413 VPB.n411 13.276
R305 VPB.n102 VPB.n84 13.276
R306 VPB.n84 VPB.n82 13.276
R307 VPB.n125 VPB.n107 13.276
R308 VPB.n107 VPB.n105 13.276
R309 VPB.n271 VPB.n253 13.276
R310 VPB.n253 VPB.n251 13.276
R311 VPB.n201 VPB.n197 13.276
R312 VPB.n276 VPB.n272 13.276
R313 VPB.n130 VPB.n126 13.276
R314 VPB.n133 VPB.n130 13.276
R315 VPB.n141 VPB.n137 13.276
R316 VPB.n145 VPB.n141 13.276
R317 VPB.n154 VPB.n150 13.276
R318 VPB.n163 VPB.n159 13.276
R319 VPB.n166 VPB.n163 13.276
R320 VPB.n348 VPB.n170 13.276
R321 VPB.n349 VPB.n348 13.276
R322 VPB.n353 VPB.n349 13.276
R323 VPB.n436 VPB.n432 13.276
R324 VPB.n41 VPB.n37 13.276
R325 VPB.n44 VPB.n41 13.276
R326 VPB.n52 VPB.n48 13.276
R327 VPB.n56 VPB.n52 13.276
R328 VPB.n65 VPB.n61 13.276
R329 VPB.n74 VPB.n70 13.276
R330 VPB.n77 VPB.n74 13.276
R331 VPB.n506 VPB.n81 13.276
R332 VPB.n191 VPB.n173 13.276
R333 VPB.n173 VPB.n171 13.276
R334 VPB.n178 VPB.n176 12.796
R335 VPB.n178 VPB.n177 12.564
R336 VPB.n170 VPB.n167 12.558
R337 VPB.n81 VPB.n78 12.558
R338 VPB.n205 VPB.n202 12.2
R339 VPB.n134 VPB.n133 12.2
R340 VPB.n45 VPB.n44 12.2
R341 VPB.n186 VPB.n185 12.198
R342 VPB.n184 VPB.n183 12.198
R343 VPB.n181 VPB.n180 12.198
R344 VPB.n150 VPB.n146 9.329
R345 VPB.n61 VPB.n57 9.329
R346 VPB.n155 VPB.n154 8.97
R347 VPB.n66 VPB.n65 8.97
R348 VPB.n191 VPB.n190 7.5
R349 VPB.n176 VPB.n175 7.5
R350 VPB.n180 VPB.n179 7.5
R351 VPB.n183 VPB.n182 7.5
R352 VPB.n173 VPB.n172 7.5
R353 VPB.n188 VPB.n174 7.5
R354 VPB.n253 VPB.n252 7.5
R355 VPB.n266 VPB.n265 7.5
R356 VPB.n260 VPB.n259 7.5
R357 VPB.n262 VPB.n261 7.5
R358 VPB.n255 VPB.n254 7.5
R359 VPB.n271 VPB.n270 7.5
R360 VPB.n107 VPB.n106 7.5
R361 VPB.n120 VPB.n119 7.5
R362 VPB.n114 VPB.n113 7.5
R363 VPB.n116 VPB.n115 7.5
R364 VPB.n109 VPB.n108 7.5
R365 VPB.n125 VPB.n124 7.5
R366 VPB.n84 VPB.n83 7.5
R367 VPB.n97 VPB.n96 7.5
R368 VPB.n91 VPB.n90 7.5
R369 VPB.n93 VPB.n92 7.5
R370 VPB.n86 VPB.n85 7.5
R371 VPB.n102 VPB.n101 7.5
R372 VPB.n413 VPB.n412 7.5
R373 VPB.n426 VPB.n425 7.5
R374 VPB.n420 VPB.n419 7.5
R375 VPB.n422 VPB.n421 7.5
R376 VPB.n415 VPB.n414 7.5
R377 VPB.n431 VPB.n430 7.5
R378 VPB.n18 VPB.n17 7.5
R379 VPB.n31 VPB.n30 7.5
R380 VPB.n25 VPB.n24 7.5
R381 VPB.n27 VPB.n26 7.5
R382 VPB.n20 VPB.n19 7.5
R383 VPB.n36 VPB.n35 7.5
R384 VPB.n509 VPB.n508 7.5
R385 VPB.n12 VPB.n11 7.5
R386 VPB.n6 VPB.n5 7.5
R387 VPB.n8 VPB.n7 7.5
R388 VPB.n2 VPB.n1 7.5
R389 VPB.n511 VPB.n510 7.5
R390 VPB.n37 VPB.n36 7.176
R391 VPB.n432 VPB.n431 7.176
R392 VPB.n349 VPB.n102 7.176
R393 VPB.n126 VPB.n125 7.176
R394 VPB.n272 VPB.n271 7.176
R395 VPB.n267 VPB.n264 6.729
R396 VPB.n263 VPB.n260 6.729
R397 VPB.n258 VPB.n255 6.729
R398 VPB.n121 VPB.n118 6.729
R399 VPB.n117 VPB.n114 6.729
R400 VPB.n112 VPB.n109 6.729
R401 VPB.n98 VPB.n95 6.729
R402 VPB.n94 VPB.n91 6.729
R403 VPB.n89 VPB.n86 6.729
R404 VPB.n427 VPB.n424 6.729
R405 VPB.n423 VPB.n420 6.729
R406 VPB.n418 VPB.n415 6.729
R407 VPB.n32 VPB.n29 6.729
R408 VPB.n28 VPB.n25 6.729
R409 VPB.n23 VPB.n20 6.729
R410 VPB.n13 VPB.n10 6.729
R411 VPB.n9 VPB.n6 6.729
R412 VPB.n4 VPB.n2 6.729
R413 VPB.n258 VPB.n257 6.728
R414 VPB.n263 VPB.n262 6.728
R415 VPB.n267 VPB.n266 6.728
R416 VPB.n270 VPB.n269 6.728
R417 VPB.n112 VPB.n111 6.728
R418 VPB.n117 VPB.n116 6.728
R419 VPB.n121 VPB.n120 6.728
R420 VPB.n124 VPB.n123 6.728
R421 VPB.n89 VPB.n88 6.728
R422 VPB.n94 VPB.n93 6.728
R423 VPB.n98 VPB.n97 6.728
R424 VPB.n101 VPB.n100 6.728
R425 VPB.n418 VPB.n417 6.728
R426 VPB.n423 VPB.n422 6.728
R427 VPB.n427 VPB.n426 6.728
R428 VPB.n430 VPB.n429 6.728
R429 VPB.n23 VPB.n22 6.728
R430 VPB.n28 VPB.n27 6.728
R431 VPB.n32 VPB.n31 6.728
R432 VPB.n35 VPB.n34 6.728
R433 VPB.n4 VPB.n3 6.728
R434 VPB.n9 VPB.n8 6.728
R435 VPB.n13 VPB.n12 6.728
R436 VPB.n512 VPB.n511 6.728
R437 VPB.n190 VPB.n189 6.398
R438 VPB.n206 VPB.n194 6.112
R439 VPB.n206 VPB.n205 6.101
R440 VPB.n231 VPB.n227 4.305
R441 VPB.n314 VPB.n310 4.305
R442 VPB.n159 VPB.n155 4.305
R443 VPB.n391 VPB.n387 4.305
R444 VPB.n474 VPB.n470 4.305
R445 VPB.n70 VPB.n66 4.305
R446 VPB.n214 VPB.n210 3.947
R447 VPB.n297 VPB.n293 3.947
R448 VPB.n146 VPB.n145 3.947
R449 VPB.n374 VPB.n370 3.947
R450 VPB.n457 VPB.n453 3.947
R451 VPB.n57 VPB.n56 3.947
R452 VPB.n188 VPB.n181 1.402
R453 VPB.n188 VPB.n184 1.402
R454 VPB.n188 VPB.n186 1.402
R455 VPB.n188 VPB.n187 1.402
R456 VPB.n202 VPB.n201 1.076
R457 VPB.n285 VPB.n282 1.076
R458 VPB.n137 VPB.n134 1.076
R459 VPB.n362 VPB.n359 1.076
R460 VPB.n445 VPB.n442 1.076
R461 VPB.n48 VPB.n45 1.076
R462 VPB.n189 VPB.n188 0.735
R463 VPB.n188 VPB.n178 0.735
R464 VPB.n241 VPB.n238 0.717
R465 VPB.n324 VPB.n321 0.717
R466 VPB.n167 VPB.n166 0.717
R467 VPB.n401 VPB.n398 0.717
R468 VPB.n484 VPB.n481 0.717
R469 VPB.n78 VPB.n77 0.717
R470 VPB.n268 VPB.n267 0.387
R471 VPB.n268 VPB.n263 0.387
R472 VPB.n268 VPB.n258 0.387
R473 VPB.n269 VPB.n268 0.387
R474 VPB.n122 VPB.n121 0.387
R475 VPB.n122 VPB.n117 0.387
R476 VPB.n122 VPB.n112 0.387
R477 VPB.n123 VPB.n122 0.387
R478 VPB.n99 VPB.n98 0.387
R479 VPB.n99 VPB.n94 0.387
R480 VPB.n99 VPB.n89 0.387
R481 VPB.n100 VPB.n99 0.387
R482 VPB.n428 VPB.n427 0.387
R483 VPB.n428 VPB.n423 0.387
R484 VPB.n428 VPB.n418 0.387
R485 VPB.n429 VPB.n428 0.387
R486 VPB.n33 VPB.n32 0.387
R487 VPB.n33 VPB.n28 0.387
R488 VPB.n33 VPB.n23 0.387
R489 VPB.n34 VPB.n33 0.387
R490 VPB.n513 VPB.n13 0.387
R491 VPB.n513 VPB.n9 0.387
R492 VPB.n513 VPB.n4 0.387
R493 VPB.n513 VPB.n512 0.387
R494 VPB.n277 VPB.n250 0.272
R495 VPB.n334 VPB.n333 0.272
R496 VPB.n437 VPB.n410 0.272
R497 VPB.n494 VPB.n493 0.272
R498 VPB.n505 VPB 0.198
R499 VPB.n208 VPB.n207 0.136
R500 VPB.n215 VPB.n208 0.136
R501 VPB.n220 VPB.n215 0.136
R502 VPB.n225 VPB.n220 0.136
R503 VPB.n232 VPB.n225 0.136
R504 VPB.n237 VPB.n232 0.136
R505 VPB.n242 VPB.n237 0.136
R506 VPB.n246 VPB.n242 0.136
R507 VPB.n250 VPB.n246 0.136
R508 VPB.n281 VPB.n277 0.136
R509 VPB.n286 VPB.n281 0.136
R510 VPB.n291 VPB.n286 0.136
R511 VPB.n298 VPB.n291 0.136
R512 VPB.n303 VPB.n298 0.136
R513 VPB.n308 VPB.n303 0.136
R514 VPB.n315 VPB.n308 0.136
R515 VPB.n320 VPB.n315 0.136
R516 VPB.n325 VPB.n320 0.136
R517 VPB.n329 VPB.n325 0.136
R518 VPB.n333 VPB.n329 0.136
R519 VPB.n335 VPB.n334 0.136
R520 VPB.n336 VPB.n335 0.136
R521 VPB.n337 VPB.n336 0.136
R522 VPB.n338 VPB.n337 0.136
R523 VPB.n339 VPB.n338 0.136
R524 VPB.n340 VPB.n339 0.136
R525 VPB.n341 VPB.n340 0.136
R526 VPB.n342 VPB.n341 0.136
R527 VPB.n343 VPB.n342 0.136
R528 VPB.n344 VPB.n343 0.136
R529 VPB.n345 VPB.n344 0.136
R530 VPB.n345 VPB 0.136
R531 VPB.n354 VPB 0.136
R532 VPB.n358 VPB.n354 0.136
R533 VPB.n363 VPB.n358 0.136
R534 VPB.n368 VPB.n363 0.136
R535 VPB.n375 VPB.n368 0.136
R536 VPB.n380 VPB.n375 0.136
R537 VPB.n385 VPB.n380 0.136
R538 VPB.n392 VPB.n385 0.136
R539 VPB.n397 VPB.n392 0.136
R540 VPB.n402 VPB.n397 0.136
R541 VPB.n406 VPB.n402 0.136
R542 VPB.n410 VPB.n406 0.136
R543 VPB.n441 VPB.n437 0.136
R544 VPB.n446 VPB.n441 0.136
R545 VPB.n451 VPB.n446 0.136
R546 VPB.n458 VPB.n451 0.136
R547 VPB.n463 VPB.n458 0.136
R548 VPB.n468 VPB.n463 0.136
R549 VPB.n475 VPB.n468 0.136
R550 VPB.n480 VPB.n475 0.136
R551 VPB.n485 VPB.n480 0.136
R552 VPB.n489 VPB.n485 0.136
R553 VPB.n493 VPB.n489 0.136
R554 VPB.n495 VPB.n494 0.136
R555 VPB.n496 VPB.n495 0.136
R556 VPB.n497 VPB.n496 0.136
R557 VPB.n498 VPB.n497 0.136
R558 VPB.n499 VPB.n498 0.136
R559 VPB.n500 VPB.n499 0.136
R560 VPB.n501 VPB.n500 0.136
R561 VPB.n502 VPB.n501 0.136
R562 VPB.n503 VPB.n502 0.136
R563 VPB.n504 VPB.n503 0.136
R564 VPB.n505 VPB.n504 0.136
R565 a_4447_943.n5 a_4447_943.t8 454.685
R566 a_4447_943.n5 a_4447_943.t9 428.979
R567 a_4447_943.n6 a_4447_943.t7 248.006
R568 a_4447_943.n9 a_4447_943.n7 229.673
R569 a_4447_943.n7 a_4447_943.n6 156.035
R570 a_4447_943.n7 a_4447_943.n4 154.293
R571 a_4447_943.n6 a_4447_943.n5 81.941
R572 a_4447_943.n3 a_4447_943.n2 79.232
R573 a_4447_943.n4 a_4447_943.n3 63.152
R574 a_4447_943.n4 a_4447_943.n0 16.08
R575 a_4447_943.n3 a_4447_943.n1 16.08
R576 a_4447_943.n9 a_4447_943.n8 15.218
R577 a_4447_943.n0 a_4447_943.t5 14.282
R578 a_4447_943.n0 a_4447_943.t6 14.282
R579 a_4447_943.n1 a_4447_943.t0 14.282
R580 a_4447_943.n1 a_4447_943.t1 14.282
R581 a_4447_943.n2 a_4447_943.t3 14.282
R582 a_4447_943.n2 a_4447_943.t2 14.282
R583 a_4447_943.n10 a_4447_943.n9 12.014
R584 a_277_1004.n7 a_277_1004.t10 512.525
R585 a_277_1004.n5 a_277_1004.t7 512.525
R586 a_277_1004.n7 a_277_1004.t11 371.139
R587 a_277_1004.n5 a_277_1004.t12 371.139
R588 a_277_1004.n8 a_277_1004.t9 244.968
R589 a_277_1004.n6 a_277_1004.t8 244.968
R590 a_277_1004.n10 a_277_1004.n4 207.04
R591 a_277_1004.n8 a_277_1004.n7 198.954
R592 a_277_1004.n6 a_277_1004.n5 198.954
R593 a_277_1004.n12 a_277_1004.n10 176.926
R594 a_277_1004.n9 a_277_1004.n6 79.491
R595 a_277_1004.n3 a_277_1004.n2 79.232
R596 a_277_1004.n10 a_277_1004.n9 77.315
R597 a_277_1004.n9 a_277_1004.n8 76
R598 a_277_1004.n4 a_277_1004.n3 63.152
R599 a_277_1004.n4 a_277_1004.n0 16.08
R600 a_277_1004.n3 a_277_1004.n1 16.08
R601 a_277_1004.n12 a_277_1004.n11 15.218
R602 a_277_1004.n0 a_277_1004.t4 14.282
R603 a_277_1004.n0 a_277_1004.t2 14.282
R604 a_277_1004.n1 a_277_1004.t1 14.282
R605 a_277_1004.n1 a_277_1004.t0 14.282
R606 a_277_1004.n2 a_277_1004.t6 14.282
R607 a_277_1004.n2 a_277_1004.t5 14.282
R608 a_277_1004.n13 a_277_1004.n12 12.014
R609 a_599_943.n5 a_599_943.t12 512.525
R610 a_599_943.n7 a_599_943.t10 454.685
R611 a_599_943.n7 a_599_943.t8 428.979
R612 a_599_943.n5 a_599_943.t7 371.139
R613 a_599_943.n6 a_599_943.t9 297.715
R614 a_599_943.n8 a_599_943.t11 248.006
R615 a_599_943.n12 a_599_943.n10 229.673
R616 a_599_943.n10 a_599_943.n4 154.293
R617 a_599_943.n6 a_599_943.n5 146.207
R618 a_599_943.n9 a_599_943.n6 84.388
R619 a_599_943.n8 a_599_943.n7 81.941
R620 a_599_943.n9 a_599_943.n8 80.035
R621 a_599_943.n3 a_599_943.n2 79.232
R622 a_599_943.n10 a_599_943.n9 76
R623 a_599_943.n4 a_599_943.n3 63.152
R624 a_599_943.n4 a_599_943.n0 16.08
R625 a_599_943.n3 a_599_943.n1 16.08
R626 a_599_943.n12 a_599_943.n11 15.218
R627 a_599_943.n0 a_599_943.t2 14.282
R628 a_599_943.n0 a_599_943.t4 14.282
R629 a_599_943.n1 a_599_943.t5 14.282
R630 a_599_943.n1 a_599_943.t6 14.282
R631 a_599_943.n2 a_599_943.t1 14.282
R632 a_599_943.n2 a_599_943.t0 14.282
R633 a_599_943.n13 a_599_943.n12 12.014
R634 a_1561_943.n8 a_1561_943.t14 454.685
R635 a_1561_943.n10 a_1561_943.t8 454.685
R636 a_1561_943.n6 a_1561_943.t15 454.685
R637 a_1561_943.n8 a_1561_943.t11 428.979
R638 a_1561_943.n10 a_1561_943.t12 428.979
R639 a_1561_943.n6 a_1561_943.t13 428.979
R640 a_1561_943.n9 a_1561_943.t7 274.559
R641 a_1561_943.n7 a_1561_943.t10 274.559
R642 a_1561_943.n11 a_1561_943.t9 274.22
R643 a_1561_943.n16 a_1561_943.n14 249.704
R644 a_1561_943.n14 a_1561_943.n5 127.74
R645 a_1561_943.n13 a_1561_943.n7 82.484
R646 a_1561_943.n12 a_1561_943.n11 79.495
R647 a_1561_943.n4 a_1561_943.n3 79.232
R648 a_1561_943.n12 a_1561_943.n9 76
R649 a_1561_943.n14 a_1561_943.n13 76
R650 a_1561_943.n5 a_1561_943.n4 63.152
R651 a_1561_943.n9 a_1561_943.n8 55.388
R652 a_1561_943.n7 a_1561_943.n6 55.388
R653 a_1561_943.n11 a_1561_943.n10 55.049
R654 a_1561_943.n16 a_1561_943.n15 30
R655 a_1561_943.n17 a_1561_943.n0 24.383
R656 a_1561_943.n17 a_1561_943.n16 23.684
R657 a_1561_943.n5 a_1561_943.n1 16.08
R658 a_1561_943.n4 a_1561_943.n2 16.08
R659 a_1561_943.n1 a_1561_943.t2 14.282
R660 a_1561_943.n1 a_1561_943.t1 14.282
R661 a_1561_943.n2 a_1561_943.t6 14.282
R662 a_1561_943.n2 a_1561_943.t5 14.282
R663 a_1561_943.n3 a_1561_943.t4 14.282
R664 a_1561_943.n3 a_1561_943.t3 14.282
R665 a_1561_943.n13 a_1561_943.n12 4.035
R666 a_91_75.t0 a_91_75.n0 117.777
R667 a_91_75.n2 a_91_75.n1 55.228
R668 a_91_75.n4 a_91_75.n3 9.111
R669 a_91_75.n8 a_91_75.n6 7.859
R670 a_91_75.t0 a_91_75.n2 4.04
R671 a_91_75.t0 a_91_75.n8 3.034
R672 a_91_75.n6 a_91_75.n4 1.964
R673 a_91_75.n6 a_91_75.n5 1.964
R674 a_91_75.n8 a_91_75.n7 0.443
R675 a_372_182.n10 a_372_182.n8 82.852
R676 a_372_182.n11 a_372_182.n0 49.6
R677 a_372_182.n7 a_372_182.n6 32.833
R678 a_372_182.n8 a_372_182.t1 32.416
R679 a_372_182.n10 a_372_182.n9 27.2
R680 a_372_182.n3 a_372_182.n2 23.284
R681 a_372_182.n11 a_372_182.n10 22.4
R682 a_372_182.n7 a_372_182.n4 19.017
R683 a_372_182.n6 a_372_182.n5 13.494
R684 a_372_182.t1 a_372_182.n1 7.04
R685 a_372_182.t1 a_372_182.n3 5.727
R686 a_372_182.n8 a_372_182.n7 1.435
R687 a_2296_182.n12 a_2296_182.n10 82.852
R688 a_2296_182.t1 a_2296_182.n2 46.91
R689 a_2296_182.n7 a_2296_182.n5 34.805
R690 a_2296_182.n7 a_2296_182.n6 32.622
R691 a_2296_182.n10 a_2296_182.t1 32.416
R692 a_2296_182.n12 a_2296_182.n11 27.2
R693 a_2296_182.n13 a_2296_182.n0 23.498
R694 a_2296_182.n13 a_2296_182.n12 22.4
R695 a_2296_182.n9 a_2296_182.n7 19.017
R696 a_2296_182.n2 a_2296_182.n1 17.006
R697 a_2296_182.n5 a_2296_182.n4 7.5
R698 a_2296_182.n9 a_2296_182.n8 7.5
R699 a_2296_182.t1 a_2296_182.n3 7.04
R700 a_2296_182.n10 a_2296_182.n9 1.435
R701 a_2201_1004.n5 a_2201_1004.t9 512.525
R702 a_2201_1004.n5 a_2201_1004.t8 371.139
R703 a_2201_1004.n6 a_2201_1004.t7 244.609
R704 a_2201_1004.n7 a_2201_1004.n4 207.399
R705 a_2201_1004.n6 a_2201_1004.n5 199.313
R706 a_2201_1004.n9 a_2201_1004.n7 176.567
R707 a_2201_1004.n7 a_2201_1004.n6 153.315
R708 a_2201_1004.n3 a_2201_1004.n2 79.232
R709 a_2201_1004.n4 a_2201_1004.n3 63.152
R710 a_2201_1004.n4 a_2201_1004.n0 16.08
R711 a_2201_1004.n3 a_2201_1004.n1 16.08
R712 a_2201_1004.n9 a_2201_1004.n8 15.218
R713 a_2201_1004.n0 a_2201_1004.t5 14.282
R714 a_2201_1004.n0 a_2201_1004.t4 14.282
R715 a_2201_1004.n1 a_2201_1004.t3 14.282
R716 a_2201_1004.n1 a_2201_1004.t2 14.282
R717 a_2201_1004.n2 a_2201_1004.t1 14.282
R718 a_2201_1004.n2 a_2201_1004.t0 14.282
R719 a_2201_1004.n10 a_2201_1004.n9 12.014
R720 a_4220_182.n10 a_4220_182.n8 82.852
R721 a_4220_182.n7 a_4220_182.n6 32.833
R722 a_4220_182.n8 a_4220_182.t1 32.416
R723 a_4220_182.n10 a_4220_182.n9 27.2
R724 a_4220_182.n11 a_4220_182.n0 23.498
R725 a_4220_182.n3 a_4220_182.n2 23.284
R726 a_4220_182.n11 a_4220_182.n10 22.4
R727 a_4220_182.n7 a_4220_182.n4 19.017
R728 a_4220_182.n6 a_4220_182.n5 13.494
R729 a_4220_182.t1 a_4220_182.n1 7.04
R730 a_4220_182.t1 a_4220_182.n3 5.727
R731 a_4220_182.n8 a_4220_182.n7 1.435
R732 a_1334_182.n9 a_1334_182.n7 82.852
R733 a_1334_182.n3 a_1334_182.n1 44.628
R734 a_1334_182.t0 a_1334_182.n9 32.417
R735 a_1334_182.n7 a_1334_182.n6 27.2
R736 a_1334_182.n5 a_1334_182.n4 23.498
R737 a_1334_182.n3 a_1334_182.n2 23.284
R738 a_1334_182.n7 a_1334_182.n5 22.4
R739 a_1334_182.t0 a_1334_182.n11 20.241
R740 a_1334_182.n11 a_1334_182.n10 13.494
R741 a_1334_182.t0 a_1334_182.n0 8.137
R742 a_1334_182.t0 a_1334_182.n3 5.727
R743 a_1334_182.n9 a_1334_182.n8 1.435
R744 a_2015_75.t0 a_2015_75.n3 117.777
R745 a_2015_75.n6 a_2015_75.n5 45.444
R746 a_2015_75.t0 a_2015_75.n6 21.213
R747 a_2015_75.t0 a_2015_75.n4 11.595
R748 a_2015_75.n2 a_2015_75.n1 2.455
R749 a_2015_75.n2 a_2015_75.n0 1.32
R750 a_2015_75.t0 a_2015_75.n2 0.246
R751 VNB.n159 VNB.n158 199.897
R752 VNB.n30 VNB.n29 199.897
R753 VNB.n10 VNB.n9 199.897
R754 VNB.n299 VNB.n298 199.897
R755 VNB.n374 VNB.n373 199.897
R756 VNB.n39 VNB.n37 154.509
R757 VNB.n168 VNB.n166 154.509
R758 VNB.n308 VNB.n306 154.509
R759 VNB.n240 VNB.n238 154.509
R760 VNB.n383 VNB.n381 154.509
R761 VNB.n125 VNB.n124 147.75
R762 VNB.n200 VNB.n199 147.75
R763 VNB.n63 VNB.n62 147.75
R764 VNB.n340 VNB.n339 147.75
R765 VNB.n132 VNB.n129 121.366
R766 VNB.n207 VNB.n204 121.366
R767 VNB.n68 VNB.n66 121.366
R768 VNB.n347 VNB.n344 121.366
R769 VNB.n278 VNB.n277 85.559
R770 VNB.n421 VNB.n420 85.559
R771 VNB.n447 VNB.n446 76
R772 VNB.n111 VNB.n110 76
R773 VNB.n115 VNB.n114 76
R774 VNB.n119 VNB.n118 76
R775 VNB.n123 VNB.n122 76
R776 VNB.n128 VNB.n127 76
R777 VNB.n140 VNB.n139 76
R778 VNB.n144 VNB.n143 76
R779 VNB.n148 VNB.n147 76
R780 VNB.n170 VNB.n169 76
R781 VNB.n174 VNB.n173 76
R782 VNB.n178 VNB.n177 76
R783 VNB.n182 VNB.n181 76
R784 VNB.n186 VNB.n185 76
R785 VNB.n190 VNB.n189 76
R786 VNB.n194 VNB.n193 76
R787 VNB.n198 VNB.n197 76
R788 VNB.n203 VNB.n202 76
R789 VNB.n215 VNB.n214 76
R790 VNB.n219 VNB.n218 76
R791 VNB.n223 VNB.n222 76
R792 VNB.n236 VNB.n235 76
R793 VNB.n242 VNB.n241 76
R794 VNB.n246 VNB.n245 76
R795 VNB.n250 VNB.n249 76
R796 VNB.n254 VNB.n253 76
R797 VNB.n258 VNB.n257 76
R798 VNB.n262 VNB.n261 76
R799 VNB.n266 VNB.n265 76
R800 VNB.n270 VNB.n269 76
R801 VNB.n274 VNB.n273 76
R802 VNB.n280 VNB.n279 76
R803 VNB.n284 VNB.n283 76
R804 VNB.n288 VNB.n287 76
R805 VNB.n310 VNB.n309 76
R806 VNB.n314 VNB.n313 76
R807 VNB.n318 VNB.n317 76
R808 VNB.n322 VNB.n321 76
R809 VNB.n326 VNB.n325 76
R810 VNB.n330 VNB.n329 76
R811 VNB.n334 VNB.n333 76
R812 VNB.n338 VNB.n337 76
R813 VNB.n343 VNB.n342 76
R814 VNB.n355 VNB.n354 76
R815 VNB.n359 VNB.n358 76
R816 VNB.n363 VNB.n362 76
R817 VNB.n385 VNB.n384 76
R818 VNB.n389 VNB.n388 76
R819 VNB.n393 VNB.n392 76
R820 VNB.n397 VNB.n396 76
R821 VNB.n401 VNB.n400 76
R822 VNB.n405 VNB.n404 76
R823 VNB.n409 VNB.n408 76
R824 VNB.n413 VNB.n412 76
R825 VNB.n417 VNB.n416 76
R826 VNB.n423 VNB.n422 76
R827 VNB.n427 VNB.n426 76
R828 VNB.n73 VNB.n72 73.875
R829 VNB.n138 VNB.n137 64.552
R830 VNB.n213 VNB.n212 64.552
R831 VNB.n71 VNB.n19 64.552
R832 VNB.n353 VNB.n352 64.552
R833 VNB.n276 VNB.n275 41.971
R834 VNB.n419 VNB.n418 41.971
R835 VNB.n132 VNB.n131 36.937
R836 VNB.n207 VNB.n206 36.937
R837 VNB.n68 VNB.n67 36.937
R838 VNB.n347 VNB.n346 36.937
R839 VNB.n106 VNB.n105 35.118
R840 VNB.n131 VNB.n130 29.844
R841 VNB.n206 VNB.n205 29.844
R842 VNB.n346 VNB.n345 29.844
R843 VNB.n137 VNB.n136 28.421
R844 VNB.n212 VNB.n211 28.421
R845 VNB.n19 VNB.n18 28.421
R846 VNB.n352 VNB.n351 28.421
R847 VNB.n137 VNB.n135 25.263
R848 VNB.n212 VNB.n210 25.263
R849 VNB.n19 VNB.n17 25.263
R850 VNB.n352 VNB.n350 25.263
R851 VNB.n135 VNB.n134 24.383
R852 VNB.n210 VNB.n209 24.383
R853 VNB.n17 VNB.n16 24.383
R854 VNB.n350 VNB.n349 24.383
R855 VNB.n95 VNB.n92 20.452
R856 VNB.n446 VNB.n443 20.452
R857 VNB.n446 VNB.n445 13.653
R858 VNB.n445 VNB.n444 13.653
R859 VNB.n426 VNB.n425 13.653
R860 VNB.n425 VNB.n424 13.653
R861 VNB.n422 VNB.n419 13.653
R862 VNB.n416 VNB.n415 13.653
R863 VNB.n415 VNB.n414 13.653
R864 VNB.n412 VNB.n411 13.653
R865 VNB.n411 VNB.n410 13.653
R866 VNB.n408 VNB.n407 13.653
R867 VNB.n407 VNB.n406 13.653
R868 VNB.n404 VNB.n403 13.653
R869 VNB.n403 VNB.n402 13.653
R870 VNB.n400 VNB.n399 13.653
R871 VNB.n399 VNB.n398 13.653
R872 VNB.n396 VNB.n395 13.653
R873 VNB.n395 VNB.n394 13.653
R874 VNB.n392 VNB.n391 13.653
R875 VNB.n391 VNB.n390 13.653
R876 VNB.n388 VNB.n387 13.653
R877 VNB.n387 VNB.n386 13.653
R878 VNB.n384 VNB.n383 13.653
R879 VNB.n383 VNB.n382 13.653
R880 VNB.n362 VNB.n361 13.653
R881 VNB.n361 VNB.n360 13.653
R882 VNB.n358 VNB.n357 13.653
R883 VNB.n357 VNB.n356 13.653
R884 VNB.n354 VNB.n348 13.653
R885 VNB.n348 VNB.n347 13.653
R886 VNB.n342 VNB.n341 13.653
R887 VNB.n341 VNB.n340 13.653
R888 VNB.n337 VNB.n336 13.653
R889 VNB.n336 VNB.n335 13.653
R890 VNB.n333 VNB.n332 13.653
R891 VNB.n332 VNB.n331 13.653
R892 VNB.n329 VNB.n328 13.653
R893 VNB.n328 VNB.n327 13.653
R894 VNB.n325 VNB.n324 13.653
R895 VNB.n324 VNB.n323 13.653
R896 VNB.n321 VNB.n320 13.653
R897 VNB.n320 VNB.n319 13.653
R898 VNB.n317 VNB.n316 13.653
R899 VNB.n316 VNB.n315 13.653
R900 VNB.n313 VNB.n312 13.653
R901 VNB.n312 VNB.n311 13.653
R902 VNB.n309 VNB.n308 13.653
R903 VNB.n308 VNB.n307 13.653
R904 VNB.n287 VNB.n286 13.653
R905 VNB.n286 VNB.n285 13.653
R906 VNB.n283 VNB.n282 13.653
R907 VNB.n282 VNB.n281 13.653
R908 VNB.n279 VNB.n276 13.653
R909 VNB.n273 VNB.n272 13.653
R910 VNB.n272 VNB.n271 13.653
R911 VNB.n269 VNB.n268 13.653
R912 VNB.n268 VNB.n267 13.653
R913 VNB.n265 VNB.n264 13.653
R914 VNB.n264 VNB.n263 13.653
R915 VNB.n261 VNB.n260 13.653
R916 VNB.n260 VNB.n259 13.653
R917 VNB.n257 VNB.n256 13.653
R918 VNB.n256 VNB.n255 13.653
R919 VNB.n253 VNB.n252 13.653
R920 VNB.n252 VNB.n251 13.653
R921 VNB.n249 VNB.n248 13.653
R922 VNB.n248 VNB.n247 13.653
R923 VNB.n245 VNB.n244 13.653
R924 VNB.n244 VNB.n243 13.653
R925 VNB.n241 VNB.n240 13.653
R926 VNB.n240 VNB.n239 13.653
R927 VNB.n236 VNB.n77 13.653
R928 VNB.n77 VNB.n76 13.653
R929 VNB.n75 VNB.n74 13.653
R930 VNB.n74 VNB.n73 13.653
R931 VNB.n70 VNB.n69 13.653
R932 VNB.n69 VNB.n68 13.653
R933 VNB.n65 VNB.n64 13.653
R934 VNB.n64 VNB.n63 13.653
R935 VNB.n61 VNB.n60 13.653
R936 VNB.n60 VNB.n59 13.653
R937 VNB.n58 VNB.n57 13.653
R938 VNB.n57 VNB.n56 13.653
R939 VNB.n55 VNB.n54 13.653
R940 VNB.n54 VNB.n53 13.653
R941 VNB.n52 VNB.n51 13.653
R942 VNB.n51 VNB.n50 13.653
R943 VNB.n49 VNB.n48 13.653
R944 VNB.n48 VNB.n47 13.653
R945 VNB.n46 VNB.n45 13.653
R946 VNB.n45 VNB.n44 13.653
R947 VNB.n43 VNB.n42 13.653
R948 VNB.n42 VNB.n41 13.653
R949 VNB.n40 VNB.n39 13.653
R950 VNB.n39 VNB.n38 13.653
R951 VNB.n222 VNB.n221 13.653
R952 VNB.n221 VNB.n220 13.653
R953 VNB.n218 VNB.n217 13.653
R954 VNB.n217 VNB.n216 13.653
R955 VNB.n214 VNB.n208 13.653
R956 VNB.n208 VNB.n207 13.653
R957 VNB.n202 VNB.n201 13.653
R958 VNB.n201 VNB.n200 13.653
R959 VNB.n197 VNB.n196 13.653
R960 VNB.n196 VNB.n195 13.653
R961 VNB.n193 VNB.n192 13.653
R962 VNB.n192 VNB.n191 13.653
R963 VNB.n189 VNB.n188 13.653
R964 VNB.n188 VNB.n187 13.653
R965 VNB.n185 VNB.n184 13.653
R966 VNB.n184 VNB.n183 13.653
R967 VNB.n181 VNB.n180 13.653
R968 VNB.n180 VNB.n179 13.653
R969 VNB.n177 VNB.n176 13.653
R970 VNB.n176 VNB.n175 13.653
R971 VNB.n173 VNB.n172 13.653
R972 VNB.n172 VNB.n171 13.653
R973 VNB.n169 VNB.n168 13.653
R974 VNB.n168 VNB.n167 13.653
R975 VNB.n147 VNB.n146 13.653
R976 VNB.n146 VNB.n145 13.653
R977 VNB.n143 VNB.n142 13.653
R978 VNB.n142 VNB.n141 13.653
R979 VNB.n139 VNB.n133 13.653
R980 VNB.n133 VNB.n132 13.653
R981 VNB.n127 VNB.n126 13.653
R982 VNB.n126 VNB.n125 13.653
R983 VNB.n122 VNB.n121 13.653
R984 VNB.n121 VNB.n120 13.653
R985 VNB.n118 VNB.n117 13.653
R986 VNB.n117 VNB.n116 13.653
R987 VNB.n114 VNB.n113 13.653
R988 VNB.n113 VNB.n112 13.653
R989 VNB.n110 VNB.n109 13.653
R990 VNB.n109 VNB.n108 13.653
R991 VNB.n102 VNB.n101 13.653
R992 VNB.n101 VNB.n100 13.653
R993 VNB.n103 VNB.n99 13.653
R994 VNB.n99 VNB.n98 13.653
R995 VNB.n104 VNB.n97 13.653
R996 VNB.n97 VNB.n96 13.653
R997 VNB.n95 VNB.n94 13.653
R998 VNB.n94 VNB.n93 13.653
R999 VNB.n435 VNB.n432 13.577
R1000 VNB.n366 VNB.n364 13.276
R1001 VNB.n379 VNB.n366 13.276
R1002 VNB.n291 VNB.n289 13.276
R1003 VNB.n304 VNB.n291 13.276
R1004 VNB.n2 VNB.n0 13.276
R1005 VNB.n15 VNB.n2 13.276
R1006 VNB.n22 VNB.n20 13.276
R1007 VNB.n35 VNB.n22 13.276
R1008 VNB.n151 VNB.n149 13.276
R1009 VNB.n164 VNB.n151 13.276
R1010 VNB.n80 VNB.n78 13.276
R1011 VNB.n92 VNB.n80 13.276
R1012 VNB.n430 VNB.n428 13.276
R1013 VNB.n443 VNB.n430 13.276
R1014 VNB.n104 VNB.n103 13.276
R1015 VNB.n103 VNB.n102 13.276
R1016 VNB.n169 VNB.n165 13.276
R1017 VNB.n40 VNB.n36 13.276
R1018 VNB.n43 VNB.n40 13.276
R1019 VNB.n46 VNB.n43 13.276
R1020 VNB.n49 VNB.n46 13.276
R1021 VNB.n52 VNB.n49 13.276
R1022 VNB.n55 VNB.n52 13.276
R1023 VNB.n58 VNB.n55 13.276
R1024 VNB.n61 VNB.n58 13.276
R1025 VNB.n65 VNB.n61 13.276
R1026 VNB.n70 VNB.n65 13.276
R1027 VNB.n236 VNB.n75 13.276
R1028 VNB.n237 VNB.n236 13.276
R1029 VNB.n241 VNB.n237 13.276
R1030 VNB.n309 VNB.n305 13.276
R1031 VNB.n384 VNB.n380 13.276
R1032 VNB.n75 VNB.n71 12.02
R1033 VNB.n92 VNB.n91 7.5
R1034 VNB.n83 VNB.n82 7.5
R1035 VNB.n86 VNB.n85 7.5
R1036 VNB.n80 VNB.n79 7.5
R1037 VNB.n164 VNB.n163 7.5
R1038 VNB.n157 VNB.n156 7.5
R1039 VNB.n153 VNB.n152 7.5
R1040 VNB.n151 VNB.n150 7.5
R1041 VNB.n35 VNB.n34 7.5
R1042 VNB.n28 VNB.n27 7.5
R1043 VNB.n24 VNB.n23 7.5
R1044 VNB.n22 VNB.n21 7.5
R1045 VNB.n15 VNB.n14 7.5
R1046 VNB.n8 VNB.n7 7.5
R1047 VNB.n4 VNB.n3 7.5
R1048 VNB.n2 VNB.n1 7.5
R1049 VNB.n304 VNB.n303 7.5
R1050 VNB.n297 VNB.n296 7.5
R1051 VNB.n293 VNB.n292 7.5
R1052 VNB.n291 VNB.n290 7.5
R1053 VNB.n379 VNB.n378 7.5
R1054 VNB.n372 VNB.n371 7.5
R1055 VNB.n368 VNB.n367 7.5
R1056 VNB.n366 VNB.n365 7.5
R1057 VNB.n437 VNB.n436 7.5
R1058 VNB.n443 VNB.n442 7.5
R1059 VNB.n430 VNB.n429 7.5
R1060 VNB.n434 VNB.n433 7.5
R1061 VNB.n380 VNB.n379 7.176
R1062 VNB.n305 VNB.n304 7.176
R1063 VNB.n237 VNB.n15 7.176
R1064 VNB.n36 VNB.n35 7.176
R1065 VNB.n165 VNB.n164 7.176
R1066 VNB.n160 VNB.n157 7.011
R1067 VNB.n155 VNB.n153 7.011
R1068 VNB.n31 VNB.n28 7.011
R1069 VNB.n26 VNB.n24 7.011
R1070 VNB.n11 VNB.n8 7.011
R1071 VNB.n6 VNB.n4 7.011
R1072 VNB.n300 VNB.n297 7.011
R1073 VNB.n295 VNB.n293 7.011
R1074 VNB.n375 VNB.n372 7.011
R1075 VNB.n370 VNB.n368 7.011
R1076 VNB.n439 VNB.n437 7.011
R1077 VNB.n163 VNB.n162 7.01
R1078 VNB.n155 VNB.n154 7.01
R1079 VNB.n160 VNB.n159 7.01
R1080 VNB.n34 VNB.n33 7.01
R1081 VNB.n26 VNB.n25 7.01
R1082 VNB.n31 VNB.n30 7.01
R1083 VNB.n14 VNB.n13 7.01
R1084 VNB.n6 VNB.n5 7.01
R1085 VNB.n11 VNB.n10 7.01
R1086 VNB.n303 VNB.n302 7.01
R1087 VNB.n295 VNB.n294 7.01
R1088 VNB.n300 VNB.n299 7.01
R1089 VNB.n378 VNB.n377 7.01
R1090 VNB.n370 VNB.n369 7.01
R1091 VNB.n375 VNB.n374 7.01
R1092 VNB.n439 VNB.n438 7.01
R1093 VNB.n84 VNB.n81 7.01
R1094 VNB.n88 VNB.n86 7.01
R1095 VNB.n91 VNB.n90 7.01
R1096 VNB.n88 VNB.n87 7.01
R1097 VNB.n84 VNB.n83 7.01
R1098 VNB.n435 VNB.n434 6.788
R1099 VNB.n442 VNB.n441 6.788
R1100 VNB.n105 VNB.n95 6.111
R1101 VNB.n105 VNB.n104 6.1
R1102 VNB.n139 VNB.n138 1.255
R1103 VNB.n214 VNB.n213 1.255
R1104 VNB.n71 VNB.n70 1.255
R1105 VNB.n279 VNB.n278 1.255
R1106 VNB.n354 VNB.n353 1.255
R1107 VNB.n422 VNB.n421 1.255
R1108 VNB.n440 VNB.n431 0.921
R1109 VNB.n440 VNB.n435 0.476
R1110 VNB.n441 VNB.n440 0.475
R1111 VNB.n170 VNB.n148 0.272
R1112 VNB.n224 VNB.n223 0.272
R1113 VNB.n310 VNB.n288 0.272
R1114 VNB.n385 VNB.n363 0.272
R1115 VNB.n161 VNB.n155 0.246
R1116 VNB.n162 VNB.n161 0.246
R1117 VNB.n161 VNB.n160 0.246
R1118 VNB.n32 VNB.n26 0.246
R1119 VNB.n33 VNB.n32 0.246
R1120 VNB.n32 VNB.n31 0.246
R1121 VNB.n12 VNB.n6 0.246
R1122 VNB.n13 VNB.n12 0.246
R1123 VNB.n12 VNB.n11 0.246
R1124 VNB.n301 VNB.n295 0.246
R1125 VNB.n302 VNB.n301 0.246
R1126 VNB.n301 VNB.n300 0.246
R1127 VNB.n376 VNB.n370 0.246
R1128 VNB.n377 VNB.n376 0.246
R1129 VNB.n376 VNB.n375 0.246
R1130 VNB.n440 VNB.n439 0.246
R1131 VNB.n90 VNB.n89 0.246
R1132 VNB.n89 VNB.n88 0.246
R1133 VNB.n89 VNB.n84 0.246
R1134 VNB.n107 VNB.n106 0.136
R1135 VNB.n111 VNB.n107 0.136
R1136 VNB.n115 VNB.n111 0.136
R1137 VNB.n119 VNB.n115 0.136
R1138 VNB.n123 VNB.n119 0.136
R1139 VNB.n128 VNB.n123 0.136
R1140 VNB.n140 VNB.n128 0.136
R1141 VNB.n144 VNB.n140 0.136
R1142 VNB.n148 VNB.n144 0.136
R1143 VNB.n174 VNB.n170 0.136
R1144 VNB.n178 VNB.n174 0.136
R1145 VNB.n182 VNB.n178 0.136
R1146 VNB.n186 VNB.n182 0.136
R1147 VNB.n190 VNB.n186 0.136
R1148 VNB.n194 VNB.n190 0.136
R1149 VNB.n198 VNB.n194 0.136
R1150 VNB.n203 VNB.n198 0.136
R1151 VNB.n215 VNB.n203 0.136
R1152 VNB.n219 VNB.n215 0.136
R1153 VNB.n223 VNB.n219 0.136
R1154 VNB.n225 VNB.n224 0.136
R1155 VNB.n226 VNB.n225 0.136
R1156 VNB.n227 VNB.n226 0.136
R1157 VNB.n228 VNB.n227 0.136
R1158 VNB.n229 VNB.n228 0.136
R1159 VNB.n230 VNB.n229 0.136
R1160 VNB.n231 VNB.n230 0.136
R1161 VNB.n232 VNB.n231 0.136
R1162 VNB.n233 VNB.n232 0.136
R1163 VNB.n234 VNB.n233 0.136
R1164 VNB.n235 VNB.n234 0.136
R1165 VNB.n235 VNB 0.136
R1166 VNB.n242 VNB 0.136
R1167 VNB.n246 VNB.n242 0.136
R1168 VNB.n250 VNB.n246 0.136
R1169 VNB.n254 VNB.n250 0.136
R1170 VNB.n258 VNB.n254 0.136
R1171 VNB.n262 VNB.n258 0.136
R1172 VNB.n266 VNB.n262 0.136
R1173 VNB.n270 VNB.n266 0.136
R1174 VNB.n274 VNB.n270 0.136
R1175 VNB.n280 VNB.n274 0.136
R1176 VNB.n284 VNB.n280 0.136
R1177 VNB.n288 VNB.n284 0.136
R1178 VNB.n314 VNB.n310 0.136
R1179 VNB.n318 VNB.n314 0.136
R1180 VNB.n322 VNB.n318 0.136
R1181 VNB.n326 VNB.n322 0.136
R1182 VNB.n330 VNB.n326 0.136
R1183 VNB.n334 VNB.n330 0.136
R1184 VNB.n338 VNB.n334 0.136
R1185 VNB.n343 VNB.n338 0.136
R1186 VNB.n355 VNB.n343 0.136
R1187 VNB.n359 VNB.n355 0.136
R1188 VNB.n363 VNB.n359 0.136
R1189 VNB.n389 VNB.n385 0.136
R1190 VNB.n393 VNB.n389 0.136
R1191 VNB.n397 VNB.n393 0.136
R1192 VNB.n401 VNB.n397 0.136
R1193 VNB.n405 VNB.n401 0.136
R1194 VNB.n409 VNB.n405 0.136
R1195 VNB.n413 VNB.n409 0.136
R1196 VNB.n417 VNB.n413 0.136
R1197 VNB.n423 VNB.n417 0.136
R1198 VNB.n427 VNB.n423 0.136
R1199 VNB.n447 VNB.n427 0.136
R1200 VNB.n447 VNB 0.031
R1201 a_3258_182.n9 a_3258_182.n7 82.852
R1202 a_3258_182.n3 a_3258_182.n1 44.628
R1203 a_3258_182.t0 a_3258_182.n9 32.417
R1204 a_3258_182.n7 a_3258_182.n6 27.2
R1205 a_3258_182.n5 a_3258_182.n4 23.498
R1206 a_3258_182.n3 a_3258_182.n2 23.284
R1207 a_3258_182.n7 a_3258_182.n5 22.4
R1208 a_3258_182.t0 a_3258_182.n11 20.241
R1209 a_3258_182.n11 a_3258_182.n10 13.494
R1210 a_3258_182.t0 a_3258_182.n0 8.137
R1211 a_3258_182.t0 a_3258_182.n3 5.727
R1212 a_3258_182.n9 a_3258_182.n8 1.435
R1213 a_5182_182.n10 a_5182_182.n8 82.852
R1214 a_5182_182.n7 a_5182_182.n6 32.833
R1215 a_5182_182.n8 a_5182_182.t1 32.416
R1216 a_5182_182.n10 a_5182_182.n9 27.2
R1217 a_5182_182.n11 a_5182_182.n0 23.498
R1218 a_5182_182.n3 a_5182_182.n2 23.284
R1219 a_5182_182.n11 a_5182_182.n10 22.4
R1220 a_5182_182.n7 a_5182_182.n4 19.017
R1221 a_5182_182.n6 a_5182_182.n5 13.494
R1222 a_5182_182.t1 a_5182_182.n1 7.04
R1223 a_5182_182.t1 a_5182_182.n3 5.727
R1224 a_5182_182.n8 a_5182_182.n7 1.435
R1225 a_2977_75.n5 a_2977_75.n4 19.724
R1226 a_2977_75.t0 a_2977_75.n3 11.595
R1227 a_2977_75.t0 a_2977_75.n5 9.207
R1228 a_2977_75.n2 a_2977_75.n1 2.455
R1229 a_2977_75.n2 a_2977_75.n0 1.32
R1230 a_2977_75.t0 a_2977_75.n2 0.246
R1231 a_1053_75.n5 a_1053_75.n4 19.724
R1232 a_1053_75.t0 a_1053_75.n3 11.595
R1233 a_1053_75.t0 a_1053_75.n5 9.207
R1234 a_1053_75.n2 a_1053_75.n1 2.455
R1235 a_1053_75.n2 a_1053_75.n0 1.32
R1236 a_1053_75.t0 a_1053_75.n2 0.246
R1237 a_3939_75.n1 a_3939_75.n0 25.576
R1238 a_3939_75.n3 a_3939_75.n2 9.111
R1239 a_3939_75.n7 a_3939_75.n6 2.455
R1240 a_3939_75.n5 a_3939_75.n3 1.964
R1241 a_3939_75.n5 a_3939_75.n4 1.964
R1242 a_3939_75.t0 a_3939_75.n1 1.871
R1243 a_3939_75.n7 a_3939_75.n5 0.636
R1244 a_3939_75.t0 a_3939_75.n7 0.246
R1245 a_4901_75.n1 a_4901_75.n0 25.576
R1246 a_4901_75.n3 a_4901_75.n2 9.111
R1247 a_4901_75.n7 a_4901_75.n6 2.455
R1248 a_4901_75.n5 a_4901_75.n3 1.964
R1249 a_4901_75.n5 a_4901_75.n4 1.964
R1250 a_4901_75.t0 a_4901_75.n1 1.871
R1251 a_4901_75.n7 a_4901_75.n5 0.636
R1252 a_4901_75.t0 a_4901_75.n7 0.246














































































































































































































































































































































































































































































































































































































































































































.ends
