magic
tech sky130A
magscale 1 2
timestamp 1648061063
<< nwell >>
rect 52 -436 352 36
<< pmos >>
rect 144 -400 174 0
rect 232 -400 262 0
<< pdiff >>
rect 88 -38 144 0
rect 88 -72 98 -38
rect 132 -72 144 -38
rect 88 -106 144 -72
rect 88 -140 98 -106
rect 132 -140 144 -106
rect 88 -174 144 -140
rect 88 -208 98 -174
rect 132 -208 144 -174
rect 88 -242 144 -208
rect 88 -276 98 -242
rect 132 -276 144 -242
rect 88 -400 144 -276
rect 174 -38 232 0
rect 174 -72 186 -38
rect 220 -72 232 -38
rect 174 -106 232 -72
rect 174 -140 186 -106
rect 220 -140 232 -106
rect 174 -174 232 -140
rect 174 -208 186 -174
rect 220 -208 232 -174
rect 174 -242 232 -208
rect 174 -276 186 -242
rect 220 -276 232 -242
rect 174 -400 232 -276
rect 262 -38 316 0
rect 262 -72 274 -38
rect 308 -72 316 -38
rect 262 -106 316 -72
rect 262 -140 274 -106
rect 308 -140 316 -106
rect 262 -174 316 -140
rect 262 -208 274 -174
rect 308 -208 316 -174
rect 262 -242 316 -208
rect 262 -276 274 -242
rect 308 -276 316 -242
rect 262 -400 316 -276
<< pdiffc >>
rect 98 -72 132 -38
rect 98 -140 132 -106
rect 98 -208 132 -174
rect 98 -276 132 -242
rect 186 -72 220 -38
rect 186 -140 220 -106
rect 186 -208 220 -174
rect 186 -276 220 -242
rect 274 -72 308 -38
rect 274 -140 308 -106
rect 274 -208 308 -174
rect 274 -276 308 -242
<< poly >>
rect 144 0 174 26
rect 232 0 262 26
rect 144 -431 174 -400
rect 232 -431 262 -400
rect 144 -461 262 -431
<< locali >>
rect 98 -38 132 42
rect 98 -106 132 -72
rect 98 -174 132 -140
rect 98 -242 132 -208
rect 98 -293 132 -276
rect 186 -38 220 0
rect 186 -106 220 -72
rect 186 -174 220 -140
rect 186 -242 220 -208
rect 186 -293 220 -276
rect 274 -38 308 42
rect 274 -106 308 -72
rect 274 -174 308 -140
rect 274 -242 308 -208
rect 274 -293 308 -276
<< end >>
