* SPICE3 file created from TMRDFFSNQNX1.ext - technology: sky130A

.subckt TMRDFFSNQNX1 QN D CLK SN
X0 a_1905_1004 a_217_1004 w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.714e+13p ps=3.0114e+08u w=2e+06u l=150000u M=2
X1  �� a_217_1004 a_757_75  �� sky130_fd_pr__nfet_01v8 ad=3.7611e+12p pd=3.297e+07u as=0p ps=0u w=3e+06u l=150000u
X2 a_5227_383 a_6149_943 a_5922_182  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3 w_n87_786 a_11673_1004 a_11033_943 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X4 QN a_8357_1004 a_16096_73  �� sky130_fd_pr__nfet_01v8 ad=5.373e+11p pd=4.72e+06u as=0p ps=0u w=3.01e+06u l=150000u
X5 a_5101_1004 a_5227_383 a_4996_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X6  �� D a_112_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X7 a_14869_1005 a_13241_1004 a_15533_1005 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X8 w_n87_786 a_343_383 a_217_1004 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X9 w_n87_786 a_5227_383 a_5101_1004 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X10 a_9178_182 SN a_8897_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X11  �� a_343_383 a_3368_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X12 w_n87_786 a_217_1004 a_343_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X13 a_11673_1004 a_11033_943 w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X14  �� a_8357_1004 a_8897_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X15 w_n87_786 a_13241_1004 a_13367_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X16 a_3473_1004 a_3599_383 w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X17 a_10111_383 CLK w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X18 a_6789_1004 a_6149_943 a_6884_182  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X19 a_5227_383 a_6149_943 w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X20 a_13241_1004 a_13367_383 w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X21 w_n87_786 a_11033_943 a_10111_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X22 w_n87_786 a_5227_383 a_8357_1004 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X23 a_6149_943 CLK w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X24 a_14869_1005 a_13241_1004 w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X25 w_n87_786 a_6149_943 a_8483_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X26 w_n87_786 CLK a_343_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X27 w_n87_786 a_8357_1004 a_14869_1005 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X28 a_3473_1004 a_343_383 w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X29  �� D a_9880_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X30 a_8483_383 SN w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X31 w_n87_786 SN a_13367_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X32 a_10111_383 a_9985_1004 w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X33 w_n87_786 a_1905_1004 a_1265_943 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X34  �� a_217_1004 a_1719_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X35 w_n87_786 a_10111_383 a_9985_1004 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X36 a_11033_943 CLK a_12470_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X37 w_n87_786 SN a_11673_1004 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X38 a_10111_383 a_11033_943 a_10806_182  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X39 a_6149_943 a_6789_1004 w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X40 a_9985_1004 a_10111_383 a_9880_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X41 w_n87_786 a_3473_1004 a_3599_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X42 QN a_3473_1004 a_15430_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X43 w_n87_786 a_1265_943 a_3599_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X44 a_14062_182 SN a_13781_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X45 a_1038_182 CLK a_757_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X46 w_n87_786 a_1265_943 a_343_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X47 a_8483_383 a_8357_1004 w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X48 w_n87_786 a_11033_943 a_13367_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X49 w_n87_786 a_5101_1004 a_5227_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X50 a_15533_1005 a_3473_1004 a_14869_1005 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X51 a_217_1004 D w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X52  �� a_10111_383 a_13136_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X53  �� a_1905_1004 a_2702_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X54 w_n87_786 D a_9985_1004 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X55 a_1905_1004 a_1265_943 w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X56  �� a_13241_1004 a_13781_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X57 a_6789_1004 a_5101_1004 w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X58  �� a_5227_383 a_8252_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X59 w_n87_786 a_9985_1004 a_11673_1004 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X60 a_217_1004 a_343_383 a_112_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X61 a_3599_383 a_1265_943 a_4294_182  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X62 a_11673_1004 a_11033_943 a_11768_182  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X63  �� a_5101_1004 a_5641_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X64 QN a_8357_1004 a_15533_1005 w_n87_786 sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=9.16e+06u as=0p ps=0u w=2e+06u l=150000u M=2
X65 a_2000_182 SN a_1719_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X66 w_n87_786 SN a_3599_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X67 w_n87_786 SN a_6789_1004 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X68  �� a_13241_1004 a_14764_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X69 a_3473_1004 a_3599_383 a_3368_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X70 a_1905_1004 SN w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X71 QN a_3473_1004 a_15533_1005 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X72 w_n87_786 a_8483_383 a_8357_1004 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X73  �� a_5101_1004 a_6603_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X74 w_n87_786 a_6149_943 a_6789_1004 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X75  �� a_3473_1004 a_4013_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X76 w_n87_786 a_10111_383 a_13241_1004 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X77 QN a_8357_1004 a_14764_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X78 a_5922_182 CLK a_5641_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X79 a_11033_943 CLK w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X80 a_5101_1004 D w_n87_786 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X81  �� a_6789_1004 a_7586_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X82  �� a_3473_1004 a_16096_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X83  �� a_9985_1004 a_10525_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X84  �� D a_4996_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X85 w_n87_786 CLK a_1265_943 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X86 a_1265_943 CLK a_2702_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X87 a_8483_383 a_6149_943 a_9178_182  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X88 a_8357_1004 a_8483_383 a_8252_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X89 a_6884_182 SN a_6603_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X90 a_13241_1004 a_13367_383 a_13136_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X91 a_4294_182 SN a_4013_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X92  �� a_9985_1004 a_11487_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X93 w_n87_786 CLK a_5227_383 w_n87_786 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X94 a_1905_1004 a_1265_943 a_2000_182  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X95 a_10806_182 CLK a_10525_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X96  �� a_11673_1004 a_12470_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X97  �� a_13241_1004 a_15430_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X98 a_343_383 a_1265_943 a_1038_182  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X99 a_13367_383 a_11033_943 a_14062_182  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X100 a_11768_182 SN a_11487_75  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X101 a_6149_943 CLK a_7586_73  �� sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
C0 w_n87_786 a_13367_383 2.34fF
C1 CLK a_10111_383 3.20fF
C2 CLK a_343_383 2.96fF
C3 a_6149_943 a_3473_1004 3.75fF
C4 w_n87_786 a_8357_1004 2.72fF
C5 a_11033_943 a_10111_383 2.89fF
C6 w_n87_786 a_11673_1004 2.09fF
C7 w_n87_786 a_5227_383 3.07fF
C8 CLK w_n87_786 5.44fF
C9 w_n87_786 a_8483_383 2.36fF
C10 CLK a_5227_383 3.80fF
C11 D a_3473_1004 7.04fF
C12 SN D 3.25fF
C13 a_8357_1004 a_3473_1004 6.70fF
C14 SN a_8357_1004 3.52fF
C15 w_n87_786 a_11033_943 2.18fF
C16 w_n87_786 a_3473_1004 2.77fF
C17 w_n87_786 a_6789_1004 2.09fF
C18 CLK a_3473_1004 2.26fF
C19 a_343_383 a_1265_943 2.89fF
C20 w_n87_786 a_3599_383 2.36fF
C21 a_11033_943 a_3473_1004 3.76fF
C22 w_n87_786 a_13241_1004 2.81fF
C23 SN a_3473_1004 2.72fF
C24 w_n87_786 a_6149_943 2.17fF
C25 w_n87_786 a_1265_943 2.17fF
C26 a_6149_943 a_5227_383 2.89fF
C27 w_n87_786 a_10111_383 3.07fF
C28 w_n87_786 a_1905_1004 2.09fF
C29 a_343_383 w_n87_786 3.07fF
C30 SN  �� 3.93fF
C31 D  �� 2.83fF
C32 a_8357_1004  �� 2.34fF **FLOATING
C33 a_3473_1004  �� 3.54fF **FLOATING
C34 w_n87_786  �� 39.51fF **FLOATING
.ends
