magic
tech sky130A
magscale 1 2
timestamp 1652319931
<< nwell >>
rect 87 1099 875 1550
rect 87 1093 220 1099
rect 87 1059 205 1093
rect 229 1059 263 1093
rect 87 1056 220 1059
rect 279 1056 875 1099
rect 87 786 875 1056
<< pwell >>
rect 34 -34 928 544
<< pdiffc >>
rect 201 1059 235 1093
rect 289 1059 323 1093
rect 465 1059 499 1093
rect 641 1059 675 1093
<< psubdiff >>
rect 34 482 928 544
rect 34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 928 17
rect 34 -34 928 -17
<< nsubdiff >>
rect 34 1497 928 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 928 1497
rect 34 822 928 884
<< psubdiffcont >>
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
<< poly >>
rect 147 383 195 413
rect 471 383 477 413
rect 147 377 177 383
rect 447 377 477 383
<< locali >>
rect 34 1497 928 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 928 1497
rect 34 1446 928 1463
rect 201 1093 235 1116
rect 201 1043 235 1059
rect 289 1093 323 1111
rect 289 1048 323 1059
rect 465 1093 499 1111
rect 465 1048 499 1059
rect 641 1093 675 1111
rect 641 1048 675 1059
rect 289 1014 831 1048
rect 205 433 239 908
rect 427 433 461 908
rect 649 449 683 940
rect 797 350 831 1014
rect 700 316 831 350
rect 700 235 734 316
rect 393 182 603 216
rect 198 34 232 167
rect 34 17 928 34
rect 34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 928 17
rect 34 -34 928 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
<< metal1 >>
rect 34 1497 928 1514
rect 34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 928 1497
rect 34 1446 928 1463
rect 34 17 928 34
rect 34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 928 17
rect 34 -34 928 -17
use poly_li1_contact  poly_li1_contact_0
timestamp 1648060378
transform 0 1 223 -1 0 941
box -32 -28 34 26
use pmos2  pmos2_0
timestamp 1648061063
transform 1 0 103 0 1 1404
box 52 -461 352 42
use nmos_bottom  nmos_bottom_0
timestamp 1651256857
transform -1 0 339 0 1 75
box 0 0 248 302
use poly_li1_contact  poly_li1_contact_1
timestamp 1648060378
transform 0 -1 221 1 0 415
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_3
timestamp 1648060378
transform 0 -1 443 1 0 939
box -32 -28 34 26
use pmos2  pmos2_2
timestamp 1648061063
transform 1 0 455 0 1 1404
box 52 -461 352 42
use pmos2  pmos2_1
timestamp 1648061063
transform 1 0 279 0 1 1404
box 52 -461 352 42
use nmos_side_left  nmos_side_left_0
timestamp 1651256873
transform 1 0 285 0 1 75
box 0 0 248 302
use poly_li1_contact  poly_li1_contact_2
timestamp 1648060378
transform 0 -1 443 1 0 415
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_5
timestamp 1648060378
transform 0 1 667 -1 0 941
box -32 -28 34 26
use nmos_top_trim1  nmos_top_trim1_0
timestamp 1651256895
transform -1 0 841 0 1 75
box 0 0 248 309
use poly_li1_contact  poly_li1_contact_4
timestamp 1648060378
transform 0 -1 665 1 0 415
box -32 -28 34 26
use diff_ring_side  diff_ring_side_1
timestamp 1652319726
transform 1 0 0 0 1 0
box -87 -34 87 1550
use diff_ring_side  diff_ring_side_0
timestamp 1652319726
transform 1 0 962 0 1 0
box -87 -34 87 1550
<< end >>
