* SPICE3 file created from DFFQX1.ext - technology: sky130A

.subckt DFFQX1 Q D CLK VDD GND
X0 GND dffx1_pcell_0/m1_2165_649# dffx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X1 dffx1_pcell_0/m1_258_797# CLK dffx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X2 VDD dffx1_pcell_0/m1_2165_649# dffx1_pcell_0/m1_258_797# VDD pshort w=2 l=0.15
X3 VDD CLK dffx1_pcell_0/m1_258_797# VDD pshort w=2 l=0.15
X4 GND dffx1_pcell_0/m1_833_723# dffx1_pcell_0/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X5 m1_3531_649# Q dffx1_pcell_0/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X6 VDD dffx1_pcell_0/m1_833_723# m1_3531_649# VDD pshort w=2 l=0.15
X7 VDD Q m1_3531_649# VDD pshort w=2 l=0.15
X8 GND m1_3531_649# dffx1_pcell_0/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X9 Q dffx1_pcell_0/m1_258_797# dffx1_pcell_0/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X10 VDD m1_3531_649# Q VDD pshort w=2 l=0.15
X11 VDD dffx1_pcell_0/m1_258_797# Q VDD pshort w=2 l=0.15
X12 GND dffx1_pcell_0/m1_258_797# dffx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X13 dffx1_pcell_0/m1_833_723# dffx1_pcell_0/m1_685_649# dffx1_pcell_0/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X14 dffx1_pcell_0/nand3x1_pcell_0/li_393_182# CLK dffx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X15 VDD dffx1_pcell_0/m1_258_797# dffx1_pcell_0/m1_833_723# VDD pshort w=2 l=0.15
X16 VDD CLK dffx1_pcell_0/m1_833_723# VDD pshort w=2 l=0.15
X17 VDD dffx1_pcell_0/m1_685_649# dffx1_pcell_0/m1_833_723# VDD pshort w=2 l=0.15
X18 GND dffx1_pcell_0/m1_833_723# dffx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X19 dffx1_pcell_0/m1_685_649# D dffx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X20 VDD dffx1_pcell_0/m1_833_723# dffx1_pcell_0/m1_685_649# VDD pshort w=2 l=0.15
X21 VDD D dffx1_pcell_0/m1_685_649# VDD pshort w=2 l=0.15
X22 GND dffx1_pcell_0/m1_685_649# dffx1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X23 dffx1_pcell_0/m1_2165_649# dffx1_pcell_0/m1_258_797# dffx1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X24 VDD dffx1_pcell_0/m1_685_649# dffx1_pcell_0/m1_2165_649# VDD pshort w=2 l=0.15
X25 VDD dffx1_pcell_0/m1_258_797# dffx1_pcell_0/m1_2165_649# VDD pshort w=2 l=0.15
C0 VDD dffx1_pcell_0/m1_258_797# 2.41fF
.ends
