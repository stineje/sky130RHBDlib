* SPICE3 file created from AOA4X1.ext - technology: sky130A

.subckt AOA4X1 Y A B C D VPB VNB
M1000 VNB a_168_157# a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=3.4356p pd=24.18u as=0p ps=0u
M1001 VNB a_864_181.t6 a_1444_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_1549_1004.t1 a_1675_383# VPB.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t10 a_168_157# a_217_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPB.t2 a_217_1004.t5 a_797_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPB.t5 a_343_383# a_217_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPB.t8 a_864_181.t4 a_1549_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPB.t0 a_1549_1004.t5 a_2183_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_797_1005.t2 a_1009_383# a_864_181.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_217_1004.t3 a_168_157# VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t6 a_1675_383# a_1549_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_217_1004.t1 a_343_383# VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_797_1005.t0 a_217_1004.t6 VPB.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1549_1004.t0 a_864_181.t5 VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_2183_182.t0 a_1549_1004.t7 VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_864_181.t1 a_1009_383# a_797_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VPB a_1009_383# 0.07fF
C1 VPB a_168_157# 0.08fF
C2 VPB a_343_383# 0.07fF
C3 VPB a_1675_383# 0.07fF
C4 a_343_383# a_168_157# 0.26fF
R0 a_1444_73.t0 a_1444_73.n1 34.62
R1 a_1444_73.t0 a_1444_73.n0 8.137
R2 a_1444_73.t0 a_1444_73.n2 4.69
R3 a_1549_1004.n4 a_1549_1004.t5 512.525
R4 a_1549_1004.n4 a_1549_1004.t7 371.139
R5 a_1549_1004.n6 a_1549_1004.n3 215.652
R6 a_1549_1004.n5 a_1549_1004.n4 211.406
R7 a_1549_1004.n5 a_1549_1004.t6 167.157
R8 a_1549_1004.n6 a_1549_1004.n5 153.043
R9 a_1549_1004.n8 a_1549_1004.n6 140.981
R10 a_1549_1004.n3 a_1549_1004.n2 76.002
R11 a_1549_1004.n9 a_1549_1004.n0 55.263
R12 a_1549_1004.n8 a_1549_1004.n7 30
R13 a_1549_1004.n9 a_1549_1004.n8 23.684
R14 a_1549_1004.n1 a_1549_1004.t2 14.282
R15 a_1549_1004.n1 a_1549_1004.t1 14.282
R16 a_1549_1004.n2 a_1549_1004.t4 14.282
R17 a_1549_1004.n2 a_1549_1004.t0 14.282
R18 a_1549_1004.n3 a_1549_1004.n1 12.85
R19 VPB VPB.n247 126.832
R20 VPB.n51 VPB.n49 94.117
R21 VPB.n210 VPB.n208 94.117
R22 VPB.n127 VPB.n125 94.117
R23 VPB.n187 VPB.n181 76.136
R24 VPB.n187 VPB.n186 76
R25 VPB.n191 VPB.n190 76
R26 VPB.n197 VPB.n196 76
R27 VPB.n211 VPB.n207 76
R28 VPB.n215 VPB.n214 76
R29 VPB.n219 VPB.n218 76
R30 VPB.n223 VPB.n222 76
R31 VPB.n228 VPB.n227 76
R32 VPB.n240 VPB.n239 76
R33 VPB.n194 VPB.n193 68.979
R34 VPB.n184 VPB.n183 64.528
R35 VPB.n21 VPB.n20 61.764
R36 VPB.n84 VPB.n83 61.764
R37 VPB.n106 VPB.n105 61.764
R38 VPB.n74 VPB.t11 55.106
R39 VPB.n150 VPB.t3 55.106
R40 VPB.n192 VPB.t1 55.106
R41 VPB.n182 VPB.t0 55.106
R42 VPB.n56 VPB.t5 55.106
R43 VPB.n132 VPB.t6 55.106
R44 VPB.n134 VPB.n133 48.952
R45 VPB.n58 VPB.n57 48.952
R46 VPB.n147 VPB.n146 44.502
R47 VPB.n39 VPB.n38 44.502
R48 VPB.n71 VPB.n70 44.502
R49 VPB.n37 VPB.n36 41.183
R50 VPB.n65 VPB.n14 40.824
R51 VPB.n141 VPB.n99 40.824
R52 VPB.n244 VPB.n240 20.452
R53 VPB.n181 VPB.n178 20.452
R54 VPB.n138 VPB.n137 17.801
R55 VPB.n62 VPB.n61 17.801
R56 VPB.n14 VPB.t4 14.282
R57 VPB.n14 VPB.t10 14.282
R58 VPB.n36 VPB.t9 14.282
R59 VPB.n36 VPB.t2 14.282
R60 VPB.n99 VPB.t7 14.282
R61 VPB.n99 VPB.t8 14.282
R62 VPB.n181 VPB.n180 13.653
R63 VPB.n180 VPB.n179 13.653
R64 VPB.n186 VPB.n185 13.653
R65 VPB.n185 VPB.n184 13.653
R66 VPB.n190 VPB.n189 13.653
R67 VPB.n189 VPB.n188 13.653
R68 VPB.n196 VPB.n195 13.653
R69 VPB.n195 VPB.n194 13.653
R70 VPB.n123 VPB.n122 13.653
R71 VPB.n122 VPB.n121 13.653
R72 VPB.n128 VPB.n127 13.653
R73 VPB.n127 VPB.n126 13.653
R74 VPB.n131 VPB.n130 13.653
R75 VPB.n130 VPB.n129 13.653
R76 VPB.n136 VPB.n135 13.653
R77 VPB.n135 VPB.n134 13.653
R78 VPB.n140 VPB.n139 13.653
R79 VPB.n139 VPB.n138 13.653
R80 VPB.n145 VPB.n144 13.653
R81 VPB.n144 VPB.n143 13.653
R82 VPB.n149 VPB.n148 13.653
R83 VPB.n148 VPB.n147 13.653
R84 VPB.n153 VPB.n152 13.653
R85 VPB.n152 VPB.n151 13.653
R86 VPB.n156 VPB.n155 13.653
R87 VPB.n155 VPB.n154 13.653
R88 VPB.n211 VPB.n210 13.653
R89 VPB.n210 VPB.n209 13.653
R90 VPB.n214 VPB.n213 13.653
R91 VPB.n213 VPB.n212 13.653
R92 VPB.n218 VPB.n217 13.653
R93 VPB.n217 VPB.n216 13.653
R94 VPB.n222 VPB.n221 13.653
R95 VPB.n221 VPB.n220 13.653
R96 VPB.n227 VPB.n226 13.653
R97 VPB.n226 VPB.n225 13.653
R98 VPB.n41 VPB.n40 13.653
R99 VPB.n40 VPB.n39 13.653
R100 VPB.n44 VPB.n43 13.653
R101 VPB.n43 VPB.n42 13.653
R102 VPB.n47 VPB.n46 13.653
R103 VPB.n46 VPB.n45 13.653
R104 VPB.n52 VPB.n51 13.653
R105 VPB.n51 VPB.n50 13.653
R106 VPB.n55 VPB.n54 13.653
R107 VPB.n54 VPB.n53 13.653
R108 VPB.n60 VPB.n59 13.653
R109 VPB.n59 VPB.n58 13.653
R110 VPB.n64 VPB.n63 13.653
R111 VPB.n63 VPB.n62 13.653
R112 VPB.n69 VPB.n68 13.653
R113 VPB.n68 VPB.n67 13.653
R114 VPB.n73 VPB.n72 13.653
R115 VPB.n72 VPB.n71 13.653
R116 VPB.n77 VPB.n76 13.653
R117 VPB.n76 VPB.n75 13.653
R118 VPB.n240 VPB.n0 13.653
R119 VPB VPB.n0 13.653
R120 VPB.n143 VPB.n142 13.35
R121 VPB.n225 VPB.n224 13.35
R122 VPB.n67 VPB.n66 13.35
R123 VPB.n244 VPB.n243 13.276
R124 VPB.n243 VPB.n241 13.276
R125 VPB.n35 VPB.n17 13.276
R126 VPB.n17 VPB.n15 13.276
R127 VPB.n98 VPB.n80 13.276
R128 VPB.n80 VPB.n78 13.276
R129 VPB.n120 VPB.n102 13.276
R130 VPB.n102 VPB.n100 13.276
R131 VPB.n124 VPB.n123 13.276
R132 VPB.n128 VPB.n124 13.276
R133 VPB.n131 VPB.n128 13.276
R134 VPB.n140 VPB.n136 13.276
R135 VPB.n149 VPB.n145 13.276
R136 VPB.n156 VPB.n153 13.276
R137 VPB.n157 VPB.n156 13.276
R138 VPB.n211 VPB.n157 13.276
R139 VPB.n214 VPB.n211 13.276
R140 VPB.n44 VPB.n41 13.276
R141 VPB.n47 VPB.n44 13.276
R142 VPB.n48 VPB.n47 13.276
R143 VPB.n52 VPB.n48 13.276
R144 VPB.n55 VPB.n52 13.276
R145 VPB.n64 VPB.n60 13.276
R146 VPB.n73 VPB.n69 13.276
R147 VPB.n240 VPB.n77 13.276
R148 VPB.n178 VPB.n160 13.276
R149 VPB.n160 VPB.n158 13.276
R150 VPB.n165 VPB.n163 12.796
R151 VPB.n165 VPB.n164 12.564
R152 VPB.n171 VPB.n170 12.198
R153 VPB.n173 VPB.n172 12.198
R154 VPB.n171 VPB.n168 12.198
R155 VPB.n136 VPB.n132 11.841
R156 VPB.n60 VPB.n56 11.841
R157 VPB.n150 VPB.n149 11.482
R158 VPB.n74 VPB.n73 11.482
R159 VPB.n178 VPB.n177 7.5
R160 VPB.n163 VPB.n162 7.5
R161 VPB.n170 VPB.n169 7.5
R162 VPB.n168 VPB.n167 7.5
R163 VPB.n160 VPB.n159 7.5
R164 VPB.n175 VPB.n161 7.5
R165 VPB.n102 VPB.n101 7.5
R166 VPB.n115 VPB.n114 7.5
R167 VPB.n109 VPB.n108 7.5
R168 VPB.n111 VPB.n110 7.5
R169 VPB.n104 VPB.n103 7.5
R170 VPB.n120 VPB.n119 7.5
R171 VPB.n80 VPB.n79 7.5
R172 VPB.n93 VPB.n92 7.5
R173 VPB.n87 VPB.n86 7.5
R174 VPB.n89 VPB.n88 7.5
R175 VPB.n82 VPB.n81 7.5
R176 VPB.n98 VPB.n97 7.5
R177 VPB.n17 VPB.n16 7.5
R178 VPB.n30 VPB.n29 7.5
R179 VPB.n24 VPB.n23 7.5
R180 VPB.n26 VPB.n25 7.5
R181 VPB.n19 VPB.n18 7.5
R182 VPB.n35 VPB.n34 7.5
R183 VPB.n243 VPB.n242 7.5
R184 VPB.n12 VPB.n11 7.5
R185 VPB.n6 VPB.n5 7.5
R186 VPB.n8 VPB.n7 7.5
R187 VPB.n2 VPB.n1 7.5
R188 VPB.n245 VPB.n244 7.5
R189 VPB.n48 VPB.n35 7.176
R190 VPB.n157 VPB.n98 7.176
R191 VPB.n124 VPB.n120 7.176
R192 VPB.n145 VPB.n141 6.817
R193 VPB.n69 VPB.n65 6.817
R194 VPB.n116 VPB.n113 6.729
R195 VPB.n112 VPB.n109 6.729
R196 VPB.n107 VPB.n104 6.729
R197 VPB.n94 VPB.n91 6.729
R198 VPB.n90 VPB.n87 6.729
R199 VPB.n85 VPB.n82 6.729
R200 VPB.n31 VPB.n28 6.729
R201 VPB.n27 VPB.n24 6.729
R202 VPB.n22 VPB.n19 6.729
R203 VPB.n13 VPB.n10 6.729
R204 VPB.n9 VPB.n6 6.729
R205 VPB.n4 VPB.n2 6.729
R206 VPB.n107 VPB.n106 6.728
R207 VPB.n112 VPB.n111 6.728
R208 VPB.n116 VPB.n115 6.728
R209 VPB.n119 VPB.n118 6.728
R210 VPB.n85 VPB.n84 6.728
R211 VPB.n90 VPB.n89 6.728
R212 VPB.n94 VPB.n93 6.728
R213 VPB.n97 VPB.n96 6.728
R214 VPB.n22 VPB.n21 6.728
R215 VPB.n27 VPB.n26 6.728
R216 VPB.n31 VPB.n30 6.728
R217 VPB.n34 VPB.n33 6.728
R218 VPB.n4 VPB.n3 6.728
R219 VPB.n9 VPB.n8 6.728
R220 VPB.n13 VPB.n12 6.728
R221 VPB.n246 VPB.n245 6.728
R222 VPB.n141 VPB.n140 6.458
R223 VPB.n65 VPB.n64 6.458
R224 VPB.n177 VPB.n176 6.398
R225 VPB.n41 VPB.n37 4.305
R226 VPB.n186 VPB.n182 2.691
R227 VPB.n196 VPB.n192 2.332
R228 VPB.n153 VPB.n150 1.794
R229 VPB.n77 VPB.n74 1.794
R230 VPB.n132 VPB.n131 1.435
R231 VPB.n56 VPB.n55 1.435
R232 VPB.n175 VPB.n166 1.402
R233 VPB.n175 VPB.n171 1.402
R234 VPB.n175 VPB.n173 1.402
R235 VPB.n175 VPB.n174 1.402
R236 VPB.n176 VPB.n175 0.735
R237 VPB.n175 VPB.n165 0.735
R238 VPB.n117 VPB.n116 0.387
R239 VPB.n117 VPB.n112 0.387
R240 VPB.n117 VPB.n107 0.387
R241 VPB.n118 VPB.n117 0.387
R242 VPB.n95 VPB.n94 0.387
R243 VPB.n95 VPB.n90 0.387
R244 VPB.n95 VPB.n85 0.387
R245 VPB.n96 VPB.n95 0.387
R246 VPB.n32 VPB.n31 0.387
R247 VPB.n32 VPB.n27 0.387
R248 VPB.n32 VPB.n22 0.387
R249 VPB.n33 VPB.n32 0.387
R250 VPB.n247 VPB.n13 0.387
R251 VPB.n247 VPB.n9 0.387
R252 VPB.n247 VPB.n4 0.387
R253 VPB.n247 VPB.n246 0.387
R254 VPB.n199 VPB.n198 0.272
R255 VPB.n207 VPB.n206 0.272
R256 VPB.n232 VPB.n231 0.272
R257 VPB.n239 VPB 0.198
R258 VPB.n191 VPB.n187 0.136
R259 VPB.n197 VPB.n191 0.136
R260 VPB.n198 VPB.n197 0.136
R261 VPB.n200 VPB.n199 0.136
R262 VPB.n201 VPB.n200 0.136
R263 VPB.n202 VPB.n201 0.136
R264 VPB.n203 VPB.n202 0.136
R265 VPB.n204 VPB.n203 0.136
R266 VPB.n205 VPB.n204 0.136
R267 VPB.n206 VPB.n205 0.136
R268 VPB.n219 VPB.n215 0.136
R269 VPB.n223 VPB.n219 0.136
R270 VPB.n228 VPB.n223 0.136
R271 VPB.n229 VPB.n228 0.136
R272 VPB.n230 VPB.n229 0.136
R273 VPB.n231 VPB.n230 0.136
R274 VPB.n233 VPB.n232 0.136
R275 VPB.n234 VPB.n233 0.136
R276 VPB.n235 VPB.n234 0.136
R277 VPB.n236 VPB.n235 0.136
R278 VPB.n237 VPB.n236 0.136
R279 VPB.n238 VPB.n237 0.136
R280 VPB.n239 VPB.n238 0.136
R281 VPB.n207 VPB 0.068
R282 VPB.n215 VPB 0.068
R283 a_217_1004.n4 a_217_1004.t6 486.819
R284 a_217_1004.n4 a_217_1004.t5 384.527
R285 a_217_1004.n6 a_217_1004.n3 215.652
R286 a_217_1004.n5 a_217_1004.t7 207.443
R287 a_217_1004.n5 a_217_1004.n4 169.7
R288 a_217_1004.n6 a_217_1004.n5 153.315
R289 a_217_1004.n8 a_217_1004.n6 140.981
R290 a_217_1004.n3 a_217_1004.n2 76.002
R291 a_217_1004.n8 a_217_1004.n7 30
R292 a_217_1004.n9 a_217_1004.n0 24.383
R293 a_217_1004.n9 a_217_1004.n8 23.684
R294 a_217_1004.n1 a_217_1004.t2 14.282
R295 a_217_1004.n1 a_217_1004.t1 14.282
R296 a_217_1004.n2 a_217_1004.t4 14.282
R297 a_217_1004.n2 a_217_1004.t3 14.282
R298 a_217_1004.n3 a_217_1004.n1 12.85
R299 a_797_1005.t1 a_797_1005.n0 101.66
R300 a_797_1005.n0 a_797_1005.t2 101.659
R301 a_797_1005.n0 a_797_1005.t3 14.294
R302 a_797_1005.n0 a_797_1005.t0 14.282
R303 a_864_181.n2 a_864_181.t4 480.392
R304 a_864_181.n2 a_864_181.t5 403.272
R305 a_864_181.n4 a_864_181.n1 228.489
R306 a_864_181.n3 a_864_181.t6 213.869
R307 a_864_181.n3 a_864_181.n2 161.6
R308 a_864_181.n4 a_864_181.n3 153.315
R309 a_864_181.n9 a_864_181.n8 118.016
R310 a_864_181.n9 a_864_181.n4 92.576
R311 a_864_181.n12 a_864_181.n0 55.263
R312 a_864_181.n11 a_864_181.n9 48.405
R313 a_864_181.n8 a_864_181.n7 30
R314 a_864_181.n11 a_864_181.n10 30
R315 a_864_181.n12 a_864_181.n11 25.263
R316 a_864_181.n6 a_864_181.n5 24.383
R317 a_864_181.n8 a_864_181.n6 23.684
R318 a_864_181.n1 a_864_181.t2 14.282
R319 a_864_181.n1 a_864_181.t1 14.282
R320 a_112_73.t0 a_112_73.n1 93.333
R321 a_112_73.n4 a_112_73.n2 55.07
R322 a_112_73.t0 a_112_73.n0 8.137
R323 a_112_73.n4 a_112_73.n3 4.619
R324 a_112_73.t0 a_112_73.n4 0.071
R325 VNB VNB.n238 300.778
R326 VNB.n89 VNB.n88 199.897
R327 VNB.n72 VNB.n71 199.897
R328 VNB.n15 VNB.n14 199.897
R329 VNB.n167 VNB.n166 158.304
R330 VNB.n188 VNB.n186 154.509
R331 VNB.n107 VNB.n105 154.509
R332 VNB.n38 VNB.n36 154.509
R333 VNB.n156 VNB.n155 105.536
R334 VNB.n121 VNB.n78 84.842
R335 VNB.n52 VNB.n4 84.842
R336 VNB.n159 VNB.n149 76.136
R337 VNB.n159 VNB.n158 76
R338 VNB.n225 VNB.n224 76
R339 VNB.n213 VNB.n212 76
R340 VNB.n205 VNB.n204 76
R341 VNB.n201 VNB.n200 76
R342 VNB.n194 VNB.n193 76
R343 VNB.n189 VNB.n185 76
R344 VNB.n175 VNB.n174 76
R345 VNB.n171 VNB.n170 76
R346 VNB.n98 VNB.t0 39.412
R347 VNB.n210 VNB.n209 36.937
R348 VNB.n123 VNB.n122 36.678
R349 VNB.n54 VNB.n53 36.678
R350 VNB.n199 VNB.n198 36.267
R351 VNB.n153 VNB.n152 35.01
R352 VNB.n168 VNB.n165 27.855
R353 VNB.n149 VNB.n146 20.452
R354 VNB.n226 VNB.n225 20.452
R355 VNB.n154 VNB.n153 20.094
R356 VNB.n164 VNB.n163 20.094
R357 VNB.n100 VNB.n99 20.094
R358 VNB.n25 VNB.n24 19.735
R359 VNB.n208 VNB.n207 19.735
R360 VNB.n197 VNB.n196 19.735
R361 VNB.n190 VNB.n61 19.735
R362 VNB.n31 VNB.n23 19.735
R363 VNB.n196 VNB.t3 19.724
R364 VNB.n153 VNB.n151 19.017
R365 VNB.n22 VNB.t1 17.353
R366 VNB.n98 VNB.n97 17.185
R367 VNB.n169 VNB.n168 16.721
R368 VNB.n158 VNB.n157 13.653
R369 VNB.n157 VNB.n156 13.653
R370 VNB.n170 VNB.n169 13.653
R371 VNB.n174 VNB.n173 13.653
R372 VNB.n173 VNB.n172 13.653
R373 VNB.n103 VNB.n102 13.653
R374 VNB.n102 VNB.n101 13.653
R375 VNB.n108 VNB.n107 13.653
R376 VNB.n107 VNB.n106 13.653
R377 VNB.n111 VNB.n110 13.653
R378 VNB.n110 VNB.n109 13.653
R379 VNB.n114 VNB.n113 13.653
R380 VNB.n113 VNB.n112 13.653
R381 VNB.n117 VNB.n116 13.653
R382 VNB.n116 VNB.n115 13.653
R383 VNB.n120 VNB.n119 13.653
R384 VNB.n119 VNB.n118 13.653
R385 VNB.n124 VNB.n123 13.653
R386 VNB.n127 VNB.n126 13.653
R387 VNB.n126 VNB.n125 13.653
R388 VNB.n130 VNB.n129 13.653
R389 VNB.n129 VNB.n128 13.653
R390 VNB.n189 VNB.n188 13.653
R391 VNB.n188 VNB.n187 13.653
R392 VNB.n193 VNB.n192 13.653
R393 VNB.n192 VNB.n191 13.653
R394 VNB.n200 VNB.n199 13.653
R395 VNB.n204 VNB.n203 13.653
R396 VNB.n203 VNB.n202 13.653
R397 VNB.n212 VNB.n211 13.653
R398 VNB.n211 VNB.n210 13.653
R399 VNB.n27 VNB.n26 13.653
R400 VNB.n30 VNB.n29 13.653
R401 VNB.n29 VNB.n28 13.653
R402 VNB.n34 VNB.n33 13.653
R403 VNB.n33 VNB.n32 13.653
R404 VNB.n39 VNB.n38 13.653
R405 VNB.n38 VNB.n37 13.653
R406 VNB.n42 VNB.n41 13.653
R407 VNB.n41 VNB.n40 13.653
R408 VNB.n45 VNB.n44 13.653
R409 VNB.n44 VNB.n43 13.653
R410 VNB.n48 VNB.n47 13.653
R411 VNB.n47 VNB.n46 13.653
R412 VNB.n51 VNB.n50 13.653
R413 VNB.n50 VNB.n49 13.653
R414 VNB.n55 VNB.n54 13.653
R415 VNB.n58 VNB.n57 13.653
R416 VNB.n57 VNB.n56 13.653
R417 VNB.n225 VNB.n0 13.653
R418 VNB VNB.n0 13.653
R419 VNB.n149 VNB.n148 13.653
R420 VNB.n148 VNB.n147 13.653
R421 VNB.n233 VNB.n230 13.577
R422 VNB.n134 VNB.n132 13.276
R423 VNB.n146 VNB.n134 13.276
R424 VNB.n81 VNB.n79 13.276
R425 VNB.n94 VNB.n81 13.276
R426 VNB.n64 VNB.n62 13.276
R427 VNB.n77 VNB.n64 13.276
R428 VNB.n7 VNB.n5 13.276
R429 VNB.n20 VNB.n7 13.276
R430 VNB.n104 VNB.n103 13.276
R431 VNB.n108 VNB.n104 13.276
R432 VNB.n111 VNB.n108 13.276
R433 VNB.n114 VNB.n111 13.276
R434 VNB.n117 VNB.n114 13.276
R435 VNB.n120 VNB.n117 13.276
R436 VNB.n127 VNB.n124 13.276
R437 VNB.n130 VNB.n127 13.276
R438 VNB.n131 VNB.n130 13.276
R439 VNB.n189 VNB.n131 13.276
R440 VNB.n30 VNB.n27 13.276
R441 VNB.n35 VNB.n34 13.276
R442 VNB.n39 VNB.n35 13.276
R443 VNB.n42 VNB.n39 13.276
R444 VNB.n45 VNB.n42 13.276
R445 VNB.n48 VNB.n45 13.276
R446 VNB.n51 VNB.n48 13.276
R447 VNB.n58 VNB.n55 13.276
R448 VNB.n225 VNB.n58 13.276
R449 VNB.n3 VNB.n1 13.276
R450 VNB.n226 VNB.n3 13.276
R451 VNB.n23 VNB.n22 12.837
R452 VNB.n190 VNB.n189 11.661
R453 VNB.n34 VNB.n31 11.661
R454 VNB.n61 VNB.n60 11.605
R455 VNB.n121 VNB.n120 10.764
R456 VNB.n52 VNB.n51 10.764
R457 VNB.n60 VNB.n59 9.809
R458 VNB.n103 VNB.n100 9.329
R459 VNB.n22 VNB.n21 7.566
R460 VNB.n151 VNB.n150 7.5
R461 VNB.n162 VNB.n161 7.5
R462 VNB.n235 VNB.n234 7.5
R463 VNB.n87 VNB.n86 7.5
R464 VNB.n83 VNB.n82 7.5
R465 VNB.n81 VNB.n80 7.5
R466 VNB.n94 VNB.n93 7.5
R467 VNB.n70 VNB.n69 7.5
R468 VNB.n66 VNB.n65 7.5
R469 VNB.n64 VNB.n63 7.5
R470 VNB.n77 VNB.n76 7.5
R471 VNB.n13 VNB.n12 7.5
R472 VNB.n9 VNB.n8 7.5
R473 VNB.n7 VNB.n6 7.5
R474 VNB.n20 VNB.n19 7.5
R475 VNB.n227 VNB.n226 7.5
R476 VNB.n3 VNB.n2 7.5
R477 VNB.n232 VNB.n231 7.5
R478 VNB.n140 VNB.n139 7.5
R479 VNB.n136 VNB.n135 7.5
R480 VNB.n134 VNB.n133 7.5
R481 VNB.n146 VNB.n145 7.5
R482 VNB.n104 VNB.n94 7.176
R483 VNB.n131 VNB.n77 7.176
R484 VNB.n35 VNB.n20 7.176
R485 VNB.t3 VNB.n195 7.04
R486 VNB.n237 VNB.n235 7.011
R487 VNB.n90 VNB.n87 7.011
R488 VNB.n85 VNB.n83 7.011
R489 VNB.n73 VNB.n70 7.011
R490 VNB.n68 VNB.n66 7.011
R491 VNB.n16 VNB.n13 7.011
R492 VNB.n11 VNB.n9 7.011
R493 VNB.n142 VNB.n140 7.011
R494 VNB.n138 VNB.n136 7.011
R495 VNB.n93 VNB.n92 7.01
R496 VNB.n85 VNB.n84 7.01
R497 VNB.n90 VNB.n89 7.01
R498 VNB.n76 VNB.n75 7.01
R499 VNB.n68 VNB.n67 7.01
R500 VNB.n73 VNB.n72 7.01
R501 VNB.n19 VNB.n18 7.01
R502 VNB.n11 VNB.n10 7.01
R503 VNB.n16 VNB.n15 7.01
R504 VNB.n145 VNB.n144 7.01
R505 VNB.n138 VNB.n137 7.01
R506 VNB.n142 VNB.n141 7.01
R507 VNB.n237 VNB.n236 7.01
R508 VNB.n233 VNB.n232 6.788
R509 VNB.n228 VNB.n227 6.788
R510 VNB.n212 VNB.n208 6.638
R511 VNB.n99 VNB.n98 6.139
R512 VNB.n207 VNB.n206 5.774
R513 VNB.n96 VNB.n95 4.551
R514 VNB.n158 VNB.n154 4.305
R515 VNB.n124 VNB.n121 2.511
R516 VNB.n200 VNB.n197 2.511
R517 VNB.n27 VNB.n25 2.511
R518 VNB.n55 VNB.n52 2.511
R519 VNB.t0 VNB.n96 2.238
R520 VNB.n168 VNB.n167 1.99
R521 VNB.n161 VNB.n160 1.935
R522 VNB.n193 VNB.n190 1.614
R523 VNB.n31 VNB.n30 1.614
R524 VNB.n238 VNB.n229 0.921
R525 VNB.n238 VNB.n233 0.476
R526 VNB.n238 VNB.n228 0.475
R527 VNB.n163 VNB.n162 0.358
R528 VNB.n177 VNB.n176 0.272
R529 VNB.n185 VNB.n184 0.272
R530 VNB.n217 VNB.n216 0.272
R531 VNB.n91 VNB.n85 0.246
R532 VNB.n92 VNB.n91 0.246
R533 VNB.n91 VNB.n90 0.246
R534 VNB.n74 VNB.n68 0.246
R535 VNB.n75 VNB.n74 0.246
R536 VNB.n74 VNB.n73 0.246
R537 VNB.n17 VNB.n11 0.246
R538 VNB.n18 VNB.n17 0.246
R539 VNB.n17 VNB.n16 0.246
R540 VNB.n143 VNB.n138 0.246
R541 VNB.n144 VNB.n143 0.246
R542 VNB.n143 VNB.n142 0.246
R543 VNB.n238 VNB.n237 0.246
R544 VNB.n224 VNB 0.198
R545 VNB.n170 VNB.n164 0.179
R546 VNB.n171 VNB.n159 0.136
R547 VNB.n175 VNB.n171 0.136
R548 VNB.n176 VNB.n175 0.136
R549 VNB.n178 VNB.n177 0.136
R550 VNB.n179 VNB.n178 0.136
R551 VNB.n180 VNB.n179 0.136
R552 VNB.n181 VNB.n180 0.136
R553 VNB.n182 VNB.n181 0.136
R554 VNB.n183 VNB.n182 0.136
R555 VNB.n184 VNB.n183 0.136
R556 VNB.n201 VNB.n194 0.136
R557 VNB.n205 VNB.n201 0.136
R558 VNB.n213 VNB.n205 0.136
R559 VNB.n214 VNB.n213 0.136
R560 VNB.n215 VNB.n214 0.136
R561 VNB.n216 VNB.n215 0.136
R562 VNB.n218 VNB.n217 0.136
R563 VNB.n219 VNB.n218 0.136
R564 VNB.n220 VNB.n219 0.136
R565 VNB.n221 VNB.n220 0.136
R566 VNB.n222 VNB.n221 0.136
R567 VNB.n223 VNB.n222 0.136
R568 VNB.n224 VNB.n223 0.136
R569 VNB.n185 VNB 0.068
R570 VNB.n194 VNB 0.068
R571 a_2183_182.n2 a_2183_182.n0 362.371
R572 a_2183_182.n2 a_2183_182.n1 15.218
R573 a_2183_182.n0 a_2183_182.t1 14.282
R574 a_2183_182.n0 a_2183_182.t0 14.282
R575 a_2183_182.n3 a_2183_182.n2 12.014
C5 VPB VNB 10.40fF
C6 a_2183_182.n0 VNB 1.03fF
C7 a_2183_182.n1 VNB 0.09fF
C8 a_2183_182.n2 VNB 0.49fF
C9 a_2183_182.n3 VNB 0.05fF
C10 a_112_73.n0 VNB 0.05fF
C11 a_112_73.n1 VNB 0.02fF
C12 a_112_73.n2 VNB 0.12fF
C13 a_112_73.n3 VNB 0.04fF
C14 a_112_73.n4 VNB 0.16fF
C15 a_864_181.n0 VNB 0.04fF
C16 a_864_181.n1 VNB 0.62fF
C17 a_864_181.n2 VNB 0.38fF
C18 a_864_181.n3 VNB 0.46fF
C19 a_864_181.n4 VNB 0.46fF
C20 a_864_181.n5 VNB 0.03fF
C21 a_864_181.n6 VNB 0.05fF
C22 a_864_181.n7 VNB 0.03fF
C23 a_864_181.n8 VNB 0.15fF
C24 a_864_181.n9 VNB 0.26fF
C25 a_864_181.n10 VNB 0.03fF
C26 a_864_181.n11 VNB 0.08fF
C27 a_864_181.n12 VNB 0.04fF
C28 a_797_1005.n0 VNB 0.55fF
C29 a_217_1004.n0 VNB 0.03fF
C30 a_217_1004.n1 VNB 0.43fF
C31 a_217_1004.n2 VNB 0.51fF
C32 a_217_1004.n3 VNB 0.31fF
C33 a_217_1004.n4 VNB 0.35fF
C34 a_217_1004.t7 VNB 0.38fF
C35 a_217_1004.n5 VNB 0.45fF
C36 a_217_1004.n6 VNB 0.49fF
C37 a_217_1004.n7 VNB 0.03fF
C38 a_217_1004.n8 VNB 0.17fF
C39 a_217_1004.n9 VNB 0.04fF
C40 VPB.n0 VNB 0.03fF
C41 VPB.n1 VNB 0.03fF
C42 VPB.n2 VNB 0.02fF
C43 VPB.n3 VNB 0.13fF
C44 VPB.n5 VNB 0.02fF
C45 VPB.n6 VNB 0.02fF
C46 VPB.n7 VNB 0.02fF
C47 VPB.n8 VNB 0.02fF
C48 VPB.n10 VNB 0.02fF
C49 VPB.n11 VNB 0.02fF
C50 VPB.n12 VNB 0.02fF
C51 VPB.n14 VNB 0.10fF
C52 VPB.n15 VNB 0.02fF
C53 VPB.n16 VNB 0.02fF
C54 VPB.n17 VNB 0.02fF
C55 VPB.n18 VNB 0.03fF
C56 VPB.n19 VNB 0.02fF
C57 VPB.n20 VNB 0.19fF
C58 VPB.n21 VNB 0.04fF
C59 VPB.n23 VNB 0.02fF
C60 VPB.n24 VNB 0.02fF
C61 VPB.n25 VNB 0.02fF
C62 VPB.n26 VNB 0.02fF
C63 VPB.n28 VNB 0.02fF
C64 VPB.n29 VNB 0.02fF
C65 VPB.n30 VNB 0.02fF
C66 VPB.n32 VNB 0.26fF
C67 VPB.n34 VNB 0.02fF
C68 VPB.n35 VNB 0.02fF
C69 VPB.n36 VNB 0.10fF
C70 VPB.n37 VNB 0.02fF
C71 VPB.n38 VNB 0.13fF
C72 VPB.n39 VNB 0.15fF
C73 VPB.n40 VNB 0.02fF
C74 VPB.n41 VNB 0.02fF
C75 VPB.n42 VNB 0.23fF
C76 VPB.n43 VNB 0.02fF
C77 VPB.n44 VNB 0.02fF
C78 VPB.n45 VNB 0.26fF
C79 VPB.n46 VNB 0.01fF
C80 VPB.n47 VNB 0.02fF
C81 VPB.n48 VNB 0.03fF
C82 VPB.n49 VNB 0.03fF
C83 VPB.n50 VNB 0.26fF
C84 VPB.n51 VNB 0.01fF
C85 VPB.n52 VNB 0.02fF
C86 VPB.n53 VNB 0.22fF
C87 VPB.n54 VNB 0.02fF
C88 VPB.n55 VNB 0.01fF
C89 VPB.n56 VNB 0.05fF
C90 VPB.n57 VNB 0.13fF
C91 VPB.n58 VNB 0.15fF
C92 VPB.n59 VNB 0.02fF
C93 VPB.n60 VNB 0.02fF
C94 VPB.n61 VNB 0.13fF
C95 VPB.n62 VNB 0.14fF
C96 VPB.n63 VNB 0.02fF
C97 VPB.n64 VNB 0.02fF
C98 VPB.n65 VNB 0.02fF
C99 VPB.n66 VNB 0.13fF
C100 VPB.n67 VNB 0.14fF
C101 VPB.n68 VNB 0.02fF
C102 VPB.n69 VNB 0.02fF
C103 VPB.n70 VNB 0.13fF
C104 VPB.n71 VNB 0.15fF
C105 VPB.n72 VNB 0.02fF
C106 VPB.n73 VNB 0.02fF
C107 VPB.n74 VNB 0.06fF
C108 VPB.n75 VNB 0.23fF
C109 VPB.n76 VNB 0.02fF
C110 VPB.n77 VNB 0.01fF
C111 VPB.n78 VNB 0.02fF
C112 VPB.n79 VNB 0.02fF
C113 VPB.n80 VNB 0.02fF
C114 VPB.n81 VNB 0.03fF
C115 VPB.n82 VNB 0.02fF
C116 VPB.n83 VNB 0.19fF
C117 VPB.n84 VNB 0.04fF
C118 VPB.n86 VNB 0.02fF
C119 VPB.n87 VNB 0.02fF
C120 VPB.n88 VNB 0.02fF
C121 VPB.n89 VNB 0.02fF
C122 VPB.n91 VNB 0.02fF
C123 VPB.n92 VNB 0.02fF
C124 VPB.n93 VNB 0.02fF
C125 VPB.n95 VNB 0.26fF
C126 VPB.n97 VNB 0.02fF
C127 VPB.n98 VNB 0.02fF
C128 VPB.n99 VNB 0.10fF
C129 VPB.n100 VNB 0.02fF
C130 VPB.n101 VNB 0.02fF
C131 VPB.n102 VNB 0.02fF
C132 VPB.n103 VNB 0.03fF
C133 VPB.n104 VNB 0.02fF
C134 VPB.n105 VNB 0.16fF
C135 VPB.n106 VNB 0.04fF
C136 VPB.n108 VNB 0.02fF
C137 VPB.n109 VNB 0.02fF
C138 VPB.n110 VNB 0.02fF
C139 VPB.n111 VNB 0.02fF
C140 VPB.n113 VNB 0.02fF
C141 VPB.n114 VNB 0.02fF
C142 VPB.n115 VNB 0.02fF
C143 VPB.n117 VNB 0.26fF
C144 VPB.n119 VNB 0.02fF
C145 VPB.n120 VNB 0.02fF
C146 VPB.n121 VNB 0.26fF
C147 VPB.n122 VNB 0.01fF
C148 VPB.n123 VNB 0.02fF
C149 VPB.n124 VNB 0.03fF
C150 VPB.n125 VNB 0.03fF
C151 VPB.n126 VNB 0.26fF
C152 VPB.n127 VNB 0.01fF
C153 VPB.n128 VNB 0.02fF
C154 VPB.n129 VNB 0.22fF
C155 VPB.n130 VNB 0.02fF
C156 VPB.n131 VNB 0.01fF
C157 VPB.n132 VNB 0.05fF
C158 VPB.n133 VNB 0.13fF
C159 VPB.n134 VNB 0.15fF
C160 VPB.n135 VNB 0.02fF
C161 VPB.n136 VNB 0.02fF
C162 VPB.n137 VNB 0.13fF
C163 VPB.n138 VNB 0.14fF
C164 VPB.n139 VNB 0.02fF
C165 VPB.n140 VNB 0.02fF
C166 VPB.n141 VNB 0.02fF
C167 VPB.n142 VNB 0.13fF
C168 VPB.n143 VNB 0.14fF
C169 VPB.n144 VNB 0.02fF
C170 VPB.n145 VNB 0.02fF
C171 VPB.n146 VNB 0.13fF
C172 VPB.n147 VNB 0.15fF
C173 VPB.n148 VNB 0.02fF
C174 VPB.n149 VNB 0.02fF
C175 VPB.n150 VNB 0.06fF
C176 VPB.n151 VNB 0.23fF
C177 VPB.n152 VNB 0.02fF
C178 VPB.n153 VNB 0.01fF
C179 VPB.n154 VNB 0.26fF
C180 VPB.n155 VNB 0.01fF
C181 VPB.n156 VNB 0.02fF
C182 VPB.n157 VNB 0.03fF
C183 VPB.n158 VNB 0.02fF
C184 VPB.n159 VNB 0.02fF
C185 VPB.n160 VNB 0.02fF
C186 VPB.n161 VNB 0.10fF
C187 VPB.n162 VNB 0.03fF
C188 VPB.n163 VNB 0.02fF
C189 VPB.n164 VNB 0.04fF
C190 VPB.n165 VNB 0.01fF
C191 VPB.n167 VNB 0.02fF
C192 VPB.n168 VNB 0.02fF
C193 VPB.n169 VNB 0.02fF
C194 VPB.n170 VNB 0.02fF
C195 VPB.n172 VNB 0.02fF
C196 VPB.n175 VNB 0.44fF
C197 VPB.n177 VNB 0.03fF
C198 VPB.n178 VNB 0.04fF
C199 VPB.n179 VNB 0.26fF
C200 VPB.n180 VNB 0.03fF
C201 VPB.n181 VNB 0.03fF
C202 VPB.n182 VNB 0.05fF
C203 VPB.n183 VNB 0.13fF
C204 VPB.n184 VNB 0.18fF
C205 VPB.n185 VNB 0.02fF
C206 VPB.n186 VNB 0.01fF
C207 VPB.n187 VNB 0.07fF
C208 VPB.n188 VNB 0.15fF
C209 VPB.n189 VNB 0.02fF
C210 VPB.n190 VNB 0.02fF
C211 VPB.n191 VNB 0.02fF
C212 VPB.n192 VNB 0.06fF
C213 VPB.n193 VNB 0.13fF
C214 VPB.n194 VNB 0.18fF
C215 VPB.n195 VNB 0.02fF
C216 VPB.n196 VNB 0.01fF
C217 VPB.n197 VNB 0.02fF
C218 VPB.n198 VNB 0.03fF
C219 VPB.n199 VNB 0.03fF
C220 VPB.n200 VNB 0.02fF
C221 VPB.n201 VNB 0.02fF
C222 VPB.n202 VNB 0.02fF
C223 VPB.n203 VNB 0.02fF
C224 VPB.n204 VNB 0.02fF
C225 VPB.n205 VNB 0.02fF
C226 VPB.n206 VNB 0.03fF
C227 VPB.n207 VNB 0.03fF
C228 VPB.n208 VNB 0.03fF
C229 VPB.n209 VNB 0.26fF
C230 VPB.n210 VNB 0.01fF
C231 VPB.n211 VNB 0.02fF
C232 VPB.n212 VNB 0.26fF
C233 VPB.n213 VNB 0.02fF
C234 VPB.n214 VNB 0.02fF
C235 VPB.n215 VNB 0.02fF
C236 VPB.n216 VNB 0.26fF
C237 VPB.n217 VNB 0.02fF
C238 VPB.n218 VNB 0.02fF
C239 VPB.n219 VNB 0.02fF
C240 VPB.n220 VNB 0.26fF
C241 VPB.n221 VNB 0.02fF
C242 VPB.n222 VNB 0.02fF
C243 VPB.n223 VNB 0.02fF
C244 VPB.n224 VNB 0.13fF
C245 VPB.n225 VNB 0.14fF
C246 VPB.n226 VNB 0.02fF
C247 VPB.n227 VNB 0.02fF
C248 VPB.n228 VNB 0.02fF
C249 VPB.n229 VNB 0.02fF
C250 VPB.n230 VNB 0.02fF
C251 VPB.n231 VNB 0.03fF
C252 VPB.n232 VNB 0.03fF
C253 VPB.n233 VNB 0.02fF
C254 VPB.n234 VNB 0.02fF
C255 VPB.n235 VNB 0.02fF
C256 VPB.n236 VNB 0.02fF
C257 VPB.n237 VNB 0.02fF
C258 VPB.n238 VNB 0.02fF
C259 VPB.n239 VNB 0.03fF
C260 VPB.n240 VNB 0.03fF
C261 VPB.n241 VNB 0.02fF
C262 VPB.n242 VNB 0.02fF
C263 VPB.n243 VNB 0.02fF
C264 VPB.n244 VNB 0.04fF
C265 VPB.n245 VNB 0.03fF
C266 VPB.n247 VNB 0.41fF
C267 a_1549_1004.n0 VNB 0.05fF
C268 a_1549_1004.n1 VNB 0.42fF
C269 a_1549_1004.n2 VNB 0.50fF
C270 a_1549_1004.n3 VNB 0.30fF
C271 a_1549_1004.n4 VNB 0.33fF
C272 a_1549_1004.t6 VNB 0.37fF
C273 a_1549_1004.n5 VNB 0.45fF
C274 a_1549_1004.n6 VNB 0.45fF
C275 a_1549_1004.n7 VNB 0.02fF
C276 a_1549_1004.n8 VNB 0.17fF
C277 a_1549_1004.n9 VNB 0.04fF
C278 a_1444_73.n0 VNB 0.05fF
C279 a_1444_73.n1 VNB 0.12fF
C280 a_1444_73.n2 VNB 0.04fF
.ends
