// File: nor3x1_pcell.spi.pex
// Created: Tue Oct 15 15:59:36 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_NOR3X1_PCELL\%noxref_1 ( 9 21 25 33 37 45 49 60 63 90 )
c51 ( 90 0 ) capacitor c=0.0964353f //x=0.56 //y=0.365
c52 ( 63 0 ) capacitor c=0.203672f //x=0.695 //y=0
c53 ( 60 0 ) capacitor c=0.250916f //x=4.07 //y=0
c54 ( 58 0 ) capacitor c=0.095941f //x=3.69 //y=0
c55 ( 52 0 ) capacitor c=0.00803396f //x=3.605 //y=0.445
c56 ( 49 0 ) capacitor c=0.00510317f //x=3.52 //y=0.53
c57 ( 48 0 ) capacitor c=0.00468234f //x=3.12 //y=0.445
c58 ( 45 0 ) capacitor c=0.00514697f //x=3.035 //y=0.53
c59 ( 40 0 ) capacitor c=0.00468234f //x=2.635 //y=0.445
c60 ( 37 0 ) capacitor c=0.00556167f //x=2.55 //y=0.53
c61 ( 36 0 ) capacitor c=0.00468234f //x=2.15 //y=0.445
c62 ( 33 0 ) capacitor c=0.00556167f //x=2.065 //y=0.53
c63 ( 28 0 ) capacitor c=0.00468234f //x=1.665 //y=0.445
c64 ( 25 0 ) capacitor c=0.00556167f //x=1.58 //y=0.53
c65 ( 24 0 ) capacitor c=0.00468234f //x=1.18 //y=0.445
c66 ( 21 0 ) capacitor c=0.00709092f //x=1.095 //y=0.53
c67 ( 16 0 ) capacitor c=0.00609805f //x=0.695 //y=0.445
c68 ( 9 0 ) capacitor c=0.207649f //x=4.07 //y=0
r69 (  74 75 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.12 //y=0 //x2=3.605 //y2=0
r70 (  73 74 ) resistor r=5.73669 //w=0.357 //l=0.16 //layer=li \
 //thickness=0.1 //x=2.96 //y=0 //x2=3.12 //y2=0
r71 (  71 73 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=2.635 //y=0 //x2=2.96 //y2=0
r72 (  70 71 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.15 //y=0 //x2=2.635 //y2=0
r73 (  69 70 ) resistor r=10.7563 //w=0.357 //l=0.3 //layer=li //thickness=0.1 \
 //x=1.85 //y=0 //x2=2.15 //y2=0
r74 (  67 69 ) resistor r=6.63305 //w=0.357 //l=0.185 //layer=li \
 //thickness=0.1 //x=1.665 //y=0 //x2=1.85 //y2=0
r75 (  66 67 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.18 //y=0 //x2=1.665 //y2=0
r76 (  65 66 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.18 //y2=0
r77 (  63 65 ) resistor r=1.61345 //w=0.357 //l=0.045 //layer=li \
 //thickness=0.1 //x=0.695 //y=0 //x2=0.74 //y2=0
r78 (  58 75 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.69 //y=0 //x2=3.605 //y2=0
r79 (  58 60 ) resistor r=13.6247 //w=0.357 //l=0.38 //layer=li \
 //thickness=0.1 //x=3.69 //y=0 //x2=4.07 //y2=0
r80 (  53 90 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.605 //y=0.615 //x2=3.605 //y2=0.53
r81 (  53 90 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=3.605 //y=0.615 //x2=3.605 //y2=0.88
r82 (  52 90 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.605 //y=0.445 //x2=3.605 //y2=0.53
r83 (  51 75 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.605 //y=0.17 //x2=3.605 //y2=0
r84 (  51 52 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=3.605 //y=0.17 //x2=3.605 //y2=0.445
r85 (  50 90 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.205 //y=0.53 //x2=3.12 //y2=0.53
r86 (  49 90 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.52 //y=0.53 //x2=3.605 //y2=0.53
r87 (  49 50 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.52 //y=0.53 //x2=3.205 //y2=0.53
r88 (  48 90 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.12 //y=0.445 //x2=3.12 //y2=0.53
r89 (  47 74 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.12 //y=0.17 //x2=3.12 //y2=0
r90 (  47 48 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=3.12 //y=0.17 //x2=3.12 //y2=0.445
r91 (  46 90 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.72 //y=0.53 //x2=2.635 //y2=0.53
r92 (  45 90 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.035 //y=0.53 //x2=3.12 //y2=0.53
r93 (  45 46 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.035 //y=0.53 //x2=2.72 //y2=0.53
r94 (  41 90 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.635 //y=0.615 //x2=2.635 //y2=0.53
r95 (  41 90 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r96 (  40 90 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.635 //y=0.445 //x2=2.635 //y2=0.53
r97 (  39 71 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.635 //y=0.17 //x2=2.635 //y2=0
r98 (  39 40 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.17 //x2=2.635 //y2=0.445
r99 (  38 90 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.235 //y=0.53 //x2=2.15 //y2=0.53
r100 (  37 90 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.55 //y=0.53 //x2=2.635 //y2=0.53
r101 (  37 38 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.235 //y2=0.53
r102 (  36 90 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.445 //x2=2.15 //y2=0.53
r103 (  35 70 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.17 //x2=2.15 //y2=0
r104 (  35 36 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.17 //x2=2.15 //y2=0.445
r105 (  34 90 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=1.665 //y2=0.53
r106 (  33 90 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.065 //y=0.53 //x2=2.15 //y2=0.53
r107 (  33 34 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=2.065 //y=0.53 //x2=1.75 //y2=0.53
r108 (  29 90 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.53
r109 (  29 90 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r110 (  28 90 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.445 //x2=1.665 //y2=0.53
r111 (  27 67 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.17 //x2=1.665 //y2=0
r112 (  27 28 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.17 //x2=1.665 //y2=0.445
r113 (  26 90 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0.53 //x2=1.18 //y2=0.53
r114 (  25 90 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.58 //y=0.53 //x2=1.665 //y2=0.53
r115 (  25 26 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.58 //y=0.53 //x2=1.265 //y2=0.53
r116 (  24 90 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.445 //x2=1.18 //y2=0.53
r117 (  23 66 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r118 (  23 24 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.445
r119 (  22 90 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.78 //y=0.53 //x2=0.695 //y2=0.53
r120 (  21 90 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0.53 //x2=1.18 //y2=0.53
r121 (  21 22 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.095 //y=0.53 //x2=0.78 //y2=0.53
r122 (  17 90 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.615 //x2=0.695 //y2=0.53
r123 (  17 90 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.615 //x2=0.695 //y2=1.22
r124 (  16 90 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.445 //x2=0.695 //y2=0.53
r125 (  15 63 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.17 //x2=0.695 //y2=0
r126 (  15 16 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.17 //x2=0.695 //y2=0.445
r127 (  9 60 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r128 (  7 73 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r129 (  7 9 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.07 //y2=0
r130 (  5 69 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r131 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r132 (  2 65 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r133 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
ends PM_NOR3X1_PCELL\%noxref_1

subckt PM_NOR3X1_PCELL\%noxref_2 ( 9 13 16 30 34 )
c42 ( 34 0 ) capacitor c=0.0267864f //x=1.085 //y=5.025
c43 ( 33 0 ) capacitor c=0.00591168f //x=1.23 //y=7.4
c44 ( 30 0 ) capacitor c=0.351373f //x=4.07 //y=7.4
c45 ( 16 0 ) capacitor c=0.211583f //x=0.74 //y=7.4
c46 ( 13 0 ) capacitor c=0.0465804f //x=1.145 //y=7.4
c47 ( 9 0 ) capacitor c=0.203056f //x=4.07 //y=7.4
r48 (  28 30 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r49 (  26 28 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r50 (  24 33 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.315 //y=7.4 //x2=1.23 //y2=7.4
r51 (  24 26 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=1.315 //y=7.4 //x2=1.85 //y2=7.4
r52 (  17 33 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.23 //y=7.23 //x2=1.23 //y2=7.4
r53 (  17 34 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=1.23 //y=7.23 //x2=1.23 //y2=6.74
r54 (  13 33 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.145 //y=7.4 //x2=1.23 //y2=7.4
r55 (  13 16 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=1.145 //y=7.4 //x2=0.74 //y2=7.4
r56 (  9 30 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=4.07 \
 //y=7.4 //x2=4.07 //y2=7.4
r57 (  7 28 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=2.96 \
 //y=7.4 //x2=2.96 //y2=7.4
r58 (  7 9 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r59 (  5 26 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=1.85 \
 //y=7.4 //x2=1.85 //y2=7.4
r60 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r61 (  2 16 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=0.74 \
 //y=7.4 //x2=0.74 //y2=7.4
r62 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_NOR3X1_PCELL\%noxref_2

subckt PM_NOR3X1_PCELL\%noxref_3 ( 3 6 8 9 10 11 12 13 14 18 20 23 25 26 31 )
c65 ( 31 0 ) capacitor c=0.04214f //x=0.955 //y=4.705
c66 ( 26 0 ) capacitor c=0.0321911f //x=1.445 //y=1.25
c67 ( 25 0 ) capacitor c=0.0185201f //x=1.445 //y=0.905
c68 ( 23 0 ) capacitor c=0.0344254f //x=1.375 //y=4.795
c69 ( 20 0 ) capacitor c=0.0133656f //x=1.29 //y=1.405
c70 ( 18 0 ) capacitor c=0.0157804f //x=1.29 //y=0.75
c71 ( 14 0 ) capacitor c=0.0828832f //x=0.915 //y=1.915
c72 ( 13 0 ) capacitor c=0.022867f //x=0.915 //y=1.56
c73 ( 12 0 ) capacitor c=0.0234318f //x=0.915 //y=1.25
c74 ( 11 0 ) capacitor c=0.0192004f //x=0.915 //y=0.905
c75 ( 10 0 ) capacitor c=0.110795f //x=1.45 //y=6.025
c76 ( 9 0 ) capacitor c=0.153847f //x=1.01 //y=6.025
c77 ( 6 0 ) capacitor c=0.00995068f //x=0.955 //y=4.705
c78 ( 3 0 ) capacitor c=0.112895f //x=1.11 //y=2.08
r79 (  33 34 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=0.955 //y=4.795 //x2=0.955 //y2=4.87
r80 (  31 33 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=0.955 //y=4.705 //x2=0.955 //y2=4.795
r81 (  26 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.25 //x2=1.405 //y2=1.405
r82 (  25 39 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.905 //x2=1.405 //y2=0.75
r83 (  25 26 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.905 //x2=1.445 //y2=1.25
r84 (  24 33 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=1.09 //y=4.795 //x2=0.955 //y2=4.795
r85 (  23 27 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.375 //y=4.795 //x2=1.45 //y2=4.87
r86 (  23 24 ) resistor r=146.138 //w=0.094 //l=0.285 //layer=ply \
 //thickness=0.18 //x=1.375 //y=4.795 //x2=1.09 //y2=4.795
r87 (  21 38 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.405 //x2=0.955 //y2=1.405
r88 (  20 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.405 //x2=1.405 //y2=1.405
r89 (  19 37 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.75 //x2=0.955 //y2=0.75
r90 (  18 39 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.75 //x2=1.405 //y2=0.75
r91 (  18 19 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.75 //x2=1.07 //y2=0.75
r92 (  14 36 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r93 (  13 38 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.56 //x2=0.955 //y2=1.405
r94 (  13 14 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.56 //x2=0.915 //y2=1.915
r95 (  12 38 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.25 //x2=0.955 //y2=1.405
r96 (  11 37 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.905 //x2=0.955 //y2=0.75
r97 (  11 12 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.905 //x2=0.915 //y2=1.25
r98 (  10 27 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.025 //x2=1.45 //y2=4.87
r99 (  9 34 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.025 //x2=1.01 //y2=4.87
r100 (  8 20 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.405 //x2=1.29 //y2=1.405
r101 (  8 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.405 //x2=1.07 //y2=1.405
r102 (  6 31 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.955 //y=4.705 //x2=0.955 //y2=4.705
r103 (  6 7 ) resistor r=7.81102 //w=0.254 //l=0.155 //layer=li \
 //thickness=0.1 //x=0.955 //y=4.705 //x2=1.11 //y2=4.705
r104 (  3 36 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r105 (  1 7 ) resistor r=3.23951 //w=0.254 //l=0.165 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.54 //x2=1.11 //y2=4.705
r106 (  1 3 ) resistor r=168.385 //w=0.187 //l=2.46 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.54 //x2=1.11 //y2=2.08
ends PM_NOR3X1_PCELL\%noxref_3

subckt PM_NOR3X1_PCELL\%noxref_4 ( 1 3 7 8 9 10 11 12 17 19 21 27 28 30 31 34 )
c80 ( 34 0 ) capacitor c=0.0366246f //x=1.885 //y=4.705
c81 ( 31 0 ) capacitor c=0.0260062f //x=1.85 //y=1.915
c82 ( 30 0 ) capacitor c=0.0407292f //x=1.85 //y=2.08
c83 ( 28 0 ) capacitor c=0.0170937f //x=2.415 //y=1.255
c84 ( 27 0 ) capacitor c=0.0176605f //x=2.415 //y=0.905
c85 ( 21 0 ) capacitor c=0.0305703f //x=2.26 //y=1.405
c86 ( 19 0 ) capacitor c=0.0157804f //x=2.26 //y=0.75
c87 ( 17 0 ) capacitor c=0.0337811f //x=2.255 //y=4.795
c88 ( 12 0 ) capacitor c=0.0189312f //x=1.885 //y=1.56
c89 ( 11 0 ) capacitor c=0.0169608f //x=1.885 //y=1.255
c90 ( 10 0 ) capacitor c=0.0176782f //x=1.885 //y=0.905
c91 ( 9 0 ) capacitor c=0.13968f //x=2.33 //y=6.025
c92 ( 8 0 ) capacitor c=0.110232f //x=1.89 //y=6.025
c93 ( 3 0 ) capacitor c=0.092194f //x=1.85 //y=2.08
c94 ( 1 0 ) capacitor c=0.00580576f //x=1.85 //y=4.54
r95 (  36 37 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.885 //y=4.795 //x2=1.885 //y2=4.87
r96 (  34 36 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.885 //y=4.705 //x2=1.885 //y2=4.795
r97 (  30 31 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r98 (  28 41 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.255 //x2=2.415 //y2=1.367
r99 (  27 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r100 (  27 28 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.255
r101 (  22 39 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r102 (  21 41 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.415 //y2=1.367
r103 (  20 38 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r104 (  19 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r105 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r106 (  18 36 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.02 //y=4.795 //x2=1.885 //y2=4.795
r107 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.795 //x2=2.33 //y2=4.87
r108 (  17 18 ) resistor r=120.5 //w=0.094 //l=0.235 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.795 //x2=2.02 //y2=4.795
r109 (  12 39 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r110 (  12 31 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r111 (  11 39 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.255 //x2=1.925 //y2=1.405
r112 (  10 38 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r113 (  10 11 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.255
r114 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.025 //x2=2.33 //y2=4.87
r115 (  8 37 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.025 //x2=1.89 //y2=4.87
r116 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r117 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r118 (  6 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.885 //y=4.705 //x2=1.885 //y2=4.705
r119 (  3 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r120 (  1 6 ) resistor r=11.332 //w=0.189 //l=0.173292 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.54 //x2=1.867 //y2=4.705
r121 (  1 3 ) resistor r=168.385 //w=0.187 //l=2.46 //layer=li //thickness=0.1 \
 //x=1.85 //y=4.54 //x2=1.85 //y2=2.08
ends PM_NOR3X1_PCELL\%noxref_4

subckt PM_NOR3X1_PCELL\%noxref_5 ( 7 8 15 16 23 24 25 )
c43 ( 25 0 ) capacitor c=0.0202519f //x=2.405 //y=5.025
c44 ( 24 0 ) capacitor c=0.0185379f //x=1.525 //y=5.025
c45 ( 23 0 ) capacitor c=0.0408953f //x=0.655 //y=5.025
c46 ( 16 0 ) capacitor c=0.00193672f //x=1.755 //y=6.91
c47 ( 15 0 ) capacitor c=0.0126253f //x=2.465 //y=6.91
c48 ( 8 0 ) capacitor c=0.00844339f //x=0.875 //y=5.21
c49 ( 7 0 ) capacitor c=0.0252644f //x=1.585 //y=5.21
r50 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.55 //y=6.825 //x2=2.55 //y2=6.74
r51 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.465 //y=6.91 //x2=2.55 //y2=6.825
r52 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.465 //y=6.91 //x2=1.755 //y2=6.91
r53 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.67 //y=6.825 //x2=1.755 //y2=6.91
r54 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.67 //y=6.825 //x2=1.67 //y2=6.4
r55 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.67 //y=5.295 //x2=1.67 //y2=5.72
r56 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.585 //y=5.21 //x2=1.67 //y2=5.295
r57 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=1.585 //y=5.21 //x2=0.875 //y2=5.21
r58 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=0.79 //y=5.295 //x2=0.875 //y2=5.21
r59 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=0.79 //y=5.295 //x2=0.79 //y2=5.72
ends PM_NOR3X1_PCELL\%noxref_5

subckt PM_NOR3X1_PCELL\%noxref_6 ( 2 7 8 9 10 11 12 13 14 16 24 25 26 31 35 )
c67 ( 41 0 ) capacitor c=0.011077f //x=3.37 //y=4.795
c68 ( 35 0 ) capacitor c=0.0431417f //x=2.96 //y=4.705
c69 ( 31 0 ) capacitor c=0.0492905f //x=2.855 //y=2.08
c70 ( 26 0 ) capacitor c=0.0363749f //x=3.735 //y=4.795
c71 ( 25 0 ) capacitor c=0.0237734f //x=3.385 //y=1.255
c72 ( 24 0 ) capacitor c=0.0191782f //x=3.385 //y=0.905
c73 ( 19 0 ) capacitor c=0.0202859f //x=3.295 //y=4.795
c74 ( 16 0 ) capacitor c=0.033152f //x=3.23 //y=1.405
c75 ( 14 0 ) capacitor c=0.0157803f //x=3.23 //y=0.75
c76 ( 13 0 ) capacitor c=0.0280515f //x=2.855 //y=1.915
c77 ( 12 0 ) capacitor c=0.0189445f //x=2.855 //y=1.56
c78 ( 11 0 ) capacitor c=0.0170937f //x=2.855 //y=1.255
c79 ( 10 0 ) capacitor c=0.0185081f //x=2.855 //y=0.905
c80 ( 9 0 ) capacitor c=0.154473f //x=3.81 //y=6.025
c81 ( 8 0 ) capacitor c=0.139411f //x=3.37 //y=6.025
c82 ( 2 0 ) capacitor c=0.0965855f //x=2.96 //y=2.08
r83 (  35 37 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.96 //y=4.705 //x2=2.96 //y2=4.795
r84 (  31 33 ) resistor r=16.5934 //w=0.305 //l=0.105 //layer=ply \
 //thickness=0.18 //x=2.855 //y=2.08 //x2=2.96 //y2=2.08
r85 (  27 41 ) resistor r=20.4101 //w=0.15 //l=0.075 //layer=ply \
 //thickness=0.18 //x=3.445 //y=4.795 //x2=3.37 //y2=4.795
r86 (  26 28 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=3.735 //y=4.795 //x2=3.81 //y2=4.87
r87 (  26 27 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=3.735 //y=4.795 //x2=3.445 //y2=4.795
r88 (  25 43 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=3.385 //y=1.255 //x2=3.385 //y2=1.367
r89 (  24 42 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.385 //y=0.905 //x2=3.345 //y2=0.75
r90 (  24 25 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=3.385 //y=0.905 //x2=3.385 //y2=1.255
r91 (  21 41 ) resistor r=5.30422 //w=0.3 //l=0.075 //layer=ply \
 //thickness=0.18 //x=3.37 //y=4.87 //x2=3.37 //y2=4.795
r92 (  20 37 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=3.095 //y=4.795 //x2=2.96 //y2=4.795
r93 (  19 41 ) resistor r=20.4101 //w=0.15 //l=0.075 //layer=ply \
 //thickness=0.18 //x=3.295 //y=4.795 //x2=3.37 //y2=4.795
r94 (  19 20 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=3.295 //y=4.795 //x2=3.095 //y2=4.795
r95 (  17 40 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.01 //y=1.405 //x2=2.895 //y2=1.405
r96 (  16 43 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=3.23 //y=1.405 //x2=3.385 //y2=1.367
r97 (  15 39 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.01 //y=0.75 //x2=2.895 //y2=0.75
r98 (  14 42 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.23 //y=0.75 //x2=3.345 //y2=0.75
r99 (  14 15 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.23 //y=0.75 //x2=3.01 //y2=0.75
r100 (  13 31 ) resistor r=19.3576 //w=0.305 //l=0.165 //layer=ply \
 //thickness=0.18 //x=2.855 //y=1.915 //x2=2.855 //y2=2.08
r101 (  12 40 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.855 //y=1.56 //x2=2.895 //y2=1.405
r102 (  12 13 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=2.855 //y=1.56 //x2=2.855 //y2=1.915
r103 (  11 40 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=2.855 //y=1.255 //x2=2.895 //y2=1.405
r104 (  10 39 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.855 //y=0.905 //x2=2.895 //y2=0.75
r105 (  10 11 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=2.855 //y=0.905 //x2=2.855 //y2=1.255
r106 (  9 28 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.81 //y=6.025 //x2=3.81 //y2=4.87
r107 (  8 21 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.37 //y=6.025 //x2=3.37 //y2=4.87
r108 (  7 16 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.12 //y=1.405 //x2=3.23 //y2=1.405
r109 (  7 17 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.12 //y=1.405 //x2=3.01 //y2=1.405
r110 (  5 35 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.96 //y=4.705 //x2=2.96 //y2=4.705
r111 (  2 33 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.96 //y=2.08 //x2=2.96 //y2=2.08
r112 (  2 5 ) resistor r=179.679 //w=0.187 //l=2.625 //layer=li \
 //thickness=0.1 //x=2.96 //y=2.08 //x2=2.96 //y2=4.705
ends PM_NOR3X1_PCELL\%noxref_6

subckt PM_NOR3X1_PCELL\%noxref_7 ( 5 6 11 17 24 26 29 31 32 33 37 )
c83 ( 37 0 ) capacitor c=0.0159625f //x=3.445 //y=5.025
c84 ( 33 0 ) capacitor c=0.00969064f //x=2.93 //y=0.905
c85 ( 32 0 ) capacitor c=0.00860823f //x=1.96 //y=0.905
c86 ( 31 0 ) capacitor c=0.007684f //x=0.99 //y=0.905
c87 ( 29 0 ) capacitor c=0.00603509f //x=3.7 //y=5.21
c88 ( 26 0 ) capacitor c=0.00544799f //x=3.12 //y=1.655
c89 ( 25 0 ) capacitor c=0.00710337f //x=2.15 //y=1.655
c90 ( 24 0 ) capacitor c=0.14166f //x=3.7 //y=5.125
c91 ( 17 0 ) capacitor c=0.0260487f //x=3.615 //y=1.655
c92 ( 11 0 ) capacitor c=0.0281501f //x=3.035 //y=1.655
c93 ( 6 0 ) capacitor c=0.00277859f //x=1.265 //y=1.655
c94 ( 5 0 ) capacitor c=0.0280953f //x=2.065 //y=1.655
r95 (  27 29 ) resistor r=7.52941 //w=0.187 //l=0.11 //layer=li \
 //thickness=0.1 //x=3.59 //y=5.21 //x2=3.7 //y2=5.21
r96 (  24 29 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.7 //y=5.125 //x2=3.7 //y2=5.21
r97 (  23 24 ) resistor r=231.701 //w=0.187 //l=3.385 //layer=li \
 //thickness=0.1 //x=3.7 //y=1.74 //x2=3.7 //y2=5.125
r98 (  19 27 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.59 //y=5.295 //x2=3.59 //y2=5.21
r99 (  19 37 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=3.59 //y=5.295 //x2=3.59 //y2=6.06
r100 (  18 26 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.205 //y=1.655 //x2=3.12 //y2=1.655
r101 (  17 23 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.615 //y=1.655 //x2=3.7 //y2=1.74
r102 (  17 18 ) resistor r=28.0642 //w=0.187 //l=0.41 //layer=li \
 //thickness=0.1 //x=3.615 //y=1.655 //x2=3.205 //y2=1.655
r103 (  13 26 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.12 //y=1.57 //x2=3.12 //y2=1.655
r104 (  13 33 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=3.12 //y=1.57 //x2=3.12 //y2=1
r105 (  12 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.235 //y=1.655 //x2=2.15 //y2=1.655
r106 (  11 26 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.035 //y=1.655 //x2=3.12 //y2=1.655
r107 (  11 12 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li \
 //thickness=0.1 //x=3.035 //y=1.655 //x2=2.235 //y2=1.655
r108 (  7 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1.655
r109 (  7 32 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r110 (  5 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.065 //y=1.655 //x2=2.15 //y2=1.655
r111 (  5 6 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li //thickness=0.1 \
 //x=2.065 //y=1.655 //x2=1.265 //y2=1.655
r112 (  1 6 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.18 //y=1.57 //x2=1.265 //y2=1.655
r113 (  1 31 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=1.18 //y=1.57 //x2=1.18 //y2=1
ends PM_NOR3X1_PCELL\%noxref_7

subckt PM_NOR3X1_PCELL\%noxref_8 ( 7 8 15 16 23 24 25 )
c37 ( 25 0 ) capacitor c=0.0362595f //x=3.885 //y=5.025
c38 ( 24 0 ) capacitor c=0.023843f //x=3.015 //y=5.025
c39 ( 23 0 ) capacitor c=0.0167469f //x=1.965 //y=5.025
c40 ( 16 0 ) capacitor c=0.00239377f //x=3.235 //y=6.91
c41 ( 15 0 ) capacitor c=0.0145111f //x=3.945 //y=6.91
c42 ( 8 0 ) capacitor c=0.00499653f //x=2.195 //y=5.21
c43 ( 7 0 ) capacitor c=0.0417267f //x=3.065 //y=5.21
r44 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.03 //y=6.825 //x2=4.03 //y2=6.74
r45 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.945 //y=6.91 //x2=4.03 //y2=6.825
r46 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.945 //y=6.91 //x2=3.235 //y2=6.91
r47 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.15 //y=6.825 //x2=3.235 //y2=6.91
r48 (  10 24 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.15 //y=6.825 //x2=3.15 //y2=6.74
r49 (  9 24 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=3.15 //y=5.295 //x2=3.15 //y2=6.06
r50 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.065 //y=5.21 //x2=3.15 //y2=5.295
r51 (  7 8 ) resistor r=59.5508 //w=0.187 //l=0.87 //layer=li //thickness=0.1 \
 //x=3.065 //y=5.21 //x2=2.195 //y2=5.21
r52 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.295 //x2=2.195 //y2=5.21
r53 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.295 //x2=2.11 //y2=5.72
ends PM_NOR3X1_PCELL\%noxref_8

