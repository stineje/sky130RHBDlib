// File: xor2X1_pcell.spi.XOR2X1_PCELL.pxi
// Created: Tue Oct 15 16:01:28 2024
// 
simulator lang=spectre
x_PM_XOR2X1_PCELL\%noxref_1 ( N_noxref_1_c_6_p N_noxref_1_c_11_p \
 N_noxref_1_c_20_p N_noxref_1_c_136_p N_noxref_1_c_36_p N_noxref_1_c_23_p \
 N_noxref_1_c_29_p N_noxref_1_c_39_p N_noxref_1_c_40_p N_noxref_1_c_96_p \
 N_noxref_1_c_156_p N_noxref_1_c_77_p N_noxref_1_c_104_p N_noxref_1_c_1_p \
 N_noxref_1_c_2_p N_noxref_1_c_3_p N_noxref_1_c_4_p N_noxref_1_c_5_p \
 N_noxref_1_M0_noxref_s N_noxref_1_M1_noxref_d N_noxref_1_M3_noxref_d \
 N_noxref_1_M5_noxref_s )  PM_XOR2X1_PCELL\%noxref_1
x_PM_XOR2X1_PCELL\%noxref_2 ( N_noxref_2_c_171_p N_noxref_2_c_172_p \
 N_noxref_2_c_173_p N_noxref_2_c_174_p N_noxref_2_c_193_p N_noxref_2_c_234_p \
 N_noxref_2_c_208_p N_noxref_2_c_257_p N_noxref_2_c_244_p N_noxref_2_c_166_n \
 N_noxref_2_c_167_n N_noxref_2_c_168_n N_noxref_2_c_169_n N_noxref_2_c_170_n \
 N_noxref_2_M6_noxref_s N_noxref_2_M7_noxref_d N_noxref_2_M8_noxref_d \
 N_noxref_2_M12_noxref_d N_noxref_2_M16_noxref_s N_noxref_2_M17_noxref_d )  \
 PM_XOR2X1_PCELL\%noxref_2
x_PM_XOR2X1_PCELL\%noxref_3 ( N_noxref_3_c_322_n N_noxref_3_c_324_n \
 N_noxref_3_c_326_n N_noxref_3_c_331_n N_noxref_3_M0_noxref_g \
 N_noxref_3_M1_noxref_g N_noxref_3_M6_noxref_g N_noxref_3_M7_noxref_g \
 N_noxref_3_M8_noxref_g N_noxref_3_M9_noxref_g N_noxref_3_c_332_n \
 N_noxref_3_c_398_p N_noxref_3_c_399_p N_noxref_3_c_334_n N_noxref_3_c_375_n \
 N_noxref_3_c_376_n N_noxref_3_c_335_n N_noxref_3_c_385_p N_noxref_3_c_336_n \
 N_noxref_3_c_338_n N_noxref_3_c_339_n N_noxref_3_c_341_n N_noxref_3_c_428_p \
 N_noxref_3_c_342_n N_noxref_3_c_343_n N_noxref_3_c_344_n N_noxref_3_c_345_n \
 N_noxref_3_c_347_n N_noxref_3_c_348_n N_noxref_3_c_378_n )  \
 PM_XOR2X1_PCELL\%noxref_3
x_PM_XOR2X1_PCELL\%noxref_4 ( N_noxref_4_c_455_n N_noxref_4_c_464_n \
 N_noxref_4_c_467_n N_noxref_4_c_506_n N_noxref_4_c_482_n N_noxref_4_c_485_n \
 N_noxref_4_c_470_n N_noxref_4_c_473_n N_noxref_4_M4_noxref_g \
 N_noxref_4_M14_noxref_g N_noxref_4_M15_noxref_g N_noxref_4_c_555_p \
 N_noxref_4_c_556_p N_noxref_4_c_557_p N_noxref_4_c_545_p N_noxref_4_c_559_p \
 N_noxref_4_c_546_p N_noxref_4_c_561_p N_noxref_4_c_547_p N_noxref_4_c_540_p \
 N_noxref_4_M0_noxref_d N_noxref_4_M6_noxref_d )  PM_XOR2X1_PCELL\%noxref_4
x_PM_XOR2X1_PCELL\%noxref_5 ( N_noxref_5_c_653_n N_noxref_5_c_651_n \
 N_noxref_5_c_636_n N_noxref_5_c_638_n N_noxref_5_c_624_n N_noxref_5_c_659_n \
 N_noxref_5_c_625_n N_noxref_5_c_641_n N_noxref_5_c_643_n N_noxref_5_c_626_n \
 N_noxref_5_c_672_n N_noxref_5_c_628_n N_noxref_5_M2_noxref_d \
 N_noxref_5_M4_noxref_d N_noxref_5_M10_noxref_d N_noxref_5_M14_noxref_d )  \
 PM_XOR2X1_PCELL\%noxref_5
x_PM_XOR2X1_PCELL\%noxref_6 ( N_noxref_6_c_794_n N_noxref_6_c_799_n \
 N_noxref_6_c_831_n N_noxref_6_c_833_n N_noxref_6_c_800_n N_noxref_6_c_773_n \
 N_noxref_6_c_774_n N_noxref_6_c_775_n N_noxref_6_c_776_n N_noxref_6_c_804_n \
 N_noxref_6_c_805_n N_noxref_6_M3_noxref_g N_noxref_6_M10_noxref_g \
 N_noxref_6_M11_noxref_g N_noxref_6_c_780_n N_noxref_6_c_782_n \
 N_noxref_6_c_783_n N_noxref_6_c_784_n N_noxref_6_c_785_n N_noxref_6_c_786_n \
 N_noxref_6_c_787_n N_noxref_6_c_789_n N_noxref_6_c_826_n \
 N_noxref_6_M5_noxref_d N_noxref_6_M16_noxref_d )  PM_XOR2X1_PCELL\%noxref_6
x_PM_XOR2X1_PCELL\%noxref_7 ( N_noxref_7_c_938_n N_noxref_7_c_991_n \
 N_noxref_7_c_962_n N_noxref_7_c_970_n N_noxref_7_c_945_n N_noxref_7_c_972_n \
 N_noxref_7_c_947_n N_noxref_7_M2_noxref_g N_noxref_7_M5_noxref_g \
 N_noxref_7_M12_noxref_g N_noxref_7_M13_noxref_g N_noxref_7_M16_noxref_g \
 N_noxref_7_M17_noxref_g N_noxref_7_c_994_n N_noxref_7_c_997_n \
 N_noxref_7_c_999_n N_noxref_7_c_1002_n N_noxref_7_c_1045_n \
 N_noxref_7_c_1046_n N_noxref_7_c_1004_n N_noxref_7_c_1005_n \
 N_noxref_7_c_952_n N_noxref_7_c_954_n N_noxref_7_c_1081_n N_noxref_7_c_987_n \
 N_noxref_7_c_955_n N_noxref_7_c_1085_n N_noxref_7_c_988_n N_noxref_7_c_956_n \
 N_noxref_7_c_1089_n N_noxref_7_c_1090_n N_noxref_7_c_958_n N_noxref_7_c_990_n \
 N_noxref_7_c_959_n )  PM_XOR2X1_PCELL\%noxref_7
x_PM_XOR2X1_PCELL\%noxref_8 ( N_noxref_8_c_1111_n N_noxref_8_c_1116_n \
 N_noxref_8_c_1118_n N_noxref_8_c_1119_n N_noxref_8_M8_noxref_s \
 N_noxref_8_M9_noxref_d N_noxref_8_M11_noxref_d )  PM_XOR2X1_PCELL\%noxref_8
x_PM_XOR2X1_PCELL\%noxref_9 ( N_noxref_9_c_1151_n N_noxref_9_c_1152_n \
 N_noxref_9_c_1156_n N_noxref_9_c_1160_n N_noxref_9_c_1161_n \
 N_noxref_9_c_1164_n N_noxref_9_M1_noxref_s )  PM_XOR2X1_PCELL\%noxref_9
x_PM_XOR2X1_PCELL\%noxref_10 ( N_noxref_10_c_1203_n N_noxref_10_c_1208_n \
 N_noxref_10_c_1209_n N_noxref_10_c_1210_n N_noxref_10_M12_noxref_s \
 N_noxref_10_M13_noxref_d N_noxref_10_M15_noxref_d )  PM_XOR2X1_PCELL\%noxref_10
x_PM_XOR2X1_PCELL\%noxref_11 ( N_noxref_11_c_1270_n N_noxref_11_c_1246_n \
 N_noxref_11_c_1250_n N_noxref_11_c_1254_n N_noxref_11_c_1255_n \
 N_noxref_11_c_1258_n N_noxref_11_M3_noxref_s )  PM_XOR2X1_PCELL\%noxref_11
cc_1 ( N_noxref_1_c_1_p N_noxref_2_c_166_n ) capacitor c=0.00989031f //x=0.63 \
 //y=0 //x2=0.74 //y2=7.4
cc_2 ( N_noxref_1_c_2_p N_noxref_2_c_167_n ) capacitor c=0.00582097f //x=2.22 \
 //y=0 //x2=2.22 //y2=7.4
cc_3 ( N_noxref_1_c_3_p N_noxref_2_c_168_n ) capacitor c=0.0057235f //x=5.55 \
 //y=0 //x2=5.55 //y2=7.4
cc_4 ( N_noxref_1_c_4_p N_noxref_2_c_169_n ) capacitor c=0.00478842f //x=8.88 \
 //y=0 //x2=8.88 //y2=7.4
cc_5 ( N_noxref_1_c_5_p N_noxref_2_c_170_n ) capacitor c=0.00989031f //x=10.47 \
 //y=0 //x2=10.36 //y2=7.4
cc_6 ( N_noxref_1_c_6_p N_noxref_3_c_322_n ) capacitor c=0.00375415f //x=10.36 \
 //y=0 //x2=3.215 //y2=4.07
cc_7 ( N_noxref_1_c_2_p N_noxref_3_c_322_n ) capacitor c=0.00249386f //x=2.22 \
 //y=0 //x2=3.215 //y2=4.07
cc_8 ( N_noxref_1_c_6_p N_noxref_3_c_324_n ) capacitor c=0.00155455f //x=10.36 \
 //y=0 //x2=0.855 //y2=4.07
cc_9 ( N_noxref_1_M0_noxref_s N_noxref_3_c_324_n ) capacitor c=5.91312e-19 \
 //x=0.495 //y=0.37 //x2=0.855 //y2=4.07
cc_10 ( N_noxref_1_c_6_p N_noxref_3_c_326_n ) capacitor c=0.00187124f \
 //x=10.36 //y=0 //x2=0.74 //y2=2.085
cc_11 ( N_noxref_1_c_11_p N_noxref_3_c_326_n ) capacitor c=8.01092e-19 \
 //x=1.03 //y=0.535 //x2=0.74 //y2=2.085
cc_12 ( N_noxref_1_c_1_p N_noxref_3_c_326_n ) capacitor c=0.028767f //x=0.63 \
 //y=0 //x2=0.74 //y2=2.085
cc_13 ( N_noxref_1_c_2_p N_noxref_3_c_326_n ) capacitor c=0.00133655f //x=2.22 \
 //y=0 //x2=0.74 //y2=2.085
cc_14 ( N_noxref_1_M0_noxref_s N_noxref_3_c_326_n ) capacitor c=0.0110965f \
 //x=0.495 //y=0.37 //x2=0.74 //y2=2.085
cc_15 ( N_noxref_1_c_2_p N_noxref_3_c_331_n ) capacitor c=0.0151398f //x=2.22 \
 //y=0 //x2=3.33 //y2=2.085
cc_16 ( N_noxref_1_c_11_p N_noxref_3_c_332_n ) capacitor c=0.0120496f //x=1.03 \
 //y=0.535 //x2=0.85 //y2=0.91
cc_17 ( N_noxref_1_M0_noxref_s N_noxref_3_c_332_n ) capacitor c=0.0316686f \
 //x=0.495 //y=0.37 //x2=0.85 //y2=0.91
cc_18 ( N_noxref_1_c_1_p N_noxref_3_c_334_n ) capacitor c=0.0124051f //x=0.63 \
 //y=0 //x2=0.85 //y2=1.92
cc_19 ( N_noxref_1_M0_noxref_s N_noxref_3_c_335_n ) capacitor c=0.00483274f \
 //x=0.495 //y=0.37 //x2=1.225 //y2=0.755
cc_20 ( N_noxref_1_c_20_p N_noxref_3_c_336_n ) capacitor c=0.0118602f \
 //x=1.515 //y=0.535 //x2=1.38 //y2=0.91
cc_21 ( N_noxref_1_M0_noxref_s N_noxref_3_c_336_n ) capacitor c=0.0143355f \
 //x=0.495 //y=0.37 //x2=1.38 //y2=0.91
cc_22 ( N_noxref_1_M0_noxref_s N_noxref_3_c_338_n ) capacitor c=0.0074042f \
 //x=0.495 //y=0.37 //x2=1.38 //y2=1.255
cc_23 ( N_noxref_1_c_23_p N_noxref_3_c_339_n ) capacitor c=0.00134217f \
 //x=3.315 //y=0 //x2=3.135 //y2=0.87
cc_24 ( N_noxref_1_M1_noxref_d N_noxref_3_c_339_n ) capacitor c=0.00220047f \
 //x=3.21 //y=0.87 //x2=3.135 //y2=0.87
cc_25 ( N_noxref_1_M1_noxref_d N_noxref_3_c_341_n ) capacitor c=0.00255985f \
 //x=3.21 //y=0.87 //x2=3.135 //y2=1.215
cc_26 ( N_noxref_1_c_2_p N_noxref_3_c_342_n ) capacitor c=0.0114882f //x=2.22 \
 //y=0 //x2=3.135 //y2=1.92
cc_27 ( N_noxref_1_M1_noxref_d N_noxref_3_c_343_n ) capacitor c=0.013135f \
 //x=3.21 //y=0.87 //x2=3.51 //y2=0.715
cc_28 ( N_noxref_1_M1_noxref_d N_noxref_3_c_344_n ) capacitor c=0.00193136f \
 //x=3.21 //y=0.87 //x2=3.51 //y2=1.37
cc_29 ( N_noxref_1_c_29_p N_noxref_3_c_345_n ) capacitor c=0.00129817f \
 //x=5.38 //y=0 //x2=3.665 //y2=0.87
cc_30 ( N_noxref_1_M1_noxref_d N_noxref_3_c_345_n ) capacitor c=0.00257848f \
 //x=3.21 //y=0.87 //x2=3.665 //y2=0.87
cc_31 ( N_noxref_1_M1_noxref_d N_noxref_3_c_347_n ) capacitor c=0.00255985f \
 //x=3.21 //y=0.87 //x2=3.665 //y2=1.215
cc_32 ( N_noxref_1_c_11_p N_noxref_3_c_348_n ) capacitor c=2.1838e-19 //x=1.03 \
 //y=0.535 //x2=0.74 //y2=2.085
cc_33 ( N_noxref_1_c_1_p N_noxref_3_c_348_n ) capacitor c=0.0108179f //x=0.63 \
 //y=0 //x2=0.74 //y2=2.085
cc_34 ( N_noxref_1_M0_noxref_s N_noxref_3_c_348_n ) capacitor c=0.00655738f \
 //x=0.495 //y=0.37 //x2=0.74 //y2=2.085
cc_35 ( N_noxref_1_c_6_p N_noxref_4_c_455_n ) capacitor c=0.0533505f //x=10.36 \
 //y=0 //x2=7.655 //y2=2.59
cc_36 ( N_noxref_1_c_36_p N_noxref_4_c_455_n ) capacitor c=0.0015622f //x=2.05 \
 //y=0 //x2=7.655 //y2=2.59
cc_37 ( N_noxref_1_c_23_p N_noxref_4_c_455_n ) capacitor c=0.00281115f \
 //x=3.315 //y=0 //x2=7.655 //y2=2.59
cc_38 ( N_noxref_1_c_29_p N_noxref_4_c_455_n ) capacitor c=0.00346399f \
 //x=5.38 //y=0 //x2=7.655 //y2=2.59
cc_39 ( N_noxref_1_c_39_p N_noxref_4_c_455_n ) capacitor c=0.00281115f \
 //x=6.645 //y=0 //x2=7.655 //y2=2.59
cc_40 ( N_noxref_1_c_40_p N_noxref_4_c_455_n ) capacitor c=9.27524e-19 \
 //x=8.71 //y=0 //x2=7.655 //y2=2.59
cc_41 ( N_noxref_1_c_2_p N_noxref_4_c_455_n ) capacitor c=0.038878f //x=2.22 \
 //y=0 //x2=7.655 //y2=2.59
cc_42 ( N_noxref_1_c_3_p N_noxref_4_c_455_n ) capacitor c=0.0338055f //x=5.55 \
 //y=0 //x2=7.655 //y2=2.59
cc_43 ( N_noxref_1_M0_noxref_s N_noxref_4_c_455_n ) capacitor c=0.00248261f \
 //x=0.495 //y=0.37 //x2=7.655 //y2=2.59
cc_44 ( N_noxref_1_c_6_p N_noxref_4_c_464_n ) capacitor c=0.00231366f \
 //x=10.36 //y=0 //x2=1.595 //y2=2.59
cc_45 ( N_noxref_1_c_2_p N_noxref_4_c_464_n ) capacitor c=0.00209945f //x=2.22 \
 //y=0 //x2=1.595 //y2=2.59
cc_46 ( N_noxref_1_M0_noxref_s N_noxref_4_c_464_n ) capacitor c=0.00120637f \
 //x=0.495 //y=0.37 //x2=1.595 //y2=2.59
cc_47 ( N_noxref_1_c_6_p N_noxref_4_c_467_n ) capacitor c=0.00129718f \
 //x=10.36 //y=0 //x2=1.395 //y2=2.08
cc_48 ( N_noxref_1_c_2_p N_noxref_4_c_467_n ) capacitor c=0.0263587f //x=2.22 \
 //y=0 //x2=1.395 //y2=2.08
cc_49 ( N_noxref_1_M0_noxref_s N_noxref_4_c_467_n ) capacitor c=0.00949589f \
 //x=0.495 //y=0.37 //x2=1.395 //y2=2.08
cc_50 ( N_noxref_1_c_1_p N_noxref_4_c_470_n ) capacitor c=9.71e-19 //x=0.63 \
 //y=0 //x2=1.48 //y2=2.59
cc_51 ( N_noxref_1_c_2_p N_noxref_4_c_470_n ) capacitor c=5.56859e-19 //x=2.22 \
 //y=0 //x2=1.48 //y2=2.59
cc_52 ( N_noxref_1_M0_noxref_s N_noxref_4_c_470_n ) capacitor c=2.30929e-19 \
 //x=0.495 //y=0.37 //x2=1.48 //y2=2.59
cc_53 ( N_noxref_1_c_3_p N_noxref_4_c_473_n ) capacitor c=6.8921e-19 //x=5.55 \
 //y=0 //x2=7.77 //y2=2.085
cc_54 ( N_noxref_1_c_4_p N_noxref_4_c_473_n ) capacitor c=0.00183906f //x=8.88 \
 //y=0 //x2=7.77 //y2=2.085
cc_55 ( N_noxref_1_c_6_p N_noxref_4_M0_noxref_d ) capacitor c=0.00136354f \
 //x=10.36 //y=0 //x2=0.925 //y2=0.91
cc_56 ( N_noxref_1_c_11_p N_noxref_4_M0_noxref_d ) capacitor c=0.0151737f \
 //x=1.03 //y=0.535 //x2=0.925 //y2=0.91
cc_57 ( N_noxref_1_c_1_p N_noxref_4_M0_noxref_d ) capacitor c=0.0094373f \
 //x=0.63 //y=0 //x2=0.925 //y2=0.91
cc_58 ( N_noxref_1_c_2_p N_noxref_4_M0_noxref_d ) capacitor c=0.00949341f \
 //x=2.22 //y=0 //x2=0.925 //y2=0.91
cc_59 ( N_noxref_1_c_5_p N_noxref_4_M0_noxref_d ) capacitor c=2.29264e-19 \
 //x=10.47 //y=0 //x2=0.925 //y2=0.91
cc_60 ( N_noxref_1_M0_noxref_s N_noxref_4_M0_noxref_d ) capacitor c=0.076995f \
 //x=0.495 //y=0.37 //x2=0.925 //y2=0.91
cc_61 ( N_noxref_1_c_3_p N_noxref_5_c_624_n ) capacitor c=0.0428968f //x=5.55 \
 //y=0 //x2=4.725 //y2=1.655
cc_62 ( N_noxref_1_c_2_p N_noxref_5_c_625_n ) capacitor c=0.00105873f //x=2.22 \
 //y=0 //x2=4.81 //y2=3.7
cc_63 ( N_noxref_1_c_4_p N_noxref_5_c_626_n ) capacitor c=0.0446773f //x=8.88 \
 //y=0 //x2=8.055 //y2=1.655
cc_64 ( N_noxref_1_M5_noxref_s N_noxref_5_c_626_n ) capacitor c=3.42693e-19 \
 //x=9.375 //y=0.37 //x2=8.055 //y2=1.655
cc_65 ( N_noxref_1_c_3_p N_noxref_5_c_628_n ) capacitor c=0.00100332f //x=5.55 \
 //y=0 //x2=8.14 //y2=3.7
cc_66 ( N_noxref_1_c_2_p N_noxref_5_M2_noxref_d ) capacitor c=8.60262e-19 \
 //x=2.22 //y=0 //x2=4.18 //y2=0.91
cc_67 ( N_noxref_1_c_3_p N_noxref_5_M2_noxref_d ) capacitor c=0.00605305f \
 //x=5.55 //y=0 //x2=4.18 //y2=0.91
cc_68 ( N_noxref_1_M1_noxref_d N_noxref_5_M2_noxref_d ) capacitor \
 c=0.00143464f //x=3.21 //y=0.87 //x2=4.18 //y2=0.91
cc_69 ( N_noxref_1_c_3_p N_noxref_5_M4_noxref_d ) capacitor c=8.60262e-19 \
 //x=5.55 //y=0 //x2=7.51 //y2=0.91
cc_70 ( N_noxref_1_c_4_p N_noxref_5_M4_noxref_d ) capacitor c=0.00605305f \
 //x=8.88 //y=0 //x2=7.51 //y2=0.91
cc_71 ( N_noxref_1_M3_noxref_d N_noxref_5_M4_noxref_d ) capacitor \
 c=0.00143464f //x=6.54 //y=0.87 //x2=7.51 //y2=0.91
cc_72 ( N_noxref_1_M5_noxref_s N_noxref_5_M4_noxref_d ) capacitor \
 c=2.07711e-19 //x=9.375 //y=0.37 //x2=7.51 //y2=0.91
cc_73 ( N_noxref_1_c_3_p N_noxref_6_c_773_n ) capacitor c=0.0151475f //x=5.55 \
 //y=0 //x2=6.66 //y2=2.085
cc_74 ( N_noxref_1_c_5_p N_noxref_6_c_774_n ) capacitor c=0.00114558f \
 //x=10.47 //y=0 //x2=9.62 //y2=3.33
cc_75 ( N_noxref_1_M5_noxref_s N_noxref_6_c_775_n ) capacitor c=0.00178356f \
 //x=9.375 //y=0.37 //x2=9.905 //y2=2.08
cc_76 ( N_noxref_1_c_6_p N_noxref_6_c_776_n ) capacitor c=0.00128495f \
 //x=10.36 //y=0 //x2=9.705 //y2=2.08
cc_77 ( N_noxref_1_c_77_p N_noxref_6_c_776_n ) capacitor c=0.00178356f //x=9.9 \
 //y=0.535 //x2=9.705 //y2=2.08
cc_78 ( N_noxref_1_c_4_p N_noxref_6_c_776_n ) capacitor c=0.0291959f //x=8.88 \
 //y=0 //x2=9.705 //y2=2.08
cc_79 ( N_noxref_1_M5_noxref_s N_noxref_6_c_776_n ) capacitor c=0.00610757f \
 //x=9.375 //y=0.37 //x2=9.705 //y2=2.08
cc_80 ( N_noxref_1_c_39_p N_noxref_6_c_780_n ) capacitor c=0.00134217f \
 //x=6.645 //y=0 //x2=6.465 //y2=0.87
cc_81 ( N_noxref_1_M3_noxref_d N_noxref_6_c_780_n ) capacitor c=0.00220047f \
 //x=6.54 //y=0.87 //x2=6.465 //y2=0.87
cc_82 ( N_noxref_1_M3_noxref_d N_noxref_6_c_782_n ) capacitor c=0.00255985f \
 //x=6.54 //y=0.87 //x2=6.465 //y2=1.215
cc_83 ( N_noxref_1_c_3_p N_noxref_6_c_783_n ) capacitor c=0.00176175f //x=5.55 \
 //y=0 //x2=6.465 //y2=1.525
cc_84 ( N_noxref_1_c_3_p N_noxref_6_c_784_n ) capacitor c=0.0114882f //x=5.55 \
 //y=0 //x2=6.465 //y2=1.92
cc_85 ( N_noxref_1_M3_noxref_d N_noxref_6_c_785_n ) capacitor c=0.013135f \
 //x=6.54 //y=0.87 //x2=6.84 //y2=0.715
cc_86 ( N_noxref_1_M3_noxref_d N_noxref_6_c_786_n ) capacitor c=0.00193136f \
 //x=6.54 //y=0.87 //x2=6.84 //y2=1.37
cc_87 ( N_noxref_1_c_40_p N_noxref_6_c_787_n ) capacitor c=0.00129817f \
 //x=8.71 //y=0 //x2=6.995 //y2=0.87
cc_88 ( N_noxref_1_M3_noxref_d N_noxref_6_c_787_n ) capacitor c=0.00257848f \
 //x=6.54 //y=0.87 //x2=6.995 //y2=0.87
cc_89 ( N_noxref_1_M3_noxref_d N_noxref_6_c_789_n ) capacitor c=0.00255985f \
 //x=6.54 //y=0.87 //x2=6.995 //y2=1.215
cc_90 ( N_noxref_1_c_6_p N_noxref_6_M5_noxref_d ) capacitor c=0.00124113f \
 //x=10.36 //y=0 //x2=9.795 //y2=0.91
cc_91 ( N_noxref_1_c_4_p N_noxref_6_M5_noxref_d ) capacitor c=0.00945919f \
 //x=8.88 //y=0 //x2=9.795 //y2=0.91
cc_92 ( N_noxref_1_c_5_p N_noxref_6_M5_noxref_d ) capacitor c=0.00966656f \
 //x=10.47 //y=0 //x2=9.795 //y2=0.91
cc_93 ( N_noxref_1_M5_noxref_s N_noxref_6_M5_noxref_d ) capacitor c=0.0920431f \
 //x=9.375 //y=0.37 //x2=9.795 //y2=0.91
cc_94 ( N_noxref_1_c_6_p N_noxref_7_c_938_n ) capacitor c=0.0344763f //x=10.36 \
 //y=0 //x2=10.245 //y2=2.96
cc_95 ( N_noxref_1_c_40_p N_noxref_7_c_938_n ) capacitor c=0.00209087f \
 //x=8.71 //y=0 //x2=10.245 //y2=2.96
cc_96 ( N_noxref_1_c_96_p N_noxref_7_c_938_n ) capacitor c=0.00129597f \
 //x=9.415 //y=0 //x2=10.245 //y2=2.96
cc_97 ( N_noxref_1_c_77_p N_noxref_7_c_938_n ) capacitor c=0.00114872f //x=9.9 \
 //y=0.535 //x2=10.245 //y2=2.96
cc_98 ( N_noxref_1_c_3_p N_noxref_7_c_938_n ) capacitor c=0.00750857f //x=5.55 \
 //y=0 //x2=10.245 //y2=2.96
cc_99 ( N_noxref_1_c_4_p N_noxref_7_c_938_n ) capacitor c=0.0144849f //x=8.88 \
 //y=0 //x2=10.245 //y2=2.96
cc_100 ( N_noxref_1_M5_noxref_s N_noxref_7_c_938_n ) capacitor c=0.00405051f \
 //x=9.375 //y=0.37 //x2=10.245 //y2=2.96
cc_101 ( N_noxref_1_c_2_p N_noxref_7_c_945_n ) capacitor c=6.9974e-19 //x=2.22 \
 //y=0 //x2=4.44 //y2=2.085
cc_102 ( N_noxref_1_c_3_p N_noxref_7_c_945_n ) capacitor c=0.00164431f \
 //x=5.55 //y=0 //x2=4.44 //y2=2.085
cc_103 ( N_noxref_1_c_6_p N_noxref_7_c_947_n ) capacitor c=0.00183756f \
 //x=10.36 //y=0 //x2=10.36 //y2=2.085
cc_104 ( N_noxref_1_c_104_p N_noxref_7_c_947_n ) capacitor c=7.8474e-19 \
 //x=10.385 //y=0.535 //x2=10.36 //y2=2.085
cc_105 ( N_noxref_1_c_4_p N_noxref_7_c_947_n ) capacitor c=0.00146529f \
 //x=8.88 //y=0 //x2=10.36 //y2=2.085
cc_106 ( N_noxref_1_c_5_p N_noxref_7_c_947_n ) capacitor c=0.0290276f \
 //x=10.47 //y=0 //x2=10.36 //y2=2.085
cc_107 ( N_noxref_1_M5_noxref_s N_noxref_7_c_947_n ) capacitor c=0.0102424f \
 //x=9.375 //y=0.37 //x2=10.36 //y2=2.085
cc_108 ( N_noxref_1_c_77_p N_noxref_7_c_952_n ) capacitor c=0.0119174f //x=9.9 \
 //y=0.535 //x2=9.72 //y2=0.91
cc_109 ( N_noxref_1_M5_noxref_s N_noxref_7_c_952_n ) capacitor c=0.0143355f \
 //x=9.375 //y=0.37 //x2=9.72 //y2=0.91
cc_110 ( N_noxref_1_M5_noxref_s N_noxref_7_c_954_n ) capacitor c=0.0074042f \
 //x=9.375 //y=0.37 //x2=9.72 //y2=1.255
cc_111 ( N_noxref_1_M5_noxref_s N_noxref_7_c_955_n ) capacitor c=0.00489f \
 //x=9.375 //y=0.37 //x2=10.095 //y2=0.755
cc_112 ( N_noxref_1_c_104_p N_noxref_7_c_956_n ) capacitor c=0.0123171f \
 //x=10.385 //y=0.535 //x2=10.25 //y2=0.91
cc_113 ( N_noxref_1_M5_noxref_s N_noxref_7_c_956_n ) capacitor c=0.0317181f \
 //x=9.375 //y=0.37 //x2=10.25 //y2=0.91
cc_114 ( N_noxref_1_c_5_p N_noxref_7_c_958_n ) capacitor c=0.0124051f \
 //x=10.47 //y=0 //x2=10.25 //y2=1.92
cc_115 ( N_noxref_1_c_104_p N_noxref_7_c_959_n ) capacitor c=2.1838e-19 \
 //x=10.385 //y=0.535 //x2=10.25 //y2=2.085
cc_116 ( N_noxref_1_c_5_p N_noxref_7_c_959_n ) capacitor c=0.0108179f \
 //x=10.47 //y=0 //x2=10.25 //y2=2.085
cc_117 ( N_noxref_1_M5_noxref_s N_noxref_7_c_959_n ) capacitor c=0.00652836f \
 //x=9.375 //y=0.37 //x2=10.25 //y2=2.085
cc_118 ( N_noxref_1_M0_noxref_s N_noxref_9_c_1151_n ) capacitor c=0.0013253f \
 //x=0.495 //y=0.37 //x2=2.915 //y2=1.5
cc_119 ( N_noxref_1_c_6_p N_noxref_9_c_1152_n ) capacitor c=0.00529166f \
 //x=10.36 //y=0 //x2=3.8 //y2=1.585
cc_120 ( N_noxref_1_c_23_p N_noxref_9_c_1152_n ) capacitor c=0.00112205f \
 //x=3.315 //y=0 //x2=3.8 //y2=1.585
cc_121 ( N_noxref_1_c_29_p N_noxref_9_c_1152_n ) capacitor c=0.00181496f \
 //x=5.38 //y=0 //x2=3.8 //y2=1.585
cc_122 ( N_noxref_1_M1_noxref_d N_noxref_9_c_1152_n ) capacitor c=0.00879196f \
 //x=3.21 //y=0.87 //x2=3.8 //y2=1.585
cc_123 ( N_noxref_1_c_6_p N_noxref_9_c_1156_n ) capacitor c=0.0026904f \
 //x=10.36 //y=0 //x2=3.885 //y2=0.62
cc_124 ( N_noxref_1_c_29_p N_noxref_9_c_1156_n ) capacitor c=0.0144735f \
 //x=5.38 //y=0 //x2=3.885 //y2=0.62
cc_125 ( N_noxref_1_c_5_p N_noxref_9_c_1156_n ) capacitor c=0.00141889f \
 //x=10.47 //y=0 //x2=3.885 //y2=0.62
cc_126 ( N_noxref_1_M1_noxref_d N_noxref_9_c_1156_n ) capacitor c=0.033812f \
 //x=3.21 //y=0.87 //x2=3.885 //y2=0.62
cc_127 ( N_noxref_1_c_2_p N_noxref_9_c_1160_n ) capacitor c=2.91423e-19 \
 //x=2.22 //y=0 //x2=3.885 //y2=1.5
cc_128 ( N_noxref_1_c_6_p N_noxref_9_c_1161_n ) capacitor c=0.0111125f \
 //x=10.36 //y=0 //x2=4.77 //y2=0.535
cc_129 ( N_noxref_1_c_29_p N_noxref_9_c_1161_n ) capacitor c=0.0370011f \
 //x=5.38 //y=0 //x2=4.77 //y2=0.535
cc_130 ( N_noxref_1_c_5_p N_noxref_9_c_1161_n ) capacitor c=0.00194827f \
 //x=10.47 //y=0 //x2=4.77 //y2=0.535
cc_131 ( N_noxref_1_c_6_p N_noxref_9_c_1164_n ) capacitor c=0.00268883f \
 //x=10.36 //y=0 //x2=4.855 //y2=0.62
cc_132 ( N_noxref_1_c_29_p N_noxref_9_c_1164_n ) capacitor c=0.0144105f \
 //x=5.38 //y=0 //x2=4.855 //y2=0.62
cc_133 ( N_noxref_1_c_3_p N_noxref_9_c_1164_n ) capacitor c=0.0431718f \
 //x=5.55 //y=0 //x2=4.855 //y2=0.62
cc_134 ( N_noxref_1_c_5_p N_noxref_9_c_1164_n ) capacitor c=0.00141054f \
 //x=10.47 //y=0 //x2=4.855 //y2=0.62
cc_135 ( N_noxref_1_c_6_p N_noxref_9_M1_noxref_s ) capacitor c=0.0026904f \
 //x=10.36 //y=0 //x2=2.78 //y2=0.37
cc_136 ( N_noxref_1_c_136_p N_noxref_9_M1_noxref_s ) capacitor c=0.0013253f \
 //x=1.6 //y=0.45 //x2=2.78 //y2=0.37
cc_137 ( N_noxref_1_c_23_p N_noxref_9_M1_noxref_s ) capacitor c=0.0144735f \
 //x=3.315 //y=0 //x2=2.78 //y2=0.37
cc_138 ( N_noxref_1_c_2_p N_noxref_9_M1_noxref_s ) capacitor c=0.058339f \
 //x=2.22 //y=0 //x2=2.78 //y2=0.37
cc_139 ( N_noxref_1_c_3_p N_noxref_9_M1_noxref_s ) capacitor c=0.00200438f \
 //x=5.55 //y=0 //x2=2.78 //y2=0.37
cc_140 ( N_noxref_1_c_5_p N_noxref_9_M1_noxref_s ) capacitor c=0.00141889f \
 //x=10.47 //y=0 //x2=2.78 //y2=0.37
cc_141 ( N_noxref_1_M1_noxref_d N_noxref_9_M1_noxref_s ) capacitor \
 c=0.0334197f //x=3.21 //y=0.87 //x2=2.78 //y2=0.37
cc_142 ( N_noxref_1_c_6_p N_noxref_11_c_1246_n ) capacitor c=0.00529166f \
 //x=10.36 //y=0 //x2=7.13 //y2=1.585
cc_143 ( N_noxref_1_c_39_p N_noxref_11_c_1246_n ) capacitor c=0.00112205f \
 //x=6.645 //y=0 //x2=7.13 //y2=1.585
cc_144 ( N_noxref_1_c_40_p N_noxref_11_c_1246_n ) capacitor c=0.00181496f \
 //x=8.71 //y=0 //x2=7.13 //y2=1.585
cc_145 ( N_noxref_1_M3_noxref_d N_noxref_11_c_1246_n ) capacitor c=0.00879196f \
 //x=6.54 //y=0.87 //x2=7.13 //y2=1.585
cc_146 ( N_noxref_1_c_6_p N_noxref_11_c_1250_n ) capacitor c=0.0026904f \
 //x=10.36 //y=0 //x2=7.215 //y2=0.62
cc_147 ( N_noxref_1_c_40_p N_noxref_11_c_1250_n ) capacitor c=0.0144735f \
 //x=8.71 //y=0 //x2=7.215 //y2=0.62
cc_148 ( N_noxref_1_c_5_p N_noxref_11_c_1250_n ) capacitor c=0.00141889f \
 //x=10.47 //y=0 //x2=7.215 //y2=0.62
cc_149 ( N_noxref_1_M3_noxref_d N_noxref_11_c_1250_n ) capacitor c=0.033812f \
 //x=6.54 //y=0.87 //x2=7.215 //y2=0.62
cc_150 ( N_noxref_1_c_3_p N_noxref_11_c_1254_n ) capacitor c=2.91423e-19 \
 //x=5.55 //y=0 //x2=7.215 //y2=1.5
cc_151 ( N_noxref_1_c_6_p N_noxref_11_c_1255_n ) capacitor c=0.0112038f \
 //x=10.36 //y=0 //x2=8.1 //y2=0.535
cc_152 ( N_noxref_1_c_40_p N_noxref_11_c_1255_n ) capacitor c=0.0370216f \
 //x=8.71 //y=0 //x2=8.1 //y2=0.535
cc_153 ( N_noxref_1_c_5_p N_noxref_11_c_1255_n ) capacitor c=0.00194827f \
 //x=10.47 //y=0 //x2=8.1 //y2=0.535
cc_154 ( N_noxref_1_c_6_p N_noxref_11_c_1258_n ) capacitor c=0.00280093f \
 //x=10.36 //y=0 //x2=8.185 //y2=0.62
cc_155 ( N_noxref_1_c_40_p N_noxref_11_c_1258_n ) capacitor c=0.0144899f \
 //x=8.71 //y=0 //x2=8.185 //y2=0.62
cc_156 ( N_noxref_1_c_156_p N_noxref_11_c_1258_n ) capacitor c=9.92084e-19 \
 //x=9.5 //y=0.45 //x2=8.185 //y2=0.62
cc_157 ( N_noxref_1_c_4_p N_noxref_11_c_1258_n ) capacitor c=0.0431718f \
 //x=8.88 //y=0 //x2=8.185 //y2=0.62
cc_158 ( N_noxref_1_c_5_p N_noxref_11_c_1258_n ) capacitor c=0.00141054f \
 //x=10.47 //y=0 //x2=8.185 //y2=0.62
cc_159 ( N_noxref_1_c_6_p N_noxref_11_M3_noxref_s ) capacitor c=0.0026904f \
 //x=10.36 //y=0 //x2=6.11 //y2=0.37
cc_160 ( N_noxref_1_c_39_p N_noxref_11_M3_noxref_s ) capacitor c=0.0144735f \
 //x=6.645 //y=0 //x2=6.11 //y2=0.37
cc_161 ( N_noxref_1_c_3_p N_noxref_11_M3_noxref_s ) capacitor c=0.058339f \
 //x=5.55 //y=0 //x2=6.11 //y2=0.37
cc_162 ( N_noxref_1_c_4_p N_noxref_11_M3_noxref_s ) capacitor c=0.00200548f \
 //x=8.88 //y=0 //x2=6.11 //y2=0.37
cc_163 ( N_noxref_1_c_5_p N_noxref_11_M3_noxref_s ) capacitor c=0.00141889f \
 //x=10.47 //y=0 //x2=6.11 //y2=0.37
cc_164 ( N_noxref_1_M3_noxref_d N_noxref_11_M3_noxref_s ) capacitor \
 c=0.0334197f //x=6.54 //y=0.87 //x2=6.11 //y2=0.37
cc_165 ( N_noxref_1_M5_noxref_s N_noxref_11_M3_noxref_s ) capacitor \
 c=9.92084e-19 //x=9.375 //y=0.37 //x2=6.11 //y2=0.37
cc_166 ( N_noxref_2_c_171_p N_noxref_3_c_322_n ) capacitor c=0.0179155f \
 //x=10.36 //y=7.4 //x2=3.215 //y2=4.07
cc_167 ( N_noxref_2_c_172_p N_noxref_3_c_322_n ) capacitor c=9.77842e-19 \
 //x=1.47 //y=7.4 //x2=3.215 //y2=4.07
cc_168 ( N_noxref_2_c_173_p N_noxref_3_c_322_n ) capacitor c=0.00124367f \
 //x=2.05 //y=7.4 //x2=3.215 //y2=4.07
cc_169 ( N_noxref_2_c_174_p N_noxref_3_c_322_n ) capacitor c=0.00216965f \
 //x=3.365 //y=7.4 //x2=3.215 //y2=4.07
cc_170 ( N_noxref_2_c_167_n N_noxref_3_c_322_n ) capacitor c=0.0280406f \
 //x=2.22 //y=7.4 //x2=3.215 //y2=4.07
cc_171 ( N_noxref_2_M7_noxref_d N_noxref_3_c_322_n ) capacitor c=0.00213856f \
 //x=1.41 //y=5.02 //x2=3.215 //y2=4.07
cc_172 ( N_noxref_2_c_171_p N_noxref_3_c_324_n ) capacitor c=0.00188164f \
 //x=10.36 //y=7.4 //x2=0.855 //y2=4.07
cc_173 ( N_noxref_2_c_166_n N_noxref_3_c_324_n ) capacitor c=0.00208272f \
 //x=0.74 //y=7.4 //x2=0.855 //y2=4.07
cc_174 ( N_noxref_2_M6_noxref_s N_noxref_3_c_324_n ) capacitor c=0.00185024f \
 //x=0.54 //y=5.02 //x2=0.855 //y2=4.07
cc_175 ( N_noxref_2_c_171_p N_noxref_3_c_326_n ) capacitor c=0.00157744f \
 //x=10.36 //y=7.4 //x2=0.74 //y2=2.085
cc_176 ( N_noxref_2_c_166_n N_noxref_3_c_326_n ) capacitor c=0.0272385f \
 //x=0.74 //y=7.4 //x2=0.74 //y2=2.085
cc_177 ( N_noxref_2_c_167_n N_noxref_3_c_326_n ) capacitor c=0.00139956f \
 //x=2.22 //y=7.4 //x2=0.74 //y2=2.085
cc_178 ( N_noxref_2_M6_noxref_s N_noxref_3_c_326_n ) capacitor c=0.00896093f \
 //x=0.54 //y=5.02 //x2=0.74 //y2=2.085
cc_179 ( N_noxref_2_c_167_n N_noxref_3_c_331_n ) capacitor c=0.0160048f \
 //x=2.22 //y=7.4 //x2=3.33 //y2=2.085
cc_180 ( N_noxref_2_c_172_p N_noxref_3_M6_noxref_g ) capacitor c=0.00748034f \
 //x=1.47 //y=7.4 //x2=0.895 //y2=6.02
cc_181 ( N_noxref_2_c_166_n N_noxref_3_M6_noxref_g ) capacitor c=0.0241676f \
 //x=0.74 //y=7.4 //x2=0.895 //y2=6.02
cc_182 ( N_noxref_2_M6_noxref_s N_noxref_3_M6_noxref_g ) capacitor \
 c=0.0528676f //x=0.54 //y=5.02 //x2=0.895 //y2=6.02
cc_183 ( N_noxref_2_c_172_p N_noxref_3_M7_noxref_g ) capacitor c=0.00697478f \
 //x=1.47 //y=7.4 //x2=1.335 //y2=6.02
cc_184 ( N_noxref_2_M7_noxref_d N_noxref_3_M7_noxref_g ) capacitor \
 c=0.0528676f //x=1.41 //y=5.02 //x2=1.335 //y2=6.02
cc_185 ( N_noxref_2_c_174_p N_noxref_3_M8_noxref_g ) capacitor c=0.00673447f \
 //x=3.365 //y=7.4 //x2=3.23 //y2=6.02
cc_186 ( N_noxref_2_c_167_n N_noxref_3_M8_noxref_g ) capacitor c=0.00449901f \
 //x=2.22 //y=7.4 //x2=3.23 //y2=6.02
cc_187 ( N_noxref_2_M8_noxref_d N_noxref_3_M8_noxref_g ) capacitor \
 c=0.0166176f //x=3.305 //y=5.02 //x2=3.23 //y2=6.02
cc_188 ( N_noxref_2_c_193_p N_noxref_3_M9_noxref_g ) capacitor c=0.006727f \
 //x=5.38 //y=7.4 //x2=3.67 //y2=6.02
cc_189 ( N_noxref_2_M8_noxref_d N_noxref_3_M9_noxref_g ) capacitor \
 c=0.0186652f //x=3.305 //y=5.02 //x2=3.67 //y2=6.02
cc_190 ( N_noxref_2_c_167_n N_noxref_3_c_375_n ) capacitor c=0.0132667f \
 //x=2.22 //y=7.4 //x2=1.26 //y2=4.79
cc_191 ( N_noxref_2_c_166_n N_noxref_3_c_376_n ) capacitor c=0.011132f \
 //x=0.74 //y=7.4 //x2=0.97 //y2=4.79
cc_192 ( N_noxref_2_M6_noxref_s N_noxref_3_c_376_n ) capacitor c=0.00524527f \
 //x=0.54 //y=5.02 //x2=0.97 //y2=4.79
cc_193 ( N_noxref_2_c_167_n N_noxref_3_c_378_n ) capacitor c=0.0125867f \
 //x=2.22 //y=7.4 //x2=3.33 //y2=4.7
cc_194 ( N_noxref_2_c_167_n N_noxref_4_c_455_n ) capacitor c=0.00137387f \
 //x=2.22 //y=7.4 //x2=7.655 //y2=2.59
cc_195 ( N_noxref_2_c_171_p N_noxref_4_c_482_n ) capacitor c=0.0012271f \
 //x=10.36 //y=7.4 //x2=1.395 //y2=4.58
cc_196 ( N_noxref_2_c_172_p N_noxref_4_c_482_n ) capacitor c=9.08147e-19 \
 //x=1.47 //y=7.4 //x2=1.395 //y2=4.58
cc_197 ( N_noxref_2_M7_noxref_d N_noxref_4_c_482_n ) capacitor c=0.00609088f \
 //x=1.41 //y=5.02 //x2=1.395 //y2=4.58
cc_198 ( N_noxref_2_c_166_n N_noxref_4_c_485_n ) capacitor c=0.0179238f \
 //x=0.74 //y=7.4 //x2=1.2 //y2=4.58
cc_199 ( N_noxref_2_c_166_n N_noxref_4_c_470_n ) capacitor c=5.65246e-19 \
 //x=0.74 //y=7.4 //x2=1.48 //y2=2.59
cc_200 ( N_noxref_2_c_167_n N_noxref_4_c_470_n ) capacitor c=0.0220651f \
 //x=2.22 //y=7.4 //x2=1.48 //y2=2.59
cc_201 ( N_noxref_2_c_168_n N_noxref_4_c_473_n ) capacitor c=0.00210246f \
 //x=5.55 //y=7.4 //x2=7.77 //y2=2.085
cc_202 ( N_noxref_2_c_169_n N_noxref_4_c_473_n ) capacitor c=0.00147528f \
 //x=8.88 //y=7.4 //x2=7.77 //y2=2.085
cc_203 ( N_noxref_2_c_208_p N_noxref_4_M14_noxref_g ) capacitor c=0.00510247f \
 //x=8.71 //y=7.4 //x2=7.44 //y2=6.02
cc_204 ( N_noxref_2_c_208_p N_noxref_4_M15_noxref_g ) capacitor c=0.00510919f \
 //x=8.71 //y=7.4 //x2=7.88 //y2=6.02
cc_205 ( N_noxref_2_c_169_n N_noxref_4_M15_noxref_g ) capacitor c=0.00788519f \
 //x=8.88 //y=7.4 //x2=7.88 //y2=6.02
cc_206 ( N_noxref_2_c_171_p N_noxref_4_M6_noxref_d ) capacitor c=0.00285171f \
 //x=10.36 //y=7.4 //x2=0.97 //y2=5.02
cc_207 ( N_noxref_2_c_172_p N_noxref_4_M6_noxref_d ) capacitor c=0.0141332f \
 //x=1.47 //y=7.4 //x2=0.97 //y2=5.02
cc_208 ( N_noxref_2_c_167_n N_noxref_4_M6_noxref_d ) capacitor c=0.0204646f \
 //x=2.22 //y=7.4 //x2=0.97 //y2=5.02
cc_209 ( N_noxref_2_c_170_n N_noxref_4_M6_noxref_d ) capacitor c=0.00135976f \
 //x=10.36 //y=7.4 //x2=0.97 //y2=5.02
cc_210 ( N_noxref_2_M6_noxref_s N_noxref_4_M6_noxref_d ) capacitor \
 c=0.0843065f //x=0.54 //y=5.02 //x2=0.97 //y2=5.02
cc_211 ( N_noxref_2_M7_noxref_d N_noxref_4_M6_noxref_d ) capacitor \
 c=0.0832641f //x=1.41 //y=5.02 //x2=0.97 //y2=5.02
cc_212 ( N_noxref_2_c_171_p N_noxref_5_c_636_n ) capacitor c=0.00114115f \
 //x=10.36 //y=7.4 //x2=4.725 //y2=5.205
cc_213 ( N_noxref_2_c_193_p N_noxref_5_c_636_n ) capacitor c=0.00139027f \
 //x=5.38 //y=7.4 //x2=4.725 //y2=5.205
cc_214 ( N_noxref_2_c_167_n N_noxref_5_c_638_n ) capacitor c=8.9933e-19 \
 //x=2.22 //y=7.4 //x2=4.415 //y2=5.205
cc_215 ( N_noxref_2_c_167_n N_noxref_5_c_625_n ) capacitor c=0.00163766f \
 //x=2.22 //y=7.4 //x2=4.81 //y2=3.7
cc_216 ( N_noxref_2_c_168_n N_noxref_5_c_625_n ) capacitor c=0.0445615f \
 //x=5.55 //y=7.4 //x2=4.81 //y2=3.7
cc_217 ( N_noxref_2_c_171_p N_noxref_5_c_641_n ) capacitor c=0.00113725f \
 //x=10.36 //y=7.4 //x2=8.055 //y2=5.205
cc_218 ( N_noxref_2_c_208_p N_noxref_5_c_641_n ) capacitor c=0.00138968f \
 //x=8.71 //y=7.4 //x2=8.055 //y2=5.205
cc_219 ( N_noxref_2_c_168_n N_noxref_5_c_643_n ) capacitor c=8.9933e-19 \
 //x=5.55 //y=7.4 //x2=7.745 //y2=5.205
cc_220 ( N_noxref_2_c_168_n N_noxref_5_c_628_n ) capacitor c=0.00177938f \
 //x=5.55 //y=7.4 //x2=8.14 //y2=3.7
cc_221 ( N_noxref_2_c_169_n N_noxref_5_c_628_n ) capacitor c=0.0420891f \
 //x=8.88 //y=7.4 //x2=8.14 //y2=3.7
cc_222 ( N_noxref_2_c_168_n N_noxref_5_M10_noxref_d ) capacitor c=0.00966019f \
 //x=5.55 //y=7.4 //x2=4.185 //y2=5.02
cc_223 ( N_noxref_2_M8_noxref_d N_noxref_5_M10_noxref_d ) capacitor \
 c=0.00561178f //x=3.305 //y=5.02 //x2=4.185 //y2=5.02
cc_224 ( N_noxref_2_c_169_n N_noxref_5_M14_noxref_d ) capacitor c=0.00966019f \
 //x=8.88 //y=7.4 //x2=7.515 //y2=5.02
cc_225 ( N_noxref_2_M12_noxref_d N_noxref_5_M14_noxref_d ) capacitor \
 c=0.00561178f //x=6.635 //y=5.02 //x2=7.515 //y2=5.02
cc_226 ( N_noxref_2_M16_noxref_s N_noxref_5_M14_noxref_d ) capacitor \
 c=5.00921e-19 //x=9.42 //y=5.02 //x2=7.515 //y2=5.02
cc_227 ( N_noxref_2_c_171_p N_noxref_6_c_794_n ) capacitor c=0.0245984f \
 //x=10.36 //y=7.4 //x2=9.505 //y2=4.07
cc_228 ( N_noxref_2_c_193_p N_noxref_6_c_794_n ) capacitor c=0.00187833f \
 //x=5.38 //y=7.4 //x2=9.505 //y2=4.07
cc_229 ( N_noxref_2_c_234_p N_noxref_6_c_794_n ) capacitor c=0.00213804f \
 //x=6.695 //y=7.4 //x2=9.505 //y2=4.07
cc_230 ( N_noxref_2_c_168_n N_noxref_6_c_794_n ) capacitor c=0.0272145f \
 //x=5.55 //y=7.4 //x2=9.505 //y2=4.07
cc_231 ( N_noxref_2_c_169_n N_noxref_6_c_794_n ) capacitor c=0.0150593f \
 //x=8.88 //y=7.4 //x2=9.505 //y2=4.07
cc_232 ( N_noxref_2_c_171_p N_noxref_6_c_799_n ) capacitor c=0.00164816f \
 //x=10.36 //y=7.4 //x2=4.555 //y2=4.07
cc_233 ( N_noxref_2_c_167_n N_noxref_6_c_800_n ) capacitor c=7.20931e-19 \
 //x=2.22 //y=7.4 //x2=4.44 //y2=4.07
cc_234 ( N_noxref_2_c_168_n N_noxref_6_c_800_n ) capacitor c=0.00211919f \
 //x=5.55 //y=7.4 //x2=4.44 //y2=4.07
cc_235 ( N_noxref_2_c_169_n N_noxref_6_c_774_n ) capacitor c=0.0195394f \
 //x=8.88 //y=7.4 //x2=9.62 //y2=3.33
cc_236 ( N_noxref_2_c_170_n N_noxref_6_c_774_n ) capacitor c=6.39704e-19 \
 //x=10.36 //y=7.4 //x2=9.62 //y2=3.33
cc_237 ( N_noxref_2_c_170_n N_noxref_6_c_804_n ) capacitor c=0.017898f \
 //x=10.36 //y=7.4 //x2=9.9 //y2=4.58
cc_238 ( N_noxref_2_c_171_p N_noxref_6_c_805_n ) capacitor c=0.00119381f \
 //x=10.36 //y=7.4 //x2=9.705 //y2=4.58
cc_239 ( N_noxref_2_c_244_p N_noxref_6_c_805_n ) capacitor c=0.0010061f \
 //x=10.34 //y=7.4 //x2=9.705 //y2=4.58
cc_240 ( N_noxref_2_M16_noxref_s N_noxref_6_c_805_n ) capacitor c=0.00562155f \
 //x=9.42 //y=5.02 //x2=9.705 //y2=4.58
cc_241 ( N_noxref_2_c_193_p N_noxref_6_M10_noxref_g ) capacitor c=0.00510247f \
 //x=5.38 //y=7.4 //x2=4.11 //y2=6.02
cc_242 ( N_noxref_2_c_193_p N_noxref_6_M11_noxref_g ) capacitor c=0.00510919f \
 //x=5.38 //y=7.4 //x2=4.55 //y2=6.02
cc_243 ( N_noxref_2_c_168_n N_noxref_6_M11_noxref_g ) capacitor c=0.0122307f \
 //x=5.55 //y=7.4 //x2=4.55 //y2=6.02
cc_244 ( N_noxref_2_c_171_p N_noxref_6_M16_noxref_d ) capacitor c=0.00275339f \
 //x=10.36 //y=7.4 //x2=9.84 //y2=5.02
cc_245 ( N_noxref_2_c_244_p N_noxref_6_M16_noxref_d ) capacitor c=0.0140667f \
 //x=10.34 //y=7.4 //x2=9.84 //y2=5.02
cc_246 ( N_noxref_2_c_169_n N_noxref_6_M16_noxref_d ) capacitor c=0.0201812f \
 //x=8.88 //y=7.4 //x2=9.84 //y2=5.02
cc_247 ( N_noxref_2_c_170_n N_noxref_6_M16_noxref_d ) capacitor c=0.00135976f \
 //x=10.36 //y=7.4 //x2=9.84 //y2=5.02
cc_248 ( N_noxref_2_M16_noxref_s N_noxref_6_M16_noxref_d ) capacitor \
 c=0.0832641f //x=9.42 //y=5.02 //x2=9.84 //y2=5.02
cc_249 ( N_noxref_2_M17_noxref_d N_noxref_6_M16_noxref_d ) capacitor \
 c=0.0843065f //x=10.28 //y=5.02 //x2=9.84 //y2=5.02
cc_250 ( N_noxref_2_c_171_p N_noxref_7_c_962_n ) capacitor c=0.0251462f \
 //x=10.36 //y=7.4 //x2=10.245 //y2=4.44
cc_251 ( N_noxref_2_c_208_p N_noxref_7_c_962_n ) capacitor c=0.00304371f \
 //x=8.71 //y=7.4 //x2=10.245 //y2=4.44
cc_252 ( N_noxref_2_c_257_p N_noxref_7_c_962_n ) capacitor c=0.00151604f \
 //x=9.46 //y=7.4 //x2=10.245 //y2=4.44
cc_253 ( N_noxref_2_c_244_p N_noxref_7_c_962_n ) capacitor c=0.00205064f \
 //x=10.34 //y=7.4 //x2=10.245 //y2=4.44
cc_254 ( N_noxref_2_c_169_n N_noxref_7_c_962_n ) capacitor c=0.0377357f \
 //x=8.88 //y=7.4 //x2=10.245 //y2=4.44
cc_255 ( N_noxref_2_c_170_n N_noxref_7_c_962_n ) capacitor c=0.00754285f \
 //x=10.36 //y=7.4 //x2=10.245 //y2=4.44
cc_256 ( N_noxref_2_M16_noxref_s N_noxref_7_c_962_n ) capacitor c=0.00317238f \
 //x=9.42 //y=5.02 //x2=10.245 //y2=4.44
cc_257 ( N_noxref_2_M17_noxref_d N_noxref_7_c_962_n ) capacitor c=0.00289303f \
 //x=10.28 //y=5.02 //x2=10.245 //y2=4.44
cc_258 ( N_noxref_2_c_171_p N_noxref_7_c_970_n ) capacitor c=0.00150124f \
 //x=10.36 //y=7.4 //x2=6.775 //y2=4.44
cc_259 ( N_noxref_2_c_168_n N_noxref_7_c_970_n ) capacitor c=0.00665137f \
 //x=5.55 //y=7.4 //x2=6.775 //y2=4.44
cc_260 ( N_noxref_2_c_168_n N_noxref_7_c_972_n ) capacitor c=0.0112651f \
 //x=5.55 //y=7.4 //x2=6.66 //y2=4.44
cc_261 ( N_noxref_2_c_171_p N_noxref_7_c_947_n ) capacitor c=0.00156416f \
 //x=10.36 //y=7.4 //x2=10.36 //y2=2.085
cc_262 ( N_noxref_2_c_169_n N_noxref_7_c_947_n ) capacitor c=9.21978e-19 \
 //x=8.88 //y=7.4 //x2=10.36 //y2=2.085
cc_263 ( N_noxref_2_c_170_n N_noxref_7_c_947_n ) capacitor c=0.0251635f \
 //x=10.36 //y=7.4 //x2=10.36 //y2=2.085
cc_264 ( N_noxref_2_M17_noxref_d N_noxref_7_c_947_n ) capacitor c=0.00892989f \
 //x=10.28 //y=5.02 //x2=10.36 //y2=2.085
cc_265 ( N_noxref_2_c_234_p N_noxref_7_M12_noxref_g ) capacitor c=0.00673447f \
 //x=6.695 //y=7.4 //x2=6.56 //y2=6.02
cc_266 ( N_noxref_2_c_168_n N_noxref_7_M12_noxref_g ) capacitor c=0.00661226f \
 //x=5.55 //y=7.4 //x2=6.56 //y2=6.02
cc_267 ( N_noxref_2_M12_noxref_d N_noxref_7_M12_noxref_g ) capacitor \
 c=0.0166176f //x=6.635 //y=5.02 //x2=6.56 //y2=6.02
cc_268 ( N_noxref_2_c_208_p N_noxref_7_M13_noxref_g ) capacitor c=0.006727f \
 //x=8.71 //y=7.4 //x2=7 //y2=6.02
cc_269 ( N_noxref_2_M12_noxref_d N_noxref_7_M13_noxref_g ) capacitor \
 c=0.0186652f //x=6.635 //y=5.02 //x2=7 //y2=6.02
cc_270 ( N_noxref_2_c_244_p N_noxref_7_M16_noxref_g ) capacitor c=0.00697478f \
 //x=10.34 //y=7.4 //x2=9.765 //y2=6.02
cc_271 ( N_noxref_2_M16_noxref_s N_noxref_7_M16_noxref_g ) capacitor \
 c=0.0528676f //x=9.42 //y=5.02 //x2=9.765 //y2=6.02
cc_272 ( N_noxref_2_c_244_p N_noxref_7_M17_noxref_g ) capacitor c=0.00748034f \
 //x=10.34 //y=7.4 //x2=10.205 //y2=6.02
cc_273 ( N_noxref_2_c_170_n N_noxref_7_M17_noxref_g ) capacitor c=0.0241676f \
 //x=10.36 //y=7.4 //x2=10.205 //y2=6.02
cc_274 ( N_noxref_2_M17_noxref_d N_noxref_7_M17_noxref_g ) capacitor \
 c=0.0528676f //x=10.28 //y=5.02 //x2=10.205 //y2=6.02
cc_275 ( N_noxref_2_c_169_n N_noxref_7_c_987_n ) capacitor c=0.0148045f \
 //x=8.88 //y=7.4 //x2=9.84 //y2=4.79
cc_276 ( N_noxref_2_c_170_n N_noxref_7_c_988_n ) capacitor c=0.0109438f \
 //x=10.36 //y=7.4 //x2=10.205 //y2=4.865
cc_277 ( N_noxref_2_M17_noxref_d N_noxref_7_c_988_n ) capacitor c=0.00523962f \
 //x=10.28 //y=5.02 //x2=10.205 //y2=4.865
cc_278 ( N_noxref_2_c_168_n N_noxref_7_c_990_n ) capacitor c=0.0124704f \
 //x=5.55 //y=7.4 //x2=6.66 //y2=4.7
cc_279 ( N_noxref_2_c_171_p N_noxref_8_c_1111_n ) capacitor c=0.00494742f \
 //x=10.36 //y=7.4 //x2=3.805 //y2=5.205
cc_280 ( N_noxref_2_c_174_p N_noxref_8_c_1111_n ) capacitor c=4.50595e-19 \
 //x=3.365 //y=7.4 //x2=3.805 //y2=5.205
cc_281 ( N_noxref_2_c_193_p N_noxref_8_c_1111_n ) capacitor c=4.35755e-19 \
 //x=5.38 //y=7.4 //x2=3.805 //y2=5.205
cc_282 ( N_noxref_2_c_168_n N_noxref_8_c_1111_n ) capacitor c=0.00289291f \
 //x=5.55 //y=7.4 //x2=3.805 //y2=5.205
cc_283 ( N_noxref_2_M8_noxref_d N_noxref_8_c_1111_n ) capacitor c=0.0127094f \
 //x=3.305 //y=5.02 //x2=3.805 //y2=5.205
cc_284 ( N_noxref_2_c_167_n N_noxref_8_c_1116_n ) capacitor c=0.0628444f \
 //x=2.22 //y=7.4 //x2=3.095 //y2=5.205
cc_285 ( N_noxref_2_M7_noxref_d N_noxref_8_c_1116_n ) capacitor c=0.00269577f \
 //x=1.41 //y=5.02 //x2=3.095 //y2=5.205
cc_286 ( N_noxref_2_c_170_n N_noxref_8_c_1118_n ) capacitor c=0.00351514f \
 //x=10.36 //y=7.4 //x2=4.685 //y2=6.905
cc_287 ( N_noxref_2_c_171_p N_noxref_8_c_1119_n ) capacitor c=0.0260915f \
 //x=10.36 //y=7.4 //x2=3.975 //y2=6.905
cc_288 ( N_noxref_2_c_193_p N_noxref_8_c_1119_n ) capacitor c=0.0593394f \
 //x=5.38 //y=7.4 //x2=3.975 //y2=6.905
cc_289 ( N_noxref_2_c_170_n N_noxref_8_c_1119_n ) capacitor c=0.00115705f \
 //x=10.36 //y=7.4 //x2=3.975 //y2=6.905
cc_290 ( N_noxref_2_c_171_p N_noxref_8_M8_noxref_s ) capacitor c=0.00242367f \
 //x=10.36 //y=7.4 //x2=2.875 //y2=5.02
cc_291 ( N_noxref_2_c_174_p N_noxref_8_M8_noxref_s ) capacitor c=0.0100244f \
 //x=3.365 //y=7.4 //x2=2.875 //y2=5.02
cc_292 ( N_noxref_2_c_170_n N_noxref_8_M8_noxref_s ) capacitor c=7.63704e-19 \
 //x=10.36 //y=7.4 //x2=2.875 //y2=5.02
cc_293 ( N_noxref_2_M8_noxref_d N_noxref_8_M8_noxref_s ) capacitor c=0.061257f \
 //x=3.305 //y=5.02 //x2=2.875 //y2=5.02
cc_294 ( N_noxref_2_c_167_n N_noxref_8_M9_noxref_d ) capacitor c=0.00130916f \
 //x=2.22 //y=7.4 //x2=3.745 //y2=5.02
cc_295 ( N_noxref_2_M8_noxref_d N_noxref_8_M9_noxref_d ) capacitor \
 c=0.0659925f //x=3.305 //y=5.02 //x2=3.745 //y2=5.02
cc_296 ( N_noxref_2_c_168_n N_noxref_8_M11_noxref_d ) capacitor c=0.0520312f \
 //x=5.55 //y=7.4 //x2=4.625 //y2=5.02
cc_297 ( N_noxref_2_M8_noxref_d N_noxref_8_M11_noxref_d ) capacitor \
 c=0.00107819f //x=3.305 //y=5.02 //x2=4.625 //y2=5.02
cc_298 ( N_noxref_2_c_171_p N_noxref_10_c_1203_n ) capacitor c=0.00445614f \
 //x=10.36 //y=7.4 //x2=7.135 //y2=5.205
cc_299 ( N_noxref_2_c_234_p N_noxref_10_c_1203_n ) capacitor c=4.50436e-19 \
 //x=6.695 //y=7.4 //x2=7.135 //y2=5.205
cc_300 ( N_noxref_2_c_208_p N_noxref_10_c_1203_n ) capacitor c=4.50291e-19 \
 //x=8.71 //y=7.4 //x2=7.135 //y2=5.205
cc_301 ( N_noxref_2_c_169_n N_noxref_10_c_1203_n ) capacitor c=0.00289291f \
 //x=8.88 //y=7.4 //x2=7.135 //y2=5.205
cc_302 ( N_noxref_2_M12_noxref_d N_noxref_10_c_1203_n ) capacitor c=0.0123249f \
 //x=6.635 //y=5.02 //x2=7.135 //y2=5.205
cc_303 ( N_noxref_2_c_168_n N_noxref_10_c_1208_n ) capacitor c=0.0628444f \
 //x=5.55 //y=7.4 //x2=6.425 //y2=5.205
cc_304 ( N_noxref_2_c_170_n N_noxref_10_c_1209_n ) capacitor c=0.00351514f \
 //x=10.36 //y=7.4 //x2=8.015 //y2=6.905
cc_305 ( N_noxref_2_c_171_p N_noxref_10_c_1210_n ) capacitor c=0.0164961f \
 //x=10.36 //y=7.4 //x2=7.305 //y2=6.905
cc_306 ( N_noxref_2_c_208_p N_noxref_10_c_1210_n ) capacitor c=0.0608014f \
 //x=8.71 //y=7.4 //x2=7.305 //y2=6.905
cc_307 ( N_noxref_2_c_170_n N_noxref_10_c_1210_n ) capacitor c=0.00115705f \
 //x=10.36 //y=7.4 //x2=7.305 //y2=6.905
cc_308 ( N_noxref_2_c_171_p N_noxref_10_M12_noxref_s ) capacitor c=0.00242367f \
 //x=10.36 //y=7.4 //x2=6.205 //y2=5.02
cc_309 ( N_noxref_2_c_234_p N_noxref_10_M12_noxref_s ) capacitor c=0.0100244f \
 //x=6.695 //y=7.4 //x2=6.205 //y2=5.02
cc_310 ( N_noxref_2_c_170_n N_noxref_10_M12_noxref_s ) capacitor c=7.63704e-19 \
 //x=10.36 //y=7.4 //x2=6.205 //y2=5.02
cc_311 ( N_noxref_2_M12_noxref_d N_noxref_10_M12_noxref_s ) capacitor \
 c=0.061257f //x=6.635 //y=5.02 //x2=6.205 //y2=5.02
cc_312 ( N_noxref_2_c_168_n N_noxref_10_M13_noxref_d ) capacitor c=0.00130916f \
 //x=5.55 //y=7.4 //x2=7.075 //y2=5.02
cc_313 ( N_noxref_2_M12_noxref_d N_noxref_10_M13_noxref_d ) capacitor \
 c=0.0659925f //x=6.635 //y=5.02 //x2=7.075 //y2=5.02
cc_314 ( N_noxref_2_c_169_n N_noxref_10_M15_noxref_d ) capacitor c=0.0520312f \
 //x=8.88 //y=7.4 //x2=7.955 //y2=5.02
cc_315 ( N_noxref_2_M12_noxref_d N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00107819f //x=6.635 //y=5.02 //x2=7.955 //y2=5.02
cc_316 ( N_noxref_2_M16_noxref_s N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00230193f //x=9.42 //y=5.02 //x2=7.955 //y2=5.02
cc_317 ( N_noxref_3_c_322_n N_noxref_4_c_455_n ) capacitor c=0.0423762f \
 //x=3.215 //y=4.07 //x2=7.655 //y2=2.59
cc_318 ( N_noxref_3_c_331_n N_noxref_4_c_455_n ) capacitor c=0.0272208f \
 //x=3.33 //y=2.085 //x2=7.655 //y2=2.59
cc_319 ( N_noxref_3_c_342_n N_noxref_4_c_455_n ) capacitor c=0.00398285f \
 //x=3.135 //y=1.92 //x2=7.655 //y2=2.59
cc_320 ( N_noxref_3_c_322_n N_noxref_4_c_464_n ) capacitor c=0.00521938f \
 //x=3.215 //y=4.07 //x2=1.595 //y2=2.59
cc_321 ( N_noxref_3_c_326_n N_noxref_4_c_464_n ) capacitor c=0.00735597f \
 //x=0.74 //y=2.085 //x2=1.595 //y2=2.59
cc_322 ( N_noxref_3_c_331_n N_noxref_4_c_467_n ) capacitor c=0.0160774f \
 //x=3.33 //y=2.085 //x2=1.395 //y2=2.08
cc_323 ( N_noxref_3_c_385_p N_noxref_4_c_467_n ) capacitor c=0.0023507f \
 //x=1.225 //y=1.41 //x2=1.395 //y2=2.08
cc_324 ( N_noxref_3_c_322_n N_noxref_4_c_506_n ) capacitor c=0.0023373f \
 //x=3.215 //y=4.07 //x2=1.195 //y2=2.08
cc_325 ( N_noxref_3_c_348_n N_noxref_4_c_506_n ) capacitor c=0.0167852f \
 //x=0.74 //y=2.085 //x2=1.195 //y2=2.08
cc_326 ( N_noxref_3_c_375_n N_noxref_4_c_482_n ) capacitor c=0.0099173f \
 //x=1.26 //y=4.79 //x2=1.395 //y2=4.58
cc_327 ( N_noxref_3_c_322_n N_noxref_4_c_485_n ) capacitor c=0.0123666f \
 //x=3.215 //y=4.07 //x2=1.2 //y2=4.58
cc_328 ( N_noxref_3_c_326_n N_noxref_4_c_485_n ) capacitor c=0.0250789f \
 //x=0.74 //y=2.085 //x2=1.2 //y2=4.58
cc_329 ( N_noxref_3_c_376_n N_noxref_4_c_485_n ) capacitor c=0.00962086f \
 //x=0.97 //y=4.79 //x2=1.2 //y2=4.58
cc_330 ( N_noxref_3_c_322_n N_noxref_4_c_470_n ) capacitor c=0.0269755f \
 //x=3.215 //y=4.07 //x2=1.48 //y2=2.59
cc_331 ( N_noxref_3_c_324_n N_noxref_4_c_470_n ) capacitor c=0.00101501f \
 //x=0.855 //y=4.07 //x2=1.48 //y2=2.59
cc_332 ( N_noxref_3_c_326_n N_noxref_4_c_470_n ) capacitor c=0.068675f \
 //x=0.74 //y=2.085 //x2=1.48 //y2=2.59
cc_333 ( N_noxref_3_c_348_n N_noxref_4_c_470_n ) capacitor c=8.49451e-19 \
 //x=0.74 //y=2.085 //x2=1.48 //y2=2.59
cc_334 ( N_noxref_3_c_326_n N_noxref_4_M0_noxref_d ) capacitor c=0.0175773f \
 //x=0.74 //y=2.085 //x2=0.925 //y2=0.91
cc_335 ( N_noxref_3_c_332_n N_noxref_4_M0_noxref_d ) capacitor c=0.00218556f \
 //x=0.85 //y=0.91 //x2=0.925 //y2=0.91
cc_336 ( N_noxref_3_c_398_p N_noxref_4_M0_noxref_d ) capacitor c=0.00347355f \
 //x=0.85 //y=1.255 //x2=0.925 //y2=0.91
cc_337 ( N_noxref_3_c_399_p N_noxref_4_M0_noxref_d ) capacitor c=0.00742431f \
 //x=0.85 //y=1.565 //x2=0.925 //y2=0.91
cc_338 ( N_noxref_3_c_334_n N_noxref_4_M0_noxref_d ) capacitor c=0.00957707f \
 //x=0.85 //y=1.92 //x2=0.925 //y2=0.91
cc_339 ( N_noxref_3_c_335_n N_noxref_4_M0_noxref_d ) capacitor c=0.00220879f \
 //x=1.225 //y=0.755 //x2=0.925 //y2=0.91
cc_340 ( N_noxref_3_c_385_p N_noxref_4_M0_noxref_d ) capacitor c=0.0138447f \
 //x=1.225 //y=1.41 //x2=0.925 //y2=0.91
cc_341 ( N_noxref_3_c_336_n N_noxref_4_M0_noxref_d ) capacitor c=0.00218624f \
 //x=1.38 //y=0.91 //x2=0.925 //y2=0.91
cc_342 ( N_noxref_3_c_338_n N_noxref_4_M0_noxref_d ) capacitor c=0.00601286f \
 //x=1.38 //y=1.255 //x2=0.925 //y2=0.91
cc_343 ( N_noxref_3_M6_noxref_g N_noxref_4_M6_noxref_d ) capacitor \
 c=0.0219309f //x=0.895 //y=6.02 //x2=0.97 //y2=5.02
cc_344 ( N_noxref_3_M7_noxref_g N_noxref_4_M6_noxref_d ) capacitor c=0.021902f \
 //x=1.335 //y=6.02 //x2=0.97 //y2=5.02
cc_345 ( N_noxref_3_c_375_n N_noxref_4_M6_noxref_d ) capacitor c=0.0146106f \
 //x=1.26 //y=4.79 //x2=0.97 //y2=5.02
cc_346 ( N_noxref_3_c_376_n N_noxref_4_M6_noxref_d ) capacitor c=0.00307344f \
 //x=0.97 //y=4.79 //x2=0.97 //y2=5.02
cc_347 ( N_noxref_3_c_331_n N_noxref_5_c_651_n ) capacitor c=0.00382062f \
 //x=3.33 //y=2.085 //x2=4.925 //y2=3.7
cc_348 ( N_noxref_3_c_331_n N_noxref_5_c_625_n ) capacitor c=0.0153974f \
 //x=3.33 //y=2.085 //x2=4.81 //y2=3.7
cc_349 ( N_noxref_3_c_322_n N_noxref_6_c_799_n ) capacitor c=0.0159617f \
 //x=3.215 //y=4.07 //x2=4.555 //y2=4.07
cc_350 ( N_noxref_3_c_331_n N_noxref_6_c_799_n ) capacitor c=0.00187343f \
 //x=3.33 //y=2.085 //x2=4.555 //y2=4.07
cc_351 ( N_noxref_3_c_322_n N_noxref_6_c_800_n ) capacitor c=0.00186775f \
 //x=3.215 //y=4.07 //x2=4.44 //y2=4.07
cc_352 ( N_noxref_3_c_331_n N_noxref_6_c_800_n ) capacitor c=0.0166316f \
 //x=3.33 //y=2.085 //x2=4.44 //y2=4.07
cc_353 ( N_noxref_3_c_378_n N_noxref_6_c_800_n ) capacitor c=0.0022916f \
 //x=3.33 //y=4.7 //x2=4.44 //y2=4.07
cc_354 ( N_noxref_3_c_331_n N_noxref_6_c_773_n ) capacitor c=2.12957e-19 \
 //x=3.33 //y=2.085 //x2=6.66 //y2=2.085
cc_355 ( N_noxref_3_M8_noxref_g N_noxref_6_M10_noxref_g ) capacitor \
 c=0.0100243f //x=3.23 //y=6.02 //x2=4.11 //y2=6.02
cc_356 ( N_noxref_3_M9_noxref_g N_noxref_6_M10_noxref_g ) capacitor \
 c=0.0610135f //x=3.67 //y=6.02 //x2=4.11 //y2=6.02
cc_357 ( N_noxref_3_M9_noxref_g N_noxref_6_M11_noxref_g ) capacitor \
 c=0.0094155f //x=3.67 //y=6.02 //x2=4.55 //y2=6.02
cc_358 ( N_noxref_3_c_331_n N_noxref_6_c_826_n ) capacitor c=0.00227843f \
 //x=3.33 //y=2.085 //x2=4.44 //y2=4.7
cc_359 ( N_noxref_3_c_378_n N_noxref_6_c_826_n ) capacitor c=0.066749f \
 //x=3.33 //y=4.7 //x2=4.44 //y2=4.7
cc_360 ( N_noxref_3_c_331_n N_noxref_7_c_991_n ) capacitor c=0.00526349f \
 //x=3.33 //y=2.085 //x2=4.555 //y2=2.96
cc_361 ( N_noxref_3_c_331_n N_noxref_7_c_945_n ) capacitor c=0.019701f \
 //x=3.33 //y=2.085 //x2=4.44 //y2=2.085
cc_362 ( N_noxref_3_c_342_n N_noxref_7_c_945_n ) capacitor c=0.00220284f \
 //x=3.135 //y=1.92 //x2=4.44 //y2=2.085
cc_363 ( N_noxref_3_c_339_n N_noxref_7_c_994_n ) capacitor c=4.86506e-19 \
 //x=3.135 //y=0.87 //x2=4.105 //y2=0.91
cc_364 ( N_noxref_3_c_341_n N_noxref_7_c_994_n ) capacitor c=0.00152104f \
 //x=3.135 //y=1.215 //x2=4.105 //y2=0.91
cc_365 ( N_noxref_3_c_345_n N_noxref_7_c_994_n ) capacitor c=0.0157772f \
 //x=3.665 //y=0.87 //x2=4.105 //y2=0.91
cc_366 ( N_noxref_3_c_428_p N_noxref_7_c_997_n ) capacitor c=0.00109982f \
 //x=3.135 //y=1.525 //x2=4.105 //y2=1.255
cc_367 ( N_noxref_3_c_347_n N_noxref_7_c_997_n ) capacitor c=0.0117362f \
 //x=3.665 //y=1.215 //x2=4.105 //y2=1.255
cc_368 ( N_noxref_3_c_428_p N_noxref_7_c_999_n ) capacitor c=9.57794e-19 \
 //x=3.135 //y=1.525 //x2=4.105 //y2=1.565
cc_369 ( N_noxref_3_c_342_n N_noxref_7_c_999_n ) capacitor c=0.00662747f \
 //x=3.135 //y=1.92 //x2=4.105 //y2=1.565
cc_370 ( N_noxref_3_c_347_n N_noxref_7_c_999_n ) capacitor c=0.00862358f \
 //x=3.665 //y=1.215 //x2=4.105 //y2=1.565
cc_371 ( N_noxref_3_c_331_n N_noxref_7_c_1002_n ) capacitor c=0.00251238f \
 //x=3.33 //y=2.085 //x2=4.105 //y2=1.92
cc_372 ( N_noxref_3_c_342_n N_noxref_7_c_1002_n ) capacitor c=0.012079f \
 //x=3.135 //y=1.92 //x2=4.105 //y2=1.92
cc_373 ( N_noxref_3_c_345_n N_noxref_7_c_1004_n ) capacitor c=0.00124821f \
 //x=3.665 //y=0.87 //x2=4.635 //y2=0.91
cc_374 ( N_noxref_3_c_347_n N_noxref_7_c_1005_n ) capacitor c=0.00200715f \
 //x=3.665 //y=1.215 //x2=4.635 //y2=1.255
cc_375 ( N_noxref_3_c_322_n N_noxref_8_c_1111_n ) capacitor c=0.00305144f \
 //x=3.215 //y=4.07 //x2=3.805 //y2=5.205
cc_376 ( N_noxref_3_c_331_n N_noxref_8_c_1111_n ) capacitor c=0.0120071f \
 //x=3.33 //y=2.085 //x2=3.805 //y2=5.205
cc_377 ( N_noxref_3_M8_noxref_g N_noxref_8_c_1111_n ) capacitor c=0.019052f \
 //x=3.23 //y=6.02 //x2=3.805 //y2=5.205
cc_378 ( N_noxref_3_M9_noxref_g N_noxref_8_c_1111_n ) capacitor c=0.0198429f \
 //x=3.67 //y=6.02 //x2=3.805 //y2=5.205
cc_379 ( N_noxref_3_c_378_n N_noxref_8_c_1111_n ) capacitor c=0.00525548f \
 //x=3.33 //y=4.7 //x2=3.805 //y2=5.205
cc_380 ( N_noxref_3_c_322_n N_noxref_8_c_1116_n ) capacitor c=0.00704018f \
 //x=3.215 //y=4.07 //x2=3.095 //y2=5.205
cc_381 ( N_noxref_3_M8_noxref_g N_noxref_8_M8_noxref_s ) capacitor \
 c=0.0441361f //x=3.23 //y=6.02 //x2=2.875 //y2=5.02
cc_382 ( N_noxref_3_M9_noxref_g N_noxref_8_M9_noxref_d ) capacitor \
 c=0.0170604f //x=3.67 //y=6.02 //x2=3.745 //y2=5.02
cc_383 ( N_noxref_3_c_342_n N_noxref_9_c_1151_n ) capacitor c=0.0034165f \
 //x=3.135 //y=1.92 //x2=2.915 //y2=1.5
cc_384 ( N_noxref_3_c_331_n N_noxref_9_c_1152_n ) capacitor c=0.0114213f \
 //x=3.33 //y=2.085 //x2=3.8 //y2=1.585
cc_385 ( N_noxref_3_c_428_p N_noxref_9_c_1152_n ) capacitor c=0.00704065f \
 //x=3.135 //y=1.525 //x2=3.8 //y2=1.585
cc_386 ( N_noxref_3_c_342_n N_noxref_9_c_1152_n ) capacitor c=0.0185489f \
 //x=3.135 //y=1.92 //x2=3.8 //y2=1.585
cc_387 ( N_noxref_3_c_344_n N_noxref_9_c_1152_n ) capacitor c=0.00780802f \
 //x=3.51 //y=1.37 //x2=3.8 //y2=1.585
cc_388 ( N_noxref_3_c_347_n N_noxref_9_c_1152_n ) capacitor c=0.0034036f \
 //x=3.665 //y=1.215 //x2=3.8 //y2=1.585
cc_389 ( N_noxref_3_c_342_n N_noxref_9_c_1160_n ) capacitor c=6.71402e-19 \
 //x=3.135 //y=1.92 //x2=3.885 //y2=1.5
cc_390 ( N_noxref_3_c_339_n N_noxref_9_M1_noxref_s ) capacitor c=0.0326577f \
 //x=3.135 //y=0.87 //x2=2.78 //y2=0.37
cc_391 ( N_noxref_3_c_428_p N_noxref_9_M1_noxref_s ) capacitor c=3.48408e-19 \
 //x=3.135 //y=1.525 //x2=2.78 //y2=0.37
cc_392 ( N_noxref_3_c_345_n N_noxref_9_M1_noxref_s ) capacitor c=0.0120759f \
 //x=3.665 //y=0.87 //x2=2.78 //y2=0.37
cc_393 ( N_noxref_4_c_455_n N_noxref_5_c_653_n ) capacitor c=0.00619185f \
 //x=7.655 //y=2.59 //x2=8.025 //y2=3.7
cc_394 ( N_noxref_4_c_473_n N_noxref_5_c_653_n ) capacitor c=0.0182357f \
 //x=7.77 //y=2.085 //x2=8.025 //y2=3.7
cc_395 ( N_noxref_4_c_455_n N_noxref_5_c_651_n ) capacitor c=6.30506e-19 \
 //x=7.655 //y=2.59 //x2=4.925 //y2=3.7
cc_396 ( N_noxref_4_c_473_n N_noxref_5_c_651_n ) capacitor c=2.02744e-19 \
 //x=7.77 //y=2.085 //x2=4.925 //y2=3.7
cc_397 ( N_noxref_4_c_455_n N_noxref_5_c_638_n ) capacitor c=4.14299e-19 \
 //x=7.655 //y=2.59 //x2=4.415 //y2=5.205
cc_398 ( N_noxref_4_c_455_n N_noxref_5_c_624_n ) capacitor c=0.00452983f \
 //x=7.655 //y=2.59 //x2=4.725 //y2=1.655
cc_399 ( N_noxref_4_c_455_n N_noxref_5_c_659_n ) capacitor c=0.00179594f \
 //x=7.655 //y=2.59 //x2=4.455 //y2=1.655
cc_400 ( N_noxref_4_c_455_n N_noxref_5_c_625_n ) capacitor c=0.0188614f \
 //x=7.655 //y=2.59 //x2=4.81 //y2=3.7
cc_401 ( N_noxref_4_c_470_n N_noxref_5_c_625_n ) capacitor c=2.79968e-19 \
 //x=1.48 //y=2.59 //x2=4.81 //y2=3.7
cc_402 ( N_noxref_4_c_473_n N_noxref_5_c_625_n ) capacitor c=0.00277451f \
 //x=7.77 //y=2.085 //x2=4.81 //y2=3.7
cc_403 ( N_noxref_4_M15_noxref_g N_noxref_5_c_641_n ) capacitor c=0.0180846f \
 //x=7.88 //y=6.02 //x2=8.055 //y2=5.205
cc_404 ( N_noxref_4_c_540_p N_noxref_5_c_641_n ) capacitor c=0.00161455f \
 //x=7.77 //y=4.7 //x2=8.055 //y2=5.205
cc_405 ( N_noxref_4_c_473_n N_noxref_5_c_643_n ) capacitor c=0.0129715f \
 //x=7.77 //y=2.085 //x2=7.745 //y2=5.205
cc_406 ( N_noxref_4_M14_noxref_g N_noxref_5_c_643_n ) capacitor c=0.0132788f \
 //x=7.44 //y=6.02 //x2=7.745 //y2=5.205
cc_407 ( N_noxref_4_c_540_p N_noxref_5_c_643_n ) capacitor c=0.00554627f \
 //x=7.77 //y=4.7 //x2=7.745 //y2=5.205
cc_408 ( N_noxref_4_c_455_n N_noxref_5_c_626_n ) capacitor c=0.00140545f \
 //x=7.655 //y=2.59 //x2=8.055 //y2=1.655
cc_409 ( N_noxref_4_c_545_p N_noxref_5_c_626_n ) capacitor c=0.00363601f \
 //x=7.435 //y=1.92 //x2=8.055 //y2=1.655
cc_410 ( N_noxref_4_c_546_p N_noxref_5_c_626_n ) capacitor c=0.00196666f \
 //x=7.81 //y=1.41 //x2=8.055 //y2=1.655
cc_411 ( N_noxref_4_c_547_p N_noxref_5_c_626_n ) capacitor c=0.00423452f \
 //x=7.965 //y=1.255 //x2=8.055 //y2=1.655
cc_412 ( N_noxref_4_c_455_n N_noxref_5_c_672_n ) capacitor c=0.00185456f \
 //x=7.655 //y=2.59 //x2=7.785 //y2=1.655
cc_413 ( N_noxref_4_c_473_n N_noxref_5_c_672_n ) capacitor c=0.0170992f \
 //x=7.77 //y=2.085 //x2=7.785 //y2=1.655
cc_414 ( N_noxref_4_c_545_p N_noxref_5_c_672_n ) capacitor c=0.00637984f \
 //x=7.435 //y=1.92 //x2=7.785 //y2=1.655
cc_415 ( N_noxref_4_c_455_n N_noxref_5_c_628_n ) capacitor c=0.0100753f \
 //x=7.655 //y=2.59 //x2=8.14 //y2=3.7
cc_416 ( N_noxref_4_c_473_n N_noxref_5_c_628_n ) capacitor c=0.187239f \
 //x=7.77 //y=2.085 //x2=8.14 //y2=3.7
cc_417 ( N_noxref_4_c_545_p N_noxref_5_c_628_n ) capacitor c=0.0185661f \
 //x=7.435 //y=1.92 //x2=8.14 //y2=3.7
cc_418 ( N_noxref_4_c_540_p N_noxref_5_c_628_n ) capacitor c=0.0232466f \
 //x=7.77 //y=4.7 //x2=8.14 //y2=3.7
cc_419 ( N_noxref_4_c_555_p N_noxref_5_M4_noxref_d ) capacitor c=0.00217566f \
 //x=7.435 //y=0.91 //x2=7.51 //y2=0.91
cc_420 ( N_noxref_4_c_556_p N_noxref_5_M4_noxref_d ) capacitor c=0.0034598f \
 //x=7.435 //y=1.255 //x2=7.51 //y2=0.91
cc_421 ( N_noxref_4_c_557_p N_noxref_5_M4_noxref_d ) capacitor c=0.00522042f \
 //x=7.435 //y=1.565 //x2=7.51 //y2=0.91
cc_422 ( N_noxref_4_c_545_p N_noxref_5_M4_noxref_d ) capacitor c=0.00643086f \
 //x=7.435 //y=1.92 //x2=7.51 //y2=0.91
cc_423 ( N_noxref_4_c_559_p N_noxref_5_M4_noxref_d ) capacitor c=0.00241053f \
 //x=7.81 //y=0.755 //x2=7.51 //y2=0.91
cc_424 ( N_noxref_4_c_546_p N_noxref_5_M4_noxref_d ) capacitor c=0.0124466f \
 //x=7.81 //y=1.41 //x2=7.51 //y2=0.91
cc_425 ( N_noxref_4_c_561_p N_noxref_5_M4_noxref_d ) capacitor c=0.00132245f \
 //x=7.965 //y=0.91 //x2=7.51 //y2=0.91
cc_426 ( N_noxref_4_c_547_p N_noxref_5_M4_noxref_d ) capacitor c=0.00566463f \
 //x=7.965 //y=1.255 //x2=7.51 //y2=0.91
cc_427 ( N_noxref_4_M15_noxref_g N_noxref_5_M14_noxref_d ) capacitor \
 c=0.0136385f //x=7.88 //y=6.02 //x2=7.515 //y2=5.02
cc_428 ( N_noxref_4_c_455_n N_noxref_6_c_794_n ) capacitor c=7.67045e-19 \
 //x=7.655 //y=2.59 //x2=9.505 //y2=4.07
cc_429 ( N_noxref_4_c_473_n N_noxref_6_c_794_n ) capacitor c=0.0166527f \
 //x=7.77 //y=2.085 //x2=9.505 //y2=4.07
cc_430 ( N_noxref_4_c_455_n N_noxref_6_c_799_n ) capacitor c=6.56372e-19 \
 //x=7.655 //y=2.59 //x2=4.555 //y2=4.07
cc_431 ( N_noxref_4_c_455_n N_noxref_6_c_831_n ) capacitor c=0.00949286f \
 //x=7.655 //y=2.59 //x2=9.505 //y2=3.33
cc_432 ( N_noxref_4_c_473_n N_noxref_6_c_831_n ) capacitor c=0.0158195f \
 //x=7.77 //y=2.085 //x2=9.505 //y2=3.33
cc_433 ( N_noxref_4_c_455_n N_noxref_6_c_833_n ) capacitor c=9.78991e-19 \
 //x=7.655 //y=2.59 //x2=6.775 //y2=3.33
cc_434 ( N_noxref_4_c_473_n N_noxref_6_c_833_n ) capacitor c=7.52994e-19 \
 //x=7.77 //y=2.085 //x2=6.775 //y2=3.33
cc_435 ( N_noxref_4_c_455_n N_noxref_6_c_773_n ) capacitor c=0.023629f \
 //x=7.655 //y=2.59 //x2=6.66 //y2=2.085
cc_436 ( N_noxref_4_c_473_n N_noxref_6_c_773_n ) capacitor c=0.0240469f \
 //x=7.77 //y=2.085 //x2=6.66 //y2=2.085
cc_437 ( N_noxref_4_c_545_p N_noxref_6_c_773_n ) capacitor c=0.00251238f \
 //x=7.435 //y=1.92 //x2=6.66 //y2=2.085
cc_438 ( N_noxref_4_c_473_n N_noxref_6_c_774_n ) capacitor c=0.00201026f \
 //x=7.77 //y=2.085 //x2=9.62 //y2=3.33
cc_439 ( N_noxref_4_c_555_p N_noxref_6_c_780_n ) capacitor c=4.86506e-19 \
 //x=7.435 //y=0.91 //x2=6.465 //y2=0.87
cc_440 ( N_noxref_4_c_555_p N_noxref_6_c_782_n ) capacitor c=0.00152104f \
 //x=7.435 //y=0.91 //x2=6.465 //y2=1.215
cc_441 ( N_noxref_4_c_556_p N_noxref_6_c_783_n ) capacitor c=0.00109982f \
 //x=7.435 //y=1.255 //x2=6.465 //y2=1.525
cc_442 ( N_noxref_4_c_557_p N_noxref_6_c_783_n ) capacitor c=9.57794e-19 \
 //x=7.435 //y=1.565 //x2=6.465 //y2=1.525
cc_443 ( N_noxref_4_c_455_n N_noxref_6_c_784_n ) capacitor c=0.00523252f \
 //x=7.655 //y=2.59 //x2=6.465 //y2=1.92
cc_444 ( N_noxref_4_c_473_n N_noxref_6_c_784_n ) capacitor c=0.00220284f \
 //x=7.77 //y=2.085 //x2=6.465 //y2=1.92
cc_445 ( N_noxref_4_c_557_p N_noxref_6_c_784_n ) capacitor c=0.00662747f \
 //x=7.435 //y=1.565 //x2=6.465 //y2=1.92
cc_446 ( N_noxref_4_c_545_p N_noxref_6_c_784_n ) capacitor c=0.012079f \
 //x=7.435 //y=1.92 //x2=6.465 //y2=1.92
cc_447 ( N_noxref_4_c_555_p N_noxref_6_c_787_n ) capacitor c=0.0157772f \
 //x=7.435 //y=0.91 //x2=6.995 //y2=0.87
cc_448 ( N_noxref_4_c_561_p N_noxref_6_c_787_n ) capacitor c=0.00124821f \
 //x=7.965 //y=0.91 //x2=6.995 //y2=0.87
cc_449 ( N_noxref_4_c_556_p N_noxref_6_c_789_n ) capacitor c=0.0117362f \
 //x=7.435 //y=1.255 //x2=6.995 //y2=1.215
cc_450 ( N_noxref_4_c_557_p N_noxref_6_c_789_n ) capacitor c=0.00862358f \
 //x=7.435 //y=1.565 //x2=6.995 //y2=1.215
cc_451 ( N_noxref_4_c_547_p N_noxref_6_c_789_n ) capacitor c=0.00200715f \
 //x=7.965 //y=1.255 //x2=6.995 //y2=1.215
cc_452 ( N_noxref_4_c_455_n N_noxref_7_c_938_n ) capacitor c=0.300234f \
 //x=7.655 //y=2.59 //x2=10.245 //y2=2.96
cc_453 ( N_noxref_4_c_473_n N_noxref_7_c_938_n ) capacitor c=0.0176337f \
 //x=7.77 //y=2.085 //x2=10.245 //y2=2.96
cc_454 ( N_noxref_4_c_455_n N_noxref_7_c_991_n ) capacitor c=0.0290321f \
 //x=7.655 //y=2.59 //x2=4.555 //y2=2.96
cc_455 ( N_noxref_4_c_473_n N_noxref_7_c_962_n ) capacitor c=0.01781f //x=7.77 \
 //y=2.085 //x2=10.245 //y2=4.44
cc_456 ( N_noxref_4_c_540_p N_noxref_7_c_962_n ) capacitor c=0.0105048f \
 //x=7.77 //y=4.7 //x2=10.245 //y2=4.44
cc_457 ( N_noxref_4_c_473_n N_noxref_7_c_970_n ) capacitor c=9.41499e-19 \
 //x=7.77 //y=2.085 //x2=6.775 //y2=4.44
cc_458 ( N_noxref_4_c_455_n N_noxref_7_c_945_n ) capacitor c=0.0210072f \
 //x=7.655 //y=2.59 //x2=4.44 //y2=2.085
cc_459 ( N_noxref_4_c_470_n N_noxref_7_c_945_n ) capacitor c=2.14844e-19 \
 //x=1.48 //y=2.59 //x2=4.44 //y2=2.085
cc_460 ( N_noxref_4_c_473_n N_noxref_7_c_972_n ) capacitor c=0.0082518f \
 //x=7.77 //y=2.085 //x2=6.66 //y2=4.44
cc_461 ( N_noxref_4_c_540_p N_noxref_7_c_972_n ) capacitor c=0.00226398f \
 //x=7.77 //y=4.7 //x2=6.66 //y2=4.44
cc_462 ( N_noxref_4_M14_noxref_g N_noxref_7_M12_noxref_g ) capacitor \
 c=0.0100243f //x=7.44 //y=6.02 //x2=6.56 //y2=6.02
cc_463 ( N_noxref_4_M14_noxref_g N_noxref_7_M13_noxref_g ) capacitor \
 c=0.0610135f //x=7.44 //y=6.02 //x2=7 //y2=6.02
cc_464 ( N_noxref_4_M15_noxref_g N_noxref_7_M13_noxref_g ) capacitor \
 c=0.0094155f //x=7.88 //y=6.02 //x2=7 //y2=6.02
cc_465 ( N_noxref_4_c_455_n N_noxref_7_c_1002_n ) capacitor c=0.0077643f \
 //x=7.655 //y=2.59 //x2=4.105 //y2=1.92
cc_466 ( N_noxref_4_c_473_n N_noxref_7_c_990_n ) capacitor c=0.0022916f \
 //x=7.77 //y=2.085 //x2=6.66 //y2=4.7
cc_467 ( N_noxref_4_c_540_p N_noxref_7_c_990_n ) capacitor c=0.066749f \
 //x=7.77 //y=4.7 //x2=6.66 //y2=4.7
cc_468 ( N_noxref_4_c_455_n N_noxref_8_c_1111_n ) capacitor c=0.00649037f \
 //x=7.655 //y=2.59 //x2=3.805 //y2=5.205
cc_469 ( N_noxref_4_c_455_n N_noxref_9_c_1151_n ) capacitor c=0.00446497f \
 //x=7.655 //y=2.59 //x2=2.915 //y2=1.5
cc_470 ( N_noxref_4_c_455_n N_noxref_9_c_1152_n ) capacitor c=0.0162406f \
 //x=7.655 //y=2.59 //x2=3.8 //y2=1.585
cc_471 ( N_noxref_4_c_455_n N_noxref_9_c_1160_n ) capacitor c=0.00435275f \
 //x=7.655 //y=2.59 //x2=3.885 //y2=1.5
cc_472 ( N_noxref_4_c_455_n N_noxref_9_c_1161_n ) capacitor c=0.00192639f \
 //x=7.655 //y=2.59 //x2=4.77 //y2=0.535
cc_473 ( N_noxref_4_c_455_n N_noxref_9_M1_noxref_s ) capacitor c=8.27974e-19 \
 //x=7.655 //y=2.59 //x2=2.78 //y2=0.37
cc_474 ( N_noxref_4_M14_noxref_g N_noxref_10_c_1203_n ) capacitor c=0.0170604f \
 //x=7.44 //y=6.02 //x2=7.135 //y2=5.205
cc_475 ( N_noxref_4_M14_noxref_g N_noxref_10_c_1209_n ) capacitor c=0.0144401f \
 //x=7.44 //y=6.02 //x2=8.015 //y2=6.905
cc_476 ( N_noxref_4_M15_noxref_g N_noxref_10_c_1209_n ) capacitor c=0.0163317f \
 //x=7.88 //y=6.02 //x2=8.015 //y2=6.905
cc_477 ( N_noxref_4_M15_noxref_g N_noxref_10_M15_noxref_d ) capacitor \
 c=0.0351101f //x=7.88 //y=6.02 //x2=7.955 //y2=5.02
cc_478 ( N_noxref_4_c_455_n N_noxref_11_c_1270_n ) capacitor c=0.00446497f \
 //x=7.655 //y=2.59 //x2=6.245 //y2=1.5
cc_479 ( N_noxref_4_c_455_n N_noxref_11_c_1246_n ) capacitor c=0.0162828f \
 //x=7.655 //y=2.59 //x2=7.13 //y2=1.585
cc_480 ( N_noxref_4_c_455_n N_noxref_11_c_1254_n ) capacitor c=0.00446497f \
 //x=7.655 //y=2.59 //x2=7.215 //y2=1.5
cc_481 ( N_noxref_4_c_557_p N_noxref_11_c_1254_n ) capacitor c=0.00628626f \
 //x=7.435 //y=1.565 //x2=7.215 //y2=1.5
cc_482 ( N_noxref_4_c_455_n N_noxref_11_c_1255_n ) capacitor c=0.00230651f \
 //x=7.655 //y=2.59 //x2=8.1 //y2=0.535
cc_483 ( N_noxref_4_c_555_p N_noxref_11_c_1255_n ) capacitor c=0.0197911f \
 //x=7.435 //y=0.91 //x2=8.1 //y2=0.535
cc_484 ( N_noxref_4_c_561_p N_noxref_11_c_1255_n ) capacitor c=0.00655813f \
 //x=7.965 //y=0.91 //x2=8.1 //y2=0.535
cc_485 ( N_noxref_4_c_555_p N_noxref_11_M3_noxref_s ) capacitor c=0.00628626f \
 //x=7.435 //y=0.91 //x2=6.11 //y2=0.37
cc_486 ( N_noxref_4_c_561_p N_noxref_11_M3_noxref_s ) capacitor c=0.0143002f \
 //x=7.965 //y=0.91 //x2=6.11 //y2=0.37
cc_487 ( N_noxref_4_c_547_p N_noxref_11_M3_noxref_s ) capacitor c=0.00290153f \
 //x=7.965 //y=1.255 //x2=6.11 //y2=0.37
cc_488 ( N_noxref_5_c_653_n N_noxref_6_c_794_n ) capacitor c=0.304758f \
 //x=8.025 //y=3.7 //x2=9.505 //y2=4.07
cc_489 ( N_noxref_5_c_651_n N_noxref_6_c_794_n ) capacitor c=0.0293663f \
 //x=4.925 //y=3.7 //x2=9.505 //y2=4.07
cc_490 ( N_noxref_5_c_636_n N_noxref_6_c_794_n ) capacitor c=0.00431193f \
 //x=4.725 //y=5.205 //x2=9.505 //y2=4.07
cc_491 ( N_noxref_5_c_625_n N_noxref_6_c_794_n ) capacitor c=0.0229481f \
 //x=4.81 //y=3.7 //x2=9.505 //y2=4.07
cc_492 ( N_noxref_5_c_628_n N_noxref_6_c_794_n ) capacitor c=0.0181107f \
 //x=8.14 //y=3.7 //x2=9.505 //y2=4.07
cc_493 ( N_noxref_5_c_636_n N_noxref_6_c_799_n ) capacitor c=0.00102585f \
 //x=4.725 //y=5.205 //x2=4.555 //y2=4.07
cc_494 ( N_noxref_5_c_638_n N_noxref_6_c_799_n ) capacitor c=0.00142608f \
 //x=4.415 //y=5.205 //x2=4.555 //y2=4.07
cc_495 ( N_noxref_5_c_625_n N_noxref_6_c_799_n ) capacitor c=0.00168517f \
 //x=4.81 //y=3.7 //x2=4.555 //y2=4.07
cc_496 ( N_noxref_5_c_653_n N_noxref_6_c_831_n ) capacitor c=0.139118f \
 //x=8.025 //y=3.7 //x2=9.505 //y2=3.33
cc_497 ( N_noxref_5_c_628_n N_noxref_6_c_831_n ) capacitor c=0.0186917f \
 //x=8.14 //y=3.7 //x2=9.505 //y2=3.33
cc_498 ( N_noxref_5_c_653_n N_noxref_6_c_833_n ) capacitor c=0.0286715f \
 //x=8.025 //y=3.7 //x2=6.775 //y2=3.33
cc_499 ( N_noxref_5_c_625_n N_noxref_6_c_833_n ) capacitor c=0.00286172f \
 //x=4.81 //y=3.7 //x2=6.775 //y2=3.33
cc_500 ( N_noxref_5_c_638_n N_noxref_6_c_800_n ) capacitor c=0.0123412f \
 //x=4.415 //y=5.205 //x2=4.44 //y2=4.07
cc_501 ( N_noxref_5_c_625_n N_noxref_6_c_800_n ) capacitor c=0.0637046f \
 //x=4.81 //y=3.7 //x2=4.44 //y2=4.07
cc_502 ( N_noxref_5_c_653_n N_noxref_6_c_773_n ) capacitor c=0.00490264f \
 //x=8.025 //y=3.7 //x2=6.66 //y2=2.085
cc_503 ( N_noxref_5_c_625_n N_noxref_6_c_773_n ) capacitor c=0.00705097f \
 //x=4.81 //y=3.7 //x2=6.66 //y2=2.085
cc_504 ( N_noxref_5_c_628_n N_noxref_6_c_773_n ) capacitor c=0.00341764f \
 //x=8.14 //y=3.7 //x2=6.66 //y2=2.085
cc_505 ( N_noxref_5_c_653_n N_noxref_6_c_774_n ) capacitor c=0.00382062f \
 //x=8.025 //y=3.7 //x2=9.62 //y2=3.33
cc_506 ( N_noxref_5_c_628_n N_noxref_6_c_776_n ) capacitor c=0.0155349f \
 //x=8.14 //y=3.7 //x2=9.705 //y2=2.08
cc_507 ( N_noxref_5_c_638_n N_noxref_6_M10_noxref_g ) capacitor c=0.0132788f \
 //x=4.415 //y=5.205 //x2=4.11 //y2=6.02
cc_508 ( N_noxref_5_c_636_n N_noxref_6_M11_noxref_g ) capacitor c=0.0187432f \
 //x=4.725 //y=5.205 //x2=4.55 //y2=6.02
cc_509 ( N_noxref_5_M10_noxref_d N_noxref_6_M11_noxref_g ) capacitor \
 c=0.0136385f //x=4.185 //y=5.02 //x2=4.55 //y2=6.02
cc_510 ( N_noxref_5_c_636_n N_noxref_6_c_826_n ) capacitor c=0.00161455f \
 //x=4.725 //y=5.205 //x2=4.44 //y2=4.7
cc_511 ( N_noxref_5_c_638_n N_noxref_6_c_826_n ) capacitor c=0.00557817f \
 //x=4.415 //y=5.205 //x2=4.44 //y2=4.7
cc_512 ( N_noxref_5_c_625_n N_noxref_6_c_826_n ) capacitor c=0.0232466f \
 //x=4.81 //y=3.7 //x2=4.44 //y2=4.7
cc_513 ( N_noxref_5_c_628_n N_noxref_6_M5_noxref_d ) capacitor c=2.78794e-19 \
 //x=8.14 //y=3.7 //x2=9.795 //y2=0.91
cc_514 ( N_noxref_5_c_628_n N_noxref_6_M16_noxref_d ) capacitor c=7.99492e-19 \
 //x=8.14 //y=3.7 //x2=9.84 //y2=5.02
cc_515 ( N_noxref_5_c_653_n N_noxref_7_c_938_n ) capacitor c=0.085016f \
 //x=8.025 //y=3.7 //x2=10.245 //y2=2.96
cc_516 ( N_noxref_5_c_651_n N_noxref_7_c_938_n ) capacitor c=0.0133597f \
 //x=4.925 //y=3.7 //x2=10.245 //y2=2.96
cc_517 ( N_noxref_5_c_625_n N_noxref_7_c_938_n ) capacitor c=0.0192028f \
 //x=4.81 //y=3.7 //x2=10.245 //y2=2.96
cc_518 ( N_noxref_5_c_626_n N_noxref_7_c_938_n ) capacitor c=0.00229609f \
 //x=8.055 //y=1.655 //x2=10.245 //y2=2.96
cc_519 ( N_noxref_5_c_628_n N_noxref_7_c_938_n ) capacitor c=0.0214051f \
 //x=8.14 //y=3.7 //x2=10.245 //y2=2.96
cc_520 ( N_noxref_5_c_625_n N_noxref_7_c_991_n ) capacitor c=0.00244604f \
 //x=4.81 //y=3.7 //x2=4.555 //y2=2.96
cc_521 ( N_noxref_5_c_653_n N_noxref_7_c_962_n ) capacitor c=0.0110294f \
 //x=8.025 //y=3.7 //x2=10.245 //y2=4.44
cc_522 ( N_noxref_5_c_641_n N_noxref_7_c_962_n ) capacitor c=0.00665427f \
 //x=8.055 //y=5.205 //x2=10.245 //y2=4.44
cc_523 ( N_noxref_5_c_643_n N_noxref_7_c_962_n ) capacitor c=0.00351988f \
 //x=7.745 //y=5.205 //x2=10.245 //y2=4.44
cc_524 ( N_noxref_5_c_628_n N_noxref_7_c_962_n ) capacitor c=0.0186407f \
 //x=8.14 //y=3.7 //x2=10.245 //y2=4.44
cc_525 ( N_noxref_5_c_653_n N_noxref_7_c_970_n ) capacitor c=0.00181512f \
 //x=8.025 //y=3.7 //x2=6.775 //y2=4.44
cc_526 ( N_noxref_5_c_659_n N_noxref_7_c_945_n ) capacitor c=0.0163885f \
 //x=4.455 //y=1.655 //x2=4.44 //y2=2.085
cc_527 ( N_noxref_5_c_625_n N_noxref_7_c_945_n ) capacitor c=0.0790313f \
 //x=4.81 //y=3.7 //x2=4.44 //y2=2.085
cc_528 ( N_noxref_5_c_625_n N_noxref_7_c_972_n ) capacitor c=7.44407e-19 \
 //x=4.81 //y=3.7 //x2=6.66 //y2=4.44
cc_529 ( N_noxref_5_c_628_n N_noxref_7_c_972_n ) capacitor c=0.00138227f \
 //x=8.14 //y=3.7 //x2=6.66 //y2=4.44
cc_530 ( N_noxref_5_c_628_n N_noxref_7_c_947_n ) capacitor c=0.0015583f \
 //x=8.14 //y=3.7 //x2=10.36 //y2=2.085
cc_531 ( N_noxref_5_M2_noxref_d N_noxref_7_c_994_n ) capacitor c=0.00217566f \
 //x=4.18 //y=0.91 //x2=4.105 //y2=0.91
cc_532 ( N_noxref_5_M2_noxref_d N_noxref_7_c_997_n ) capacitor c=0.0034598f \
 //x=4.18 //y=0.91 //x2=4.105 //y2=1.255
cc_533 ( N_noxref_5_M2_noxref_d N_noxref_7_c_999_n ) capacitor c=0.00522042f \
 //x=4.18 //y=0.91 //x2=4.105 //y2=1.565
cc_534 ( N_noxref_5_c_624_n N_noxref_7_c_1002_n ) capacitor c=0.00363601f \
 //x=4.725 //y=1.655 //x2=4.105 //y2=1.92
cc_535 ( N_noxref_5_c_659_n N_noxref_7_c_1002_n ) capacitor c=0.00637984f \
 //x=4.455 //y=1.655 //x2=4.105 //y2=1.92
cc_536 ( N_noxref_5_c_625_n N_noxref_7_c_1002_n ) capacitor c=0.0185661f \
 //x=4.81 //y=3.7 //x2=4.105 //y2=1.92
cc_537 ( N_noxref_5_M2_noxref_d N_noxref_7_c_1002_n ) capacitor c=0.00643086f \
 //x=4.18 //y=0.91 //x2=4.105 //y2=1.92
cc_538 ( N_noxref_5_M2_noxref_d N_noxref_7_c_1045_n ) capacitor c=0.00241053f \
 //x=4.18 //y=0.91 //x2=4.48 //y2=0.755
cc_539 ( N_noxref_5_c_624_n N_noxref_7_c_1046_n ) capacitor c=0.00196666f \
 //x=4.725 //y=1.655 //x2=4.48 //y2=1.41
cc_540 ( N_noxref_5_M2_noxref_d N_noxref_7_c_1046_n ) capacitor c=0.0124466f \
 //x=4.18 //y=0.91 //x2=4.48 //y2=1.41
cc_541 ( N_noxref_5_M2_noxref_d N_noxref_7_c_1004_n ) capacitor c=0.00132245f \
 //x=4.18 //y=0.91 //x2=4.635 //y2=0.91
cc_542 ( N_noxref_5_c_624_n N_noxref_7_c_1005_n ) capacitor c=0.00423452f \
 //x=4.725 //y=1.655 //x2=4.635 //y2=1.255
cc_543 ( N_noxref_5_M2_noxref_d N_noxref_7_c_1005_n ) capacitor c=0.00566463f \
 //x=4.18 //y=0.91 //x2=4.635 //y2=1.255
cc_544 ( N_noxref_5_c_638_n N_noxref_8_c_1111_n ) capacitor c=0.0348754f \
 //x=4.415 //y=5.205 //x2=3.805 //y2=5.205
cc_545 ( N_noxref_5_c_636_n N_noxref_8_c_1118_n ) capacitor c=0.0015978f \
 //x=4.725 //y=5.205 //x2=4.685 //y2=6.905
cc_546 ( N_noxref_5_M10_noxref_d N_noxref_8_c_1118_n ) capacitor c=0.01159f \
 //x=4.185 //y=5.02 //x2=4.685 //y2=6.905
cc_547 ( N_noxref_5_M10_noxref_d N_noxref_8_M8_noxref_s ) capacitor \
 c=0.00107541f //x=4.185 //y=5.02 //x2=2.875 //y2=5.02
cc_548 ( N_noxref_5_M10_noxref_d N_noxref_8_M9_noxref_d ) capacitor \
 c=0.0348754f //x=4.185 //y=5.02 //x2=3.745 //y2=5.02
cc_549 ( N_noxref_5_c_636_n N_noxref_8_M11_noxref_d ) capacitor c=0.0154556f \
 //x=4.725 //y=5.205 //x2=4.625 //y2=5.02
cc_550 ( N_noxref_5_M10_noxref_d N_noxref_8_M11_noxref_d ) capacitor \
 c=0.0458293f //x=4.185 //y=5.02 //x2=4.625 //y2=5.02
cc_551 ( N_noxref_5_c_659_n N_noxref_9_c_1151_n ) capacitor c=2.94752e-19 \
 //x=4.455 //y=1.655 //x2=2.915 //y2=1.5
cc_552 ( N_noxref_5_c_659_n N_noxref_9_c_1160_n ) capacitor c=0.0200666f \
 //x=4.455 //y=1.655 //x2=3.885 //y2=1.5
cc_553 ( N_noxref_5_c_624_n N_noxref_9_c_1161_n ) capacitor c=0.00457193f \
 //x=4.725 //y=1.655 //x2=4.77 //y2=0.535
cc_554 ( N_noxref_5_M2_noxref_d N_noxref_9_c_1161_n ) capacitor c=0.0113706f \
 //x=4.18 //y=0.91 //x2=4.77 //y2=0.535
cc_555 ( N_noxref_5_c_624_n N_noxref_9_M1_noxref_s ) capacitor c=0.0141081f \
 //x=4.725 //y=1.655 //x2=2.78 //y2=0.37
cc_556 ( N_noxref_5_M2_noxref_d N_noxref_9_M1_noxref_s ) capacitor \
 c=0.0436902f //x=4.18 //y=0.91 //x2=2.78 //y2=0.37
cc_557 ( N_noxref_5_c_643_n N_noxref_10_c_1203_n ) capacitor c=0.0348754f \
 //x=7.745 //y=5.205 //x2=7.135 //y2=5.205
cc_558 ( N_noxref_5_c_636_n N_noxref_10_c_1208_n ) capacitor c=2.91997e-19 \
 //x=4.725 //y=5.205 //x2=6.425 //y2=5.205
cc_559 ( N_noxref_5_c_641_n N_noxref_10_c_1209_n ) capacitor c=0.00157156f \
 //x=8.055 //y=5.205 //x2=8.015 //y2=6.905
cc_560 ( N_noxref_5_M14_noxref_d N_noxref_10_c_1209_n ) capacitor c=0.011538f \
 //x=7.515 //y=5.02 //x2=8.015 //y2=6.905
cc_561 ( N_noxref_5_M10_noxref_d N_noxref_10_M12_noxref_s ) capacitor \
 c=4.36987e-19 //x=4.185 //y=5.02 //x2=6.205 //y2=5.02
cc_562 ( N_noxref_5_M14_noxref_d N_noxref_10_M12_noxref_s ) capacitor \
 c=0.00107541f //x=7.515 //y=5.02 //x2=6.205 //y2=5.02
cc_563 ( N_noxref_5_M14_noxref_d N_noxref_10_M13_noxref_d ) capacitor \
 c=0.0348754f //x=7.515 //y=5.02 //x2=7.075 //y2=5.02
cc_564 ( N_noxref_5_c_641_n N_noxref_10_M15_noxref_d ) capacitor c=0.0151538f \
 //x=8.055 //y=5.205 //x2=7.955 //y2=5.02
cc_565 ( N_noxref_5_M14_noxref_d N_noxref_10_M15_noxref_d ) capacitor \
 c=0.0458293f //x=7.515 //y=5.02 //x2=7.955 //y2=5.02
cc_566 ( N_noxref_5_c_624_n N_noxref_11_c_1270_n ) capacitor c=3.32751e-19 \
 //x=4.725 //y=1.655 //x2=6.245 //y2=1.5
cc_567 ( N_noxref_5_c_672_n N_noxref_11_c_1270_n ) capacitor c=2.94752e-19 \
 //x=7.785 //y=1.655 //x2=6.245 //y2=1.5
cc_568 ( N_noxref_5_c_672_n N_noxref_11_c_1254_n ) capacitor c=0.0202508f \
 //x=7.785 //y=1.655 //x2=7.215 //y2=1.5
cc_569 ( N_noxref_5_c_626_n N_noxref_11_c_1255_n ) capacitor c=0.00458523f \
 //x=8.055 //y=1.655 //x2=8.1 //y2=0.535
cc_570 ( N_noxref_5_M4_noxref_d N_noxref_11_c_1255_n ) capacitor c=0.0113663f \
 //x=7.51 //y=0.91 //x2=8.1 //y2=0.535
cc_571 ( N_noxref_5_c_626_n N_noxref_11_M3_noxref_s ) capacitor c=0.0143532f \
 //x=8.055 //y=1.655 //x2=6.11 //y2=0.37
cc_572 ( N_noxref_5_M4_noxref_d N_noxref_11_M3_noxref_s ) capacitor \
 c=0.0438744f //x=7.51 //y=0.91 //x2=6.11 //y2=0.37
cc_573 ( N_noxref_6_c_794_n N_noxref_7_c_938_n ) capacitor c=0.0166896f \
 //x=9.505 //y=4.07 //x2=10.245 //y2=2.96
cc_574 ( N_noxref_6_c_831_n N_noxref_7_c_938_n ) capacitor c=0.269397f \
 //x=9.505 //y=3.33 //x2=10.245 //y2=2.96
cc_575 ( N_noxref_6_c_833_n N_noxref_7_c_938_n ) capacitor c=0.0291219f \
 //x=6.775 //y=3.33 //x2=10.245 //y2=2.96
cc_576 ( N_noxref_6_c_773_n N_noxref_7_c_938_n ) capacitor c=0.0215791f \
 //x=6.66 //y=2.085 //x2=10.245 //y2=2.96
cc_577 ( N_noxref_6_c_774_n N_noxref_7_c_938_n ) capacitor c=0.0267634f \
 //x=9.62 //y=3.33 //x2=10.245 //y2=2.96
cc_578 ( N_noxref_6_c_775_n N_noxref_7_c_938_n ) capacitor c=0.00763858f \
 //x=9.905 //y=2.08 //x2=10.245 //y2=2.96
cc_579 ( N_noxref_6_c_804_n N_noxref_7_c_938_n ) capacitor c=0.00159282f \
 //x=9.9 //y=4.58 //x2=10.245 //y2=2.96
cc_580 ( N_noxref_6_c_799_n N_noxref_7_c_991_n ) capacitor c=0.00956028f \
 //x=4.555 //y=4.07 //x2=4.555 //y2=2.96
cc_581 ( N_noxref_6_c_800_n N_noxref_7_c_991_n ) capacitor c=2.06418e-19 \
 //x=4.44 //y=4.07 //x2=4.555 //y2=2.96
cc_582 ( N_noxref_6_c_794_n N_noxref_7_c_962_n ) capacitor c=0.267726f \
 //x=9.505 //y=4.07 //x2=10.245 //y2=4.44
cc_583 ( N_noxref_6_c_831_n N_noxref_7_c_962_n ) capacitor c=0.00450734f \
 //x=9.505 //y=3.33 //x2=10.245 //y2=4.44
cc_584 ( N_noxref_6_c_774_n N_noxref_7_c_962_n ) capacitor c=0.0131307f \
 //x=9.62 //y=3.33 //x2=10.245 //y2=4.44
cc_585 ( N_noxref_6_c_804_n N_noxref_7_c_962_n ) capacitor c=0.0204817f \
 //x=9.9 //y=4.58 //x2=10.245 //y2=4.44
cc_586 ( N_noxref_6_c_805_n N_noxref_7_c_962_n ) capacitor c=0.00582322f \
 //x=9.705 //y=4.58 //x2=10.245 //y2=4.44
cc_587 ( N_noxref_6_c_794_n N_noxref_7_c_970_n ) capacitor c=0.0286083f \
 //x=9.505 //y=4.07 //x2=6.775 //y2=4.44
cc_588 ( N_noxref_6_c_799_n N_noxref_7_c_945_n ) capacitor c=2.06418e-19 \
 //x=4.555 //y=4.07 //x2=4.44 //y2=2.085
cc_589 ( N_noxref_6_c_800_n N_noxref_7_c_945_n ) capacitor c=0.00912271f \
 //x=4.44 //y=4.07 //x2=4.44 //y2=2.085
cc_590 ( N_noxref_6_c_773_n N_noxref_7_c_945_n ) capacitor c=3.72011e-19 \
 //x=6.66 //y=2.085 //x2=4.44 //y2=2.085
cc_591 ( N_noxref_6_c_794_n N_noxref_7_c_972_n ) capacitor c=0.00480464f \
 //x=9.505 //y=4.07 //x2=6.66 //y2=4.44
cc_592 ( N_noxref_6_c_773_n N_noxref_7_c_972_n ) capacitor c=0.00883142f \
 //x=6.66 //y=2.085 //x2=6.66 //y2=4.44
cc_593 ( N_noxref_6_c_794_n N_noxref_7_c_947_n ) capacitor c=0.00642908f \
 //x=9.505 //y=4.07 //x2=10.36 //y2=2.085
cc_594 ( N_noxref_6_c_831_n N_noxref_7_c_947_n ) capacitor c=0.00598101f \
 //x=9.505 //y=3.33 //x2=10.36 //y2=2.085
cc_595 ( N_noxref_6_c_774_n N_noxref_7_c_947_n ) capacitor c=0.0642592f \
 //x=9.62 //y=3.33 //x2=10.36 //y2=2.085
cc_596 ( N_noxref_6_c_804_n N_noxref_7_c_947_n ) capacitor c=0.0265353f \
 //x=9.9 //y=4.58 //x2=10.36 //y2=2.085
cc_597 ( N_noxref_6_M5_noxref_d N_noxref_7_c_947_n ) capacitor c=0.0175773f \
 //x=9.795 //y=0.91 //x2=10.36 //y2=2.085
cc_598 ( N_noxref_6_M16_noxref_d N_noxref_7_M16_noxref_g ) capacitor \
 c=0.021902f //x=9.84 //y=5.02 //x2=9.765 //y2=6.02
cc_599 ( N_noxref_6_M16_noxref_d N_noxref_7_M17_noxref_g ) capacitor \
 c=0.0219309f //x=9.84 //y=5.02 //x2=10.205 //y2=6.02
cc_600 ( N_noxref_6_M5_noxref_d N_noxref_7_c_952_n ) capacitor c=0.00216577f \
 //x=9.795 //y=0.91 //x2=9.72 //y2=0.91
cc_601 ( N_noxref_6_c_775_n N_noxref_7_c_954_n ) capacitor c=0.0023507f \
 //x=9.905 //y=2.08 //x2=9.72 //y2=1.255
cc_602 ( N_noxref_6_M5_noxref_d N_noxref_7_c_954_n ) capacitor c=0.00599232f \
 //x=9.795 //y=0.91 //x2=9.72 //y2=1.255
cc_603 ( N_noxref_6_c_804_n N_noxref_7_c_1081_n ) capacitor c=0.00491319f \
 //x=9.9 //y=4.58 //x2=10.13 //y2=4.79
cc_604 ( N_noxref_6_M16_noxref_d N_noxref_7_c_1081_n ) capacitor c=0.0146106f \
 //x=9.84 //y=5.02 //x2=10.13 //y2=4.79
cc_605 ( N_noxref_6_c_805_n N_noxref_7_c_987_n ) capacitor c=0.00491319f \
 //x=9.705 //y=4.58 //x2=9.84 //y2=4.79
cc_606 ( N_noxref_6_M5_noxref_d N_noxref_7_c_955_n ) capacitor c=0.00220879f \
 //x=9.795 //y=0.91 //x2=10.095 //y2=0.755
cc_607 ( N_noxref_6_M5_noxref_d N_noxref_7_c_1085_n ) capacitor c=0.0138447f \
 //x=9.795 //y=0.91 //x2=10.095 //y2=1.41
cc_608 ( N_noxref_6_c_804_n N_noxref_7_c_988_n ) capacitor c=0.00941483f \
 //x=9.9 //y=4.58 //x2=10.205 //y2=4.865
cc_609 ( N_noxref_6_M16_noxref_d N_noxref_7_c_988_n ) capacitor c=0.00307344f \
 //x=9.84 //y=5.02 //x2=10.205 //y2=4.865
cc_610 ( N_noxref_6_M5_noxref_d N_noxref_7_c_956_n ) capacitor c=0.00220616f \
 //x=9.795 //y=0.91 //x2=10.25 //y2=0.91
cc_611 ( N_noxref_6_M5_noxref_d N_noxref_7_c_1089_n ) capacitor c=0.00347355f \
 //x=9.795 //y=0.91 //x2=10.25 //y2=1.255
cc_612 ( N_noxref_6_M5_noxref_d N_noxref_7_c_1090_n ) capacitor c=0.007449f \
 //x=9.795 //y=0.91 //x2=10.25 //y2=1.565
cc_613 ( N_noxref_6_M5_noxref_d N_noxref_7_c_958_n ) capacitor c=0.00957707f \
 //x=9.795 //y=0.91 //x2=10.25 //y2=1.92
cc_614 ( N_noxref_6_c_794_n N_noxref_7_c_990_n ) capacitor c=6.08197e-19 \
 //x=9.505 //y=4.07 //x2=6.66 //y2=4.7
cc_615 ( N_noxref_6_c_774_n N_noxref_7_c_959_n ) capacitor c=8.49451e-19 \
 //x=9.62 //y=3.33 //x2=10.25 //y2=2.085
cc_616 ( N_noxref_6_c_775_n N_noxref_7_c_959_n ) capacitor c=0.0167852f \
 //x=9.905 //y=2.08 //x2=10.25 //y2=2.085
cc_617 ( N_noxref_6_M10_noxref_g N_noxref_8_c_1111_n ) capacitor c=0.0170604f \
 //x=4.11 //y=6.02 //x2=3.805 //y2=5.205
cc_618 ( N_noxref_6_M10_noxref_g N_noxref_8_c_1118_n ) capacitor c=0.0150677f \
 //x=4.11 //y=6.02 //x2=4.685 //y2=6.905
cc_619 ( N_noxref_6_M11_noxref_g N_noxref_8_c_1118_n ) capacitor c=0.016333f \
 //x=4.55 //y=6.02 //x2=4.685 //y2=6.905
cc_620 ( N_noxref_6_M11_noxref_g N_noxref_8_M11_noxref_d ) capacitor \
 c=0.0351101f //x=4.55 //y=6.02 //x2=4.625 //y2=5.02
cc_621 ( N_noxref_6_c_794_n N_noxref_10_c_1208_n ) capacitor c=0.0060417f \
 //x=9.505 //y=4.07 //x2=6.425 //y2=5.205
cc_622 ( N_noxref_6_c_784_n N_noxref_11_c_1270_n ) capacitor c=0.0034165f \
 //x=6.465 //y=1.92 //x2=6.245 //y2=1.5
cc_623 ( N_noxref_6_c_773_n N_noxref_11_c_1246_n ) capacitor c=0.0113444f \
 //x=6.66 //y=2.085 //x2=7.13 //y2=1.585
cc_624 ( N_noxref_6_c_783_n N_noxref_11_c_1246_n ) capacitor c=0.00704065f \
 //x=6.465 //y=1.525 //x2=7.13 //y2=1.585
cc_625 ( N_noxref_6_c_784_n N_noxref_11_c_1246_n ) capacitor c=0.0185489f \
 //x=6.465 //y=1.92 //x2=7.13 //y2=1.585
cc_626 ( N_noxref_6_c_786_n N_noxref_11_c_1246_n ) capacitor c=0.00780802f \
 //x=6.84 //y=1.37 //x2=7.13 //y2=1.585
cc_627 ( N_noxref_6_c_789_n N_noxref_11_c_1246_n ) capacitor c=0.0034036f \
 //x=6.995 //y=1.215 //x2=7.13 //y2=1.585
cc_628 ( N_noxref_6_c_784_n N_noxref_11_c_1254_n ) capacitor c=6.71402e-19 \
 //x=6.465 //y=1.92 //x2=7.215 //y2=1.5
cc_629 ( N_noxref_6_c_780_n N_noxref_11_M3_noxref_s ) capacitor c=0.0326577f \
 //x=6.465 //y=0.87 //x2=6.11 //y2=0.37
cc_630 ( N_noxref_6_c_783_n N_noxref_11_M3_noxref_s ) capacitor c=3.48408e-19 \
 //x=6.465 //y=1.525 //x2=6.11 //y2=0.37
cc_631 ( N_noxref_6_c_787_n N_noxref_11_M3_noxref_s ) capacitor c=0.0120759f \
 //x=6.995 //y=0.87 //x2=6.11 //y2=0.37
cc_632 ( N_noxref_7_c_999_n N_noxref_9_c_1160_n ) capacitor c=0.00628626f \
 //x=4.105 //y=1.565 //x2=3.885 //y2=1.5
cc_633 ( N_noxref_7_c_994_n N_noxref_9_c_1161_n ) capacitor c=0.0197911f \
 //x=4.105 //y=0.91 //x2=4.77 //y2=0.535
cc_634 ( N_noxref_7_c_1004_n N_noxref_9_c_1161_n ) capacitor c=0.00655813f \
 //x=4.635 //y=0.91 //x2=4.77 //y2=0.535
cc_635 ( N_noxref_7_c_994_n N_noxref_9_M1_noxref_s ) capacitor c=0.00628626f \
 //x=4.105 //y=0.91 //x2=2.78 //y2=0.37
cc_636 ( N_noxref_7_c_1004_n N_noxref_9_M1_noxref_s ) capacitor c=0.0143002f \
 //x=4.635 //y=0.91 //x2=2.78 //y2=0.37
cc_637 ( N_noxref_7_c_1005_n N_noxref_9_M1_noxref_s ) capacitor c=0.00290153f \
 //x=4.635 //y=1.255 //x2=2.78 //y2=0.37
cc_638 ( N_noxref_7_c_962_n N_noxref_10_c_1203_n ) capacitor c=0.0172642f \
 //x=10.245 //y=4.44 //x2=7.135 //y2=5.205
cc_639 ( N_noxref_7_c_970_n N_noxref_10_c_1203_n ) capacitor c=0.00485884f \
 //x=6.775 //y=4.44 //x2=7.135 //y2=5.205
cc_640 ( N_noxref_7_c_972_n N_noxref_10_c_1203_n ) capacitor c=0.0111238f \
 //x=6.66 //y=4.44 //x2=7.135 //y2=5.205
cc_641 ( N_noxref_7_M12_noxref_g N_noxref_10_c_1203_n ) capacitor c=0.018644f \
 //x=6.56 //y=6.02 //x2=7.135 //y2=5.205
cc_642 ( N_noxref_7_M13_noxref_g N_noxref_10_c_1203_n ) capacitor c=0.0169648f \
 //x=7 //y=6.02 //x2=7.135 //y2=5.205
cc_643 ( N_noxref_7_c_990_n N_noxref_10_c_1203_n ) capacitor c=0.00531676f \
 //x=6.66 //y=4.7 //x2=7.135 //y2=5.205
cc_644 ( N_noxref_7_c_962_n N_noxref_10_c_1209_n ) capacitor c=0.00389598f \
 //x=10.245 //y=4.44 //x2=8.015 //y2=6.905
cc_645 ( N_noxref_7_M12_noxref_g N_noxref_10_M12_noxref_s ) capacitor \
 c=0.0441361f //x=6.56 //y=6.02 //x2=6.205 //y2=5.02
cc_646 ( N_noxref_7_M13_noxref_g N_noxref_10_M13_noxref_d ) capacitor \
 c=0.0170604f //x=7 //y=6.02 //x2=7.075 //y2=5.02
cc_647 ( N_noxref_7_c_938_n N_noxref_11_M3_noxref_s ) capacitor c=6.22885e-19 \
 //x=10.245 //y=2.96 //x2=6.11 //y2=0.37
cc_648 ( N_noxref_8_M11_noxref_d N_noxref_10_M12_noxref_s ) capacitor \
 c=0.00181587f //x=4.625 //y=5.02 //x2=6.205 //y2=5.02
cc_649 ( N_noxref_9_c_1164_n N_noxref_11_M3_noxref_s ) capacitor c=0.00174327f \
 //x=4.855 //y=0.62 //x2=6.11 //y2=0.37
