* SPICE3 file created from DFFX1.ext - technology: sky130A

.subckt DFFX1 Q QN D CLK VPB VNB
M1000 QN Q a_3072_73.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1001 VPB.t21 a_147_159.t5 a_1845_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPB.t23 a_147_159.t6 a_277_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t7 a_1845_1004.t5 a_147_159.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 QN a_277_1004.t7 VPB.t8 pshort w=2u l=0.15u
+  ad=1.16p pd=9.16u as=0p ps=0u
M1005 VNB a_599_943.t5 a_1740_73.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1006 VPB.t16 CLK a_277_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPB.t19 CLK a_147_159.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 QN Q VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VNB a_147_159.t13 a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t2 a_599_943.t6 a_277_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPB.t3 a_277_1004.t8 a_599_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 Q QN VPB.t15 pshort w=2u l=0.15u
+  ad=1.16p pd=9.16u as=0p ps=0u
M1013 VNB QN a_3738_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPB.t25 a_147_159.t7 Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1845_1004.t2 a_147_159.t8 VPB.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 VNB a_277_1004.t9 a_1074_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1017 Q a_147_159.t9 VPB.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_277_1004.t5 a_147_159.t11 VPB.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPB.t1 a_1305_383# a_599_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPB.t13 a_599_943.t7 a_1845_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_277_1004.t3 CLK VPB.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VNB a_277_1004.t10 a_3072_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_147_159.t2 CLK VPB.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPB.t5 a_277_1004.t11 QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q a_147_159.t12 a_3738_73.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1026 a_277_1004.t1 a_599_943.t8 VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_599_943.t3 a_277_1004.t12 VPB.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_147_159.t1 a_1845_1004.t6 VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPB.t11 Q QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPB.t14 QN Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 VNB a_1845_1004.t7 a_2406_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_599_943.t1 a_1305_383# VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1845_1004.t0 a_599_943.t10 VPB.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u






R0 a_147_159.n8 a_147_159.t6 512.525
R1 a_147_159.n6 a_147_159.t5 472.359
R2 a_147_159.n4 a_147_159.t7 472.359
R3 a_147_159.n6 a_147_159.t8 384.527
R4 a_147_159.n4 a_147_159.t9 384.527
R5 a_147_159.n8 a_147_159.t11 371.139
R6 a_147_159.n9 a_147_159.t13 324.268
R7 a_147_159.n7 a_147_159.t10 277.772
R8 a_147_159.n5 a_147_159.t12 277.772
R9 a_147_159.n14 a_147_159.n12 247.192
R10 a_147_159.n9 a_147_159.n8 119.654
R11 a_147_159.n12 a_147_159.n3 109.441
R12 a_147_159.n10 a_147_159.n9 82.484
R13 a_147_159.n11 a_147_159.n5 80.307
R14 a_147_159.n3 a_147_159.n2 76.002
R15 a_147_159.n10 a_147_159.n7 76
R16 a_147_159.n12 a_147_159.n11 76
R17 a_147_159.n7 a_147_159.n6 67.001
R18 a_147_159.n5 a_147_159.n4 67.001
R19 a_147_159.n14 a_147_159.n13 30
R20 a_147_159.n15 a_147_159.n0 24.383
R21 a_147_159.n15 a_147_159.n14 23.684
R22 a_147_159.n1 a_147_159.t3 14.282
R23 a_147_159.n1 a_147_159.t2 14.282
R24 a_147_159.n2 a_147_159.t0 14.282
R25 a_147_159.n2 a_147_159.t1 14.282
R26 a_147_159.n3 a_147_159.n1 12.85
R27 a_147_159.n11 a_147_159.n10 2.947
R28 a_1845_1004.n4 a_1845_1004.t5 480.392
R29 a_1845_1004.n4 a_1845_1004.t6 403.272
R30 a_1845_1004.n5 a_1845_1004.t7 266.974
R31 a_1845_1004.n8 a_1845_1004.n6 194.086
R32 a_1845_1004.n6 a_1845_1004.n3 162.547
R33 a_1845_1004.n6 a_1845_1004.n5 153.315
R34 a_1845_1004.n5 a_1845_1004.n4 108.494
R35 a_1845_1004.n3 a_1845_1004.n2 76.002
R36 a_1845_1004.n8 a_1845_1004.n7 30
R37 a_1845_1004.n9 a_1845_1004.n0 24.383
R38 a_1845_1004.n9 a_1845_1004.n8 23.684
R39 a_1845_1004.n1 a_1845_1004.t4 14.282
R40 a_1845_1004.n1 a_1845_1004.t2 14.282
R41 a_1845_1004.n2 a_1845_1004.t1 14.282
R42 a_1845_1004.n2 a_1845_1004.t0 14.282
R43 a_1845_1004.n3 a_1845_1004.n1 12.85
R44 VPB VPB.n413 126.832
R45 VPB.n40 VPB.n38 94.117
R46 VPB.n355 VPB.n353 94.117
R47 VPB.n294 VPB.n292 94.117
R48 VPB.n132 VPB.n130 94.117
R49 VPB.n247 VPB.n245 94.117
R50 VPB.n50 VPB.n49 80.104
R51 VPB.n298 VPB.n82 76
R52 VPB.n208 VPB.n207 76
R53 VPB.n213 VPB.n212 76
R54 VPB.n218 VPB.n217 76
R55 VPB.n222 VPB.n221 76
R56 VPB.n249 VPB.n248 76
R57 VPB.n254 VPB.n253 76
R58 VPB.n259 VPB.n258 76
R59 VPB.n266 VPB.n265 76
R60 VPB.n271 VPB.n270 76
R61 VPB.n276 VPB.n275 76
R62 VPB.n281 VPB.n280 76
R63 VPB.n295 VPB.n291 76
R64 VPB.n304 VPB.n303 76
R65 VPB.n311 VPB.n310 76
R66 VPB.n316 VPB.n315 76
R67 VPB.n321 VPB.n320 76
R68 VPB.n326 VPB.n325 76
R69 VPB.n330 VPB.n329 76
R70 VPB.n357 VPB.n356 76
R71 VPB.n362 VPB.n361 76
R72 VPB.n367 VPB.n366 76
R73 VPB.n374 VPB.n373 76
R74 VPB.n379 VPB.n378 76
R75 VPB.n384 VPB.n383 76
R76 VPB.n389 VPB.n388 76
R77 VPB.n393 VPB.n392 76
R78 VPB.n406 VPB.n405 76
R79 VPB.n72 VPB.n71 75.654
R80 VPB.n22 VPB.n21 61.764
R81 VPB.n337 VPB.n336 61.764
R82 VPB.n89 VPB.n88 61.764
R83 VPB.n111 VPB.n110 61.764
R84 VPB.n229 VPB.n228 61.764
R85 VPB.n78 VPB.t22 55.106
R86 VPB.n385 VPB.t10 55.106
R87 VPB.n322 VPB.t9 55.106
R88 VPB.n155 VPB.t6 55.106
R89 VPB.n277 VPB.t8 55.106
R90 VPB.n214 VPB.t15 55.106
R91 VPB.n45 VPB.t2 55.106
R92 VPB.n358 VPB.t1 55.106
R93 VPB.n299 VPB.t21 55.106
R94 VPB.n137 VPB.t19 55.106
R95 VPB.n250 VPB.t11 55.106
R96 VPB.n197 VPB.t25 55.106
R97 VPB.n194 VPB.n193 48.952
R98 VPB.n256 VPB.n255 48.952
R99 VPB.n139 VPB.n138 48.952
R100 VPB.n301 VPB.n300 48.952
R101 VPB.n364 VPB.n363 48.952
R102 VPB.n54 VPB.n53 48.952
R103 VPB.n210 VPB.n209 44.502
R104 VPB.n273 VPB.n272 44.502
R105 VPB.n152 VPB.n151 44.502
R106 VPB.n318 VPB.n317 44.502
R107 VPB.n381 VPB.n380 44.502
R108 VPB.n68 VPB.n67 44.502
R109 VPB.n66 VPB.n14 40.824
R110 VPB.n57 VPB.n15 40.824
R111 VPB.n369 VPB.n368 40.824
R112 VPB.n306 VPB.n305 40.824
R113 VPB.n146 VPB.n104 40.824
R114 VPB.n261 VPB.n260 40.824
R115 VPB.n188 VPB.n187 40.824
R116 VPB.n202 VPB.n201 35.116
R117 VPB.n410 VPB.n406 20.452
R118 VPB.n186 VPB.n183 20.452
R119 VPB.n190 VPB.n189 17.801
R120 VPB.n263 VPB.n262 17.801
R121 VPB.n143 VPB.n142 17.801
R122 VPB.n308 VPB.n307 17.801
R123 VPB.n371 VPB.n370 17.801
R124 VPB.n59 VPB.n58 17.801
R125 VPB.n14 VPB.t17 14.282
R126 VPB.n14 VPB.t23 14.282
R127 VPB.n15 VPB.t4 14.282
R128 VPB.n15 VPB.t16 14.282
R129 VPB.n368 VPB.t0 14.282
R130 VPB.n368 VPB.t3 14.282
R131 VPB.n305 VPB.t20 14.282
R132 VPB.n305 VPB.t13 14.282
R133 VPB.n104 VPB.t18 14.282
R134 VPB.n104 VPB.t7 14.282
R135 VPB.n260 VPB.t12 14.282
R136 VPB.n260 VPB.t5 14.282
R137 VPB.n187 VPB.t24 14.282
R138 VPB.n187 VPB.t14 14.282
R139 VPB.n186 VPB.n185 13.653
R140 VPB.n185 VPB.n184 13.653
R141 VPB.n200 VPB.n199 13.653
R142 VPB.n199 VPB.n198 13.653
R143 VPB.n196 VPB.n195 13.653
R144 VPB.n195 VPB.n194 13.653
R145 VPB.n192 VPB.n191 13.653
R146 VPB.n191 VPB.n190 13.653
R147 VPB.n207 VPB.n206 13.653
R148 VPB.n206 VPB.n205 13.653
R149 VPB.n212 VPB.n211 13.653
R150 VPB.n211 VPB.n210 13.653
R151 VPB.n217 VPB.n216 13.653
R152 VPB.n216 VPB.n215 13.653
R153 VPB.n221 VPB.n220 13.653
R154 VPB.n220 VPB.n219 13.653
R155 VPB.n248 VPB.n247 13.653
R156 VPB.n247 VPB.n246 13.653
R157 VPB.n253 VPB.n252 13.653
R158 VPB.n252 VPB.n251 13.653
R159 VPB.n258 VPB.n257 13.653
R160 VPB.n257 VPB.n256 13.653
R161 VPB.n265 VPB.n264 13.653
R162 VPB.n264 VPB.n263 13.653
R163 VPB.n270 VPB.n269 13.653
R164 VPB.n269 VPB.n268 13.653
R165 VPB.n275 VPB.n274 13.653
R166 VPB.n274 VPB.n273 13.653
R167 VPB.n280 VPB.n279 13.653
R168 VPB.n279 VPB.n278 13.653
R169 VPB.n128 VPB.n127 13.653
R170 VPB.n127 VPB.n126 13.653
R171 VPB.n133 VPB.n132 13.653
R172 VPB.n132 VPB.n131 13.653
R173 VPB.n136 VPB.n135 13.653
R174 VPB.n135 VPB.n134 13.653
R175 VPB.n141 VPB.n140 13.653
R176 VPB.n140 VPB.n139 13.653
R177 VPB.n145 VPB.n144 13.653
R178 VPB.n144 VPB.n143 13.653
R179 VPB.n150 VPB.n149 13.653
R180 VPB.n149 VPB.n148 13.653
R181 VPB.n154 VPB.n153 13.653
R182 VPB.n153 VPB.n152 13.653
R183 VPB.n158 VPB.n157 13.653
R184 VPB.n157 VPB.n156 13.653
R185 VPB.n161 VPB.n160 13.653
R186 VPB.n160 VPB.n159 13.653
R187 VPB.n295 VPB.n294 13.653
R188 VPB.n294 VPB.n293 13.653
R189 VPB.n298 VPB.n297 13.653
R190 VPB.n297 VPB.n296 13.653
R191 VPB.n303 VPB.n302 13.653
R192 VPB.n302 VPB.n301 13.653
R193 VPB.n310 VPB.n309 13.653
R194 VPB.n309 VPB.n308 13.653
R195 VPB.n315 VPB.n314 13.653
R196 VPB.n314 VPB.n313 13.653
R197 VPB.n320 VPB.n319 13.653
R198 VPB.n319 VPB.n318 13.653
R199 VPB.n325 VPB.n324 13.653
R200 VPB.n324 VPB.n323 13.653
R201 VPB.n329 VPB.n328 13.653
R202 VPB.n328 VPB.n327 13.653
R203 VPB.n356 VPB.n355 13.653
R204 VPB.n355 VPB.n354 13.653
R205 VPB.n361 VPB.n360 13.653
R206 VPB.n360 VPB.n359 13.653
R207 VPB.n366 VPB.n365 13.653
R208 VPB.n365 VPB.n364 13.653
R209 VPB.n373 VPB.n372 13.653
R210 VPB.n372 VPB.n371 13.653
R211 VPB.n378 VPB.n377 13.653
R212 VPB.n377 VPB.n376 13.653
R213 VPB.n383 VPB.n382 13.653
R214 VPB.n382 VPB.n381 13.653
R215 VPB.n388 VPB.n387 13.653
R216 VPB.n387 VPB.n386 13.653
R217 VPB.n392 VPB.n391 13.653
R218 VPB.n391 VPB.n390 13.653
R219 VPB.n41 VPB.n40 13.653
R220 VPB.n40 VPB.n39 13.653
R221 VPB.n44 VPB.n43 13.653
R222 VPB.n43 VPB.n42 13.653
R223 VPB.n48 VPB.n47 13.653
R224 VPB.n47 VPB.n46 13.653
R225 VPB.n52 VPB.n51 13.653
R226 VPB.n51 VPB.n50 13.653
R227 VPB.n56 VPB.n55 13.653
R228 VPB.n55 VPB.n54 13.653
R229 VPB.n61 VPB.n60 13.653
R230 VPB.n60 VPB.n59 13.653
R231 VPB.n65 VPB.n64 13.653
R232 VPB.n64 VPB.n63 13.653
R233 VPB.n70 VPB.n69 13.653
R234 VPB.n69 VPB.n68 13.653
R235 VPB.n74 VPB.n73 13.653
R236 VPB.n73 VPB.n72 13.653
R237 VPB.n77 VPB.n76 13.653
R238 VPB.n76 VPB.n75 13.653
R239 VPB.n81 VPB.n80 13.653
R240 VPB.n80 VPB.n79 13.653
R241 VPB.n406 VPB.n0 13.653
R242 VPB VPB.n0 13.653
R243 VPB.n205 VPB.n204 13.35
R244 VPB.n268 VPB.n267 13.35
R245 VPB.n148 VPB.n147 13.35
R246 VPB.n313 VPB.n312 13.35
R247 VPB.n376 VPB.n375 13.35
R248 VPB.n63 VPB.n62 13.35
R249 VPB.n410 VPB.n409 13.276
R250 VPB.n409 VPB.n407 13.276
R251 VPB.n36 VPB.n18 13.276
R252 VPB.n18 VPB.n16 13.276
R253 VPB.n351 VPB.n333 13.276
R254 VPB.n333 VPB.n331 13.276
R255 VPB.n103 VPB.n85 13.276
R256 VPB.n85 VPB.n83 13.276
R257 VPB.n125 VPB.n107 13.276
R258 VPB.n107 VPB.n105 13.276
R259 VPB.n243 VPB.n225 13.276
R260 VPB.n225 VPB.n223 13.276
R261 VPB.n196 VPB.n192 13.276
R262 VPB.n248 VPB.n244 13.276
R263 VPB.n129 VPB.n128 13.276
R264 VPB.n133 VPB.n129 13.276
R265 VPB.n136 VPB.n133 13.276
R266 VPB.n145 VPB.n141 13.276
R267 VPB.n154 VPB.n150 13.276
R268 VPB.n161 VPB.n158 13.276
R269 VPB.n162 VPB.n161 13.276
R270 VPB.n295 VPB.n162 13.276
R271 VPB.n298 VPB.n295 13.276
R272 VPB.n356 VPB.n352 13.276
R273 VPB.n41 VPB.n37 13.276
R274 VPB.n44 VPB.n41 13.276
R275 VPB.n52 VPB.n48 13.276
R276 VPB.n56 VPB.n52 13.276
R277 VPB.n65 VPB.n61 13.276
R278 VPB.n74 VPB.n70 13.276
R279 VPB.n77 VPB.n74 13.276
R280 VPB.n406 VPB.n81 13.276
R281 VPB.n183 VPB.n165 13.276
R282 VPB.n165 VPB.n163 13.276
R283 VPB.n170 VPB.n168 12.796
R284 VPB.n170 VPB.n169 12.564
R285 VPB.n81 VPB.n78 12.558
R286 VPB.n45 VPB.n44 12.2
R287 VPB.n178 VPB.n177 12.198
R288 VPB.n174 VPB.n173 12.198
R289 VPB.n178 VPB.n175 12.198
R290 VPB.n197 VPB.n196 11.841
R291 VPB.n141 VPB.n137 11.841
R292 VPB.n303 VPB.n299 11.841
R293 VPB.n155 VPB.n154 11.482
R294 VPB.n61 VPB.n57 9.329
R295 VPB.n66 VPB.n65 8.97
R296 VPB.n183 VPB.n182 7.5
R297 VPB.n168 VPB.n167 7.5
R298 VPB.n173 VPB.n172 7.5
R299 VPB.n177 VPB.n176 7.5
R300 VPB.n165 VPB.n164 7.5
R301 VPB.n180 VPB.n166 7.5
R302 VPB.n225 VPB.n224 7.5
R303 VPB.n238 VPB.n237 7.5
R304 VPB.n232 VPB.n231 7.5
R305 VPB.n234 VPB.n233 7.5
R306 VPB.n227 VPB.n226 7.5
R307 VPB.n243 VPB.n242 7.5
R308 VPB.n107 VPB.n106 7.5
R309 VPB.n120 VPB.n119 7.5
R310 VPB.n114 VPB.n113 7.5
R311 VPB.n116 VPB.n115 7.5
R312 VPB.n109 VPB.n108 7.5
R313 VPB.n125 VPB.n124 7.5
R314 VPB.n85 VPB.n84 7.5
R315 VPB.n98 VPB.n97 7.5
R316 VPB.n92 VPB.n91 7.5
R317 VPB.n94 VPB.n93 7.5
R318 VPB.n87 VPB.n86 7.5
R319 VPB.n103 VPB.n102 7.5
R320 VPB.n333 VPB.n332 7.5
R321 VPB.n346 VPB.n345 7.5
R322 VPB.n340 VPB.n339 7.5
R323 VPB.n342 VPB.n341 7.5
R324 VPB.n335 VPB.n334 7.5
R325 VPB.n351 VPB.n350 7.5
R326 VPB.n18 VPB.n17 7.5
R327 VPB.n31 VPB.n30 7.5
R328 VPB.n25 VPB.n24 7.5
R329 VPB.n27 VPB.n26 7.5
R330 VPB.n20 VPB.n19 7.5
R331 VPB.n36 VPB.n35 7.5
R332 VPB.n409 VPB.n408 7.5
R333 VPB.n12 VPB.n11 7.5
R334 VPB.n6 VPB.n5 7.5
R335 VPB.n8 VPB.n7 7.5
R336 VPB.n2 VPB.n1 7.5
R337 VPB.n411 VPB.n410 7.5
R338 VPB.n37 VPB.n36 7.176
R339 VPB.n352 VPB.n351 7.176
R340 VPB.n162 VPB.n103 7.176
R341 VPB.n129 VPB.n125 7.176
R342 VPB.n244 VPB.n243 7.176
R343 VPB.n150 VPB.n146 6.817
R344 VPB.n239 VPB.n236 6.729
R345 VPB.n235 VPB.n232 6.729
R346 VPB.n230 VPB.n227 6.729
R347 VPB.n121 VPB.n118 6.729
R348 VPB.n117 VPB.n114 6.729
R349 VPB.n112 VPB.n109 6.729
R350 VPB.n99 VPB.n96 6.729
R351 VPB.n95 VPB.n92 6.729
R352 VPB.n90 VPB.n87 6.729
R353 VPB.n347 VPB.n344 6.729
R354 VPB.n343 VPB.n340 6.729
R355 VPB.n338 VPB.n335 6.729
R356 VPB.n32 VPB.n29 6.729
R357 VPB.n28 VPB.n25 6.729
R358 VPB.n23 VPB.n20 6.729
R359 VPB.n13 VPB.n10 6.729
R360 VPB.n9 VPB.n6 6.729
R361 VPB.n4 VPB.n2 6.729
R362 VPB.n230 VPB.n229 6.728
R363 VPB.n235 VPB.n234 6.728
R364 VPB.n239 VPB.n238 6.728
R365 VPB.n242 VPB.n241 6.728
R366 VPB.n112 VPB.n111 6.728
R367 VPB.n117 VPB.n116 6.728
R368 VPB.n121 VPB.n120 6.728
R369 VPB.n124 VPB.n123 6.728
R370 VPB.n90 VPB.n89 6.728
R371 VPB.n95 VPB.n94 6.728
R372 VPB.n99 VPB.n98 6.728
R373 VPB.n102 VPB.n101 6.728
R374 VPB.n338 VPB.n337 6.728
R375 VPB.n343 VPB.n342 6.728
R376 VPB.n347 VPB.n346 6.728
R377 VPB.n350 VPB.n349 6.728
R378 VPB.n23 VPB.n22 6.728
R379 VPB.n28 VPB.n27 6.728
R380 VPB.n32 VPB.n31 6.728
R381 VPB.n35 VPB.n34 6.728
R382 VPB.n4 VPB.n3 6.728
R383 VPB.n9 VPB.n8 6.728
R384 VPB.n13 VPB.n12 6.728
R385 VPB.n412 VPB.n411 6.728
R386 VPB.n192 VPB.n188 6.458
R387 VPB.n265 VPB.n261 6.458
R388 VPB.n146 VPB.n145 6.458
R389 VPB.n310 VPB.n306 6.458
R390 VPB.n373 VPB.n369 6.458
R391 VPB.n182 VPB.n181 6.398
R392 VPB.n201 VPB.n186 6.112
R393 VPB.n201 VPB.n200 6.101
R394 VPB.n70 VPB.n66 4.305
R395 VPB.n57 VPB.n56 3.947
R396 VPB.n217 VPB.n214 1.794
R397 VPB.n280 VPB.n277 1.794
R398 VPB.n158 VPB.n155 1.794
R399 VPB.n325 VPB.n322 1.794
R400 VPB.n388 VPB.n385 1.794
R401 VPB.n200 VPB.n197 1.435
R402 VPB.n253 VPB.n250 1.435
R403 VPB.n137 VPB.n136 1.435
R404 VPB.n299 VPB.n298 1.435
R405 VPB.n361 VPB.n358 1.435
R406 VPB.n180 VPB.n171 1.402
R407 VPB.n180 VPB.n174 1.402
R408 VPB.n180 VPB.n178 1.402
R409 VPB.n180 VPB.n179 1.402
R410 VPB.n48 VPB.n45 1.076
R411 VPB.n181 VPB.n180 0.735
R412 VPB.n180 VPB.n170 0.735
R413 VPB.n78 VPB.n77 0.717
R414 VPB.n240 VPB.n239 0.387
R415 VPB.n240 VPB.n235 0.387
R416 VPB.n240 VPB.n230 0.387
R417 VPB.n241 VPB.n240 0.387
R418 VPB.n122 VPB.n121 0.387
R419 VPB.n122 VPB.n117 0.387
R420 VPB.n122 VPB.n112 0.387
R421 VPB.n123 VPB.n122 0.387
R422 VPB.n100 VPB.n99 0.387
R423 VPB.n100 VPB.n95 0.387
R424 VPB.n100 VPB.n90 0.387
R425 VPB.n101 VPB.n100 0.387
R426 VPB.n348 VPB.n347 0.387
R427 VPB.n348 VPB.n343 0.387
R428 VPB.n348 VPB.n338 0.387
R429 VPB.n349 VPB.n348 0.387
R430 VPB.n33 VPB.n32 0.387
R431 VPB.n33 VPB.n28 0.387
R432 VPB.n33 VPB.n23 0.387
R433 VPB.n34 VPB.n33 0.387
R434 VPB.n413 VPB.n13 0.387
R435 VPB.n413 VPB.n9 0.387
R436 VPB.n413 VPB.n4 0.387
R437 VPB.n413 VPB.n412 0.387
R438 VPB.n249 VPB.n222 0.268
R439 VPB.n283 VPB.n282 0.268
R440 VPB.n291 VPB.n290 0.268
R441 VPB.n357 VPB.n330 0.268
R442 VPB.n394 VPB.n393 0.268
R443 VPB.n405 VPB 0.195
R444 VPB.n203 VPB.n202 0.134
R445 VPB.n208 VPB.n203 0.134
R446 VPB.n213 VPB.n208 0.134
R447 VPB.n218 VPB.n213 0.134
R448 VPB.n222 VPB.n218 0.134
R449 VPB.n254 VPB.n249 0.134
R450 VPB.n259 VPB.n254 0.134
R451 VPB.n266 VPB.n259 0.134
R452 VPB.n271 VPB.n266 0.134
R453 VPB.n276 VPB.n271 0.134
R454 VPB.n281 VPB.n276 0.134
R455 VPB.n282 VPB.n281 0.134
R456 VPB.n284 VPB.n283 0.134
R457 VPB.n285 VPB.n284 0.134
R458 VPB.n286 VPB.n285 0.134
R459 VPB.n287 VPB.n286 0.134
R460 VPB.n288 VPB.n287 0.134
R461 VPB.n289 VPB.n288 0.134
R462 VPB.n290 VPB.n289 0.134
R463 VPB.n291 VPB.n82 0.134
R464 VPB.n304 VPB.n82 0.134
R465 VPB.n311 VPB.n304 0.134
R466 VPB.n316 VPB.n311 0.134
R467 VPB.n321 VPB.n316 0.134
R468 VPB.n326 VPB.n321 0.134
R469 VPB.n330 VPB.n326 0.134
R470 VPB.n362 VPB.n357 0.134
R471 VPB.n367 VPB.n362 0.134
R472 VPB.n374 VPB.n367 0.134
R473 VPB.n379 VPB.n374 0.134
R474 VPB.n384 VPB.n379 0.134
R475 VPB.n389 VPB.n384 0.134
R476 VPB.n393 VPB.n389 0.134
R477 VPB.n395 VPB.n394 0.134
R478 VPB.n396 VPB.n395 0.134
R479 VPB.n397 VPB.n396 0.134
R480 VPB.n398 VPB.n397 0.134
R481 VPB.n399 VPB.n398 0.134
R482 VPB.n400 VPB.n399 0.134
R483 VPB.n401 VPB.n400 0.134
R484 VPB.n402 VPB.n401 0.134
R485 VPB.n403 VPB.n402 0.134
R486 VPB.n404 VPB.n403 0.134
R487 VPB.n405 VPB.n404 0.134
R488 a_277_1004.n8 a_277_1004.t8 480.392
R489 a_277_1004.n6 a_277_1004.t11 480.392
R490 a_277_1004.n8 a_277_1004.t12 403.272
R491 a_277_1004.n6 a_277_1004.t7 403.272
R492 a_277_1004.n9 a_277_1004.t9 293.527
R493 a_277_1004.n7 a_277_1004.t10 293.527
R494 a_277_1004.n13 a_277_1004.n11 223.151
R495 a_277_1004.n11 a_277_1004.n5 154.293
R496 a_277_1004.n10 a_277_1004.n7 83.3
R497 a_277_1004.n9 a_277_1004.n8 81.941
R498 a_277_1004.n7 a_277_1004.n6 81.941
R499 a_277_1004.n4 a_277_1004.n3 79.232
R500 a_277_1004.n11 a_277_1004.n10 77.315
R501 a_277_1004.n10 a_277_1004.n9 76
R502 a_277_1004.n5 a_277_1004.n4 63.152
R503 a_277_1004.n13 a_277_1004.n12 30
R504 a_277_1004.n14 a_277_1004.n0 24.383
R505 a_277_1004.n14 a_277_1004.n13 23.684
R506 a_277_1004.n5 a_277_1004.n1 16.08
R507 a_277_1004.n4 a_277_1004.n2 16.08
R508 a_277_1004.n1 a_277_1004.t0 14.282
R509 a_277_1004.n1 a_277_1004.t1 14.282
R510 a_277_1004.n2 a_277_1004.t4 14.282
R511 a_277_1004.n2 a_277_1004.t3 14.282
R512 a_277_1004.n3 a_277_1004.t6 14.282
R513 a_277_1004.n3 a_277_1004.t5 14.282
R514 a_91_75.t0 a_91_75.n0 117.777
R515 a_91_75.n2 a_91_75.n1 55.228
R516 a_91_75.n4 a_91_75.n3 9.111
R517 a_91_75.n8 a_91_75.n6 7.859
R518 a_91_75.t0 a_91_75.n2 4.04
R519 a_91_75.t0 a_91_75.n8 3.034
R520 a_91_75.n6 a_91_75.n4 1.964
R521 a_91_75.n6 a_91_75.n5 1.964
R522 a_91_75.n8 a_91_75.n7 0.443
R523 a_372_182.n8 a_372_182.n6 96.467
R524 a_372_182.n3 a_372_182.n1 44.628
R525 a_372_182.t0 a_372_182.n8 32.417
R526 a_372_182.n3 a_372_182.n2 23.284
R527 a_372_182.n6 a_372_182.n5 22.349
R528 a_372_182.t0 a_372_182.n10 20.241
R529 a_372_182.n10 a_372_182.n9 13.494
R530 a_372_182.n6 a_372_182.n4 8.443
R531 a_372_182.t0 a_372_182.n0 8.137
R532 a_372_182.t0 a_372_182.n3 5.727
R533 a_372_182.n8 a_372_182.n7 1.435
R534 a_599_943.n4 a_599_943.t7 480.392
R535 a_599_943.n6 a_599_943.t8 454.685
R536 a_599_943.n6 a_599_943.t6 428.979
R537 a_599_943.n4 a_599_943.t10 403.272
R538 a_599_943.n5 a_599_943.t5 266.974
R539 a_599_943.n7 a_599_943.t9 221.453
R540 a_599_943.n11 a_599_943.n9 194.086
R541 a_599_943.n9 a_599_943.n3 162.547
R542 a_599_943.n7 a_599_943.n6 108.494
R543 a_599_943.n5 a_599_943.n4 108.494
R544 a_599_943.n8 a_599_943.n7 78.947
R545 a_599_943.n8 a_599_943.n5 77.315
R546 a_599_943.n3 a_599_943.n2 76.002
R547 a_599_943.n9 a_599_943.n8 76
R548 a_599_943.n11 a_599_943.n10 30
R549 a_599_943.n12 a_599_943.n0 24.383
R550 a_599_943.n12 a_599_943.n11 23.684
R551 a_599_943.n1 a_599_943.t2 14.282
R552 a_599_943.n1 a_599_943.t1 14.282
R553 a_599_943.n2 a_599_943.t4 14.282
R554 a_599_943.n2 a_599_943.t3 14.282
R555 a_599_943.n3 a_599_943.n1 12.85
R556 a_1740_73.n10 a_1740_73.n9 93.333
R557 a_1740_73.n2 a_1740_73.n1 41.622
R558 a_1740_73.n13 a_1740_73.n12 26.667
R559 a_1740_73.n6 a_1740_73.n5 24.977
R560 a_1740_73.t0 a_1740_73.n2 21.209
R561 a_1740_73.t0 a_1740_73.n3 11.595
R562 a_1740_73.t1 a_1740_73.n8 8.137
R563 a_1740_73.t0 a_1740_73.n0 6.109
R564 a_1740_73.t1 a_1740_73.n7 4.864
R565 a_1740_73.t0 a_1740_73.n4 3.871
R566 a_1740_73.t0 a_1740_73.n13 2.535
R567 a_1740_73.n13 a_1740_73.t1 1.145
R568 a_1740_73.n7 a_1740_73.n6 1.13
R569 a_1740_73.t1 a_1740_73.n11 0.804
R570 a_1740_73.n11 a_1740_73.n10 0.136
R571 VNB VNB.n366 300.778
R572 VNB.n194 VNB.n193 199.897
R573 VNB.n88 VNB.n87 199.897
R574 VNB.n68 VNB.n67 199.897
R575 VNB.n292 VNB.n291 199.897
R576 VNB.n15 VNB.n14 199.897
R577 VNB.n100 VNB.n98 154.509
R578 VNB.n203 VNB.n201 154.509
R579 VNB.n301 VNB.n299 154.509
R580 VNB.n251 VNB.n249 154.509
R581 VNB.n24 VNB.n22 154.509
R582 VNB.n160 VNB.n159 121.366
R583 VNB.n219 VNB.n218 121.366
R584 VNB.n112 VNB.n111 121.366
R585 VNB.n317 VNB.n316 121.366
R586 VNB.n53 VNB.n4 85.559
R587 VNB.n269 VNB.n268 84.842
R588 VNB.n255 VNB.n57 76
R589 VNB.n353 VNB.n352 76
R590 VNB.n340 VNB.n339 76
R591 VNB.n336 VNB.n335 76
R592 VNB.n332 VNB.n331 76
R593 VNB.n321 VNB.n320 76
R594 VNB.n315 VNB.n314 76
R595 VNB.n311 VNB.n310 76
R596 VNB.n307 VNB.n306 76
R597 VNB.n303 VNB.n302 76
R598 VNB.n281 VNB.n280 76
R599 VNB.n277 VNB.n276 76
R600 VNB.n273 VNB.n272 76
R601 VNB.n267 VNB.n266 76
R602 VNB.n263 VNB.n262 76
R603 VNB.n259 VNB.n258 76
R604 VNB.n252 VNB.n248 76
R605 VNB.n238 VNB.n237 76
R606 VNB.n234 VNB.n233 76
R607 VNB.n223 VNB.n222 76
R608 VNB.n217 VNB.n216 76
R609 VNB.n213 VNB.n212 76
R610 VNB.n209 VNB.n208 76
R611 VNB.n205 VNB.n204 76
R612 VNB.n183 VNB.n182 76
R613 VNB.n179 VNB.n178 76
R614 VNB.n175 VNB.n174 76
R615 VNB.n164 VNB.n163 76
R616 VNB.n169 VNB.n168 63.835
R617 VNB.n228 VNB.n227 63.835
R618 VNB.n116 VNB.n77 63.835
R619 VNB.n326 VNB.n325 63.835
R620 VNB.n51 VNB.n50 41.971
R621 VNB.n161 VNB.n160 36.937
R622 VNB.n220 VNB.n219 36.937
R623 VNB.n113 VNB.n112 36.937
R624 VNB.n318 VNB.n317 36.937
R625 VNB.n271 VNB.n270 36.678
R626 VNB.n157 VNB.n156 35.118
R627 VNB.n168 VNB.n167 28.421
R628 VNB.n227 VNB.n226 28.421
R629 VNB.n77 VNB.n76 28.421
R630 VNB.n325 VNB.n324 28.421
R631 VNB.n172 VNB.n171 27.855
R632 VNB.n231 VNB.n230 27.855
R633 VNB.n119 VNB.n118 27.855
R634 VNB.n329 VNB.n328 27.855
R635 VNB.n168 VNB.n166 25.263
R636 VNB.n227 VNB.n225 25.263
R637 VNB.n77 VNB.n75 25.263
R638 VNB.n325 VNB.n323 25.263
R639 VNB.n166 VNB.n165 24.383
R640 VNB.n225 VNB.n224 24.383
R641 VNB.n75 VNB.n74 24.383
R642 VNB.n323 VNB.n322 24.383
R643 VNB.n146 VNB.n143 20.452
R644 VNB.n354 VNB.n353 20.452
R645 VNB.n173 VNB.n172 16.721
R646 VNB.n232 VNB.n231 16.721
R647 VNB.n120 VNB.n119 16.721
R648 VNB.n330 VNB.n329 16.721
R649 VNB.n155 VNB.n154 13.653
R650 VNB.n154 VNB.n153 13.653
R651 VNB.n152 VNB.n151 13.653
R652 VNB.n151 VNB.n150 13.653
R653 VNB.n149 VNB.n148 13.653
R654 VNB.n148 VNB.n147 13.653
R655 VNB.n163 VNB.n162 13.653
R656 VNB.n162 VNB.n161 13.653
R657 VNB.n174 VNB.n173 13.653
R658 VNB.n178 VNB.n177 13.653
R659 VNB.n177 VNB.n176 13.653
R660 VNB.n182 VNB.n181 13.653
R661 VNB.n181 VNB.n180 13.653
R662 VNB.n204 VNB.n203 13.653
R663 VNB.n203 VNB.n202 13.653
R664 VNB.n208 VNB.n207 13.653
R665 VNB.n207 VNB.n206 13.653
R666 VNB.n212 VNB.n211 13.653
R667 VNB.n211 VNB.n210 13.653
R668 VNB.n216 VNB.n215 13.653
R669 VNB.n215 VNB.n214 13.653
R670 VNB.n222 VNB.n221 13.653
R671 VNB.n221 VNB.n220 13.653
R672 VNB.n233 VNB.n232 13.653
R673 VNB.n237 VNB.n236 13.653
R674 VNB.n236 VNB.n235 13.653
R675 VNB.n96 VNB.n95 13.653
R676 VNB.n95 VNB.n94 13.653
R677 VNB.n101 VNB.n100 13.653
R678 VNB.n100 VNB.n99 13.653
R679 VNB.n104 VNB.n103 13.653
R680 VNB.n103 VNB.n102 13.653
R681 VNB.n107 VNB.n106 13.653
R682 VNB.n106 VNB.n105 13.653
R683 VNB.n110 VNB.n109 13.653
R684 VNB.n109 VNB.n108 13.653
R685 VNB.n115 VNB.n114 13.653
R686 VNB.n114 VNB.n113 13.653
R687 VNB.n121 VNB.n120 13.653
R688 VNB.n124 VNB.n123 13.653
R689 VNB.n123 VNB.n122 13.653
R690 VNB.n127 VNB.n126 13.653
R691 VNB.n126 VNB.n125 13.653
R692 VNB.n252 VNB.n251 13.653
R693 VNB.n251 VNB.n250 13.653
R694 VNB.n255 VNB.n254 13.653
R695 VNB.n254 VNB.n253 13.653
R696 VNB.n258 VNB.n257 13.653
R697 VNB.n257 VNB.n256 13.653
R698 VNB.n262 VNB.n261 13.653
R699 VNB.n261 VNB.n260 13.653
R700 VNB.n266 VNB.n265 13.653
R701 VNB.n265 VNB.n264 13.653
R702 VNB.n272 VNB.n271 13.653
R703 VNB.n276 VNB.n275 13.653
R704 VNB.n275 VNB.n274 13.653
R705 VNB.n280 VNB.n279 13.653
R706 VNB.n279 VNB.n278 13.653
R707 VNB.n302 VNB.n301 13.653
R708 VNB.n301 VNB.n300 13.653
R709 VNB.n306 VNB.n305 13.653
R710 VNB.n305 VNB.n304 13.653
R711 VNB.n310 VNB.n309 13.653
R712 VNB.n309 VNB.n308 13.653
R713 VNB.n314 VNB.n313 13.653
R714 VNB.n313 VNB.n312 13.653
R715 VNB.n320 VNB.n319 13.653
R716 VNB.n319 VNB.n318 13.653
R717 VNB.n331 VNB.n330 13.653
R718 VNB.n335 VNB.n334 13.653
R719 VNB.n334 VNB.n333 13.653
R720 VNB.n339 VNB.n338 13.653
R721 VNB.n338 VNB.n337 13.653
R722 VNB.n25 VNB.n24 13.653
R723 VNB.n24 VNB.n23 13.653
R724 VNB.n28 VNB.n27 13.653
R725 VNB.n27 VNB.n26 13.653
R726 VNB.n31 VNB.n30 13.653
R727 VNB.n30 VNB.n29 13.653
R728 VNB.n34 VNB.n33 13.653
R729 VNB.n33 VNB.n32 13.653
R730 VNB.n37 VNB.n36 13.653
R731 VNB.n36 VNB.n35 13.653
R732 VNB.n40 VNB.n39 13.653
R733 VNB.n39 VNB.n38 13.653
R734 VNB.n43 VNB.n42 13.653
R735 VNB.n42 VNB.n41 13.653
R736 VNB.n46 VNB.n45 13.653
R737 VNB.n45 VNB.n44 13.653
R738 VNB.n49 VNB.n48 13.653
R739 VNB.n48 VNB.n47 13.653
R740 VNB.n52 VNB.n51 13.653
R741 VNB.n56 VNB.n55 13.653
R742 VNB.n55 VNB.n54 13.653
R743 VNB.n353 VNB.n0 13.653
R744 VNB VNB.n0 13.653
R745 VNB.n146 VNB.n145 13.653
R746 VNB.n145 VNB.n144 13.653
R747 VNB.n361 VNB.n358 13.577
R748 VNB.n131 VNB.n129 13.276
R749 VNB.n143 VNB.n131 13.276
R750 VNB.n186 VNB.n184 13.276
R751 VNB.n199 VNB.n186 13.276
R752 VNB.n80 VNB.n78 13.276
R753 VNB.n93 VNB.n80 13.276
R754 VNB.n60 VNB.n58 13.276
R755 VNB.n73 VNB.n60 13.276
R756 VNB.n284 VNB.n282 13.276
R757 VNB.n297 VNB.n284 13.276
R758 VNB.n7 VNB.n5 13.276
R759 VNB.n20 VNB.n7 13.276
R760 VNB.n155 VNB.n152 13.276
R761 VNB.n152 VNB.n149 13.276
R762 VNB.n204 VNB.n200 13.276
R763 VNB.n97 VNB.n96 13.276
R764 VNB.n101 VNB.n97 13.276
R765 VNB.n104 VNB.n101 13.276
R766 VNB.n107 VNB.n104 13.276
R767 VNB.n110 VNB.n107 13.276
R768 VNB.n115 VNB.n110 13.276
R769 VNB.n124 VNB.n121 13.276
R770 VNB.n127 VNB.n124 13.276
R771 VNB.n128 VNB.n127 13.276
R772 VNB.n252 VNB.n128 13.276
R773 VNB.n255 VNB.n252 13.276
R774 VNB.n258 VNB.n255 13.276
R775 VNB.n302 VNB.n298 13.276
R776 VNB.n25 VNB.n21 13.276
R777 VNB.n28 VNB.n25 13.276
R778 VNB.n31 VNB.n28 13.276
R779 VNB.n34 VNB.n31 13.276
R780 VNB.n37 VNB.n34 13.276
R781 VNB.n40 VNB.n37 13.276
R782 VNB.n43 VNB.n40 13.276
R783 VNB.n46 VNB.n43 13.276
R784 VNB.n49 VNB.n46 13.276
R785 VNB.n52 VNB.n49 13.276
R786 VNB.n353 VNB.n56 13.276
R787 VNB.n3 VNB.n1 13.276
R788 VNB.n354 VNB.n3 13.276
R789 VNB.n56 VNB.n53 12.02
R790 VNB.n116 VNB.n115 10.764
R791 VNB.n363 VNB.n362 7.5
R792 VNB.n192 VNB.n191 7.5
R793 VNB.n188 VNB.n187 7.5
R794 VNB.n186 VNB.n185 7.5
R795 VNB.n199 VNB.n198 7.5
R796 VNB.n86 VNB.n85 7.5
R797 VNB.n82 VNB.n81 7.5
R798 VNB.n80 VNB.n79 7.5
R799 VNB.n93 VNB.n92 7.5
R800 VNB.n66 VNB.n65 7.5
R801 VNB.n62 VNB.n61 7.5
R802 VNB.n60 VNB.n59 7.5
R803 VNB.n73 VNB.n72 7.5
R804 VNB.n290 VNB.n289 7.5
R805 VNB.n286 VNB.n285 7.5
R806 VNB.n284 VNB.n283 7.5
R807 VNB.n297 VNB.n296 7.5
R808 VNB.n13 VNB.n12 7.5
R809 VNB.n9 VNB.n8 7.5
R810 VNB.n7 VNB.n6 7.5
R811 VNB.n20 VNB.n19 7.5
R812 VNB.n355 VNB.n354 7.5
R813 VNB.n3 VNB.n2 7.5
R814 VNB.n360 VNB.n359 7.5
R815 VNB.n137 VNB.n136 7.5
R816 VNB.n133 VNB.n132 7.5
R817 VNB.n131 VNB.n130 7.5
R818 VNB.n143 VNB.n142 7.5
R819 VNB.n200 VNB.n199 7.176
R820 VNB.n97 VNB.n93 7.176
R821 VNB.n128 VNB.n73 7.176
R822 VNB.n298 VNB.n297 7.176
R823 VNB.n21 VNB.n20 7.176
R824 VNB.n365 VNB.n363 7.011
R825 VNB.n195 VNB.n192 7.011
R826 VNB.n190 VNB.n188 7.011
R827 VNB.n89 VNB.n86 7.011
R828 VNB.n84 VNB.n82 7.011
R829 VNB.n69 VNB.n66 7.011
R830 VNB.n64 VNB.n62 7.011
R831 VNB.n293 VNB.n290 7.011
R832 VNB.n288 VNB.n286 7.011
R833 VNB.n16 VNB.n13 7.011
R834 VNB.n11 VNB.n9 7.011
R835 VNB.n139 VNB.n137 7.011
R836 VNB.n135 VNB.n133 7.011
R837 VNB.n198 VNB.n197 7.01
R838 VNB.n190 VNB.n189 7.01
R839 VNB.n195 VNB.n194 7.01
R840 VNB.n92 VNB.n91 7.01
R841 VNB.n84 VNB.n83 7.01
R842 VNB.n89 VNB.n88 7.01
R843 VNB.n72 VNB.n71 7.01
R844 VNB.n64 VNB.n63 7.01
R845 VNB.n69 VNB.n68 7.01
R846 VNB.n296 VNB.n295 7.01
R847 VNB.n288 VNB.n287 7.01
R848 VNB.n293 VNB.n292 7.01
R849 VNB.n19 VNB.n18 7.01
R850 VNB.n11 VNB.n10 7.01
R851 VNB.n16 VNB.n15 7.01
R852 VNB.n142 VNB.n141 7.01
R853 VNB.n135 VNB.n134 7.01
R854 VNB.n139 VNB.n138 7.01
R855 VNB.n365 VNB.n364 7.01
R856 VNB.n361 VNB.n360 6.788
R857 VNB.n356 VNB.n355 6.788
R858 VNB.n156 VNB.n146 6.111
R859 VNB.n156 VNB.n155 6.1
R860 VNB.n174 VNB.n169 2.511
R861 VNB.n233 VNB.n228 2.511
R862 VNB.n121 VNB.n116 2.511
R863 VNB.n272 VNB.n269 2.511
R864 VNB.n331 VNB.n326 2.511
R865 VNB.n172 VNB.n170 1.99
R866 VNB.n231 VNB.n229 1.99
R867 VNB.n119 VNB.n117 1.99
R868 VNB.n329 VNB.n327 1.99
R869 VNB.n53 VNB.n52 1.255
R870 VNB.n366 VNB.n357 0.921
R871 VNB.n366 VNB.n361 0.476
R872 VNB.n366 VNB.n356 0.475
R873 VNB.n205 VNB.n183 0.272
R874 VNB.n240 VNB.n239 0.272
R875 VNB.n248 VNB.n247 0.272
R876 VNB.n303 VNB.n281 0.272
R877 VNB.n341 VNB.n340 0.272
R878 VNB.n196 VNB.n190 0.246
R879 VNB.n197 VNB.n196 0.246
R880 VNB.n196 VNB.n195 0.246
R881 VNB.n90 VNB.n84 0.246
R882 VNB.n91 VNB.n90 0.246
R883 VNB.n90 VNB.n89 0.246
R884 VNB.n70 VNB.n64 0.246
R885 VNB.n71 VNB.n70 0.246
R886 VNB.n70 VNB.n69 0.246
R887 VNB.n294 VNB.n288 0.246
R888 VNB.n295 VNB.n294 0.246
R889 VNB.n294 VNB.n293 0.246
R890 VNB.n17 VNB.n11 0.246
R891 VNB.n18 VNB.n17 0.246
R892 VNB.n17 VNB.n16 0.246
R893 VNB.n140 VNB.n135 0.246
R894 VNB.n141 VNB.n140 0.246
R895 VNB.n140 VNB.n139 0.246
R896 VNB.n366 VNB.n365 0.246
R897 VNB.n352 VNB 0.198
R898 VNB.n158 VNB.n157 0.136
R899 VNB.n164 VNB.n158 0.136
R900 VNB.n175 VNB.n164 0.136
R901 VNB.n179 VNB.n175 0.136
R902 VNB.n183 VNB.n179 0.136
R903 VNB.n209 VNB.n205 0.136
R904 VNB.n213 VNB.n209 0.136
R905 VNB.n217 VNB.n213 0.136
R906 VNB.n223 VNB.n217 0.136
R907 VNB.n234 VNB.n223 0.136
R908 VNB.n238 VNB.n234 0.136
R909 VNB.n239 VNB.n238 0.136
R910 VNB.n241 VNB.n240 0.136
R911 VNB.n242 VNB.n241 0.136
R912 VNB.n243 VNB.n242 0.136
R913 VNB.n244 VNB.n243 0.136
R914 VNB.n245 VNB.n244 0.136
R915 VNB.n246 VNB.n245 0.136
R916 VNB.n247 VNB.n246 0.136
R917 VNB.n248 VNB.n57 0.136
R918 VNB.n259 VNB.n57 0.136
R919 VNB.n263 VNB.n259 0.136
R920 VNB.n267 VNB.n263 0.136
R921 VNB.n273 VNB.n267 0.136
R922 VNB.n277 VNB.n273 0.136
R923 VNB.n281 VNB.n277 0.136
R924 VNB.n307 VNB.n303 0.136
R925 VNB.n311 VNB.n307 0.136
R926 VNB.n315 VNB.n311 0.136
R927 VNB.n321 VNB.n315 0.136
R928 VNB.n332 VNB.n321 0.136
R929 VNB.n336 VNB.n332 0.136
R930 VNB.n340 VNB.n336 0.136
R931 VNB.n342 VNB.n341 0.136
R932 VNB.n343 VNB.n342 0.136
R933 VNB.n344 VNB.n343 0.136
R934 VNB.n345 VNB.n344 0.136
R935 VNB.n346 VNB.n345 0.136
R936 VNB.n347 VNB.n346 0.136
R937 VNB.n348 VNB.n347 0.136
R938 VNB.n349 VNB.n348 0.136
R939 VNB.n350 VNB.n349 0.136
R940 VNB.n351 VNB.n350 0.136
R941 VNB.n352 VNB.n351 0.136
R942 a_2406_73.n12 a_2406_73.n11 26.811
R943 a_2406_73.n6 a_2406_73.n5 24.977
R944 a_2406_73.n2 a_2406_73.n1 24.877
R945 a_2406_73.t0 a_2406_73.n2 12.677
R946 a_2406_73.t0 a_2406_73.n3 11.595
R947 a_2406_73.t1 a_2406_73.n8 8.137
R948 a_2406_73.t0 a_2406_73.n4 7.273
R949 a_2406_73.t0 a_2406_73.n0 6.109
R950 a_2406_73.t1 a_2406_73.n7 4.864
R951 a_2406_73.t0 a_2406_73.n12 2.074
R952 a_2406_73.n7 a_2406_73.n6 1.13
R953 a_2406_73.n12 a_2406_73.t1 0.937
R954 a_2406_73.t1 a_2406_73.n10 0.804
R955 a_2406_73.n10 a_2406_73.n9 0.136
R956 a_3738_73.n12 a_3738_73.n11 26.811
R957 a_3738_73.n6 a_3738_73.n5 24.977
R958 a_3738_73.n2 a_3738_73.n1 24.877
R959 a_3738_73.t0 a_3738_73.n2 12.677
R960 a_3738_73.t0 a_3738_73.n3 11.595
R961 a_3738_73.t1 a_3738_73.n8 8.137
R962 a_3738_73.t0 a_3738_73.n4 7.273
R963 a_3738_73.t0 a_3738_73.n0 6.109
R964 a_3738_73.t1 a_3738_73.n7 4.864
R965 a_3738_73.t0 a_3738_73.n12 2.074
R966 a_3738_73.n7 a_3738_73.n6 1.13
R967 a_3738_73.n12 a_3738_73.t1 0.937
R968 a_3738_73.t1 a_3738_73.n10 0.804
R969 a_3738_73.n10 a_3738_73.n9 0.136
R970 a_1074_73.t0 a_1074_73.n1 34.62
R971 a_1074_73.t0 a_1074_73.n0 8.137
R972 a_1074_73.t0 a_1074_73.n2 4.69
R973 a_3072_73.n12 a_3072_73.n11 26.811
R974 a_3072_73.n6 a_3072_73.n5 24.977
R975 a_3072_73.n2 a_3072_73.n1 24.877
R976 a_3072_73.t0 a_3072_73.n2 12.677
R977 a_3072_73.t0 a_3072_73.n3 11.595
R978 a_3072_73.t1 a_3072_73.n8 8.137
R979 a_3072_73.t0 a_3072_73.n4 7.273
R980 a_3072_73.t0 a_3072_73.n0 6.109
R981 a_3072_73.t1 a_3072_73.n7 4.864
R982 a_3072_73.t0 a_3072_73.n12 2.074
R983 a_3072_73.n7 a_3072_73.n6 1.13
R984 a_3072_73.n12 a_3072_73.t1 0.937
R985 a_3072_73.t1 a_3072_73.n10 0.804
R986 a_3072_73.n10 a_3072_73.n9 0.136








































































































































































































































































































































































































































































































































.ends
