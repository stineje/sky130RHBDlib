magic
tech sky130A
magscale 1 2
timestamp 1669564320
<< nwell >>
rect -87 786 18069 1550
<< pwell >>
rect -34 -34 18016 544
<< nmos >>
rect 147 290 177 351
tri 177 290 193 306 sw
rect 447 290 477 351
rect 147 260 253 290
tri 253 260 283 290 sw
rect 147 159 177 260
tri 177 244 193 260 nw
tri 237 244 253 260 ne
tri 177 159 193 175 sw
tri 237 159 253 175 se
rect 253 159 283 260
tri 342 260 372 290 se
rect 372 260 477 290
rect 342 166 372 260
tri 372 244 388 260 nw
tri 431 244 447 260 ne
tri 372 166 388 182 sw
tri 431 166 447 182 se
rect 447 166 477 260
tri 147 129 177 159 ne
rect 177 129 253 159
tri 253 129 283 159 nw
tri 342 136 372 166 ne
rect 372 136 447 166
tri 447 136 477 166 nw
rect 649 298 679 351
tri 679 298 695 314 sw
rect 649 268 755 298
tri 755 268 785 298 sw
rect 649 167 679 268
tri 679 252 695 268 nw
tri 739 252 755 268 ne
tri 679 167 695 183 sw
tri 739 167 755 183 se
rect 755 167 785 268
tri 649 137 679 167 ne
rect 679 137 755 167
tri 755 137 785 167 nw
rect 1109 290 1139 351
tri 1139 290 1155 306 sw
rect 1409 290 1439 351
rect 1109 260 1215 290
tri 1215 260 1245 290 sw
rect 1109 159 1139 260
tri 1139 244 1155 260 nw
tri 1199 244 1215 260 ne
tri 1139 159 1155 175 sw
tri 1199 159 1215 175 se
rect 1215 159 1245 260
tri 1304 260 1334 290 se
rect 1334 260 1439 290
rect 1304 166 1334 260
tri 1334 244 1350 260 nw
tri 1393 244 1409 260 ne
tri 1334 166 1350 182 sw
tri 1393 166 1409 182 se
rect 1409 166 1439 260
tri 1109 129 1139 159 ne
rect 1139 129 1215 159
tri 1215 129 1245 159 nw
tri 1304 136 1334 166 ne
rect 1334 136 1409 166
tri 1409 136 1439 166 nw
rect 1611 298 1641 351
tri 1641 298 1657 314 sw
rect 1611 268 1717 298
tri 1717 268 1747 298 sw
rect 1611 167 1641 268
tri 1641 252 1657 268 nw
tri 1701 252 1717 268 ne
tri 1641 167 1657 183 sw
tri 1701 167 1717 183 se
rect 1717 167 1747 268
tri 1611 137 1641 167 ne
rect 1641 137 1717 167
tri 1717 137 1747 167 nw
rect 2092 288 2122 349
tri 2122 288 2138 304 sw
rect 2286 296 2316 349
tri 2316 296 2332 312 sw
rect 2092 258 2198 288
tri 2198 258 2228 288 sw
rect 2286 266 2392 296
tri 2392 266 2422 296 sw
rect 2092 157 2122 258
tri 2122 242 2138 258 nw
tri 2182 242 2198 258 ne
tri 2122 157 2138 173 sw
tri 2182 157 2198 173 se
rect 2198 157 2228 258
rect 2286 165 2316 266
tri 2316 250 2332 266 nw
tri 2376 250 2392 266 ne
tri 2316 165 2332 181 sw
tri 2376 165 2392 181 se
rect 2392 165 2422 266
tri 2092 127 2122 157 ne
rect 2122 127 2198 157
tri 2198 127 2228 157 nw
tri 2286 135 2316 165 ne
rect 2316 135 2392 165
tri 2392 135 2422 165 nw
rect 2737 290 2767 351
tri 2767 290 2783 306 sw
rect 3037 290 3067 351
rect 2737 260 2843 290
tri 2843 260 2873 290 sw
rect 2737 159 2767 260
tri 2767 244 2783 260 nw
tri 2827 244 2843 260 ne
tri 2767 159 2783 175 sw
tri 2827 159 2843 175 se
rect 2843 159 2873 260
tri 2932 260 2962 290 se
rect 2962 260 3067 290
rect 2932 166 2962 260
tri 2962 244 2978 260 nw
tri 3021 244 3037 260 ne
tri 2962 166 2978 182 sw
tri 3021 166 3037 182 se
rect 3037 166 3067 260
tri 2737 129 2767 159 ne
rect 2767 129 2843 159
tri 2843 129 2873 159 nw
tri 2932 136 2962 166 ne
rect 2962 136 3037 166
tri 3037 136 3067 166 nw
rect 3239 298 3269 351
tri 3269 298 3285 314 sw
rect 3239 268 3345 298
tri 3345 268 3375 298 sw
rect 3239 167 3269 268
tri 3269 252 3285 268 nw
tri 3329 252 3345 268 ne
tri 3269 167 3285 183 sw
tri 3329 167 3345 183 se
rect 3345 167 3375 268
tri 3239 137 3269 167 ne
rect 3269 137 3345 167
tri 3345 137 3375 167 nw
rect 3699 290 3729 351
tri 3729 290 3745 306 sw
rect 3999 290 4029 351
rect 3699 260 3805 290
tri 3805 260 3835 290 sw
rect 3699 159 3729 260
tri 3729 244 3745 260 nw
tri 3789 244 3805 260 ne
tri 3729 159 3745 175 sw
tri 3789 159 3805 175 se
rect 3805 159 3835 260
tri 3894 260 3924 290 se
rect 3924 260 4029 290
rect 3894 166 3924 260
tri 3924 244 3940 260 nw
tri 3983 244 3999 260 ne
tri 3924 166 3940 182 sw
tri 3983 166 3999 182 se
rect 3999 166 4029 260
tri 3699 129 3729 159 ne
rect 3729 129 3805 159
tri 3805 129 3835 159 nw
tri 3894 136 3924 166 ne
rect 3924 136 3999 166
tri 3999 136 4029 166 nw
rect 4201 298 4231 351
tri 4231 298 4247 314 sw
rect 4201 268 4307 298
tri 4307 268 4337 298 sw
rect 4201 167 4231 268
tri 4231 252 4247 268 nw
tri 4291 252 4307 268 ne
tri 4231 167 4247 183 sw
tri 4291 167 4307 183 se
rect 4307 167 4337 268
tri 4201 137 4231 167 ne
rect 4231 137 4307 167
tri 4307 137 4337 167 nw
rect 4682 288 4712 349
tri 4712 288 4728 304 sw
rect 4876 296 4906 349
tri 4906 296 4922 312 sw
rect 4682 258 4788 288
tri 4788 258 4818 288 sw
rect 4876 266 4982 296
tri 4982 266 5012 296 sw
rect 4682 157 4712 258
tri 4712 242 4728 258 nw
tri 4772 242 4788 258 ne
tri 4712 157 4728 173 sw
tri 4772 157 4788 173 se
rect 4788 157 4818 258
rect 4876 165 4906 266
tri 4906 250 4922 266 nw
tri 4966 250 4982 266 ne
tri 4906 165 4922 181 sw
tri 4966 165 4982 181 se
rect 4982 165 5012 266
tri 4682 127 4712 157 ne
rect 4712 127 4788 157
tri 4788 127 4818 157 nw
tri 4876 135 4906 165 ne
rect 4906 135 4982 165
tri 4982 135 5012 165 nw
rect 5327 290 5357 351
tri 5357 290 5373 306 sw
rect 5627 290 5657 351
rect 5327 260 5433 290
tri 5433 260 5463 290 sw
rect 5327 159 5357 260
tri 5357 244 5373 260 nw
tri 5417 244 5433 260 ne
tri 5357 159 5373 175 sw
tri 5417 159 5433 175 se
rect 5433 159 5463 260
tri 5522 260 5552 290 se
rect 5552 260 5657 290
rect 5522 166 5552 260
tri 5552 244 5568 260 nw
tri 5611 244 5627 260 ne
tri 5552 166 5568 182 sw
tri 5611 166 5627 182 se
rect 5627 166 5657 260
tri 5327 129 5357 159 ne
rect 5357 129 5433 159
tri 5433 129 5463 159 nw
tri 5522 136 5552 166 ne
rect 5552 136 5627 166
tri 5627 136 5657 166 nw
rect 5829 298 5859 351
tri 5859 298 5875 314 sw
rect 5829 268 5935 298
tri 5935 268 5965 298 sw
rect 5829 167 5859 268
tri 5859 252 5875 268 nw
tri 5919 252 5935 268 ne
tri 5859 167 5875 183 sw
tri 5919 167 5935 183 se
rect 5935 167 5965 268
tri 5829 137 5859 167 ne
rect 5859 137 5935 167
tri 5935 137 5965 167 nw
rect 6289 290 6319 351
tri 6319 290 6335 306 sw
rect 6589 290 6619 351
rect 6289 260 6395 290
tri 6395 260 6425 290 sw
rect 6289 159 6319 260
tri 6319 244 6335 260 nw
tri 6379 244 6395 260 ne
tri 6319 159 6335 175 sw
tri 6379 159 6395 175 se
rect 6395 159 6425 260
tri 6484 260 6514 290 se
rect 6514 260 6619 290
rect 6484 166 6514 260
tri 6514 244 6530 260 nw
tri 6573 244 6589 260 ne
tri 6514 166 6530 182 sw
tri 6573 166 6589 182 se
rect 6589 166 6619 260
tri 6289 129 6319 159 ne
rect 6319 129 6395 159
tri 6395 129 6425 159 nw
tri 6484 136 6514 166 ne
rect 6514 136 6589 166
tri 6589 136 6619 166 nw
rect 6791 298 6821 351
tri 6821 298 6837 314 sw
rect 6791 268 6897 298
tri 6897 268 6927 298 sw
rect 6791 167 6821 268
tri 6821 252 6837 268 nw
tri 6881 252 6897 268 ne
tri 6821 167 6837 183 sw
tri 6881 167 6897 183 se
rect 6897 167 6927 268
tri 6791 137 6821 167 ne
rect 6821 137 6897 167
tri 6897 137 6927 167 nw
rect 7272 288 7302 349
tri 7302 288 7318 304 sw
rect 7466 296 7496 349
tri 7496 296 7512 312 sw
rect 7272 258 7378 288
tri 7378 258 7408 288 sw
rect 7466 266 7572 296
tri 7572 266 7602 296 sw
rect 7272 157 7302 258
tri 7302 242 7318 258 nw
tri 7362 242 7378 258 ne
tri 7302 157 7318 173 sw
tri 7362 157 7378 173 se
rect 7378 157 7408 258
rect 7466 165 7496 266
tri 7496 250 7512 266 nw
tri 7556 250 7572 266 ne
tri 7496 165 7512 181 sw
tri 7556 165 7572 181 se
rect 7572 165 7602 266
tri 7272 127 7302 157 ne
rect 7302 127 7378 157
tri 7378 127 7408 157 nw
tri 7466 135 7496 165 ne
rect 7496 135 7572 165
tri 7572 135 7602 165 nw
rect 7917 290 7947 351
tri 7947 290 7963 306 sw
rect 8217 290 8247 351
rect 7917 260 8023 290
tri 8023 260 8053 290 sw
rect 7917 159 7947 260
tri 7947 244 7963 260 nw
tri 8007 244 8023 260 ne
tri 7947 159 7963 175 sw
tri 8007 159 8023 175 se
rect 8023 159 8053 260
tri 8112 260 8142 290 se
rect 8142 260 8247 290
rect 8112 166 8142 260
tri 8142 244 8158 260 nw
tri 8201 244 8217 260 ne
tri 8142 166 8158 182 sw
tri 8201 166 8217 182 se
rect 8217 166 8247 260
tri 7917 129 7947 159 ne
rect 7947 129 8023 159
tri 8023 129 8053 159 nw
tri 8112 136 8142 166 ne
rect 8142 136 8217 166
tri 8217 136 8247 166 nw
rect 8419 298 8449 351
tri 8449 298 8465 314 sw
rect 8419 268 8525 298
tri 8525 268 8555 298 sw
rect 8419 167 8449 268
tri 8449 252 8465 268 nw
tri 8509 252 8525 268 ne
tri 8449 167 8465 183 sw
tri 8509 167 8525 183 se
rect 8525 167 8555 268
tri 8419 137 8449 167 ne
rect 8449 137 8525 167
tri 8525 137 8555 167 nw
rect 8879 290 8909 351
tri 8909 290 8925 306 sw
rect 9179 290 9209 351
rect 8879 260 8985 290
tri 8985 260 9015 290 sw
rect 8879 159 8909 260
tri 8909 244 8925 260 nw
tri 8969 244 8985 260 ne
tri 8909 159 8925 175 sw
tri 8969 159 8985 175 se
rect 8985 159 9015 260
tri 9074 260 9104 290 se
rect 9104 260 9209 290
rect 9074 166 9104 260
tri 9104 244 9120 260 nw
tri 9163 244 9179 260 ne
tri 9104 166 9120 182 sw
tri 9163 166 9179 182 se
rect 9179 166 9209 260
tri 8879 129 8909 159 ne
rect 8909 129 8985 159
tri 8985 129 9015 159 nw
tri 9074 136 9104 166 ne
rect 9104 136 9179 166
tri 9179 136 9209 166 nw
rect 9381 298 9411 351
tri 9411 298 9427 314 sw
rect 9381 268 9487 298
tri 9487 268 9517 298 sw
rect 9381 167 9411 268
tri 9411 252 9427 268 nw
tri 9471 252 9487 268 ne
tri 9411 167 9427 183 sw
tri 9471 167 9487 183 se
rect 9487 167 9517 268
tri 9381 137 9411 167 ne
rect 9411 137 9487 167
tri 9487 137 9517 167 nw
rect 9862 288 9892 349
tri 9892 288 9908 304 sw
rect 10056 296 10086 349
tri 10086 296 10102 312 sw
rect 9862 258 9968 288
tri 9968 258 9998 288 sw
rect 10056 266 10162 296
tri 10162 266 10192 296 sw
rect 9862 157 9892 258
tri 9892 242 9908 258 nw
tri 9952 242 9968 258 ne
tri 9892 157 9908 173 sw
tri 9952 157 9968 173 se
rect 9968 157 9998 258
rect 10056 165 10086 266
tri 10086 250 10102 266 nw
tri 10146 250 10162 266 ne
tri 10086 165 10102 181 sw
tri 10146 165 10162 181 se
rect 10162 165 10192 266
tri 9862 127 9892 157 ne
rect 9892 127 9968 157
tri 9968 127 9998 157 nw
tri 10056 135 10086 165 ne
rect 10086 135 10162 165
tri 10162 135 10192 165 nw
rect 10507 290 10537 351
tri 10537 290 10553 306 sw
rect 10807 290 10837 351
rect 10507 260 10613 290
tri 10613 260 10643 290 sw
rect 10507 159 10537 260
tri 10537 244 10553 260 nw
tri 10597 244 10613 260 ne
tri 10537 159 10553 175 sw
tri 10597 159 10613 175 se
rect 10613 159 10643 260
tri 10702 260 10732 290 se
rect 10732 260 10837 290
rect 10702 166 10732 260
tri 10732 244 10748 260 nw
tri 10791 244 10807 260 ne
tri 10732 166 10748 182 sw
tri 10791 166 10807 182 se
rect 10807 166 10837 260
tri 10507 129 10537 159 ne
rect 10537 129 10613 159
tri 10613 129 10643 159 nw
tri 10702 136 10732 166 ne
rect 10732 136 10807 166
tri 10807 136 10837 166 nw
rect 11009 298 11039 351
tri 11039 298 11055 314 sw
rect 11009 268 11115 298
tri 11115 268 11145 298 sw
rect 11009 167 11039 268
tri 11039 252 11055 268 nw
tri 11099 252 11115 268 ne
tri 11039 167 11055 183 sw
tri 11099 167 11115 183 se
rect 11115 167 11145 268
tri 11009 137 11039 167 ne
rect 11039 137 11115 167
tri 11115 137 11145 167 nw
rect 11469 290 11499 351
tri 11499 290 11515 306 sw
rect 11769 290 11799 351
rect 11469 260 11575 290
tri 11575 260 11605 290 sw
rect 11469 159 11499 260
tri 11499 244 11515 260 nw
tri 11559 244 11575 260 ne
tri 11499 159 11515 175 sw
tri 11559 159 11575 175 se
rect 11575 159 11605 260
tri 11664 260 11694 290 se
rect 11694 260 11799 290
rect 11664 166 11694 260
tri 11694 244 11710 260 nw
tri 11753 244 11769 260 ne
tri 11694 166 11710 182 sw
tri 11753 166 11769 182 se
rect 11769 166 11799 260
tri 11469 129 11499 159 ne
rect 11499 129 11575 159
tri 11575 129 11605 159 nw
tri 11664 136 11694 166 ne
rect 11694 136 11769 166
tri 11769 136 11799 166 nw
rect 11971 298 12001 351
tri 12001 298 12017 314 sw
rect 11971 268 12077 298
tri 12077 268 12107 298 sw
rect 11971 167 12001 268
tri 12001 252 12017 268 nw
tri 12061 252 12077 268 ne
tri 12001 167 12017 183 sw
tri 12061 167 12077 183 se
rect 12077 167 12107 268
tri 11971 137 12001 167 ne
rect 12001 137 12077 167
tri 12077 137 12107 167 nw
rect 12452 288 12482 349
tri 12482 288 12498 304 sw
rect 12646 296 12676 349
tri 12676 296 12692 312 sw
rect 12452 258 12558 288
tri 12558 258 12588 288 sw
rect 12646 266 12752 296
tri 12752 266 12782 296 sw
rect 12452 157 12482 258
tri 12482 242 12498 258 nw
tri 12542 242 12558 258 ne
tri 12482 157 12498 173 sw
tri 12542 157 12558 173 se
rect 12558 157 12588 258
rect 12646 165 12676 266
tri 12676 250 12692 266 nw
tri 12736 250 12752 266 ne
tri 12676 165 12692 181 sw
tri 12736 165 12752 181 se
rect 12752 165 12782 266
tri 12452 127 12482 157 ne
rect 12482 127 12558 157
tri 12558 127 12588 157 nw
tri 12646 135 12676 165 ne
rect 12676 135 12752 165
tri 12752 135 12782 165 nw
rect 13097 290 13127 351
tri 13127 290 13143 306 sw
rect 13397 290 13427 351
rect 13097 260 13203 290
tri 13203 260 13233 290 sw
rect 13097 159 13127 260
tri 13127 244 13143 260 nw
tri 13187 244 13203 260 ne
tri 13127 159 13143 175 sw
tri 13187 159 13203 175 se
rect 13203 159 13233 260
tri 13292 260 13322 290 se
rect 13322 260 13427 290
rect 13292 166 13322 260
tri 13322 244 13338 260 nw
tri 13381 244 13397 260 ne
tri 13322 166 13338 182 sw
tri 13381 166 13397 182 se
rect 13397 166 13427 260
tri 13097 129 13127 159 ne
rect 13127 129 13203 159
tri 13203 129 13233 159 nw
tri 13292 136 13322 166 ne
rect 13322 136 13397 166
tri 13397 136 13427 166 nw
rect 13599 298 13629 351
tri 13629 298 13645 314 sw
rect 13599 268 13705 298
tri 13705 268 13735 298 sw
rect 13599 167 13629 268
tri 13629 252 13645 268 nw
tri 13689 252 13705 268 ne
tri 13629 167 13645 183 sw
tri 13689 167 13705 183 se
rect 13705 167 13735 268
tri 13599 137 13629 167 ne
rect 13629 137 13705 167
tri 13705 137 13735 167 nw
rect 14059 290 14089 351
tri 14089 290 14105 306 sw
rect 14359 290 14389 351
rect 14059 260 14165 290
tri 14165 260 14195 290 sw
rect 14059 159 14089 260
tri 14089 244 14105 260 nw
tri 14149 244 14165 260 ne
tri 14089 159 14105 175 sw
tri 14149 159 14165 175 se
rect 14165 159 14195 260
tri 14254 260 14284 290 se
rect 14284 260 14389 290
rect 14254 166 14284 260
tri 14284 244 14300 260 nw
tri 14343 244 14359 260 ne
tri 14284 166 14300 182 sw
tri 14343 166 14359 182 se
rect 14359 166 14389 260
tri 14059 129 14089 159 ne
rect 14089 129 14165 159
tri 14165 129 14195 159 nw
tri 14254 136 14284 166 ne
rect 14284 136 14359 166
tri 14359 136 14389 166 nw
rect 14561 298 14591 351
tri 14591 298 14607 314 sw
rect 14561 268 14667 298
tri 14667 268 14697 298 sw
rect 14561 167 14591 268
tri 14591 252 14607 268 nw
tri 14651 252 14667 268 ne
tri 14591 167 14607 183 sw
tri 14651 167 14667 183 se
rect 14667 167 14697 268
tri 14561 137 14591 167 ne
rect 14591 137 14667 167
tri 14667 137 14697 167 nw
rect 15042 288 15072 349
tri 15072 288 15088 304 sw
rect 15236 296 15266 349
tri 15266 296 15282 312 sw
rect 15042 258 15148 288
tri 15148 258 15178 288 sw
rect 15236 266 15342 296
tri 15342 266 15372 296 sw
rect 15042 157 15072 258
tri 15072 242 15088 258 nw
tri 15132 242 15148 258 ne
tri 15072 157 15088 173 sw
tri 15132 157 15148 173 se
rect 15148 157 15178 258
rect 15236 165 15266 266
tri 15266 250 15282 266 nw
tri 15326 250 15342 266 ne
tri 15266 165 15282 181 sw
tri 15326 165 15342 181 se
rect 15342 165 15372 266
tri 15042 127 15072 157 ne
rect 15072 127 15148 157
tri 15148 127 15178 157 nw
tri 15236 135 15266 165 ne
rect 15266 135 15342 165
tri 15342 135 15372 165 nw
rect 15708 288 15738 349
tri 15738 288 15754 304 sw
rect 15902 296 15932 349
tri 15932 296 15948 312 sw
rect 15708 258 15814 288
tri 15814 258 15844 288 sw
rect 15902 266 16008 296
tri 16008 266 16038 296 sw
rect 15708 157 15738 258
tri 15738 242 15754 258 nw
tri 15798 242 15814 258 ne
tri 15738 157 15754 173 sw
tri 15798 157 15814 173 se
rect 15814 157 15844 258
rect 15902 165 15932 266
tri 15932 250 15948 266 nw
tri 15992 250 16008 266 ne
tri 15932 165 15948 181 sw
tri 15992 165 16008 181 se
rect 16008 165 16038 266
tri 15708 127 15738 157 ne
rect 15738 127 15814 157
tri 15814 127 15844 157 nw
tri 15902 135 15932 165 ne
rect 15932 135 16008 165
tri 16008 135 16038 165 nw
rect 16374 288 16404 349
tri 16404 288 16420 304 sw
tri 16658 296 16674 312 se
rect 16674 296 16704 349
rect 16374 258 16480 288
tri 16480 258 16510 288 sw
tri 16568 266 16598 296 se
rect 16598 266 16704 296
rect 16374 157 16404 258
tri 16404 242 16420 258 nw
tri 16464 242 16480 258 ne
tri 16404 157 16420 173 sw
tri 16464 157 16480 173 se
rect 16480 157 16510 258
rect 16568 165 16598 266
tri 16598 250 16614 266 nw
tri 16658 250 16674 266 ne
tri 16598 165 16614 181 sw
tri 16658 165 16674 181 se
rect 16674 165 16704 266
tri 16374 127 16404 157 ne
rect 16404 127 16480 157
tri 16480 127 16510 157 nw
tri 16568 135 16598 165 ne
rect 16598 135 16674 165
tri 16674 135 16704 165 nw
rect 17040 288 17070 349
tri 17070 288 17086 304 sw
rect 17234 296 17264 349
tri 17264 296 17280 312 sw
rect 17040 258 17146 288
tri 17146 258 17176 288 sw
rect 17234 266 17340 296
tri 17340 266 17370 296 sw
rect 17040 157 17070 258
tri 17070 242 17086 258 nw
tri 17130 242 17146 258 ne
tri 17070 157 17086 173 sw
tri 17130 157 17146 173 se
rect 17146 157 17176 258
rect 17234 251 17265 266
tri 17265 251 17280 266 nw
tri 17324 251 17339 266 ne
rect 17339 251 17370 266
rect 17234 165 17264 251
tri 17264 165 17280 181 sw
tri 17324 165 17340 181 se
rect 17340 165 17370 251
tri 17040 127 17070 157 ne
rect 17070 127 17146 157
tri 17146 127 17176 157 nw
tri 17234 135 17264 165 ne
rect 17264 135 17340 165
tri 17340 135 17370 165 nw
rect 17693 297 17723 350
tri 17723 297 17739 313 sw
rect 17693 267 17799 297
tri 17799 267 17829 297 sw
rect 17693 166 17723 267
tri 17723 251 17739 267 nw
tri 17783 251 17799 267 ne
tri 17723 166 17739 182 sw
tri 17783 166 17799 182 se
rect 17799 166 17829 267
tri 17693 136 17723 166 ne
rect 17723 136 17799 166
tri 17799 136 17829 166 nw
<< pmos >>
rect 247 1004 277 1404
rect 335 1004 365 1404
rect 423 1004 453 1404
rect 511 1004 541 1404
rect 599 1004 629 1404
rect 687 1004 717 1404
rect 1209 1004 1239 1404
rect 1297 1004 1327 1404
rect 1385 1004 1415 1404
rect 1473 1004 1503 1404
rect 1561 1004 1591 1404
rect 1649 1004 1679 1404
rect 2111 1004 2141 1404
rect 2199 1004 2229 1404
rect 2287 1004 2317 1404
rect 2375 1004 2405 1404
rect 2837 1004 2867 1404
rect 2925 1004 2955 1404
rect 3013 1004 3043 1404
rect 3101 1004 3131 1404
rect 3189 1004 3219 1404
rect 3277 1004 3307 1404
rect 3799 1004 3829 1404
rect 3887 1004 3917 1404
rect 3975 1004 4005 1404
rect 4063 1004 4093 1404
rect 4151 1004 4181 1404
rect 4239 1004 4269 1404
rect 4701 1004 4731 1404
rect 4789 1004 4819 1404
rect 4877 1004 4907 1404
rect 4965 1004 4995 1404
rect 5427 1004 5457 1404
rect 5515 1004 5545 1404
rect 5603 1004 5633 1404
rect 5691 1004 5721 1404
rect 5779 1004 5809 1404
rect 5867 1004 5897 1404
rect 6389 1004 6419 1404
rect 6477 1004 6507 1404
rect 6565 1004 6595 1404
rect 6653 1004 6683 1404
rect 6741 1004 6771 1404
rect 6829 1004 6859 1404
rect 7291 1004 7321 1404
rect 7379 1004 7409 1404
rect 7467 1004 7497 1404
rect 7555 1004 7585 1404
rect 8017 1004 8047 1404
rect 8105 1004 8135 1404
rect 8193 1004 8223 1404
rect 8281 1004 8311 1404
rect 8369 1004 8399 1404
rect 8457 1004 8487 1404
rect 8979 1004 9009 1404
rect 9067 1004 9097 1404
rect 9155 1004 9185 1404
rect 9243 1004 9273 1404
rect 9331 1004 9361 1404
rect 9419 1004 9449 1404
rect 9881 1004 9911 1404
rect 9969 1004 9999 1404
rect 10057 1004 10087 1404
rect 10145 1004 10175 1404
rect 10607 1004 10637 1404
rect 10695 1004 10725 1404
rect 10783 1004 10813 1404
rect 10871 1004 10901 1404
rect 10959 1004 10989 1404
rect 11047 1004 11077 1404
rect 11569 1004 11599 1404
rect 11657 1004 11687 1404
rect 11745 1004 11775 1404
rect 11833 1004 11863 1404
rect 11921 1004 11951 1404
rect 12009 1004 12039 1404
rect 12471 1004 12501 1404
rect 12559 1004 12589 1404
rect 12647 1004 12677 1404
rect 12735 1004 12765 1404
rect 13197 1004 13227 1404
rect 13285 1004 13315 1404
rect 13373 1004 13403 1404
rect 13461 1004 13491 1404
rect 13549 1004 13579 1404
rect 13637 1004 13667 1404
rect 14159 1004 14189 1404
rect 14247 1004 14277 1404
rect 14335 1004 14365 1404
rect 14423 1004 14453 1404
rect 14511 1004 14541 1404
rect 14599 1004 14629 1404
rect 15061 1004 15091 1404
rect 15149 1004 15179 1404
rect 15237 1004 15267 1404
rect 15325 1004 15355 1404
rect 15727 1005 15757 1405
rect 15815 1005 15845 1405
rect 15903 1005 15933 1405
rect 15991 1005 16021 1405
rect 16391 1005 16421 1405
rect 16479 1005 16509 1405
rect 16567 1005 16597 1405
rect 16655 1005 16685 1405
rect 17059 1005 17089 1405
rect 17147 1005 17177 1405
rect 17235 1005 17265 1405
rect 17323 1005 17353 1405
rect 17702 1004 17732 1404
rect 17790 1004 17820 1404
<< ndiff >>
rect 91 335 147 351
rect 91 301 101 335
rect 135 301 147 335
rect 91 263 147 301
rect 177 335 447 351
rect 177 306 198 335
tri 177 290 193 306 ne
rect 193 301 198 306
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 447 335
rect 193 290 447 301
rect 477 335 533 351
rect 477 301 489 335
rect 523 301 533 335
rect 91 229 101 263
rect 135 229 147 263
tri 253 260 283 290 ne
rect 283 263 342 290
rect 91 195 147 229
rect 91 161 101 195
rect 135 161 147 195
rect 91 129 147 161
tri 177 244 193 260 se
rect 193 244 237 260
tri 237 244 253 260 sw
rect 177 210 253 244
rect 177 176 198 210
rect 232 176 253 210
rect 177 175 253 176
tri 177 159 193 175 ne
rect 193 159 237 175
tri 237 159 253 175 nw
rect 283 229 295 263
rect 329 229 342 263
tri 342 260 372 290 nw
rect 283 195 342 229
rect 283 161 295 195
rect 329 161 342 195
tri 372 244 388 260 se
rect 388 244 431 260
tri 431 244 447 260 sw
rect 372 216 447 244
rect 372 182 393 216
rect 427 182 447 216
tri 372 166 388 182 ne
rect 388 166 431 182
tri 431 166 447 182 nw
tri 147 129 177 159 sw
tri 253 129 283 159 se
rect 283 136 342 161
tri 342 136 372 166 sw
tri 447 136 477 166 se
rect 477 136 533 301
rect 283 129 533 136
rect 91 125 533 129
rect 91 91 101 125
rect 135 91 295 125
rect 329 91 392 125
rect 426 91 489 125
rect 523 91 533 125
rect 91 75 533 91
rect 593 335 649 351
rect 593 301 603 335
rect 637 301 649 335
rect 593 263 649 301
rect 679 314 841 351
tri 679 298 695 314 ne
rect 695 298 841 314
tri 755 268 785 298 ne
rect 593 229 603 263
rect 637 229 649 263
rect 593 195 649 229
rect 593 161 603 195
rect 637 161 649 195
tri 679 252 695 268 se
rect 695 252 739 268
tri 739 252 755 268 sw
rect 679 219 755 252
rect 679 185 700 219
rect 734 185 755 219
rect 679 183 755 185
tri 679 167 695 183 ne
rect 695 167 739 183
tri 739 167 755 183 nw
rect 785 263 841 298
rect 785 229 797 263
rect 831 229 841 263
rect 785 195 841 229
rect 593 137 649 161
tri 649 137 679 167 sw
tri 755 137 785 167 se
rect 785 161 797 195
rect 831 161 841 195
rect 785 137 841 161
rect 593 125 841 137
rect 593 91 603 125
rect 637 91 700 125
rect 734 91 797 125
rect 831 91 841 125
rect 593 75 841 91
rect 1053 335 1109 351
rect 1053 301 1063 335
rect 1097 301 1109 335
rect 1053 263 1109 301
rect 1139 335 1409 351
rect 1139 306 1160 335
tri 1139 290 1155 306 ne
rect 1155 301 1160 306
rect 1194 301 1257 335
rect 1291 301 1354 335
rect 1388 301 1409 335
rect 1155 290 1409 301
rect 1439 335 1495 351
rect 1439 301 1451 335
rect 1485 301 1495 335
rect 1053 229 1063 263
rect 1097 229 1109 263
tri 1215 260 1245 290 ne
rect 1245 263 1304 290
rect 1053 195 1109 229
rect 1053 161 1063 195
rect 1097 161 1109 195
rect 1053 129 1109 161
tri 1139 244 1155 260 se
rect 1155 244 1199 260
tri 1199 244 1215 260 sw
rect 1139 210 1215 244
rect 1139 176 1160 210
rect 1194 176 1215 210
rect 1139 175 1215 176
tri 1139 159 1155 175 ne
rect 1155 159 1199 175
tri 1199 159 1215 175 nw
rect 1245 229 1257 263
rect 1291 229 1304 263
tri 1304 260 1334 290 nw
rect 1245 195 1304 229
rect 1245 161 1257 195
rect 1291 161 1304 195
tri 1334 244 1350 260 se
rect 1350 244 1393 260
tri 1393 244 1409 260 sw
rect 1334 216 1409 244
rect 1334 182 1355 216
rect 1389 182 1409 216
tri 1334 166 1350 182 ne
rect 1350 166 1393 182
tri 1393 166 1409 182 nw
tri 1109 129 1139 159 sw
tri 1215 129 1245 159 se
rect 1245 136 1304 161
tri 1304 136 1334 166 sw
tri 1409 136 1439 166 se
rect 1439 136 1495 301
rect 1245 129 1495 136
rect 1053 125 1495 129
rect 1053 91 1063 125
rect 1097 91 1257 125
rect 1291 91 1354 125
rect 1388 91 1451 125
rect 1485 91 1495 125
rect 1053 75 1495 91
rect 1555 335 1611 351
rect 1555 301 1565 335
rect 1599 301 1611 335
rect 1555 263 1611 301
rect 1641 314 1803 351
tri 1641 298 1657 314 ne
rect 1657 298 1803 314
tri 1717 268 1747 298 ne
rect 1555 229 1565 263
rect 1599 229 1611 263
rect 1555 195 1611 229
rect 1555 161 1565 195
rect 1599 161 1611 195
tri 1641 252 1657 268 se
rect 1657 252 1701 268
tri 1701 252 1717 268 sw
rect 1641 219 1717 252
rect 1641 185 1662 219
rect 1696 185 1717 219
rect 1641 183 1717 185
tri 1641 167 1657 183 ne
rect 1657 167 1701 183
tri 1701 167 1717 183 nw
rect 1747 263 1803 298
rect 1747 229 1759 263
rect 1793 229 1803 263
rect 1747 195 1803 229
rect 1555 137 1611 161
tri 1611 137 1641 167 sw
tri 1717 137 1747 167 se
rect 1747 161 1759 195
rect 1793 161 1803 195
rect 1747 137 1803 161
rect 1555 125 1803 137
rect 1555 91 1565 125
rect 1599 91 1662 125
rect 1696 91 1759 125
rect 1793 91 1803 125
rect 1555 75 1803 91
rect 2036 333 2092 349
rect 2036 299 2046 333
rect 2080 299 2092 333
rect 2036 261 2092 299
rect 2122 333 2286 349
rect 2122 304 2143 333
tri 2122 288 2138 304 ne
rect 2138 299 2143 304
rect 2177 299 2240 333
rect 2274 299 2286 333
rect 2138 288 2286 299
rect 2316 312 2478 349
tri 2316 296 2332 312 ne
rect 2332 296 2478 312
rect 2036 227 2046 261
rect 2080 227 2092 261
tri 2198 258 2228 288 ne
rect 2228 261 2286 288
tri 2392 266 2422 296 ne
rect 2036 193 2092 227
rect 2036 159 2046 193
rect 2080 159 2092 193
rect 2036 127 2092 159
tri 2122 242 2138 258 se
rect 2138 242 2182 258
tri 2182 242 2198 258 sw
rect 2122 208 2198 242
rect 2122 174 2143 208
rect 2177 174 2198 208
rect 2122 173 2198 174
tri 2122 157 2138 173 ne
rect 2138 157 2182 173
tri 2182 157 2198 173 nw
rect 2228 227 2240 261
rect 2274 227 2286 261
rect 2228 193 2286 227
rect 2228 159 2240 193
rect 2274 159 2286 193
tri 2316 250 2332 266 se
rect 2332 250 2376 266
tri 2376 250 2392 266 sw
rect 2316 217 2392 250
rect 2316 183 2337 217
rect 2371 183 2392 217
rect 2316 181 2392 183
tri 2316 165 2332 181 ne
rect 2332 165 2376 181
tri 2376 165 2392 181 nw
rect 2422 261 2478 296
rect 2422 227 2434 261
rect 2468 227 2478 261
rect 2422 193 2478 227
tri 2092 127 2122 157 sw
tri 2198 127 2228 157 se
rect 2228 135 2286 159
tri 2286 135 2316 165 sw
tri 2392 135 2422 165 se
rect 2422 159 2434 193
rect 2468 159 2478 193
rect 2422 135 2478 159
rect 2228 127 2478 135
rect 2036 123 2478 127
rect 2036 89 2046 123
rect 2080 89 2240 123
rect 2274 89 2337 123
rect 2371 89 2434 123
rect 2468 89 2478 123
rect 2036 73 2478 89
rect 2681 335 2737 351
rect 2681 301 2691 335
rect 2725 301 2737 335
rect 2681 263 2737 301
rect 2767 335 3037 351
rect 2767 306 2788 335
tri 2767 290 2783 306 ne
rect 2783 301 2788 306
rect 2822 301 2885 335
rect 2919 301 2982 335
rect 3016 301 3037 335
rect 2783 290 3037 301
rect 3067 335 3123 351
rect 3067 301 3079 335
rect 3113 301 3123 335
rect 2681 229 2691 263
rect 2725 229 2737 263
tri 2843 260 2873 290 ne
rect 2873 263 2932 290
rect 2681 195 2737 229
rect 2681 161 2691 195
rect 2725 161 2737 195
rect 2681 129 2737 161
tri 2767 244 2783 260 se
rect 2783 244 2827 260
tri 2827 244 2843 260 sw
rect 2767 210 2843 244
rect 2767 176 2788 210
rect 2822 176 2843 210
rect 2767 175 2843 176
tri 2767 159 2783 175 ne
rect 2783 159 2827 175
tri 2827 159 2843 175 nw
rect 2873 229 2885 263
rect 2919 229 2932 263
tri 2932 260 2962 290 nw
rect 2873 195 2932 229
rect 2873 161 2885 195
rect 2919 161 2932 195
tri 2962 244 2978 260 se
rect 2978 244 3021 260
tri 3021 244 3037 260 sw
rect 2962 216 3037 244
rect 2962 182 2983 216
rect 3017 182 3037 216
tri 2962 166 2978 182 ne
rect 2978 166 3021 182
tri 3021 166 3037 182 nw
tri 2737 129 2767 159 sw
tri 2843 129 2873 159 se
rect 2873 136 2932 161
tri 2932 136 2962 166 sw
tri 3037 136 3067 166 se
rect 3067 136 3123 301
rect 2873 129 3123 136
rect 2681 125 3123 129
rect 2681 91 2691 125
rect 2725 91 2885 125
rect 2919 91 2982 125
rect 3016 91 3079 125
rect 3113 91 3123 125
rect 2681 75 3123 91
rect 3183 335 3239 351
rect 3183 301 3193 335
rect 3227 301 3239 335
rect 3183 263 3239 301
rect 3269 314 3431 351
tri 3269 298 3285 314 ne
rect 3285 298 3431 314
tri 3345 268 3375 298 ne
rect 3183 229 3193 263
rect 3227 229 3239 263
rect 3183 195 3239 229
rect 3183 161 3193 195
rect 3227 161 3239 195
tri 3269 252 3285 268 se
rect 3285 252 3329 268
tri 3329 252 3345 268 sw
rect 3269 219 3345 252
rect 3269 185 3290 219
rect 3324 185 3345 219
rect 3269 183 3345 185
tri 3269 167 3285 183 ne
rect 3285 167 3329 183
tri 3329 167 3345 183 nw
rect 3375 263 3431 298
rect 3375 229 3387 263
rect 3421 229 3431 263
rect 3375 195 3431 229
rect 3183 137 3239 161
tri 3239 137 3269 167 sw
tri 3345 137 3375 167 se
rect 3375 161 3387 195
rect 3421 161 3431 195
rect 3375 137 3431 161
rect 3183 125 3431 137
rect 3183 91 3193 125
rect 3227 91 3290 125
rect 3324 91 3387 125
rect 3421 91 3431 125
rect 3183 75 3431 91
rect 3643 335 3699 351
rect 3643 301 3653 335
rect 3687 301 3699 335
rect 3643 263 3699 301
rect 3729 335 3999 351
rect 3729 306 3750 335
tri 3729 290 3745 306 ne
rect 3745 301 3750 306
rect 3784 301 3847 335
rect 3881 301 3944 335
rect 3978 301 3999 335
rect 3745 290 3999 301
rect 4029 335 4085 351
rect 4029 301 4041 335
rect 4075 301 4085 335
rect 3643 229 3653 263
rect 3687 229 3699 263
tri 3805 260 3835 290 ne
rect 3835 263 3894 290
rect 3643 195 3699 229
rect 3643 161 3653 195
rect 3687 161 3699 195
rect 3643 129 3699 161
tri 3729 244 3745 260 se
rect 3745 244 3789 260
tri 3789 244 3805 260 sw
rect 3729 210 3805 244
rect 3729 176 3750 210
rect 3784 176 3805 210
rect 3729 175 3805 176
tri 3729 159 3745 175 ne
rect 3745 159 3789 175
tri 3789 159 3805 175 nw
rect 3835 229 3847 263
rect 3881 229 3894 263
tri 3894 260 3924 290 nw
rect 3835 195 3894 229
rect 3835 161 3847 195
rect 3881 161 3894 195
tri 3924 244 3940 260 se
rect 3940 244 3983 260
tri 3983 244 3999 260 sw
rect 3924 216 3999 244
rect 3924 182 3945 216
rect 3979 182 3999 216
tri 3924 166 3940 182 ne
rect 3940 166 3983 182
tri 3983 166 3999 182 nw
tri 3699 129 3729 159 sw
tri 3805 129 3835 159 se
rect 3835 136 3894 161
tri 3894 136 3924 166 sw
tri 3999 136 4029 166 se
rect 4029 136 4085 301
rect 3835 129 4085 136
rect 3643 125 4085 129
rect 3643 91 3653 125
rect 3687 91 3847 125
rect 3881 91 3944 125
rect 3978 91 4041 125
rect 4075 91 4085 125
rect 3643 75 4085 91
rect 4145 335 4201 351
rect 4145 301 4155 335
rect 4189 301 4201 335
rect 4145 263 4201 301
rect 4231 314 4393 351
tri 4231 298 4247 314 ne
rect 4247 298 4393 314
tri 4307 268 4337 298 ne
rect 4145 229 4155 263
rect 4189 229 4201 263
rect 4145 195 4201 229
rect 4145 161 4155 195
rect 4189 161 4201 195
tri 4231 252 4247 268 se
rect 4247 252 4291 268
tri 4291 252 4307 268 sw
rect 4231 219 4307 252
rect 4231 185 4252 219
rect 4286 185 4307 219
rect 4231 183 4307 185
tri 4231 167 4247 183 ne
rect 4247 167 4291 183
tri 4291 167 4307 183 nw
rect 4337 263 4393 298
rect 4337 229 4349 263
rect 4383 229 4393 263
rect 4337 195 4393 229
rect 4145 137 4201 161
tri 4201 137 4231 167 sw
tri 4307 137 4337 167 se
rect 4337 161 4349 195
rect 4383 161 4393 195
rect 4337 137 4393 161
rect 4145 125 4393 137
rect 4145 91 4155 125
rect 4189 91 4252 125
rect 4286 91 4349 125
rect 4383 91 4393 125
rect 4145 75 4393 91
rect 4626 333 4682 349
rect 4626 299 4636 333
rect 4670 299 4682 333
rect 4626 261 4682 299
rect 4712 333 4876 349
rect 4712 304 4733 333
tri 4712 288 4728 304 ne
rect 4728 299 4733 304
rect 4767 299 4830 333
rect 4864 299 4876 333
rect 4728 288 4876 299
rect 4906 312 5068 349
tri 4906 296 4922 312 ne
rect 4922 296 5068 312
rect 4626 227 4636 261
rect 4670 227 4682 261
tri 4788 258 4818 288 ne
rect 4818 261 4876 288
tri 4982 266 5012 296 ne
rect 4626 193 4682 227
rect 4626 159 4636 193
rect 4670 159 4682 193
rect 4626 127 4682 159
tri 4712 242 4728 258 se
rect 4728 242 4772 258
tri 4772 242 4788 258 sw
rect 4712 208 4788 242
rect 4712 174 4733 208
rect 4767 174 4788 208
rect 4712 173 4788 174
tri 4712 157 4728 173 ne
rect 4728 157 4772 173
tri 4772 157 4788 173 nw
rect 4818 227 4830 261
rect 4864 227 4876 261
rect 4818 193 4876 227
rect 4818 159 4830 193
rect 4864 159 4876 193
tri 4906 250 4922 266 se
rect 4922 250 4966 266
tri 4966 250 4982 266 sw
rect 4906 217 4982 250
rect 4906 183 4927 217
rect 4961 183 4982 217
rect 4906 181 4982 183
tri 4906 165 4922 181 ne
rect 4922 165 4966 181
tri 4966 165 4982 181 nw
rect 5012 261 5068 296
rect 5012 227 5024 261
rect 5058 227 5068 261
rect 5012 193 5068 227
tri 4682 127 4712 157 sw
tri 4788 127 4818 157 se
rect 4818 135 4876 159
tri 4876 135 4906 165 sw
tri 4982 135 5012 165 se
rect 5012 159 5024 193
rect 5058 159 5068 193
rect 5012 135 5068 159
rect 4818 127 5068 135
rect 4626 123 5068 127
rect 4626 89 4636 123
rect 4670 89 4830 123
rect 4864 89 4927 123
rect 4961 89 5024 123
rect 5058 89 5068 123
rect 4626 73 5068 89
rect 5271 335 5327 351
rect 5271 301 5281 335
rect 5315 301 5327 335
rect 5271 263 5327 301
rect 5357 335 5627 351
rect 5357 306 5378 335
tri 5357 290 5373 306 ne
rect 5373 301 5378 306
rect 5412 301 5475 335
rect 5509 301 5572 335
rect 5606 301 5627 335
rect 5373 290 5627 301
rect 5657 335 5713 351
rect 5657 301 5669 335
rect 5703 301 5713 335
rect 5271 229 5281 263
rect 5315 229 5327 263
tri 5433 260 5463 290 ne
rect 5463 263 5522 290
rect 5271 195 5327 229
rect 5271 161 5281 195
rect 5315 161 5327 195
rect 5271 129 5327 161
tri 5357 244 5373 260 se
rect 5373 244 5417 260
tri 5417 244 5433 260 sw
rect 5357 210 5433 244
rect 5357 176 5378 210
rect 5412 176 5433 210
rect 5357 175 5433 176
tri 5357 159 5373 175 ne
rect 5373 159 5417 175
tri 5417 159 5433 175 nw
rect 5463 229 5475 263
rect 5509 229 5522 263
tri 5522 260 5552 290 nw
rect 5463 195 5522 229
rect 5463 161 5475 195
rect 5509 161 5522 195
tri 5552 244 5568 260 se
rect 5568 244 5611 260
tri 5611 244 5627 260 sw
rect 5552 216 5627 244
rect 5552 182 5573 216
rect 5607 182 5627 216
tri 5552 166 5568 182 ne
rect 5568 166 5611 182
tri 5611 166 5627 182 nw
tri 5327 129 5357 159 sw
tri 5433 129 5463 159 se
rect 5463 136 5522 161
tri 5522 136 5552 166 sw
tri 5627 136 5657 166 se
rect 5657 136 5713 301
rect 5463 129 5713 136
rect 5271 125 5713 129
rect 5271 91 5281 125
rect 5315 91 5475 125
rect 5509 91 5572 125
rect 5606 91 5669 125
rect 5703 91 5713 125
rect 5271 75 5713 91
rect 5773 335 5829 351
rect 5773 301 5783 335
rect 5817 301 5829 335
rect 5773 263 5829 301
rect 5859 314 6021 351
tri 5859 298 5875 314 ne
rect 5875 298 6021 314
tri 5935 268 5965 298 ne
rect 5773 229 5783 263
rect 5817 229 5829 263
rect 5773 195 5829 229
rect 5773 161 5783 195
rect 5817 161 5829 195
tri 5859 252 5875 268 se
rect 5875 252 5919 268
tri 5919 252 5935 268 sw
rect 5859 219 5935 252
rect 5859 185 5880 219
rect 5914 185 5935 219
rect 5859 183 5935 185
tri 5859 167 5875 183 ne
rect 5875 167 5919 183
tri 5919 167 5935 183 nw
rect 5965 263 6021 298
rect 5965 229 5977 263
rect 6011 229 6021 263
rect 5965 195 6021 229
rect 5773 137 5829 161
tri 5829 137 5859 167 sw
tri 5935 137 5965 167 se
rect 5965 161 5977 195
rect 6011 161 6021 195
rect 5965 137 6021 161
rect 5773 125 6021 137
rect 5773 91 5783 125
rect 5817 91 5880 125
rect 5914 91 5977 125
rect 6011 91 6021 125
rect 5773 75 6021 91
rect 6233 335 6289 351
rect 6233 301 6243 335
rect 6277 301 6289 335
rect 6233 263 6289 301
rect 6319 335 6589 351
rect 6319 306 6340 335
tri 6319 290 6335 306 ne
rect 6335 301 6340 306
rect 6374 301 6437 335
rect 6471 301 6534 335
rect 6568 301 6589 335
rect 6335 290 6589 301
rect 6619 335 6675 351
rect 6619 301 6631 335
rect 6665 301 6675 335
rect 6233 229 6243 263
rect 6277 229 6289 263
tri 6395 260 6425 290 ne
rect 6425 263 6484 290
rect 6233 195 6289 229
rect 6233 161 6243 195
rect 6277 161 6289 195
rect 6233 129 6289 161
tri 6319 244 6335 260 se
rect 6335 244 6379 260
tri 6379 244 6395 260 sw
rect 6319 210 6395 244
rect 6319 176 6340 210
rect 6374 176 6395 210
rect 6319 175 6395 176
tri 6319 159 6335 175 ne
rect 6335 159 6379 175
tri 6379 159 6395 175 nw
rect 6425 229 6437 263
rect 6471 229 6484 263
tri 6484 260 6514 290 nw
rect 6425 195 6484 229
rect 6425 161 6437 195
rect 6471 161 6484 195
tri 6514 244 6530 260 se
rect 6530 244 6573 260
tri 6573 244 6589 260 sw
rect 6514 216 6589 244
rect 6514 182 6535 216
rect 6569 182 6589 216
tri 6514 166 6530 182 ne
rect 6530 166 6573 182
tri 6573 166 6589 182 nw
tri 6289 129 6319 159 sw
tri 6395 129 6425 159 se
rect 6425 136 6484 161
tri 6484 136 6514 166 sw
tri 6589 136 6619 166 se
rect 6619 136 6675 301
rect 6425 129 6675 136
rect 6233 125 6675 129
rect 6233 91 6243 125
rect 6277 91 6437 125
rect 6471 91 6534 125
rect 6568 91 6631 125
rect 6665 91 6675 125
rect 6233 75 6675 91
rect 6735 335 6791 351
rect 6735 301 6745 335
rect 6779 301 6791 335
rect 6735 263 6791 301
rect 6821 314 6983 351
tri 6821 298 6837 314 ne
rect 6837 298 6983 314
tri 6897 268 6927 298 ne
rect 6735 229 6745 263
rect 6779 229 6791 263
rect 6735 195 6791 229
rect 6735 161 6745 195
rect 6779 161 6791 195
tri 6821 252 6837 268 se
rect 6837 252 6881 268
tri 6881 252 6897 268 sw
rect 6821 219 6897 252
rect 6821 185 6842 219
rect 6876 185 6897 219
rect 6821 183 6897 185
tri 6821 167 6837 183 ne
rect 6837 167 6881 183
tri 6881 167 6897 183 nw
rect 6927 263 6983 298
rect 6927 229 6939 263
rect 6973 229 6983 263
rect 6927 195 6983 229
rect 6735 137 6791 161
tri 6791 137 6821 167 sw
tri 6897 137 6927 167 se
rect 6927 161 6939 195
rect 6973 161 6983 195
rect 6927 137 6983 161
rect 6735 125 6983 137
rect 6735 91 6745 125
rect 6779 91 6842 125
rect 6876 91 6939 125
rect 6973 91 6983 125
rect 6735 75 6983 91
rect 7216 333 7272 349
rect 7216 299 7226 333
rect 7260 299 7272 333
rect 7216 261 7272 299
rect 7302 333 7466 349
rect 7302 304 7323 333
tri 7302 288 7318 304 ne
rect 7318 299 7323 304
rect 7357 299 7420 333
rect 7454 299 7466 333
rect 7318 288 7466 299
rect 7496 312 7658 349
tri 7496 296 7512 312 ne
rect 7512 296 7658 312
rect 7216 227 7226 261
rect 7260 227 7272 261
tri 7378 258 7408 288 ne
rect 7408 261 7466 288
tri 7572 266 7602 296 ne
rect 7216 193 7272 227
rect 7216 159 7226 193
rect 7260 159 7272 193
rect 7216 127 7272 159
tri 7302 242 7318 258 se
rect 7318 242 7362 258
tri 7362 242 7378 258 sw
rect 7302 208 7378 242
rect 7302 174 7323 208
rect 7357 174 7378 208
rect 7302 173 7378 174
tri 7302 157 7318 173 ne
rect 7318 157 7362 173
tri 7362 157 7378 173 nw
rect 7408 227 7420 261
rect 7454 227 7466 261
rect 7408 193 7466 227
rect 7408 159 7420 193
rect 7454 159 7466 193
tri 7496 250 7512 266 se
rect 7512 250 7556 266
tri 7556 250 7572 266 sw
rect 7496 217 7572 250
rect 7496 183 7517 217
rect 7551 183 7572 217
rect 7496 181 7572 183
tri 7496 165 7512 181 ne
rect 7512 165 7556 181
tri 7556 165 7572 181 nw
rect 7602 261 7658 296
rect 7602 227 7614 261
rect 7648 227 7658 261
rect 7602 193 7658 227
tri 7272 127 7302 157 sw
tri 7378 127 7408 157 se
rect 7408 135 7466 159
tri 7466 135 7496 165 sw
tri 7572 135 7602 165 se
rect 7602 159 7614 193
rect 7648 159 7658 193
rect 7602 135 7658 159
rect 7408 127 7658 135
rect 7216 123 7658 127
rect 7216 89 7226 123
rect 7260 89 7420 123
rect 7454 89 7517 123
rect 7551 89 7614 123
rect 7648 89 7658 123
rect 7216 73 7658 89
rect 7861 335 7917 351
rect 7861 301 7871 335
rect 7905 301 7917 335
rect 7861 263 7917 301
rect 7947 335 8217 351
rect 7947 306 7968 335
tri 7947 290 7963 306 ne
rect 7963 301 7968 306
rect 8002 301 8065 335
rect 8099 301 8162 335
rect 8196 301 8217 335
rect 7963 290 8217 301
rect 8247 335 8303 351
rect 8247 301 8259 335
rect 8293 301 8303 335
rect 7861 229 7871 263
rect 7905 229 7917 263
tri 8023 260 8053 290 ne
rect 8053 263 8112 290
rect 7861 195 7917 229
rect 7861 161 7871 195
rect 7905 161 7917 195
rect 7861 129 7917 161
tri 7947 244 7963 260 se
rect 7963 244 8007 260
tri 8007 244 8023 260 sw
rect 7947 210 8023 244
rect 7947 176 7968 210
rect 8002 176 8023 210
rect 7947 175 8023 176
tri 7947 159 7963 175 ne
rect 7963 159 8007 175
tri 8007 159 8023 175 nw
rect 8053 229 8065 263
rect 8099 229 8112 263
tri 8112 260 8142 290 nw
rect 8053 195 8112 229
rect 8053 161 8065 195
rect 8099 161 8112 195
tri 8142 244 8158 260 se
rect 8158 244 8201 260
tri 8201 244 8217 260 sw
rect 8142 216 8217 244
rect 8142 182 8163 216
rect 8197 182 8217 216
tri 8142 166 8158 182 ne
rect 8158 166 8201 182
tri 8201 166 8217 182 nw
tri 7917 129 7947 159 sw
tri 8023 129 8053 159 se
rect 8053 136 8112 161
tri 8112 136 8142 166 sw
tri 8217 136 8247 166 se
rect 8247 136 8303 301
rect 8053 129 8303 136
rect 7861 125 8303 129
rect 7861 91 7871 125
rect 7905 91 8065 125
rect 8099 91 8162 125
rect 8196 91 8259 125
rect 8293 91 8303 125
rect 7861 75 8303 91
rect 8363 335 8419 351
rect 8363 301 8373 335
rect 8407 301 8419 335
rect 8363 263 8419 301
rect 8449 314 8611 351
tri 8449 298 8465 314 ne
rect 8465 298 8611 314
tri 8525 268 8555 298 ne
rect 8363 229 8373 263
rect 8407 229 8419 263
rect 8363 195 8419 229
rect 8363 161 8373 195
rect 8407 161 8419 195
tri 8449 252 8465 268 se
rect 8465 252 8509 268
tri 8509 252 8525 268 sw
rect 8449 219 8525 252
rect 8449 185 8470 219
rect 8504 185 8525 219
rect 8449 183 8525 185
tri 8449 167 8465 183 ne
rect 8465 167 8509 183
tri 8509 167 8525 183 nw
rect 8555 263 8611 298
rect 8555 229 8567 263
rect 8601 229 8611 263
rect 8555 195 8611 229
rect 8363 137 8419 161
tri 8419 137 8449 167 sw
tri 8525 137 8555 167 se
rect 8555 161 8567 195
rect 8601 161 8611 195
rect 8555 137 8611 161
rect 8363 125 8611 137
rect 8363 91 8373 125
rect 8407 91 8470 125
rect 8504 91 8567 125
rect 8601 91 8611 125
rect 8363 75 8611 91
rect 8823 335 8879 351
rect 8823 301 8833 335
rect 8867 301 8879 335
rect 8823 263 8879 301
rect 8909 335 9179 351
rect 8909 306 8930 335
tri 8909 290 8925 306 ne
rect 8925 301 8930 306
rect 8964 301 9027 335
rect 9061 301 9124 335
rect 9158 301 9179 335
rect 8925 290 9179 301
rect 9209 335 9265 351
rect 9209 301 9221 335
rect 9255 301 9265 335
rect 8823 229 8833 263
rect 8867 229 8879 263
tri 8985 260 9015 290 ne
rect 9015 263 9074 290
rect 8823 195 8879 229
rect 8823 161 8833 195
rect 8867 161 8879 195
rect 8823 129 8879 161
tri 8909 244 8925 260 se
rect 8925 244 8969 260
tri 8969 244 8985 260 sw
rect 8909 210 8985 244
rect 8909 176 8930 210
rect 8964 176 8985 210
rect 8909 175 8985 176
tri 8909 159 8925 175 ne
rect 8925 159 8969 175
tri 8969 159 8985 175 nw
rect 9015 229 9027 263
rect 9061 229 9074 263
tri 9074 260 9104 290 nw
rect 9015 195 9074 229
rect 9015 161 9027 195
rect 9061 161 9074 195
tri 9104 244 9120 260 se
rect 9120 244 9163 260
tri 9163 244 9179 260 sw
rect 9104 216 9179 244
rect 9104 182 9125 216
rect 9159 182 9179 216
tri 9104 166 9120 182 ne
rect 9120 166 9163 182
tri 9163 166 9179 182 nw
tri 8879 129 8909 159 sw
tri 8985 129 9015 159 se
rect 9015 136 9074 161
tri 9074 136 9104 166 sw
tri 9179 136 9209 166 se
rect 9209 136 9265 301
rect 9015 129 9265 136
rect 8823 125 9265 129
rect 8823 91 8833 125
rect 8867 91 9027 125
rect 9061 91 9124 125
rect 9158 91 9221 125
rect 9255 91 9265 125
rect 8823 75 9265 91
rect 9325 335 9381 351
rect 9325 301 9335 335
rect 9369 301 9381 335
rect 9325 263 9381 301
rect 9411 314 9573 351
tri 9411 298 9427 314 ne
rect 9427 298 9573 314
tri 9487 268 9517 298 ne
rect 9325 229 9335 263
rect 9369 229 9381 263
rect 9325 195 9381 229
rect 9325 161 9335 195
rect 9369 161 9381 195
tri 9411 252 9427 268 se
rect 9427 252 9471 268
tri 9471 252 9487 268 sw
rect 9411 219 9487 252
rect 9411 185 9432 219
rect 9466 185 9487 219
rect 9411 183 9487 185
tri 9411 167 9427 183 ne
rect 9427 167 9471 183
tri 9471 167 9487 183 nw
rect 9517 263 9573 298
rect 9517 229 9529 263
rect 9563 229 9573 263
rect 9517 195 9573 229
rect 9325 137 9381 161
tri 9381 137 9411 167 sw
tri 9487 137 9517 167 se
rect 9517 161 9529 195
rect 9563 161 9573 195
rect 9517 137 9573 161
rect 9325 125 9573 137
rect 9325 91 9335 125
rect 9369 91 9432 125
rect 9466 91 9529 125
rect 9563 91 9573 125
rect 9325 75 9573 91
rect 9806 333 9862 349
rect 9806 299 9816 333
rect 9850 299 9862 333
rect 9806 261 9862 299
rect 9892 333 10056 349
rect 9892 304 9913 333
tri 9892 288 9908 304 ne
rect 9908 299 9913 304
rect 9947 299 10010 333
rect 10044 299 10056 333
rect 9908 288 10056 299
rect 10086 312 10248 349
tri 10086 296 10102 312 ne
rect 10102 296 10248 312
rect 9806 227 9816 261
rect 9850 227 9862 261
tri 9968 258 9998 288 ne
rect 9998 261 10056 288
tri 10162 266 10192 296 ne
rect 9806 193 9862 227
rect 9806 159 9816 193
rect 9850 159 9862 193
rect 9806 127 9862 159
tri 9892 242 9908 258 se
rect 9908 242 9952 258
tri 9952 242 9968 258 sw
rect 9892 208 9968 242
rect 9892 174 9913 208
rect 9947 174 9968 208
rect 9892 173 9968 174
tri 9892 157 9908 173 ne
rect 9908 157 9952 173
tri 9952 157 9968 173 nw
rect 9998 227 10010 261
rect 10044 227 10056 261
rect 9998 193 10056 227
rect 9998 159 10010 193
rect 10044 159 10056 193
tri 10086 250 10102 266 se
rect 10102 250 10146 266
tri 10146 250 10162 266 sw
rect 10086 217 10162 250
rect 10086 183 10107 217
rect 10141 183 10162 217
rect 10086 181 10162 183
tri 10086 165 10102 181 ne
rect 10102 165 10146 181
tri 10146 165 10162 181 nw
rect 10192 261 10248 296
rect 10192 227 10204 261
rect 10238 227 10248 261
rect 10192 193 10248 227
tri 9862 127 9892 157 sw
tri 9968 127 9998 157 se
rect 9998 135 10056 159
tri 10056 135 10086 165 sw
tri 10162 135 10192 165 se
rect 10192 159 10204 193
rect 10238 159 10248 193
rect 10192 135 10248 159
rect 9998 127 10248 135
rect 9806 123 10248 127
rect 9806 89 9816 123
rect 9850 89 10010 123
rect 10044 89 10107 123
rect 10141 89 10204 123
rect 10238 89 10248 123
rect 9806 73 10248 89
rect 10451 335 10507 351
rect 10451 301 10461 335
rect 10495 301 10507 335
rect 10451 263 10507 301
rect 10537 335 10807 351
rect 10537 306 10558 335
tri 10537 290 10553 306 ne
rect 10553 301 10558 306
rect 10592 301 10655 335
rect 10689 301 10752 335
rect 10786 301 10807 335
rect 10553 290 10807 301
rect 10837 335 10893 351
rect 10837 301 10849 335
rect 10883 301 10893 335
rect 10451 229 10461 263
rect 10495 229 10507 263
tri 10613 260 10643 290 ne
rect 10643 263 10702 290
rect 10451 195 10507 229
rect 10451 161 10461 195
rect 10495 161 10507 195
rect 10451 129 10507 161
tri 10537 244 10553 260 se
rect 10553 244 10597 260
tri 10597 244 10613 260 sw
rect 10537 210 10613 244
rect 10537 176 10558 210
rect 10592 176 10613 210
rect 10537 175 10613 176
tri 10537 159 10553 175 ne
rect 10553 159 10597 175
tri 10597 159 10613 175 nw
rect 10643 229 10655 263
rect 10689 229 10702 263
tri 10702 260 10732 290 nw
rect 10643 195 10702 229
rect 10643 161 10655 195
rect 10689 161 10702 195
tri 10732 244 10748 260 se
rect 10748 244 10791 260
tri 10791 244 10807 260 sw
rect 10732 216 10807 244
rect 10732 182 10753 216
rect 10787 182 10807 216
tri 10732 166 10748 182 ne
rect 10748 166 10791 182
tri 10791 166 10807 182 nw
tri 10507 129 10537 159 sw
tri 10613 129 10643 159 se
rect 10643 136 10702 161
tri 10702 136 10732 166 sw
tri 10807 136 10837 166 se
rect 10837 136 10893 301
rect 10643 129 10893 136
rect 10451 125 10893 129
rect 10451 91 10461 125
rect 10495 91 10655 125
rect 10689 91 10752 125
rect 10786 91 10849 125
rect 10883 91 10893 125
rect 10451 75 10893 91
rect 10953 335 11009 351
rect 10953 301 10963 335
rect 10997 301 11009 335
rect 10953 263 11009 301
rect 11039 314 11201 351
tri 11039 298 11055 314 ne
rect 11055 298 11201 314
tri 11115 268 11145 298 ne
rect 10953 229 10963 263
rect 10997 229 11009 263
rect 10953 195 11009 229
rect 10953 161 10963 195
rect 10997 161 11009 195
tri 11039 252 11055 268 se
rect 11055 252 11099 268
tri 11099 252 11115 268 sw
rect 11039 219 11115 252
rect 11039 185 11060 219
rect 11094 185 11115 219
rect 11039 183 11115 185
tri 11039 167 11055 183 ne
rect 11055 167 11099 183
tri 11099 167 11115 183 nw
rect 11145 263 11201 298
rect 11145 229 11157 263
rect 11191 229 11201 263
rect 11145 195 11201 229
rect 10953 137 11009 161
tri 11009 137 11039 167 sw
tri 11115 137 11145 167 se
rect 11145 161 11157 195
rect 11191 161 11201 195
rect 11145 137 11201 161
rect 10953 125 11201 137
rect 10953 91 10963 125
rect 10997 91 11060 125
rect 11094 91 11157 125
rect 11191 91 11201 125
rect 10953 75 11201 91
rect 11413 335 11469 351
rect 11413 301 11423 335
rect 11457 301 11469 335
rect 11413 263 11469 301
rect 11499 335 11769 351
rect 11499 306 11520 335
tri 11499 290 11515 306 ne
rect 11515 301 11520 306
rect 11554 301 11617 335
rect 11651 301 11714 335
rect 11748 301 11769 335
rect 11515 290 11769 301
rect 11799 335 11855 351
rect 11799 301 11811 335
rect 11845 301 11855 335
rect 11413 229 11423 263
rect 11457 229 11469 263
tri 11575 260 11605 290 ne
rect 11605 263 11664 290
rect 11413 195 11469 229
rect 11413 161 11423 195
rect 11457 161 11469 195
rect 11413 129 11469 161
tri 11499 244 11515 260 se
rect 11515 244 11559 260
tri 11559 244 11575 260 sw
rect 11499 210 11575 244
rect 11499 176 11520 210
rect 11554 176 11575 210
rect 11499 175 11575 176
tri 11499 159 11515 175 ne
rect 11515 159 11559 175
tri 11559 159 11575 175 nw
rect 11605 229 11617 263
rect 11651 229 11664 263
tri 11664 260 11694 290 nw
rect 11605 195 11664 229
rect 11605 161 11617 195
rect 11651 161 11664 195
tri 11694 244 11710 260 se
rect 11710 244 11753 260
tri 11753 244 11769 260 sw
rect 11694 216 11769 244
rect 11694 182 11715 216
rect 11749 182 11769 216
tri 11694 166 11710 182 ne
rect 11710 166 11753 182
tri 11753 166 11769 182 nw
tri 11469 129 11499 159 sw
tri 11575 129 11605 159 se
rect 11605 136 11664 161
tri 11664 136 11694 166 sw
tri 11769 136 11799 166 se
rect 11799 136 11855 301
rect 11605 129 11855 136
rect 11413 125 11855 129
rect 11413 91 11423 125
rect 11457 91 11617 125
rect 11651 91 11714 125
rect 11748 91 11811 125
rect 11845 91 11855 125
rect 11413 75 11855 91
rect 11915 335 11971 351
rect 11915 301 11925 335
rect 11959 301 11971 335
rect 11915 263 11971 301
rect 12001 314 12163 351
tri 12001 298 12017 314 ne
rect 12017 298 12163 314
tri 12077 268 12107 298 ne
rect 11915 229 11925 263
rect 11959 229 11971 263
rect 11915 195 11971 229
rect 11915 161 11925 195
rect 11959 161 11971 195
tri 12001 252 12017 268 se
rect 12017 252 12061 268
tri 12061 252 12077 268 sw
rect 12001 219 12077 252
rect 12001 185 12022 219
rect 12056 185 12077 219
rect 12001 183 12077 185
tri 12001 167 12017 183 ne
rect 12017 167 12061 183
tri 12061 167 12077 183 nw
rect 12107 263 12163 298
rect 12107 229 12119 263
rect 12153 229 12163 263
rect 12107 195 12163 229
rect 11915 137 11971 161
tri 11971 137 12001 167 sw
tri 12077 137 12107 167 se
rect 12107 161 12119 195
rect 12153 161 12163 195
rect 12107 137 12163 161
rect 11915 125 12163 137
rect 11915 91 11925 125
rect 11959 91 12022 125
rect 12056 91 12119 125
rect 12153 91 12163 125
rect 11915 75 12163 91
rect 12396 333 12452 349
rect 12396 299 12406 333
rect 12440 299 12452 333
rect 12396 261 12452 299
rect 12482 333 12646 349
rect 12482 304 12503 333
tri 12482 288 12498 304 ne
rect 12498 299 12503 304
rect 12537 299 12600 333
rect 12634 299 12646 333
rect 12498 288 12646 299
rect 12676 312 12838 349
tri 12676 296 12692 312 ne
rect 12692 296 12838 312
rect 12396 227 12406 261
rect 12440 227 12452 261
tri 12558 258 12588 288 ne
rect 12588 261 12646 288
tri 12752 266 12782 296 ne
rect 12396 193 12452 227
rect 12396 159 12406 193
rect 12440 159 12452 193
rect 12396 127 12452 159
tri 12482 242 12498 258 se
rect 12498 242 12542 258
tri 12542 242 12558 258 sw
rect 12482 208 12558 242
rect 12482 174 12503 208
rect 12537 174 12558 208
rect 12482 173 12558 174
tri 12482 157 12498 173 ne
rect 12498 157 12542 173
tri 12542 157 12558 173 nw
rect 12588 227 12600 261
rect 12634 227 12646 261
rect 12588 193 12646 227
rect 12588 159 12600 193
rect 12634 159 12646 193
tri 12676 250 12692 266 se
rect 12692 250 12736 266
tri 12736 250 12752 266 sw
rect 12676 217 12752 250
rect 12676 183 12697 217
rect 12731 183 12752 217
rect 12676 181 12752 183
tri 12676 165 12692 181 ne
rect 12692 165 12736 181
tri 12736 165 12752 181 nw
rect 12782 261 12838 296
rect 12782 227 12794 261
rect 12828 227 12838 261
rect 12782 193 12838 227
tri 12452 127 12482 157 sw
tri 12558 127 12588 157 se
rect 12588 135 12646 159
tri 12646 135 12676 165 sw
tri 12752 135 12782 165 se
rect 12782 159 12794 193
rect 12828 159 12838 193
rect 12782 135 12838 159
rect 12588 127 12838 135
rect 12396 123 12838 127
rect 12396 89 12406 123
rect 12440 89 12600 123
rect 12634 89 12697 123
rect 12731 89 12794 123
rect 12828 89 12838 123
rect 12396 73 12838 89
rect 13041 335 13097 351
rect 13041 301 13051 335
rect 13085 301 13097 335
rect 13041 263 13097 301
rect 13127 335 13397 351
rect 13127 306 13148 335
tri 13127 290 13143 306 ne
rect 13143 301 13148 306
rect 13182 301 13245 335
rect 13279 301 13342 335
rect 13376 301 13397 335
rect 13143 290 13397 301
rect 13427 335 13483 351
rect 13427 301 13439 335
rect 13473 301 13483 335
rect 13041 229 13051 263
rect 13085 229 13097 263
tri 13203 260 13233 290 ne
rect 13233 263 13292 290
rect 13041 195 13097 229
rect 13041 161 13051 195
rect 13085 161 13097 195
rect 13041 129 13097 161
tri 13127 244 13143 260 se
rect 13143 244 13187 260
tri 13187 244 13203 260 sw
rect 13127 210 13203 244
rect 13127 176 13148 210
rect 13182 176 13203 210
rect 13127 175 13203 176
tri 13127 159 13143 175 ne
rect 13143 159 13187 175
tri 13187 159 13203 175 nw
rect 13233 229 13245 263
rect 13279 229 13292 263
tri 13292 260 13322 290 nw
rect 13233 195 13292 229
rect 13233 161 13245 195
rect 13279 161 13292 195
tri 13322 244 13338 260 se
rect 13338 244 13381 260
tri 13381 244 13397 260 sw
rect 13322 216 13397 244
rect 13322 182 13343 216
rect 13377 182 13397 216
tri 13322 166 13338 182 ne
rect 13338 166 13381 182
tri 13381 166 13397 182 nw
tri 13097 129 13127 159 sw
tri 13203 129 13233 159 se
rect 13233 136 13292 161
tri 13292 136 13322 166 sw
tri 13397 136 13427 166 se
rect 13427 136 13483 301
rect 13233 129 13483 136
rect 13041 125 13483 129
rect 13041 91 13051 125
rect 13085 91 13245 125
rect 13279 91 13342 125
rect 13376 91 13439 125
rect 13473 91 13483 125
rect 13041 75 13483 91
rect 13543 335 13599 351
rect 13543 301 13553 335
rect 13587 301 13599 335
rect 13543 263 13599 301
rect 13629 314 13791 351
tri 13629 298 13645 314 ne
rect 13645 298 13791 314
tri 13705 268 13735 298 ne
rect 13543 229 13553 263
rect 13587 229 13599 263
rect 13543 195 13599 229
rect 13543 161 13553 195
rect 13587 161 13599 195
tri 13629 252 13645 268 se
rect 13645 252 13689 268
tri 13689 252 13705 268 sw
rect 13629 219 13705 252
rect 13629 185 13650 219
rect 13684 185 13705 219
rect 13629 183 13705 185
tri 13629 167 13645 183 ne
rect 13645 167 13689 183
tri 13689 167 13705 183 nw
rect 13735 263 13791 298
rect 13735 229 13747 263
rect 13781 229 13791 263
rect 13735 195 13791 229
rect 13543 137 13599 161
tri 13599 137 13629 167 sw
tri 13705 137 13735 167 se
rect 13735 161 13747 195
rect 13781 161 13791 195
rect 13735 137 13791 161
rect 13543 125 13791 137
rect 13543 91 13553 125
rect 13587 91 13650 125
rect 13684 91 13747 125
rect 13781 91 13791 125
rect 13543 75 13791 91
rect 14003 335 14059 351
rect 14003 301 14013 335
rect 14047 301 14059 335
rect 14003 263 14059 301
rect 14089 335 14359 351
rect 14089 306 14110 335
tri 14089 290 14105 306 ne
rect 14105 301 14110 306
rect 14144 301 14207 335
rect 14241 301 14304 335
rect 14338 301 14359 335
rect 14105 290 14359 301
rect 14389 335 14445 351
rect 14389 301 14401 335
rect 14435 301 14445 335
rect 14003 229 14013 263
rect 14047 229 14059 263
tri 14165 260 14195 290 ne
rect 14195 263 14254 290
rect 14003 195 14059 229
rect 14003 161 14013 195
rect 14047 161 14059 195
rect 14003 129 14059 161
tri 14089 244 14105 260 se
rect 14105 244 14149 260
tri 14149 244 14165 260 sw
rect 14089 210 14165 244
rect 14089 176 14110 210
rect 14144 176 14165 210
rect 14089 175 14165 176
tri 14089 159 14105 175 ne
rect 14105 159 14149 175
tri 14149 159 14165 175 nw
rect 14195 229 14207 263
rect 14241 229 14254 263
tri 14254 260 14284 290 nw
rect 14195 195 14254 229
rect 14195 161 14207 195
rect 14241 161 14254 195
tri 14284 244 14300 260 se
rect 14300 244 14343 260
tri 14343 244 14359 260 sw
rect 14284 216 14359 244
rect 14284 182 14305 216
rect 14339 182 14359 216
tri 14284 166 14300 182 ne
rect 14300 166 14343 182
tri 14343 166 14359 182 nw
tri 14059 129 14089 159 sw
tri 14165 129 14195 159 se
rect 14195 136 14254 161
tri 14254 136 14284 166 sw
tri 14359 136 14389 166 se
rect 14389 136 14445 301
rect 14195 129 14445 136
rect 14003 125 14445 129
rect 14003 91 14013 125
rect 14047 91 14207 125
rect 14241 91 14304 125
rect 14338 91 14401 125
rect 14435 91 14445 125
rect 14003 75 14445 91
rect 14505 335 14561 351
rect 14505 301 14515 335
rect 14549 301 14561 335
rect 14505 263 14561 301
rect 14591 314 14753 351
tri 14591 298 14607 314 ne
rect 14607 298 14753 314
tri 14667 268 14697 298 ne
rect 14505 229 14515 263
rect 14549 229 14561 263
rect 14505 195 14561 229
rect 14505 161 14515 195
rect 14549 161 14561 195
tri 14591 252 14607 268 se
rect 14607 252 14651 268
tri 14651 252 14667 268 sw
rect 14591 219 14667 252
rect 14591 185 14612 219
rect 14646 185 14667 219
rect 14591 183 14667 185
tri 14591 167 14607 183 ne
rect 14607 167 14651 183
tri 14651 167 14667 183 nw
rect 14697 263 14753 298
rect 14697 229 14709 263
rect 14743 229 14753 263
rect 14697 195 14753 229
rect 14505 137 14561 161
tri 14561 137 14591 167 sw
tri 14667 137 14697 167 se
rect 14697 161 14709 195
rect 14743 161 14753 195
rect 14697 137 14753 161
rect 14505 125 14753 137
rect 14505 91 14515 125
rect 14549 91 14612 125
rect 14646 91 14709 125
rect 14743 91 14753 125
rect 14505 75 14753 91
rect 14986 333 15042 349
rect 14986 299 14996 333
rect 15030 299 15042 333
rect 14986 261 15042 299
rect 15072 333 15236 349
rect 15072 304 15093 333
tri 15072 288 15088 304 ne
rect 15088 299 15093 304
rect 15127 299 15190 333
rect 15224 299 15236 333
rect 15088 288 15236 299
rect 15266 312 15428 349
tri 15266 296 15282 312 ne
rect 15282 296 15428 312
rect 14986 227 14996 261
rect 15030 227 15042 261
tri 15148 258 15178 288 ne
rect 15178 261 15236 288
tri 15342 266 15372 296 ne
rect 14986 193 15042 227
rect 14986 159 14996 193
rect 15030 159 15042 193
rect 14986 127 15042 159
tri 15072 242 15088 258 se
rect 15088 242 15132 258
tri 15132 242 15148 258 sw
rect 15072 208 15148 242
rect 15072 174 15093 208
rect 15127 174 15148 208
rect 15072 173 15148 174
tri 15072 157 15088 173 ne
rect 15088 157 15132 173
tri 15132 157 15148 173 nw
rect 15178 227 15190 261
rect 15224 227 15236 261
rect 15178 193 15236 227
rect 15178 159 15190 193
rect 15224 159 15236 193
tri 15266 250 15282 266 se
rect 15282 250 15326 266
tri 15326 250 15342 266 sw
rect 15266 217 15342 250
rect 15266 183 15287 217
rect 15321 183 15342 217
rect 15266 181 15342 183
tri 15266 165 15282 181 ne
rect 15282 165 15326 181
tri 15326 165 15342 181 nw
rect 15372 261 15428 296
rect 15372 227 15384 261
rect 15418 227 15428 261
rect 15372 193 15428 227
tri 15042 127 15072 157 sw
tri 15148 127 15178 157 se
rect 15178 135 15236 159
tri 15236 135 15266 165 sw
tri 15342 135 15372 165 se
rect 15372 159 15384 193
rect 15418 159 15428 193
rect 15372 135 15428 159
rect 15178 127 15428 135
rect 14986 123 15428 127
rect 14986 89 14996 123
rect 15030 89 15190 123
rect 15224 89 15287 123
rect 15321 89 15384 123
rect 15418 89 15428 123
rect 14986 73 15428 89
rect 15652 333 15708 349
rect 15652 299 15662 333
rect 15696 299 15708 333
rect 15652 261 15708 299
rect 15738 333 15902 349
rect 15738 304 15759 333
tri 15738 288 15754 304 ne
rect 15754 299 15759 304
rect 15793 299 15856 333
rect 15890 299 15902 333
rect 15754 288 15902 299
rect 15932 333 16092 349
rect 15932 312 16050 333
tri 15932 296 15948 312 ne
rect 15948 299 16050 312
rect 16084 299 16092 333
rect 15948 296 16092 299
rect 15652 227 15662 261
rect 15696 227 15708 261
tri 15814 258 15844 288 ne
rect 15844 261 15902 288
tri 16008 266 16038 296 ne
rect 15652 193 15708 227
rect 15652 159 15662 193
rect 15696 159 15708 193
rect 15652 127 15708 159
tri 15738 242 15754 258 se
rect 15754 242 15798 258
tri 15798 242 15814 258 sw
rect 15738 208 15814 242
rect 15738 174 15759 208
rect 15793 174 15814 208
rect 15738 173 15814 174
tri 15738 157 15754 173 ne
rect 15754 157 15798 173
tri 15798 157 15814 173 nw
rect 15844 227 15856 261
rect 15890 227 15902 261
rect 15844 193 15902 227
rect 15844 159 15856 193
rect 15890 159 15902 193
tri 15932 250 15948 266 se
rect 15948 250 15992 266
tri 15992 250 16008 266 sw
rect 15932 217 16008 250
rect 15932 183 15952 217
rect 15986 183 16008 217
rect 15932 181 16008 183
tri 15932 165 15948 181 ne
rect 15948 165 15992 181
tri 15992 165 16008 181 nw
rect 16038 261 16092 296
rect 16038 227 16050 261
rect 16084 227 16092 261
rect 16038 193 16092 227
tri 15708 127 15738 157 sw
tri 15814 127 15844 157 se
rect 15844 135 15902 159
tri 15902 135 15932 165 sw
tri 16008 135 16038 165 se
rect 16038 159 16050 193
rect 16084 159 16092 193
rect 16038 135 16092 159
rect 15844 127 16092 135
rect 15652 123 16092 127
rect 15652 89 15662 123
rect 15696 89 15856 123
rect 15890 89 15952 123
rect 15986 89 16050 123
rect 16084 89 16092 123
rect 15652 73 16092 89
rect 16318 333 16374 349
rect 16318 299 16328 333
rect 16362 299 16374 333
rect 16318 261 16374 299
rect 16404 333 16674 349
rect 16404 304 16425 333
tri 16404 288 16420 304 ne
rect 16420 299 16425 304
rect 16459 299 16522 333
rect 16556 312 16674 333
rect 16556 299 16658 312
rect 16420 296 16658 299
tri 16658 296 16674 312 nw
rect 16704 333 16760 349
rect 16704 299 16716 333
rect 16750 299 16760 333
rect 16420 288 16568 296
rect 16318 227 16328 261
rect 16362 227 16374 261
tri 16480 258 16510 288 ne
rect 16510 261 16568 288
tri 16568 266 16598 296 nw
rect 16318 193 16374 227
rect 16318 159 16328 193
rect 16362 159 16374 193
rect 16318 127 16374 159
tri 16404 242 16420 258 se
rect 16420 242 16464 258
tri 16464 242 16480 258 sw
rect 16404 208 16480 242
rect 16404 174 16425 208
rect 16459 174 16480 208
rect 16404 173 16480 174
tri 16404 157 16420 173 ne
rect 16420 157 16464 173
tri 16464 157 16480 173 nw
rect 16510 227 16522 261
rect 16556 227 16568 261
rect 16510 193 16568 227
rect 16510 159 16522 193
rect 16556 159 16568 193
tri 16598 250 16614 266 se
rect 16614 250 16658 266
tri 16658 250 16674 266 sw
rect 16598 217 16674 250
rect 16598 183 16619 217
rect 16653 183 16674 217
rect 16598 181 16674 183
tri 16598 165 16614 181 ne
rect 16614 165 16658 181
tri 16658 165 16674 181 nw
rect 16704 261 16760 299
rect 16704 227 16716 261
rect 16750 227 16760 261
rect 16704 193 16760 227
tri 16374 127 16404 157 sw
tri 16480 127 16510 157 se
rect 16510 135 16568 159
tri 16568 135 16598 165 sw
tri 16674 135 16704 165 se
rect 16704 159 16716 193
rect 16750 159 16760 193
rect 16704 135 16760 159
rect 16510 127 16760 135
rect 16318 123 16760 127
rect 16318 89 16328 123
rect 16362 89 16522 123
rect 16556 89 16619 123
rect 16653 89 16716 123
rect 16750 89 16760 123
rect 16318 73 16760 89
rect 16984 333 17040 349
rect 16984 299 16994 333
rect 17028 299 17040 333
rect 16984 261 17040 299
rect 17070 333 17234 349
rect 17070 304 17091 333
tri 17070 288 17086 304 ne
rect 17086 299 17091 304
rect 17125 299 17188 333
rect 17222 299 17234 333
rect 17086 288 17234 299
rect 17264 312 17426 349
tri 17264 296 17280 312 ne
rect 17280 296 17426 312
rect 16984 227 16994 261
rect 17028 227 17040 261
tri 17146 258 17176 288 ne
rect 17176 261 17234 288
tri 17340 266 17370 296 ne
rect 16984 193 17040 227
rect 16984 159 16994 193
rect 17028 159 17040 193
rect 16984 127 17040 159
tri 17070 242 17086 258 se
rect 17086 242 17130 258
tri 17130 242 17146 258 sw
rect 17070 208 17146 242
rect 17070 174 17091 208
rect 17125 174 17146 208
rect 17070 173 17146 174
tri 17070 157 17086 173 ne
rect 17086 157 17130 173
tri 17130 157 17146 173 nw
rect 17176 227 17188 261
rect 17222 227 17234 261
tri 17265 251 17280 266 se
rect 17280 251 17324 266
tri 17324 251 17339 266 sw
rect 17370 261 17426 296
rect 17176 193 17234 227
rect 17176 159 17188 193
rect 17222 159 17234 193
rect 17264 217 17340 251
rect 17264 183 17285 217
rect 17319 183 17340 217
rect 17264 181 17340 183
tri 17264 165 17280 181 ne
rect 17280 165 17324 181
tri 17324 165 17340 181 nw
rect 17370 227 17382 261
rect 17416 227 17426 261
rect 17370 193 17426 227
tri 17040 127 17070 157 sw
tri 17146 127 17176 157 se
rect 17176 135 17234 159
tri 17234 135 17264 165 sw
tri 17340 135 17370 165 se
rect 17370 159 17382 193
rect 17416 159 17426 193
rect 17370 135 17426 159
rect 17176 127 17426 135
rect 16984 123 17426 127
rect 16984 89 16994 123
rect 17028 89 17188 123
rect 17222 89 17285 123
rect 17319 89 17382 123
rect 17416 89 17426 123
rect 16984 73 17426 89
rect 17637 334 17693 350
rect 17637 300 17647 334
rect 17681 300 17693 334
rect 17637 262 17693 300
rect 17723 334 17883 350
rect 17723 313 17841 334
tri 17723 297 17739 313 ne
rect 17739 300 17841 313
rect 17875 300 17883 334
rect 17739 297 17883 300
tri 17799 267 17829 297 ne
rect 17637 228 17647 262
rect 17681 228 17693 262
rect 17637 194 17693 228
rect 17637 160 17647 194
rect 17681 160 17693 194
tri 17723 251 17739 267 se
rect 17739 251 17783 267
tri 17783 251 17799 267 sw
rect 17723 218 17799 251
rect 17723 184 17743 218
rect 17777 184 17799 218
rect 17723 182 17799 184
tri 17723 166 17739 182 ne
rect 17739 166 17783 182
tri 17783 166 17799 182 nw
rect 17829 262 17883 297
rect 17829 228 17841 262
rect 17875 228 17883 262
rect 17829 194 17883 228
rect 17637 136 17693 160
tri 17693 136 17723 166 sw
tri 17799 136 17829 166 se
rect 17829 160 17841 194
rect 17875 160 17883 194
rect 17829 136 17883 160
rect 17637 124 17883 136
rect 17637 90 17647 124
rect 17681 90 17743 124
rect 17777 90 17841 124
rect 17875 90 17883 124
rect 17637 74 17883 90
<< pdiff >>
rect 191 1366 247 1404
rect 191 1332 201 1366
rect 235 1332 247 1366
rect 191 1298 247 1332
rect 191 1264 201 1298
rect 235 1264 247 1298
rect 191 1230 247 1264
rect 191 1196 201 1230
rect 235 1196 247 1230
rect 191 1162 247 1196
rect 191 1128 201 1162
rect 235 1128 247 1162
rect 191 1093 247 1128
rect 191 1059 201 1093
rect 235 1059 247 1093
rect 191 1004 247 1059
rect 277 1366 335 1404
rect 277 1332 289 1366
rect 323 1332 335 1366
rect 277 1298 335 1332
rect 277 1264 289 1298
rect 323 1264 335 1298
rect 277 1230 335 1264
rect 277 1196 289 1230
rect 323 1196 335 1230
rect 277 1162 335 1196
rect 277 1128 289 1162
rect 323 1128 335 1162
rect 277 1093 335 1128
rect 277 1059 289 1093
rect 323 1059 335 1093
rect 277 1004 335 1059
rect 365 1366 423 1404
rect 365 1332 377 1366
rect 411 1332 423 1366
rect 365 1298 423 1332
rect 365 1264 377 1298
rect 411 1264 423 1298
rect 365 1230 423 1264
rect 365 1196 377 1230
rect 411 1196 423 1230
rect 365 1162 423 1196
rect 365 1128 377 1162
rect 411 1128 423 1162
rect 365 1004 423 1128
rect 453 1366 511 1404
rect 453 1332 465 1366
rect 499 1332 511 1366
rect 453 1298 511 1332
rect 453 1264 465 1298
rect 499 1264 511 1298
rect 453 1230 511 1264
rect 453 1196 465 1230
rect 499 1196 511 1230
rect 453 1162 511 1196
rect 453 1128 465 1162
rect 499 1128 511 1162
rect 453 1093 511 1128
rect 453 1059 465 1093
rect 499 1059 511 1093
rect 453 1004 511 1059
rect 541 1366 599 1404
rect 541 1332 553 1366
rect 587 1332 599 1366
rect 541 1298 599 1332
rect 541 1264 553 1298
rect 587 1264 599 1298
rect 541 1230 599 1264
rect 541 1196 553 1230
rect 587 1196 599 1230
rect 541 1162 599 1196
rect 541 1128 553 1162
rect 587 1128 599 1162
rect 541 1004 599 1128
rect 629 1366 687 1404
rect 629 1332 641 1366
rect 675 1332 687 1366
rect 629 1298 687 1332
rect 629 1264 641 1298
rect 675 1264 687 1298
rect 629 1230 687 1264
rect 629 1196 641 1230
rect 675 1196 687 1230
rect 629 1162 687 1196
rect 629 1128 641 1162
rect 675 1128 687 1162
rect 629 1093 687 1128
rect 629 1059 641 1093
rect 675 1059 687 1093
rect 629 1004 687 1059
rect 717 1366 771 1404
rect 717 1332 729 1366
rect 763 1332 771 1366
rect 717 1298 771 1332
rect 717 1264 729 1298
rect 763 1264 771 1298
rect 717 1230 771 1264
rect 717 1196 729 1230
rect 763 1196 771 1230
rect 717 1162 771 1196
rect 717 1128 729 1162
rect 763 1128 771 1162
rect 717 1004 771 1128
rect 1153 1366 1209 1404
rect 1153 1332 1163 1366
rect 1197 1332 1209 1366
rect 1153 1298 1209 1332
rect 1153 1264 1163 1298
rect 1197 1264 1209 1298
rect 1153 1230 1209 1264
rect 1153 1196 1163 1230
rect 1197 1196 1209 1230
rect 1153 1162 1209 1196
rect 1153 1128 1163 1162
rect 1197 1128 1209 1162
rect 1153 1093 1209 1128
rect 1153 1059 1163 1093
rect 1197 1059 1209 1093
rect 1153 1004 1209 1059
rect 1239 1366 1297 1404
rect 1239 1332 1251 1366
rect 1285 1332 1297 1366
rect 1239 1298 1297 1332
rect 1239 1264 1251 1298
rect 1285 1264 1297 1298
rect 1239 1230 1297 1264
rect 1239 1196 1251 1230
rect 1285 1196 1297 1230
rect 1239 1162 1297 1196
rect 1239 1128 1251 1162
rect 1285 1128 1297 1162
rect 1239 1093 1297 1128
rect 1239 1059 1251 1093
rect 1285 1059 1297 1093
rect 1239 1004 1297 1059
rect 1327 1366 1385 1404
rect 1327 1332 1339 1366
rect 1373 1332 1385 1366
rect 1327 1298 1385 1332
rect 1327 1264 1339 1298
rect 1373 1264 1385 1298
rect 1327 1230 1385 1264
rect 1327 1196 1339 1230
rect 1373 1196 1385 1230
rect 1327 1162 1385 1196
rect 1327 1128 1339 1162
rect 1373 1128 1385 1162
rect 1327 1004 1385 1128
rect 1415 1366 1473 1404
rect 1415 1332 1427 1366
rect 1461 1332 1473 1366
rect 1415 1298 1473 1332
rect 1415 1264 1427 1298
rect 1461 1264 1473 1298
rect 1415 1230 1473 1264
rect 1415 1196 1427 1230
rect 1461 1196 1473 1230
rect 1415 1162 1473 1196
rect 1415 1128 1427 1162
rect 1461 1128 1473 1162
rect 1415 1093 1473 1128
rect 1415 1059 1427 1093
rect 1461 1059 1473 1093
rect 1415 1004 1473 1059
rect 1503 1366 1561 1404
rect 1503 1332 1515 1366
rect 1549 1332 1561 1366
rect 1503 1298 1561 1332
rect 1503 1264 1515 1298
rect 1549 1264 1561 1298
rect 1503 1230 1561 1264
rect 1503 1196 1515 1230
rect 1549 1196 1561 1230
rect 1503 1162 1561 1196
rect 1503 1128 1515 1162
rect 1549 1128 1561 1162
rect 1503 1004 1561 1128
rect 1591 1366 1649 1404
rect 1591 1332 1603 1366
rect 1637 1332 1649 1366
rect 1591 1298 1649 1332
rect 1591 1264 1603 1298
rect 1637 1264 1649 1298
rect 1591 1230 1649 1264
rect 1591 1196 1603 1230
rect 1637 1196 1649 1230
rect 1591 1162 1649 1196
rect 1591 1128 1603 1162
rect 1637 1128 1649 1162
rect 1591 1093 1649 1128
rect 1591 1059 1603 1093
rect 1637 1059 1649 1093
rect 1591 1004 1649 1059
rect 1679 1366 1733 1404
rect 1679 1332 1691 1366
rect 1725 1332 1733 1366
rect 1679 1298 1733 1332
rect 1679 1264 1691 1298
rect 1725 1264 1733 1298
rect 1679 1230 1733 1264
rect 1679 1196 1691 1230
rect 1725 1196 1733 1230
rect 1679 1162 1733 1196
rect 1679 1128 1691 1162
rect 1725 1128 1733 1162
rect 1679 1004 1733 1128
rect 2055 1366 2111 1404
rect 2055 1332 2065 1366
rect 2099 1332 2111 1366
rect 2055 1298 2111 1332
rect 2055 1264 2065 1298
rect 2099 1264 2111 1298
rect 2055 1230 2111 1264
rect 2055 1196 2065 1230
rect 2099 1196 2111 1230
rect 2055 1162 2111 1196
rect 2055 1128 2065 1162
rect 2099 1128 2111 1162
rect 2055 1093 2111 1128
rect 2055 1059 2065 1093
rect 2099 1059 2111 1093
rect 2055 1004 2111 1059
rect 2141 1366 2199 1404
rect 2141 1332 2153 1366
rect 2187 1332 2199 1366
rect 2141 1298 2199 1332
rect 2141 1264 2153 1298
rect 2187 1264 2199 1298
rect 2141 1230 2199 1264
rect 2141 1196 2153 1230
rect 2187 1196 2199 1230
rect 2141 1162 2199 1196
rect 2141 1128 2153 1162
rect 2187 1128 2199 1162
rect 2141 1093 2199 1128
rect 2141 1059 2153 1093
rect 2187 1059 2199 1093
rect 2141 1004 2199 1059
rect 2229 1366 2287 1404
rect 2229 1332 2241 1366
rect 2275 1332 2287 1366
rect 2229 1298 2287 1332
rect 2229 1264 2241 1298
rect 2275 1264 2287 1298
rect 2229 1230 2287 1264
rect 2229 1196 2241 1230
rect 2275 1196 2287 1230
rect 2229 1162 2287 1196
rect 2229 1128 2241 1162
rect 2275 1128 2287 1162
rect 2229 1004 2287 1128
rect 2317 1366 2375 1404
rect 2317 1332 2329 1366
rect 2363 1332 2375 1366
rect 2317 1298 2375 1332
rect 2317 1264 2329 1298
rect 2363 1264 2375 1298
rect 2317 1230 2375 1264
rect 2317 1196 2329 1230
rect 2363 1196 2375 1230
rect 2317 1162 2375 1196
rect 2317 1128 2329 1162
rect 2363 1128 2375 1162
rect 2317 1093 2375 1128
rect 2317 1059 2329 1093
rect 2363 1059 2375 1093
rect 2317 1004 2375 1059
rect 2405 1366 2459 1404
rect 2405 1332 2417 1366
rect 2451 1332 2459 1366
rect 2405 1298 2459 1332
rect 2405 1264 2417 1298
rect 2451 1264 2459 1298
rect 2405 1230 2459 1264
rect 2405 1196 2417 1230
rect 2451 1196 2459 1230
rect 2405 1162 2459 1196
rect 2405 1128 2417 1162
rect 2451 1128 2459 1162
rect 2405 1004 2459 1128
rect 2781 1366 2837 1404
rect 2781 1332 2791 1366
rect 2825 1332 2837 1366
rect 2781 1298 2837 1332
rect 2781 1264 2791 1298
rect 2825 1264 2837 1298
rect 2781 1230 2837 1264
rect 2781 1196 2791 1230
rect 2825 1196 2837 1230
rect 2781 1162 2837 1196
rect 2781 1128 2791 1162
rect 2825 1128 2837 1162
rect 2781 1093 2837 1128
rect 2781 1059 2791 1093
rect 2825 1059 2837 1093
rect 2781 1004 2837 1059
rect 2867 1366 2925 1404
rect 2867 1332 2879 1366
rect 2913 1332 2925 1366
rect 2867 1298 2925 1332
rect 2867 1264 2879 1298
rect 2913 1264 2925 1298
rect 2867 1230 2925 1264
rect 2867 1196 2879 1230
rect 2913 1196 2925 1230
rect 2867 1162 2925 1196
rect 2867 1128 2879 1162
rect 2913 1128 2925 1162
rect 2867 1093 2925 1128
rect 2867 1059 2879 1093
rect 2913 1059 2925 1093
rect 2867 1004 2925 1059
rect 2955 1366 3013 1404
rect 2955 1332 2967 1366
rect 3001 1332 3013 1366
rect 2955 1298 3013 1332
rect 2955 1264 2967 1298
rect 3001 1264 3013 1298
rect 2955 1230 3013 1264
rect 2955 1196 2967 1230
rect 3001 1196 3013 1230
rect 2955 1162 3013 1196
rect 2955 1128 2967 1162
rect 3001 1128 3013 1162
rect 2955 1004 3013 1128
rect 3043 1366 3101 1404
rect 3043 1332 3055 1366
rect 3089 1332 3101 1366
rect 3043 1298 3101 1332
rect 3043 1264 3055 1298
rect 3089 1264 3101 1298
rect 3043 1230 3101 1264
rect 3043 1196 3055 1230
rect 3089 1196 3101 1230
rect 3043 1162 3101 1196
rect 3043 1128 3055 1162
rect 3089 1128 3101 1162
rect 3043 1093 3101 1128
rect 3043 1059 3055 1093
rect 3089 1059 3101 1093
rect 3043 1004 3101 1059
rect 3131 1366 3189 1404
rect 3131 1332 3143 1366
rect 3177 1332 3189 1366
rect 3131 1298 3189 1332
rect 3131 1264 3143 1298
rect 3177 1264 3189 1298
rect 3131 1230 3189 1264
rect 3131 1196 3143 1230
rect 3177 1196 3189 1230
rect 3131 1162 3189 1196
rect 3131 1128 3143 1162
rect 3177 1128 3189 1162
rect 3131 1004 3189 1128
rect 3219 1366 3277 1404
rect 3219 1332 3231 1366
rect 3265 1332 3277 1366
rect 3219 1298 3277 1332
rect 3219 1264 3231 1298
rect 3265 1264 3277 1298
rect 3219 1230 3277 1264
rect 3219 1196 3231 1230
rect 3265 1196 3277 1230
rect 3219 1162 3277 1196
rect 3219 1128 3231 1162
rect 3265 1128 3277 1162
rect 3219 1093 3277 1128
rect 3219 1059 3231 1093
rect 3265 1059 3277 1093
rect 3219 1004 3277 1059
rect 3307 1366 3361 1404
rect 3307 1332 3319 1366
rect 3353 1332 3361 1366
rect 3307 1298 3361 1332
rect 3307 1264 3319 1298
rect 3353 1264 3361 1298
rect 3307 1230 3361 1264
rect 3307 1196 3319 1230
rect 3353 1196 3361 1230
rect 3307 1162 3361 1196
rect 3307 1128 3319 1162
rect 3353 1128 3361 1162
rect 3307 1004 3361 1128
rect 3743 1366 3799 1404
rect 3743 1332 3753 1366
rect 3787 1332 3799 1366
rect 3743 1298 3799 1332
rect 3743 1264 3753 1298
rect 3787 1264 3799 1298
rect 3743 1230 3799 1264
rect 3743 1196 3753 1230
rect 3787 1196 3799 1230
rect 3743 1162 3799 1196
rect 3743 1128 3753 1162
rect 3787 1128 3799 1162
rect 3743 1093 3799 1128
rect 3743 1059 3753 1093
rect 3787 1059 3799 1093
rect 3743 1004 3799 1059
rect 3829 1366 3887 1404
rect 3829 1332 3841 1366
rect 3875 1332 3887 1366
rect 3829 1298 3887 1332
rect 3829 1264 3841 1298
rect 3875 1264 3887 1298
rect 3829 1230 3887 1264
rect 3829 1196 3841 1230
rect 3875 1196 3887 1230
rect 3829 1162 3887 1196
rect 3829 1128 3841 1162
rect 3875 1128 3887 1162
rect 3829 1093 3887 1128
rect 3829 1059 3841 1093
rect 3875 1059 3887 1093
rect 3829 1004 3887 1059
rect 3917 1366 3975 1404
rect 3917 1332 3929 1366
rect 3963 1332 3975 1366
rect 3917 1298 3975 1332
rect 3917 1264 3929 1298
rect 3963 1264 3975 1298
rect 3917 1230 3975 1264
rect 3917 1196 3929 1230
rect 3963 1196 3975 1230
rect 3917 1162 3975 1196
rect 3917 1128 3929 1162
rect 3963 1128 3975 1162
rect 3917 1004 3975 1128
rect 4005 1366 4063 1404
rect 4005 1332 4017 1366
rect 4051 1332 4063 1366
rect 4005 1298 4063 1332
rect 4005 1264 4017 1298
rect 4051 1264 4063 1298
rect 4005 1230 4063 1264
rect 4005 1196 4017 1230
rect 4051 1196 4063 1230
rect 4005 1162 4063 1196
rect 4005 1128 4017 1162
rect 4051 1128 4063 1162
rect 4005 1093 4063 1128
rect 4005 1059 4017 1093
rect 4051 1059 4063 1093
rect 4005 1004 4063 1059
rect 4093 1366 4151 1404
rect 4093 1332 4105 1366
rect 4139 1332 4151 1366
rect 4093 1298 4151 1332
rect 4093 1264 4105 1298
rect 4139 1264 4151 1298
rect 4093 1230 4151 1264
rect 4093 1196 4105 1230
rect 4139 1196 4151 1230
rect 4093 1162 4151 1196
rect 4093 1128 4105 1162
rect 4139 1128 4151 1162
rect 4093 1004 4151 1128
rect 4181 1366 4239 1404
rect 4181 1332 4193 1366
rect 4227 1332 4239 1366
rect 4181 1298 4239 1332
rect 4181 1264 4193 1298
rect 4227 1264 4239 1298
rect 4181 1230 4239 1264
rect 4181 1196 4193 1230
rect 4227 1196 4239 1230
rect 4181 1162 4239 1196
rect 4181 1128 4193 1162
rect 4227 1128 4239 1162
rect 4181 1093 4239 1128
rect 4181 1059 4193 1093
rect 4227 1059 4239 1093
rect 4181 1004 4239 1059
rect 4269 1366 4323 1404
rect 4269 1332 4281 1366
rect 4315 1332 4323 1366
rect 4269 1298 4323 1332
rect 4269 1264 4281 1298
rect 4315 1264 4323 1298
rect 4269 1230 4323 1264
rect 4269 1196 4281 1230
rect 4315 1196 4323 1230
rect 4269 1162 4323 1196
rect 4269 1128 4281 1162
rect 4315 1128 4323 1162
rect 4269 1004 4323 1128
rect 4645 1366 4701 1404
rect 4645 1332 4655 1366
rect 4689 1332 4701 1366
rect 4645 1298 4701 1332
rect 4645 1264 4655 1298
rect 4689 1264 4701 1298
rect 4645 1230 4701 1264
rect 4645 1196 4655 1230
rect 4689 1196 4701 1230
rect 4645 1162 4701 1196
rect 4645 1128 4655 1162
rect 4689 1128 4701 1162
rect 4645 1093 4701 1128
rect 4645 1059 4655 1093
rect 4689 1059 4701 1093
rect 4645 1004 4701 1059
rect 4731 1366 4789 1404
rect 4731 1332 4743 1366
rect 4777 1332 4789 1366
rect 4731 1298 4789 1332
rect 4731 1264 4743 1298
rect 4777 1264 4789 1298
rect 4731 1230 4789 1264
rect 4731 1196 4743 1230
rect 4777 1196 4789 1230
rect 4731 1162 4789 1196
rect 4731 1128 4743 1162
rect 4777 1128 4789 1162
rect 4731 1093 4789 1128
rect 4731 1059 4743 1093
rect 4777 1059 4789 1093
rect 4731 1004 4789 1059
rect 4819 1366 4877 1404
rect 4819 1332 4831 1366
rect 4865 1332 4877 1366
rect 4819 1298 4877 1332
rect 4819 1264 4831 1298
rect 4865 1264 4877 1298
rect 4819 1230 4877 1264
rect 4819 1196 4831 1230
rect 4865 1196 4877 1230
rect 4819 1162 4877 1196
rect 4819 1128 4831 1162
rect 4865 1128 4877 1162
rect 4819 1004 4877 1128
rect 4907 1366 4965 1404
rect 4907 1332 4919 1366
rect 4953 1332 4965 1366
rect 4907 1298 4965 1332
rect 4907 1264 4919 1298
rect 4953 1264 4965 1298
rect 4907 1230 4965 1264
rect 4907 1196 4919 1230
rect 4953 1196 4965 1230
rect 4907 1162 4965 1196
rect 4907 1128 4919 1162
rect 4953 1128 4965 1162
rect 4907 1093 4965 1128
rect 4907 1059 4919 1093
rect 4953 1059 4965 1093
rect 4907 1004 4965 1059
rect 4995 1366 5049 1404
rect 4995 1332 5007 1366
rect 5041 1332 5049 1366
rect 4995 1298 5049 1332
rect 4995 1264 5007 1298
rect 5041 1264 5049 1298
rect 4995 1230 5049 1264
rect 4995 1196 5007 1230
rect 5041 1196 5049 1230
rect 4995 1162 5049 1196
rect 4995 1128 5007 1162
rect 5041 1128 5049 1162
rect 4995 1004 5049 1128
rect 5371 1366 5427 1404
rect 5371 1332 5381 1366
rect 5415 1332 5427 1366
rect 5371 1298 5427 1332
rect 5371 1264 5381 1298
rect 5415 1264 5427 1298
rect 5371 1230 5427 1264
rect 5371 1196 5381 1230
rect 5415 1196 5427 1230
rect 5371 1162 5427 1196
rect 5371 1128 5381 1162
rect 5415 1128 5427 1162
rect 5371 1093 5427 1128
rect 5371 1059 5381 1093
rect 5415 1059 5427 1093
rect 5371 1004 5427 1059
rect 5457 1366 5515 1404
rect 5457 1332 5469 1366
rect 5503 1332 5515 1366
rect 5457 1298 5515 1332
rect 5457 1264 5469 1298
rect 5503 1264 5515 1298
rect 5457 1230 5515 1264
rect 5457 1196 5469 1230
rect 5503 1196 5515 1230
rect 5457 1162 5515 1196
rect 5457 1128 5469 1162
rect 5503 1128 5515 1162
rect 5457 1093 5515 1128
rect 5457 1059 5469 1093
rect 5503 1059 5515 1093
rect 5457 1004 5515 1059
rect 5545 1366 5603 1404
rect 5545 1332 5557 1366
rect 5591 1332 5603 1366
rect 5545 1298 5603 1332
rect 5545 1264 5557 1298
rect 5591 1264 5603 1298
rect 5545 1230 5603 1264
rect 5545 1196 5557 1230
rect 5591 1196 5603 1230
rect 5545 1162 5603 1196
rect 5545 1128 5557 1162
rect 5591 1128 5603 1162
rect 5545 1004 5603 1128
rect 5633 1366 5691 1404
rect 5633 1332 5645 1366
rect 5679 1332 5691 1366
rect 5633 1298 5691 1332
rect 5633 1264 5645 1298
rect 5679 1264 5691 1298
rect 5633 1230 5691 1264
rect 5633 1196 5645 1230
rect 5679 1196 5691 1230
rect 5633 1162 5691 1196
rect 5633 1128 5645 1162
rect 5679 1128 5691 1162
rect 5633 1093 5691 1128
rect 5633 1059 5645 1093
rect 5679 1059 5691 1093
rect 5633 1004 5691 1059
rect 5721 1366 5779 1404
rect 5721 1332 5733 1366
rect 5767 1332 5779 1366
rect 5721 1298 5779 1332
rect 5721 1264 5733 1298
rect 5767 1264 5779 1298
rect 5721 1230 5779 1264
rect 5721 1196 5733 1230
rect 5767 1196 5779 1230
rect 5721 1162 5779 1196
rect 5721 1128 5733 1162
rect 5767 1128 5779 1162
rect 5721 1004 5779 1128
rect 5809 1366 5867 1404
rect 5809 1332 5821 1366
rect 5855 1332 5867 1366
rect 5809 1298 5867 1332
rect 5809 1264 5821 1298
rect 5855 1264 5867 1298
rect 5809 1230 5867 1264
rect 5809 1196 5821 1230
rect 5855 1196 5867 1230
rect 5809 1162 5867 1196
rect 5809 1128 5821 1162
rect 5855 1128 5867 1162
rect 5809 1093 5867 1128
rect 5809 1059 5821 1093
rect 5855 1059 5867 1093
rect 5809 1004 5867 1059
rect 5897 1366 5951 1404
rect 5897 1332 5909 1366
rect 5943 1332 5951 1366
rect 5897 1298 5951 1332
rect 5897 1264 5909 1298
rect 5943 1264 5951 1298
rect 5897 1230 5951 1264
rect 5897 1196 5909 1230
rect 5943 1196 5951 1230
rect 5897 1162 5951 1196
rect 5897 1128 5909 1162
rect 5943 1128 5951 1162
rect 5897 1004 5951 1128
rect 6333 1366 6389 1404
rect 6333 1332 6343 1366
rect 6377 1332 6389 1366
rect 6333 1298 6389 1332
rect 6333 1264 6343 1298
rect 6377 1264 6389 1298
rect 6333 1230 6389 1264
rect 6333 1196 6343 1230
rect 6377 1196 6389 1230
rect 6333 1162 6389 1196
rect 6333 1128 6343 1162
rect 6377 1128 6389 1162
rect 6333 1093 6389 1128
rect 6333 1059 6343 1093
rect 6377 1059 6389 1093
rect 6333 1004 6389 1059
rect 6419 1366 6477 1404
rect 6419 1332 6431 1366
rect 6465 1332 6477 1366
rect 6419 1298 6477 1332
rect 6419 1264 6431 1298
rect 6465 1264 6477 1298
rect 6419 1230 6477 1264
rect 6419 1196 6431 1230
rect 6465 1196 6477 1230
rect 6419 1162 6477 1196
rect 6419 1128 6431 1162
rect 6465 1128 6477 1162
rect 6419 1093 6477 1128
rect 6419 1059 6431 1093
rect 6465 1059 6477 1093
rect 6419 1004 6477 1059
rect 6507 1366 6565 1404
rect 6507 1332 6519 1366
rect 6553 1332 6565 1366
rect 6507 1298 6565 1332
rect 6507 1264 6519 1298
rect 6553 1264 6565 1298
rect 6507 1230 6565 1264
rect 6507 1196 6519 1230
rect 6553 1196 6565 1230
rect 6507 1162 6565 1196
rect 6507 1128 6519 1162
rect 6553 1128 6565 1162
rect 6507 1004 6565 1128
rect 6595 1366 6653 1404
rect 6595 1332 6607 1366
rect 6641 1332 6653 1366
rect 6595 1298 6653 1332
rect 6595 1264 6607 1298
rect 6641 1264 6653 1298
rect 6595 1230 6653 1264
rect 6595 1196 6607 1230
rect 6641 1196 6653 1230
rect 6595 1162 6653 1196
rect 6595 1128 6607 1162
rect 6641 1128 6653 1162
rect 6595 1093 6653 1128
rect 6595 1059 6607 1093
rect 6641 1059 6653 1093
rect 6595 1004 6653 1059
rect 6683 1366 6741 1404
rect 6683 1332 6695 1366
rect 6729 1332 6741 1366
rect 6683 1298 6741 1332
rect 6683 1264 6695 1298
rect 6729 1264 6741 1298
rect 6683 1230 6741 1264
rect 6683 1196 6695 1230
rect 6729 1196 6741 1230
rect 6683 1162 6741 1196
rect 6683 1128 6695 1162
rect 6729 1128 6741 1162
rect 6683 1004 6741 1128
rect 6771 1366 6829 1404
rect 6771 1332 6783 1366
rect 6817 1332 6829 1366
rect 6771 1298 6829 1332
rect 6771 1264 6783 1298
rect 6817 1264 6829 1298
rect 6771 1230 6829 1264
rect 6771 1196 6783 1230
rect 6817 1196 6829 1230
rect 6771 1162 6829 1196
rect 6771 1128 6783 1162
rect 6817 1128 6829 1162
rect 6771 1093 6829 1128
rect 6771 1059 6783 1093
rect 6817 1059 6829 1093
rect 6771 1004 6829 1059
rect 6859 1366 6913 1404
rect 6859 1332 6871 1366
rect 6905 1332 6913 1366
rect 6859 1298 6913 1332
rect 6859 1264 6871 1298
rect 6905 1264 6913 1298
rect 6859 1230 6913 1264
rect 6859 1196 6871 1230
rect 6905 1196 6913 1230
rect 6859 1162 6913 1196
rect 6859 1128 6871 1162
rect 6905 1128 6913 1162
rect 6859 1004 6913 1128
rect 7235 1366 7291 1404
rect 7235 1332 7245 1366
rect 7279 1332 7291 1366
rect 7235 1298 7291 1332
rect 7235 1264 7245 1298
rect 7279 1264 7291 1298
rect 7235 1230 7291 1264
rect 7235 1196 7245 1230
rect 7279 1196 7291 1230
rect 7235 1162 7291 1196
rect 7235 1128 7245 1162
rect 7279 1128 7291 1162
rect 7235 1093 7291 1128
rect 7235 1059 7245 1093
rect 7279 1059 7291 1093
rect 7235 1004 7291 1059
rect 7321 1366 7379 1404
rect 7321 1332 7333 1366
rect 7367 1332 7379 1366
rect 7321 1298 7379 1332
rect 7321 1264 7333 1298
rect 7367 1264 7379 1298
rect 7321 1230 7379 1264
rect 7321 1196 7333 1230
rect 7367 1196 7379 1230
rect 7321 1162 7379 1196
rect 7321 1128 7333 1162
rect 7367 1128 7379 1162
rect 7321 1093 7379 1128
rect 7321 1059 7333 1093
rect 7367 1059 7379 1093
rect 7321 1004 7379 1059
rect 7409 1366 7467 1404
rect 7409 1332 7421 1366
rect 7455 1332 7467 1366
rect 7409 1298 7467 1332
rect 7409 1264 7421 1298
rect 7455 1264 7467 1298
rect 7409 1230 7467 1264
rect 7409 1196 7421 1230
rect 7455 1196 7467 1230
rect 7409 1162 7467 1196
rect 7409 1128 7421 1162
rect 7455 1128 7467 1162
rect 7409 1004 7467 1128
rect 7497 1366 7555 1404
rect 7497 1332 7509 1366
rect 7543 1332 7555 1366
rect 7497 1298 7555 1332
rect 7497 1264 7509 1298
rect 7543 1264 7555 1298
rect 7497 1230 7555 1264
rect 7497 1196 7509 1230
rect 7543 1196 7555 1230
rect 7497 1162 7555 1196
rect 7497 1128 7509 1162
rect 7543 1128 7555 1162
rect 7497 1093 7555 1128
rect 7497 1059 7509 1093
rect 7543 1059 7555 1093
rect 7497 1004 7555 1059
rect 7585 1366 7639 1404
rect 7585 1332 7597 1366
rect 7631 1332 7639 1366
rect 7585 1298 7639 1332
rect 7585 1264 7597 1298
rect 7631 1264 7639 1298
rect 7585 1230 7639 1264
rect 7585 1196 7597 1230
rect 7631 1196 7639 1230
rect 7585 1162 7639 1196
rect 7585 1128 7597 1162
rect 7631 1128 7639 1162
rect 7585 1004 7639 1128
rect 7961 1366 8017 1404
rect 7961 1332 7971 1366
rect 8005 1332 8017 1366
rect 7961 1298 8017 1332
rect 7961 1264 7971 1298
rect 8005 1264 8017 1298
rect 7961 1230 8017 1264
rect 7961 1196 7971 1230
rect 8005 1196 8017 1230
rect 7961 1162 8017 1196
rect 7961 1128 7971 1162
rect 8005 1128 8017 1162
rect 7961 1093 8017 1128
rect 7961 1059 7971 1093
rect 8005 1059 8017 1093
rect 7961 1004 8017 1059
rect 8047 1366 8105 1404
rect 8047 1332 8059 1366
rect 8093 1332 8105 1366
rect 8047 1298 8105 1332
rect 8047 1264 8059 1298
rect 8093 1264 8105 1298
rect 8047 1230 8105 1264
rect 8047 1196 8059 1230
rect 8093 1196 8105 1230
rect 8047 1162 8105 1196
rect 8047 1128 8059 1162
rect 8093 1128 8105 1162
rect 8047 1093 8105 1128
rect 8047 1059 8059 1093
rect 8093 1059 8105 1093
rect 8047 1004 8105 1059
rect 8135 1366 8193 1404
rect 8135 1332 8147 1366
rect 8181 1332 8193 1366
rect 8135 1298 8193 1332
rect 8135 1264 8147 1298
rect 8181 1264 8193 1298
rect 8135 1230 8193 1264
rect 8135 1196 8147 1230
rect 8181 1196 8193 1230
rect 8135 1162 8193 1196
rect 8135 1128 8147 1162
rect 8181 1128 8193 1162
rect 8135 1004 8193 1128
rect 8223 1366 8281 1404
rect 8223 1332 8235 1366
rect 8269 1332 8281 1366
rect 8223 1298 8281 1332
rect 8223 1264 8235 1298
rect 8269 1264 8281 1298
rect 8223 1230 8281 1264
rect 8223 1196 8235 1230
rect 8269 1196 8281 1230
rect 8223 1162 8281 1196
rect 8223 1128 8235 1162
rect 8269 1128 8281 1162
rect 8223 1093 8281 1128
rect 8223 1059 8235 1093
rect 8269 1059 8281 1093
rect 8223 1004 8281 1059
rect 8311 1366 8369 1404
rect 8311 1332 8323 1366
rect 8357 1332 8369 1366
rect 8311 1298 8369 1332
rect 8311 1264 8323 1298
rect 8357 1264 8369 1298
rect 8311 1230 8369 1264
rect 8311 1196 8323 1230
rect 8357 1196 8369 1230
rect 8311 1162 8369 1196
rect 8311 1128 8323 1162
rect 8357 1128 8369 1162
rect 8311 1004 8369 1128
rect 8399 1366 8457 1404
rect 8399 1332 8411 1366
rect 8445 1332 8457 1366
rect 8399 1298 8457 1332
rect 8399 1264 8411 1298
rect 8445 1264 8457 1298
rect 8399 1230 8457 1264
rect 8399 1196 8411 1230
rect 8445 1196 8457 1230
rect 8399 1162 8457 1196
rect 8399 1128 8411 1162
rect 8445 1128 8457 1162
rect 8399 1093 8457 1128
rect 8399 1059 8411 1093
rect 8445 1059 8457 1093
rect 8399 1004 8457 1059
rect 8487 1366 8541 1404
rect 8487 1332 8499 1366
rect 8533 1332 8541 1366
rect 8487 1298 8541 1332
rect 8487 1264 8499 1298
rect 8533 1264 8541 1298
rect 8487 1230 8541 1264
rect 8487 1196 8499 1230
rect 8533 1196 8541 1230
rect 8487 1162 8541 1196
rect 8487 1128 8499 1162
rect 8533 1128 8541 1162
rect 8487 1004 8541 1128
rect 8923 1366 8979 1404
rect 8923 1332 8933 1366
rect 8967 1332 8979 1366
rect 8923 1298 8979 1332
rect 8923 1264 8933 1298
rect 8967 1264 8979 1298
rect 8923 1230 8979 1264
rect 8923 1196 8933 1230
rect 8967 1196 8979 1230
rect 8923 1162 8979 1196
rect 8923 1128 8933 1162
rect 8967 1128 8979 1162
rect 8923 1093 8979 1128
rect 8923 1059 8933 1093
rect 8967 1059 8979 1093
rect 8923 1004 8979 1059
rect 9009 1366 9067 1404
rect 9009 1332 9021 1366
rect 9055 1332 9067 1366
rect 9009 1298 9067 1332
rect 9009 1264 9021 1298
rect 9055 1264 9067 1298
rect 9009 1230 9067 1264
rect 9009 1196 9021 1230
rect 9055 1196 9067 1230
rect 9009 1162 9067 1196
rect 9009 1128 9021 1162
rect 9055 1128 9067 1162
rect 9009 1093 9067 1128
rect 9009 1059 9021 1093
rect 9055 1059 9067 1093
rect 9009 1004 9067 1059
rect 9097 1366 9155 1404
rect 9097 1332 9109 1366
rect 9143 1332 9155 1366
rect 9097 1298 9155 1332
rect 9097 1264 9109 1298
rect 9143 1264 9155 1298
rect 9097 1230 9155 1264
rect 9097 1196 9109 1230
rect 9143 1196 9155 1230
rect 9097 1162 9155 1196
rect 9097 1128 9109 1162
rect 9143 1128 9155 1162
rect 9097 1004 9155 1128
rect 9185 1366 9243 1404
rect 9185 1332 9197 1366
rect 9231 1332 9243 1366
rect 9185 1298 9243 1332
rect 9185 1264 9197 1298
rect 9231 1264 9243 1298
rect 9185 1230 9243 1264
rect 9185 1196 9197 1230
rect 9231 1196 9243 1230
rect 9185 1162 9243 1196
rect 9185 1128 9197 1162
rect 9231 1128 9243 1162
rect 9185 1093 9243 1128
rect 9185 1059 9197 1093
rect 9231 1059 9243 1093
rect 9185 1004 9243 1059
rect 9273 1366 9331 1404
rect 9273 1332 9285 1366
rect 9319 1332 9331 1366
rect 9273 1298 9331 1332
rect 9273 1264 9285 1298
rect 9319 1264 9331 1298
rect 9273 1230 9331 1264
rect 9273 1196 9285 1230
rect 9319 1196 9331 1230
rect 9273 1162 9331 1196
rect 9273 1128 9285 1162
rect 9319 1128 9331 1162
rect 9273 1004 9331 1128
rect 9361 1366 9419 1404
rect 9361 1332 9373 1366
rect 9407 1332 9419 1366
rect 9361 1298 9419 1332
rect 9361 1264 9373 1298
rect 9407 1264 9419 1298
rect 9361 1230 9419 1264
rect 9361 1196 9373 1230
rect 9407 1196 9419 1230
rect 9361 1162 9419 1196
rect 9361 1128 9373 1162
rect 9407 1128 9419 1162
rect 9361 1093 9419 1128
rect 9361 1059 9373 1093
rect 9407 1059 9419 1093
rect 9361 1004 9419 1059
rect 9449 1366 9503 1404
rect 9449 1332 9461 1366
rect 9495 1332 9503 1366
rect 9449 1298 9503 1332
rect 9449 1264 9461 1298
rect 9495 1264 9503 1298
rect 9449 1230 9503 1264
rect 9449 1196 9461 1230
rect 9495 1196 9503 1230
rect 9449 1162 9503 1196
rect 9449 1128 9461 1162
rect 9495 1128 9503 1162
rect 9449 1004 9503 1128
rect 9825 1366 9881 1404
rect 9825 1332 9835 1366
rect 9869 1332 9881 1366
rect 9825 1298 9881 1332
rect 9825 1264 9835 1298
rect 9869 1264 9881 1298
rect 9825 1230 9881 1264
rect 9825 1196 9835 1230
rect 9869 1196 9881 1230
rect 9825 1162 9881 1196
rect 9825 1128 9835 1162
rect 9869 1128 9881 1162
rect 9825 1093 9881 1128
rect 9825 1059 9835 1093
rect 9869 1059 9881 1093
rect 9825 1004 9881 1059
rect 9911 1366 9969 1404
rect 9911 1332 9923 1366
rect 9957 1332 9969 1366
rect 9911 1298 9969 1332
rect 9911 1264 9923 1298
rect 9957 1264 9969 1298
rect 9911 1230 9969 1264
rect 9911 1196 9923 1230
rect 9957 1196 9969 1230
rect 9911 1162 9969 1196
rect 9911 1128 9923 1162
rect 9957 1128 9969 1162
rect 9911 1093 9969 1128
rect 9911 1059 9923 1093
rect 9957 1059 9969 1093
rect 9911 1004 9969 1059
rect 9999 1366 10057 1404
rect 9999 1332 10011 1366
rect 10045 1332 10057 1366
rect 9999 1298 10057 1332
rect 9999 1264 10011 1298
rect 10045 1264 10057 1298
rect 9999 1230 10057 1264
rect 9999 1196 10011 1230
rect 10045 1196 10057 1230
rect 9999 1162 10057 1196
rect 9999 1128 10011 1162
rect 10045 1128 10057 1162
rect 9999 1004 10057 1128
rect 10087 1366 10145 1404
rect 10087 1332 10099 1366
rect 10133 1332 10145 1366
rect 10087 1298 10145 1332
rect 10087 1264 10099 1298
rect 10133 1264 10145 1298
rect 10087 1230 10145 1264
rect 10087 1196 10099 1230
rect 10133 1196 10145 1230
rect 10087 1162 10145 1196
rect 10087 1128 10099 1162
rect 10133 1128 10145 1162
rect 10087 1093 10145 1128
rect 10087 1059 10099 1093
rect 10133 1059 10145 1093
rect 10087 1004 10145 1059
rect 10175 1366 10229 1404
rect 10175 1332 10187 1366
rect 10221 1332 10229 1366
rect 10175 1298 10229 1332
rect 10175 1264 10187 1298
rect 10221 1264 10229 1298
rect 10175 1230 10229 1264
rect 10175 1196 10187 1230
rect 10221 1196 10229 1230
rect 10175 1162 10229 1196
rect 10175 1128 10187 1162
rect 10221 1128 10229 1162
rect 10175 1004 10229 1128
rect 10551 1366 10607 1404
rect 10551 1332 10561 1366
rect 10595 1332 10607 1366
rect 10551 1298 10607 1332
rect 10551 1264 10561 1298
rect 10595 1264 10607 1298
rect 10551 1230 10607 1264
rect 10551 1196 10561 1230
rect 10595 1196 10607 1230
rect 10551 1162 10607 1196
rect 10551 1128 10561 1162
rect 10595 1128 10607 1162
rect 10551 1093 10607 1128
rect 10551 1059 10561 1093
rect 10595 1059 10607 1093
rect 10551 1004 10607 1059
rect 10637 1366 10695 1404
rect 10637 1332 10649 1366
rect 10683 1332 10695 1366
rect 10637 1298 10695 1332
rect 10637 1264 10649 1298
rect 10683 1264 10695 1298
rect 10637 1230 10695 1264
rect 10637 1196 10649 1230
rect 10683 1196 10695 1230
rect 10637 1162 10695 1196
rect 10637 1128 10649 1162
rect 10683 1128 10695 1162
rect 10637 1093 10695 1128
rect 10637 1059 10649 1093
rect 10683 1059 10695 1093
rect 10637 1004 10695 1059
rect 10725 1366 10783 1404
rect 10725 1332 10737 1366
rect 10771 1332 10783 1366
rect 10725 1298 10783 1332
rect 10725 1264 10737 1298
rect 10771 1264 10783 1298
rect 10725 1230 10783 1264
rect 10725 1196 10737 1230
rect 10771 1196 10783 1230
rect 10725 1162 10783 1196
rect 10725 1128 10737 1162
rect 10771 1128 10783 1162
rect 10725 1004 10783 1128
rect 10813 1366 10871 1404
rect 10813 1332 10825 1366
rect 10859 1332 10871 1366
rect 10813 1298 10871 1332
rect 10813 1264 10825 1298
rect 10859 1264 10871 1298
rect 10813 1230 10871 1264
rect 10813 1196 10825 1230
rect 10859 1196 10871 1230
rect 10813 1162 10871 1196
rect 10813 1128 10825 1162
rect 10859 1128 10871 1162
rect 10813 1093 10871 1128
rect 10813 1059 10825 1093
rect 10859 1059 10871 1093
rect 10813 1004 10871 1059
rect 10901 1366 10959 1404
rect 10901 1332 10913 1366
rect 10947 1332 10959 1366
rect 10901 1298 10959 1332
rect 10901 1264 10913 1298
rect 10947 1264 10959 1298
rect 10901 1230 10959 1264
rect 10901 1196 10913 1230
rect 10947 1196 10959 1230
rect 10901 1162 10959 1196
rect 10901 1128 10913 1162
rect 10947 1128 10959 1162
rect 10901 1004 10959 1128
rect 10989 1366 11047 1404
rect 10989 1332 11001 1366
rect 11035 1332 11047 1366
rect 10989 1298 11047 1332
rect 10989 1264 11001 1298
rect 11035 1264 11047 1298
rect 10989 1230 11047 1264
rect 10989 1196 11001 1230
rect 11035 1196 11047 1230
rect 10989 1162 11047 1196
rect 10989 1128 11001 1162
rect 11035 1128 11047 1162
rect 10989 1093 11047 1128
rect 10989 1059 11001 1093
rect 11035 1059 11047 1093
rect 10989 1004 11047 1059
rect 11077 1366 11131 1404
rect 11077 1332 11089 1366
rect 11123 1332 11131 1366
rect 11077 1298 11131 1332
rect 11077 1264 11089 1298
rect 11123 1264 11131 1298
rect 11077 1230 11131 1264
rect 11077 1196 11089 1230
rect 11123 1196 11131 1230
rect 11077 1162 11131 1196
rect 11077 1128 11089 1162
rect 11123 1128 11131 1162
rect 11077 1004 11131 1128
rect 11513 1366 11569 1404
rect 11513 1332 11523 1366
rect 11557 1332 11569 1366
rect 11513 1298 11569 1332
rect 11513 1264 11523 1298
rect 11557 1264 11569 1298
rect 11513 1230 11569 1264
rect 11513 1196 11523 1230
rect 11557 1196 11569 1230
rect 11513 1162 11569 1196
rect 11513 1128 11523 1162
rect 11557 1128 11569 1162
rect 11513 1093 11569 1128
rect 11513 1059 11523 1093
rect 11557 1059 11569 1093
rect 11513 1004 11569 1059
rect 11599 1366 11657 1404
rect 11599 1332 11611 1366
rect 11645 1332 11657 1366
rect 11599 1298 11657 1332
rect 11599 1264 11611 1298
rect 11645 1264 11657 1298
rect 11599 1230 11657 1264
rect 11599 1196 11611 1230
rect 11645 1196 11657 1230
rect 11599 1162 11657 1196
rect 11599 1128 11611 1162
rect 11645 1128 11657 1162
rect 11599 1093 11657 1128
rect 11599 1059 11611 1093
rect 11645 1059 11657 1093
rect 11599 1004 11657 1059
rect 11687 1366 11745 1404
rect 11687 1332 11699 1366
rect 11733 1332 11745 1366
rect 11687 1298 11745 1332
rect 11687 1264 11699 1298
rect 11733 1264 11745 1298
rect 11687 1230 11745 1264
rect 11687 1196 11699 1230
rect 11733 1196 11745 1230
rect 11687 1162 11745 1196
rect 11687 1128 11699 1162
rect 11733 1128 11745 1162
rect 11687 1004 11745 1128
rect 11775 1366 11833 1404
rect 11775 1332 11787 1366
rect 11821 1332 11833 1366
rect 11775 1298 11833 1332
rect 11775 1264 11787 1298
rect 11821 1264 11833 1298
rect 11775 1230 11833 1264
rect 11775 1196 11787 1230
rect 11821 1196 11833 1230
rect 11775 1162 11833 1196
rect 11775 1128 11787 1162
rect 11821 1128 11833 1162
rect 11775 1093 11833 1128
rect 11775 1059 11787 1093
rect 11821 1059 11833 1093
rect 11775 1004 11833 1059
rect 11863 1366 11921 1404
rect 11863 1332 11875 1366
rect 11909 1332 11921 1366
rect 11863 1298 11921 1332
rect 11863 1264 11875 1298
rect 11909 1264 11921 1298
rect 11863 1230 11921 1264
rect 11863 1196 11875 1230
rect 11909 1196 11921 1230
rect 11863 1162 11921 1196
rect 11863 1128 11875 1162
rect 11909 1128 11921 1162
rect 11863 1004 11921 1128
rect 11951 1366 12009 1404
rect 11951 1332 11963 1366
rect 11997 1332 12009 1366
rect 11951 1298 12009 1332
rect 11951 1264 11963 1298
rect 11997 1264 12009 1298
rect 11951 1230 12009 1264
rect 11951 1196 11963 1230
rect 11997 1196 12009 1230
rect 11951 1162 12009 1196
rect 11951 1128 11963 1162
rect 11997 1128 12009 1162
rect 11951 1093 12009 1128
rect 11951 1059 11963 1093
rect 11997 1059 12009 1093
rect 11951 1004 12009 1059
rect 12039 1366 12093 1404
rect 12039 1332 12051 1366
rect 12085 1332 12093 1366
rect 12039 1298 12093 1332
rect 12039 1264 12051 1298
rect 12085 1264 12093 1298
rect 12039 1230 12093 1264
rect 12039 1196 12051 1230
rect 12085 1196 12093 1230
rect 12039 1162 12093 1196
rect 12039 1128 12051 1162
rect 12085 1128 12093 1162
rect 12039 1004 12093 1128
rect 12415 1366 12471 1404
rect 12415 1332 12425 1366
rect 12459 1332 12471 1366
rect 12415 1298 12471 1332
rect 12415 1264 12425 1298
rect 12459 1264 12471 1298
rect 12415 1230 12471 1264
rect 12415 1196 12425 1230
rect 12459 1196 12471 1230
rect 12415 1162 12471 1196
rect 12415 1128 12425 1162
rect 12459 1128 12471 1162
rect 12415 1093 12471 1128
rect 12415 1059 12425 1093
rect 12459 1059 12471 1093
rect 12415 1004 12471 1059
rect 12501 1366 12559 1404
rect 12501 1332 12513 1366
rect 12547 1332 12559 1366
rect 12501 1298 12559 1332
rect 12501 1264 12513 1298
rect 12547 1264 12559 1298
rect 12501 1230 12559 1264
rect 12501 1196 12513 1230
rect 12547 1196 12559 1230
rect 12501 1162 12559 1196
rect 12501 1128 12513 1162
rect 12547 1128 12559 1162
rect 12501 1093 12559 1128
rect 12501 1059 12513 1093
rect 12547 1059 12559 1093
rect 12501 1004 12559 1059
rect 12589 1366 12647 1404
rect 12589 1332 12601 1366
rect 12635 1332 12647 1366
rect 12589 1298 12647 1332
rect 12589 1264 12601 1298
rect 12635 1264 12647 1298
rect 12589 1230 12647 1264
rect 12589 1196 12601 1230
rect 12635 1196 12647 1230
rect 12589 1162 12647 1196
rect 12589 1128 12601 1162
rect 12635 1128 12647 1162
rect 12589 1004 12647 1128
rect 12677 1366 12735 1404
rect 12677 1332 12689 1366
rect 12723 1332 12735 1366
rect 12677 1298 12735 1332
rect 12677 1264 12689 1298
rect 12723 1264 12735 1298
rect 12677 1230 12735 1264
rect 12677 1196 12689 1230
rect 12723 1196 12735 1230
rect 12677 1162 12735 1196
rect 12677 1128 12689 1162
rect 12723 1128 12735 1162
rect 12677 1093 12735 1128
rect 12677 1059 12689 1093
rect 12723 1059 12735 1093
rect 12677 1004 12735 1059
rect 12765 1366 12819 1404
rect 12765 1332 12777 1366
rect 12811 1332 12819 1366
rect 12765 1298 12819 1332
rect 12765 1264 12777 1298
rect 12811 1264 12819 1298
rect 12765 1230 12819 1264
rect 12765 1196 12777 1230
rect 12811 1196 12819 1230
rect 12765 1162 12819 1196
rect 12765 1128 12777 1162
rect 12811 1128 12819 1162
rect 12765 1004 12819 1128
rect 13141 1366 13197 1404
rect 13141 1332 13151 1366
rect 13185 1332 13197 1366
rect 13141 1298 13197 1332
rect 13141 1264 13151 1298
rect 13185 1264 13197 1298
rect 13141 1230 13197 1264
rect 13141 1196 13151 1230
rect 13185 1196 13197 1230
rect 13141 1162 13197 1196
rect 13141 1128 13151 1162
rect 13185 1128 13197 1162
rect 13141 1093 13197 1128
rect 13141 1059 13151 1093
rect 13185 1059 13197 1093
rect 13141 1004 13197 1059
rect 13227 1366 13285 1404
rect 13227 1332 13239 1366
rect 13273 1332 13285 1366
rect 13227 1298 13285 1332
rect 13227 1264 13239 1298
rect 13273 1264 13285 1298
rect 13227 1230 13285 1264
rect 13227 1196 13239 1230
rect 13273 1196 13285 1230
rect 13227 1162 13285 1196
rect 13227 1128 13239 1162
rect 13273 1128 13285 1162
rect 13227 1093 13285 1128
rect 13227 1059 13239 1093
rect 13273 1059 13285 1093
rect 13227 1004 13285 1059
rect 13315 1366 13373 1404
rect 13315 1332 13327 1366
rect 13361 1332 13373 1366
rect 13315 1298 13373 1332
rect 13315 1264 13327 1298
rect 13361 1264 13373 1298
rect 13315 1230 13373 1264
rect 13315 1196 13327 1230
rect 13361 1196 13373 1230
rect 13315 1162 13373 1196
rect 13315 1128 13327 1162
rect 13361 1128 13373 1162
rect 13315 1004 13373 1128
rect 13403 1366 13461 1404
rect 13403 1332 13415 1366
rect 13449 1332 13461 1366
rect 13403 1298 13461 1332
rect 13403 1264 13415 1298
rect 13449 1264 13461 1298
rect 13403 1230 13461 1264
rect 13403 1196 13415 1230
rect 13449 1196 13461 1230
rect 13403 1162 13461 1196
rect 13403 1128 13415 1162
rect 13449 1128 13461 1162
rect 13403 1093 13461 1128
rect 13403 1059 13415 1093
rect 13449 1059 13461 1093
rect 13403 1004 13461 1059
rect 13491 1366 13549 1404
rect 13491 1332 13503 1366
rect 13537 1332 13549 1366
rect 13491 1298 13549 1332
rect 13491 1264 13503 1298
rect 13537 1264 13549 1298
rect 13491 1230 13549 1264
rect 13491 1196 13503 1230
rect 13537 1196 13549 1230
rect 13491 1162 13549 1196
rect 13491 1128 13503 1162
rect 13537 1128 13549 1162
rect 13491 1004 13549 1128
rect 13579 1366 13637 1404
rect 13579 1332 13591 1366
rect 13625 1332 13637 1366
rect 13579 1298 13637 1332
rect 13579 1264 13591 1298
rect 13625 1264 13637 1298
rect 13579 1230 13637 1264
rect 13579 1196 13591 1230
rect 13625 1196 13637 1230
rect 13579 1162 13637 1196
rect 13579 1128 13591 1162
rect 13625 1128 13637 1162
rect 13579 1093 13637 1128
rect 13579 1059 13591 1093
rect 13625 1059 13637 1093
rect 13579 1004 13637 1059
rect 13667 1366 13721 1404
rect 13667 1332 13679 1366
rect 13713 1332 13721 1366
rect 13667 1298 13721 1332
rect 13667 1264 13679 1298
rect 13713 1264 13721 1298
rect 13667 1230 13721 1264
rect 13667 1196 13679 1230
rect 13713 1196 13721 1230
rect 13667 1162 13721 1196
rect 13667 1128 13679 1162
rect 13713 1128 13721 1162
rect 13667 1004 13721 1128
rect 14103 1366 14159 1404
rect 14103 1332 14113 1366
rect 14147 1332 14159 1366
rect 14103 1298 14159 1332
rect 14103 1264 14113 1298
rect 14147 1264 14159 1298
rect 14103 1230 14159 1264
rect 14103 1196 14113 1230
rect 14147 1196 14159 1230
rect 14103 1162 14159 1196
rect 14103 1128 14113 1162
rect 14147 1128 14159 1162
rect 14103 1093 14159 1128
rect 14103 1059 14113 1093
rect 14147 1059 14159 1093
rect 14103 1004 14159 1059
rect 14189 1366 14247 1404
rect 14189 1332 14201 1366
rect 14235 1332 14247 1366
rect 14189 1298 14247 1332
rect 14189 1264 14201 1298
rect 14235 1264 14247 1298
rect 14189 1230 14247 1264
rect 14189 1196 14201 1230
rect 14235 1196 14247 1230
rect 14189 1162 14247 1196
rect 14189 1128 14201 1162
rect 14235 1128 14247 1162
rect 14189 1093 14247 1128
rect 14189 1059 14201 1093
rect 14235 1059 14247 1093
rect 14189 1004 14247 1059
rect 14277 1366 14335 1404
rect 14277 1332 14289 1366
rect 14323 1332 14335 1366
rect 14277 1298 14335 1332
rect 14277 1264 14289 1298
rect 14323 1264 14335 1298
rect 14277 1230 14335 1264
rect 14277 1196 14289 1230
rect 14323 1196 14335 1230
rect 14277 1162 14335 1196
rect 14277 1128 14289 1162
rect 14323 1128 14335 1162
rect 14277 1004 14335 1128
rect 14365 1366 14423 1404
rect 14365 1332 14377 1366
rect 14411 1332 14423 1366
rect 14365 1298 14423 1332
rect 14365 1264 14377 1298
rect 14411 1264 14423 1298
rect 14365 1230 14423 1264
rect 14365 1196 14377 1230
rect 14411 1196 14423 1230
rect 14365 1162 14423 1196
rect 14365 1128 14377 1162
rect 14411 1128 14423 1162
rect 14365 1093 14423 1128
rect 14365 1059 14377 1093
rect 14411 1059 14423 1093
rect 14365 1004 14423 1059
rect 14453 1366 14511 1404
rect 14453 1332 14465 1366
rect 14499 1332 14511 1366
rect 14453 1298 14511 1332
rect 14453 1264 14465 1298
rect 14499 1264 14511 1298
rect 14453 1230 14511 1264
rect 14453 1196 14465 1230
rect 14499 1196 14511 1230
rect 14453 1162 14511 1196
rect 14453 1128 14465 1162
rect 14499 1128 14511 1162
rect 14453 1004 14511 1128
rect 14541 1366 14599 1404
rect 14541 1332 14553 1366
rect 14587 1332 14599 1366
rect 14541 1298 14599 1332
rect 14541 1264 14553 1298
rect 14587 1264 14599 1298
rect 14541 1230 14599 1264
rect 14541 1196 14553 1230
rect 14587 1196 14599 1230
rect 14541 1162 14599 1196
rect 14541 1128 14553 1162
rect 14587 1128 14599 1162
rect 14541 1093 14599 1128
rect 14541 1059 14553 1093
rect 14587 1059 14599 1093
rect 14541 1004 14599 1059
rect 14629 1366 14683 1404
rect 14629 1332 14641 1366
rect 14675 1332 14683 1366
rect 14629 1298 14683 1332
rect 14629 1264 14641 1298
rect 14675 1264 14683 1298
rect 14629 1230 14683 1264
rect 14629 1196 14641 1230
rect 14675 1196 14683 1230
rect 14629 1162 14683 1196
rect 14629 1128 14641 1162
rect 14675 1128 14683 1162
rect 14629 1004 14683 1128
rect 15005 1366 15061 1404
rect 15005 1332 15015 1366
rect 15049 1332 15061 1366
rect 15005 1298 15061 1332
rect 15005 1264 15015 1298
rect 15049 1264 15061 1298
rect 15005 1230 15061 1264
rect 15005 1196 15015 1230
rect 15049 1196 15061 1230
rect 15005 1162 15061 1196
rect 15005 1128 15015 1162
rect 15049 1128 15061 1162
rect 15005 1093 15061 1128
rect 15005 1059 15015 1093
rect 15049 1059 15061 1093
rect 15005 1004 15061 1059
rect 15091 1366 15149 1404
rect 15091 1332 15103 1366
rect 15137 1332 15149 1366
rect 15091 1298 15149 1332
rect 15091 1264 15103 1298
rect 15137 1264 15149 1298
rect 15091 1230 15149 1264
rect 15091 1196 15103 1230
rect 15137 1196 15149 1230
rect 15091 1162 15149 1196
rect 15091 1128 15103 1162
rect 15137 1128 15149 1162
rect 15091 1093 15149 1128
rect 15091 1059 15103 1093
rect 15137 1059 15149 1093
rect 15091 1004 15149 1059
rect 15179 1366 15237 1404
rect 15179 1332 15191 1366
rect 15225 1332 15237 1366
rect 15179 1298 15237 1332
rect 15179 1264 15191 1298
rect 15225 1264 15237 1298
rect 15179 1230 15237 1264
rect 15179 1196 15191 1230
rect 15225 1196 15237 1230
rect 15179 1162 15237 1196
rect 15179 1128 15191 1162
rect 15225 1128 15237 1162
rect 15179 1004 15237 1128
rect 15267 1366 15325 1404
rect 15267 1332 15279 1366
rect 15313 1332 15325 1366
rect 15267 1298 15325 1332
rect 15267 1264 15279 1298
rect 15313 1264 15325 1298
rect 15267 1230 15325 1264
rect 15267 1196 15279 1230
rect 15313 1196 15325 1230
rect 15267 1162 15325 1196
rect 15267 1128 15279 1162
rect 15313 1128 15325 1162
rect 15267 1093 15325 1128
rect 15267 1059 15279 1093
rect 15313 1059 15325 1093
rect 15267 1004 15325 1059
rect 15355 1366 15409 1404
rect 15355 1332 15367 1366
rect 15401 1332 15409 1366
rect 15355 1298 15409 1332
rect 15355 1264 15367 1298
rect 15401 1264 15409 1298
rect 15355 1230 15409 1264
rect 15355 1196 15367 1230
rect 15401 1196 15409 1230
rect 15355 1162 15409 1196
rect 15355 1128 15367 1162
rect 15401 1128 15409 1162
rect 15355 1004 15409 1128
rect 15671 1365 15727 1405
rect 15671 1331 15681 1365
rect 15715 1331 15727 1365
rect 15671 1297 15727 1331
rect 15671 1263 15681 1297
rect 15715 1263 15727 1297
rect 15671 1229 15727 1263
rect 15671 1195 15681 1229
rect 15715 1195 15727 1229
rect 15671 1161 15727 1195
rect 15671 1127 15681 1161
rect 15715 1127 15727 1161
rect 15671 1093 15727 1127
rect 15671 1059 15681 1093
rect 15715 1059 15727 1093
rect 15671 1005 15727 1059
rect 15757 1365 15815 1405
rect 15757 1331 15769 1365
rect 15803 1331 15815 1365
rect 15757 1297 15815 1331
rect 15757 1263 15769 1297
rect 15803 1263 15815 1297
rect 15757 1229 15815 1263
rect 15757 1195 15769 1229
rect 15803 1195 15815 1229
rect 15757 1161 15815 1195
rect 15757 1127 15769 1161
rect 15803 1127 15815 1161
rect 15757 1093 15815 1127
rect 15757 1059 15769 1093
rect 15803 1059 15815 1093
rect 15757 1005 15815 1059
rect 15845 1365 15903 1405
rect 15845 1331 15857 1365
rect 15891 1331 15903 1365
rect 15845 1297 15903 1331
rect 15845 1263 15857 1297
rect 15891 1263 15903 1297
rect 15845 1229 15903 1263
rect 15845 1195 15857 1229
rect 15891 1195 15903 1229
rect 15845 1161 15903 1195
rect 15845 1127 15857 1161
rect 15891 1127 15903 1161
rect 15845 1005 15903 1127
rect 15933 1365 15991 1405
rect 15933 1331 15945 1365
rect 15979 1331 15991 1365
rect 15933 1297 15991 1331
rect 15933 1263 15945 1297
rect 15979 1263 15991 1297
rect 15933 1229 15991 1263
rect 15933 1195 15945 1229
rect 15979 1195 15991 1229
rect 15933 1161 15991 1195
rect 15933 1127 15945 1161
rect 15979 1127 15991 1161
rect 15933 1005 15991 1127
rect 16021 1365 16075 1405
rect 16021 1331 16033 1365
rect 16067 1331 16075 1365
rect 16021 1297 16075 1331
rect 16021 1263 16033 1297
rect 16067 1263 16075 1297
rect 16021 1229 16075 1263
rect 16021 1195 16033 1229
rect 16067 1195 16075 1229
rect 16021 1161 16075 1195
rect 16021 1127 16033 1161
rect 16067 1127 16075 1161
rect 16021 1093 16075 1127
rect 16021 1059 16033 1093
rect 16067 1059 16075 1093
rect 16021 1005 16075 1059
rect 16337 1365 16391 1405
rect 16337 1331 16345 1365
rect 16379 1331 16391 1365
rect 16337 1297 16391 1331
rect 16337 1263 16345 1297
rect 16379 1263 16391 1297
rect 16337 1229 16391 1263
rect 16337 1195 16345 1229
rect 16379 1195 16391 1229
rect 16337 1161 16391 1195
rect 16337 1127 16345 1161
rect 16379 1127 16391 1161
rect 16337 1005 16391 1127
rect 16421 1297 16479 1405
rect 16421 1263 16433 1297
rect 16467 1263 16479 1297
rect 16421 1229 16479 1263
rect 16421 1195 16433 1229
rect 16467 1195 16479 1229
rect 16421 1161 16479 1195
rect 16421 1127 16433 1161
rect 16467 1127 16479 1161
rect 16421 1093 16479 1127
rect 16421 1059 16433 1093
rect 16467 1059 16479 1093
rect 16421 1005 16479 1059
rect 16509 1365 16567 1405
rect 16509 1331 16521 1365
rect 16555 1331 16567 1365
rect 16509 1297 16567 1331
rect 16509 1263 16521 1297
rect 16555 1263 16567 1297
rect 16509 1229 16567 1263
rect 16509 1195 16521 1229
rect 16555 1195 16567 1229
rect 16509 1161 16567 1195
rect 16509 1127 16521 1161
rect 16555 1127 16567 1161
rect 16509 1005 16567 1127
rect 16597 1297 16655 1405
rect 16597 1263 16609 1297
rect 16643 1263 16655 1297
rect 16597 1229 16655 1263
rect 16597 1195 16609 1229
rect 16643 1195 16655 1229
rect 16597 1161 16655 1195
rect 16597 1127 16609 1161
rect 16643 1127 16655 1161
rect 16597 1005 16655 1127
rect 16685 1365 16741 1405
rect 16685 1331 16697 1365
rect 16731 1331 16741 1365
rect 16685 1297 16741 1331
rect 16685 1263 16697 1297
rect 16731 1263 16741 1297
rect 16685 1229 16741 1263
rect 16685 1195 16697 1229
rect 16731 1195 16741 1229
rect 16685 1161 16741 1195
rect 16685 1127 16697 1161
rect 16731 1127 16741 1161
rect 16685 1005 16741 1127
rect 17003 1365 17059 1405
rect 17003 1331 17013 1365
rect 17047 1331 17059 1365
rect 17003 1297 17059 1331
rect 17003 1263 17013 1297
rect 17047 1263 17059 1297
rect 17003 1229 17059 1263
rect 17003 1195 17013 1229
rect 17047 1195 17059 1229
rect 17003 1161 17059 1195
rect 17003 1127 17013 1161
rect 17047 1127 17059 1161
rect 17003 1005 17059 1127
rect 17089 1297 17147 1405
rect 17089 1263 17101 1297
rect 17135 1263 17147 1297
rect 17089 1229 17147 1263
rect 17089 1195 17101 1229
rect 17135 1195 17147 1229
rect 17089 1161 17147 1195
rect 17089 1127 17101 1161
rect 17135 1127 17147 1161
rect 17089 1093 17147 1127
rect 17089 1059 17101 1093
rect 17135 1059 17147 1093
rect 17089 1005 17147 1059
rect 17177 1365 17235 1405
rect 17177 1331 17189 1365
rect 17223 1331 17235 1365
rect 17177 1297 17235 1331
rect 17177 1263 17189 1297
rect 17223 1263 17235 1297
rect 17177 1229 17235 1263
rect 17177 1195 17189 1229
rect 17223 1195 17235 1229
rect 17177 1161 17235 1195
rect 17177 1127 17189 1161
rect 17223 1127 17235 1161
rect 17177 1005 17235 1127
rect 17265 1297 17323 1405
rect 17265 1263 17277 1297
rect 17311 1263 17323 1297
rect 17265 1229 17323 1263
rect 17265 1195 17277 1229
rect 17311 1195 17323 1229
rect 17265 1161 17323 1195
rect 17265 1127 17277 1161
rect 17311 1127 17323 1161
rect 17265 1093 17323 1127
rect 17265 1059 17277 1093
rect 17311 1059 17323 1093
rect 17265 1005 17323 1059
rect 17353 1365 17407 1405
rect 17353 1331 17365 1365
rect 17399 1331 17407 1365
rect 17353 1297 17407 1331
rect 17353 1263 17365 1297
rect 17399 1263 17407 1297
rect 17353 1229 17407 1263
rect 17353 1195 17365 1229
rect 17399 1195 17407 1229
rect 17353 1161 17407 1195
rect 17353 1127 17365 1161
rect 17399 1127 17407 1161
rect 17353 1005 17407 1127
rect 17646 1366 17702 1404
rect 17646 1332 17656 1366
rect 17690 1332 17702 1366
rect 17646 1298 17702 1332
rect 17646 1264 17656 1298
rect 17690 1264 17702 1298
rect 17646 1230 17702 1264
rect 17646 1196 17656 1230
rect 17690 1196 17702 1230
rect 17646 1162 17702 1196
rect 17646 1128 17656 1162
rect 17690 1128 17702 1162
rect 17646 1093 17702 1128
rect 17646 1059 17656 1093
rect 17690 1059 17702 1093
rect 17646 1004 17702 1059
rect 17732 1366 17790 1404
rect 17732 1332 17744 1366
rect 17778 1332 17790 1366
rect 17732 1298 17790 1332
rect 17732 1264 17744 1298
rect 17778 1264 17790 1298
rect 17732 1230 17790 1264
rect 17732 1196 17744 1230
rect 17778 1196 17790 1230
rect 17732 1162 17790 1196
rect 17732 1128 17744 1162
rect 17778 1128 17790 1162
rect 17732 1093 17790 1128
rect 17732 1059 17744 1093
rect 17778 1059 17790 1093
rect 17732 1004 17790 1059
rect 17820 1366 17874 1404
rect 17820 1332 17832 1366
rect 17866 1332 17874 1366
rect 17820 1298 17874 1332
rect 17820 1264 17832 1298
rect 17866 1264 17874 1298
rect 17820 1230 17874 1264
rect 17820 1196 17832 1230
rect 17866 1196 17874 1230
rect 17820 1162 17874 1196
rect 17820 1128 17832 1162
rect 17866 1128 17874 1162
rect 17820 1093 17874 1128
rect 17820 1059 17832 1093
rect 17866 1059 17874 1093
rect 17820 1004 17874 1059
<< ndiffc >>
rect 101 301 135 335
rect 198 301 232 335
rect 295 301 329 335
rect 392 301 426 335
rect 489 301 523 335
rect 101 229 135 263
rect 101 161 135 195
rect 198 176 232 210
rect 295 229 329 263
rect 295 161 329 195
rect 393 182 427 216
rect 101 91 135 125
rect 295 91 329 125
rect 392 91 426 125
rect 489 91 523 125
rect 603 301 637 335
rect 603 229 637 263
rect 603 161 637 195
rect 700 185 734 219
rect 797 229 831 263
rect 797 161 831 195
rect 603 91 637 125
rect 700 91 734 125
rect 797 91 831 125
rect 1063 301 1097 335
rect 1160 301 1194 335
rect 1257 301 1291 335
rect 1354 301 1388 335
rect 1451 301 1485 335
rect 1063 229 1097 263
rect 1063 161 1097 195
rect 1160 176 1194 210
rect 1257 229 1291 263
rect 1257 161 1291 195
rect 1355 182 1389 216
rect 1063 91 1097 125
rect 1257 91 1291 125
rect 1354 91 1388 125
rect 1451 91 1485 125
rect 1565 301 1599 335
rect 1565 229 1599 263
rect 1565 161 1599 195
rect 1662 185 1696 219
rect 1759 229 1793 263
rect 1759 161 1793 195
rect 1565 91 1599 125
rect 1662 91 1696 125
rect 1759 91 1793 125
rect 2046 299 2080 333
rect 2143 299 2177 333
rect 2240 299 2274 333
rect 2046 227 2080 261
rect 2046 159 2080 193
rect 2143 174 2177 208
rect 2240 227 2274 261
rect 2240 159 2274 193
rect 2337 183 2371 217
rect 2434 227 2468 261
rect 2434 159 2468 193
rect 2046 89 2080 123
rect 2240 89 2274 123
rect 2337 89 2371 123
rect 2434 89 2468 123
rect 2691 301 2725 335
rect 2788 301 2822 335
rect 2885 301 2919 335
rect 2982 301 3016 335
rect 3079 301 3113 335
rect 2691 229 2725 263
rect 2691 161 2725 195
rect 2788 176 2822 210
rect 2885 229 2919 263
rect 2885 161 2919 195
rect 2983 182 3017 216
rect 2691 91 2725 125
rect 2885 91 2919 125
rect 2982 91 3016 125
rect 3079 91 3113 125
rect 3193 301 3227 335
rect 3193 229 3227 263
rect 3193 161 3227 195
rect 3290 185 3324 219
rect 3387 229 3421 263
rect 3387 161 3421 195
rect 3193 91 3227 125
rect 3290 91 3324 125
rect 3387 91 3421 125
rect 3653 301 3687 335
rect 3750 301 3784 335
rect 3847 301 3881 335
rect 3944 301 3978 335
rect 4041 301 4075 335
rect 3653 229 3687 263
rect 3653 161 3687 195
rect 3750 176 3784 210
rect 3847 229 3881 263
rect 3847 161 3881 195
rect 3945 182 3979 216
rect 3653 91 3687 125
rect 3847 91 3881 125
rect 3944 91 3978 125
rect 4041 91 4075 125
rect 4155 301 4189 335
rect 4155 229 4189 263
rect 4155 161 4189 195
rect 4252 185 4286 219
rect 4349 229 4383 263
rect 4349 161 4383 195
rect 4155 91 4189 125
rect 4252 91 4286 125
rect 4349 91 4383 125
rect 4636 299 4670 333
rect 4733 299 4767 333
rect 4830 299 4864 333
rect 4636 227 4670 261
rect 4636 159 4670 193
rect 4733 174 4767 208
rect 4830 227 4864 261
rect 4830 159 4864 193
rect 4927 183 4961 217
rect 5024 227 5058 261
rect 5024 159 5058 193
rect 4636 89 4670 123
rect 4830 89 4864 123
rect 4927 89 4961 123
rect 5024 89 5058 123
rect 5281 301 5315 335
rect 5378 301 5412 335
rect 5475 301 5509 335
rect 5572 301 5606 335
rect 5669 301 5703 335
rect 5281 229 5315 263
rect 5281 161 5315 195
rect 5378 176 5412 210
rect 5475 229 5509 263
rect 5475 161 5509 195
rect 5573 182 5607 216
rect 5281 91 5315 125
rect 5475 91 5509 125
rect 5572 91 5606 125
rect 5669 91 5703 125
rect 5783 301 5817 335
rect 5783 229 5817 263
rect 5783 161 5817 195
rect 5880 185 5914 219
rect 5977 229 6011 263
rect 5977 161 6011 195
rect 5783 91 5817 125
rect 5880 91 5914 125
rect 5977 91 6011 125
rect 6243 301 6277 335
rect 6340 301 6374 335
rect 6437 301 6471 335
rect 6534 301 6568 335
rect 6631 301 6665 335
rect 6243 229 6277 263
rect 6243 161 6277 195
rect 6340 176 6374 210
rect 6437 229 6471 263
rect 6437 161 6471 195
rect 6535 182 6569 216
rect 6243 91 6277 125
rect 6437 91 6471 125
rect 6534 91 6568 125
rect 6631 91 6665 125
rect 6745 301 6779 335
rect 6745 229 6779 263
rect 6745 161 6779 195
rect 6842 185 6876 219
rect 6939 229 6973 263
rect 6939 161 6973 195
rect 6745 91 6779 125
rect 6842 91 6876 125
rect 6939 91 6973 125
rect 7226 299 7260 333
rect 7323 299 7357 333
rect 7420 299 7454 333
rect 7226 227 7260 261
rect 7226 159 7260 193
rect 7323 174 7357 208
rect 7420 227 7454 261
rect 7420 159 7454 193
rect 7517 183 7551 217
rect 7614 227 7648 261
rect 7614 159 7648 193
rect 7226 89 7260 123
rect 7420 89 7454 123
rect 7517 89 7551 123
rect 7614 89 7648 123
rect 7871 301 7905 335
rect 7968 301 8002 335
rect 8065 301 8099 335
rect 8162 301 8196 335
rect 8259 301 8293 335
rect 7871 229 7905 263
rect 7871 161 7905 195
rect 7968 176 8002 210
rect 8065 229 8099 263
rect 8065 161 8099 195
rect 8163 182 8197 216
rect 7871 91 7905 125
rect 8065 91 8099 125
rect 8162 91 8196 125
rect 8259 91 8293 125
rect 8373 301 8407 335
rect 8373 229 8407 263
rect 8373 161 8407 195
rect 8470 185 8504 219
rect 8567 229 8601 263
rect 8567 161 8601 195
rect 8373 91 8407 125
rect 8470 91 8504 125
rect 8567 91 8601 125
rect 8833 301 8867 335
rect 8930 301 8964 335
rect 9027 301 9061 335
rect 9124 301 9158 335
rect 9221 301 9255 335
rect 8833 229 8867 263
rect 8833 161 8867 195
rect 8930 176 8964 210
rect 9027 229 9061 263
rect 9027 161 9061 195
rect 9125 182 9159 216
rect 8833 91 8867 125
rect 9027 91 9061 125
rect 9124 91 9158 125
rect 9221 91 9255 125
rect 9335 301 9369 335
rect 9335 229 9369 263
rect 9335 161 9369 195
rect 9432 185 9466 219
rect 9529 229 9563 263
rect 9529 161 9563 195
rect 9335 91 9369 125
rect 9432 91 9466 125
rect 9529 91 9563 125
rect 9816 299 9850 333
rect 9913 299 9947 333
rect 10010 299 10044 333
rect 9816 227 9850 261
rect 9816 159 9850 193
rect 9913 174 9947 208
rect 10010 227 10044 261
rect 10010 159 10044 193
rect 10107 183 10141 217
rect 10204 227 10238 261
rect 10204 159 10238 193
rect 9816 89 9850 123
rect 10010 89 10044 123
rect 10107 89 10141 123
rect 10204 89 10238 123
rect 10461 301 10495 335
rect 10558 301 10592 335
rect 10655 301 10689 335
rect 10752 301 10786 335
rect 10849 301 10883 335
rect 10461 229 10495 263
rect 10461 161 10495 195
rect 10558 176 10592 210
rect 10655 229 10689 263
rect 10655 161 10689 195
rect 10753 182 10787 216
rect 10461 91 10495 125
rect 10655 91 10689 125
rect 10752 91 10786 125
rect 10849 91 10883 125
rect 10963 301 10997 335
rect 10963 229 10997 263
rect 10963 161 10997 195
rect 11060 185 11094 219
rect 11157 229 11191 263
rect 11157 161 11191 195
rect 10963 91 10997 125
rect 11060 91 11094 125
rect 11157 91 11191 125
rect 11423 301 11457 335
rect 11520 301 11554 335
rect 11617 301 11651 335
rect 11714 301 11748 335
rect 11811 301 11845 335
rect 11423 229 11457 263
rect 11423 161 11457 195
rect 11520 176 11554 210
rect 11617 229 11651 263
rect 11617 161 11651 195
rect 11715 182 11749 216
rect 11423 91 11457 125
rect 11617 91 11651 125
rect 11714 91 11748 125
rect 11811 91 11845 125
rect 11925 301 11959 335
rect 11925 229 11959 263
rect 11925 161 11959 195
rect 12022 185 12056 219
rect 12119 229 12153 263
rect 12119 161 12153 195
rect 11925 91 11959 125
rect 12022 91 12056 125
rect 12119 91 12153 125
rect 12406 299 12440 333
rect 12503 299 12537 333
rect 12600 299 12634 333
rect 12406 227 12440 261
rect 12406 159 12440 193
rect 12503 174 12537 208
rect 12600 227 12634 261
rect 12600 159 12634 193
rect 12697 183 12731 217
rect 12794 227 12828 261
rect 12794 159 12828 193
rect 12406 89 12440 123
rect 12600 89 12634 123
rect 12697 89 12731 123
rect 12794 89 12828 123
rect 13051 301 13085 335
rect 13148 301 13182 335
rect 13245 301 13279 335
rect 13342 301 13376 335
rect 13439 301 13473 335
rect 13051 229 13085 263
rect 13051 161 13085 195
rect 13148 176 13182 210
rect 13245 229 13279 263
rect 13245 161 13279 195
rect 13343 182 13377 216
rect 13051 91 13085 125
rect 13245 91 13279 125
rect 13342 91 13376 125
rect 13439 91 13473 125
rect 13553 301 13587 335
rect 13553 229 13587 263
rect 13553 161 13587 195
rect 13650 185 13684 219
rect 13747 229 13781 263
rect 13747 161 13781 195
rect 13553 91 13587 125
rect 13650 91 13684 125
rect 13747 91 13781 125
rect 14013 301 14047 335
rect 14110 301 14144 335
rect 14207 301 14241 335
rect 14304 301 14338 335
rect 14401 301 14435 335
rect 14013 229 14047 263
rect 14013 161 14047 195
rect 14110 176 14144 210
rect 14207 229 14241 263
rect 14207 161 14241 195
rect 14305 182 14339 216
rect 14013 91 14047 125
rect 14207 91 14241 125
rect 14304 91 14338 125
rect 14401 91 14435 125
rect 14515 301 14549 335
rect 14515 229 14549 263
rect 14515 161 14549 195
rect 14612 185 14646 219
rect 14709 229 14743 263
rect 14709 161 14743 195
rect 14515 91 14549 125
rect 14612 91 14646 125
rect 14709 91 14743 125
rect 14996 299 15030 333
rect 15093 299 15127 333
rect 15190 299 15224 333
rect 14996 227 15030 261
rect 14996 159 15030 193
rect 15093 174 15127 208
rect 15190 227 15224 261
rect 15190 159 15224 193
rect 15287 183 15321 217
rect 15384 227 15418 261
rect 15384 159 15418 193
rect 14996 89 15030 123
rect 15190 89 15224 123
rect 15287 89 15321 123
rect 15384 89 15418 123
rect 15662 299 15696 333
rect 15759 299 15793 333
rect 15856 299 15890 333
rect 16050 299 16084 333
rect 15662 227 15696 261
rect 15662 159 15696 193
rect 15759 174 15793 208
rect 15856 227 15890 261
rect 15856 159 15890 193
rect 15952 183 15986 217
rect 16050 227 16084 261
rect 16050 159 16084 193
rect 15662 89 15696 123
rect 15856 89 15890 123
rect 15952 89 15986 123
rect 16050 89 16084 123
rect 16328 299 16362 333
rect 16425 299 16459 333
rect 16522 299 16556 333
rect 16716 299 16750 333
rect 16328 227 16362 261
rect 16328 159 16362 193
rect 16425 174 16459 208
rect 16522 227 16556 261
rect 16522 159 16556 193
rect 16619 183 16653 217
rect 16716 227 16750 261
rect 16716 159 16750 193
rect 16328 89 16362 123
rect 16522 89 16556 123
rect 16619 89 16653 123
rect 16716 89 16750 123
rect 16994 299 17028 333
rect 17091 299 17125 333
rect 17188 299 17222 333
rect 16994 227 17028 261
rect 16994 159 17028 193
rect 17091 174 17125 208
rect 17188 227 17222 261
rect 17188 159 17222 193
rect 17285 183 17319 217
rect 17382 227 17416 261
rect 17382 159 17416 193
rect 16994 89 17028 123
rect 17188 89 17222 123
rect 17285 89 17319 123
rect 17382 89 17416 123
rect 17647 300 17681 334
rect 17841 300 17875 334
rect 17647 228 17681 262
rect 17647 160 17681 194
rect 17743 184 17777 218
rect 17841 228 17875 262
rect 17841 160 17875 194
rect 17647 90 17681 124
rect 17743 90 17777 124
rect 17841 90 17875 124
<< pdiffc >>
rect 201 1332 235 1366
rect 201 1264 235 1298
rect 201 1196 235 1230
rect 201 1128 235 1162
rect 201 1059 235 1093
rect 289 1332 323 1366
rect 289 1264 323 1298
rect 289 1196 323 1230
rect 289 1128 323 1162
rect 289 1059 323 1093
rect 377 1332 411 1366
rect 377 1264 411 1298
rect 377 1196 411 1230
rect 377 1128 411 1162
rect 465 1332 499 1366
rect 465 1264 499 1298
rect 465 1196 499 1230
rect 465 1128 499 1162
rect 465 1059 499 1093
rect 553 1332 587 1366
rect 553 1264 587 1298
rect 553 1196 587 1230
rect 553 1128 587 1162
rect 641 1332 675 1366
rect 641 1264 675 1298
rect 641 1196 675 1230
rect 641 1128 675 1162
rect 641 1059 675 1093
rect 729 1332 763 1366
rect 729 1264 763 1298
rect 729 1196 763 1230
rect 729 1128 763 1162
rect 1163 1332 1197 1366
rect 1163 1264 1197 1298
rect 1163 1196 1197 1230
rect 1163 1128 1197 1162
rect 1163 1059 1197 1093
rect 1251 1332 1285 1366
rect 1251 1264 1285 1298
rect 1251 1196 1285 1230
rect 1251 1128 1285 1162
rect 1251 1059 1285 1093
rect 1339 1332 1373 1366
rect 1339 1264 1373 1298
rect 1339 1196 1373 1230
rect 1339 1128 1373 1162
rect 1427 1332 1461 1366
rect 1427 1264 1461 1298
rect 1427 1196 1461 1230
rect 1427 1128 1461 1162
rect 1427 1059 1461 1093
rect 1515 1332 1549 1366
rect 1515 1264 1549 1298
rect 1515 1196 1549 1230
rect 1515 1128 1549 1162
rect 1603 1332 1637 1366
rect 1603 1264 1637 1298
rect 1603 1196 1637 1230
rect 1603 1128 1637 1162
rect 1603 1059 1637 1093
rect 1691 1332 1725 1366
rect 1691 1264 1725 1298
rect 1691 1196 1725 1230
rect 1691 1128 1725 1162
rect 2065 1332 2099 1366
rect 2065 1264 2099 1298
rect 2065 1196 2099 1230
rect 2065 1128 2099 1162
rect 2065 1059 2099 1093
rect 2153 1332 2187 1366
rect 2153 1264 2187 1298
rect 2153 1196 2187 1230
rect 2153 1128 2187 1162
rect 2153 1059 2187 1093
rect 2241 1332 2275 1366
rect 2241 1264 2275 1298
rect 2241 1196 2275 1230
rect 2241 1128 2275 1162
rect 2329 1332 2363 1366
rect 2329 1264 2363 1298
rect 2329 1196 2363 1230
rect 2329 1128 2363 1162
rect 2329 1059 2363 1093
rect 2417 1332 2451 1366
rect 2417 1264 2451 1298
rect 2417 1196 2451 1230
rect 2417 1128 2451 1162
rect 2791 1332 2825 1366
rect 2791 1264 2825 1298
rect 2791 1196 2825 1230
rect 2791 1128 2825 1162
rect 2791 1059 2825 1093
rect 2879 1332 2913 1366
rect 2879 1264 2913 1298
rect 2879 1196 2913 1230
rect 2879 1128 2913 1162
rect 2879 1059 2913 1093
rect 2967 1332 3001 1366
rect 2967 1264 3001 1298
rect 2967 1196 3001 1230
rect 2967 1128 3001 1162
rect 3055 1332 3089 1366
rect 3055 1264 3089 1298
rect 3055 1196 3089 1230
rect 3055 1128 3089 1162
rect 3055 1059 3089 1093
rect 3143 1332 3177 1366
rect 3143 1264 3177 1298
rect 3143 1196 3177 1230
rect 3143 1128 3177 1162
rect 3231 1332 3265 1366
rect 3231 1264 3265 1298
rect 3231 1196 3265 1230
rect 3231 1128 3265 1162
rect 3231 1059 3265 1093
rect 3319 1332 3353 1366
rect 3319 1264 3353 1298
rect 3319 1196 3353 1230
rect 3319 1128 3353 1162
rect 3753 1332 3787 1366
rect 3753 1264 3787 1298
rect 3753 1196 3787 1230
rect 3753 1128 3787 1162
rect 3753 1059 3787 1093
rect 3841 1332 3875 1366
rect 3841 1264 3875 1298
rect 3841 1196 3875 1230
rect 3841 1128 3875 1162
rect 3841 1059 3875 1093
rect 3929 1332 3963 1366
rect 3929 1264 3963 1298
rect 3929 1196 3963 1230
rect 3929 1128 3963 1162
rect 4017 1332 4051 1366
rect 4017 1264 4051 1298
rect 4017 1196 4051 1230
rect 4017 1128 4051 1162
rect 4017 1059 4051 1093
rect 4105 1332 4139 1366
rect 4105 1264 4139 1298
rect 4105 1196 4139 1230
rect 4105 1128 4139 1162
rect 4193 1332 4227 1366
rect 4193 1264 4227 1298
rect 4193 1196 4227 1230
rect 4193 1128 4227 1162
rect 4193 1059 4227 1093
rect 4281 1332 4315 1366
rect 4281 1264 4315 1298
rect 4281 1196 4315 1230
rect 4281 1128 4315 1162
rect 4655 1332 4689 1366
rect 4655 1264 4689 1298
rect 4655 1196 4689 1230
rect 4655 1128 4689 1162
rect 4655 1059 4689 1093
rect 4743 1332 4777 1366
rect 4743 1264 4777 1298
rect 4743 1196 4777 1230
rect 4743 1128 4777 1162
rect 4743 1059 4777 1093
rect 4831 1332 4865 1366
rect 4831 1264 4865 1298
rect 4831 1196 4865 1230
rect 4831 1128 4865 1162
rect 4919 1332 4953 1366
rect 4919 1264 4953 1298
rect 4919 1196 4953 1230
rect 4919 1128 4953 1162
rect 4919 1059 4953 1093
rect 5007 1332 5041 1366
rect 5007 1264 5041 1298
rect 5007 1196 5041 1230
rect 5007 1128 5041 1162
rect 5381 1332 5415 1366
rect 5381 1264 5415 1298
rect 5381 1196 5415 1230
rect 5381 1128 5415 1162
rect 5381 1059 5415 1093
rect 5469 1332 5503 1366
rect 5469 1264 5503 1298
rect 5469 1196 5503 1230
rect 5469 1128 5503 1162
rect 5469 1059 5503 1093
rect 5557 1332 5591 1366
rect 5557 1264 5591 1298
rect 5557 1196 5591 1230
rect 5557 1128 5591 1162
rect 5645 1332 5679 1366
rect 5645 1264 5679 1298
rect 5645 1196 5679 1230
rect 5645 1128 5679 1162
rect 5645 1059 5679 1093
rect 5733 1332 5767 1366
rect 5733 1264 5767 1298
rect 5733 1196 5767 1230
rect 5733 1128 5767 1162
rect 5821 1332 5855 1366
rect 5821 1264 5855 1298
rect 5821 1196 5855 1230
rect 5821 1128 5855 1162
rect 5821 1059 5855 1093
rect 5909 1332 5943 1366
rect 5909 1264 5943 1298
rect 5909 1196 5943 1230
rect 5909 1128 5943 1162
rect 6343 1332 6377 1366
rect 6343 1264 6377 1298
rect 6343 1196 6377 1230
rect 6343 1128 6377 1162
rect 6343 1059 6377 1093
rect 6431 1332 6465 1366
rect 6431 1264 6465 1298
rect 6431 1196 6465 1230
rect 6431 1128 6465 1162
rect 6431 1059 6465 1093
rect 6519 1332 6553 1366
rect 6519 1264 6553 1298
rect 6519 1196 6553 1230
rect 6519 1128 6553 1162
rect 6607 1332 6641 1366
rect 6607 1264 6641 1298
rect 6607 1196 6641 1230
rect 6607 1128 6641 1162
rect 6607 1059 6641 1093
rect 6695 1332 6729 1366
rect 6695 1264 6729 1298
rect 6695 1196 6729 1230
rect 6695 1128 6729 1162
rect 6783 1332 6817 1366
rect 6783 1264 6817 1298
rect 6783 1196 6817 1230
rect 6783 1128 6817 1162
rect 6783 1059 6817 1093
rect 6871 1332 6905 1366
rect 6871 1264 6905 1298
rect 6871 1196 6905 1230
rect 6871 1128 6905 1162
rect 7245 1332 7279 1366
rect 7245 1264 7279 1298
rect 7245 1196 7279 1230
rect 7245 1128 7279 1162
rect 7245 1059 7279 1093
rect 7333 1332 7367 1366
rect 7333 1264 7367 1298
rect 7333 1196 7367 1230
rect 7333 1128 7367 1162
rect 7333 1059 7367 1093
rect 7421 1332 7455 1366
rect 7421 1264 7455 1298
rect 7421 1196 7455 1230
rect 7421 1128 7455 1162
rect 7509 1332 7543 1366
rect 7509 1264 7543 1298
rect 7509 1196 7543 1230
rect 7509 1128 7543 1162
rect 7509 1059 7543 1093
rect 7597 1332 7631 1366
rect 7597 1264 7631 1298
rect 7597 1196 7631 1230
rect 7597 1128 7631 1162
rect 7971 1332 8005 1366
rect 7971 1264 8005 1298
rect 7971 1196 8005 1230
rect 7971 1128 8005 1162
rect 7971 1059 8005 1093
rect 8059 1332 8093 1366
rect 8059 1264 8093 1298
rect 8059 1196 8093 1230
rect 8059 1128 8093 1162
rect 8059 1059 8093 1093
rect 8147 1332 8181 1366
rect 8147 1264 8181 1298
rect 8147 1196 8181 1230
rect 8147 1128 8181 1162
rect 8235 1332 8269 1366
rect 8235 1264 8269 1298
rect 8235 1196 8269 1230
rect 8235 1128 8269 1162
rect 8235 1059 8269 1093
rect 8323 1332 8357 1366
rect 8323 1264 8357 1298
rect 8323 1196 8357 1230
rect 8323 1128 8357 1162
rect 8411 1332 8445 1366
rect 8411 1264 8445 1298
rect 8411 1196 8445 1230
rect 8411 1128 8445 1162
rect 8411 1059 8445 1093
rect 8499 1332 8533 1366
rect 8499 1264 8533 1298
rect 8499 1196 8533 1230
rect 8499 1128 8533 1162
rect 8933 1332 8967 1366
rect 8933 1264 8967 1298
rect 8933 1196 8967 1230
rect 8933 1128 8967 1162
rect 8933 1059 8967 1093
rect 9021 1332 9055 1366
rect 9021 1264 9055 1298
rect 9021 1196 9055 1230
rect 9021 1128 9055 1162
rect 9021 1059 9055 1093
rect 9109 1332 9143 1366
rect 9109 1264 9143 1298
rect 9109 1196 9143 1230
rect 9109 1128 9143 1162
rect 9197 1332 9231 1366
rect 9197 1264 9231 1298
rect 9197 1196 9231 1230
rect 9197 1128 9231 1162
rect 9197 1059 9231 1093
rect 9285 1332 9319 1366
rect 9285 1264 9319 1298
rect 9285 1196 9319 1230
rect 9285 1128 9319 1162
rect 9373 1332 9407 1366
rect 9373 1264 9407 1298
rect 9373 1196 9407 1230
rect 9373 1128 9407 1162
rect 9373 1059 9407 1093
rect 9461 1332 9495 1366
rect 9461 1264 9495 1298
rect 9461 1196 9495 1230
rect 9461 1128 9495 1162
rect 9835 1332 9869 1366
rect 9835 1264 9869 1298
rect 9835 1196 9869 1230
rect 9835 1128 9869 1162
rect 9835 1059 9869 1093
rect 9923 1332 9957 1366
rect 9923 1264 9957 1298
rect 9923 1196 9957 1230
rect 9923 1128 9957 1162
rect 9923 1059 9957 1093
rect 10011 1332 10045 1366
rect 10011 1264 10045 1298
rect 10011 1196 10045 1230
rect 10011 1128 10045 1162
rect 10099 1332 10133 1366
rect 10099 1264 10133 1298
rect 10099 1196 10133 1230
rect 10099 1128 10133 1162
rect 10099 1059 10133 1093
rect 10187 1332 10221 1366
rect 10187 1264 10221 1298
rect 10187 1196 10221 1230
rect 10187 1128 10221 1162
rect 10561 1332 10595 1366
rect 10561 1264 10595 1298
rect 10561 1196 10595 1230
rect 10561 1128 10595 1162
rect 10561 1059 10595 1093
rect 10649 1332 10683 1366
rect 10649 1264 10683 1298
rect 10649 1196 10683 1230
rect 10649 1128 10683 1162
rect 10649 1059 10683 1093
rect 10737 1332 10771 1366
rect 10737 1264 10771 1298
rect 10737 1196 10771 1230
rect 10737 1128 10771 1162
rect 10825 1332 10859 1366
rect 10825 1264 10859 1298
rect 10825 1196 10859 1230
rect 10825 1128 10859 1162
rect 10825 1059 10859 1093
rect 10913 1332 10947 1366
rect 10913 1264 10947 1298
rect 10913 1196 10947 1230
rect 10913 1128 10947 1162
rect 11001 1332 11035 1366
rect 11001 1264 11035 1298
rect 11001 1196 11035 1230
rect 11001 1128 11035 1162
rect 11001 1059 11035 1093
rect 11089 1332 11123 1366
rect 11089 1264 11123 1298
rect 11089 1196 11123 1230
rect 11089 1128 11123 1162
rect 11523 1332 11557 1366
rect 11523 1264 11557 1298
rect 11523 1196 11557 1230
rect 11523 1128 11557 1162
rect 11523 1059 11557 1093
rect 11611 1332 11645 1366
rect 11611 1264 11645 1298
rect 11611 1196 11645 1230
rect 11611 1128 11645 1162
rect 11611 1059 11645 1093
rect 11699 1332 11733 1366
rect 11699 1264 11733 1298
rect 11699 1196 11733 1230
rect 11699 1128 11733 1162
rect 11787 1332 11821 1366
rect 11787 1264 11821 1298
rect 11787 1196 11821 1230
rect 11787 1128 11821 1162
rect 11787 1059 11821 1093
rect 11875 1332 11909 1366
rect 11875 1264 11909 1298
rect 11875 1196 11909 1230
rect 11875 1128 11909 1162
rect 11963 1332 11997 1366
rect 11963 1264 11997 1298
rect 11963 1196 11997 1230
rect 11963 1128 11997 1162
rect 11963 1059 11997 1093
rect 12051 1332 12085 1366
rect 12051 1264 12085 1298
rect 12051 1196 12085 1230
rect 12051 1128 12085 1162
rect 12425 1332 12459 1366
rect 12425 1264 12459 1298
rect 12425 1196 12459 1230
rect 12425 1128 12459 1162
rect 12425 1059 12459 1093
rect 12513 1332 12547 1366
rect 12513 1264 12547 1298
rect 12513 1196 12547 1230
rect 12513 1128 12547 1162
rect 12513 1059 12547 1093
rect 12601 1332 12635 1366
rect 12601 1264 12635 1298
rect 12601 1196 12635 1230
rect 12601 1128 12635 1162
rect 12689 1332 12723 1366
rect 12689 1264 12723 1298
rect 12689 1196 12723 1230
rect 12689 1128 12723 1162
rect 12689 1059 12723 1093
rect 12777 1332 12811 1366
rect 12777 1264 12811 1298
rect 12777 1196 12811 1230
rect 12777 1128 12811 1162
rect 13151 1332 13185 1366
rect 13151 1264 13185 1298
rect 13151 1196 13185 1230
rect 13151 1128 13185 1162
rect 13151 1059 13185 1093
rect 13239 1332 13273 1366
rect 13239 1264 13273 1298
rect 13239 1196 13273 1230
rect 13239 1128 13273 1162
rect 13239 1059 13273 1093
rect 13327 1332 13361 1366
rect 13327 1264 13361 1298
rect 13327 1196 13361 1230
rect 13327 1128 13361 1162
rect 13415 1332 13449 1366
rect 13415 1264 13449 1298
rect 13415 1196 13449 1230
rect 13415 1128 13449 1162
rect 13415 1059 13449 1093
rect 13503 1332 13537 1366
rect 13503 1264 13537 1298
rect 13503 1196 13537 1230
rect 13503 1128 13537 1162
rect 13591 1332 13625 1366
rect 13591 1264 13625 1298
rect 13591 1196 13625 1230
rect 13591 1128 13625 1162
rect 13591 1059 13625 1093
rect 13679 1332 13713 1366
rect 13679 1264 13713 1298
rect 13679 1196 13713 1230
rect 13679 1128 13713 1162
rect 14113 1332 14147 1366
rect 14113 1264 14147 1298
rect 14113 1196 14147 1230
rect 14113 1128 14147 1162
rect 14113 1059 14147 1093
rect 14201 1332 14235 1366
rect 14201 1264 14235 1298
rect 14201 1196 14235 1230
rect 14201 1128 14235 1162
rect 14201 1059 14235 1093
rect 14289 1332 14323 1366
rect 14289 1264 14323 1298
rect 14289 1196 14323 1230
rect 14289 1128 14323 1162
rect 14377 1332 14411 1366
rect 14377 1264 14411 1298
rect 14377 1196 14411 1230
rect 14377 1128 14411 1162
rect 14377 1059 14411 1093
rect 14465 1332 14499 1366
rect 14465 1264 14499 1298
rect 14465 1196 14499 1230
rect 14465 1128 14499 1162
rect 14553 1332 14587 1366
rect 14553 1264 14587 1298
rect 14553 1196 14587 1230
rect 14553 1128 14587 1162
rect 14553 1059 14587 1093
rect 14641 1332 14675 1366
rect 14641 1264 14675 1298
rect 14641 1196 14675 1230
rect 14641 1128 14675 1162
rect 15015 1332 15049 1366
rect 15015 1264 15049 1298
rect 15015 1196 15049 1230
rect 15015 1128 15049 1162
rect 15015 1059 15049 1093
rect 15103 1332 15137 1366
rect 15103 1264 15137 1298
rect 15103 1196 15137 1230
rect 15103 1128 15137 1162
rect 15103 1059 15137 1093
rect 15191 1332 15225 1366
rect 15191 1264 15225 1298
rect 15191 1196 15225 1230
rect 15191 1128 15225 1162
rect 15279 1332 15313 1366
rect 15279 1264 15313 1298
rect 15279 1196 15313 1230
rect 15279 1128 15313 1162
rect 15279 1059 15313 1093
rect 15367 1332 15401 1366
rect 15367 1264 15401 1298
rect 15367 1196 15401 1230
rect 15367 1128 15401 1162
rect 15681 1331 15715 1365
rect 15681 1263 15715 1297
rect 15681 1195 15715 1229
rect 15681 1127 15715 1161
rect 15681 1059 15715 1093
rect 15769 1331 15803 1365
rect 15769 1263 15803 1297
rect 15769 1195 15803 1229
rect 15769 1127 15803 1161
rect 15769 1059 15803 1093
rect 15857 1331 15891 1365
rect 15857 1263 15891 1297
rect 15857 1195 15891 1229
rect 15857 1127 15891 1161
rect 15945 1331 15979 1365
rect 15945 1263 15979 1297
rect 15945 1195 15979 1229
rect 15945 1127 15979 1161
rect 16033 1331 16067 1365
rect 16033 1263 16067 1297
rect 16033 1195 16067 1229
rect 16033 1127 16067 1161
rect 16033 1059 16067 1093
rect 16345 1331 16379 1365
rect 16345 1263 16379 1297
rect 16345 1195 16379 1229
rect 16345 1127 16379 1161
rect 16433 1263 16467 1297
rect 16433 1195 16467 1229
rect 16433 1127 16467 1161
rect 16433 1059 16467 1093
rect 16521 1331 16555 1365
rect 16521 1263 16555 1297
rect 16521 1195 16555 1229
rect 16521 1127 16555 1161
rect 16609 1263 16643 1297
rect 16609 1195 16643 1229
rect 16609 1127 16643 1161
rect 16697 1331 16731 1365
rect 16697 1263 16731 1297
rect 16697 1195 16731 1229
rect 16697 1127 16731 1161
rect 17013 1331 17047 1365
rect 17013 1263 17047 1297
rect 17013 1195 17047 1229
rect 17013 1127 17047 1161
rect 17101 1263 17135 1297
rect 17101 1195 17135 1229
rect 17101 1127 17135 1161
rect 17101 1059 17135 1093
rect 17189 1331 17223 1365
rect 17189 1263 17223 1297
rect 17189 1195 17223 1229
rect 17189 1127 17223 1161
rect 17277 1263 17311 1297
rect 17277 1195 17311 1229
rect 17277 1127 17311 1161
rect 17277 1059 17311 1093
rect 17365 1331 17399 1365
rect 17365 1263 17399 1297
rect 17365 1195 17399 1229
rect 17365 1127 17399 1161
rect 17656 1332 17690 1366
rect 17656 1264 17690 1298
rect 17656 1196 17690 1230
rect 17656 1128 17690 1162
rect 17656 1059 17690 1093
rect 17744 1332 17778 1366
rect 17744 1264 17778 1298
rect 17744 1196 17778 1230
rect 17744 1128 17778 1162
rect 17744 1059 17778 1093
rect 17832 1332 17866 1366
rect 17832 1264 17866 1298
rect 17832 1196 17866 1230
rect 17832 1128 17866 1162
rect 17832 1059 17866 1093
<< psubdiff >>
rect -34 482 18016 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 928 461 996 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 928 427 945 461
rect 979 427 996 461
rect 1890 461 1958 482
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 928 313 996 353
rect 1890 427 1907 461
rect 1941 427 1958 461
rect 2556 461 2624 482
rect 1890 387 1958 427
rect 1890 353 1907 387
rect 1941 353 1958 387
rect 928 279 945 313
rect 979 279 996 313
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect -34 17 34 57
rect 928 57 945 91
rect 979 57 996 91
rect 1890 313 1958 353
rect 2556 427 2573 461
rect 2607 427 2624 461
rect 3518 461 3586 482
rect 2556 387 2624 427
rect 2556 353 2573 387
rect 2607 353 2624 387
rect 1890 279 1907 313
rect 1941 279 1958 313
rect 1890 239 1958 279
rect 1890 205 1907 239
rect 1941 205 1958 239
rect 1890 165 1958 205
rect 1890 131 1907 165
rect 1941 131 1958 165
rect 1890 91 1958 131
rect 928 17 996 57
rect 1890 57 1907 91
rect 1941 57 1958 91
rect 2556 313 2624 353
rect 3518 427 3535 461
rect 3569 427 3586 461
rect 4480 461 4548 482
rect 3518 387 3586 427
rect 3518 353 3535 387
rect 3569 353 3586 387
rect 2556 279 2573 313
rect 2607 279 2624 313
rect 2556 239 2624 279
rect 2556 205 2573 239
rect 2607 205 2624 239
rect 2556 165 2624 205
rect 2556 131 2573 165
rect 2607 131 2624 165
rect 2556 91 2624 131
rect 1890 17 1958 57
rect 2556 57 2573 91
rect 2607 57 2624 91
rect 3518 313 3586 353
rect 4480 427 4497 461
rect 4531 427 4548 461
rect 5146 461 5214 482
rect 4480 387 4548 427
rect 4480 353 4497 387
rect 4531 353 4548 387
rect 3518 279 3535 313
rect 3569 279 3586 313
rect 3518 239 3586 279
rect 3518 205 3535 239
rect 3569 205 3586 239
rect 3518 165 3586 205
rect 3518 131 3535 165
rect 3569 131 3586 165
rect 3518 91 3586 131
rect 2556 17 2624 57
rect 3518 57 3535 91
rect 3569 57 3586 91
rect 4480 313 4548 353
rect 5146 427 5163 461
rect 5197 427 5214 461
rect 6108 461 6176 482
rect 5146 387 5214 427
rect 5146 353 5163 387
rect 5197 353 5214 387
rect 4480 279 4497 313
rect 4531 279 4548 313
rect 4480 239 4548 279
rect 4480 205 4497 239
rect 4531 205 4548 239
rect 4480 165 4548 205
rect 4480 131 4497 165
rect 4531 131 4548 165
rect 4480 91 4548 131
rect 3518 17 3586 57
rect 4480 57 4497 91
rect 4531 57 4548 91
rect 5146 313 5214 353
rect 6108 427 6125 461
rect 6159 427 6176 461
rect 7070 461 7138 482
rect 6108 387 6176 427
rect 6108 353 6125 387
rect 6159 353 6176 387
rect 5146 279 5163 313
rect 5197 279 5214 313
rect 5146 239 5214 279
rect 5146 205 5163 239
rect 5197 205 5214 239
rect 5146 165 5214 205
rect 5146 131 5163 165
rect 5197 131 5214 165
rect 5146 91 5214 131
rect 4480 17 4548 57
rect 5146 57 5163 91
rect 5197 57 5214 91
rect 6108 313 6176 353
rect 7070 427 7087 461
rect 7121 427 7138 461
rect 7736 461 7804 482
rect 7070 387 7138 427
rect 7070 353 7087 387
rect 7121 353 7138 387
rect 6108 279 6125 313
rect 6159 279 6176 313
rect 6108 239 6176 279
rect 6108 205 6125 239
rect 6159 205 6176 239
rect 6108 165 6176 205
rect 6108 131 6125 165
rect 6159 131 6176 165
rect 6108 91 6176 131
rect 5146 17 5214 57
rect 6108 57 6125 91
rect 6159 57 6176 91
rect 7070 313 7138 353
rect 7736 427 7753 461
rect 7787 427 7804 461
rect 8698 461 8766 482
rect 7736 387 7804 427
rect 7736 353 7753 387
rect 7787 353 7804 387
rect 7070 279 7087 313
rect 7121 279 7138 313
rect 7070 239 7138 279
rect 7070 205 7087 239
rect 7121 205 7138 239
rect 7070 165 7138 205
rect 7070 131 7087 165
rect 7121 131 7138 165
rect 7070 91 7138 131
rect 6108 17 6176 57
rect 7070 57 7087 91
rect 7121 57 7138 91
rect 7736 313 7804 353
rect 8698 427 8715 461
rect 8749 427 8766 461
rect 9660 461 9728 482
rect 8698 387 8766 427
rect 8698 353 8715 387
rect 8749 353 8766 387
rect 7736 279 7753 313
rect 7787 279 7804 313
rect 7736 239 7804 279
rect 7736 205 7753 239
rect 7787 205 7804 239
rect 7736 165 7804 205
rect 7736 131 7753 165
rect 7787 131 7804 165
rect 7736 91 7804 131
rect 7070 17 7138 57
rect 7736 57 7753 91
rect 7787 57 7804 91
rect 8698 313 8766 353
rect 9660 427 9677 461
rect 9711 427 9728 461
rect 10326 461 10394 482
rect 9660 387 9728 427
rect 9660 353 9677 387
rect 9711 353 9728 387
rect 8698 279 8715 313
rect 8749 279 8766 313
rect 8698 239 8766 279
rect 8698 205 8715 239
rect 8749 205 8766 239
rect 8698 165 8766 205
rect 8698 131 8715 165
rect 8749 131 8766 165
rect 8698 91 8766 131
rect 7736 17 7804 57
rect 8698 57 8715 91
rect 8749 57 8766 91
rect 9660 313 9728 353
rect 10326 427 10343 461
rect 10377 427 10394 461
rect 11288 461 11356 482
rect 10326 387 10394 427
rect 10326 353 10343 387
rect 10377 353 10394 387
rect 9660 279 9677 313
rect 9711 279 9728 313
rect 9660 239 9728 279
rect 9660 205 9677 239
rect 9711 205 9728 239
rect 9660 165 9728 205
rect 9660 131 9677 165
rect 9711 131 9728 165
rect 9660 91 9728 131
rect 8698 17 8766 57
rect 9660 57 9677 91
rect 9711 57 9728 91
rect 10326 313 10394 353
rect 11288 427 11305 461
rect 11339 427 11356 461
rect 12250 461 12318 482
rect 11288 387 11356 427
rect 11288 353 11305 387
rect 11339 353 11356 387
rect 10326 279 10343 313
rect 10377 279 10394 313
rect 10326 239 10394 279
rect 10326 205 10343 239
rect 10377 205 10394 239
rect 10326 165 10394 205
rect 10326 131 10343 165
rect 10377 131 10394 165
rect 10326 91 10394 131
rect 9660 17 9728 57
rect 10326 57 10343 91
rect 10377 57 10394 91
rect 11288 313 11356 353
rect 12250 427 12267 461
rect 12301 427 12318 461
rect 12916 461 12984 482
rect 12250 387 12318 427
rect 12250 353 12267 387
rect 12301 353 12318 387
rect 11288 279 11305 313
rect 11339 279 11356 313
rect 11288 239 11356 279
rect 11288 205 11305 239
rect 11339 205 11356 239
rect 11288 165 11356 205
rect 11288 131 11305 165
rect 11339 131 11356 165
rect 11288 91 11356 131
rect 10326 17 10394 57
rect 11288 57 11305 91
rect 11339 57 11356 91
rect 12250 313 12318 353
rect 12916 427 12933 461
rect 12967 427 12984 461
rect 13878 461 13946 482
rect 12916 387 12984 427
rect 12916 353 12933 387
rect 12967 353 12984 387
rect 12250 279 12267 313
rect 12301 279 12318 313
rect 12250 239 12318 279
rect 12250 205 12267 239
rect 12301 205 12318 239
rect 12250 165 12318 205
rect 12250 131 12267 165
rect 12301 131 12318 165
rect 12250 91 12318 131
rect 11288 17 11356 57
rect 12250 57 12267 91
rect 12301 57 12318 91
rect 12916 313 12984 353
rect 13878 427 13895 461
rect 13929 427 13946 461
rect 14840 461 14908 482
rect 13878 387 13946 427
rect 13878 353 13895 387
rect 13929 353 13946 387
rect 12916 279 12933 313
rect 12967 279 12984 313
rect 12916 239 12984 279
rect 12916 205 12933 239
rect 12967 205 12984 239
rect 12916 165 12984 205
rect 12916 131 12933 165
rect 12967 131 12984 165
rect 12916 91 12984 131
rect 12250 17 12318 57
rect 12916 57 12933 91
rect 12967 57 12984 91
rect 13878 313 13946 353
rect 14840 427 14857 461
rect 14891 427 14908 461
rect 15506 461 15574 482
rect 14840 387 14908 427
rect 14840 353 14857 387
rect 14891 353 14908 387
rect 13878 279 13895 313
rect 13929 279 13946 313
rect 13878 239 13946 279
rect 13878 205 13895 239
rect 13929 205 13946 239
rect 13878 165 13946 205
rect 13878 131 13895 165
rect 13929 131 13946 165
rect 13878 91 13946 131
rect 12916 17 12984 57
rect 13878 57 13895 91
rect 13929 57 13946 91
rect 14840 313 14908 353
rect 15506 427 15523 461
rect 15557 427 15574 461
rect 16172 461 16240 482
rect 15506 387 15574 427
rect 15506 353 15523 387
rect 15557 353 15574 387
rect 16172 427 16189 461
rect 16223 427 16240 461
rect 16838 461 16906 482
rect 16172 387 16240 427
rect 14840 279 14857 313
rect 14891 279 14908 313
rect 14840 239 14908 279
rect 14840 205 14857 239
rect 14891 205 14908 239
rect 14840 165 14908 205
rect 14840 131 14857 165
rect 14891 131 14908 165
rect 14840 91 14908 131
rect 13878 17 13946 57
rect 14840 57 14857 91
rect 14891 57 14908 91
rect 15506 313 15574 353
rect 16172 353 16189 387
rect 16223 353 16240 387
rect 15506 279 15523 313
rect 15557 279 15574 313
rect 15506 239 15574 279
rect 15506 205 15523 239
rect 15557 205 15574 239
rect 15506 165 15574 205
rect 15506 131 15523 165
rect 15557 131 15574 165
rect 15506 91 15574 131
rect 14840 17 14908 57
rect 15506 57 15523 91
rect 15557 57 15574 91
rect 16172 313 16240 353
rect 16838 427 16855 461
rect 16889 427 16906 461
rect 17504 461 17572 482
rect 16838 387 16906 427
rect 16838 353 16855 387
rect 16889 353 16906 387
rect 17504 427 17521 461
rect 17555 427 17572 461
rect 17948 461 18016 482
rect 17504 387 17572 427
rect 16172 279 16189 313
rect 16223 279 16240 313
rect 16172 239 16240 279
rect 16172 205 16189 239
rect 16223 205 16240 239
rect 16172 165 16240 205
rect 16172 131 16189 165
rect 16223 131 16240 165
rect 16172 91 16240 131
rect 15506 17 15574 57
rect 16172 57 16189 91
rect 16223 57 16240 91
rect 16838 313 16906 353
rect 17504 353 17521 387
rect 17555 353 17572 387
rect 17948 427 17965 461
rect 17999 427 18016 461
rect 16838 279 16855 313
rect 16889 279 16906 313
rect 16838 239 16906 279
rect 16838 205 16855 239
rect 16889 205 16906 239
rect 16838 165 16906 205
rect 16838 131 16855 165
rect 16889 131 16906 165
rect 16838 91 16906 131
rect 16172 17 16240 57
rect 16838 57 16855 91
rect 16889 57 16906 91
rect 17504 313 17572 353
rect 17948 387 18016 427
rect 17948 353 17965 387
rect 17999 353 18016 387
rect 17504 279 17521 313
rect 17555 279 17572 313
rect 17504 239 17572 279
rect 17504 205 17521 239
rect 17555 205 17572 239
rect 17504 165 17572 205
rect 17504 131 17521 165
rect 17555 131 17572 165
rect 17504 91 17572 131
rect 16838 17 16906 57
rect 17504 57 17521 91
rect 17555 57 17572 91
rect 17948 313 18016 353
rect 17948 279 17965 313
rect 17999 279 18016 313
rect 17948 239 18016 279
rect 17948 205 17965 239
rect 17999 205 18016 239
rect 17948 165 18016 205
rect 17948 131 17965 165
rect 17999 131 18016 165
rect 17948 91 18016 131
rect 17504 17 17572 57
rect 17948 57 17965 91
rect 17999 57 18016 91
rect 17948 17 18016 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5533 17
rect 5567 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5755 17
rect 5789 -17 5829 17
rect 5863 -17 5903 17
rect 5937 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6199 17
rect 6233 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6495 17
rect 6529 -17 6569 17
rect 6603 -17 6643 17
rect 6677 -17 6717 17
rect 6751 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7161 17
rect 7195 -17 7235 17
rect 7269 -17 7309 17
rect 7343 -17 7383 17
rect 7417 -17 7457 17
rect 7491 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7679 17
rect 7713 -17 7827 17
rect 7861 -17 7901 17
rect 7935 -17 7975 17
rect 8009 -17 8049 17
rect 8083 -17 8123 17
rect 8157 -17 8197 17
rect 8231 -17 8271 17
rect 8305 -17 8345 17
rect 8379 -17 8419 17
rect 8453 -17 8493 17
rect 8527 -17 8567 17
rect 8601 -17 8641 17
rect 8675 -17 8789 17
rect 8823 -17 8863 17
rect 8897 -17 8937 17
rect 8971 -17 9011 17
rect 9045 -17 9085 17
rect 9119 -17 9159 17
rect 9193 -17 9233 17
rect 9267 -17 9307 17
rect 9341 -17 9381 17
rect 9415 -17 9455 17
rect 9489 -17 9529 17
rect 9563 -17 9603 17
rect 9637 -17 9751 17
rect 9785 -17 9825 17
rect 9859 -17 9899 17
rect 9933 -17 9973 17
rect 10007 -17 10047 17
rect 10081 -17 10121 17
rect 10155 -17 10195 17
rect 10229 -17 10269 17
rect 10303 -17 10417 17
rect 10451 -17 10491 17
rect 10525 -17 10565 17
rect 10599 -17 10639 17
rect 10673 -17 10713 17
rect 10747 -17 10787 17
rect 10821 -17 10861 17
rect 10895 -17 10935 17
rect 10969 -17 11009 17
rect 11043 -17 11083 17
rect 11117 -17 11157 17
rect 11191 -17 11231 17
rect 11265 -17 11379 17
rect 11413 -17 11453 17
rect 11487 -17 11527 17
rect 11561 -17 11601 17
rect 11635 -17 11675 17
rect 11709 -17 11749 17
rect 11783 -17 11823 17
rect 11857 -17 11897 17
rect 11931 -17 11971 17
rect 12005 -17 12045 17
rect 12079 -17 12119 17
rect 12153 -17 12193 17
rect 12227 -17 12341 17
rect 12375 -17 12415 17
rect 12449 -17 12489 17
rect 12523 -17 12563 17
rect 12597 -17 12637 17
rect 12671 -17 12711 17
rect 12745 -17 12785 17
rect 12819 -17 12859 17
rect 12893 -17 13007 17
rect 13041 -17 13081 17
rect 13115 -17 13155 17
rect 13189 -17 13229 17
rect 13263 -17 13303 17
rect 13337 -17 13377 17
rect 13411 -17 13451 17
rect 13485 -17 13525 17
rect 13559 -17 13599 17
rect 13633 -17 13673 17
rect 13707 -17 13747 17
rect 13781 -17 13821 17
rect 13855 -17 13969 17
rect 14003 -17 14043 17
rect 14077 -17 14117 17
rect 14151 -17 14191 17
rect 14225 -17 14265 17
rect 14299 -17 14339 17
rect 14373 -17 14413 17
rect 14447 -17 14487 17
rect 14521 -17 14561 17
rect 14595 -17 14635 17
rect 14669 -17 14709 17
rect 14743 -17 14783 17
rect 14817 -17 14931 17
rect 14965 -17 15005 17
rect 15039 -17 15079 17
rect 15113 -17 15153 17
rect 15187 -17 15227 17
rect 15261 -17 15301 17
rect 15335 -17 15375 17
rect 15409 -17 15449 17
rect 15483 -17 15597 17
rect 15631 -17 15671 17
rect 15705 -17 15745 17
rect 15779 -17 15819 17
rect 15853 -17 15893 17
rect 15927 -17 15967 17
rect 16001 -17 16041 17
rect 16075 -17 16115 17
rect 16149 -17 16263 17
rect 16297 -17 16337 17
rect 16371 -17 16411 17
rect 16445 -17 16485 17
rect 16519 -17 16559 17
rect 16593 -17 16633 17
rect 16667 -17 16707 17
rect 16741 -17 16781 17
rect 16815 -17 16929 17
rect 16963 -17 17003 17
rect 17037 -17 17077 17
rect 17111 -17 17151 17
rect 17185 -17 17225 17
rect 17259 -17 17299 17
rect 17333 -17 17373 17
rect 17407 -17 17447 17
rect 17481 -17 17595 17
rect 17629 -17 17669 17
rect 17703 -17 17743 17
rect 17777 -17 17817 17
rect 17851 -17 17891 17
rect 17925 -17 18016 17
rect -34 -34 18016 -17
<< nsubdiff >>
rect -34 1497 18016 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5533 1497
rect 5567 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5755 1497
rect 5789 1463 5829 1497
rect 5863 1463 5903 1497
rect 5937 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6199 1497
rect 6233 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6495 1497
rect 6529 1463 6569 1497
rect 6603 1463 6643 1497
rect 6677 1463 6717 1497
rect 6751 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7161 1497
rect 7195 1463 7235 1497
rect 7269 1463 7309 1497
rect 7343 1463 7383 1497
rect 7417 1463 7457 1497
rect 7491 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7679 1497
rect 7713 1463 7827 1497
rect 7861 1463 7901 1497
rect 7935 1463 7975 1497
rect 8009 1463 8049 1497
rect 8083 1463 8123 1497
rect 8157 1463 8197 1497
rect 8231 1463 8271 1497
rect 8305 1463 8345 1497
rect 8379 1463 8419 1497
rect 8453 1463 8493 1497
rect 8527 1463 8567 1497
rect 8601 1463 8641 1497
rect 8675 1463 8789 1497
rect 8823 1463 8863 1497
rect 8897 1463 8937 1497
rect 8971 1463 9011 1497
rect 9045 1463 9085 1497
rect 9119 1463 9159 1497
rect 9193 1463 9233 1497
rect 9267 1463 9307 1497
rect 9341 1463 9381 1497
rect 9415 1463 9455 1497
rect 9489 1463 9529 1497
rect 9563 1463 9603 1497
rect 9637 1463 9751 1497
rect 9785 1463 9825 1497
rect 9859 1463 9899 1497
rect 9933 1463 9973 1497
rect 10007 1463 10047 1497
rect 10081 1463 10121 1497
rect 10155 1463 10195 1497
rect 10229 1463 10269 1497
rect 10303 1463 10417 1497
rect 10451 1463 10491 1497
rect 10525 1463 10565 1497
rect 10599 1463 10639 1497
rect 10673 1463 10713 1497
rect 10747 1463 10787 1497
rect 10821 1463 10861 1497
rect 10895 1463 10935 1497
rect 10969 1463 11009 1497
rect 11043 1463 11083 1497
rect 11117 1463 11157 1497
rect 11191 1463 11231 1497
rect 11265 1463 11379 1497
rect 11413 1463 11453 1497
rect 11487 1463 11527 1497
rect 11561 1463 11601 1497
rect 11635 1463 11675 1497
rect 11709 1463 11749 1497
rect 11783 1463 11823 1497
rect 11857 1463 11897 1497
rect 11931 1463 11971 1497
rect 12005 1463 12045 1497
rect 12079 1463 12119 1497
rect 12153 1463 12193 1497
rect 12227 1463 12341 1497
rect 12375 1463 12415 1497
rect 12449 1463 12489 1497
rect 12523 1463 12563 1497
rect 12597 1463 12637 1497
rect 12671 1463 12711 1497
rect 12745 1463 12785 1497
rect 12819 1463 12859 1497
rect 12893 1463 13007 1497
rect 13041 1463 13081 1497
rect 13115 1463 13155 1497
rect 13189 1463 13229 1497
rect 13263 1463 13303 1497
rect 13337 1463 13377 1497
rect 13411 1463 13451 1497
rect 13485 1463 13525 1497
rect 13559 1463 13599 1497
rect 13633 1463 13673 1497
rect 13707 1463 13747 1497
rect 13781 1463 13821 1497
rect 13855 1463 13969 1497
rect 14003 1463 14043 1497
rect 14077 1463 14117 1497
rect 14151 1463 14191 1497
rect 14225 1463 14265 1497
rect 14299 1463 14339 1497
rect 14373 1463 14413 1497
rect 14447 1463 14487 1497
rect 14521 1463 14561 1497
rect 14595 1463 14635 1497
rect 14669 1463 14709 1497
rect 14743 1463 14783 1497
rect 14817 1463 14931 1497
rect 14965 1463 15005 1497
rect 15039 1463 15079 1497
rect 15113 1463 15153 1497
rect 15187 1463 15227 1497
rect 15261 1463 15301 1497
rect 15335 1463 15375 1497
rect 15409 1463 15449 1497
rect 15483 1463 15597 1497
rect 15631 1463 15671 1497
rect 15705 1463 15745 1497
rect 15779 1463 15819 1497
rect 15853 1463 15893 1497
rect 15927 1463 15967 1497
rect 16001 1463 16041 1497
rect 16075 1463 16115 1497
rect 16149 1463 16263 1497
rect 16297 1463 16337 1497
rect 16371 1463 16411 1497
rect 16445 1463 16485 1497
rect 16519 1463 16559 1497
rect 16593 1463 16633 1497
rect 16667 1463 16707 1497
rect 16741 1463 16781 1497
rect 16815 1463 16929 1497
rect 16963 1463 17003 1497
rect 17037 1463 17077 1497
rect 17111 1463 17151 1497
rect 17185 1463 17225 1497
rect 17259 1463 17299 1497
rect 17333 1463 17373 1497
rect 17407 1463 17447 1497
rect 17481 1463 17595 1497
rect 17629 1463 17669 1497
rect 17703 1463 17743 1497
rect 17777 1463 17817 1497
rect 17851 1463 17891 1497
rect 17925 1463 18016 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 928 1423 996 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 1890 1423 1958 1463
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect 928 1019 945 1053
rect 979 1019 996 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 928 979 996 1019
rect 1890 1389 1907 1423
rect 1941 1389 1958 1423
rect 2556 1423 2624 1463
rect 1890 1349 1958 1389
rect 1890 1315 1907 1349
rect 1941 1315 1958 1349
rect 1890 1275 1958 1315
rect 1890 1241 1907 1275
rect 1941 1241 1958 1275
rect 1890 1201 1958 1241
rect 1890 1167 1907 1201
rect 1941 1167 1958 1201
rect 1890 1127 1958 1167
rect 1890 1093 1907 1127
rect 1941 1093 1958 1127
rect 1890 1053 1958 1093
rect 1890 1019 1907 1053
rect 1941 1019 1958 1053
rect 928 945 945 979
rect 979 945 996 979
rect -34 871 -17 905
rect 17 884 34 905
rect 928 905 996 945
rect 1890 979 1958 1019
rect 2556 1389 2573 1423
rect 2607 1389 2624 1423
rect 3518 1423 3586 1463
rect 2556 1349 2624 1389
rect 2556 1315 2573 1349
rect 2607 1315 2624 1349
rect 2556 1275 2624 1315
rect 2556 1241 2573 1275
rect 2607 1241 2624 1275
rect 2556 1201 2624 1241
rect 2556 1167 2573 1201
rect 2607 1167 2624 1201
rect 2556 1127 2624 1167
rect 2556 1093 2573 1127
rect 2607 1093 2624 1127
rect 2556 1053 2624 1093
rect 2556 1019 2573 1053
rect 2607 1019 2624 1053
rect 1890 945 1907 979
rect 1941 945 1958 979
rect 928 884 945 905
rect 17 871 945 884
rect 979 884 996 905
rect 1890 905 1958 945
rect 2556 979 2624 1019
rect 3518 1389 3535 1423
rect 3569 1389 3586 1423
rect 4480 1423 4548 1463
rect 3518 1349 3586 1389
rect 3518 1315 3535 1349
rect 3569 1315 3586 1349
rect 3518 1275 3586 1315
rect 3518 1241 3535 1275
rect 3569 1241 3586 1275
rect 3518 1201 3586 1241
rect 3518 1167 3535 1201
rect 3569 1167 3586 1201
rect 3518 1127 3586 1167
rect 3518 1093 3535 1127
rect 3569 1093 3586 1127
rect 3518 1053 3586 1093
rect 3518 1019 3535 1053
rect 3569 1019 3586 1053
rect 2556 945 2573 979
rect 2607 945 2624 979
rect 1890 884 1907 905
rect 979 871 1907 884
rect 1941 884 1958 905
rect 2556 905 2624 945
rect 3518 979 3586 1019
rect 4480 1389 4497 1423
rect 4531 1389 4548 1423
rect 5146 1423 5214 1463
rect 4480 1349 4548 1389
rect 4480 1315 4497 1349
rect 4531 1315 4548 1349
rect 4480 1275 4548 1315
rect 4480 1241 4497 1275
rect 4531 1241 4548 1275
rect 4480 1201 4548 1241
rect 4480 1167 4497 1201
rect 4531 1167 4548 1201
rect 4480 1127 4548 1167
rect 4480 1093 4497 1127
rect 4531 1093 4548 1127
rect 4480 1053 4548 1093
rect 4480 1019 4497 1053
rect 4531 1019 4548 1053
rect 3518 945 3535 979
rect 3569 945 3586 979
rect 2556 884 2573 905
rect 1941 871 2573 884
rect 2607 884 2624 905
rect 3518 905 3586 945
rect 4480 979 4548 1019
rect 5146 1389 5163 1423
rect 5197 1389 5214 1423
rect 6108 1423 6176 1463
rect 5146 1349 5214 1389
rect 5146 1315 5163 1349
rect 5197 1315 5214 1349
rect 5146 1275 5214 1315
rect 5146 1241 5163 1275
rect 5197 1241 5214 1275
rect 5146 1201 5214 1241
rect 5146 1167 5163 1201
rect 5197 1167 5214 1201
rect 5146 1127 5214 1167
rect 5146 1093 5163 1127
rect 5197 1093 5214 1127
rect 5146 1053 5214 1093
rect 5146 1019 5163 1053
rect 5197 1019 5214 1053
rect 4480 945 4497 979
rect 4531 945 4548 979
rect 3518 884 3535 905
rect 2607 871 3535 884
rect 3569 884 3586 905
rect 4480 905 4548 945
rect 5146 979 5214 1019
rect 6108 1389 6125 1423
rect 6159 1389 6176 1423
rect 7070 1423 7138 1463
rect 6108 1349 6176 1389
rect 6108 1315 6125 1349
rect 6159 1315 6176 1349
rect 6108 1275 6176 1315
rect 6108 1241 6125 1275
rect 6159 1241 6176 1275
rect 6108 1201 6176 1241
rect 6108 1167 6125 1201
rect 6159 1167 6176 1201
rect 6108 1127 6176 1167
rect 6108 1093 6125 1127
rect 6159 1093 6176 1127
rect 6108 1053 6176 1093
rect 6108 1019 6125 1053
rect 6159 1019 6176 1053
rect 5146 945 5163 979
rect 5197 945 5214 979
rect 4480 884 4497 905
rect 3569 871 4497 884
rect 4531 884 4548 905
rect 5146 905 5214 945
rect 6108 979 6176 1019
rect 7070 1389 7087 1423
rect 7121 1389 7138 1423
rect 7736 1423 7804 1463
rect 7070 1349 7138 1389
rect 7070 1315 7087 1349
rect 7121 1315 7138 1349
rect 7070 1275 7138 1315
rect 7070 1241 7087 1275
rect 7121 1241 7138 1275
rect 7070 1201 7138 1241
rect 7070 1167 7087 1201
rect 7121 1167 7138 1201
rect 7070 1127 7138 1167
rect 7070 1093 7087 1127
rect 7121 1093 7138 1127
rect 7070 1053 7138 1093
rect 7070 1019 7087 1053
rect 7121 1019 7138 1053
rect 6108 945 6125 979
rect 6159 945 6176 979
rect 5146 884 5163 905
rect 4531 871 5163 884
rect 5197 884 5214 905
rect 6108 905 6176 945
rect 7070 979 7138 1019
rect 7736 1389 7753 1423
rect 7787 1389 7804 1423
rect 8698 1423 8766 1463
rect 7736 1349 7804 1389
rect 7736 1315 7753 1349
rect 7787 1315 7804 1349
rect 7736 1275 7804 1315
rect 7736 1241 7753 1275
rect 7787 1241 7804 1275
rect 7736 1201 7804 1241
rect 7736 1167 7753 1201
rect 7787 1167 7804 1201
rect 7736 1127 7804 1167
rect 7736 1093 7753 1127
rect 7787 1093 7804 1127
rect 7736 1053 7804 1093
rect 7736 1019 7753 1053
rect 7787 1019 7804 1053
rect 7070 945 7087 979
rect 7121 945 7138 979
rect 6108 884 6125 905
rect 5197 871 6125 884
rect 6159 884 6176 905
rect 7070 905 7138 945
rect 7736 979 7804 1019
rect 8698 1389 8715 1423
rect 8749 1389 8766 1423
rect 9660 1423 9728 1463
rect 8698 1349 8766 1389
rect 8698 1315 8715 1349
rect 8749 1315 8766 1349
rect 8698 1275 8766 1315
rect 8698 1241 8715 1275
rect 8749 1241 8766 1275
rect 8698 1201 8766 1241
rect 8698 1167 8715 1201
rect 8749 1167 8766 1201
rect 8698 1127 8766 1167
rect 8698 1093 8715 1127
rect 8749 1093 8766 1127
rect 8698 1053 8766 1093
rect 8698 1019 8715 1053
rect 8749 1019 8766 1053
rect 7736 945 7753 979
rect 7787 945 7804 979
rect 7070 884 7087 905
rect 6159 871 7087 884
rect 7121 884 7138 905
rect 7736 905 7804 945
rect 8698 979 8766 1019
rect 9660 1389 9677 1423
rect 9711 1389 9728 1423
rect 10326 1423 10394 1463
rect 9660 1349 9728 1389
rect 9660 1315 9677 1349
rect 9711 1315 9728 1349
rect 9660 1275 9728 1315
rect 9660 1241 9677 1275
rect 9711 1241 9728 1275
rect 9660 1201 9728 1241
rect 9660 1167 9677 1201
rect 9711 1167 9728 1201
rect 9660 1127 9728 1167
rect 9660 1093 9677 1127
rect 9711 1093 9728 1127
rect 9660 1053 9728 1093
rect 9660 1019 9677 1053
rect 9711 1019 9728 1053
rect 8698 945 8715 979
rect 8749 945 8766 979
rect 7736 884 7753 905
rect 7121 871 7753 884
rect 7787 884 7804 905
rect 8698 905 8766 945
rect 9660 979 9728 1019
rect 10326 1389 10343 1423
rect 10377 1389 10394 1423
rect 11288 1423 11356 1463
rect 10326 1349 10394 1389
rect 10326 1315 10343 1349
rect 10377 1315 10394 1349
rect 10326 1275 10394 1315
rect 10326 1241 10343 1275
rect 10377 1241 10394 1275
rect 10326 1201 10394 1241
rect 10326 1167 10343 1201
rect 10377 1167 10394 1201
rect 10326 1127 10394 1167
rect 10326 1093 10343 1127
rect 10377 1093 10394 1127
rect 10326 1053 10394 1093
rect 10326 1019 10343 1053
rect 10377 1019 10394 1053
rect 9660 945 9677 979
rect 9711 945 9728 979
rect 8698 884 8715 905
rect 7787 871 8715 884
rect 8749 884 8766 905
rect 9660 905 9728 945
rect 10326 979 10394 1019
rect 11288 1389 11305 1423
rect 11339 1389 11356 1423
rect 12250 1423 12318 1463
rect 11288 1349 11356 1389
rect 11288 1315 11305 1349
rect 11339 1315 11356 1349
rect 11288 1275 11356 1315
rect 11288 1241 11305 1275
rect 11339 1241 11356 1275
rect 11288 1201 11356 1241
rect 11288 1167 11305 1201
rect 11339 1167 11356 1201
rect 11288 1127 11356 1167
rect 11288 1093 11305 1127
rect 11339 1093 11356 1127
rect 11288 1053 11356 1093
rect 11288 1019 11305 1053
rect 11339 1019 11356 1053
rect 10326 945 10343 979
rect 10377 945 10394 979
rect 9660 884 9677 905
rect 8749 871 9677 884
rect 9711 884 9728 905
rect 10326 905 10394 945
rect 11288 979 11356 1019
rect 12250 1389 12267 1423
rect 12301 1389 12318 1423
rect 12916 1423 12984 1463
rect 12250 1349 12318 1389
rect 12250 1315 12267 1349
rect 12301 1315 12318 1349
rect 12250 1275 12318 1315
rect 12250 1241 12267 1275
rect 12301 1241 12318 1275
rect 12250 1201 12318 1241
rect 12250 1167 12267 1201
rect 12301 1167 12318 1201
rect 12250 1127 12318 1167
rect 12250 1093 12267 1127
rect 12301 1093 12318 1127
rect 12250 1053 12318 1093
rect 12250 1019 12267 1053
rect 12301 1019 12318 1053
rect 11288 945 11305 979
rect 11339 945 11356 979
rect 10326 884 10343 905
rect 9711 871 10343 884
rect 10377 884 10394 905
rect 11288 905 11356 945
rect 12250 979 12318 1019
rect 12916 1389 12933 1423
rect 12967 1389 12984 1423
rect 13878 1423 13946 1463
rect 12916 1349 12984 1389
rect 12916 1315 12933 1349
rect 12967 1315 12984 1349
rect 12916 1275 12984 1315
rect 12916 1241 12933 1275
rect 12967 1241 12984 1275
rect 12916 1201 12984 1241
rect 12916 1167 12933 1201
rect 12967 1167 12984 1201
rect 12916 1127 12984 1167
rect 12916 1093 12933 1127
rect 12967 1093 12984 1127
rect 12916 1053 12984 1093
rect 12916 1019 12933 1053
rect 12967 1019 12984 1053
rect 12250 945 12267 979
rect 12301 945 12318 979
rect 11288 884 11305 905
rect 10377 871 11305 884
rect 11339 884 11356 905
rect 12250 905 12318 945
rect 12916 979 12984 1019
rect 13878 1389 13895 1423
rect 13929 1389 13946 1423
rect 14840 1423 14908 1463
rect 13878 1349 13946 1389
rect 13878 1315 13895 1349
rect 13929 1315 13946 1349
rect 13878 1275 13946 1315
rect 13878 1241 13895 1275
rect 13929 1241 13946 1275
rect 13878 1201 13946 1241
rect 13878 1167 13895 1201
rect 13929 1167 13946 1201
rect 13878 1127 13946 1167
rect 13878 1093 13895 1127
rect 13929 1093 13946 1127
rect 13878 1053 13946 1093
rect 13878 1019 13895 1053
rect 13929 1019 13946 1053
rect 12916 945 12933 979
rect 12967 945 12984 979
rect 12250 884 12267 905
rect 11339 871 12267 884
rect 12301 884 12318 905
rect 12916 905 12984 945
rect 13878 979 13946 1019
rect 14840 1389 14857 1423
rect 14891 1389 14908 1423
rect 15506 1423 15574 1463
rect 14840 1349 14908 1389
rect 14840 1315 14857 1349
rect 14891 1315 14908 1349
rect 14840 1275 14908 1315
rect 14840 1241 14857 1275
rect 14891 1241 14908 1275
rect 14840 1201 14908 1241
rect 14840 1167 14857 1201
rect 14891 1167 14908 1201
rect 14840 1127 14908 1167
rect 14840 1093 14857 1127
rect 14891 1093 14908 1127
rect 14840 1053 14908 1093
rect 14840 1019 14857 1053
rect 14891 1019 14908 1053
rect 13878 945 13895 979
rect 13929 945 13946 979
rect 12916 884 12933 905
rect 12301 871 12933 884
rect 12967 884 12984 905
rect 13878 905 13946 945
rect 14840 979 14908 1019
rect 15506 1389 15523 1423
rect 15557 1389 15574 1423
rect 16172 1423 16240 1463
rect 15506 1349 15574 1389
rect 15506 1315 15523 1349
rect 15557 1315 15574 1349
rect 15506 1275 15574 1315
rect 15506 1241 15523 1275
rect 15557 1241 15574 1275
rect 15506 1201 15574 1241
rect 15506 1167 15523 1201
rect 15557 1167 15574 1201
rect 15506 1127 15574 1167
rect 15506 1093 15523 1127
rect 15557 1093 15574 1127
rect 15506 1053 15574 1093
rect 15506 1019 15523 1053
rect 15557 1019 15574 1053
rect 14840 945 14857 979
rect 14891 945 14908 979
rect 13878 884 13895 905
rect 12967 871 13895 884
rect 13929 884 13946 905
rect 14840 905 14908 945
rect 15506 979 15574 1019
rect 16172 1389 16189 1423
rect 16223 1389 16240 1423
rect 16838 1423 16906 1463
rect 17486 1459 17572 1463
rect 16172 1349 16240 1389
rect 16172 1315 16189 1349
rect 16223 1315 16240 1349
rect 16172 1275 16240 1315
rect 16172 1241 16189 1275
rect 16223 1241 16240 1275
rect 16172 1201 16240 1241
rect 16172 1167 16189 1201
rect 16223 1167 16240 1201
rect 16172 1127 16240 1167
rect 16172 1093 16189 1127
rect 16223 1093 16240 1127
rect 16172 1053 16240 1093
rect 16172 1019 16189 1053
rect 16223 1019 16240 1053
rect 15506 945 15523 979
rect 15557 945 15574 979
rect 14840 884 14857 905
rect 13929 871 14857 884
rect 14891 884 14908 905
rect 15506 905 15574 945
rect 16172 979 16240 1019
rect 16838 1389 16855 1423
rect 16889 1389 16906 1423
rect 17504 1423 17572 1459
rect 16838 1349 16906 1389
rect 16838 1315 16855 1349
rect 16889 1315 16906 1349
rect 16838 1275 16906 1315
rect 16838 1241 16855 1275
rect 16889 1241 16906 1275
rect 16838 1201 16906 1241
rect 16838 1167 16855 1201
rect 16889 1167 16906 1201
rect 16838 1127 16906 1167
rect 16838 1093 16855 1127
rect 16889 1093 16906 1127
rect 16838 1053 16906 1093
rect 16838 1019 16855 1053
rect 16889 1019 16906 1053
rect 16172 945 16189 979
rect 16223 945 16240 979
rect 15506 884 15523 905
rect 14891 871 15523 884
rect 15557 884 15574 905
rect 16172 905 16240 945
rect 16838 979 16906 1019
rect 17504 1389 17521 1423
rect 17555 1389 17572 1423
rect 17948 1423 18016 1463
rect 17504 1349 17572 1389
rect 17504 1315 17521 1349
rect 17555 1315 17572 1349
rect 17504 1275 17572 1315
rect 17504 1241 17521 1275
rect 17555 1241 17572 1275
rect 17504 1201 17572 1241
rect 17504 1167 17521 1201
rect 17555 1167 17572 1201
rect 17504 1127 17572 1167
rect 17504 1093 17521 1127
rect 17555 1093 17572 1127
rect 17504 1053 17572 1093
rect 17504 1019 17521 1053
rect 17555 1019 17572 1053
rect 16838 945 16855 979
rect 16889 945 16906 979
rect 16172 884 16189 905
rect 15557 871 16189 884
rect 16223 884 16240 905
rect 16838 905 16906 945
rect 17504 979 17572 1019
rect 17948 1389 17965 1423
rect 17999 1389 18016 1423
rect 17948 1349 18016 1389
rect 17948 1315 17965 1349
rect 17999 1315 18016 1349
rect 17948 1275 18016 1315
rect 17948 1241 17965 1275
rect 17999 1241 18016 1275
rect 17948 1201 18016 1241
rect 17948 1167 17965 1201
rect 17999 1167 18016 1201
rect 17948 1127 18016 1167
rect 17948 1093 17965 1127
rect 17999 1093 18016 1127
rect 17948 1053 18016 1093
rect 17948 1019 17965 1053
rect 17999 1019 18016 1053
rect 17504 945 17521 979
rect 17555 945 17572 979
rect 16838 884 16855 905
rect 16223 871 16855 884
rect 16889 884 16906 905
rect 17504 905 17572 945
rect 17948 979 18016 1019
rect 17948 945 17965 979
rect 17999 945 18016 979
rect 17504 884 17521 905
rect 16889 871 17521 884
rect 17555 884 17572 905
rect 17948 905 18016 945
rect 17948 884 17965 905
rect 17555 871 17965 884
rect 17999 871 18016 905
rect -34 822 18016 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 945 427 979 461
rect 945 353 979 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1907 427 1941 461
rect 1907 353 1941 387
rect 945 279 979 313
rect 945 205 979 239
rect 945 131 979 165
rect 945 57 979 91
rect 2573 427 2607 461
rect 2573 353 2607 387
rect 1907 279 1941 313
rect 1907 205 1941 239
rect 1907 131 1941 165
rect 1907 57 1941 91
rect 3535 427 3569 461
rect 3535 353 3569 387
rect 2573 279 2607 313
rect 2573 205 2607 239
rect 2573 131 2607 165
rect 2573 57 2607 91
rect 4497 427 4531 461
rect 4497 353 4531 387
rect 3535 279 3569 313
rect 3535 205 3569 239
rect 3535 131 3569 165
rect 3535 57 3569 91
rect 5163 427 5197 461
rect 5163 353 5197 387
rect 4497 279 4531 313
rect 4497 205 4531 239
rect 4497 131 4531 165
rect 4497 57 4531 91
rect 6125 427 6159 461
rect 6125 353 6159 387
rect 5163 279 5197 313
rect 5163 205 5197 239
rect 5163 131 5197 165
rect 5163 57 5197 91
rect 7087 427 7121 461
rect 7087 353 7121 387
rect 6125 279 6159 313
rect 6125 205 6159 239
rect 6125 131 6159 165
rect 6125 57 6159 91
rect 7753 427 7787 461
rect 7753 353 7787 387
rect 7087 279 7121 313
rect 7087 205 7121 239
rect 7087 131 7121 165
rect 7087 57 7121 91
rect 8715 427 8749 461
rect 8715 353 8749 387
rect 7753 279 7787 313
rect 7753 205 7787 239
rect 7753 131 7787 165
rect 7753 57 7787 91
rect 9677 427 9711 461
rect 9677 353 9711 387
rect 8715 279 8749 313
rect 8715 205 8749 239
rect 8715 131 8749 165
rect 8715 57 8749 91
rect 10343 427 10377 461
rect 10343 353 10377 387
rect 9677 279 9711 313
rect 9677 205 9711 239
rect 9677 131 9711 165
rect 9677 57 9711 91
rect 11305 427 11339 461
rect 11305 353 11339 387
rect 10343 279 10377 313
rect 10343 205 10377 239
rect 10343 131 10377 165
rect 10343 57 10377 91
rect 12267 427 12301 461
rect 12267 353 12301 387
rect 11305 279 11339 313
rect 11305 205 11339 239
rect 11305 131 11339 165
rect 11305 57 11339 91
rect 12933 427 12967 461
rect 12933 353 12967 387
rect 12267 279 12301 313
rect 12267 205 12301 239
rect 12267 131 12301 165
rect 12267 57 12301 91
rect 13895 427 13929 461
rect 13895 353 13929 387
rect 12933 279 12967 313
rect 12933 205 12967 239
rect 12933 131 12967 165
rect 12933 57 12967 91
rect 14857 427 14891 461
rect 14857 353 14891 387
rect 13895 279 13929 313
rect 13895 205 13929 239
rect 13895 131 13929 165
rect 13895 57 13929 91
rect 15523 427 15557 461
rect 15523 353 15557 387
rect 16189 427 16223 461
rect 14857 279 14891 313
rect 14857 205 14891 239
rect 14857 131 14891 165
rect 14857 57 14891 91
rect 16189 353 16223 387
rect 15523 279 15557 313
rect 15523 205 15557 239
rect 15523 131 15557 165
rect 15523 57 15557 91
rect 16855 427 16889 461
rect 16855 353 16889 387
rect 17521 427 17555 461
rect 16189 279 16223 313
rect 16189 205 16223 239
rect 16189 131 16223 165
rect 16189 57 16223 91
rect 17521 353 17555 387
rect 17965 427 17999 461
rect 16855 279 16889 313
rect 16855 205 16889 239
rect 16855 131 16889 165
rect 16855 57 16889 91
rect 17965 353 17999 387
rect 17521 279 17555 313
rect 17521 205 17555 239
rect 17521 131 17555 165
rect 17521 57 17555 91
rect 17965 279 17999 313
rect 17965 205 17999 239
rect 17965 131 17999 165
rect 17965 57 17999 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4793 -17 4827 17
rect 4867 -17 4901 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5089 -17 5123 17
rect 5237 -17 5271 17
rect 5311 -17 5345 17
rect 5385 -17 5419 17
rect 5459 -17 5493 17
rect 5533 -17 5567 17
rect 5607 -17 5641 17
rect 5681 -17 5715 17
rect 5755 -17 5789 17
rect 5829 -17 5863 17
rect 5903 -17 5937 17
rect 5977 -17 6011 17
rect 6051 -17 6085 17
rect 6199 -17 6233 17
rect 6273 -17 6307 17
rect 6347 -17 6381 17
rect 6421 -17 6455 17
rect 6495 -17 6529 17
rect 6569 -17 6603 17
rect 6643 -17 6677 17
rect 6717 -17 6751 17
rect 6791 -17 6825 17
rect 6865 -17 6899 17
rect 6939 -17 6973 17
rect 7013 -17 7047 17
rect 7161 -17 7195 17
rect 7235 -17 7269 17
rect 7309 -17 7343 17
rect 7383 -17 7417 17
rect 7457 -17 7491 17
rect 7531 -17 7565 17
rect 7605 -17 7639 17
rect 7679 -17 7713 17
rect 7827 -17 7861 17
rect 7901 -17 7935 17
rect 7975 -17 8009 17
rect 8049 -17 8083 17
rect 8123 -17 8157 17
rect 8197 -17 8231 17
rect 8271 -17 8305 17
rect 8345 -17 8379 17
rect 8419 -17 8453 17
rect 8493 -17 8527 17
rect 8567 -17 8601 17
rect 8641 -17 8675 17
rect 8789 -17 8823 17
rect 8863 -17 8897 17
rect 8937 -17 8971 17
rect 9011 -17 9045 17
rect 9085 -17 9119 17
rect 9159 -17 9193 17
rect 9233 -17 9267 17
rect 9307 -17 9341 17
rect 9381 -17 9415 17
rect 9455 -17 9489 17
rect 9529 -17 9563 17
rect 9603 -17 9637 17
rect 9751 -17 9785 17
rect 9825 -17 9859 17
rect 9899 -17 9933 17
rect 9973 -17 10007 17
rect 10047 -17 10081 17
rect 10121 -17 10155 17
rect 10195 -17 10229 17
rect 10269 -17 10303 17
rect 10417 -17 10451 17
rect 10491 -17 10525 17
rect 10565 -17 10599 17
rect 10639 -17 10673 17
rect 10713 -17 10747 17
rect 10787 -17 10821 17
rect 10861 -17 10895 17
rect 10935 -17 10969 17
rect 11009 -17 11043 17
rect 11083 -17 11117 17
rect 11157 -17 11191 17
rect 11231 -17 11265 17
rect 11379 -17 11413 17
rect 11453 -17 11487 17
rect 11527 -17 11561 17
rect 11601 -17 11635 17
rect 11675 -17 11709 17
rect 11749 -17 11783 17
rect 11823 -17 11857 17
rect 11897 -17 11931 17
rect 11971 -17 12005 17
rect 12045 -17 12079 17
rect 12119 -17 12153 17
rect 12193 -17 12227 17
rect 12341 -17 12375 17
rect 12415 -17 12449 17
rect 12489 -17 12523 17
rect 12563 -17 12597 17
rect 12637 -17 12671 17
rect 12711 -17 12745 17
rect 12785 -17 12819 17
rect 12859 -17 12893 17
rect 13007 -17 13041 17
rect 13081 -17 13115 17
rect 13155 -17 13189 17
rect 13229 -17 13263 17
rect 13303 -17 13337 17
rect 13377 -17 13411 17
rect 13451 -17 13485 17
rect 13525 -17 13559 17
rect 13599 -17 13633 17
rect 13673 -17 13707 17
rect 13747 -17 13781 17
rect 13821 -17 13855 17
rect 13969 -17 14003 17
rect 14043 -17 14077 17
rect 14117 -17 14151 17
rect 14191 -17 14225 17
rect 14265 -17 14299 17
rect 14339 -17 14373 17
rect 14413 -17 14447 17
rect 14487 -17 14521 17
rect 14561 -17 14595 17
rect 14635 -17 14669 17
rect 14709 -17 14743 17
rect 14783 -17 14817 17
rect 14931 -17 14965 17
rect 15005 -17 15039 17
rect 15079 -17 15113 17
rect 15153 -17 15187 17
rect 15227 -17 15261 17
rect 15301 -17 15335 17
rect 15375 -17 15409 17
rect 15449 -17 15483 17
rect 15597 -17 15631 17
rect 15671 -17 15705 17
rect 15745 -17 15779 17
rect 15819 -17 15853 17
rect 15893 -17 15927 17
rect 15967 -17 16001 17
rect 16041 -17 16075 17
rect 16115 -17 16149 17
rect 16263 -17 16297 17
rect 16337 -17 16371 17
rect 16411 -17 16445 17
rect 16485 -17 16519 17
rect 16559 -17 16593 17
rect 16633 -17 16667 17
rect 16707 -17 16741 17
rect 16781 -17 16815 17
rect 16929 -17 16963 17
rect 17003 -17 17037 17
rect 17077 -17 17111 17
rect 17151 -17 17185 17
rect 17225 -17 17259 17
rect 17299 -17 17333 17
rect 17373 -17 17407 17
rect 17447 -17 17481 17
rect 17595 -17 17629 17
rect 17669 -17 17703 17
rect 17743 -17 17777 17
rect 17817 -17 17851 17
rect 17891 -17 17925 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4793 1463 4827 1497
rect 4867 1463 4901 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5089 1463 5123 1497
rect 5237 1463 5271 1497
rect 5311 1463 5345 1497
rect 5385 1463 5419 1497
rect 5459 1463 5493 1497
rect 5533 1463 5567 1497
rect 5607 1463 5641 1497
rect 5681 1463 5715 1497
rect 5755 1463 5789 1497
rect 5829 1463 5863 1497
rect 5903 1463 5937 1497
rect 5977 1463 6011 1497
rect 6051 1463 6085 1497
rect 6199 1463 6233 1497
rect 6273 1463 6307 1497
rect 6347 1463 6381 1497
rect 6421 1463 6455 1497
rect 6495 1463 6529 1497
rect 6569 1463 6603 1497
rect 6643 1463 6677 1497
rect 6717 1463 6751 1497
rect 6791 1463 6825 1497
rect 6865 1463 6899 1497
rect 6939 1463 6973 1497
rect 7013 1463 7047 1497
rect 7161 1463 7195 1497
rect 7235 1463 7269 1497
rect 7309 1463 7343 1497
rect 7383 1463 7417 1497
rect 7457 1463 7491 1497
rect 7531 1463 7565 1497
rect 7605 1463 7639 1497
rect 7679 1463 7713 1497
rect 7827 1463 7861 1497
rect 7901 1463 7935 1497
rect 7975 1463 8009 1497
rect 8049 1463 8083 1497
rect 8123 1463 8157 1497
rect 8197 1463 8231 1497
rect 8271 1463 8305 1497
rect 8345 1463 8379 1497
rect 8419 1463 8453 1497
rect 8493 1463 8527 1497
rect 8567 1463 8601 1497
rect 8641 1463 8675 1497
rect 8789 1463 8823 1497
rect 8863 1463 8897 1497
rect 8937 1463 8971 1497
rect 9011 1463 9045 1497
rect 9085 1463 9119 1497
rect 9159 1463 9193 1497
rect 9233 1463 9267 1497
rect 9307 1463 9341 1497
rect 9381 1463 9415 1497
rect 9455 1463 9489 1497
rect 9529 1463 9563 1497
rect 9603 1463 9637 1497
rect 9751 1463 9785 1497
rect 9825 1463 9859 1497
rect 9899 1463 9933 1497
rect 9973 1463 10007 1497
rect 10047 1463 10081 1497
rect 10121 1463 10155 1497
rect 10195 1463 10229 1497
rect 10269 1463 10303 1497
rect 10417 1463 10451 1497
rect 10491 1463 10525 1497
rect 10565 1463 10599 1497
rect 10639 1463 10673 1497
rect 10713 1463 10747 1497
rect 10787 1463 10821 1497
rect 10861 1463 10895 1497
rect 10935 1463 10969 1497
rect 11009 1463 11043 1497
rect 11083 1463 11117 1497
rect 11157 1463 11191 1497
rect 11231 1463 11265 1497
rect 11379 1463 11413 1497
rect 11453 1463 11487 1497
rect 11527 1463 11561 1497
rect 11601 1463 11635 1497
rect 11675 1463 11709 1497
rect 11749 1463 11783 1497
rect 11823 1463 11857 1497
rect 11897 1463 11931 1497
rect 11971 1463 12005 1497
rect 12045 1463 12079 1497
rect 12119 1463 12153 1497
rect 12193 1463 12227 1497
rect 12341 1463 12375 1497
rect 12415 1463 12449 1497
rect 12489 1463 12523 1497
rect 12563 1463 12597 1497
rect 12637 1463 12671 1497
rect 12711 1463 12745 1497
rect 12785 1463 12819 1497
rect 12859 1463 12893 1497
rect 13007 1463 13041 1497
rect 13081 1463 13115 1497
rect 13155 1463 13189 1497
rect 13229 1463 13263 1497
rect 13303 1463 13337 1497
rect 13377 1463 13411 1497
rect 13451 1463 13485 1497
rect 13525 1463 13559 1497
rect 13599 1463 13633 1497
rect 13673 1463 13707 1497
rect 13747 1463 13781 1497
rect 13821 1463 13855 1497
rect 13969 1463 14003 1497
rect 14043 1463 14077 1497
rect 14117 1463 14151 1497
rect 14191 1463 14225 1497
rect 14265 1463 14299 1497
rect 14339 1463 14373 1497
rect 14413 1463 14447 1497
rect 14487 1463 14521 1497
rect 14561 1463 14595 1497
rect 14635 1463 14669 1497
rect 14709 1463 14743 1497
rect 14783 1463 14817 1497
rect 14931 1463 14965 1497
rect 15005 1463 15039 1497
rect 15079 1463 15113 1497
rect 15153 1463 15187 1497
rect 15227 1463 15261 1497
rect 15301 1463 15335 1497
rect 15375 1463 15409 1497
rect 15449 1463 15483 1497
rect 15597 1463 15631 1497
rect 15671 1463 15705 1497
rect 15745 1463 15779 1497
rect 15819 1463 15853 1497
rect 15893 1463 15927 1497
rect 15967 1463 16001 1497
rect 16041 1463 16075 1497
rect 16115 1463 16149 1497
rect 16263 1463 16297 1497
rect 16337 1463 16371 1497
rect 16411 1463 16445 1497
rect 16485 1463 16519 1497
rect 16559 1463 16593 1497
rect 16633 1463 16667 1497
rect 16707 1463 16741 1497
rect 16781 1463 16815 1497
rect 16929 1463 16963 1497
rect 17003 1463 17037 1497
rect 17077 1463 17111 1497
rect 17151 1463 17185 1497
rect 17225 1463 17259 1497
rect 17299 1463 17333 1497
rect 17373 1463 17407 1497
rect 17447 1463 17481 1497
rect 17595 1463 17629 1497
rect 17669 1463 17703 1497
rect 17743 1463 17777 1497
rect 17817 1463 17851 1497
rect 17891 1463 17925 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 945 1389 979 1423
rect 945 1315 979 1349
rect 945 1241 979 1275
rect 945 1167 979 1201
rect 945 1093 979 1127
rect 945 1019 979 1053
rect -17 945 17 979
rect 1907 1389 1941 1423
rect 1907 1315 1941 1349
rect 1907 1241 1941 1275
rect 1907 1167 1941 1201
rect 1907 1093 1941 1127
rect 1907 1019 1941 1053
rect 945 945 979 979
rect -17 871 17 905
rect 2573 1389 2607 1423
rect 2573 1315 2607 1349
rect 2573 1241 2607 1275
rect 2573 1167 2607 1201
rect 2573 1093 2607 1127
rect 2573 1019 2607 1053
rect 1907 945 1941 979
rect 945 871 979 905
rect 3535 1389 3569 1423
rect 3535 1315 3569 1349
rect 3535 1241 3569 1275
rect 3535 1167 3569 1201
rect 3535 1093 3569 1127
rect 3535 1019 3569 1053
rect 2573 945 2607 979
rect 1907 871 1941 905
rect 4497 1389 4531 1423
rect 4497 1315 4531 1349
rect 4497 1241 4531 1275
rect 4497 1167 4531 1201
rect 4497 1093 4531 1127
rect 4497 1019 4531 1053
rect 3535 945 3569 979
rect 2573 871 2607 905
rect 5163 1389 5197 1423
rect 5163 1315 5197 1349
rect 5163 1241 5197 1275
rect 5163 1167 5197 1201
rect 5163 1093 5197 1127
rect 5163 1019 5197 1053
rect 4497 945 4531 979
rect 3535 871 3569 905
rect 6125 1389 6159 1423
rect 6125 1315 6159 1349
rect 6125 1241 6159 1275
rect 6125 1167 6159 1201
rect 6125 1093 6159 1127
rect 6125 1019 6159 1053
rect 5163 945 5197 979
rect 4497 871 4531 905
rect 7087 1389 7121 1423
rect 7087 1315 7121 1349
rect 7087 1241 7121 1275
rect 7087 1167 7121 1201
rect 7087 1093 7121 1127
rect 7087 1019 7121 1053
rect 6125 945 6159 979
rect 5163 871 5197 905
rect 7753 1389 7787 1423
rect 7753 1315 7787 1349
rect 7753 1241 7787 1275
rect 7753 1167 7787 1201
rect 7753 1093 7787 1127
rect 7753 1019 7787 1053
rect 7087 945 7121 979
rect 6125 871 6159 905
rect 8715 1389 8749 1423
rect 8715 1315 8749 1349
rect 8715 1241 8749 1275
rect 8715 1167 8749 1201
rect 8715 1093 8749 1127
rect 8715 1019 8749 1053
rect 7753 945 7787 979
rect 7087 871 7121 905
rect 9677 1389 9711 1423
rect 9677 1315 9711 1349
rect 9677 1241 9711 1275
rect 9677 1167 9711 1201
rect 9677 1093 9711 1127
rect 9677 1019 9711 1053
rect 8715 945 8749 979
rect 7753 871 7787 905
rect 10343 1389 10377 1423
rect 10343 1315 10377 1349
rect 10343 1241 10377 1275
rect 10343 1167 10377 1201
rect 10343 1093 10377 1127
rect 10343 1019 10377 1053
rect 9677 945 9711 979
rect 8715 871 8749 905
rect 11305 1389 11339 1423
rect 11305 1315 11339 1349
rect 11305 1241 11339 1275
rect 11305 1167 11339 1201
rect 11305 1093 11339 1127
rect 11305 1019 11339 1053
rect 10343 945 10377 979
rect 9677 871 9711 905
rect 12267 1389 12301 1423
rect 12267 1315 12301 1349
rect 12267 1241 12301 1275
rect 12267 1167 12301 1201
rect 12267 1093 12301 1127
rect 12267 1019 12301 1053
rect 11305 945 11339 979
rect 10343 871 10377 905
rect 12933 1389 12967 1423
rect 12933 1315 12967 1349
rect 12933 1241 12967 1275
rect 12933 1167 12967 1201
rect 12933 1093 12967 1127
rect 12933 1019 12967 1053
rect 12267 945 12301 979
rect 11305 871 11339 905
rect 13895 1389 13929 1423
rect 13895 1315 13929 1349
rect 13895 1241 13929 1275
rect 13895 1167 13929 1201
rect 13895 1093 13929 1127
rect 13895 1019 13929 1053
rect 12933 945 12967 979
rect 12267 871 12301 905
rect 14857 1389 14891 1423
rect 14857 1315 14891 1349
rect 14857 1241 14891 1275
rect 14857 1167 14891 1201
rect 14857 1093 14891 1127
rect 14857 1019 14891 1053
rect 13895 945 13929 979
rect 12933 871 12967 905
rect 15523 1389 15557 1423
rect 15523 1315 15557 1349
rect 15523 1241 15557 1275
rect 15523 1167 15557 1201
rect 15523 1093 15557 1127
rect 15523 1019 15557 1053
rect 14857 945 14891 979
rect 13895 871 13929 905
rect 16189 1389 16223 1423
rect 16189 1315 16223 1349
rect 16189 1241 16223 1275
rect 16189 1167 16223 1201
rect 16189 1093 16223 1127
rect 16189 1019 16223 1053
rect 15523 945 15557 979
rect 14857 871 14891 905
rect 16855 1389 16889 1423
rect 16855 1315 16889 1349
rect 16855 1241 16889 1275
rect 16855 1167 16889 1201
rect 16855 1093 16889 1127
rect 16855 1019 16889 1053
rect 16189 945 16223 979
rect 15523 871 15557 905
rect 17521 1389 17555 1423
rect 17521 1315 17555 1349
rect 17521 1241 17555 1275
rect 17521 1167 17555 1201
rect 17521 1093 17555 1127
rect 17521 1019 17555 1053
rect 16855 945 16889 979
rect 16189 871 16223 905
rect 17965 1389 17999 1423
rect 17965 1315 17999 1349
rect 17965 1241 17999 1275
rect 17965 1167 17999 1201
rect 17965 1093 17999 1127
rect 17965 1019 17999 1053
rect 17521 945 17555 979
rect 16855 871 16889 905
rect 17965 945 17999 979
rect 17521 871 17555 905
rect 17965 871 17999 905
<< poly >>
rect 247 1404 277 1430
rect 335 1404 365 1430
rect 423 1404 453 1430
rect 511 1404 541 1430
rect 599 1404 629 1430
rect 687 1404 717 1430
rect 1209 1404 1239 1430
rect 1297 1404 1327 1430
rect 1385 1404 1415 1430
rect 1473 1404 1503 1430
rect 1561 1404 1591 1430
rect 1649 1404 1679 1430
rect 247 973 277 1004
rect 335 973 365 1004
rect 423 973 453 1004
rect 511 973 541 1004
rect 195 957 365 973
rect 195 923 205 957
rect 239 943 365 957
rect 417 957 541 973
rect 239 923 249 943
rect 195 907 249 923
rect 417 923 427 957
rect 461 943 541 957
rect 599 973 629 1004
rect 687 973 717 1004
rect 599 957 717 973
rect 599 943 649 957
rect 461 923 471 943
rect 417 907 471 923
rect 639 923 649 943
rect 683 943 717 957
rect 2111 1404 2141 1430
rect 2199 1404 2229 1430
rect 2287 1404 2317 1430
rect 2375 1404 2405 1430
rect 1209 973 1239 1004
rect 1297 973 1327 1004
rect 1385 973 1415 1004
rect 1473 973 1503 1004
rect 683 923 693 943
rect 639 907 693 923
rect 1157 957 1327 973
rect 1157 923 1167 957
rect 1201 943 1327 957
rect 1379 957 1503 973
rect 1201 923 1211 943
rect 1157 907 1211 923
rect 1379 923 1389 957
rect 1423 943 1503 957
rect 1561 973 1591 1004
rect 1649 973 1679 1004
rect 1561 957 1679 973
rect 1561 943 1611 957
rect 1423 923 1433 943
rect 1379 907 1433 923
rect 1601 923 1611 943
rect 1645 943 1679 957
rect 2837 1404 2867 1430
rect 2925 1404 2955 1430
rect 3013 1404 3043 1430
rect 3101 1404 3131 1430
rect 3189 1404 3219 1430
rect 3277 1404 3307 1430
rect 1645 923 1655 943
rect 1601 907 1655 923
rect 2111 973 2141 1004
rect 2199 973 2229 1004
rect 2287 973 2317 1004
rect 2375 973 2405 1004
rect 2111 957 2229 973
rect 2111 943 2129 957
rect 2119 923 2129 943
rect 2163 943 2229 957
rect 2273 957 2405 973
rect 2163 923 2173 943
rect 2119 907 2173 923
rect 2273 923 2283 957
rect 2317 943 2405 957
rect 3799 1404 3829 1430
rect 3887 1404 3917 1430
rect 3975 1404 4005 1430
rect 4063 1404 4093 1430
rect 4151 1404 4181 1430
rect 4239 1404 4269 1430
rect 2837 973 2867 1004
rect 2925 973 2955 1004
rect 3013 973 3043 1004
rect 3101 973 3131 1004
rect 2317 923 2327 943
rect 2273 907 2327 923
rect 2785 957 2955 973
rect 2785 923 2795 957
rect 2829 943 2955 957
rect 3007 957 3131 973
rect 2829 923 2839 943
rect 2785 907 2839 923
rect 3007 923 3017 957
rect 3051 943 3131 957
rect 3189 973 3219 1004
rect 3277 973 3307 1004
rect 3189 957 3307 973
rect 3189 943 3239 957
rect 3051 923 3061 943
rect 3007 907 3061 923
rect 3229 923 3239 943
rect 3273 943 3307 957
rect 4701 1404 4731 1430
rect 4789 1404 4819 1430
rect 4877 1404 4907 1430
rect 4965 1404 4995 1430
rect 3799 973 3829 1004
rect 3887 973 3917 1004
rect 3975 973 4005 1004
rect 4063 973 4093 1004
rect 3273 923 3283 943
rect 3229 907 3283 923
rect 3747 957 3917 973
rect 3747 923 3757 957
rect 3791 943 3917 957
rect 3969 957 4093 973
rect 3791 923 3801 943
rect 3747 907 3801 923
rect 3969 923 3979 957
rect 4013 943 4093 957
rect 4151 973 4181 1004
rect 4239 973 4269 1004
rect 4151 957 4269 973
rect 4151 943 4201 957
rect 4013 923 4023 943
rect 3969 907 4023 923
rect 4191 923 4201 943
rect 4235 943 4269 957
rect 5427 1404 5457 1430
rect 5515 1404 5545 1430
rect 5603 1404 5633 1430
rect 5691 1404 5721 1430
rect 5779 1404 5809 1430
rect 5867 1404 5897 1430
rect 4235 923 4245 943
rect 4191 907 4245 923
rect 4701 973 4731 1004
rect 4789 973 4819 1004
rect 4877 973 4907 1004
rect 4965 973 4995 1004
rect 4701 957 4819 973
rect 4701 943 4719 957
rect 4709 923 4719 943
rect 4753 943 4819 957
rect 4863 957 4995 973
rect 4753 923 4763 943
rect 4709 907 4763 923
rect 4863 923 4873 957
rect 4907 943 4995 957
rect 6389 1404 6419 1430
rect 6477 1404 6507 1430
rect 6565 1404 6595 1430
rect 6653 1404 6683 1430
rect 6741 1404 6771 1430
rect 6829 1404 6859 1430
rect 5427 973 5457 1004
rect 5515 973 5545 1004
rect 5603 973 5633 1004
rect 5691 973 5721 1004
rect 4907 923 4917 943
rect 4863 907 4917 923
rect 5375 957 5545 973
rect 5375 923 5385 957
rect 5419 943 5545 957
rect 5597 957 5721 973
rect 5419 923 5429 943
rect 5375 907 5429 923
rect 5597 923 5607 957
rect 5641 943 5721 957
rect 5779 973 5809 1004
rect 5867 973 5897 1004
rect 5779 957 5897 973
rect 5779 943 5829 957
rect 5641 923 5651 943
rect 5597 907 5651 923
rect 5819 923 5829 943
rect 5863 943 5897 957
rect 7291 1404 7321 1430
rect 7379 1404 7409 1430
rect 7467 1404 7497 1430
rect 7555 1404 7585 1430
rect 6389 973 6419 1004
rect 6477 973 6507 1004
rect 6565 973 6595 1004
rect 6653 973 6683 1004
rect 5863 923 5873 943
rect 5819 907 5873 923
rect 6337 957 6507 973
rect 6337 923 6347 957
rect 6381 943 6507 957
rect 6559 957 6683 973
rect 6381 923 6391 943
rect 6337 907 6391 923
rect 6559 923 6569 957
rect 6603 943 6683 957
rect 6741 973 6771 1004
rect 6829 973 6859 1004
rect 6741 957 6859 973
rect 6741 943 6791 957
rect 6603 923 6613 943
rect 6559 907 6613 923
rect 6781 923 6791 943
rect 6825 943 6859 957
rect 8017 1404 8047 1430
rect 8105 1404 8135 1430
rect 8193 1404 8223 1430
rect 8281 1404 8311 1430
rect 8369 1404 8399 1430
rect 8457 1404 8487 1430
rect 6825 923 6835 943
rect 6781 907 6835 923
rect 7291 973 7321 1004
rect 7379 973 7409 1004
rect 7467 973 7497 1004
rect 7555 973 7585 1004
rect 7291 957 7409 973
rect 7291 943 7309 957
rect 7299 923 7309 943
rect 7343 943 7409 957
rect 7453 957 7585 973
rect 7343 923 7353 943
rect 7299 907 7353 923
rect 7453 923 7463 957
rect 7497 943 7585 957
rect 8979 1404 9009 1430
rect 9067 1404 9097 1430
rect 9155 1404 9185 1430
rect 9243 1404 9273 1430
rect 9331 1404 9361 1430
rect 9419 1404 9449 1430
rect 8017 973 8047 1004
rect 8105 973 8135 1004
rect 8193 973 8223 1004
rect 8281 973 8311 1004
rect 7497 923 7507 943
rect 7453 907 7507 923
rect 7965 957 8135 973
rect 7965 923 7975 957
rect 8009 943 8135 957
rect 8187 957 8311 973
rect 8009 923 8019 943
rect 7965 907 8019 923
rect 8187 923 8197 957
rect 8231 943 8311 957
rect 8369 973 8399 1004
rect 8457 973 8487 1004
rect 8369 957 8487 973
rect 8369 943 8419 957
rect 8231 923 8241 943
rect 8187 907 8241 923
rect 8409 923 8419 943
rect 8453 943 8487 957
rect 9881 1404 9911 1430
rect 9969 1404 9999 1430
rect 10057 1404 10087 1430
rect 10145 1404 10175 1430
rect 8979 973 9009 1004
rect 9067 973 9097 1004
rect 9155 973 9185 1004
rect 9243 973 9273 1004
rect 8453 923 8463 943
rect 8409 907 8463 923
rect 8927 957 9097 973
rect 8927 923 8937 957
rect 8971 943 9097 957
rect 9149 957 9273 973
rect 8971 923 8981 943
rect 8927 907 8981 923
rect 9149 923 9159 957
rect 9193 943 9273 957
rect 9331 973 9361 1004
rect 9419 973 9449 1004
rect 9331 957 9449 973
rect 9331 943 9381 957
rect 9193 923 9203 943
rect 9149 907 9203 923
rect 9371 923 9381 943
rect 9415 943 9449 957
rect 10607 1404 10637 1430
rect 10695 1404 10725 1430
rect 10783 1404 10813 1430
rect 10871 1404 10901 1430
rect 10959 1404 10989 1430
rect 11047 1404 11077 1430
rect 9415 923 9425 943
rect 9371 907 9425 923
rect 9881 973 9911 1004
rect 9969 973 9999 1004
rect 10057 973 10087 1004
rect 10145 973 10175 1004
rect 9881 957 9999 973
rect 9881 943 9899 957
rect 9889 923 9899 943
rect 9933 943 9999 957
rect 10043 957 10175 973
rect 9933 923 9943 943
rect 9889 907 9943 923
rect 10043 923 10053 957
rect 10087 943 10175 957
rect 11569 1404 11599 1430
rect 11657 1404 11687 1430
rect 11745 1404 11775 1430
rect 11833 1404 11863 1430
rect 11921 1404 11951 1430
rect 12009 1404 12039 1430
rect 10607 973 10637 1004
rect 10695 973 10725 1004
rect 10783 973 10813 1004
rect 10871 973 10901 1004
rect 10087 923 10097 943
rect 10043 907 10097 923
rect 10555 957 10725 973
rect 10555 923 10565 957
rect 10599 943 10725 957
rect 10777 957 10901 973
rect 10599 923 10609 943
rect 10555 907 10609 923
rect 10777 923 10787 957
rect 10821 943 10901 957
rect 10959 973 10989 1004
rect 11047 973 11077 1004
rect 10959 957 11077 973
rect 10959 943 11009 957
rect 10821 923 10831 943
rect 10777 907 10831 923
rect 10999 923 11009 943
rect 11043 943 11077 957
rect 12471 1404 12501 1430
rect 12559 1404 12589 1430
rect 12647 1404 12677 1430
rect 12735 1404 12765 1430
rect 11569 973 11599 1004
rect 11657 973 11687 1004
rect 11745 973 11775 1004
rect 11833 973 11863 1004
rect 11043 923 11053 943
rect 10999 907 11053 923
rect 11517 957 11687 973
rect 11517 923 11527 957
rect 11561 943 11687 957
rect 11739 957 11863 973
rect 11561 923 11571 943
rect 11517 907 11571 923
rect 11739 923 11749 957
rect 11783 943 11863 957
rect 11921 973 11951 1004
rect 12009 973 12039 1004
rect 11921 957 12039 973
rect 11921 943 11971 957
rect 11783 923 11793 943
rect 11739 907 11793 923
rect 11961 923 11971 943
rect 12005 943 12039 957
rect 13197 1404 13227 1430
rect 13285 1404 13315 1430
rect 13373 1404 13403 1430
rect 13461 1404 13491 1430
rect 13549 1404 13579 1430
rect 13637 1404 13667 1430
rect 12005 923 12015 943
rect 11961 907 12015 923
rect 12471 973 12501 1004
rect 12559 973 12589 1004
rect 12647 973 12677 1004
rect 12735 973 12765 1004
rect 12471 957 12589 973
rect 12471 943 12489 957
rect 12479 923 12489 943
rect 12523 943 12589 957
rect 12633 957 12765 973
rect 12523 923 12533 943
rect 12479 907 12533 923
rect 12633 923 12643 957
rect 12677 943 12765 957
rect 14159 1404 14189 1430
rect 14247 1404 14277 1430
rect 14335 1404 14365 1430
rect 14423 1404 14453 1430
rect 14511 1404 14541 1430
rect 14599 1404 14629 1430
rect 13197 973 13227 1004
rect 13285 973 13315 1004
rect 13373 973 13403 1004
rect 13461 973 13491 1004
rect 12677 923 12687 943
rect 12633 907 12687 923
rect 13145 957 13315 973
rect 13145 923 13155 957
rect 13189 943 13315 957
rect 13367 957 13491 973
rect 13189 923 13199 943
rect 13145 907 13199 923
rect 13367 923 13377 957
rect 13411 943 13491 957
rect 13549 973 13579 1004
rect 13637 973 13667 1004
rect 13549 957 13667 973
rect 13549 943 13599 957
rect 13411 923 13421 943
rect 13367 907 13421 923
rect 13589 923 13599 943
rect 13633 943 13667 957
rect 15061 1404 15091 1430
rect 15149 1404 15179 1430
rect 15237 1404 15267 1430
rect 15325 1404 15355 1430
rect 14159 973 14189 1004
rect 14247 973 14277 1004
rect 14335 973 14365 1004
rect 14423 973 14453 1004
rect 13633 923 13643 943
rect 13589 907 13643 923
rect 14107 957 14277 973
rect 14107 923 14117 957
rect 14151 943 14277 957
rect 14329 957 14453 973
rect 14151 923 14161 943
rect 14107 907 14161 923
rect 14329 923 14339 957
rect 14373 943 14453 957
rect 14511 973 14541 1004
rect 14599 973 14629 1004
rect 14511 957 14629 973
rect 14511 943 14561 957
rect 14373 923 14383 943
rect 14329 907 14383 923
rect 14551 923 14561 943
rect 14595 943 14629 957
rect 15727 1405 15757 1431
rect 15815 1405 15845 1431
rect 15903 1405 15933 1431
rect 15991 1405 16021 1431
rect 14595 923 14605 943
rect 14551 907 14605 923
rect 15061 973 15091 1004
rect 15149 973 15179 1004
rect 15237 973 15267 1004
rect 15325 973 15355 1004
rect 15061 957 15179 973
rect 15061 943 15079 957
rect 15069 923 15079 943
rect 15113 943 15179 957
rect 15223 957 15355 973
rect 15113 923 15123 943
rect 15069 907 15123 923
rect 15223 923 15233 957
rect 15267 943 15355 957
rect 16391 1405 16421 1431
rect 16479 1405 16509 1431
rect 16567 1405 16597 1431
rect 16655 1405 16685 1431
rect 15727 974 15757 1005
rect 15815 974 15845 1005
rect 15903 974 15933 1005
rect 15991 974 16021 1005
rect 15267 923 15277 943
rect 15223 907 15277 923
rect 15661 958 15845 974
rect 15661 924 15671 958
rect 15705 944 15845 958
rect 15891 958 16021 974
rect 15705 924 15715 944
rect 15661 908 15715 924
rect 15891 924 15901 958
rect 15935 944 16021 958
rect 17059 1405 17089 1431
rect 17147 1405 17177 1431
rect 17235 1405 17265 1431
rect 17323 1405 17353 1431
rect 15935 924 15945 944
rect 15891 908 15945 924
rect 16391 974 16421 1005
rect 16479 974 16509 1005
rect 16391 958 16509 974
rect 16391 944 16411 958
rect 16401 924 16411 944
rect 16445 944 16509 958
rect 16567 974 16597 1005
rect 16655 974 16685 1005
rect 17702 1404 17732 1430
rect 17790 1404 17820 1430
rect 16567 958 16751 974
rect 16567 944 16707 958
rect 16445 924 16455 944
rect 16401 908 16455 924
rect 16697 924 16707 944
rect 16741 924 16751 958
rect 16697 908 16751 924
rect 17059 974 17089 1005
rect 17147 974 17177 1005
rect 17235 974 17265 1005
rect 17323 974 17353 1005
rect 16993 958 17177 974
rect 16993 924 17003 958
rect 17037 944 17177 958
rect 17219 958 17353 974
rect 17037 924 17047 944
rect 16993 908 17047 924
rect 17219 924 17229 958
rect 17263 944 17353 958
rect 17702 973 17732 1004
rect 17790 973 17820 1004
rect 17263 924 17273 944
rect 17219 908 17273 924
rect 17659 957 17820 973
rect 17659 923 17669 957
rect 17703 943 17820 957
rect 17703 923 17713 943
rect 17659 907 17713 923
rect 195 433 249 449
rect 195 413 205 433
rect 147 399 205 413
rect 239 399 249 433
rect 147 383 249 399
rect 417 433 471 449
rect 417 399 427 433
rect 461 413 471 433
rect 639 433 693 449
rect 461 399 477 413
rect 417 383 477 399
rect 639 399 649 433
rect 683 399 693 433
rect 639 383 693 399
rect 1157 433 1211 449
rect 1157 413 1167 433
rect 147 351 177 383
rect 447 351 477 383
rect 649 351 679 383
rect 1109 399 1167 413
rect 1201 399 1211 433
rect 1109 383 1211 399
rect 1379 433 1433 449
rect 1379 399 1389 433
rect 1423 413 1433 433
rect 1601 433 1655 449
rect 1423 399 1439 413
rect 1379 383 1439 399
rect 1601 399 1611 433
rect 1645 399 1655 433
rect 1601 383 1655 399
rect 2119 433 2173 449
rect 2119 413 2129 433
rect 1109 351 1139 383
rect 1409 351 1439 383
rect 1611 351 1641 383
rect 2092 399 2129 413
rect 2163 399 2173 433
rect 2092 383 2173 399
rect 2267 433 2321 449
rect 2267 399 2277 433
rect 2311 399 2321 433
rect 2267 383 2321 399
rect 2785 433 2839 449
rect 2785 413 2795 433
rect 2092 349 2122 383
rect 2286 349 2316 383
rect 2737 399 2795 413
rect 2829 399 2839 433
rect 2737 383 2839 399
rect 3007 433 3061 449
rect 3007 399 3017 433
rect 3051 413 3061 433
rect 3229 433 3283 449
rect 3051 399 3067 413
rect 3007 383 3067 399
rect 3229 399 3239 433
rect 3273 399 3283 433
rect 3229 383 3283 399
rect 3747 433 3801 449
rect 3747 413 3757 433
rect 2737 351 2767 383
rect 3037 351 3067 383
rect 3239 351 3269 383
rect 3699 399 3757 413
rect 3791 399 3801 433
rect 3699 383 3801 399
rect 3969 433 4023 449
rect 3969 399 3979 433
rect 4013 413 4023 433
rect 4191 433 4245 449
rect 4013 399 4029 413
rect 3969 383 4029 399
rect 4191 399 4201 433
rect 4235 399 4245 433
rect 4191 383 4245 399
rect 4709 433 4763 449
rect 4709 413 4719 433
rect 3699 351 3729 383
rect 3999 351 4029 383
rect 4201 351 4231 383
rect 4682 399 4719 413
rect 4753 399 4763 433
rect 4682 383 4763 399
rect 4857 433 4911 449
rect 4857 399 4867 433
rect 4901 399 4911 433
rect 4857 383 4911 399
rect 5375 433 5429 449
rect 5375 413 5385 433
rect 4682 349 4712 383
rect 4876 349 4906 383
rect 5327 399 5385 413
rect 5419 399 5429 433
rect 5327 383 5429 399
rect 5597 433 5651 449
rect 5597 399 5607 433
rect 5641 413 5651 433
rect 5819 433 5873 449
rect 5641 399 5657 413
rect 5597 383 5657 399
rect 5819 399 5829 433
rect 5863 399 5873 433
rect 5819 383 5873 399
rect 6337 433 6391 449
rect 6337 413 6347 433
rect 5327 351 5357 383
rect 5627 351 5657 383
rect 5829 351 5859 383
rect 6289 399 6347 413
rect 6381 399 6391 433
rect 6289 383 6391 399
rect 6559 433 6613 449
rect 6559 399 6569 433
rect 6603 413 6613 433
rect 6781 433 6835 449
rect 6603 399 6619 413
rect 6559 383 6619 399
rect 6781 399 6791 433
rect 6825 399 6835 433
rect 6781 383 6835 399
rect 7299 433 7353 449
rect 7299 413 7309 433
rect 6289 351 6319 383
rect 6589 351 6619 383
rect 6791 351 6821 383
rect 7272 399 7309 413
rect 7343 399 7353 433
rect 7272 383 7353 399
rect 7447 433 7501 449
rect 7447 399 7457 433
rect 7491 399 7501 433
rect 7447 383 7501 399
rect 7965 433 8019 449
rect 7965 413 7975 433
rect 7272 349 7302 383
rect 7466 349 7496 383
rect 7917 399 7975 413
rect 8009 399 8019 433
rect 7917 383 8019 399
rect 8187 433 8241 449
rect 8187 399 8197 433
rect 8231 413 8241 433
rect 8409 433 8463 449
rect 8231 399 8247 413
rect 8187 383 8247 399
rect 8409 399 8419 433
rect 8453 399 8463 433
rect 8409 383 8463 399
rect 8927 433 8981 449
rect 8927 413 8937 433
rect 7917 351 7947 383
rect 8217 351 8247 383
rect 8419 351 8449 383
rect 8879 399 8937 413
rect 8971 399 8981 433
rect 8879 383 8981 399
rect 9149 433 9203 449
rect 9149 399 9159 433
rect 9193 413 9203 433
rect 9371 433 9425 449
rect 9193 399 9209 413
rect 9149 383 9209 399
rect 9371 399 9381 433
rect 9415 399 9425 433
rect 9371 383 9425 399
rect 9889 433 9943 449
rect 9889 413 9899 433
rect 8879 351 8909 383
rect 9179 351 9209 383
rect 9381 351 9411 383
rect 9862 399 9899 413
rect 9933 399 9943 433
rect 9862 383 9943 399
rect 10037 433 10091 449
rect 10037 399 10047 433
rect 10081 399 10091 433
rect 10037 383 10091 399
rect 10555 433 10609 449
rect 10555 413 10565 433
rect 9862 349 9892 383
rect 10056 349 10086 383
rect 10507 399 10565 413
rect 10599 399 10609 433
rect 10507 383 10609 399
rect 10777 433 10831 449
rect 10777 399 10787 433
rect 10821 413 10831 433
rect 10999 433 11053 449
rect 10821 399 10837 413
rect 10777 383 10837 399
rect 10999 399 11009 433
rect 11043 399 11053 433
rect 10999 383 11053 399
rect 11517 433 11571 449
rect 11517 413 11527 433
rect 10507 351 10537 383
rect 10807 351 10837 383
rect 11009 351 11039 383
rect 11469 399 11527 413
rect 11561 399 11571 433
rect 11469 383 11571 399
rect 11739 433 11793 449
rect 11739 399 11749 433
rect 11783 413 11793 433
rect 11961 433 12015 449
rect 11783 399 11799 413
rect 11739 383 11799 399
rect 11961 399 11971 433
rect 12005 399 12015 433
rect 11961 383 12015 399
rect 12479 433 12533 449
rect 12479 413 12489 433
rect 11469 351 11499 383
rect 11769 351 11799 383
rect 11971 351 12001 383
rect 12452 399 12489 413
rect 12523 399 12533 433
rect 12452 383 12533 399
rect 12627 433 12681 449
rect 12627 399 12637 433
rect 12671 399 12681 433
rect 12627 383 12681 399
rect 13145 433 13199 449
rect 13145 413 13155 433
rect 12452 349 12482 383
rect 12646 349 12676 383
rect 13097 399 13155 413
rect 13189 399 13199 433
rect 13097 383 13199 399
rect 13367 433 13421 449
rect 13367 399 13377 433
rect 13411 413 13421 433
rect 13589 433 13643 449
rect 13411 399 13427 413
rect 13367 383 13427 399
rect 13589 399 13599 433
rect 13633 399 13643 433
rect 13589 383 13643 399
rect 14107 433 14161 449
rect 14107 413 14117 433
rect 13097 351 13127 383
rect 13397 351 13427 383
rect 13599 351 13629 383
rect 14059 399 14117 413
rect 14151 399 14161 433
rect 14059 383 14161 399
rect 14329 433 14383 449
rect 14329 399 14339 433
rect 14373 413 14383 433
rect 14551 433 14605 449
rect 14373 399 14389 413
rect 14329 383 14389 399
rect 14551 399 14561 433
rect 14595 399 14605 433
rect 14551 383 14605 399
rect 15069 433 15123 449
rect 15069 413 15079 433
rect 14059 351 14089 383
rect 14359 351 14389 383
rect 14561 351 14591 383
rect 15042 399 15079 413
rect 15113 399 15123 433
rect 15042 383 15123 399
rect 15217 433 15271 449
rect 15217 399 15227 433
rect 15261 399 15271 433
rect 15217 383 15271 399
rect 15042 349 15072 383
rect 15236 349 15266 383
rect 15661 433 15715 449
rect 15661 399 15671 433
rect 15705 413 15715 433
rect 15883 433 15937 449
rect 15705 399 15738 413
rect 15661 383 15738 399
rect 15883 399 15893 433
rect 15927 399 15937 433
rect 15883 383 15937 399
rect 16401 433 16455 449
rect 16401 413 16411 433
rect 15708 349 15738 383
rect 15902 349 15932 383
rect 16374 399 16411 413
rect 16445 399 16455 433
rect 16697 433 16751 449
rect 16697 413 16707 433
rect 16374 383 16455 399
rect 16674 399 16707 413
rect 16741 399 16751 433
rect 16674 383 16751 399
rect 16374 349 16404 383
rect 16674 349 16704 383
rect 16993 433 17047 449
rect 16993 399 17003 433
rect 17037 413 17047 433
rect 17215 433 17269 449
rect 17037 399 17070 413
rect 16993 383 17070 399
rect 17215 399 17225 433
rect 17259 399 17269 433
rect 17215 383 17269 399
rect 17040 349 17070 383
rect 17234 349 17264 383
rect 17659 434 17713 450
rect 17659 400 17669 434
rect 17703 413 17713 434
rect 17703 400 17723 413
rect 17659 384 17723 400
rect 17693 350 17723 384
<< polycont >>
rect 205 923 239 957
rect 427 923 461 957
rect 649 923 683 957
rect 1167 923 1201 957
rect 1389 923 1423 957
rect 1611 923 1645 957
rect 2129 923 2163 957
rect 2283 923 2317 957
rect 2795 923 2829 957
rect 3017 923 3051 957
rect 3239 923 3273 957
rect 3757 923 3791 957
rect 3979 923 4013 957
rect 4201 923 4235 957
rect 4719 923 4753 957
rect 4873 923 4907 957
rect 5385 923 5419 957
rect 5607 923 5641 957
rect 5829 923 5863 957
rect 6347 923 6381 957
rect 6569 923 6603 957
rect 6791 923 6825 957
rect 7309 923 7343 957
rect 7463 923 7497 957
rect 7975 923 8009 957
rect 8197 923 8231 957
rect 8419 923 8453 957
rect 8937 923 8971 957
rect 9159 923 9193 957
rect 9381 923 9415 957
rect 9899 923 9933 957
rect 10053 923 10087 957
rect 10565 923 10599 957
rect 10787 923 10821 957
rect 11009 923 11043 957
rect 11527 923 11561 957
rect 11749 923 11783 957
rect 11971 923 12005 957
rect 12489 923 12523 957
rect 12643 923 12677 957
rect 13155 923 13189 957
rect 13377 923 13411 957
rect 13599 923 13633 957
rect 14117 923 14151 957
rect 14339 923 14373 957
rect 14561 923 14595 957
rect 15079 923 15113 957
rect 15233 923 15267 957
rect 15671 924 15705 958
rect 15901 924 15935 958
rect 16411 924 16445 958
rect 16707 924 16741 958
rect 17003 924 17037 958
rect 17229 924 17263 958
rect 17669 923 17703 957
rect 205 399 239 433
rect 427 399 461 433
rect 649 399 683 433
rect 1167 399 1201 433
rect 1389 399 1423 433
rect 1611 399 1645 433
rect 2129 399 2163 433
rect 2277 399 2311 433
rect 2795 399 2829 433
rect 3017 399 3051 433
rect 3239 399 3273 433
rect 3757 399 3791 433
rect 3979 399 4013 433
rect 4201 399 4235 433
rect 4719 399 4753 433
rect 4867 399 4901 433
rect 5385 399 5419 433
rect 5607 399 5641 433
rect 5829 399 5863 433
rect 6347 399 6381 433
rect 6569 399 6603 433
rect 6791 399 6825 433
rect 7309 399 7343 433
rect 7457 399 7491 433
rect 7975 399 8009 433
rect 8197 399 8231 433
rect 8419 399 8453 433
rect 8937 399 8971 433
rect 9159 399 9193 433
rect 9381 399 9415 433
rect 9899 399 9933 433
rect 10047 399 10081 433
rect 10565 399 10599 433
rect 10787 399 10821 433
rect 11009 399 11043 433
rect 11527 399 11561 433
rect 11749 399 11783 433
rect 11971 399 12005 433
rect 12489 399 12523 433
rect 12637 399 12671 433
rect 13155 399 13189 433
rect 13377 399 13411 433
rect 13599 399 13633 433
rect 14117 399 14151 433
rect 14339 399 14373 433
rect 14561 399 14595 433
rect 15079 399 15113 433
rect 15227 399 15261 433
rect 15671 399 15705 433
rect 15893 399 15927 433
rect 16411 399 16445 433
rect 16707 399 16741 433
rect 17003 399 17037 433
rect 17225 399 17259 433
rect 17669 400 17703 434
<< locali >>
rect -34 1497 18016 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5533 1497
rect 5567 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5755 1497
rect 5789 1463 5829 1497
rect 5863 1463 5903 1497
rect 5937 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6199 1497
rect 6233 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6495 1497
rect 6529 1463 6569 1497
rect 6603 1463 6643 1497
rect 6677 1463 6717 1497
rect 6751 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7161 1497
rect 7195 1463 7235 1497
rect 7269 1463 7309 1497
rect 7343 1463 7383 1497
rect 7417 1463 7457 1497
rect 7491 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7679 1497
rect 7713 1463 7827 1497
rect 7861 1463 7901 1497
rect 7935 1463 7975 1497
rect 8009 1463 8049 1497
rect 8083 1463 8123 1497
rect 8157 1463 8197 1497
rect 8231 1463 8271 1497
rect 8305 1463 8345 1497
rect 8379 1463 8419 1497
rect 8453 1463 8493 1497
rect 8527 1463 8567 1497
rect 8601 1463 8641 1497
rect 8675 1463 8789 1497
rect 8823 1463 8863 1497
rect 8897 1463 8937 1497
rect 8971 1463 9011 1497
rect 9045 1463 9085 1497
rect 9119 1463 9159 1497
rect 9193 1463 9233 1497
rect 9267 1463 9307 1497
rect 9341 1463 9381 1497
rect 9415 1463 9455 1497
rect 9489 1463 9529 1497
rect 9563 1463 9603 1497
rect 9637 1463 9751 1497
rect 9785 1463 9825 1497
rect 9859 1463 9899 1497
rect 9933 1463 9973 1497
rect 10007 1463 10047 1497
rect 10081 1463 10121 1497
rect 10155 1463 10195 1497
rect 10229 1463 10269 1497
rect 10303 1463 10417 1497
rect 10451 1463 10491 1497
rect 10525 1463 10565 1497
rect 10599 1463 10639 1497
rect 10673 1463 10713 1497
rect 10747 1463 10787 1497
rect 10821 1463 10861 1497
rect 10895 1463 10935 1497
rect 10969 1463 11009 1497
rect 11043 1463 11083 1497
rect 11117 1463 11157 1497
rect 11191 1463 11231 1497
rect 11265 1463 11379 1497
rect 11413 1463 11453 1497
rect 11487 1463 11527 1497
rect 11561 1463 11601 1497
rect 11635 1463 11675 1497
rect 11709 1463 11749 1497
rect 11783 1463 11823 1497
rect 11857 1463 11897 1497
rect 11931 1463 11971 1497
rect 12005 1463 12045 1497
rect 12079 1463 12119 1497
rect 12153 1463 12193 1497
rect 12227 1463 12341 1497
rect 12375 1463 12415 1497
rect 12449 1463 12489 1497
rect 12523 1463 12563 1497
rect 12597 1463 12637 1497
rect 12671 1463 12711 1497
rect 12745 1463 12785 1497
rect 12819 1463 12859 1497
rect 12893 1463 13007 1497
rect 13041 1463 13081 1497
rect 13115 1463 13155 1497
rect 13189 1463 13229 1497
rect 13263 1463 13303 1497
rect 13337 1463 13377 1497
rect 13411 1463 13451 1497
rect 13485 1463 13525 1497
rect 13559 1463 13599 1497
rect 13633 1463 13673 1497
rect 13707 1463 13747 1497
rect 13781 1463 13821 1497
rect 13855 1463 13969 1497
rect 14003 1463 14043 1497
rect 14077 1463 14117 1497
rect 14151 1463 14191 1497
rect 14225 1463 14265 1497
rect 14299 1463 14339 1497
rect 14373 1463 14413 1497
rect 14447 1463 14487 1497
rect 14521 1463 14561 1497
rect 14595 1463 14635 1497
rect 14669 1463 14709 1497
rect 14743 1463 14783 1497
rect 14817 1463 14931 1497
rect 14965 1463 15005 1497
rect 15039 1463 15079 1497
rect 15113 1463 15153 1497
rect 15187 1463 15227 1497
rect 15261 1463 15301 1497
rect 15335 1463 15375 1497
rect 15409 1463 15449 1497
rect 15483 1463 15597 1497
rect 15631 1463 15671 1497
rect 15705 1463 15745 1497
rect 15779 1463 15819 1497
rect 15853 1463 15893 1497
rect 15927 1463 15967 1497
rect 16001 1463 16041 1497
rect 16075 1463 16115 1497
rect 16149 1463 16263 1497
rect 16297 1463 16337 1497
rect 16371 1463 16411 1497
rect 16445 1463 16485 1497
rect 16519 1463 16559 1497
rect 16593 1463 16633 1497
rect 16667 1463 16707 1497
rect 16741 1463 16781 1497
rect 16815 1463 16929 1497
rect 16963 1463 17003 1497
rect 17037 1463 17077 1497
rect 17111 1463 17151 1497
rect 17185 1463 17225 1497
rect 17259 1463 17299 1497
rect 17333 1463 17373 1497
rect 17407 1463 17447 1497
rect 17481 1463 17595 1497
rect 17629 1463 17669 1497
rect 17703 1463 17743 1497
rect 17777 1463 17817 1497
rect 17851 1463 17891 1497
rect 17925 1463 18016 1497
rect -34 1446 18016 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 201 1366 235 1446
rect 201 1298 235 1332
rect 201 1230 235 1264
rect 201 1162 235 1196
rect 201 1093 235 1128
rect 201 1043 235 1059
rect 289 1366 323 1404
rect 289 1298 323 1332
rect 289 1230 323 1264
rect 289 1162 323 1196
rect 289 1093 323 1128
rect 377 1366 411 1446
rect 377 1298 411 1332
rect 377 1230 411 1264
rect 377 1162 411 1196
rect 377 1111 411 1128
rect 465 1366 499 1404
rect 465 1298 499 1332
rect 465 1230 499 1264
rect 465 1162 499 1196
rect 289 1048 323 1059
rect 465 1093 499 1128
rect 553 1366 587 1446
rect 553 1298 587 1332
rect 553 1230 587 1264
rect 553 1162 587 1196
rect 553 1111 587 1128
rect 641 1366 675 1404
rect 641 1298 675 1332
rect 641 1230 675 1264
rect 641 1162 675 1196
rect 465 1048 499 1059
rect 641 1093 675 1128
rect 729 1366 763 1446
rect 729 1298 763 1332
rect 729 1230 763 1264
rect 729 1162 763 1196
rect 729 1111 763 1128
rect 928 1423 996 1446
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 641 1048 675 1059
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect -34 979 34 1019
rect 289 1014 831 1048
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect 205 831 239 923
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 797
rect 205 383 239 399
rect 427 957 461 973
rect 427 905 461 923
rect 427 433 461 871
rect 427 383 461 399
rect 649 957 683 973
rect 649 683 683 923
rect 649 433 683 649
rect 649 383 683 399
rect 797 757 831 1014
rect 928 1019 945 1053
rect 979 1019 996 1053
rect 1163 1366 1197 1446
rect 1163 1298 1197 1332
rect 1163 1230 1197 1264
rect 1163 1162 1197 1196
rect 1163 1093 1197 1128
rect 1163 1043 1197 1059
rect 1251 1366 1285 1404
rect 1251 1298 1285 1332
rect 1251 1230 1285 1264
rect 1251 1162 1285 1196
rect 1251 1093 1285 1128
rect 1339 1366 1373 1446
rect 1339 1298 1373 1332
rect 1339 1230 1373 1264
rect 1339 1162 1373 1196
rect 1339 1111 1373 1128
rect 1427 1366 1461 1404
rect 1427 1298 1461 1332
rect 1427 1230 1461 1264
rect 1427 1162 1461 1196
rect 1251 1048 1285 1059
rect 1427 1093 1461 1128
rect 1515 1366 1549 1446
rect 1515 1298 1549 1332
rect 1515 1230 1549 1264
rect 1515 1162 1549 1196
rect 1515 1111 1549 1128
rect 1603 1366 1637 1404
rect 1603 1298 1637 1332
rect 1603 1230 1637 1264
rect 1603 1162 1637 1196
rect 1427 1048 1461 1059
rect 1603 1093 1637 1128
rect 1691 1366 1725 1446
rect 1691 1298 1725 1332
rect 1691 1230 1725 1264
rect 1691 1162 1725 1196
rect 1691 1111 1725 1128
rect 1890 1423 1958 1446
rect 1890 1389 1907 1423
rect 1941 1389 1958 1423
rect 1890 1349 1958 1389
rect 1890 1315 1907 1349
rect 1941 1315 1958 1349
rect 1890 1275 1958 1315
rect 1890 1241 1907 1275
rect 1941 1241 1958 1275
rect 1890 1201 1958 1241
rect 1890 1167 1907 1201
rect 1941 1167 1958 1201
rect 1890 1127 1958 1167
rect 1603 1048 1637 1059
rect 1890 1093 1907 1127
rect 1941 1093 1958 1127
rect 1890 1053 1958 1093
rect 928 979 996 1019
rect 1251 1014 1793 1048
rect 928 945 945 979
rect 979 945 996 979
rect 928 905 996 945
rect 928 871 945 905
rect 979 871 996 905
rect 928 822 996 871
rect 1167 957 1201 973
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 101 335 135 351
rect 295 335 329 351
rect 489 335 523 351
rect 135 301 198 335
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 489 335
rect 101 263 135 301
rect 101 195 135 229
rect 295 263 329 301
rect 489 285 523 301
rect 603 335 637 351
rect 797 350 831 723
rect 1167 757 1201 923
rect 603 263 637 301
rect 101 125 135 161
rect 101 75 135 91
rect 198 210 232 226
rect -34 34 34 57
rect 198 34 232 176
rect 295 195 329 229
rect 393 216 427 232
rect 603 216 637 229
rect 427 195 637 216
rect 427 182 603 195
rect 393 166 427 182
rect 295 125 329 161
rect 700 316 831 350
rect 928 461 996 544
rect 928 427 945 461
rect 979 427 996 461
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect 1167 433 1201 723
rect 1167 383 1201 399
rect 1389 957 1423 973
rect 1389 535 1423 923
rect 1389 433 1423 501
rect 1389 383 1423 399
rect 1611 957 1645 973
rect 1611 461 1645 923
rect 1611 383 1645 399
rect 1759 683 1793 1014
rect 1890 1019 1907 1053
rect 1941 1019 1958 1053
rect 2065 1366 2099 1446
rect 2065 1298 2099 1332
rect 2065 1230 2099 1264
rect 2065 1162 2099 1196
rect 2065 1093 2099 1128
rect 2065 1027 2099 1059
rect 2153 1366 2187 1404
rect 2153 1298 2187 1332
rect 2153 1230 2187 1264
rect 2153 1162 2187 1196
rect 2153 1093 2187 1128
rect 2241 1366 2275 1446
rect 2241 1298 2275 1332
rect 2241 1230 2275 1264
rect 2241 1162 2275 1196
rect 2241 1111 2275 1128
rect 2329 1366 2363 1404
rect 2329 1298 2363 1332
rect 2329 1230 2363 1264
rect 2329 1162 2363 1196
rect 2153 1057 2187 1059
rect 2329 1093 2363 1128
rect 2417 1366 2451 1446
rect 2417 1298 2451 1332
rect 2417 1230 2451 1264
rect 2417 1162 2451 1196
rect 2417 1111 2451 1128
rect 2556 1423 2624 1446
rect 2556 1389 2573 1423
rect 2607 1389 2624 1423
rect 2556 1349 2624 1389
rect 2556 1315 2573 1349
rect 2607 1315 2624 1349
rect 2556 1275 2624 1315
rect 2556 1241 2573 1275
rect 2607 1241 2624 1275
rect 2556 1201 2624 1241
rect 2556 1167 2573 1201
rect 2607 1167 2624 1201
rect 2556 1127 2624 1167
rect 2329 1057 2363 1059
rect 2556 1093 2573 1127
rect 2607 1093 2624 1127
rect 2153 1023 2459 1057
rect 1890 979 1958 1019
rect 1890 945 1907 979
rect 1941 945 1958 979
rect 1890 905 1958 945
rect 1890 871 1907 905
rect 1941 871 1958 905
rect 1890 822 1958 871
rect 2129 957 2163 973
rect 2283 957 2317 973
rect 700 219 734 316
rect 928 313 996 353
rect 928 279 945 313
rect 979 279 996 313
rect 700 169 734 185
rect 797 263 831 279
rect 797 195 831 229
rect 489 125 523 141
rect 329 91 392 125
rect 426 91 489 125
rect 295 75 329 91
rect 489 75 523 91
rect 603 125 637 161
rect 797 125 831 161
rect 637 91 700 125
rect 734 91 797 125
rect 603 75 637 91
rect 797 75 831 91
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect 928 57 945 91
rect 979 57 996 91
rect 1063 335 1097 351
rect 1257 335 1291 351
rect 1451 335 1485 351
rect 1097 301 1160 335
rect 1194 301 1257 335
rect 1291 301 1354 335
rect 1388 301 1451 335
rect 1063 263 1097 301
rect 1063 195 1097 229
rect 1257 263 1291 301
rect 1451 285 1485 301
rect 1565 335 1599 351
rect 1759 350 1793 649
rect 2129 683 2163 923
rect 1565 263 1599 301
rect 1063 125 1097 161
rect 1063 75 1097 91
rect 1160 210 1194 226
rect 928 34 996 57
rect 1160 34 1194 176
rect 1257 195 1291 229
rect 1355 216 1389 232
rect 1565 216 1599 229
rect 1389 195 1599 216
rect 1389 182 1565 195
rect 1355 166 1389 182
rect 1257 125 1291 161
rect 1662 316 1793 350
rect 1890 461 1958 544
rect 1890 427 1907 461
rect 1941 427 1958 461
rect 1890 387 1958 427
rect 1890 353 1907 387
rect 1941 353 1958 387
rect 2129 433 2163 649
rect 2129 383 2163 399
rect 2277 923 2283 942
rect 2277 907 2317 923
rect 2277 831 2311 907
rect 2277 433 2311 797
rect 2277 383 2311 399
rect 2425 683 2459 1023
rect 2556 1053 2624 1093
rect 2556 1019 2573 1053
rect 2607 1019 2624 1053
rect 2791 1366 2825 1446
rect 2791 1298 2825 1332
rect 2791 1230 2825 1264
rect 2791 1162 2825 1196
rect 2791 1093 2825 1128
rect 2791 1043 2825 1059
rect 2879 1366 2913 1404
rect 2879 1298 2913 1332
rect 2879 1230 2913 1264
rect 2879 1162 2913 1196
rect 2879 1093 2913 1128
rect 2967 1366 3001 1446
rect 2967 1298 3001 1332
rect 2967 1230 3001 1264
rect 2967 1162 3001 1196
rect 2967 1111 3001 1128
rect 3055 1366 3089 1404
rect 3055 1298 3089 1332
rect 3055 1230 3089 1264
rect 3055 1162 3089 1196
rect 2879 1048 2913 1059
rect 3055 1093 3089 1128
rect 3143 1366 3177 1446
rect 3143 1298 3177 1332
rect 3143 1230 3177 1264
rect 3143 1162 3177 1196
rect 3143 1111 3177 1128
rect 3231 1366 3265 1404
rect 3231 1298 3265 1332
rect 3231 1230 3265 1264
rect 3231 1162 3265 1196
rect 3055 1048 3089 1059
rect 3231 1093 3265 1128
rect 3319 1366 3353 1446
rect 3319 1298 3353 1332
rect 3319 1230 3353 1264
rect 3319 1162 3353 1196
rect 3319 1111 3353 1128
rect 3518 1423 3586 1446
rect 3518 1389 3535 1423
rect 3569 1389 3586 1423
rect 3518 1349 3586 1389
rect 3518 1315 3535 1349
rect 3569 1315 3586 1349
rect 3518 1275 3586 1315
rect 3518 1241 3535 1275
rect 3569 1241 3586 1275
rect 3518 1201 3586 1241
rect 3518 1167 3535 1201
rect 3569 1167 3586 1201
rect 3518 1127 3586 1167
rect 3231 1048 3265 1059
rect 3518 1093 3535 1127
rect 3569 1093 3586 1127
rect 3518 1053 3586 1093
rect 2556 979 2624 1019
rect 2879 1014 3421 1048
rect 2556 945 2573 979
rect 2607 945 2624 979
rect 2556 905 2624 945
rect 2556 871 2573 905
rect 2607 871 2624 905
rect 2556 822 2624 871
rect 2795 957 2829 973
rect 1662 219 1696 316
rect 1890 313 1958 353
rect 1890 279 1907 313
rect 1941 279 1958 313
rect 1662 169 1696 185
rect 1759 263 1793 279
rect 1759 195 1793 229
rect 1451 125 1485 141
rect 1291 91 1354 125
rect 1388 91 1451 125
rect 1257 75 1291 91
rect 1451 75 1485 91
rect 1565 125 1599 161
rect 1759 125 1793 161
rect 1599 91 1662 125
rect 1696 91 1759 125
rect 1565 75 1599 91
rect 1759 75 1793 91
rect 1890 239 1958 279
rect 1890 205 1907 239
rect 1941 205 1958 239
rect 1890 165 1958 205
rect 1890 131 1907 165
rect 1941 131 1958 165
rect 1890 91 1958 131
rect 1890 57 1907 91
rect 1941 57 1958 91
rect 2046 333 2080 349
rect 2240 333 2274 349
rect 2425 348 2459 649
rect 2795 683 2829 923
rect 2080 299 2143 333
rect 2177 299 2240 333
rect 2046 261 2080 299
rect 2046 193 2080 227
rect 2240 261 2274 299
rect 2046 123 2080 159
rect 2046 73 2080 89
rect 2143 208 2177 224
rect 1890 34 1958 57
rect 2143 34 2177 174
rect 2240 193 2274 227
rect 2337 314 2459 348
rect 2556 461 2624 544
rect 2556 427 2573 461
rect 2607 427 2624 461
rect 2556 387 2624 427
rect 2556 353 2573 387
rect 2607 353 2624 387
rect 2795 433 2829 649
rect 2795 383 2829 399
rect 3017 957 3051 973
rect 3017 905 3051 923
rect 3017 433 3051 871
rect 3017 383 3051 399
rect 3239 957 3273 973
rect 3239 461 3273 923
rect 3239 383 3273 399
rect 3387 831 3421 1014
rect 3518 1019 3535 1053
rect 3569 1019 3586 1053
rect 3753 1366 3787 1446
rect 3753 1298 3787 1332
rect 3753 1230 3787 1264
rect 3753 1162 3787 1196
rect 3753 1093 3787 1128
rect 3753 1043 3787 1059
rect 3841 1366 3875 1404
rect 3841 1298 3875 1332
rect 3841 1230 3875 1264
rect 3841 1162 3875 1196
rect 3841 1093 3875 1128
rect 3929 1366 3963 1446
rect 3929 1298 3963 1332
rect 3929 1230 3963 1264
rect 3929 1162 3963 1196
rect 3929 1111 3963 1128
rect 4017 1366 4051 1404
rect 4017 1298 4051 1332
rect 4017 1230 4051 1264
rect 4017 1162 4051 1196
rect 3841 1048 3875 1059
rect 4017 1093 4051 1128
rect 4105 1366 4139 1446
rect 4105 1298 4139 1332
rect 4105 1230 4139 1264
rect 4105 1162 4139 1196
rect 4105 1111 4139 1128
rect 4193 1366 4227 1404
rect 4193 1298 4227 1332
rect 4193 1230 4227 1264
rect 4193 1162 4227 1196
rect 4017 1048 4051 1059
rect 4193 1093 4227 1128
rect 4281 1366 4315 1446
rect 4281 1298 4315 1332
rect 4281 1230 4315 1264
rect 4281 1162 4315 1196
rect 4281 1111 4315 1128
rect 4480 1423 4548 1446
rect 4480 1389 4497 1423
rect 4531 1389 4548 1423
rect 4480 1349 4548 1389
rect 4480 1315 4497 1349
rect 4531 1315 4548 1349
rect 4480 1275 4548 1315
rect 4480 1241 4497 1275
rect 4531 1241 4548 1275
rect 4480 1201 4548 1241
rect 4480 1167 4497 1201
rect 4531 1167 4548 1201
rect 4480 1127 4548 1167
rect 4193 1048 4227 1059
rect 4480 1093 4497 1127
rect 4531 1093 4548 1127
rect 4480 1053 4548 1093
rect 3518 979 3586 1019
rect 3841 1014 4383 1048
rect 3518 945 3535 979
rect 3569 945 3586 979
rect 3518 905 3586 945
rect 3518 871 3535 905
rect 3569 871 3586 905
rect 3518 822 3586 871
rect 3757 957 3791 973
rect 2337 217 2371 314
rect 2556 313 2624 353
rect 2556 279 2573 313
rect 2607 279 2624 313
rect 2337 167 2371 183
rect 2434 261 2468 277
rect 2434 193 2468 227
rect 2240 123 2274 159
rect 2434 123 2468 159
rect 2274 89 2337 123
rect 2371 89 2434 123
rect 2240 73 2274 89
rect 2434 73 2468 89
rect 2556 239 2624 279
rect 2556 205 2573 239
rect 2607 205 2624 239
rect 2556 165 2624 205
rect 2556 131 2573 165
rect 2607 131 2624 165
rect 2556 91 2624 131
rect 2556 57 2573 91
rect 2607 57 2624 91
rect 2691 335 2725 351
rect 2885 335 2919 351
rect 3079 335 3113 351
rect 2725 301 2788 335
rect 2822 301 2885 335
rect 2919 301 2982 335
rect 3016 301 3079 335
rect 2691 263 2725 301
rect 2691 195 2725 229
rect 2885 263 2919 301
rect 3079 285 3113 301
rect 3193 335 3227 351
rect 3387 350 3421 797
rect 3757 757 3791 923
rect 3193 263 3227 301
rect 2691 125 2725 161
rect 2691 75 2725 91
rect 2788 210 2822 226
rect 2556 34 2624 57
rect 2788 34 2822 176
rect 2885 195 2919 229
rect 2983 216 3017 232
rect 3193 216 3227 229
rect 3017 195 3227 216
rect 3017 182 3193 195
rect 2983 166 3017 182
rect 2885 125 2919 161
rect 3290 316 3421 350
rect 3518 461 3586 544
rect 3518 427 3535 461
rect 3569 427 3586 461
rect 3518 387 3586 427
rect 3518 353 3535 387
rect 3569 353 3586 387
rect 3757 433 3791 723
rect 3757 383 3791 399
rect 3979 957 4013 973
rect 3979 461 4013 923
rect 3979 383 4013 399
rect 4201 957 4235 973
rect 4201 609 4235 923
rect 4201 433 4235 575
rect 4201 383 4235 399
rect 4349 831 4383 1014
rect 4480 1019 4497 1053
rect 4531 1019 4548 1053
rect 4655 1366 4689 1446
rect 4655 1298 4689 1332
rect 4655 1230 4689 1264
rect 4655 1162 4689 1196
rect 4655 1093 4689 1128
rect 4655 1027 4689 1059
rect 4743 1366 4777 1404
rect 4743 1298 4777 1332
rect 4743 1230 4777 1264
rect 4743 1162 4777 1196
rect 4743 1093 4777 1128
rect 4831 1366 4865 1446
rect 4831 1298 4865 1332
rect 4831 1230 4865 1264
rect 4831 1162 4865 1196
rect 4831 1111 4865 1128
rect 4919 1366 4953 1404
rect 4919 1298 4953 1332
rect 4919 1230 4953 1264
rect 4919 1162 4953 1196
rect 4743 1057 4777 1059
rect 4919 1093 4953 1128
rect 5007 1366 5041 1446
rect 5007 1298 5041 1332
rect 5007 1230 5041 1264
rect 5007 1162 5041 1196
rect 5007 1111 5041 1128
rect 5146 1423 5214 1446
rect 5146 1389 5163 1423
rect 5197 1389 5214 1423
rect 5146 1349 5214 1389
rect 5146 1315 5163 1349
rect 5197 1315 5214 1349
rect 5146 1275 5214 1315
rect 5146 1241 5163 1275
rect 5197 1241 5214 1275
rect 5146 1201 5214 1241
rect 5146 1167 5163 1201
rect 5197 1167 5214 1201
rect 5146 1127 5214 1167
rect 4919 1057 4953 1059
rect 5146 1093 5163 1127
rect 5197 1093 5214 1127
rect 4743 1023 5049 1057
rect 4480 979 4548 1019
rect 4480 945 4497 979
rect 4531 945 4548 979
rect 4480 905 4548 945
rect 4480 871 4497 905
rect 4531 871 4548 905
rect 4480 822 4548 871
rect 4719 957 4753 973
rect 4873 957 4907 973
rect 4719 831 4753 923
rect 3290 219 3324 316
rect 3518 313 3586 353
rect 3518 279 3535 313
rect 3569 279 3586 313
rect 3290 169 3324 185
rect 3387 263 3421 279
rect 3387 195 3421 229
rect 3079 125 3113 141
rect 2919 91 2982 125
rect 3016 91 3079 125
rect 2885 75 2919 91
rect 3079 75 3113 91
rect 3193 125 3227 161
rect 3387 125 3421 161
rect 3227 91 3290 125
rect 3324 91 3387 125
rect 3193 75 3227 91
rect 3387 75 3421 91
rect 3518 239 3586 279
rect 3518 205 3535 239
rect 3569 205 3586 239
rect 3518 165 3586 205
rect 3518 131 3535 165
rect 3569 131 3586 165
rect 3518 91 3586 131
rect 3518 57 3535 91
rect 3569 57 3586 91
rect 3653 335 3687 351
rect 3847 335 3881 351
rect 4041 335 4075 351
rect 3687 301 3750 335
rect 3784 301 3847 335
rect 3881 301 3944 335
rect 3978 301 4041 335
rect 3653 263 3687 301
rect 3653 195 3687 229
rect 3847 263 3881 301
rect 4041 285 4075 301
rect 4155 335 4189 351
rect 4349 350 4383 797
rect 4155 263 4189 301
rect 3653 125 3687 161
rect 3653 75 3687 91
rect 3750 210 3784 226
rect 3518 34 3586 57
rect 3750 34 3784 176
rect 3847 195 3881 229
rect 3945 216 3979 232
rect 4155 216 4189 229
rect 3979 195 4189 216
rect 3979 182 4155 195
rect 3945 166 3979 182
rect 3847 125 3881 161
rect 4252 316 4383 350
rect 4480 461 4548 544
rect 4480 427 4497 461
rect 4531 427 4548 461
rect 4480 387 4548 427
rect 4480 353 4497 387
rect 4531 353 4548 387
rect 4719 433 4753 797
rect 4719 383 4753 399
rect 4867 923 4873 942
rect 4867 907 4907 923
rect 4867 831 4901 907
rect 4867 433 4901 797
rect 4867 383 4901 399
rect 5015 609 5049 1023
rect 5146 1053 5214 1093
rect 5146 1019 5163 1053
rect 5197 1019 5214 1053
rect 5381 1366 5415 1446
rect 5381 1298 5415 1332
rect 5381 1230 5415 1264
rect 5381 1162 5415 1196
rect 5381 1093 5415 1128
rect 5381 1043 5415 1059
rect 5469 1366 5503 1404
rect 5469 1298 5503 1332
rect 5469 1230 5503 1264
rect 5469 1162 5503 1196
rect 5469 1093 5503 1128
rect 5557 1366 5591 1446
rect 5557 1298 5591 1332
rect 5557 1230 5591 1264
rect 5557 1162 5591 1196
rect 5557 1111 5591 1128
rect 5645 1366 5679 1404
rect 5645 1298 5679 1332
rect 5645 1230 5679 1264
rect 5645 1162 5679 1196
rect 5469 1048 5503 1059
rect 5645 1093 5679 1128
rect 5733 1366 5767 1446
rect 5733 1298 5767 1332
rect 5733 1230 5767 1264
rect 5733 1162 5767 1196
rect 5733 1111 5767 1128
rect 5821 1366 5855 1404
rect 5821 1298 5855 1332
rect 5821 1230 5855 1264
rect 5821 1162 5855 1196
rect 5645 1048 5679 1059
rect 5821 1093 5855 1128
rect 5909 1366 5943 1446
rect 5909 1298 5943 1332
rect 5909 1230 5943 1264
rect 5909 1162 5943 1196
rect 5909 1111 5943 1128
rect 6108 1423 6176 1446
rect 6108 1389 6125 1423
rect 6159 1389 6176 1423
rect 6108 1349 6176 1389
rect 6108 1315 6125 1349
rect 6159 1315 6176 1349
rect 6108 1275 6176 1315
rect 6108 1241 6125 1275
rect 6159 1241 6176 1275
rect 6108 1201 6176 1241
rect 6108 1167 6125 1201
rect 6159 1167 6176 1201
rect 6108 1127 6176 1167
rect 5821 1048 5855 1059
rect 6108 1093 6125 1127
rect 6159 1093 6176 1127
rect 6108 1053 6176 1093
rect 5146 979 5214 1019
rect 5469 1014 6011 1048
rect 5146 945 5163 979
rect 5197 945 5214 979
rect 5146 905 5214 945
rect 5146 871 5163 905
rect 5197 871 5214 905
rect 5146 822 5214 871
rect 5385 957 5419 973
rect 5385 831 5419 923
rect 4252 219 4286 316
rect 4480 313 4548 353
rect 4480 279 4497 313
rect 4531 279 4548 313
rect 4252 169 4286 185
rect 4349 263 4383 279
rect 4349 195 4383 229
rect 4041 125 4075 141
rect 3881 91 3944 125
rect 3978 91 4041 125
rect 3847 75 3881 91
rect 4041 75 4075 91
rect 4155 125 4189 161
rect 4349 125 4383 161
rect 4189 91 4252 125
rect 4286 91 4349 125
rect 4155 75 4189 91
rect 4349 75 4383 91
rect 4480 239 4548 279
rect 4480 205 4497 239
rect 4531 205 4548 239
rect 4480 165 4548 205
rect 4480 131 4497 165
rect 4531 131 4548 165
rect 4480 91 4548 131
rect 4480 57 4497 91
rect 4531 57 4548 91
rect 4636 333 4670 349
rect 4830 333 4864 349
rect 5015 348 5049 575
rect 4670 299 4733 333
rect 4767 299 4830 333
rect 4636 261 4670 299
rect 4636 193 4670 227
rect 4830 261 4864 299
rect 4636 123 4670 159
rect 4636 73 4670 89
rect 4733 208 4767 224
rect 4480 34 4548 57
rect 4733 34 4767 174
rect 4830 193 4864 227
rect 4927 314 5049 348
rect 5146 461 5214 544
rect 5146 427 5163 461
rect 5197 427 5214 461
rect 5146 387 5214 427
rect 5146 353 5163 387
rect 5197 353 5214 387
rect 5385 433 5419 797
rect 5385 383 5419 399
rect 5607 957 5641 973
rect 5607 905 5641 923
rect 5607 433 5641 871
rect 5607 383 5641 399
rect 5829 957 5863 973
rect 5829 683 5863 923
rect 5829 433 5863 649
rect 5829 383 5863 399
rect 5977 757 6011 1014
rect 6108 1019 6125 1053
rect 6159 1019 6176 1053
rect 6343 1366 6377 1446
rect 6343 1298 6377 1332
rect 6343 1230 6377 1264
rect 6343 1162 6377 1196
rect 6343 1093 6377 1128
rect 6343 1043 6377 1059
rect 6431 1366 6465 1404
rect 6431 1298 6465 1332
rect 6431 1230 6465 1264
rect 6431 1162 6465 1196
rect 6431 1093 6465 1128
rect 6519 1366 6553 1446
rect 6519 1298 6553 1332
rect 6519 1230 6553 1264
rect 6519 1162 6553 1196
rect 6519 1111 6553 1128
rect 6607 1366 6641 1404
rect 6607 1298 6641 1332
rect 6607 1230 6641 1264
rect 6607 1162 6641 1196
rect 6431 1048 6465 1059
rect 6607 1093 6641 1128
rect 6695 1366 6729 1446
rect 6695 1298 6729 1332
rect 6695 1230 6729 1264
rect 6695 1162 6729 1196
rect 6695 1111 6729 1128
rect 6783 1366 6817 1404
rect 6783 1298 6817 1332
rect 6783 1230 6817 1264
rect 6783 1162 6817 1196
rect 6607 1048 6641 1059
rect 6783 1093 6817 1128
rect 6871 1366 6905 1446
rect 6871 1298 6905 1332
rect 6871 1230 6905 1264
rect 6871 1162 6905 1196
rect 6871 1111 6905 1128
rect 7070 1423 7138 1446
rect 7070 1389 7087 1423
rect 7121 1389 7138 1423
rect 7070 1349 7138 1389
rect 7070 1315 7087 1349
rect 7121 1315 7138 1349
rect 7070 1275 7138 1315
rect 7070 1241 7087 1275
rect 7121 1241 7138 1275
rect 7070 1201 7138 1241
rect 7070 1167 7087 1201
rect 7121 1167 7138 1201
rect 7070 1127 7138 1167
rect 6783 1048 6817 1059
rect 7070 1093 7087 1127
rect 7121 1093 7138 1127
rect 7070 1053 7138 1093
rect 6108 979 6176 1019
rect 6431 1014 6973 1048
rect 6108 945 6125 979
rect 6159 945 6176 979
rect 6108 905 6176 945
rect 6108 871 6125 905
rect 6159 871 6176 905
rect 6108 822 6176 871
rect 6347 957 6381 973
rect 4927 217 4961 314
rect 5146 313 5214 353
rect 5146 279 5163 313
rect 5197 279 5214 313
rect 4927 167 4961 183
rect 5024 261 5058 277
rect 5024 193 5058 227
rect 4830 123 4864 159
rect 5024 123 5058 159
rect 4864 89 4927 123
rect 4961 89 5024 123
rect 4830 73 4864 89
rect 5024 73 5058 89
rect 5146 239 5214 279
rect 5146 205 5163 239
rect 5197 205 5214 239
rect 5146 165 5214 205
rect 5146 131 5163 165
rect 5197 131 5214 165
rect 5146 91 5214 131
rect 5146 57 5163 91
rect 5197 57 5214 91
rect 5281 335 5315 351
rect 5475 335 5509 351
rect 5669 335 5703 351
rect 5315 301 5378 335
rect 5412 301 5475 335
rect 5509 301 5572 335
rect 5606 301 5669 335
rect 5281 263 5315 301
rect 5281 195 5315 229
rect 5475 263 5509 301
rect 5669 285 5703 301
rect 5783 335 5817 351
rect 5977 350 6011 723
rect 6347 757 6381 923
rect 5783 263 5817 301
rect 5281 125 5315 161
rect 5281 75 5315 91
rect 5378 210 5412 226
rect 5146 34 5214 57
rect 5378 34 5412 176
rect 5475 195 5509 229
rect 5573 216 5607 232
rect 5783 216 5817 229
rect 5607 195 5817 216
rect 5607 182 5783 195
rect 5573 166 5607 182
rect 5475 125 5509 161
rect 5880 316 6011 350
rect 6108 461 6176 544
rect 6108 427 6125 461
rect 6159 427 6176 461
rect 6108 387 6176 427
rect 6108 353 6125 387
rect 6159 353 6176 387
rect 6347 433 6381 723
rect 6347 383 6381 399
rect 6569 957 6603 973
rect 6569 535 6603 923
rect 6569 433 6603 501
rect 6569 383 6603 399
rect 6791 957 6825 973
rect 6791 461 6825 923
rect 6791 383 6825 399
rect 6939 683 6973 1014
rect 7070 1019 7087 1053
rect 7121 1019 7138 1053
rect 7245 1366 7279 1446
rect 7245 1298 7279 1332
rect 7245 1230 7279 1264
rect 7245 1162 7279 1196
rect 7245 1093 7279 1128
rect 7245 1027 7279 1059
rect 7333 1366 7367 1404
rect 7333 1298 7367 1332
rect 7333 1230 7367 1264
rect 7333 1162 7367 1196
rect 7333 1093 7367 1128
rect 7421 1366 7455 1446
rect 7421 1298 7455 1332
rect 7421 1230 7455 1264
rect 7421 1162 7455 1196
rect 7421 1111 7455 1128
rect 7509 1366 7543 1404
rect 7509 1298 7543 1332
rect 7509 1230 7543 1264
rect 7509 1162 7543 1196
rect 7333 1057 7367 1059
rect 7509 1093 7543 1128
rect 7597 1366 7631 1446
rect 7597 1298 7631 1332
rect 7597 1230 7631 1264
rect 7597 1162 7631 1196
rect 7597 1111 7631 1128
rect 7736 1423 7804 1446
rect 7736 1389 7753 1423
rect 7787 1389 7804 1423
rect 7736 1349 7804 1389
rect 7736 1315 7753 1349
rect 7787 1315 7804 1349
rect 7736 1275 7804 1315
rect 7736 1241 7753 1275
rect 7787 1241 7804 1275
rect 7736 1201 7804 1241
rect 7736 1167 7753 1201
rect 7787 1167 7804 1201
rect 7736 1127 7804 1167
rect 7509 1057 7543 1059
rect 7736 1093 7753 1127
rect 7787 1093 7804 1127
rect 7333 1023 7639 1057
rect 7070 979 7138 1019
rect 7070 945 7087 979
rect 7121 945 7138 979
rect 7070 905 7138 945
rect 7070 871 7087 905
rect 7121 871 7138 905
rect 7070 822 7138 871
rect 7309 957 7343 973
rect 7463 957 7497 973
rect 5880 219 5914 316
rect 6108 313 6176 353
rect 6108 279 6125 313
rect 6159 279 6176 313
rect 5880 169 5914 185
rect 5977 263 6011 279
rect 5977 195 6011 229
rect 5669 125 5703 141
rect 5509 91 5572 125
rect 5606 91 5669 125
rect 5475 75 5509 91
rect 5669 75 5703 91
rect 5783 125 5817 161
rect 5977 125 6011 161
rect 5817 91 5880 125
rect 5914 91 5977 125
rect 5783 75 5817 91
rect 5977 75 6011 91
rect 6108 239 6176 279
rect 6108 205 6125 239
rect 6159 205 6176 239
rect 6108 165 6176 205
rect 6108 131 6125 165
rect 6159 131 6176 165
rect 6108 91 6176 131
rect 6108 57 6125 91
rect 6159 57 6176 91
rect 6243 335 6277 351
rect 6437 335 6471 351
rect 6631 335 6665 351
rect 6277 301 6340 335
rect 6374 301 6437 335
rect 6471 301 6534 335
rect 6568 301 6631 335
rect 6243 263 6277 301
rect 6243 195 6277 229
rect 6437 263 6471 301
rect 6631 285 6665 301
rect 6745 335 6779 351
rect 6939 350 6973 649
rect 7309 683 7343 923
rect 6745 263 6779 301
rect 6243 125 6277 161
rect 6243 75 6277 91
rect 6340 210 6374 226
rect 6108 34 6176 57
rect 6340 34 6374 176
rect 6437 195 6471 229
rect 6535 216 6569 232
rect 6745 216 6779 229
rect 6569 195 6779 216
rect 6569 182 6745 195
rect 6535 166 6569 182
rect 6437 125 6471 161
rect 6842 316 6973 350
rect 7070 461 7138 544
rect 7070 427 7087 461
rect 7121 427 7138 461
rect 7070 387 7138 427
rect 7070 353 7087 387
rect 7121 353 7138 387
rect 7309 433 7343 649
rect 7309 383 7343 399
rect 7457 923 7463 942
rect 7457 907 7497 923
rect 7457 831 7491 907
rect 7457 433 7491 797
rect 7457 383 7491 399
rect 7605 683 7639 1023
rect 7736 1053 7804 1093
rect 7736 1019 7753 1053
rect 7787 1019 7804 1053
rect 7971 1366 8005 1446
rect 7971 1298 8005 1332
rect 7971 1230 8005 1264
rect 7971 1162 8005 1196
rect 7971 1093 8005 1128
rect 7971 1043 8005 1059
rect 8059 1366 8093 1404
rect 8059 1298 8093 1332
rect 8059 1230 8093 1264
rect 8059 1162 8093 1196
rect 8059 1093 8093 1128
rect 8147 1366 8181 1446
rect 8147 1298 8181 1332
rect 8147 1230 8181 1264
rect 8147 1162 8181 1196
rect 8147 1111 8181 1128
rect 8235 1366 8269 1404
rect 8235 1298 8269 1332
rect 8235 1230 8269 1264
rect 8235 1162 8269 1196
rect 8059 1048 8093 1059
rect 8235 1093 8269 1128
rect 8323 1366 8357 1446
rect 8323 1298 8357 1332
rect 8323 1230 8357 1264
rect 8323 1162 8357 1196
rect 8323 1111 8357 1128
rect 8411 1366 8445 1404
rect 8411 1298 8445 1332
rect 8411 1230 8445 1264
rect 8411 1162 8445 1196
rect 8235 1048 8269 1059
rect 8411 1093 8445 1128
rect 8499 1366 8533 1446
rect 8499 1298 8533 1332
rect 8499 1230 8533 1264
rect 8499 1162 8533 1196
rect 8499 1111 8533 1128
rect 8698 1423 8766 1446
rect 8698 1389 8715 1423
rect 8749 1389 8766 1423
rect 8698 1349 8766 1389
rect 8698 1315 8715 1349
rect 8749 1315 8766 1349
rect 8698 1275 8766 1315
rect 8698 1241 8715 1275
rect 8749 1241 8766 1275
rect 8698 1201 8766 1241
rect 8698 1167 8715 1201
rect 8749 1167 8766 1201
rect 8698 1127 8766 1167
rect 8411 1048 8445 1059
rect 8698 1093 8715 1127
rect 8749 1093 8766 1127
rect 8698 1053 8766 1093
rect 7736 979 7804 1019
rect 8059 1014 8601 1048
rect 7736 945 7753 979
rect 7787 945 7804 979
rect 7736 905 7804 945
rect 7736 871 7753 905
rect 7787 871 7804 905
rect 7736 822 7804 871
rect 7975 957 8009 973
rect 6842 219 6876 316
rect 7070 313 7138 353
rect 7070 279 7087 313
rect 7121 279 7138 313
rect 6842 169 6876 185
rect 6939 263 6973 279
rect 6939 195 6973 229
rect 6631 125 6665 141
rect 6471 91 6534 125
rect 6568 91 6631 125
rect 6437 75 6471 91
rect 6631 75 6665 91
rect 6745 125 6779 161
rect 6939 125 6973 161
rect 6779 91 6842 125
rect 6876 91 6939 125
rect 6745 75 6779 91
rect 6939 75 6973 91
rect 7070 239 7138 279
rect 7070 205 7087 239
rect 7121 205 7138 239
rect 7070 165 7138 205
rect 7070 131 7087 165
rect 7121 131 7138 165
rect 7070 91 7138 131
rect 7070 57 7087 91
rect 7121 57 7138 91
rect 7226 333 7260 349
rect 7420 333 7454 349
rect 7605 348 7639 649
rect 7975 683 8009 923
rect 7260 299 7323 333
rect 7357 299 7420 333
rect 7226 261 7260 299
rect 7226 193 7260 227
rect 7420 261 7454 299
rect 7226 123 7260 159
rect 7226 73 7260 89
rect 7323 208 7357 224
rect 7070 34 7138 57
rect 7323 34 7357 174
rect 7420 193 7454 227
rect 7517 314 7639 348
rect 7736 461 7804 544
rect 7736 427 7753 461
rect 7787 427 7804 461
rect 7736 387 7804 427
rect 7736 353 7753 387
rect 7787 353 7804 387
rect 7975 433 8009 649
rect 7975 383 8009 399
rect 8197 957 8231 973
rect 8197 905 8231 923
rect 8197 433 8231 871
rect 8197 383 8231 399
rect 8419 957 8453 973
rect 8419 461 8453 923
rect 8419 383 8453 399
rect 8567 831 8601 1014
rect 8698 1019 8715 1053
rect 8749 1019 8766 1053
rect 8933 1366 8967 1446
rect 8933 1298 8967 1332
rect 8933 1230 8967 1264
rect 8933 1162 8967 1196
rect 8933 1093 8967 1128
rect 8933 1043 8967 1059
rect 9021 1366 9055 1404
rect 9021 1298 9055 1332
rect 9021 1230 9055 1264
rect 9021 1162 9055 1196
rect 9021 1093 9055 1128
rect 9109 1366 9143 1446
rect 9109 1298 9143 1332
rect 9109 1230 9143 1264
rect 9109 1162 9143 1196
rect 9109 1111 9143 1128
rect 9197 1366 9231 1404
rect 9197 1298 9231 1332
rect 9197 1230 9231 1264
rect 9197 1162 9231 1196
rect 9021 1048 9055 1059
rect 9197 1093 9231 1128
rect 9285 1366 9319 1446
rect 9285 1298 9319 1332
rect 9285 1230 9319 1264
rect 9285 1162 9319 1196
rect 9285 1111 9319 1128
rect 9373 1366 9407 1404
rect 9373 1298 9407 1332
rect 9373 1230 9407 1264
rect 9373 1162 9407 1196
rect 9197 1048 9231 1059
rect 9373 1093 9407 1128
rect 9461 1366 9495 1446
rect 9461 1298 9495 1332
rect 9461 1230 9495 1264
rect 9461 1162 9495 1196
rect 9461 1111 9495 1128
rect 9660 1423 9728 1446
rect 9660 1389 9677 1423
rect 9711 1389 9728 1423
rect 9660 1349 9728 1389
rect 9660 1315 9677 1349
rect 9711 1315 9728 1349
rect 9660 1275 9728 1315
rect 9660 1241 9677 1275
rect 9711 1241 9728 1275
rect 9660 1201 9728 1241
rect 9660 1167 9677 1201
rect 9711 1167 9728 1201
rect 9660 1127 9728 1167
rect 9373 1048 9407 1059
rect 9660 1093 9677 1127
rect 9711 1093 9728 1127
rect 9660 1053 9728 1093
rect 8698 979 8766 1019
rect 9021 1014 9563 1048
rect 8698 945 8715 979
rect 8749 945 8766 979
rect 8698 905 8766 945
rect 8698 871 8715 905
rect 8749 871 8766 905
rect 8698 822 8766 871
rect 8937 957 8971 973
rect 7517 217 7551 314
rect 7736 313 7804 353
rect 7736 279 7753 313
rect 7787 279 7804 313
rect 7517 167 7551 183
rect 7614 261 7648 277
rect 7614 193 7648 227
rect 7420 123 7454 159
rect 7614 123 7648 159
rect 7454 89 7517 123
rect 7551 89 7614 123
rect 7420 73 7454 89
rect 7614 73 7648 89
rect 7736 239 7804 279
rect 7736 205 7753 239
rect 7787 205 7804 239
rect 7736 165 7804 205
rect 7736 131 7753 165
rect 7787 131 7804 165
rect 7736 91 7804 131
rect 7736 57 7753 91
rect 7787 57 7804 91
rect 7871 335 7905 351
rect 8065 335 8099 351
rect 8259 335 8293 351
rect 7905 301 7968 335
rect 8002 301 8065 335
rect 8099 301 8162 335
rect 8196 301 8259 335
rect 7871 263 7905 301
rect 7871 195 7905 229
rect 8065 263 8099 301
rect 8259 285 8293 301
rect 8373 335 8407 351
rect 8567 350 8601 797
rect 8937 757 8971 923
rect 8373 263 8407 301
rect 7871 125 7905 161
rect 7871 75 7905 91
rect 7968 210 8002 226
rect 7736 34 7804 57
rect 7968 34 8002 176
rect 8065 195 8099 229
rect 8163 216 8197 232
rect 8373 216 8407 229
rect 8197 195 8407 216
rect 8197 182 8373 195
rect 8163 166 8197 182
rect 8065 125 8099 161
rect 8470 316 8601 350
rect 8698 461 8766 544
rect 8698 427 8715 461
rect 8749 427 8766 461
rect 8698 387 8766 427
rect 8698 353 8715 387
rect 8749 353 8766 387
rect 8937 433 8971 723
rect 8937 383 8971 399
rect 9159 957 9193 973
rect 9159 461 9193 923
rect 9159 383 9193 399
rect 9381 957 9415 973
rect 9381 683 9415 923
rect 9381 433 9415 649
rect 9381 383 9415 399
rect 9529 757 9563 1014
rect 9660 1019 9677 1053
rect 9711 1019 9728 1053
rect 9835 1366 9869 1446
rect 9835 1298 9869 1332
rect 9835 1230 9869 1264
rect 9835 1162 9869 1196
rect 9835 1093 9869 1128
rect 9835 1027 9869 1059
rect 9923 1366 9957 1404
rect 9923 1298 9957 1332
rect 9923 1230 9957 1264
rect 9923 1162 9957 1196
rect 9923 1093 9957 1128
rect 10011 1366 10045 1446
rect 10011 1298 10045 1332
rect 10011 1230 10045 1264
rect 10011 1162 10045 1196
rect 10011 1111 10045 1128
rect 10099 1366 10133 1404
rect 10099 1298 10133 1332
rect 10099 1230 10133 1264
rect 10099 1162 10133 1196
rect 9923 1057 9957 1059
rect 10099 1093 10133 1128
rect 10187 1366 10221 1446
rect 10187 1298 10221 1332
rect 10187 1230 10221 1264
rect 10187 1162 10221 1196
rect 10187 1111 10221 1128
rect 10326 1423 10394 1446
rect 10326 1389 10343 1423
rect 10377 1389 10394 1423
rect 10326 1349 10394 1389
rect 10326 1315 10343 1349
rect 10377 1315 10394 1349
rect 10326 1275 10394 1315
rect 10326 1241 10343 1275
rect 10377 1241 10394 1275
rect 10326 1201 10394 1241
rect 10326 1167 10343 1201
rect 10377 1167 10394 1201
rect 10326 1127 10394 1167
rect 10099 1057 10133 1059
rect 10326 1093 10343 1127
rect 10377 1093 10394 1127
rect 9923 1023 10229 1057
rect 9660 979 9728 1019
rect 9660 945 9677 979
rect 9711 945 9728 979
rect 9660 905 9728 945
rect 9660 871 9677 905
rect 9711 871 9728 905
rect 9660 822 9728 871
rect 9899 957 9933 973
rect 10053 957 10087 973
rect 8470 219 8504 316
rect 8698 313 8766 353
rect 8698 279 8715 313
rect 8749 279 8766 313
rect 8470 169 8504 185
rect 8567 263 8601 279
rect 8567 195 8601 229
rect 8259 125 8293 141
rect 8099 91 8162 125
rect 8196 91 8259 125
rect 8065 75 8099 91
rect 8259 75 8293 91
rect 8373 125 8407 161
rect 8567 125 8601 161
rect 8407 91 8470 125
rect 8504 91 8567 125
rect 8373 75 8407 91
rect 8567 75 8601 91
rect 8698 239 8766 279
rect 8698 205 8715 239
rect 8749 205 8766 239
rect 8698 165 8766 205
rect 8698 131 8715 165
rect 8749 131 8766 165
rect 8698 91 8766 131
rect 8698 57 8715 91
rect 8749 57 8766 91
rect 8833 335 8867 351
rect 9027 335 9061 351
rect 9221 335 9255 351
rect 8867 301 8930 335
rect 8964 301 9027 335
rect 9061 301 9124 335
rect 9158 301 9221 335
rect 8833 263 8867 301
rect 8833 195 8867 229
rect 9027 263 9061 301
rect 9221 285 9255 301
rect 9335 335 9369 351
rect 9529 350 9563 723
rect 9899 757 9933 923
rect 9335 263 9369 301
rect 8833 125 8867 161
rect 8833 75 8867 91
rect 8930 210 8964 226
rect 8698 34 8766 57
rect 8930 34 8964 176
rect 9027 195 9061 229
rect 9125 216 9159 232
rect 9335 216 9369 229
rect 9159 195 9369 216
rect 9159 182 9335 195
rect 9125 166 9159 182
rect 9027 125 9061 161
rect 9432 316 9563 350
rect 9660 461 9728 544
rect 9660 427 9677 461
rect 9711 427 9728 461
rect 9660 387 9728 427
rect 9660 353 9677 387
rect 9711 353 9728 387
rect 9899 433 9933 723
rect 9899 383 9933 399
rect 10047 923 10053 942
rect 10047 907 10087 923
rect 10047 831 10081 907
rect 10047 433 10081 797
rect 10047 383 10081 399
rect 10195 683 10229 1023
rect 10326 1053 10394 1093
rect 10326 1019 10343 1053
rect 10377 1019 10394 1053
rect 10561 1366 10595 1446
rect 10561 1298 10595 1332
rect 10561 1230 10595 1264
rect 10561 1162 10595 1196
rect 10561 1093 10595 1128
rect 10561 1043 10595 1059
rect 10649 1366 10683 1404
rect 10649 1298 10683 1332
rect 10649 1230 10683 1264
rect 10649 1162 10683 1196
rect 10649 1093 10683 1128
rect 10737 1366 10771 1446
rect 10737 1298 10771 1332
rect 10737 1230 10771 1264
rect 10737 1162 10771 1196
rect 10737 1111 10771 1128
rect 10825 1366 10859 1404
rect 10825 1298 10859 1332
rect 10825 1230 10859 1264
rect 10825 1162 10859 1196
rect 10649 1048 10683 1059
rect 10825 1093 10859 1128
rect 10913 1366 10947 1446
rect 10913 1298 10947 1332
rect 10913 1230 10947 1264
rect 10913 1162 10947 1196
rect 10913 1111 10947 1128
rect 11001 1366 11035 1404
rect 11001 1298 11035 1332
rect 11001 1230 11035 1264
rect 11001 1162 11035 1196
rect 10825 1048 10859 1059
rect 11001 1093 11035 1128
rect 11089 1366 11123 1446
rect 11089 1298 11123 1332
rect 11089 1230 11123 1264
rect 11089 1162 11123 1196
rect 11089 1111 11123 1128
rect 11288 1423 11356 1446
rect 11288 1389 11305 1423
rect 11339 1389 11356 1423
rect 11288 1349 11356 1389
rect 11288 1315 11305 1349
rect 11339 1315 11356 1349
rect 11288 1275 11356 1315
rect 11288 1241 11305 1275
rect 11339 1241 11356 1275
rect 11288 1201 11356 1241
rect 11288 1167 11305 1201
rect 11339 1167 11356 1201
rect 11288 1127 11356 1167
rect 11001 1048 11035 1059
rect 11288 1093 11305 1127
rect 11339 1093 11356 1127
rect 11288 1053 11356 1093
rect 10326 979 10394 1019
rect 10649 1014 11191 1048
rect 10326 945 10343 979
rect 10377 945 10394 979
rect 10326 905 10394 945
rect 10326 871 10343 905
rect 10377 871 10394 905
rect 10326 822 10394 871
rect 10565 957 10599 973
rect 10565 831 10599 923
rect 9432 219 9466 316
rect 9660 313 9728 353
rect 9660 279 9677 313
rect 9711 279 9728 313
rect 9432 169 9466 185
rect 9529 263 9563 279
rect 9529 195 9563 229
rect 9221 125 9255 141
rect 9061 91 9124 125
rect 9158 91 9221 125
rect 9027 75 9061 91
rect 9221 75 9255 91
rect 9335 125 9369 161
rect 9529 125 9563 161
rect 9369 91 9432 125
rect 9466 91 9529 125
rect 9335 75 9369 91
rect 9529 75 9563 91
rect 9660 239 9728 279
rect 9660 205 9677 239
rect 9711 205 9728 239
rect 9660 165 9728 205
rect 9660 131 9677 165
rect 9711 131 9728 165
rect 9660 91 9728 131
rect 9660 57 9677 91
rect 9711 57 9728 91
rect 9816 333 9850 349
rect 10010 333 10044 349
rect 10195 348 10229 649
rect 9850 299 9913 333
rect 9947 299 10010 333
rect 9816 261 9850 299
rect 9816 193 9850 227
rect 10010 261 10044 299
rect 9816 123 9850 159
rect 9816 73 9850 89
rect 9913 208 9947 224
rect 9660 34 9728 57
rect 9913 34 9947 174
rect 10010 193 10044 227
rect 10107 314 10229 348
rect 10326 461 10394 544
rect 10326 427 10343 461
rect 10377 427 10394 461
rect 10326 387 10394 427
rect 10326 353 10343 387
rect 10377 353 10394 387
rect 10565 433 10599 797
rect 10565 383 10599 399
rect 10787 957 10821 973
rect 10787 905 10821 923
rect 10787 433 10821 871
rect 10787 383 10821 399
rect 11009 957 11043 973
rect 11009 683 11043 923
rect 11009 433 11043 649
rect 11009 383 11043 399
rect 11157 757 11191 1014
rect 11288 1019 11305 1053
rect 11339 1019 11356 1053
rect 11523 1366 11557 1446
rect 11523 1298 11557 1332
rect 11523 1230 11557 1264
rect 11523 1162 11557 1196
rect 11523 1093 11557 1128
rect 11523 1043 11557 1059
rect 11611 1366 11645 1404
rect 11611 1298 11645 1332
rect 11611 1230 11645 1264
rect 11611 1162 11645 1196
rect 11611 1093 11645 1128
rect 11699 1366 11733 1446
rect 11699 1298 11733 1332
rect 11699 1230 11733 1264
rect 11699 1162 11733 1196
rect 11699 1111 11733 1128
rect 11787 1366 11821 1404
rect 11787 1298 11821 1332
rect 11787 1230 11821 1264
rect 11787 1162 11821 1196
rect 11611 1048 11645 1059
rect 11787 1093 11821 1128
rect 11875 1366 11909 1446
rect 11875 1298 11909 1332
rect 11875 1230 11909 1264
rect 11875 1162 11909 1196
rect 11875 1111 11909 1128
rect 11963 1366 11997 1404
rect 11963 1298 11997 1332
rect 11963 1230 11997 1264
rect 11963 1162 11997 1196
rect 11787 1048 11821 1059
rect 11963 1093 11997 1128
rect 12051 1366 12085 1446
rect 12051 1298 12085 1332
rect 12051 1230 12085 1264
rect 12051 1162 12085 1196
rect 12051 1111 12085 1128
rect 12250 1423 12318 1446
rect 12250 1389 12267 1423
rect 12301 1389 12318 1423
rect 12250 1349 12318 1389
rect 12250 1315 12267 1349
rect 12301 1315 12318 1349
rect 12250 1275 12318 1315
rect 12250 1241 12267 1275
rect 12301 1241 12318 1275
rect 12250 1201 12318 1241
rect 12250 1167 12267 1201
rect 12301 1167 12318 1201
rect 12250 1127 12318 1167
rect 11963 1048 11997 1059
rect 12250 1093 12267 1127
rect 12301 1093 12318 1127
rect 12250 1053 12318 1093
rect 11288 979 11356 1019
rect 11611 1014 12153 1048
rect 11288 945 11305 979
rect 11339 945 11356 979
rect 11288 905 11356 945
rect 11288 871 11305 905
rect 11339 871 11356 905
rect 11288 822 11356 871
rect 11527 957 11561 973
rect 10107 217 10141 314
rect 10326 313 10394 353
rect 10326 279 10343 313
rect 10377 279 10394 313
rect 10107 167 10141 183
rect 10204 261 10238 277
rect 10204 193 10238 227
rect 10010 123 10044 159
rect 10204 123 10238 159
rect 10044 89 10107 123
rect 10141 89 10204 123
rect 10010 73 10044 89
rect 10204 73 10238 89
rect 10326 239 10394 279
rect 10326 205 10343 239
rect 10377 205 10394 239
rect 10326 165 10394 205
rect 10326 131 10343 165
rect 10377 131 10394 165
rect 10326 91 10394 131
rect 10326 57 10343 91
rect 10377 57 10394 91
rect 10461 335 10495 351
rect 10655 335 10689 351
rect 10849 335 10883 351
rect 10495 301 10558 335
rect 10592 301 10655 335
rect 10689 301 10752 335
rect 10786 301 10849 335
rect 10461 263 10495 301
rect 10461 195 10495 229
rect 10655 263 10689 301
rect 10849 285 10883 301
rect 10963 335 10997 351
rect 11157 350 11191 723
rect 11527 757 11561 923
rect 10963 263 10997 301
rect 10461 125 10495 161
rect 10461 75 10495 91
rect 10558 210 10592 226
rect 10326 34 10394 57
rect 10558 34 10592 176
rect 10655 195 10689 229
rect 10753 216 10787 232
rect 10963 216 10997 229
rect 10787 195 10997 216
rect 10787 182 10963 195
rect 10753 166 10787 182
rect 10655 125 10689 161
rect 11060 316 11191 350
rect 11288 461 11356 544
rect 11288 427 11305 461
rect 11339 427 11356 461
rect 11288 387 11356 427
rect 11288 353 11305 387
rect 11339 353 11356 387
rect 11527 433 11561 723
rect 11527 383 11561 399
rect 11749 957 11783 973
rect 11749 535 11783 923
rect 11749 433 11783 501
rect 11749 383 11783 399
rect 11971 957 12005 973
rect 11971 461 12005 923
rect 11971 383 12005 399
rect 12119 683 12153 1014
rect 12250 1019 12267 1053
rect 12301 1019 12318 1053
rect 12425 1366 12459 1446
rect 12425 1298 12459 1332
rect 12425 1230 12459 1264
rect 12425 1162 12459 1196
rect 12425 1093 12459 1128
rect 12425 1027 12459 1059
rect 12513 1366 12547 1404
rect 12513 1298 12547 1332
rect 12513 1230 12547 1264
rect 12513 1162 12547 1196
rect 12513 1093 12547 1128
rect 12601 1366 12635 1446
rect 12601 1298 12635 1332
rect 12601 1230 12635 1264
rect 12601 1162 12635 1196
rect 12601 1111 12635 1128
rect 12689 1366 12723 1404
rect 12689 1298 12723 1332
rect 12689 1230 12723 1264
rect 12689 1162 12723 1196
rect 12513 1057 12547 1059
rect 12689 1093 12723 1128
rect 12777 1366 12811 1446
rect 12777 1298 12811 1332
rect 12777 1230 12811 1264
rect 12777 1162 12811 1196
rect 12777 1111 12811 1128
rect 12916 1423 12984 1446
rect 12916 1389 12933 1423
rect 12967 1389 12984 1423
rect 12916 1349 12984 1389
rect 12916 1315 12933 1349
rect 12967 1315 12984 1349
rect 12916 1275 12984 1315
rect 12916 1241 12933 1275
rect 12967 1241 12984 1275
rect 12916 1201 12984 1241
rect 12916 1167 12933 1201
rect 12967 1167 12984 1201
rect 12916 1127 12984 1167
rect 12689 1057 12723 1059
rect 12916 1093 12933 1127
rect 12967 1093 12984 1127
rect 12513 1023 12819 1057
rect 12250 979 12318 1019
rect 12250 945 12267 979
rect 12301 945 12318 979
rect 12250 905 12318 945
rect 12250 871 12267 905
rect 12301 871 12318 905
rect 12250 822 12318 871
rect 12489 957 12523 973
rect 12643 957 12677 973
rect 11060 219 11094 316
rect 11288 313 11356 353
rect 11288 279 11305 313
rect 11339 279 11356 313
rect 11060 169 11094 185
rect 11157 263 11191 279
rect 11157 195 11191 229
rect 10849 125 10883 141
rect 10689 91 10752 125
rect 10786 91 10849 125
rect 10655 75 10689 91
rect 10849 75 10883 91
rect 10963 125 10997 161
rect 11157 125 11191 161
rect 10997 91 11060 125
rect 11094 91 11157 125
rect 10963 75 10997 91
rect 11157 75 11191 91
rect 11288 239 11356 279
rect 11288 205 11305 239
rect 11339 205 11356 239
rect 11288 165 11356 205
rect 11288 131 11305 165
rect 11339 131 11356 165
rect 11288 91 11356 131
rect 11288 57 11305 91
rect 11339 57 11356 91
rect 11423 335 11457 351
rect 11617 335 11651 351
rect 11811 335 11845 351
rect 11457 301 11520 335
rect 11554 301 11617 335
rect 11651 301 11714 335
rect 11748 301 11811 335
rect 11423 263 11457 301
rect 11423 195 11457 229
rect 11617 263 11651 301
rect 11811 285 11845 301
rect 11925 335 11959 351
rect 12119 350 12153 649
rect 12489 683 12523 923
rect 11925 263 11959 301
rect 11423 125 11457 161
rect 11423 75 11457 91
rect 11520 210 11554 226
rect 11288 34 11356 57
rect 11520 34 11554 176
rect 11617 195 11651 229
rect 11715 216 11749 232
rect 11925 216 11959 229
rect 11749 195 11959 216
rect 11749 182 11925 195
rect 11715 166 11749 182
rect 11617 125 11651 161
rect 12022 316 12153 350
rect 12250 461 12318 544
rect 12250 427 12267 461
rect 12301 427 12318 461
rect 12250 387 12318 427
rect 12250 353 12267 387
rect 12301 353 12318 387
rect 12489 433 12523 649
rect 12489 383 12523 399
rect 12637 923 12643 942
rect 12637 907 12677 923
rect 12637 831 12671 907
rect 12637 433 12671 797
rect 12637 383 12671 399
rect 12785 683 12819 1023
rect 12916 1053 12984 1093
rect 12916 1019 12933 1053
rect 12967 1019 12984 1053
rect 13151 1366 13185 1446
rect 13151 1298 13185 1332
rect 13151 1230 13185 1264
rect 13151 1162 13185 1196
rect 13151 1093 13185 1128
rect 13151 1043 13185 1059
rect 13239 1366 13273 1404
rect 13239 1298 13273 1332
rect 13239 1230 13273 1264
rect 13239 1162 13273 1196
rect 13239 1093 13273 1128
rect 13327 1366 13361 1446
rect 13327 1298 13361 1332
rect 13327 1230 13361 1264
rect 13327 1162 13361 1196
rect 13327 1111 13361 1128
rect 13415 1366 13449 1404
rect 13415 1298 13449 1332
rect 13415 1230 13449 1264
rect 13415 1162 13449 1196
rect 13239 1048 13273 1059
rect 13415 1093 13449 1128
rect 13503 1366 13537 1446
rect 13503 1298 13537 1332
rect 13503 1230 13537 1264
rect 13503 1162 13537 1196
rect 13503 1111 13537 1128
rect 13591 1366 13625 1404
rect 13591 1298 13625 1332
rect 13591 1230 13625 1264
rect 13591 1162 13625 1196
rect 13415 1048 13449 1059
rect 13591 1093 13625 1128
rect 13679 1366 13713 1446
rect 13679 1298 13713 1332
rect 13679 1230 13713 1264
rect 13679 1162 13713 1196
rect 13679 1111 13713 1128
rect 13878 1423 13946 1446
rect 13878 1389 13895 1423
rect 13929 1389 13946 1423
rect 13878 1349 13946 1389
rect 13878 1315 13895 1349
rect 13929 1315 13946 1349
rect 13878 1275 13946 1315
rect 13878 1241 13895 1275
rect 13929 1241 13946 1275
rect 13878 1201 13946 1241
rect 13878 1167 13895 1201
rect 13929 1167 13946 1201
rect 13878 1127 13946 1167
rect 13591 1048 13625 1059
rect 13878 1093 13895 1127
rect 13929 1093 13946 1127
rect 13878 1053 13946 1093
rect 12916 979 12984 1019
rect 13239 1014 13781 1048
rect 12916 945 12933 979
rect 12967 945 12984 979
rect 12916 905 12984 945
rect 12916 871 12933 905
rect 12967 871 12984 905
rect 12916 822 12984 871
rect 13155 957 13189 973
rect 12022 219 12056 316
rect 12250 313 12318 353
rect 12250 279 12267 313
rect 12301 279 12318 313
rect 12022 169 12056 185
rect 12119 263 12153 279
rect 12119 195 12153 229
rect 11811 125 11845 141
rect 11651 91 11714 125
rect 11748 91 11811 125
rect 11617 75 11651 91
rect 11811 75 11845 91
rect 11925 125 11959 161
rect 12119 125 12153 161
rect 11959 91 12022 125
rect 12056 91 12119 125
rect 11925 75 11959 91
rect 12119 75 12153 91
rect 12250 239 12318 279
rect 12250 205 12267 239
rect 12301 205 12318 239
rect 12250 165 12318 205
rect 12250 131 12267 165
rect 12301 131 12318 165
rect 12250 91 12318 131
rect 12250 57 12267 91
rect 12301 57 12318 91
rect 12406 333 12440 349
rect 12600 333 12634 349
rect 12785 348 12819 649
rect 13155 683 13189 923
rect 12440 299 12503 333
rect 12537 299 12600 333
rect 12406 261 12440 299
rect 12406 193 12440 227
rect 12600 261 12634 299
rect 12406 123 12440 159
rect 12406 73 12440 89
rect 12503 208 12537 224
rect 12250 34 12318 57
rect 12503 34 12537 174
rect 12600 193 12634 227
rect 12697 314 12819 348
rect 12916 461 12984 544
rect 12916 427 12933 461
rect 12967 427 12984 461
rect 12916 387 12984 427
rect 12916 353 12933 387
rect 12967 353 12984 387
rect 13155 433 13189 649
rect 13155 383 13189 399
rect 13377 957 13411 973
rect 13377 905 13411 923
rect 13377 433 13411 871
rect 13377 383 13411 399
rect 13599 957 13633 973
rect 13599 461 13633 923
rect 13599 383 13633 399
rect 13747 831 13781 1014
rect 13878 1019 13895 1053
rect 13929 1019 13946 1053
rect 14113 1366 14147 1446
rect 14113 1298 14147 1332
rect 14113 1230 14147 1264
rect 14113 1162 14147 1196
rect 14113 1093 14147 1128
rect 14113 1043 14147 1059
rect 14201 1366 14235 1404
rect 14201 1298 14235 1332
rect 14201 1230 14235 1264
rect 14201 1162 14235 1196
rect 14201 1093 14235 1128
rect 14289 1366 14323 1446
rect 14289 1298 14323 1332
rect 14289 1230 14323 1264
rect 14289 1162 14323 1196
rect 14289 1111 14323 1128
rect 14377 1366 14411 1404
rect 14377 1298 14411 1332
rect 14377 1230 14411 1264
rect 14377 1162 14411 1196
rect 14201 1048 14235 1059
rect 14377 1093 14411 1128
rect 14465 1366 14499 1446
rect 14465 1298 14499 1332
rect 14465 1230 14499 1264
rect 14465 1162 14499 1196
rect 14465 1111 14499 1128
rect 14553 1366 14587 1404
rect 14553 1298 14587 1332
rect 14553 1230 14587 1264
rect 14553 1162 14587 1196
rect 14377 1048 14411 1059
rect 14553 1093 14587 1128
rect 14641 1366 14675 1446
rect 14641 1298 14675 1332
rect 14641 1230 14675 1264
rect 14641 1162 14675 1196
rect 14641 1111 14675 1128
rect 14840 1423 14908 1446
rect 14840 1389 14857 1423
rect 14891 1389 14908 1423
rect 14840 1349 14908 1389
rect 14840 1315 14857 1349
rect 14891 1315 14908 1349
rect 14840 1275 14908 1315
rect 14840 1241 14857 1275
rect 14891 1241 14908 1275
rect 14840 1201 14908 1241
rect 14840 1167 14857 1201
rect 14891 1167 14908 1201
rect 14840 1127 14908 1167
rect 14553 1048 14587 1059
rect 14840 1093 14857 1127
rect 14891 1093 14908 1127
rect 14840 1053 14908 1093
rect 13878 979 13946 1019
rect 14201 1014 14743 1048
rect 13878 945 13895 979
rect 13929 945 13946 979
rect 13878 905 13946 945
rect 13878 871 13895 905
rect 13929 871 13946 905
rect 13878 822 13946 871
rect 14117 957 14151 973
rect 12697 217 12731 314
rect 12916 313 12984 353
rect 12916 279 12933 313
rect 12967 279 12984 313
rect 12697 167 12731 183
rect 12794 261 12828 277
rect 12794 193 12828 227
rect 12600 123 12634 159
rect 12794 123 12828 159
rect 12634 89 12697 123
rect 12731 89 12794 123
rect 12600 73 12634 89
rect 12794 73 12828 89
rect 12916 239 12984 279
rect 12916 205 12933 239
rect 12967 205 12984 239
rect 12916 165 12984 205
rect 12916 131 12933 165
rect 12967 131 12984 165
rect 12916 91 12984 131
rect 12916 57 12933 91
rect 12967 57 12984 91
rect 13051 335 13085 351
rect 13245 335 13279 351
rect 13439 335 13473 351
rect 13085 301 13148 335
rect 13182 301 13245 335
rect 13279 301 13342 335
rect 13376 301 13439 335
rect 13051 263 13085 301
rect 13051 195 13085 229
rect 13245 263 13279 301
rect 13439 285 13473 301
rect 13553 335 13587 351
rect 13747 350 13781 797
rect 14117 757 14151 923
rect 13553 263 13587 301
rect 13051 125 13085 161
rect 13051 75 13085 91
rect 13148 210 13182 226
rect 12916 34 12984 57
rect 13148 34 13182 176
rect 13245 195 13279 229
rect 13343 216 13377 232
rect 13553 216 13587 229
rect 13377 195 13587 216
rect 13377 182 13553 195
rect 13343 166 13377 182
rect 13245 125 13279 161
rect 13650 316 13781 350
rect 13878 461 13946 544
rect 13878 427 13895 461
rect 13929 427 13946 461
rect 13878 387 13946 427
rect 13878 353 13895 387
rect 13929 353 13946 387
rect 14117 433 14151 723
rect 14117 383 14151 399
rect 14339 957 14373 973
rect 14339 461 14373 923
rect 14339 383 14373 399
rect 14561 957 14595 973
rect 14561 757 14595 923
rect 14561 433 14595 723
rect 14561 383 14595 399
rect 14709 831 14743 1014
rect 14840 1019 14857 1053
rect 14891 1019 14908 1053
rect 15015 1366 15049 1446
rect 15015 1298 15049 1332
rect 15015 1230 15049 1264
rect 15015 1162 15049 1196
rect 15015 1093 15049 1128
rect 15015 1027 15049 1059
rect 15103 1366 15137 1404
rect 15103 1298 15137 1332
rect 15103 1230 15137 1264
rect 15103 1162 15137 1196
rect 15103 1093 15137 1128
rect 15191 1366 15225 1446
rect 15191 1298 15225 1332
rect 15191 1230 15225 1264
rect 15191 1162 15225 1196
rect 15191 1111 15225 1128
rect 15279 1366 15313 1404
rect 15279 1298 15313 1332
rect 15279 1230 15313 1264
rect 15279 1162 15313 1196
rect 15103 1057 15137 1059
rect 15279 1093 15313 1128
rect 15367 1366 15401 1446
rect 15367 1298 15401 1332
rect 15367 1230 15401 1264
rect 15367 1162 15401 1196
rect 15367 1111 15401 1128
rect 15506 1423 15574 1446
rect 15506 1389 15523 1423
rect 15557 1389 15574 1423
rect 15506 1349 15574 1389
rect 15506 1315 15523 1349
rect 15557 1315 15574 1349
rect 15506 1275 15574 1315
rect 15506 1241 15523 1275
rect 15557 1241 15574 1275
rect 15506 1201 15574 1241
rect 15506 1167 15523 1201
rect 15557 1167 15574 1201
rect 15506 1127 15574 1167
rect 15279 1057 15313 1059
rect 15506 1093 15523 1127
rect 15557 1093 15574 1127
rect 15103 1023 15409 1057
rect 14840 979 14908 1019
rect 14840 945 14857 979
rect 14891 945 14908 979
rect 14840 905 14908 945
rect 14840 871 14857 905
rect 14891 871 14908 905
rect 14840 822 14908 871
rect 15079 957 15113 973
rect 15233 957 15267 973
rect 15079 831 15113 923
rect 13650 219 13684 316
rect 13878 313 13946 353
rect 13878 279 13895 313
rect 13929 279 13946 313
rect 13650 169 13684 185
rect 13747 263 13781 279
rect 13747 195 13781 229
rect 13439 125 13473 141
rect 13279 91 13342 125
rect 13376 91 13439 125
rect 13245 75 13279 91
rect 13439 75 13473 91
rect 13553 125 13587 161
rect 13747 125 13781 161
rect 13587 91 13650 125
rect 13684 91 13747 125
rect 13553 75 13587 91
rect 13747 75 13781 91
rect 13878 239 13946 279
rect 13878 205 13895 239
rect 13929 205 13946 239
rect 13878 165 13946 205
rect 13878 131 13895 165
rect 13929 131 13946 165
rect 13878 91 13946 131
rect 13878 57 13895 91
rect 13929 57 13946 91
rect 14013 335 14047 351
rect 14207 335 14241 351
rect 14401 335 14435 351
rect 14047 301 14110 335
rect 14144 301 14207 335
rect 14241 301 14304 335
rect 14338 301 14401 335
rect 14013 263 14047 301
rect 14013 195 14047 229
rect 14207 263 14241 301
rect 14401 285 14435 301
rect 14515 335 14549 351
rect 14709 350 14743 797
rect 14515 263 14549 301
rect 14013 125 14047 161
rect 14013 75 14047 91
rect 14110 210 14144 226
rect 13878 34 13946 57
rect 14110 34 14144 176
rect 14207 195 14241 229
rect 14305 216 14339 232
rect 14515 216 14549 229
rect 14339 195 14549 216
rect 14339 182 14515 195
rect 14305 166 14339 182
rect 14207 125 14241 161
rect 14612 316 14743 350
rect 14840 461 14908 544
rect 14840 427 14857 461
rect 14891 427 14908 461
rect 14840 387 14908 427
rect 14840 353 14857 387
rect 14891 353 14908 387
rect 15079 433 15113 797
rect 15079 383 15113 399
rect 15227 923 15233 942
rect 15227 907 15267 923
rect 15227 831 15261 907
rect 15227 433 15261 797
rect 15227 383 15261 399
rect 15375 757 15409 1023
rect 15506 1053 15574 1093
rect 15506 1019 15523 1053
rect 15557 1019 15574 1053
rect 15681 1365 15715 1446
rect 15681 1297 15715 1331
rect 15681 1229 15715 1263
rect 15681 1161 15715 1195
rect 15681 1093 15715 1127
rect 15681 1025 15715 1059
rect 15769 1365 15805 1399
rect 15857 1365 15891 1446
rect 15769 1297 15803 1331
rect 15769 1229 15803 1263
rect 15769 1161 15803 1195
rect 15769 1093 15803 1127
rect 15857 1297 15891 1331
rect 15857 1229 15891 1263
rect 15857 1161 15891 1195
rect 15857 1111 15891 1127
rect 15945 1365 15979 1399
rect 15945 1297 15979 1331
rect 15945 1229 15979 1263
rect 15945 1161 15979 1195
rect 15945 1059 15979 1127
rect 15769 1025 15945 1059
rect 16033 1365 16067 1446
rect 16033 1297 16067 1331
rect 16033 1229 16067 1263
rect 16033 1161 16067 1195
rect 16033 1093 16067 1127
rect 16033 1025 16067 1059
rect 16172 1423 16240 1446
rect 16172 1389 16189 1423
rect 16223 1389 16240 1423
rect 16838 1423 16906 1446
rect 16172 1349 16240 1389
rect 16172 1315 16189 1349
rect 16223 1315 16240 1349
rect 16172 1275 16240 1315
rect 16172 1241 16189 1275
rect 16223 1241 16240 1275
rect 16172 1201 16240 1241
rect 16172 1167 16189 1201
rect 16223 1167 16240 1201
rect 16172 1127 16240 1167
rect 16172 1093 16189 1127
rect 16223 1093 16240 1127
rect 16172 1053 16240 1093
rect 15506 979 15574 1019
rect 15945 1009 15979 1025
rect 16172 1019 16189 1053
rect 16223 1019 16240 1053
rect 15506 945 15523 979
rect 15557 945 15574 979
rect 16172 979 16240 1019
rect 16345 1365 16731 1399
rect 16345 1297 16379 1331
rect 16345 1229 16379 1263
rect 16345 1161 16379 1195
rect 16345 1059 16379 1127
rect 16433 1297 16467 1313
rect 16433 1229 16467 1263
rect 16433 1161 16467 1195
rect 16433 1093 16467 1127
rect 16521 1297 16555 1331
rect 16521 1229 16555 1263
rect 16521 1161 16555 1195
rect 16521 1111 16555 1127
rect 16609 1297 16643 1313
rect 16609 1229 16643 1263
rect 16609 1161 16643 1195
rect 16609 1059 16643 1127
rect 16697 1297 16731 1331
rect 16697 1229 16731 1263
rect 16697 1161 16731 1195
rect 16697 1075 16731 1127
rect 16838 1389 16855 1423
rect 16889 1389 16906 1423
rect 17504 1423 17572 1446
rect 16838 1349 16906 1389
rect 16838 1315 16855 1349
rect 16889 1315 16906 1349
rect 16838 1275 16906 1315
rect 16838 1241 16855 1275
rect 16889 1241 16906 1275
rect 16838 1201 16906 1241
rect 16838 1167 16855 1201
rect 16889 1167 16906 1201
rect 16838 1127 16906 1167
rect 16838 1093 16855 1127
rect 16889 1093 16906 1127
rect 16433 1025 16609 1059
rect 16345 1009 16379 1025
rect 16609 1009 16643 1025
rect 16838 1053 16906 1093
rect 16838 1019 16855 1053
rect 16889 1019 16906 1053
rect 15506 905 15574 945
rect 15506 871 15523 905
rect 15557 871 15574 905
rect 15506 822 15574 871
rect 15671 958 15705 974
rect 15901 958 15935 974
rect 15671 905 15705 924
rect 14612 219 14646 316
rect 14840 313 14908 353
rect 14840 279 14857 313
rect 14891 279 14908 313
rect 14612 169 14646 185
rect 14709 263 14743 279
rect 14709 195 14743 229
rect 14401 125 14435 141
rect 14241 91 14304 125
rect 14338 91 14401 125
rect 14207 75 14241 91
rect 14401 75 14435 91
rect 14515 125 14549 161
rect 14709 125 14743 161
rect 14549 91 14612 125
rect 14646 91 14709 125
rect 14515 75 14549 91
rect 14709 75 14743 91
rect 14840 239 14908 279
rect 14840 205 14857 239
rect 14891 205 14908 239
rect 14840 165 14908 205
rect 14840 131 14857 165
rect 14891 131 14908 165
rect 14840 91 14908 131
rect 14840 57 14857 91
rect 14891 57 14908 91
rect 14996 333 15030 349
rect 15190 333 15224 349
rect 15375 348 15409 723
rect 15671 683 15705 871
rect 15030 299 15093 333
rect 15127 299 15190 333
rect 14996 261 15030 299
rect 14996 193 15030 227
rect 15190 261 15224 299
rect 14996 123 15030 159
rect 14996 73 15030 89
rect 15093 208 15127 224
rect 14840 34 14908 57
rect 15093 34 15127 174
rect 15190 193 15224 227
rect 15287 314 15409 348
rect 15506 461 15574 544
rect 15506 427 15523 461
rect 15557 427 15574 461
rect 15506 387 15574 427
rect 15506 353 15523 387
rect 15557 353 15574 387
rect 15671 433 15705 649
rect 15671 383 15705 399
rect 15893 924 15901 942
rect 15893 908 15935 924
rect 16172 945 16189 979
rect 16223 945 16240 979
rect 16838 979 16906 1019
rect 17013 1365 17399 1399
rect 17013 1297 17047 1331
rect 17013 1229 17047 1263
rect 17013 1161 17047 1195
rect 17013 1059 17047 1127
rect 17101 1297 17135 1313
rect 17101 1229 17135 1263
rect 17101 1161 17135 1195
rect 17101 1093 17135 1127
rect 17189 1297 17223 1331
rect 17189 1229 17223 1263
rect 17189 1161 17223 1195
rect 17189 1111 17223 1127
rect 17277 1297 17311 1313
rect 17277 1229 17311 1263
rect 17277 1161 17311 1195
rect 17277 1093 17311 1127
rect 17365 1297 17399 1331
rect 17365 1229 17399 1263
rect 17365 1161 17399 1195
rect 17365 1111 17399 1127
rect 17504 1389 17521 1423
rect 17555 1389 17572 1423
rect 17504 1349 17572 1389
rect 17504 1315 17521 1349
rect 17555 1315 17572 1349
rect 17504 1275 17572 1315
rect 17504 1241 17521 1275
rect 17555 1241 17572 1275
rect 17504 1201 17572 1241
rect 17504 1167 17521 1201
rect 17555 1167 17572 1201
rect 17504 1127 17572 1167
rect 17504 1093 17521 1127
rect 17555 1093 17572 1127
rect 17101 1025 17407 1059
rect 17013 1009 17047 1025
rect 15893 831 15927 908
rect 16172 905 16240 945
rect 16172 871 16189 905
rect 16223 871 16240 905
rect 16172 822 16240 871
rect 16411 958 16445 974
rect 16411 905 16445 924
rect 15893 757 15927 797
rect 15893 433 15927 723
rect 15893 383 15927 399
rect 16172 461 16240 544
rect 16172 427 16189 461
rect 16223 427 16240 461
rect 16172 387 16240 427
rect 15287 217 15321 314
rect 15506 313 15574 353
rect 16172 353 16189 387
rect 16223 353 16240 387
rect 16411 433 16445 871
rect 16411 383 16445 399
rect 16707 958 16741 974
rect 16707 609 16741 924
rect 16838 945 16855 979
rect 16889 945 16906 979
rect 16838 905 16906 945
rect 16838 871 16855 905
rect 16889 871 16906 905
rect 16838 822 16906 871
rect 17003 958 17037 974
rect 16707 433 16741 575
rect 16707 383 16741 399
rect 16838 461 16906 544
rect 16838 427 16855 461
rect 16889 427 16906 461
rect 16838 387 16906 427
rect 15506 279 15523 313
rect 15557 279 15574 313
rect 15287 167 15321 183
rect 15384 261 15418 277
rect 15384 193 15418 227
rect 15190 123 15224 159
rect 15384 123 15418 159
rect 15224 89 15287 123
rect 15321 89 15384 123
rect 15190 73 15224 89
rect 15384 73 15418 89
rect 15506 239 15574 279
rect 15506 205 15523 239
rect 15557 205 15574 239
rect 15506 165 15574 205
rect 15506 131 15523 165
rect 15557 131 15574 165
rect 15506 91 15574 131
rect 15506 57 15523 91
rect 15557 57 15574 91
rect 15662 333 15696 349
rect 15856 333 15890 349
rect 15696 299 15759 333
rect 15793 299 15856 333
rect 15662 261 15696 299
rect 15662 193 15696 227
rect 15856 261 15890 299
rect 16050 333 16084 349
rect 15953 253 15987 269
rect 15662 123 15696 159
rect 15662 73 15696 89
rect 15759 208 15793 224
rect 15506 34 15574 57
rect 15759 34 15793 174
rect 15856 193 15890 227
rect 15952 219 15953 234
rect 15952 217 15987 219
rect 15986 203 15987 217
rect 16050 261 16084 299
rect 15952 167 15986 183
rect 16050 193 16084 227
rect 15856 123 15890 159
rect 16050 123 16084 159
rect 15890 89 15952 123
rect 15986 89 16050 123
rect 15856 73 15890 89
rect 16050 73 16084 89
rect 16172 313 16240 353
rect 16838 353 16855 387
rect 16889 353 16906 387
rect 17003 433 17037 924
rect 17003 383 17037 399
rect 17225 958 17263 974
rect 17225 924 17229 958
rect 17225 908 17263 924
rect 17225 831 17259 908
rect 17225 433 17259 797
rect 17225 383 17259 399
rect 17373 831 17407 1025
rect 17504 1053 17572 1093
rect 17504 1019 17521 1053
rect 17555 1019 17572 1053
rect 17656 1366 17690 1446
rect 17656 1298 17690 1332
rect 17656 1230 17690 1264
rect 17656 1162 17690 1196
rect 17656 1093 17690 1128
rect 17656 1037 17690 1059
rect 17744 1366 17778 1404
rect 17744 1298 17778 1332
rect 17744 1230 17778 1264
rect 17744 1162 17778 1196
rect 17744 1093 17778 1128
rect 17504 979 17572 1019
rect 17504 945 17521 979
rect 17555 945 17572 979
rect 17504 905 17572 945
rect 17504 871 17521 905
rect 17555 871 17572 905
rect 17504 822 17572 871
rect 17669 957 17703 973
rect 17669 831 17703 923
rect 17744 933 17778 1059
rect 17832 1366 17866 1446
rect 17832 1298 17866 1332
rect 17832 1230 17866 1264
rect 17832 1162 17866 1196
rect 17832 1093 17866 1128
rect 17832 1037 17866 1059
rect 17948 1423 18016 1446
rect 17948 1389 17965 1423
rect 17999 1389 18016 1423
rect 17948 1349 18016 1389
rect 17948 1315 17965 1349
rect 17999 1315 18016 1349
rect 17948 1275 18016 1315
rect 17948 1241 17965 1275
rect 17999 1241 18016 1275
rect 17948 1201 18016 1241
rect 17948 1167 17965 1201
rect 17999 1167 18016 1201
rect 17948 1127 18016 1167
rect 17948 1093 17965 1127
rect 17999 1093 18016 1127
rect 17948 1053 18016 1093
rect 17948 1019 17965 1053
rect 17999 1019 18016 1053
rect 17948 979 18016 1019
rect 17948 945 17965 979
rect 17999 945 18016 979
rect 17744 899 17851 933
rect 16172 279 16189 313
rect 16223 279 16240 313
rect 16172 239 16240 279
rect 16172 205 16189 239
rect 16223 205 16240 239
rect 16172 165 16240 205
rect 16172 131 16189 165
rect 16223 131 16240 165
rect 16172 91 16240 131
rect 16172 57 16189 91
rect 16223 57 16240 91
rect 16328 333 16362 349
rect 16522 333 16556 349
rect 16362 299 16425 333
rect 16459 299 16522 333
rect 16328 261 16362 299
rect 16328 193 16362 227
rect 16522 261 16556 299
rect 16716 333 16750 349
rect 16328 123 16362 159
rect 16328 73 16362 89
rect 16425 208 16459 224
rect 16172 34 16240 57
rect 16425 34 16459 174
rect 16522 193 16556 227
rect 16619 253 16653 269
rect 16619 217 16653 219
rect 16619 167 16653 183
rect 16716 261 16750 299
rect 16716 193 16750 227
rect 16522 123 16556 159
rect 16716 123 16750 159
rect 16556 89 16619 123
rect 16653 89 16716 123
rect 16522 73 16556 89
rect 16716 73 16750 89
rect 16838 313 16906 353
rect 16838 279 16855 313
rect 16889 279 16906 313
rect 16838 239 16906 279
rect 16838 205 16855 239
rect 16889 205 16906 239
rect 16838 165 16906 205
rect 16838 131 16855 165
rect 16889 131 16906 165
rect 16838 91 16906 131
rect 16838 57 16855 91
rect 16889 57 16906 91
rect 16994 333 17028 349
rect 17188 333 17222 349
rect 17373 346 17407 797
rect 17028 299 17091 333
rect 17125 299 17188 333
rect 16994 261 17028 299
rect 16994 193 17028 227
rect 17188 261 17222 299
rect 16994 123 17028 159
rect 16994 73 17028 89
rect 17091 208 17125 224
rect 16838 34 16906 57
rect 17091 34 17125 174
rect 17188 193 17222 227
rect 17285 312 17407 346
rect 17504 461 17572 544
rect 17504 427 17521 461
rect 17555 427 17572 461
rect 17504 387 17572 427
rect 17504 353 17521 387
rect 17555 353 17572 387
rect 17669 434 17703 797
rect 17817 433 17851 899
rect 17948 905 18016 945
rect 17948 871 17965 905
rect 17999 871 18016 905
rect 17948 822 18016 871
rect 17669 384 17703 400
rect 17743 399 17851 433
rect 17948 461 18016 544
rect 17948 427 17965 461
rect 17999 427 18016 461
rect 17504 313 17572 353
rect 17285 253 17319 312
rect 17504 279 17521 313
rect 17555 279 17572 313
rect 17285 217 17319 219
rect 17285 167 17319 183
rect 17382 261 17416 278
rect 17382 193 17416 227
rect 17188 123 17222 159
rect 17382 123 17416 159
rect 17222 89 17285 123
rect 17319 89 17382 123
rect 17188 73 17222 89
rect 17382 73 17416 89
rect 17504 239 17572 279
rect 17504 205 17521 239
rect 17555 205 17572 239
rect 17504 165 17572 205
rect 17504 131 17521 165
rect 17555 131 17572 165
rect 17504 91 17572 131
rect 17504 57 17521 91
rect 17555 57 17572 91
rect 17504 34 17572 57
rect 17647 334 17681 350
rect 17647 262 17681 300
rect 17647 194 17681 228
rect 17743 218 17777 399
rect 17948 387 18016 427
rect 17948 353 17965 387
rect 17999 353 18016 387
rect 17743 168 17777 184
rect 17841 334 17875 350
rect 17841 262 17875 300
rect 17841 194 17875 228
rect 17647 124 17681 160
rect 17841 124 17875 160
rect 17681 90 17743 124
rect 17777 90 17841 124
rect 17647 34 17681 90
rect 17744 34 17778 90
rect 17841 34 17875 90
rect 17948 313 18016 353
rect 17948 279 17965 313
rect 17999 279 18016 313
rect 17948 239 18016 279
rect 17948 205 17965 239
rect 17999 205 18016 239
rect 17948 165 18016 205
rect 17948 131 17965 165
rect 17999 131 18016 165
rect 17948 91 18016 131
rect 17948 57 17965 91
rect 17999 57 18016 91
rect 17948 34 18016 57
rect -34 17 18016 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5533 17
rect 5567 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5755 17
rect 5789 -17 5829 17
rect 5863 -17 5903 17
rect 5937 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6199 17
rect 6233 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6495 17
rect 6529 -17 6569 17
rect 6603 -17 6643 17
rect 6677 -17 6717 17
rect 6751 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7161 17
rect 7195 -17 7235 17
rect 7269 -17 7309 17
rect 7343 -17 7383 17
rect 7417 -17 7457 17
rect 7491 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7679 17
rect 7713 -17 7827 17
rect 7861 -17 7901 17
rect 7935 -17 7975 17
rect 8009 -17 8049 17
rect 8083 -17 8123 17
rect 8157 -17 8197 17
rect 8231 -17 8271 17
rect 8305 -17 8345 17
rect 8379 -17 8419 17
rect 8453 -17 8493 17
rect 8527 -17 8567 17
rect 8601 -17 8641 17
rect 8675 -17 8789 17
rect 8823 -17 8863 17
rect 8897 -17 8937 17
rect 8971 -17 9011 17
rect 9045 -17 9085 17
rect 9119 -17 9159 17
rect 9193 -17 9233 17
rect 9267 -17 9307 17
rect 9341 -17 9381 17
rect 9415 -17 9455 17
rect 9489 -17 9529 17
rect 9563 -17 9603 17
rect 9637 -17 9751 17
rect 9785 -17 9825 17
rect 9859 -17 9899 17
rect 9933 -17 9973 17
rect 10007 -17 10047 17
rect 10081 -17 10121 17
rect 10155 -17 10195 17
rect 10229 -17 10269 17
rect 10303 -17 10417 17
rect 10451 -17 10491 17
rect 10525 -17 10565 17
rect 10599 -17 10639 17
rect 10673 -17 10713 17
rect 10747 -17 10787 17
rect 10821 -17 10861 17
rect 10895 -17 10935 17
rect 10969 -17 11009 17
rect 11043 -17 11083 17
rect 11117 -17 11157 17
rect 11191 -17 11231 17
rect 11265 -17 11379 17
rect 11413 -17 11453 17
rect 11487 -17 11527 17
rect 11561 -17 11601 17
rect 11635 -17 11675 17
rect 11709 -17 11749 17
rect 11783 -17 11823 17
rect 11857 -17 11897 17
rect 11931 -17 11971 17
rect 12005 -17 12045 17
rect 12079 -17 12119 17
rect 12153 -17 12193 17
rect 12227 -17 12341 17
rect 12375 -17 12415 17
rect 12449 -17 12489 17
rect 12523 -17 12563 17
rect 12597 -17 12637 17
rect 12671 -17 12711 17
rect 12745 -17 12785 17
rect 12819 -17 12859 17
rect 12893 -17 13007 17
rect 13041 -17 13081 17
rect 13115 -17 13155 17
rect 13189 -17 13229 17
rect 13263 -17 13303 17
rect 13337 -17 13377 17
rect 13411 -17 13451 17
rect 13485 -17 13525 17
rect 13559 -17 13599 17
rect 13633 -17 13673 17
rect 13707 -17 13747 17
rect 13781 -17 13821 17
rect 13855 -17 13969 17
rect 14003 -17 14043 17
rect 14077 -17 14117 17
rect 14151 -17 14191 17
rect 14225 -17 14265 17
rect 14299 -17 14339 17
rect 14373 -17 14413 17
rect 14447 -17 14487 17
rect 14521 -17 14561 17
rect 14595 -17 14635 17
rect 14669 -17 14709 17
rect 14743 -17 14783 17
rect 14817 -17 14931 17
rect 14965 -17 15005 17
rect 15039 -17 15079 17
rect 15113 -17 15153 17
rect 15187 -17 15227 17
rect 15261 -17 15301 17
rect 15335 -17 15375 17
rect 15409 -17 15449 17
rect 15483 -17 15597 17
rect 15631 -17 15671 17
rect 15705 -17 15745 17
rect 15779 -17 15819 17
rect 15853 -17 15893 17
rect 15927 -17 15967 17
rect 16001 -17 16041 17
rect 16075 -17 16115 17
rect 16149 -17 16263 17
rect 16297 -17 16337 17
rect 16371 -17 16411 17
rect 16445 -17 16485 17
rect 16519 -17 16559 17
rect 16593 -17 16633 17
rect 16667 -17 16707 17
rect 16741 -17 16781 17
rect 16815 -17 16929 17
rect 16963 -17 17003 17
rect 17037 -17 17077 17
rect 17111 -17 17151 17
rect 17185 -17 17225 17
rect 17259 -17 17299 17
rect 17333 -17 17373 17
rect 17407 -17 17447 17
rect 17481 -17 17595 17
rect 17629 -17 17669 17
rect 17703 -17 17743 17
rect 17777 -17 17817 17
rect 17851 -17 17891 17
rect 17925 -17 18016 17
rect -34 -34 18016 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4793 1463 4827 1497
rect 4867 1463 4901 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5089 1463 5123 1497
rect 5237 1463 5271 1497
rect 5311 1463 5345 1497
rect 5385 1463 5419 1497
rect 5459 1463 5493 1497
rect 5533 1463 5567 1497
rect 5607 1463 5641 1497
rect 5681 1463 5715 1497
rect 5755 1463 5789 1497
rect 5829 1463 5863 1497
rect 5903 1463 5937 1497
rect 5977 1463 6011 1497
rect 6051 1463 6085 1497
rect 6199 1463 6233 1497
rect 6273 1463 6307 1497
rect 6347 1463 6381 1497
rect 6421 1463 6455 1497
rect 6495 1463 6529 1497
rect 6569 1463 6603 1497
rect 6643 1463 6677 1497
rect 6717 1463 6751 1497
rect 6791 1463 6825 1497
rect 6865 1463 6899 1497
rect 6939 1463 6973 1497
rect 7013 1463 7047 1497
rect 7161 1463 7195 1497
rect 7235 1463 7269 1497
rect 7309 1463 7343 1497
rect 7383 1463 7417 1497
rect 7457 1463 7491 1497
rect 7531 1463 7565 1497
rect 7605 1463 7639 1497
rect 7679 1463 7713 1497
rect 7827 1463 7861 1497
rect 7901 1463 7935 1497
rect 7975 1463 8009 1497
rect 8049 1463 8083 1497
rect 8123 1463 8157 1497
rect 8197 1463 8231 1497
rect 8271 1463 8305 1497
rect 8345 1463 8379 1497
rect 8419 1463 8453 1497
rect 8493 1463 8527 1497
rect 8567 1463 8601 1497
rect 8641 1463 8675 1497
rect 8789 1463 8823 1497
rect 8863 1463 8897 1497
rect 8937 1463 8971 1497
rect 9011 1463 9045 1497
rect 9085 1463 9119 1497
rect 9159 1463 9193 1497
rect 9233 1463 9267 1497
rect 9307 1463 9341 1497
rect 9381 1463 9415 1497
rect 9455 1463 9489 1497
rect 9529 1463 9563 1497
rect 9603 1463 9637 1497
rect 9751 1463 9785 1497
rect 9825 1463 9859 1497
rect 9899 1463 9933 1497
rect 9973 1463 10007 1497
rect 10047 1463 10081 1497
rect 10121 1463 10155 1497
rect 10195 1463 10229 1497
rect 10269 1463 10303 1497
rect 10417 1463 10451 1497
rect 10491 1463 10525 1497
rect 10565 1463 10599 1497
rect 10639 1463 10673 1497
rect 10713 1463 10747 1497
rect 10787 1463 10821 1497
rect 10861 1463 10895 1497
rect 10935 1463 10969 1497
rect 11009 1463 11043 1497
rect 11083 1463 11117 1497
rect 11157 1463 11191 1497
rect 11231 1463 11265 1497
rect 11379 1463 11413 1497
rect 11453 1463 11487 1497
rect 11527 1463 11561 1497
rect 11601 1463 11635 1497
rect 11675 1463 11709 1497
rect 11749 1463 11783 1497
rect 11823 1463 11857 1497
rect 11897 1463 11931 1497
rect 11971 1463 12005 1497
rect 12045 1463 12079 1497
rect 12119 1463 12153 1497
rect 12193 1463 12227 1497
rect 12341 1463 12375 1497
rect 12415 1463 12449 1497
rect 12489 1463 12523 1497
rect 12563 1463 12597 1497
rect 12637 1463 12671 1497
rect 12711 1463 12745 1497
rect 12785 1463 12819 1497
rect 12859 1463 12893 1497
rect 13007 1463 13041 1497
rect 13081 1463 13115 1497
rect 13155 1463 13189 1497
rect 13229 1463 13263 1497
rect 13303 1463 13337 1497
rect 13377 1463 13411 1497
rect 13451 1463 13485 1497
rect 13525 1463 13559 1497
rect 13599 1463 13633 1497
rect 13673 1463 13707 1497
rect 13747 1463 13781 1497
rect 13821 1463 13855 1497
rect 13969 1463 14003 1497
rect 14043 1463 14077 1497
rect 14117 1463 14151 1497
rect 14191 1463 14225 1497
rect 14265 1463 14299 1497
rect 14339 1463 14373 1497
rect 14413 1463 14447 1497
rect 14487 1463 14521 1497
rect 14561 1463 14595 1497
rect 14635 1463 14669 1497
rect 14709 1463 14743 1497
rect 14783 1463 14817 1497
rect 14931 1463 14965 1497
rect 15005 1463 15039 1497
rect 15079 1463 15113 1497
rect 15153 1463 15187 1497
rect 15227 1463 15261 1497
rect 15301 1463 15335 1497
rect 15375 1463 15409 1497
rect 15449 1463 15483 1497
rect 15597 1463 15631 1497
rect 15671 1463 15705 1497
rect 15745 1463 15779 1497
rect 15819 1463 15853 1497
rect 15893 1463 15927 1497
rect 15967 1463 16001 1497
rect 16041 1463 16075 1497
rect 16115 1463 16149 1497
rect 16263 1463 16297 1497
rect 16337 1463 16371 1497
rect 16411 1463 16445 1497
rect 16485 1463 16519 1497
rect 16559 1463 16593 1497
rect 16633 1463 16667 1497
rect 16707 1463 16741 1497
rect 16781 1463 16815 1497
rect 16929 1463 16963 1497
rect 17003 1463 17037 1497
rect 17077 1463 17111 1497
rect 17151 1463 17185 1497
rect 17225 1463 17259 1497
rect 17299 1463 17333 1497
rect 17373 1463 17407 1497
rect 17447 1463 17481 1497
rect 17595 1463 17629 1497
rect 17669 1463 17703 1497
rect 17743 1463 17777 1497
rect 17817 1463 17851 1497
rect 17891 1463 17925 1497
rect 205 797 239 831
rect 427 871 461 905
rect 649 649 683 683
rect 797 723 831 757
rect 1167 723 1201 757
rect 1389 501 1423 535
rect 1611 433 1645 461
rect 1611 427 1645 433
rect 1759 649 1793 683
rect 2129 649 2163 683
rect 2277 797 2311 831
rect 2425 649 2459 683
rect 2795 649 2829 683
rect 3017 871 3051 905
rect 3239 433 3273 461
rect 3239 427 3273 433
rect 3387 797 3421 831
rect 3757 723 3791 757
rect 3979 433 4013 461
rect 3979 427 4013 433
rect 4201 575 4235 609
rect 4349 797 4383 831
rect 4719 797 4753 831
rect 4867 797 4901 831
rect 5015 575 5049 609
rect 5385 797 5419 831
rect 5607 871 5641 905
rect 5829 649 5863 683
rect 5977 723 6011 757
rect 6347 723 6381 757
rect 6569 501 6603 535
rect 6791 433 6825 461
rect 6791 427 6825 433
rect 6939 649 6973 683
rect 7309 649 7343 683
rect 7457 797 7491 831
rect 7605 649 7639 683
rect 7975 649 8009 683
rect 8197 871 8231 905
rect 8419 433 8453 461
rect 8419 427 8453 433
rect 8567 797 8601 831
rect 8937 723 8971 757
rect 9159 433 9193 461
rect 9159 427 9193 433
rect 9381 649 9415 683
rect 9529 723 9563 757
rect 9899 723 9933 757
rect 10047 797 10081 831
rect 10195 649 10229 683
rect 10565 797 10599 831
rect 10787 871 10821 905
rect 11009 649 11043 683
rect 11157 723 11191 757
rect 11527 723 11561 757
rect 11749 501 11783 535
rect 11971 433 12005 461
rect 11971 427 12005 433
rect 12119 649 12153 683
rect 12489 649 12523 683
rect 12637 797 12671 831
rect 12785 649 12819 683
rect 13155 649 13189 683
rect 13377 871 13411 905
rect 13599 433 13633 461
rect 13599 427 13633 433
rect 13747 797 13781 831
rect 14117 723 14151 757
rect 14339 433 14373 461
rect 14339 427 14373 433
rect 14561 723 14595 757
rect 14709 797 14743 831
rect 15079 797 15113 831
rect 15227 797 15261 831
rect 15945 1025 15979 1059
rect 16345 1025 16379 1059
rect 16609 1025 16643 1059
rect 15671 871 15705 905
rect 15375 723 15409 757
rect 15671 649 15705 683
rect 17013 1025 17047 1059
rect 15893 797 15927 831
rect 16411 871 16445 905
rect 15893 723 15927 757
rect 16707 575 16741 609
rect 16707 399 16741 433
rect 15953 219 15987 253
rect 17003 399 17037 433
rect 17225 797 17259 831
rect 17373 797 17407 831
rect 16619 219 16653 253
rect 17669 797 17703 831
rect 17285 219 17319 253
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4793 -17 4827 17
rect 4867 -17 4901 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5089 -17 5123 17
rect 5237 -17 5271 17
rect 5311 -17 5345 17
rect 5385 -17 5419 17
rect 5459 -17 5493 17
rect 5533 -17 5567 17
rect 5607 -17 5641 17
rect 5681 -17 5715 17
rect 5755 -17 5789 17
rect 5829 -17 5863 17
rect 5903 -17 5937 17
rect 5977 -17 6011 17
rect 6051 -17 6085 17
rect 6199 -17 6233 17
rect 6273 -17 6307 17
rect 6347 -17 6381 17
rect 6421 -17 6455 17
rect 6495 -17 6529 17
rect 6569 -17 6603 17
rect 6643 -17 6677 17
rect 6717 -17 6751 17
rect 6791 -17 6825 17
rect 6865 -17 6899 17
rect 6939 -17 6973 17
rect 7013 -17 7047 17
rect 7161 -17 7195 17
rect 7235 -17 7269 17
rect 7309 -17 7343 17
rect 7383 -17 7417 17
rect 7457 -17 7491 17
rect 7531 -17 7565 17
rect 7605 -17 7639 17
rect 7679 -17 7713 17
rect 7827 -17 7861 17
rect 7901 -17 7935 17
rect 7975 -17 8009 17
rect 8049 -17 8083 17
rect 8123 -17 8157 17
rect 8197 -17 8231 17
rect 8271 -17 8305 17
rect 8345 -17 8379 17
rect 8419 -17 8453 17
rect 8493 -17 8527 17
rect 8567 -17 8601 17
rect 8641 -17 8675 17
rect 8789 -17 8823 17
rect 8863 -17 8897 17
rect 8937 -17 8971 17
rect 9011 -17 9045 17
rect 9085 -17 9119 17
rect 9159 -17 9193 17
rect 9233 -17 9267 17
rect 9307 -17 9341 17
rect 9381 -17 9415 17
rect 9455 -17 9489 17
rect 9529 -17 9563 17
rect 9603 -17 9637 17
rect 9751 -17 9785 17
rect 9825 -17 9859 17
rect 9899 -17 9933 17
rect 9973 -17 10007 17
rect 10047 -17 10081 17
rect 10121 -17 10155 17
rect 10195 -17 10229 17
rect 10269 -17 10303 17
rect 10417 -17 10451 17
rect 10491 -17 10525 17
rect 10565 -17 10599 17
rect 10639 -17 10673 17
rect 10713 -17 10747 17
rect 10787 -17 10821 17
rect 10861 -17 10895 17
rect 10935 -17 10969 17
rect 11009 -17 11043 17
rect 11083 -17 11117 17
rect 11157 -17 11191 17
rect 11231 -17 11265 17
rect 11379 -17 11413 17
rect 11453 -17 11487 17
rect 11527 -17 11561 17
rect 11601 -17 11635 17
rect 11675 -17 11709 17
rect 11749 -17 11783 17
rect 11823 -17 11857 17
rect 11897 -17 11931 17
rect 11971 -17 12005 17
rect 12045 -17 12079 17
rect 12119 -17 12153 17
rect 12193 -17 12227 17
rect 12341 -17 12375 17
rect 12415 -17 12449 17
rect 12489 -17 12523 17
rect 12563 -17 12597 17
rect 12637 -17 12671 17
rect 12711 -17 12745 17
rect 12785 -17 12819 17
rect 12859 -17 12893 17
rect 13007 -17 13041 17
rect 13081 -17 13115 17
rect 13155 -17 13189 17
rect 13229 -17 13263 17
rect 13303 -17 13337 17
rect 13377 -17 13411 17
rect 13451 -17 13485 17
rect 13525 -17 13559 17
rect 13599 -17 13633 17
rect 13673 -17 13707 17
rect 13747 -17 13781 17
rect 13821 -17 13855 17
rect 13969 -17 14003 17
rect 14043 -17 14077 17
rect 14117 -17 14151 17
rect 14191 -17 14225 17
rect 14265 -17 14299 17
rect 14339 -17 14373 17
rect 14413 -17 14447 17
rect 14487 -17 14521 17
rect 14561 -17 14595 17
rect 14635 -17 14669 17
rect 14709 -17 14743 17
rect 14783 -17 14817 17
rect 14931 -17 14965 17
rect 15005 -17 15039 17
rect 15079 -17 15113 17
rect 15153 -17 15187 17
rect 15227 -17 15261 17
rect 15301 -17 15335 17
rect 15375 -17 15409 17
rect 15449 -17 15483 17
rect 15597 -17 15631 17
rect 15671 -17 15705 17
rect 15745 -17 15779 17
rect 15819 -17 15853 17
rect 15893 -17 15927 17
rect 15967 -17 16001 17
rect 16041 -17 16075 17
rect 16115 -17 16149 17
rect 16263 -17 16297 17
rect 16337 -17 16371 17
rect 16411 -17 16445 17
rect 16485 -17 16519 17
rect 16559 -17 16593 17
rect 16633 -17 16667 17
rect 16707 -17 16741 17
rect 16781 -17 16815 17
rect 16929 -17 16963 17
rect 17003 -17 17037 17
rect 17077 -17 17111 17
rect 17151 -17 17185 17
rect 17225 -17 17259 17
rect 17299 -17 17333 17
rect 17373 -17 17407 17
rect 17447 -17 17481 17
rect 17595 -17 17629 17
rect 17669 -17 17703 17
rect 17743 -17 17777 17
rect 17817 -17 17851 17
rect 17891 -17 17925 17
<< metal1 >>
rect -34 1497 18016 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4867 1497
rect 4901 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5533 1497
rect 5567 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5755 1497
rect 5789 1463 5829 1497
rect 5863 1463 5903 1497
rect 5937 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6199 1497
rect 6233 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6495 1497
rect 6529 1463 6569 1497
rect 6603 1463 6643 1497
rect 6677 1463 6717 1497
rect 6751 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7161 1497
rect 7195 1463 7235 1497
rect 7269 1463 7309 1497
rect 7343 1463 7383 1497
rect 7417 1463 7457 1497
rect 7491 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7679 1497
rect 7713 1463 7827 1497
rect 7861 1463 7901 1497
rect 7935 1463 7975 1497
rect 8009 1463 8049 1497
rect 8083 1463 8123 1497
rect 8157 1463 8197 1497
rect 8231 1463 8271 1497
rect 8305 1463 8345 1497
rect 8379 1463 8419 1497
rect 8453 1463 8493 1497
rect 8527 1463 8567 1497
rect 8601 1463 8641 1497
rect 8675 1463 8789 1497
rect 8823 1463 8863 1497
rect 8897 1463 8937 1497
rect 8971 1463 9011 1497
rect 9045 1463 9085 1497
rect 9119 1463 9159 1497
rect 9193 1463 9233 1497
rect 9267 1463 9307 1497
rect 9341 1463 9381 1497
rect 9415 1463 9455 1497
rect 9489 1463 9529 1497
rect 9563 1463 9603 1497
rect 9637 1463 9751 1497
rect 9785 1463 9825 1497
rect 9859 1463 9899 1497
rect 9933 1463 9973 1497
rect 10007 1463 10047 1497
rect 10081 1463 10121 1497
rect 10155 1463 10195 1497
rect 10229 1463 10269 1497
rect 10303 1463 10417 1497
rect 10451 1463 10491 1497
rect 10525 1463 10565 1497
rect 10599 1463 10639 1497
rect 10673 1463 10713 1497
rect 10747 1463 10787 1497
rect 10821 1463 10861 1497
rect 10895 1463 10935 1497
rect 10969 1463 11009 1497
rect 11043 1463 11083 1497
rect 11117 1463 11157 1497
rect 11191 1463 11231 1497
rect 11265 1463 11379 1497
rect 11413 1463 11453 1497
rect 11487 1463 11527 1497
rect 11561 1463 11601 1497
rect 11635 1463 11675 1497
rect 11709 1463 11749 1497
rect 11783 1463 11823 1497
rect 11857 1463 11897 1497
rect 11931 1463 11971 1497
rect 12005 1463 12045 1497
rect 12079 1463 12119 1497
rect 12153 1463 12193 1497
rect 12227 1463 12341 1497
rect 12375 1463 12415 1497
rect 12449 1463 12489 1497
rect 12523 1463 12563 1497
rect 12597 1463 12637 1497
rect 12671 1463 12711 1497
rect 12745 1463 12785 1497
rect 12819 1463 12859 1497
rect 12893 1463 13007 1497
rect 13041 1463 13081 1497
rect 13115 1463 13155 1497
rect 13189 1463 13229 1497
rect 13263 1463 13303 1497
rect 13337 1463 13377 1497
rect 13411 1463 13451 1497
rect 13485 1463 13525 1497
rect 13559 1463 13599 1497
rect 13633 1463 13673 1497
rect 13707 1463 13747 1497
rect 13781 1463 13821 1497
rect 13855 1463 13969 1497
rect 14003 1463 14043 1497
rect 14077 1463 14117 1497
rect 14151 1463 14191 1497
rect 14225 1463 14265 1497
rect 14299 1463 14339 1497
rect 14373 1463 14413 1497
rect 14447 1463 14487 1497
rect 14521 1463 14561 1497
rect 14595 1463 14635 1497
rect 14669 1463 14709 1497
rect 14743 1463 14783 1497
rect 14817 1463 14931 1497
rect 14965 1463 15005 1497
rect 15039 1463 15079 1497
rect 15113 1463 15153 1497
rect 15187 1463 15227 1497
rect 15261 1463 15301 1497
rect 15335 1463 15375 1497
rect 15409 1463 15449 1497
rect 15483 1463 15597 1497
rect 15631 1463 15671 1497
rect 15705 1463 15745 1497
rect 15779 1463 15819 1497
rect 15853 1463 15893 1497
rect 15927 1463 15967 1497
rect 16001 1463 16041 1497
rect 16075 1463 16115 1497
rect 16149 1463 16263 1497
rect 16297 1463 16337 1497
rect 16371 1463 16411 1497
rect 16445 1463 16485 1497
rect 16519 1463 16559 1497
rect 16593 1463 16633 1497
rect 16667 1463 16707 1497
rect 16741 1463 16781 1497
rect 16815 1463 16929 1497
rect 16963 1463 17003 1497
rect 17037 1463 17077 1497
rect 17111 1463 17151 1497
rect 17185 1463 17225 1497
rect 17259 1463 17299 1497
rect 17333 1463 17373 1497
rect 17407 1463 17447 1497
rect 17481 1463 17595 1497
rect 17629 1463 17669 1497
rect 17703 1463 17743 1497
rect 17777 1463 17817 1497
rect 17851 1463 17891 1497
rect 17925 1463 18016 1497
rect -34 1446 18016 1463
rect 15939 1059 15985 1065
rect 16339 1059 16385 1065
rect 16603 1059 16649 1065
rect 17007 1059 17053 1065
rect 15933 1025 15945 1059
rect 15979 1025 16345 1059
rect 16379 1025 16391 1059
rect 16597 1025 16609 1059
rect 16643 1025 17013 1059
rect 17047 1025 17059 1059
rect 15939 1019 15985 1025
rect 16339 1019 16385 1025
rect 16603 1019 16649 1025
rect 17007 1019 17053 1025
rect 421 905 467 911
rect 3011 905 3057 911
rect 5601 905 5647 911
rect 8191 905 8237 911
rect 10781 905 10827 911
rect 13371 905 13417 911
rect 15665 905 15711 911
rect 16405 905 16451 911
rect 415 871 427 905
rect 461 871 3017 905
rect 3051 871 5607 905
rect 5641 871 8197 905
rect 8231 871 10787 905
rect 10821 871 13377 905
rect 13411 871 13423 905
rect 15659 871 15671 905
rect 15705 871 16411 905
rect 16445 871 16457 905
rect 421 865 467 871
rect 3011 865 3057 871
rect 5601 865 5647 871
rect 8191 865 8237 871
rect 10781 865 10827 871
rect 13371 865 13417 871
rect 15665 865 15711 871
rect 16405 865 16451 871
rect 199 831 245 837
rect 2271 831 2317 837
rect 3381 831 3427 837
rect 4343 831 4389 837
rect 4713 831 4759 837
rect 4861 831 4907 837
rect 5379 831 5425 837
rect 7451 831 7497 837
rect 8561 831 8607 837
rect 10041 831 10087 837
rect 10559 831 10605 837
rect 12631 831 12677 837
rect 13741 831 13787 837
rect 14703 831 14749 837
rect 15073 831 15119 837
rect 15221 831 15267 837
rect 15887 831 15933 837
rect 17219 831 17265 837
rect 17367 831 17413 837
rect 17663 831 17709 837
rect 193 797 205 831
rect 239 797 2277 831
rect 2311 797 3387 831
rect 3421 797 4349 831
rect 4383 797 4719 831
rect 4753 797 4867 831
rect 4901 797 4913 831
rect 5373 797 5385 831
rect 5419 797 7457 831
rect 7491 797 8567 831
rect 8601 797 10047 831
rect 10081 797 10093 831
rect 10553 797 10565 831
rect 10599 797 12637 831
rect 12671 797 13747 831
rect 13781 797 14709 831
rect 14743 797 15079 831
rect 15113 797 15227 831
rect 15261 797 15273 831
rect 15881 797 15893 831
rect 15927 797 17225 831
rect 17259 797 17271 831
rect 17361 797 17373 831
rect 17407 797 17669 831
rect 17703 797 17715 831
rect 199 791 245 797
rect 2271 791 2317 797
rect 3381 791 3427 797
rect 4343 791 4389 797
rect 4713 791 4759 797
rect 4861 791 4907 797
rect 5379 791 5425 797
rect 7451 791 7497 797
rect 8561 791 8607 797
rect 10041 791 10087 797
rect 10559 791 10605 797
rect 12631 791 12677 797
rect 13741 791 13787 797
rect 14703 791 14749 797
rect 15073 791 15119 797
rect 15221 791 15267 797
rect 15887 791 15933 797
rect 17219 791 17265 797
rect 17367 791 17413 797
rect 17663 791 17709 797
rect 791 757 837 763
rect 1161 757 1207 763
rect 3751 757 3797 763
rect 5971 757 6017 763
rect 6341 757 6387 763
rect 8931 757 8977 763
rect 9523 757 9569 763
rect 9893 757 9939 763
rect 11151 757 11197 763
rect 11521 757 11567 763
rect 14111 757 14157 763
rect 14555 757 14601 763
rect 15369 757 15415 763
rect 15887 757 15933 763
rect 785 723 797 757
rect 831 723 1167 757
rect 1201 723 3757 757
rect 3791 723 3803 757
rect 5965 723 5977 757
rect 6011 723 6347 757
rect 6381 723 8937 757
rect 8971 723 8983 757
rect 9517 723 9529 757
rect 9563 723 9899 757
rect 9933 723 9945 757
rect 11145 723 11157 757
rect 11191 723 11527 757
rect 11561 723 14117 757
rect 14151 723 14163 757
rect 14549 723 14561 757
rect 14595 723 15375 757
rect 15409 723 15893 757
rect 15927 723 15939 757
rect 791 717 837 723
rect 1161 717 1207 723
rect 3751 717 3797 723
rect 5971 717 6017 723
rect 6341 717 6387 723
rect 8931 717 8977 723
rect 9523 717 9569 723
rect 9893 717 9939 723
rect 11151 717 11197 723
rect 11521 717 11567 723
rect 14111 717 14157 723
rect 14555 717 14601 723
rect 15369 717 15415 723
rect 15887 717 15933 723
rect 643 683 689 689
rect 1753 683 1799 689
rect 2123 683 2169 689
rect 2419 683 2465 689
rect 2789 683 2835 689
rect 5823 683 5869 689
rect 6933 683 6979 689
rect 7303 683 7349 689
rect 7599 683 7645 689
rect 7969 683 8015 689
rect 9375 683 9421 689
rect 10189 683 10235 689
rect 11003 683 11049 689
rect 12113 683 12159 689
rect 12483 683 12529 689
rect 12779 683 12825 689
rect 13149 683 13195 689
rect 15665 683 15711 689
rect 637 649 649 683
rect 683 649 1759 683
rect 1793 649 2129 683
rect 2163 649 2175 683
rect 2413 649 2425 683
rect 2459 649 2795 683
rect 2829 649 2841 683
rect 5817 649 5829 683
rect 5863 649 6939 683
rect 6973 649 7309 683
rect 7343 649 7355 683
rect 7593 649 7605 683
rect 7639 649 7975 683
rect 8009 649 8021 683
rect 9369 649 9381 683
rect 9415 649 10195 683
rect 10229 649 11009 683
rect 11043 649 12119 683
rect 12153 649 12489 683
rect 12523 649 12785 683
rect 12819 649 13155 683
rect 13189 649 15671 683
rect 15705 649 15717 683
rect 643 643 689 649
rect 1753 643 1799 649
rect 2123 643 2169 649
rect 2419 643 2465 649
rect 2789 643 2835 649
rect 5823 643 5869 649
rect 6933 643 6979 649
rect 7303 643 7349 649
rect 7599 643 7645 649
rect 7969 643 8015 649
rect 9375 643 9421 649
rect 10189 643 10235 649
rect 11003 643 11049 649
rect 12113 643 12159 649
rect 12483 643 12529 649
rect 12779 643 12825 649
rect 13149 643 13195 649
rect 15665 643 15711 649
rect 4195 609 4241 615
rect 5009 609 5055 615
rect 16701 609 16747 615
rect 4189 575 4201 609
rect 4235 575 5015 609
rect 5049 575 16707 609
rect 16741 575 16753 609
rect 4195 569 4241 575
rect 5009 569 5055 575
rect 16701 569 16747 575
rect 1383 535 1429 541
rect 6563 535 6609 541
rect 11743 535 11789 541
rect 1377 501 1389 535
rect 1423 501 6569 535
rect 6603 501 11749 535
rect 11783 501 11819 535
rect 1383 495 1429 501
rect 6563 495 6609 501
rect 11743 495 11789 501
rect 1605 461 1651 467
rect 3233 461 3279 467
rect 3973 461 4019 467
rect 6785 461 6831 467
rect 8413 461 8459 467
rect 9153 461 9199 467
rect 11965 461 12011 467
rect 13593 461 13639 467
rect 14333 461 14379 467
rect 1599 427 1611 461
rect 1645 427 3239 461
rect 3273 427 3979 461
rect 4013 427 6791 461
rect 6825 427 8419 461
rect 8453 427 9159 461
rect 9193 427 11971 461
rect 12005 427 13599 461
rect 13633 427 14339 461
rect 14373 427 14385 461
rect 16701 433 16747 439
rect 16997 433 17043 439
rect 1605 421 1651 427
rect 3233 421 3279 427
rect 3973 421 4019 427
rect 6785 421 6831 427
rect 8413 421 8459 427
rect 9153 421 9199 427
rect 11965 421 12011 427
rect 13593 421 13639 427
rect 14333 421 14379 427
rect 16695 399 16707 433
rect 16741 399 17003 433
rect 17037 399 17049 433
rect 16701 393 16747 399
rect 16997 393 17043 399
rect 15947 253 15993 259
rect 16613 253 16659 259
rect 17279 253 17325 259
rect 15941 219 15953 253
rect 15987 219 16619 253
rect 16653 219 17285 253
rect 17319 219 17331 253
rect 15947 213 15993 219
rect 16613 213 16659 219
rect 17279 213 17325 219
rect -34 17 18016 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4867 17
rect 4901 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5533 17
rect 5567 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5755 17
rect 5789 -17 5829 17
rect 5863 -17 5903 17
rect 5937 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6199 17
rect 6233 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6495 17
rect 6529 -17 6569 17
rect 6603 -17 6643 17
rect 6677 -17 6717 17
rect 6751 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7161 17
rect 7195 -17 7235 17
rect 7269 -17 7309 17
rect 7343 -17 7383 17
rect 7417 -17 7457 17
rect 7491 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7679 17
rect 7713 -17 7827 17
rect 7861 -17 7901 17
rect 7935 -17 7975 17
rect 8009 -17 8049 17
rect 8083 -17 8123 17
rect 8157 -17 8197 17
rect 8231 -17 8271 17
rect 8305 -17 8345 17
rect 8379 -17 8419 17
rect 8453 -17 8493 17
rect 8527 -17 8567 17
rect 8601 -17 8641 17
rect 8675 -17 8789 17
rect 8823 -17 8863 17
rect 8897 -17 8937 17
rect 8971 -17 9011 17
rect 9045 -17 9085 17
rect 9119 -17 9159 17
rect 9193 -17 9233 17
rect 9267 -17 9307 17
rect 9341 -17 9381 17
rect 9415 -17 9455 17
rect 9489 -17 9529 17
rect 9563 -17 9603 17
rect 9637 -17 9751 17
rect 9785 -17 9825 17
rect 9859 -17 9899 17
rect 9933 -17 9973 17
rect 10007 -17 10047 17
rect 10081 -17 10121 17
rect 10155 -17 10195 17
rect 10229 -17 10269 17
rect 10303 -17 10417 17
rect 10451 -17 10491 17
rect 10525 -17 10565 17
rect 10599 -17 10639 17
rect 10673 -17 10713 17
rect 10747 -17 10787 17
rect 10821 -17 10861 17
rect 10895 -17 10935 17
rect 10969 -17 11009 17
rect 11043 -17 11083 17
rect 11117 -17 11157 17
rect 11191 -17 11231 17
rect 11265 -17 11379 17
rect 11413 -17 11453 17
rect 11487 -17 11527 17
rect 11561 -17 11601 17
rect 11635 -17 11675 17
rect 11709 -17 11749 17
rect 11783 -17 11823 17
rect 11857 -17 11897 17
rect 11931 -17 11971 17
rect 12005 -17 12045 17
rect 12079 -17 12119 17
rect 12153 -17 12193 17
rect 12227 -17 12341 17
rect 12375 -17 12415 17
rect 12449 -17 12489 17
rect 12523 -17 12563 17
rect 12597 -17 12637 17
rect 12671 -17 12711 17
rect 12745 -17 12785 17
rect 12819 -17 12859 17
rect 12893 -17 13007 17
rect 13041 -17 13081 17
rect 13115 -17 13155 17
rect 13189 -17 13229 17
rect 13263 -17 13303 17
rect 13337 -17 13377 17
rect 13411 -17 13451 17
rect 13485 -17 13525 17
rect 13559 -17 13599 17
rect 13633 -17 13673 17
rect 13707 -17 13747 17
rect 13781 -17 13821 17
rect 13855 -17 13969 17
rect 14003 -17 14043 17
rect 14077 -17 14117 17
rect 14151 -17 14191 17
rect 14225 -17 14265 17
rect 14299 -17 14339 17
rect 14373 -17 14413 17
rect 14447 -17 14487 17
rect 14521 -17 14561 17
rect 14595 -17 14635 17
rect 14669 -17 14709 17
rect 14743 -17 14783 17
rect 14817 -17 14931 17
rect 14965 -17 15005 17
rect 15039 -17 15079 17
rect 15113 -17 15153 17
rect 15187 -17 15227 17
rect 15261 -17 15301 17
rect 15335 -17 15375 17
rect 15409 -17 15449 17
rect 15483 -17 15597 17
rect 15631 -17 15671 17
rect 15705 -17 15745 17
rect 15779 -17 15819 17
rect 15853 -17 15893 17
rect 15927 -17 15967 17
rect 16001 -17 16041 17
rect 16075 -17 16115 17
rect 16149 -17 16263 17
rect 16297 -17 16337 17
rect 16371 -17 16411 17
rect 16445 -17 16485 17
rect 16519 -17 16559 17
rect 16593 -17 16633 17
rect 16667 -17 16707 17
rect 16741 -17 16781 17
rect 16815 -17 16929 17
rect 16963 -17 17003 17
rect 17037 -17 17077 17
rect 17111 -17 17151 17
rect 17185 -17 17225 17
rect 17259 -17 17299 17
rect 17333 -17 17373 17
rect 17407 -17 17447 17
rect 17481 -17 17595 17
rect 17629 -17 17669 17
rect 17703 -17 17743 17
rect 17777 -17 17817 17
rect 17851 -17 17891 17
rect 17925 -17 18016 17
rect -34 -34 18016 -17
<< labels >>
rlabel metal1 17817 871 17851 905 1 Q
port 1 n
rlabel metal1 17817 797 17851 831 1 Q
port 2 n
rlabel metal1 17817 723 17851 757 1 Q
port 3 n
rlabel metal1 17817 649 17851 683 1 Q
port 4 n
rlabel metal1 17817 575 17851 609 1 Q
port 5 n
rlabel metal1 17817 501 17851 535 1 Q
port 6 n
rlabel metal1 17817 427 17851 461 1 Q
port 7 n
rlabel metal1 1389 501 1423 535 1 D
port 8 n
rlabel metal1 1389 575 1423 609 1 D
port 9 n
rlabel metal1 427 871 461 905 1 CLK
port 10 n
rlabel metal1 427 723 461 757 1 CLK
port 11 n
rlabel metal1 427 649 461 683 1 CLK
port 12 n
rlabel metal1 427 575 461 609 1 CLK
port 13 n
rlabel metal1 427 501 461 535 1 CLK
port 14 n
rlabel metal1 3017 575 3051 609 1 CLK
port 15 n
rlabel metal1 3017 649 3051 683 1 CLK
port 16 n
rlabel metal1 5607 649 5641 683 1 CLK
port 17 n
rlabel metal1 5607 723 5641 757 1 CLK
port 18 n
rlabel metal1 8197 649 8231 683 1 CLK
port 19 n
rlabel metal1 10787 723 10821 757 1 CLK
port 20 n
rlabel metal1 3017 871 3051 905 1 CLK
port 21 n
rlabel metal1 5607 871 5641 905 1 CLK
port 22 n
rlabel metal1 8197 871 8231 905 1 CLK
port 23 n
rlabel metal1 10787 871 10821 905 1 CLK
port 24 n
rlabel metal1 13377 871 13411 905 1 CLK
port 25 n
rlabel metal1 1611 575 1645 609 1 RN
port 26 n
rlabel metal1 1611 427 1645 461 1 RN
port 27 n
rlabel metal1 3239 575 3273 609 1 RN
port 28 n
rlabel metal1 3239 649 3273 683 1 RN
port 29 n
rlabel metal1 3979 649 4013 683 1 RN
port 30 n
rlabel metal1 3979 575 4013 609 1 RN
port 31 n
rlabel metal1 8419 649 8453 683 1 RN
port 32 n
rlabel metal1 9159 649 9193 683 1 RN
port 33 n
rlabel metal1 9159 723 9193 757 1 RN
port 34 n
rlabel metal1 14339 723 14373 757 1 RN
port 35 n
rlabel metal1 -34 1446 18016 1514 1 VPWR
port 36 n
rlabel metal1 -34 -34 18016 34 1 VGND
port 37 n
rlabel nwell 57 1463 91 1497 1 VPB
port 38 n
rlabel pwell 57 -17 91 17 1 VNB
port 39 n
<< end >>
