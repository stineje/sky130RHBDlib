magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< metal3 >>
rect 10151 1378 14931 2306
<< obsm3 >>
rect 120 1378 4900 2306
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 15000 10947
rect 0 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 15000 9869
rect 0 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 2304 254 2307
rect 0 2240 272 2304
rect 290 2240 354 2304
rect 372 2240 436 2304
rect 454 2240 518 2304
rect 536 2240 600 2304
rect 618 2240 682 2304
rect 699 2240 763 2304
rect 780 2240 844 2304
rect 861 2240 925 2304
rect 942 2240 1006 2304
rect 1023 2240 1087 2304
rect 1104 2240 1168 2304
rect 1185 2240 1249 2304
rect 1266 2240 1330 2304
rect 1347 2240 1411 2304
rect 1428 2240 1492 2304
rect 1509 2240 1573 2304
rect 1590 2240 1654 2304
rect 1671 2240 1735 2304
rect 1752 2240 1816 2304
rect 1833 2240 1897 2304
rect 1914 2240 1978 2304
rect 1995 2240 2059 2304
rect 2076 2240 2140 2304
rect 2157 2240 2221 2304
rect 2238 2240 2302 2304
rect 2319 2240 2383 2304
rect 2400 2240 2464 2304
rect 2481 2240 2545 2304
rect 2562 2240 2626 2304
rect 2643 2240 2707 2304
rect 2724 2240 2788 2304
rect 2805 2240 2869 2304
rect 2886 2240 2950 2304
rect 2967 2240 3031 2304
rect 3048 2240 3112 2304
rect 3129 2240 3193 2304
rect 3210 2240 3274 2304
rect 3291 2240 3355 2304
rect 3372 2240 3436 2304
rect 3453 2240 3517 2304
rect 3534 2240 3598 2304
rect 3615 2240 3679 2304
rect 3696 2240 3760 2304
rect 3777 2240 3841 2304
rect 3858 2240 3922 2304
rect 3939 2240 4003 2304
rect 4020 2240 4084 2304
rect 4101 2240 4165 2304
rect 4182 2240 4246 2304
rect 4263 2240 4327 2304
rect 4344 2240 4408 2304
rect 4425 2240 4489 2304
rect 4506 2240 4570 2304
rect 4587 2240 4651 2304
rect 4668 2240 4732 2304
rect 4749 2240 4813 2304
rect 4830 2240 4894 2304
rect 0 2218 254 2240
rect 0 2154 272 2218
rect 290 2154 354 2218
rect 372 2154 436 2218
rect 454 2154 518 2218
rect 536 2154 600 2218
rect 618 2154 682 2218
rect 699 2154 763 2218
rect 780 2154 844 2218
rect 861 2154 925 2218
rect 942 2154 1006 2218
rect 1023 2154 1087 2218
rect 1104 2154 1168 2218
rect 1185 2154 1249 2218
rect 1266 2154 1330 2218
rect 1347 2154 1411 2218
rect 1428 2154 1492 2218
rect 1509 2154 1573 2218
rect 1590 2154 1654 2218
rect 1671 2154 1735 2218
rect 1752 2154 1816 2218
rect 1833 2154 1897 2218
rect 1914 2154 1978 2218
rect 1995 2154 2059 2218
rect 2076 2154 2140 2218
rect 2157 2154 2221 2218
rect 2238 2154 2302 2218
rect 2319 2154 2383 2218
rect 2400 2154 2464 2218
rect 2481 2154 2545 2218
rect 2562 2154 2626 2218
rect 2643 2154 2707 2218
rect 2724 2154 2788 2218
rect 2805 2154 2869 2218
rect 2886 2154 2950 2218
rect 2967 2154 3031 2218
rect 3048 2154 3112 2218
rect 3129 2154 3193 2218
rect 3210 2154 3274 2218
rect 3291 2154 3355 2218
rect 3372 2154 3436 2218
rect 3453 2154 3517 2218
rect 3534 2154 3598 2218
rect 3615 2154 3679 2218
rect 3696 2154 3760 2218
rect 3777 2154 3841 2218
rect 3858 2154 3922 2218
rect 3939 2154 4003 2218
rect 4020 2154 4084 2218
rect 4101 2154 4165 2218
rect 4182 2154 4246 2218
rect 4263 2154 4327 2218
rect 4344 2154 4408 2218
rect 4425 2154 4489 2218
rect 4506 2154 4570 2218
rect 4587 2154 4651 2218
rect 4668 2154 4732 2218
rect 4749 2154 4813 2218
rect 4830 2154 4894 2218
rect 0 2132 254 2154
rect 0 2068 272 2132
rect 290 2068 354 2132
rect 372 2068 436 2132
rect 454 2068 518 2132
rect 536 2068 600 2132
rect 618 2068 682 2132
rect 699 2068 763 2132
rect 780 2068 844 2132
rect 861 2068 925 2132
rect 942 2068 1006 2132
rect 1023 2068 1087 2132
rect 1104 2068 1168 2132
rect 1185 2068 1249 2132
rect 1266 2068 1330 2132
rect 1347 2068 1411 2132
rect 1428 2068 1492 2132
rect 1509 2068 1573 2132
rect 1590 2068 1654 2132
rect 1671 2068 1735 2132
rect 1752 2068 1816 2132
rect 1833 2068 1897 2132
rect 1914 2068 1978 2132
rect 1995 2068 2059 2132
rect 2076 2068 2140 2132
rect 2157 2068 2221 2132
rect 2238 2068 2302 2132
rect 2319 2068 2383 2132
rect 2400 2068 2464 2132
rect 2481 2068 2545 2132
rect 2562 2068 2626 2132
rect 2643 2068 2707 2132
rect 2724 2068 2788 2132
rect 2805 2068 2869 2132
rect 2886 2068 2950 2132
rect 2967 2068 3031 2132
rect 3048 2068 3112 2132
rect 3129 2068 3193 2132
rect 3210 2068 3274 2132
rect 3291 2068 3355 2132
rect 3372 2068 3436 2132
rect 3453 2068 3517 2132
rect 3534 2068 3598 2132
rect 3615 2068 3679 2132
rect 3696 2068 3760 2132
rect 3777 2068 3841 2132
rect 3858 2068 3922 2132
rect 3939 2068 4003 2132
rect 4020 2068 4084 2132
rect 4101 2068 4165 2132
rect 4182 2068 4246 2132
rect 4263 2068 4327 2132
rect 4344 2068 4408 2132
rect 4425 2068 4489 2132
rect 4506 2068 4570 2132
rect 4587 2068 4651 2132
rect 4668 2068 4732 2132
rect 4749 2068 4813 2132
rect 4830 2068 4894 2132
rect 0 2046 254 2068
rect 0 1982 272 2046
rect 290 1982 354 2046
rect 372 1982 436 2046
rect 454 1982 518 2046
rect 536 1982 600 2046
rect 618 1982 682 2046
rect 699 1982 763 2046
rect 780 1982 844 2046
rect 861 1982 925 2046
rect 942 1982 1006 2046
rect 1023 1982 1087 2046
rect 1104 1982 1168 2046
rect 1185 1982 1249 2046
rect 1266 1982 1330 2046
rect 1347 1982 1411 2046
rect 1428 1982 1492 2046
rect 1509 1982 1573 2046
rect 1590 1982 1654 2046
rect 1671 1982 1735 2046
rect 1752 1982 1816 2046
rect 1833 1982 1897 2046
rect 1914 1982 1978 2046
rect 1995 1982 2059 2046
rect 2076 1982 2140 2046
rect 2157 1982 2221 2046
rect 2238 1982 2302 2046
rect 2319 1982 2383 2046
rect 2400 1982 2464 2046
rect 2481 1982 2545 2046
rect 2562 1982 2626 2046
rect 2643 1982 2707 2046
rect 2724 1982 2788 2046
rect 2805 1982 2869 2046
rect 2886 1982 2950 2046
rect 2967 1982 3031 2046
rect 3048 1982 3112 2046
rect 3129 1982 3193 2046
rect 3210 1982 3274 2046
rect 3291 1982 3355 2046
rect 3372 1982 3436 2046
rect 3453 1982 3517 2046
rect 3534 1982 3598 2046
rect 3615 1982 3679 2046
rect 3696 1982 3760 2046
rect 3777 1982 3841 2046
rect 3858 1982 3922 2046
rect 3939 1982 4003 2046
rect 4020 1982 4084 2046
rect 4101 1982 4165 2046
rect 4182 1982 4246 2046
rect 4263 1982 4327 2046
rect 4344 1982 4408 2046
rect 4425 1982 4489 2046
rect 4506 1982 4570 2046
rect 4587 1982 4651 2046
rect 4668 1982 4732 2046
rect 4749 1982 4813 2046
rect 4830 1982 4894 2046
rect 0 1960 254 1982
rect 0 1896 272 1960
rect 290 1896 354 1960
rect 372 1896 436 1960
rect 454 1896 518 1960
rect 536 1896 600 1960
rect 618 1896 682 1960
rect 699 1896 763 1960
rect 780 1896 844 1960
rect 861 1896 925 1960
rect 942 1896 1006 1960
rect 1023 1896 1087 1960
rect 1104 1896 1168 1960
rect 1185 1896 1249 1960
rect 1266 1896 1330 1960
rect 1347 1896 1411 1960
rect 1428 1896 1492 1960
rect 1509 1896 1573 1960
rect 1590 1896 1654 1960
rect 1671 1896 1735 1960
rect 1752 1896 1816 1960
rect 1833 1896 1897 1960
rect 1914 1896 1978 1960
rect 1995 1896 2059 1960
rect 2076 1896 2140 1960
rect 2157 1896 2221 1960
rect 2238 1896 2302 1960
rect 2319 1896 2383 1960
rect 2400 1896 2464 1960
rect 2481 1896 2545 1960
rect 2562 1896 2626 1960
rect 2643 1896 2707 1960
rect 2724 1896 2788 1960
rect 2805 1896 2869 1960
rect 2886 1896 2950 1960
rect 2967 1896 3031 1960
rect 3048 1896 3112 1960
rect 3129 1896 3193 1960
rect 3210 1896 3274 1960
rect 3291 1896 3355 1960
rect 3372 1896 3436 1960
rect 3453 1896 3517 1960
rect 3534 1896 3598 1960
rect 3615 1896 3679 1960
rect 3696 1896 3760 1960
rect 3777 1896 3841 1960
rect 3858 1896 3922 1960
rect 3939 1896 4003 1960
rect 4020 1896 4084 1960
rect 4101 1896 4165 1960
rect 4182 1896 4246 1960
rect 4263 1896 4327 1960
rect 4344 1896 4408 1960
rect 4425 1896 4489 1960
rect 4506 1896 4570 1960
rect 4587 1896 4651 1960
rect 4668 1896 4732 1960
rect 4749 1896 4813 1960
rect 4830 1896 4894 1960
rect 0 1874 254 1896
rect 0 1810 272 1874
rect 290 1810 354 1874
rect 372 1810 436 1874
rect 454 1810 518 1874
rect 536 1810 600 1874
rect 618 1810 682 1874
rect 699 1810 763 1874
rect 780 1810 844 1874
rect 861 1810 925 1874
rect 942 1810 1006 1874
rect 1023 1810 1087 1874
rect 1104 1810 1168 1874
rect 1185 1810 1249 1874
rect 1266 1810 1330 1874
rect 1347 1810 1411 1874
rect 1428 1810 1492 1874
rect 1509 1810 1573 1874
rect 1590 1810 1654 1874
rect 1671 1810 1735 1874
rect 1752 1810 1816 1874
rect 1833 1810 1897 1874
rect 1914 1810 1978 1874
rect 1995 1810 2059 1874
rect 2076 1810 2140 1874
rect 2157 1810 2221 1874
rect 2238 1810 2302 1874
rect 2319 1810 2383 1874
rect 2400 1810 2464 1874
rect 2481 1810 2545 1874
rect 2562 1810 2626 1874
rect 2643 1810 2707 1874
rect 2724 1810 2788 1874
rect 2805 1810 2869 1874
rect 2886 1810 2950 1874
rect 2967 1810 3031 1874
rect 3048 1810 3112 1874
rect 3129 1810 3193 1874
rect 3210 1810 3274 1874
rect 3291 1810 3355 1874
rect 3372 1810 3436 1874
rect 3453 1810 3517 1874
rect 3534 1810 3598 1874
rect 3615 1810 3679 1874
rect 3696 1810 3760 1874
rect 3777 1810 3841 1874
rect 3858 1810 3922 1874
rect 3939 1810 4003 1874
rect 4020 1810 4084 1874
rect 4101 1810 4165 1874
rect 4182 1810 4246 1874
rect 4263 1810 4327 1874
rect 4344 1810 4408 1874
rect 4425 1810 4489 1874
rect 4506 1810 4570 1874
rect 4587 1810 4651 1874
rect 4668 1810 4732 1874
rect 4749 1810 4813 1874
rect 4830 1810 4894 1874
rect 0 1788 254 1810
rect 0 1724 272 1788
rect 290 1724 354 1788
rect 372 1724 436 1788
rect 454 1724 518 1788
rect 536 1724 600 1788
rect 618 1724 682 1788
rect 699 1724 763 1788
rect 780 1724 844 1788
rect 861 1724 925 1788
rect 942 1724 1006 1788
rect 1023 1724 1087 1788
rect 1104 1724 1168 1788
rect 1185 1724 1249 1788
rect 1266 1724 1330 1788
rect 1347 1724 1411 1788
rect 1428 1724 1492 1788
rect 1509 1724 1573 1788
rect 1590 1724 1654 1788
rect 1671 1724 1735 1788
rect 1752 1724 1816 1788
rect 1833 1724 1897 1788
rect 1914 1724 1978 1788
rect 1995 1724 2059 1788
rect 2076 1724 2140 1788
rect 2157 1724 2221 1788
rect 2238 1724 2302 1788
rect 2319 1724 2383 1788
rect 2400 1724 2464 1788
rect 2481 1724 2545 1788
rect 2562 1724 2626 1788
rect 2643 1724 2707 1788
rect 2724 1724 2788 1788
rect 2805 1724 2869 1788
rect 2886 1724 2950 1788
rect 2967 1724 3031 1788
rect 3048 1724 3112 1788
rect 3129 1724 3193 1788
rect 3210 1724 3274 1788
rect 3291 1724 3355 1788
rect 3372 1724 3436 1788
rect 3453 1724 3517 1788
rect 3534 1724 3598 1788
rect 3615 1724 3679 1788
rect 3696 1724 3760 1788
rect 3777 1724 3841 1788
rect 3858 1724 3922 1788
rect 3939 1724 4003 1788
rect 4020 1724 4084 1788
rect 4101 1724 4165 1788
rect 4182 1724 4246 1788
rect 4263 1724 4327 1788
rect 4344 1724 4408 1788
rect 4425 1724 4489 1788
rect 4506 1724 4570 1788
rect 4587 1724 4651 1788
rect 4668 1724 4732 1788
rect 4749 1724 4813 1788
rect 4830 1724 4894 1788
rect 0 1702 254 1724
rect 0 1638 272 1702
rect 290 1638 354 1702
rect 372 1638 436 1702
rect 454 1638 518 1702
rect 536 1638 600 1702
rect 618 1638 682 1702
rect 699 1638 763 1702
rect 780 1638 844 1702
rect 861 1638 925 1702
rect 942 1638 1006 1702
rect 1023 1638 1087 1702
rect 1104 1638 1168 1702
rect 1185 1638 1249 1702
rect 1266 1638 1330 1702
rect 1347 1638 1411 1702
rect 1428 1638 1492 1702
rect 1509 1638 1573 1702
rect 1590 1638 1654 1702
rect 1671 1638 1735 1702
rect 1752 1638 1816 1702
rect 1833 1638 1897 1702
rect 1914 1638 1978 1702
rect 1995 1638 2059 1702
rect 2076 1638 2140 1702
rect 2157 1638 2221 1702
rect 2238 1638 2302 1702
rect 2319 1638 2383 1702
rect 2400 1638 2464 1702
rect 2481 1638 2545 1702
rect 2562 1638 2626 1702
rect 2643 1638 2707 1702
rect 2724 1638 2788 1702
rect 2805 1638 2869 1702
rect 2886 1638 2950 1702
rect 2967 1638 3031 1702
rect 3048 1638 3112 1702
rect 3129 1638 3193 1702
rect 3210 1638 3274 1702
rect 3291 1638 3355 1702
rect 3372 1638 3436 1702
rect 3453 1638 3517 1702
rect 3534 1638 3598 1702
rect 3615 1638 3679 1702
rect 3696 1638 3760 1702
rect 3777 1638 3841 1702
rect 3858 1638 3922 1702
rect 3939 1638 4003 1702
rect 4020 1638 4084 1702
rect 4101 1638 4165 1702
rect 4182 1638 4246 1702
rect 4263 1638 4327 1702
rect 4344 1638 4408 1702
rect 4425 1638 4489 1702
rect 4506 1638 4570 1702
rect 4587 1638 4651 1702
rect 4668 1638 4732 1702
rect 4749 1638 4813 1702
rect 4830 1638 4894 1702
rect 0 1616 254 1638
rect 0 1552 272 1616
rect 290 1552 354 1616
rect 372 1552 436 1616
rect 454 1552 518 1616
rect 536 1552 600 1616
rect 618 1552 682 1616
rect 699 1552 763 1616
rect 780 1552 844 1616
rect 861 1552 925 1616
rect 942 1552 1006 1616
rect 1023 1552 1087 1616
rect 1104 1552 1168 1616
rect 1185 1552 1249 1616
rect 1266 1552 1330 1616
rect 1347 1552 1411 1616
rect 1428 1552 1492 1616
rect 1509 1552 1573 1616
rect 1590 1552 1654 1616
rect 1671 1552 1735 1616
rect 1752 1552 1816 1616
rect 1833 1552 1897 1616
rect 1914 1552 1978 1616
rect 1995 1552 2059 1616
rect 2076 1552 2140 1616
rect 2157 1552 2221 1616
rect 2238 1552 2302 1616
rect 2319 1552 2383 1616
rect 2400 1552 2464 1616
rect 2481 1552 2545 1616
rect 2562 1552 2626 1616
rect 2643 1552 2707 1616
rect 2724 1552 2788 1616
rect 2805 1552 2869 1616
rect 2886 1552 2950 1616
rect 2967 1552 3031 1616
rect 3048 1552 3112 1616
rect 3129 1552 3193 1616
rect 3210 1552 3274 1616
rect 3291 1552 3355 1616
rect 3372 1552 3436 1616
rect 3453 1552 3517 1616
rect 3534 1552 3598 1616
rect 3615 1552 3679 1616
rect 3696 1552 3760 1616
rect 3777 1552 3841 1616
rect 3858 1552 3922 1616
rect 3939 1552 4003 1616
rect 4020 1552 4084 1616
rect 4101 1552 4165 1616
rect 4182 1552 4246 1616
rect 4263 1552 4327 1616
rect 4344 1552 4408 1616
rect 4425 1552 4489 1616
rect 4506 1552 4570 1616
rect 4587 1552 4651 1616
rect 4668 1552 4732 1616
rect 4749 1552 4813 1616
rect 4830 1552 4894 1616
rect 0 1530 254 1552
rect 0 1466 272 1530
rect 290 1466 354 1530
rect 372 1466 436 1530
rect 454 1466 518 1530
rect 536 1466 600 1530
rect 618 1466 682 1530
rect 699 1466 763 1530
rect 780 1466 844 1530
rect 861 1466 925 1530
rect 942 1466 1006 1530
rect 1023 1466 1087 1530
rect 1104 1466 1168 1530
rect 1185 1466 1249 1530
rect 1266 1466 1330 1530
rect 1347 1466 1411 1530
rect 1428 1466 1492 1530
rect 1509 1466 1573 1530
rect 1590 1466 1654 1530
rect 1671 1466 1735 1530
rect 1752 1466 1816 1530
rect 1833 1466 1897 1530
rect 1914 1466 1978 1530
rect 1995 1466 2059 1530
rect 2076 1466 2140 1530
rect 2157 1466 2221 1530
rect 2238 1466 2302 1530
rect 2319 1466 2383 1530
rect 2400 1466 2464 1530
rect 2481 1466 2545 1530
rect 2562 1466 2626 1530
rect 2643 1466 2707 1530
rect 2724 1466 2788 1530
rect 2805 1466 2869 1530
rect 2886 1466 2950 1530
rect 2967 1466 3031 1530
rect 3048 1466 3112 1530
rect 3129 1466 3193 1530
rect 3210 1466 3274 1530
rect 3291 1466 3355 1530
rect 3372 1466 3436 1530
rect 3453 1466 3517 1530
rect 3534 1466 3598 1530
rect 3615 1466 3679 1530
rect 3696 1466 3760 1530
rect 3777 1466 3841 1530
rect 3858 1466 3922 1530
rect 3939 1466 4003 1530
rect 4020 1466 4084 1530
rect 4101 1466 4165 1530
rect 4182 1466 4246 1530
rect 4263 1466 4327 1530
rect 4344 1466 4408 1530
rect 4425 1466 4489 1530
rect 4506 1466 4570 1530
rect 4587 1466 4651 1530
rect 4668 1466 4732 1530
rect 4749 1466 4813 1530
rect 4830 1466 4894 1530
rect 0 1444 254 1466
rect 0 1380 272 1444
rect 290 1380 354 1444
rect 372 1380 436 1444
rect 454 1380 518 1444
rect 536 1380 600 1444
rect 618 1380 682 1444
rect 699 1380 763 1444
rect 780 1380 844 1444
rect 861 1380 925 1444
rect 942 1380 1006 1444
rect 1023 1380 1087 1444
rect 1104 1380 1168 1444
rect 1185 1380 1249 1444
rect 1266 1380 1330 1444
rect 1347 1380 1411 1444
rect 1428 1380 1492 1444
rect 1509 1380 1573 1444
rect 1590 1380 1654 1444
rect 1671 1380 1735 1444
rect 1752 1380 1816 1444
rect 1833 1380 1897 1444
rect 1914 1380 1978 1444
rect 1995 1380 2059 1444
rect 2076 1380 2140 1444
rect 2157 1380 2221 1444
rect 2238 1380 2302 1444
rect 2319 1380 2383 1444
rect 2400 1380 2464 1444
rect 2481 1380 2545 1444
rect 2562 1380 2626 1444
rect 2643 1380 2707 1444
rect 2724 1380 2788 1444
rect 2805 1380 2869 1444
rect 2886 1380 2950 1444
rect 2967 1380 3031 1444
rect 3048 1380 3112 1444
rect 3129 1380 3193 1444
rect 3210 1380 3274 1444
rect 3291 1380 3355 1444
rect 3372 1380 3436 1444
rect 3453 1380 3517 1444
rect 3534 1380 3598 1444
rect 3615 1380 3679 1444
rect 3696 1380 3760 1444
rect 3777 1380 3841 1444
rect 3858 1380 3922 1444
rect 3939 1380 4003 1444
rect 4020 1380 4084 1444
rect 4101 1380 4165 1444
rect 4182 1380 4246 1444
rect 4263 1380 4327 1444
rect 4344 1380 4408 1444
rect 4425 1380 4489 1444
rect 4506 1380 4570 1444
rect 4587 1380 4651 1444
rect 4668 1380 4732 1444
rect 4749 1380 4813 1444
rect 4830 1380 4894 1444
rect 0 1377 254 1380
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< obsm4 >>
rect 334 34677 14666 39600
rect 193 18680 14807 34677
rect 334 13527 14666 18680
rect 193 13387 14807 13527
rect 334 12337 14666 13387
rect 193 12217 14807 12337
rect 334 11167 14666 12217
rect 193 11027 14807 11167
rect 334 9949 14666 10145
rect 193 8927 14807 9067
rect 334 7837 14666 8927
rect 193 7717 14807 7837
rect 334 6867 14666 7717
rect 193 6747 14807 6867
rect 334 5897 14666 6747
rect 193 5777 14807 5897
rect 334 4687 14666 5777
rect 193 4567 14807 4687
rect 334 3477 14666 4567
rect 193 3357 14807 3477
rect 273 2507 14727 3357
rect 193 2387 14807 2507
rect 334 2304 14666 2387
rect 354 2240 372 2304
rect 436 2240 454 2304
rect 518 2240 536 2304
rect 600 2240 618 2304
rect 682 2240 699 2304
rect 763 2240 780 2304
rect 844 2240 861 2304
rect 925 2240 942 2304
rect 1006 2240 1023 2304
rect 1087 2240 1104 2304
rect 1168 2240 1185 2304
rect 1249 2240 1266 2304
rect 1330 2240 1347 2304
rect 1411 2240 1428 2304
rect 1492 2240 1509 2304
rect 1573 2240 1590 2304
rect 1654 2240 1671 2304
rect 1735 2240 1752 2304
rect 1816 2240 1833 2304
rect 1897 2240 1914 2304
rect 1978 2240 1995 2304
rect 2059 2240 2076 2304
rect 2140 2240 2157 2304
rect 2221 2240 2238 2304
rect 2302 2240 2319 2304
rect 2383 2240 2400 2304
rect 2464 2240 2481 2304
rect 2545 2240 2562 2304
rect 2626 2240 2643 2304
rect 2707 2240 2724 2304
rect 2788 2240 2805 2304
rect 2869 2240 2886 2304
rect 2950 2240 2967 2304
rect 3031 2240 3048 2304
rect 3112 2240 3129 2304
rect 3193 2240 3210 2304
rect 3274 2240 3291 2304
rect 3355 2240 3372 2304
rect 3436 2240 3453 2304
rect 3517 2240 3534 2304
rect 3598 2240 3615 2304
rect 3679 2240 3696 2304
rect 3760 2240 3777 2304
rect 3841 2240 3858 2304
rect 3922 2240 3939 2304
rect 4003 2240 4020 2304
rect 4084 2240 4101 2304
rect 4165 2240 4182 2304
rect 4246 2240 4263 2304
rect 4327 2240 4344 2304
rect 4408 2240 4425 2304
rect 4489 2240 4506 2304
rect 4570 2240 4587 2304
rect 4651 2240 4668 2304
rect 4732 2240 4749 2304
rect 4813 2240 4830 2304
rect 4894 2240 14666 2304
rect 334 2218 14666 2240
rect 354 2154 372 2218
rect 436 2154 454 2218
rect 518 2154 536 2218
rect 600 2154 618 2218
rect 682 2154 699 2218
rect 763 2154 780 2218
rect 844 2154 861 2218
rect 925 2154 942 2218
rect 1006 2154 1023 2218
rect 1087 2154 1104 2218
rect 1168 2154 1185 2218
rect 1249 2154 1266 2218
rect 1330 2154 1347 2218
rect 1411 2154 1428 2218
rect 1492 2154 1509 2218
rect 1573 2154 1590 2218
rect 1654 2154 1671 2218
rect 1735 2154 1752 2218
rect 1816 2154 1833 2218
rect 1897 2154 1914 2218
rect 1978 2154 1995 2218
rect 2059 2154 2076 2218
rect 2140 2154 2157 2218
rect 2221 2154 2238 2218
rect 2302 2154 2319 2218
rect 2383 2154 2400 2218
rect 2464 2154 2481 2218
rect 2545 2154 2562 2218
rect 2626 2154 2643 2218
rect 2707 2154 2724 2218
rect 2788 2154 2805 2218
rect 2869 2154 2886 2218
rect 2950 2154 2967 2218
rect 3031 2154 3048 2218
rect 3112 2154 3129 2218
rect 3193 2154 3210 2218
rect 3274 2154 3291 2218
rect 3355 2154 3372 2218
rect 3436 2154 3453 2218
rect 3517 2154 3534 2218
rect 3598 2154 3615 2218
rect 3679 2154 3696 2218
rect 3760 2154 3777 2218
rect 3841 2154 3858 2218
rect 3922 2154 3939 2218
rect 4003 2154 4020 2218
rect 4084 2154 4101 2218
rect 4165 2154 4182 2218
rect 4246 2154 4263 2218
rect 4327 2154 4344 2218
rect 4408 2154 4425 2218
rect 4489 2154 4506 2218
rect 4570 2154 4587 2218
rect 4651 2154 4668 2218
rect 4732 2154 4749 2218
rect 4813 2154 4830 2218
rect 4894 2154 14666 2218
rect 334 2132 14666 2154
rect 354 2068 372 2132
rect 436 2068 454 2132
rect 518 2068 536 2132
rect 600 2068 618 2132
rect 682 2068 699 2132
rect 763 2068 780 2132
rect 844 2068 861 2132
rect 925 2068 942 2132
rect 1006 2068 1023 2132
rect 1087 2068 1104 2132
rect 1168 2068 1185 2132
rect 1249 2068 1266 2132
rect 1330 2068 1347 2132
rect 1411 2068 1428 2132
rect 1492 2068 1509 2132
rect 1573 2068 1590 2132
rect 1654 2068 1671 2132
rect 1735 2068 1752 2132
rect 1816 2068 1833 2132
rect 1897 2068 1914 2132
rect 1978 2068 1995 2132
rect 2059 2068 2076 2132
rect 2140 2068 2157 2132
rect 2221 2068 2238 2132
rect 2302 2068 2319 2132
rect 2383 2068 2400 2132
rect 2464 2068 2481 2132
rect 2545 2068 2562 2132
rect 2626 2068 2643 2132
rect 2707 2068 2724 2132
rect 2788 2068 2805 2132
rect 2869 2068 2886 2132
rect 2950 2068 2967 2132
rect 3031 2068 3048 2132
rect 3112 2068 3129 2132
rect 3193 2068 3210 2132
rect 3274 2068 3291 2132
rect 3355 2068 3372 2132
rect 3436 2068 3453 2132
rect 3517 2068 3534 2132
rect 3598 2068 3615 2132
rect 3679 2068 3696 2132
rect 3760 2068 3777 2132
rect 3841 2068 3858 2132
rect 3922 2068 3939 2132
rect 4003 2068 4020 2132
rect 4084 2068 4101 2132
rect 4165 2068 4182 2132
rect 4246 2068 4263 2132
rect 4327 2068 4344 2132
rect 4408 2068 4425 2132
rect 4489 2068 4506 2132
rect 4570 2068 4587 2132
rect 4651 2068 4668 2132
rect 4732 2068 4749 2132
rect 4813 2068 4830 2132
rect 4894 2068 14666 2132
rect 334 2046 14666 2068
rect 354 1982 372 2046
rect 436 1982 454 2046
rect 518 1982 536 2046
rect 600 1982 618 2046
rect 682 1982 699 2046
rect 763 1982 780 2046
rect 844 1982 861 2046
rect 925 1982 942 2046
rect 1006 1982 1023 2046
rect 1087 1982 1104 2046
rect 1168 1982 1185 2046
rect 1249 1982 1266 2046
rect 1330 1982 1347 2046
rect 1411 1982 1428 2046
rect 1492 1982 1509 2046
rect 1573 1982 1590 2046
rect 1654 1982 1671 2046
rect 1735 1982 1752 2046
rect 1816 1982 1833 2046
rect 1897 1982 1914 2046
rect 1978 1982 1995 2046
rect 2059 1982 2076 2046
rect 2140 1982 2157 2046
rect 2221 1982 2238 2046
rect 2302 1982 2319 2046
rect 2383 1982 2400 2046
rect 2464 1982 2481 2046
rect 2545 1982 2562 2046
rect 2626 1982 2643 2046
rect 2707 1982 2724 2046
rect 2788 1982 2805 2046
rect 2869 1982 2886 2046
rect 2950 1982 2967 2046
rect 3031 1982 3048 2046
rect 3112 1982 3129 2046
rect 3193 1982 3210 2046
rect 3274 1982 3291 2046
rect 3355 1982 3372 2046
rect 3436 1982 3453 2046
rect 3517 1982 3534 2046
rect 3598 1982 3615 2046
rect 3679 1982 3696 2046
rect 3760 1982 3777 2046
rect 3841 1982 3858 2046
rect 3922 1982 3939 2046
rect 4003 1982 4020 2046
rect 4084 1982 4101 2046
rect 4165 1982 4182 2046
rect 4246 1982 4263 2046
rect 4327 1982 4344 2046
rect 4408 1982 4425 2046
rect 4489 1982 4506 2046
rect 4570 1982 4587 2046
rect 4651 1982 4668 2046
rect 4732 1982 4749 2046
rect 4813 1982 4830 2046
rect 4894 1982 14666 2046
rect 334 1960 14666 1982
rect 354 1896 372 1960
rect 436 1896 454 1960
rect 518 1896 536 1960
rect 600 1896 618 1960
rect 682 1896 699 1960
rect 763 1896 780 1960
rect 844 1896 861 1960
rect 925 1896 942 1960
rect 1006 1896 1023 1960
rect 1087 1896 1104 1960
rect 1168 1896 1185 1960
rect 1249 1896 1266 1960
rect 1330 1896 1347 1960
rect 1411 1896 1428 1960
rect 1492 1896 1509 1960
rect 1573 1896 1590 1960
rect 1654 1896 1671 1960
rect 1735 1896 1752 1960
rect 1816 1896 1833 1960
rect 1897 1896 1914 1960
rect 1978 1896 1995 1960
rect 2059 1896 2076 1960
rect 2140 1896 2157 1960
rect 2221 1896 2238 1960
rect 2302 1896 2319 1960
rect 2383 1896 2400 1960
rect 2464 1896 2481 1960
rect 2545 1896 2562 1960
rect 2626 1896 2643 1960
rect 2707 1896 2724 1960
rect 2788 1896 2805 1960
rect 2869 1896 2886 1960
rect 2950 1896 2967 1960
rect 3031 1896 3048 1960
rect 3112 1896 3129 1960
rect 3193 1896 3210 1960
rect 3274 1896 3291 1960
rect 3355 1896 3372 1960
rect 3436 1896 3453 1960
rect 3517 1896 3534 1960
rect 3598 1896 3615 1960
rect 3679 1896 3696 1960
rect 3760 1896 3777 1960
rect 3841 1896 3858 1960
rect 3922 1896 3939 1960
rect 4003 1896 4020 1960
rect 4084 1896 4101 1960
rect 4165 1896 4182 1960
rect 4246 1896 4263 1960
rect 4327 1896 4344 1960
rect 4408 1896 4425 1960
rect 4489 1896 4506 1960
rect 4570 1896 4587 1960
rect 4651 1896 4668 1960
rect 4732 1896 4749 1960
rect 4813 1896 4830 1960
rect 4894 1896 14666 1960
rect 334 1874 14666 1896
rect 354 1810 372 1874
rect 436 1810 454 1874
rect 518 1810 536 1874
rect 600 1810 618 1874
rect 682 1810 699 1874
rect 763 1810 780 1874
rect 844 1810 861 1874
rect 925 1810 942 1874
rect 1006 1810 1023 1874
rect 1087 1810 1104 1874
rect 1168 1810 1185 1874
rect 1249 1810 1266 1874
rect 1330 1810 1347 1874
rect 1411 1810 1428 1874
rect 1492 1810 1509 1874
rect 1573 1810 1590 1874
rect 1654 1810 1671 1874
rect 1735 1810 1752 1874
rect 1816 1810 1833 1874
rect 1897 1810 1914 1874
rect 1978 1810 1995 1874
rect 2059 1810 2076 1874
rect 2140 1810 2157 1874
rect 2221 1810 2238 1874
rect 2302 1810 2319 1874
rect 2383 1810 2400 1874
rect 2464 1810 2481 1874
rect 2545 1810 2562 1874
rect 2626 1810 2643 1874
rect 2707 1810 2724 1874
rect 2788 1810 2805 1874
rect 2869 1810 2886 1874
rect 2950 1810 2967 1874
rect 3031 1810 3048 1874
rect 3112 1810 3129 1874
rect 3193 1810 3210 1874
rect 3274 1810 3291 1874
rect 3355 1810 3372 1874
rect 3436 1810 3453 1874
rect 3517 1810 3534 1874
rect 3598 1810 3615 1874
rect 3679 1810 3696 1874
rect 3760 1810 3777 1874
rect 3841 1810 3858 1874
rect 3922 1810 3939 1874
rect 4003 1810 4020 1874
rect 4084 1810 4101 1874
rect 4165 1810 4182 1874
rect 4246 1810 4263 1874
rect 4327 1810 4344 1874
rect 4408 1810 4425 1874
rect 4489 1810 4506 1874
rect 4570 1810 4587 1874
rect 4651 1810 4668 1874
rect 4732 1810 4749 1874
rect 4813 1810 4830 1874
rect 4894 1810 14666 1874
rect 334 1788 14666 1810
rect 354 1724 372 1788
rect 436 1724 454 1788
rect 518 1724 536 1788
rect 600 1724 618 1788
rect 682 1724 699 1788
rect 763 1724 780 1788
rect 844 1724 861 1788
rect 925 1724 942 1788
rect 1006 1724 1023 1788
rect 1087 1724 1104 1788
rect 1168 1724 1185 1788
rect 1249 1724 1266 1788
rect 1330 1724 1347 1788
rect 1411 1724 1428 1788
rect 1492 1724 1509 1788
rect 1573 1724 1590 1788
rect 1654 1724 1671 1788
rect 1735 1724 1752 1788
rect 1816 1724 1833 1788
rect 1897 1724 1914 1788
rect 1978 1724 1995 1788
rect 2059 1724 2076 1788
rect 2140 1724 2157 1788
rect 2221 1724 2238 1788
rect 2302 1724 2319 1788
rect 2383 1724 2400 1788
rect 2464 1724 2481 1788
rect 2545 1724 2562 1788
rect 2626 1724 2643 1788
rect 2707 1724 2724 1788
rect 2788 1724 2805 1788
rect 2869 1724 2886 1788
rect 2950 1724 2967 1788
rect 3031 1724 3048 1788
rect 3112 1724 3129 1788
rect 3193 1724 3210 1788
rect 3274 1724 3291 1788
rect 3355 1724 3372 1788
rect 3436 1724 3453 1788
rect 3517 1724 3534 1788
rect 3598 1724 3615 1788
rect 3679 1724 3696 1788
rect 3760 1724 3777 1788
rect 3841 1724 3858 1788
rect 3922 1724 3939 1788
rect 4003 1724 4020 1788
rect 4084 1724 4101 1788
rect 4165 1724 4182 1788
rect 4246 1724 4263 1788
rect 4327 1724 4344 1788
rect 4408 1724 4425 1788
rect 4489 1724 4506 1788
rect 4570 1724 4587 1788
rect 4651 1724 4668 1788
rect 4732 1724 4749 1788
rect 4813 1724 4830 1788
rect 4894 1724 14666 1788
rect 334 1702 14666 1724
rect 354 1638 372 1702
rect 436 1638 454 1702
rect 518 1638 536 1702
rect 600 1638 618 1702
rect 682 1638 699 1702
rect 763 1638 780 1702
rect 844 1638 861 1702
rect 925 1638 942 1702
rect 1006 1638 1023 1702
rect 1087 1638 1104 1702
rect 1168 1638 1185 1702
rect 1249 1638 1266 1702
rect 1330 1638 1347 1702
rect 1411 1638 1428 1702
rect 1492 1638 1509 1702
rect 1573 1638 1590 1702
rect 1654 1638 1671 1702
rect 1735 1638 1752 1702
rect 1816 1638 1833 1702
rect 1897 1638 1914 1702
rect 1978 1638 1995 1702
rect 2059 1638 2076 1702
rect 2140 1638 2157 1702
rect 2221 1638 2238 1702
rect 2302 1638 2319 1702
rect 2383 1638 2400 1702
rect 2464 1638 2481 1702
rect 2545 1638 2562 1702
rect 2626 1638 2643 1702
rect 2707 1638 2724 1702
rect 2788 1638 2805 1702
rect 2869 1638 2886 1702
rect 2950 1638 2967 1702
rect 3031 1638 3048 1702
rect 3112 1638 3129 1702
rect 3193 1638 3210 1702
rect 3274 1638 3291 1702
rect 3355 1638 3372 1702
rect 3436 1638 3453 1702
rect 3517 1638 3534 1702
rect 3598 1638 3615 1702
rect 3679 1638 3696 1702
rect 3760 1638 3777 1702
rect 3841 1638 3858 1702
rect 3922 1638 3939 1702
rect 4003 1638 4020 1702
rect 4084 1638 4101 1702
rect 4165 1638 4182 1702
rect 4246 1638 4263 1702
rect 4327 1638 4344 1702
rect 4408 1638 4425 1702
rect 4489 1638 4506 1702
rect 4570 1638 4587 1702
rect 4651 1638 4668 1702
rect 4732 1638 4749 1702
rect 4813 1638 4830 1702
rect 4894 1638 14666 1702
rect 334 1616 14666 1638
rect 354 1552 372 1616
rect 436 1552 454 1616
rect 518 1552 536 1616
rect 600 1552 618 1616
rect 682 1552 699 1616
rect 763 1552 780 1616
rect 844 1552 861 1616
rect 925 1552 942 1616
rect 1006 1552 1023 1616
rect 1087 1552 1104 1616
rect 1168 1552 1185 1616
rect 1249 1552 1266 1616
rect 1330 1552 1347 1616
rect 1411 1552 1428 1616
rect 1492 1552 1509 1616
rect 1573 1552 1590 1616
rect 1654 1552 1671 1616
rect 1735 1552 1752 1616
rect 1816 1552 1833 1616
rect 1897 1552 1914 1616
rect 1978 1552 1995 1616
rect 2059 1552 2076 1616
rect 2140 1552 2157 1616
rect 2221 1552 2238 1616
rect 2302 1552 2319 1616
rect 2383 1552 2400 1616
rect 2464 1552 2481 1616
rect 2545 1552 2562 1616
rect 2626 1552 2643 1616
rect 2707 1552 2724 1616
rect 2788 1552 2805 1616
rect 2869 1552 2886 1616
rect 2950 1552 2967 1616
rect 3031 1552 3048 1616
rect 3112 1552 3129 1616
rect 3193 1552 3210 1616
rect 3274 1552 3291 1616
rect 3355 1552 3372 1616
rect 3436 1552 3453 1616
rect 3517 1552 3534 1616
rect 3598 1552 3615 1616
rect 3679 1552 3696 1616
rect 3760 1552 3777 1616
rect 3841 1552 3858 1616
rect 3922 1552 3939 1616
rect 4003 1552 4020 1616
rect 4084 1552 4101 1616
rect 4165 1552 4182 1616
rect 4246 1552 4263 1616
rect 4327 1552 4344 1616
rect 4408 1552 4425 1616
rect 4489 1552 4506 1616
rect 4570 1552 4587 1616
rect 4651 1552 4668 1616
rect 4732 1552 4749 1616
rect 4813 1552 4830 1616
rect 4894 1552 14666 1616
rect 334 1530 14666 1552
rect 354 1466 372 1530
rect 436 1466 454 1530
rect 518 1466 536 1530
rect 600 1466 618 1530
rect 682 1466 699 1530
rect 763 1466 780 1530
rect 844 1466 861 1530
rect 925 1466 942 1530
rect 1006 1466 1023 1530
rect 1087 1466 1104 1530
rect 1168 1466 1185 1530
rect 1249 1466 1266 1530
rect 1330 1466 1347 1530
rect 1411 1466 1428 1530
rect 1492 1466 1509 1530
rect 1573 1466 1590 1530
rect 1654 1466 1671 1530
rect 1735 1466 1752 1530
rect 1816 1466 1833 1530
rect 1897 1466 1914 1530
rect 1978 1466 1995 1530
rect 2059 1466 2076 1530
rect 2140 1466 2157 1530
rect 2221 1466 2238 1530
rect 2302 1466 2319 1530
rect 2383 1466 2400 1530
rect 2464 1466 2481 1530
rect 2545 1466 2562 1530
rect 2626 1466 2643 1530
rect 2707 1466 2724 1530
rect 2788 1466 2805 1530
rect 2869 1466 2886 1530
rect 2950 1466 2967 1530
rect 3031 1466 3048 1530
rect 3112 1466 3129 1530
rect 3193 1466 3210 1530
rect 3274 1466 3291 1530
rect 3355 1466 3372 1530
rect 3436 1466 3453 1530
rect 3517 1466 3534 1530
rect 3598 1466 3615 1530
rect 3679 1466 3696 1530
rect 3760 1466 3777 1530
rect 3841 1466 3858 1530
rect 3922 1466 3939 1530
rect 4003 1466 4020 1530
rect 4084 1466 4101 1530
rect 4165 1466 4182 1530
rect 4246 1466 4263 1530
rect 4327 1466 4344 1530
rect 4408 1466 4425 1530
rect 4489 1466 4506 1530
rect 4570 1466 4587 1530
rect 4651 1466 4668 1530
rect 4732 1466 4749 1530
rect 4813 1466 4830 1530
rect 4894 1466 14666 1530
rect 334 1444 14666 1466
rect 354 1380 372 1444
rect 436 1380 454 1444
rect 518 1380 536 1444
rect 600 1380 618 1444
rect 682 1380 699 1444
rect 763 1380 780 1444
rect 844 1380 861 1444
rect 925 1380 942 1444
rect 1006 1380 1023 1444
rect 1087 1380 1104 1444
rect 1168 1380 1185 1444
rect 1249 1380 1266 1444
rect 1330 1380 1347 1444
rect 1411 1380 1428 1444
rect 1492 1380 1509 1444
rect 1573 1380 1590 1444
rect 1654 1380 1671 1444
rect 1735 1380 1752 1444
rect 1816 1380 1833 1444
rect 1897 1380 1914 1444
rect 1978 1380 1995 1444
rect 2059 1380 2076 1444
rect 2140 1380 2157 1444
rect 2221 1380 2238 1444
rect 2302 1380 2319 1444
rect 2383 1380 2400 1444
rect 2464 1380 2481 1444
rect 2545 1380 2562 1444
rect 2626 1380 2643 1444
rect 2707 1380 2724 1444
rect 2788 1380 2805 1444
rect 2869 1380 2886 1444
rect 2950 1380 2967 1444
rect 3031 1380 3048 1444
rect 3112 1380 3129 1444
rect 3193 1380 3210 1444
rect 3274 1380 3291 1444
rect 3355 1380 3372 1444
rect 3436 1380 3453 1444
rect 3517 1380 3534 1444
rect 3598 1380 3615 1444
rect 3679 1380 3696 1444
rect 3760 1380 3777 1444
rect 3841 1380 3858 1444
rect 3922 1380 3939 1444
rect 4003 1380 4020 1444
rect 4084 1380 4101 1444
rect 4165 1380 4182 1444
rect 4246 1380 4263 1444
rect 4327 1380 4344 1444
rect 4408 1380 4425 1444
rect 4489 1380 4506 1444
rect 4570 1380 4587 1444
rect 4651 1380 4668 1444
rect 4732 1380 4749 1444
rect 4813 1380 4830 1444
rect 4894 1380 14666 1444
rect 334 1297 14666 1380
rect 193 1177 14807 1297
rect 334 7 14666 1177
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 0 12437 254 13287
rect 0 11267 254 12117
rect 0 9147 254 10947
rect 0 7937 254 8827
rect 0 6968 254 7617
rect 14746 13607 15000 18597
rect 14746 12437 15000 13287
rect 14746 11267 15000 12117
rect 14746 9147 15000 10947
rect 14746 7937 15000 8827
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 0 4787 254 5677
rect 0 3577 254 4467
rect 14746 5997 15000 6647
rect 14746 4787 15000 5677
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 0 27 254 1077
rect 14746 1397 15000 2287
rect 14746 27 15000 1077
<< obsm5 >>
rect 574 34437 14426 39600
rect 0 18917 15000 34437
rect 574 6968 14426 18917
rect 0 6967 15000 6968
rect 574 3257 14426 6967
rect 513 2607 14487 3257
rect 574 27 14426 2607
<< labels >>
rlabel metal5 s 0 12437 254 13287 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 0 12417 254 13307 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 0 3557 254 4487 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 9147 254 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9147 15000 9213 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10881 15000 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 6947 254 7637 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 4 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 6 VCCHIB
port 4 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 6 VCCHIB
port 4 nsew power bidirectional
rlabel metal4 s 0 7 254 1097 6 VCCHIB
port 4 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 5 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 0 1377 254 2307 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10151 1378 14931 2306 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14873 2252 14913 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14873 2166 14913 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14873 2080 14913 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14873 1994 14913 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14873 1908 14913 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14873 1822 14913 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14873 1736 14913 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14873 1650 14913 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14873 1564 14913 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14873 1478 14913 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14873 1392 14913 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14792 2252 14832 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14792 2166 14832 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14792 2080 14832 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14792 1994 14832 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14792 1908 14832 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14792 1822 14832 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14792 1736 14832 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14792 1650 14832 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14792 1564 14832 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14792 1478 14832 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14792 1392 14832 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14711 2252 14751 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14711 2166 14751 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14711 2080 14751 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14711 1994 14751 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14711 1908 14751 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14711 1822 14751 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14711 1736 14751 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14711 1650 14751 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14711 1564 14751 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14711 1478 14751 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14711 1392 14751 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14630 2252 14670 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14630 2166 14670 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14630 2080 14670 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14630 1994 14670 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14630 1908 14670 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14630 1822 14670 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14630 1736 14670 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14630 1650 14670 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14630 1564 14670 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14630 1478 14670 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14630 1392 14670 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14549 2252 14589 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14549 2166 14589 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14549 2080 14589 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14549 1994 14589 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14549 1908 14589 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14549 1822 14589 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14549 1736 14589 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14549 1650 14589 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14549 1564 14589 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14549 1478 14589 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14549 1392 14589 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14468 2252 14508 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14468 2166 14508 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14468 2080 14508 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14468 1994 14508 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14468 1908 14508 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14468 1822 14508 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14468 1736 14508 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14468 1650 14508 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14468 1564 14508 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14468 1478 14508 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14468 1392 14508 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14387 2252 14427 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14387 2166 14427 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14387 2080 14427 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14387 1994 14427 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14387 1908 14427 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14387 1822 14427 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14387 1736 14427 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14387 1650 14427 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14387 1564 14427 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14387 1478 14427 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14387 1392 14427 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14306 2252 14346 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14306 2166 14346 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14306 2080 14346 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14306 1994 14346 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14306 1908 14346 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14306 1822 14346 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14306 1736 14346 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14306 1650 14346 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14306 1564 14346 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14306 1478 14346 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14306 1392 14346 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14225 2252 14265 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14225 2166 14265 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14225 2080 14265 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14225 1994 14265 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14225 1908 14265 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14225 1822 14265 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14225 1736 14265 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14225 1650 14265 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14225 1564 14265 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14225 1478 14265 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14225 1392 14265 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14144 2252 14184 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14144 2166 14184 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14144 2080 14184 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14144 1994 14184 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14144 1908 14184 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14144 1822 14184 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14144 1736 14184 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14144 1650 14184 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14144 1564 14184 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14144 1478 14184 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14144 1392 14184 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14063 2252 14103 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14063 2166 14103 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14063 2080 14103 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14063 1994 14103 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14063 1908 14103 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14063 1822 14103 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14063 1736 14103 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14063 1650 14103 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14063 1564 14103 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14063 1478 14103 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 14063 1392 14103 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13982 2252 14022 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13982 2166 14022 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13982 2080 14022 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13982 1994 14022 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13982 1908 14022 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13982 1822 14022 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13982 1736 14022 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13982 1650 14022 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13982 1564 14022 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13982 1478 14022 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13982 1392 14022 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13901 2252 13941 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13901 2166 13941 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13901 2080 13941 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13901 1994 13941 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13901 1908 13941 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13901 1822 13941 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13901 1736 13941 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13901 1650 13941 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13901 1564 13941 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13901 1478 13941 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13901 1392 13941 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13820 2252 13860 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13820 2166 13860 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13820 2080 13860 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13820 1994 13860 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13820 1908 13860 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13820 1822 13860 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13820 1736 13860 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13820 1650 13860 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13820 1564 13860 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13820 1478 13860 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13820 1392 13860 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13739 2252 13779 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13739 2166 13779 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13739 2080 13779 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13739 1994 13779 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13739 1908 13779 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13739 1822 13779 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13739 1736 13779 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13739 1650 13779 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13739 1564 13779 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13739 1478 13779 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13739 1392 13779 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13658 2252 13698 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13658 2166 13698 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13658 2080 13698 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13658 1994 13698 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13658 1908 13698 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13658 1822 13698 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13658 1736 13698 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13658 1650 13698 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13658 1564 13698 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13658 1478 13698 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13658 1392 13698 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13577 2252 13617 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13577 2166 13617 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13577 2080 13617 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13577 1994 13617 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13577 1908 13617 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13577 1822 13617 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13577 1736 13617 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13577 1650 13617 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13577 1564 13617 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13577 1478 13617 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13577 1392 13617 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13496 2252 13536 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13496 2166 13536 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13496 2080 13536 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13496 1994 13536 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13496 1908 13536 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13496 1822 13536 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13496 1736 13536 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13496 1650 13536 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13496 1564 13536 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13496 1478 13536 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13496 1392 13536 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13415 2252 13455 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13415 2166 13455 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13415 2080 13455 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13415 1994 13455 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13415 1908 13455 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13415 1822 13455 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13415 1736 13455 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13415 1650 13455 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13415 1564 13455 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13415 1478 13455 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13415 1392 13455 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13334 2252 13374 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13334 2166 13374 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13334 2080 13374 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13334 1994 13374 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13334 1908 13374 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13334 1822 13374 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13334 1736 13374 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13334 1650 13374 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13334 1564 13374 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13334 1478 13374 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13334 1392 13374 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13253 2252 13293 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13253 2166 13293 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13253 2080 13293 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13253 1994 13293 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13253 1908 13293 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13253 1822 13293 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13253 1736 13293 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13253 1650 13293 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13253 1564 13293 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13253 1478 13293 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13253 1392 13293 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13172 2252 13212 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13172 2166 13212 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13172 2080 13212 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13172 1994 13212 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13172 1908 13212 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13172 1822 13212 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13172 1736 13212 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13172 1650 13212 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13172 1564 13212 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13172 1478 13212 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13172 1392 13212 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13091 2252 13131 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13091 2166 13131 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13091 2080 13131 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13091 1994 13131 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13091 1908 13131 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13091 1822 13131 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13091 1736 13131 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13091 1650 13131 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13091 1564 13131 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13091 1478 13131 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13091 1392 13131 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13010 2252 13050 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13010 2166 13050 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13010 2080 13050 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13010 1994 13050 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13010 1908 13050 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13010 1822 13050 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13010 1736 13050 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13010 1650 13050 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13010 1564 13050 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13010 1478 13050 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 13010 1392 13050 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12929 2252 12969 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12929 2166 12969 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12929 2080 12969 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12929 1994 12969 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12929 1908 12969 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12929 1822 12969 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12929 1736 12969 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12929 1650 12969 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12929 1564 12969 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12929 1478 12969 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12929 1392 12969 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12848 2252 12888 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12848 2166 12888 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12848 2080 12888 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12848 1994 12888 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12848 1908 12888 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12848 1822 12888 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12848 1736 12888 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12848 1650 12888 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12848 1564 12888 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12848 1478 12888 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12848 1392 12888 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12767 2252 12807 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12767 2166 12807 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12767 2080 12807 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12767 1994 12807 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12767 1908 12807 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12767 1822 12807 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12767 1736 12807 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12767 1650 12807 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12767 1564 12807 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12767 1478 12807 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12767 1392 12807 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12686 2252 12726 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12686 2166 12726 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12686 2080 12726 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12686 1994 12726 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12686 1908 12726 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12686 1822 12726 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12686 1736 12726 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12686 1650 12726 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12686 1564 12726 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12686 1478 12726 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12686 1392 12726 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12605 2252 12645 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12605 2166 12645 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12605 2080 12645 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12605 1994 12645 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12605 1908 12645 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12605 1822 12645 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12605 1736 12645 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12605 1650 12645 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12605 1564 12645 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12605 1478 12645 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12605 1392 12645 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12524 2252 12564 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12524 2166 12564 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12524 2080 12564 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12524 1994 12564 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12524 1908 12564 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12524 1822 12564 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12524 1736 12564 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12524 1650 12564 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12524 1564 12564 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12524 1478 12564 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12524 1392 12564 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12443 2252 12483 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12443 2166 12483 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12443 2080 12483 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12443 1994 12483 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12443 1908 12483 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12443 1822 12483 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12443 1736 12483 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12443 1650 12483 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12443 1564 12483 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12443 1478 12483 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12443 1392 12483 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12362 2252 12402 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12362 2166 12402 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12362 2080 12402 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12362 1994 12402 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12362 1908 12402 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12362 1822 12402 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12362 1736 12402 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12362 1650 12402 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12362 1564 12402 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12362 1478 12402 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12362 1392 12402 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12281 2252 12321 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12281 2166 12321 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12281 2080 12321 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12281 1994 12321 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12281 1908 12321 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12281 1822 12321 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12281 1736 12321 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12281 1650 12321 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12281 1564 12321 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12281 1478 12321 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12281 1392 12321 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12200 2252 12240 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12200 2166 12240 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12200 2080 12240 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12200 1994 12240 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12200 1908 12240 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12200 1822 12240 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12200 1736 12240 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12200 1650 12240 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12200 1564 12240 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12200 1478 12240 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12200 1392 12240 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12119 2252 12159 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12119 2166 12159 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12119 2080 12159 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12119 1994 12159 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12119 1908 12159 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12119 1822 12159 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12119 1736 12159 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12119 1650 12159 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12119 1564 12159 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12119 1478 12159 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12119 1392 12159 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12038 2252 12078 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12038 2166 12078 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12038 2080 12078 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12038 1994 12078 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12038 1908 12078 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12038 1822 12078 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12038 1736 12078 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12038 1650 12078 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12038 1564 12078 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12038 1478 12078 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 12038 1392 12078 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11957 2252 11997 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11957 2166 11997 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11957 2080 11997 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11957 1994 11997 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11957 1908 11997 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11957 1822 11997 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11957 1736 11997 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11957 1650 11997 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11957 1564 11997 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11957 1478 11997 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11957 1392 11997 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11876 2252 11916 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11876 2166 11916 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11876 2080 11916 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11876 1994 11916 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11876 1908 11916 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11876 1822 11916 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11876 1736 11916 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11876 1650 11916 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11876 1564 11916 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11876 1478 11916 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11876 1392 11916 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11795 2252 11835 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11795 2166 11835 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11795 2080 11835 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11795 1994 11835 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11795 1908 11835 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11795 1822 11835 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11795 1736 11835 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11795 1650 11835 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11795 1564 11835 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11795 1478 11835 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11795 1392 11835 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11714 2252 11754 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11714 2166 11754 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11714 2080 11754 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11714 1994 11754 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11714 1908 11754 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11714 1822 11754 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11714 1736 11754 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11714 1650 11754 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11714 1564 11754 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11714 1478 11754 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11714 1392 11754 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11633 2252 11673 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11633 2166 11673 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11633 2080 11673 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11633 1994 11673 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11633 1908 11673 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11633 1822 11673 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11633 1736 11673 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11633 1650 11673 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11633 1564 11673 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11633 1478 11673 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11633 1392 11673 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11552 2252 11592 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11552 2166 11592 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11552 2080 11592 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11552 1994 11592 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11552 1908 11592 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11552 1822 11592 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11552 1736 11592 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11552 1650 11592 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11552 1564 11592 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11552 1478 11592 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11552 1392 11592 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11471 2252 11511 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11471 2166 11511 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11471 2080 11511 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11471 1994 11511 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11471 1908 11511 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11471 1822 11511 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11471 1736 11511 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11471 1650 11511 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11471 1564 11511 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11471 1478 11511 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11471 1392 11511 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11390 2252 11430 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11390 2166 11430 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11390 2080 11430 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11390 1994 11430 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11390 1908 11430 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11390 1822 11430 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11390 1736 11430 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11390 1650 11430 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11390 1564 11430 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11390 1478 11430 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11390 1392 11430 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11309 2252 11349 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11309 2166 11349 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11309 2080 11349 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11309 1994 11349 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11309 1908 11349 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11309 1822 11349 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11309 1736 11349 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11309 1650 11349 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11309 1564 11349 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11309 1478 11349 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11309 1392 11349 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11228 2252 11268 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11228 2166 11268 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11228 2080 11268 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11228 1994 11268 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11228 1908 11268 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11228 1822 11268 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11228 1736 11268 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11228 1650 11268 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11228 1564 11268 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11228 1478 11268 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11228 1392 11268 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11147 2252 11187 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11147 2166 11187 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11147 2080 11187 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11147 1994 11187 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11147 1908 11187 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11147 1822 11187 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11147 1736 11187 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11147 1650 11187 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11147 1564 11187 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11147 1478 11187 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11147 1392 11187 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11066 2252 11106 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11066 2166 11106 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11066 2080 11106 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11066 1994 11106 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11066 1908 11106 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11066 1822 11106 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11066 1736 11106 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11066 1650 11106 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11066 1564 11106 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11066 1478 11106 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 11066 1392 11106 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10985 2252 11025 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10985 2166 11025 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10985 2080 11025 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10985 1994 11025 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10985 1908 11025 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10985 1822 11025 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10985 1736 11025 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10985 1650 11025 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10985 1564 11025 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10985 1478 11025 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10985 1392 11025 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10904 2252 10944 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10904 2166 10944 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10904 2080 10944 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10904 1994 10944 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10904 1908 10944 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10904 1822 10944 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10904 1736 10944 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10904 1650 10944 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10904 1564 10944 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10904 1478 10944 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10904 1392 10944 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10823 2252 10863 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10823 2166 10863 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10823 2080 10863 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10823 1994 10863 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10823 1908 10863 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10823 1822 10863 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10823 1736 10863 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10823 1650 10863 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10823 1564 10863 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10823 1478 10863 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10823 1392 10863 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10742 2252 10782 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10742 2166 10782 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10742 2080 10782 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10742 1994 10782 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10742 1908 10782 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10742 1822 10782 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10742 1736 10782 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10742 1650 10782 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10742 1564 10782 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10742 1478 10782 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10742 1392 10782 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10661 2252 10701 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10661 2166 10701 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10661 2080 10701 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10661 1994 10701 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10661 1908 10701 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10661 1822 10701 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10661 1736 10701 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10661 1650 10701 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10661 1564 10701 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10661 1478 10701 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10661 1392 10701 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10579 2252 10619 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10579 2166 10619 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10579 2080 10619 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10579 1994 10619 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10579 1908 10619 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10579 1822 10619 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10579 1736 10619 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10579 1650 10619 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10579 1564 10619 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10579 1478 10619 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10579 1392 10619 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10497 2252 10537 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10497 2166 10537 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10497 2080 10537 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10497 1994 10537 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10497 1908 10537 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10497 1822 10537 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10497 1736 10537 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10497 1650 10537 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10497 1564 10537 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10497 1478 10537 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10497 1392 10537 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10415 2252 10455 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10415 2166 10455 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10415 2080 10455 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10415 1994 10455 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10415 1908 10455 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10415 1822 10455 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10415 1736 10455 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10415 1650 10455 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10415 1564 10455 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10415 1478 10455 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10415 1392 10455 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10333 2252 10373 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10333 2166 10373 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10333 2080 10373 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10333 1994 10373 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10333 1908 10373 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10333 1822 10373 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10333 1736 10373 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10333 1650 10373 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10333 1564 10373 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10333 1478 10373 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10333 1392 10373 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10251 2252 10291 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10251 2166 10291 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10251 2080 10291 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10251 1994 10291 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10251 1908 10291 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10251 1822 10291 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10251 1736 10291 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10251 1650 10291 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10251 1564 10291 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10251 1478 10291 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10251 1392 10291 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10169 2252 10209 2292 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10169 2166 10209 2206 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10169 2080 10209 2120 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10169 1994 10209 2034 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10169 1908 10209 1948 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10169 1822 10209 1862 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10169 1736 10209 1776 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10169 1650 10209 1690 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10169 1564 10209 1604 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10169 1478 10209 1518 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 10169 1392 10209 1432 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4830 2240 4894 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4830 2240 4894 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4830 2154 4894 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4830 2154 4894 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4830 2068 4894 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4830 2068 4894 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4830 1982 4894 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4830 1982 4894 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4830 1896 4894 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4830 1896 4894 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4830 1810 4894 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4830 1810 4894 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4830 1724 4894 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4830 1724 4894 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4830 1638 4894 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4830 1638 4894 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4830 1552 4894 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4830 1552 4894 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4830 1466 4894 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4830 1466 4894 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4830 1380 4894 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4830 1380 4894 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4749 2240 4813 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4749 2240 4813 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4749 2154 4813 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4749 2154 4813 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4749 2068 4813 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4749 2068 4813 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4749 1982 4813 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4749 1982 4813 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4749 1896 4813 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4749 1896 4813 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4749 1810 4813 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4749 1810 4813 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4749 1724 4813 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4749 1724 4813 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4749 1638 4813 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4749 1638 4813 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4749 1552 4813 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4749 1552 4813 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4749 1466 4813 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4749 1466 4813 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4749 1380 4813 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4749 1380 4813 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4668 2240 4732 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4668 2240 4732 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4668 2154 4732 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4668 2154 4732 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4668 2068 4732 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4668 2068 4732 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4668 1982 4732 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4668 1982 4732 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4668 1896 4732 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4668 1896 4732 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4668 1810 4732 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4668 1810 4732 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4668 1724 4732 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4668 1724 4732 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4668 1638 4732 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4668 1638 4732 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4668 1552 4732 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4668 1552 4732 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4668 1466 4732 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4668 1466 4732 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4668 1380 4732 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4668 1380 4732 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4587 2240 4651 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4587 2240 4651 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4587 2154 4651 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4587 2154 4651 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4587 2068 4651 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4587 2068 4651 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4587 1982 4651 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4587 1982 4651 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4587 1896 4651 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4587 1896 4651 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4587 1810 4651 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4587 1810 4651 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4587 1724 4651 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4587 1724 4651 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4587 1638 4651 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4587 1638 4651 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4587 1552 4651 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4587 1552 4651 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4587 1466 4651 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4587 1466 4651 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4587 1380 4651 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4587 1380 4651 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4506 2240 4570 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4506 2240 4570 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4506 2154 4570 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4506 2154 4570 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4506 2068 4570 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4506 2068 4570 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4506 1982 4570 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4506 1982 4570 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4506 1896 4570 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4506 1896 4570 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4506 1810 4570 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4506 1810 4570 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4506 1724 4570 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4506 1724 4570 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4506 1638 4570 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4506 1638 4570 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4506 1552 4570 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4506 1552 4570 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4506 1466 4570 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4506 1466 4570 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4506 1380 4570 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4506 1380 4570 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4425 2240 4489 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4425 2240 4489 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4425 2154 4489 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4425 2154 4489 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4425 2068 4489 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4425 2068 4489 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4425 1982 4489 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4425 1982 4489 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4425 1896 4489 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4425 1896 4489 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4425 1810 4489 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4425 1810 4489 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4425 1724 4489 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4425 1724 4489 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4425 1638 4489 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4425 1638 4489 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4425 1552 4489 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4425 1552 4489 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4425 1466 4489 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4425 1466 4489 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4425 1380 4489 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4425 1380 4489 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4344 2240 4408 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4344 2240 4408 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4344 2154 4408 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4344 2154 4408 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4344 2068 4408 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4344 2068 4408 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4344 1982 4408 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4344 1982 4408 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4344 1896 4408 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4344 1896 4408 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4344 1810 4408 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4344 1810 4408 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4344 1724 4408 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4344 1724 4408 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4344 1638 4408 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4344 1638 4408 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4344 1552 4408 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4344 1552 4408 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4344 1466 4408 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4344 1466 4408 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4344 1380 4408 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4344 1380 4408 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4263 2240 4327 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4263 2240 4327 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4263 2154 4327 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4263 2154 4327 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4263 2068 4327 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4263 2068 4327 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4263 1982 4327 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4263 1982 4327 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4263 1896 4327 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4263 1896 4327 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4263 1810 4327 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4263 1810 4327 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4263 1724 4327 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4263 1724 4327 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4263 1638 4327 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4263 1638 4327 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4263 1552 4327 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4263 1552 4327 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4263 1466 4327 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4263 1466 4327 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4263 1380 4327 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4263 1380 4327 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4182 2240 4246 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4182 2240 4246 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4182 2154 4246 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4182 2154 4246 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4182 2068 4246 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4182 2068 4246 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4182 1982 4246 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4182 1982 4246 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4182 1896 4246 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4182 1896 4246 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4182 1810 4246 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4182 1810 4246 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4182 1724 4246 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4182 1724 4246 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4182 1638 4246 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4182 1638 4246 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4182 1552 4246 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4182 1552 4246 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4182 1466 4246 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4182 1466 4246 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4182 1380 4246 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4182 1380 4246 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4101 2240 4165 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4101 2240 4165 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4101 2154 4165 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4101 2154 4165 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4101 2068 4165 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4101 2068 4165 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4101 1982 4165 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4101 1982 4165 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4101 1896 4165 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4101 1896 4165 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4101 1810 4165 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4101 1810 4165 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4101 1724 4165 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4101 1724 4165 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4101 1638 4165 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4101 1638 4165 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4101 1552 4165 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4101 1552 4165 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4101 1466 4165 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4101 1466 4165 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4101 1380 4165 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4101 1380 4165 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4020 2240 4084 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4020 2240 4084 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4020 2154 4084 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4020 2154 4084 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4020 2068 4084 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4020 2068 4084 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4020 1982 4084 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4020 1982 4084 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4020 1896 4084 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4020 1896 4084 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4020 1810 4084 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4020 1810 4084 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4020 1724 4084 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4020 1724 4084 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4020 1638 4084 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4020 1638 4084 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4020 1552 4084 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4020 1552 4084 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4020 1466 4084 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4020 1466 4084 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 4020 1380 4084 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 4020 1380 4084 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3939 2240 4003 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3939 2240 4003 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3939 2154 4003 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3939 2154 4003 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3939 2068 4003 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3939 2068 4003 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3939 1982 4003 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3939 1982 4003 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3939 1896 4003 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3939 1896 4003 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3939 1810 4003 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3939 1810 4003 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3939 1724 4003 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3939 1724 4003 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3939 1638 4003 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3939 1638 4003 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3939 1552 4003 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3939 1552 4003 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3939 1466 4003 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3939 1466 4003 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3939 1380 4003 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3939 1380 4003 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3858 2240 3922 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3858 2240 3922 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3858 2154 3922 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3858 2154 3922 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3858 2068 3922 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3858 2068 3922 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3858 1982 3922 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3858 1982 3922 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3858 1896 3922 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3858 1896 3922 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3858 1810 3922 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3858 1810 3922 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3858 1724 3922 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3858 1724 3922 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3858 1638 3922 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3858 1638 3922 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3858 1552 3922 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3858 1552 3922 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3858 1466 3922 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3858 1466 3922 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3858 1380 3922 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3858 1380 3922 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3777 2240 3841 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3777 2240 3841 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3777 2154 3841 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3777 2154 3841 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3777 2068 3841 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3777 2068 3841 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3777 1982 3841 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3777 1982 3841 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3777 1896 3841 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3777 1896 3841 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3777 1810 3841 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3777 1810 3841 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3777 1724 3841 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3777 1724 3841 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3777 1638 3841 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3777 1638 3841 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3777 1552 3841 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3777 1552 3841 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3777 1466 3841 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3777 1466 3841 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3777 1380 3841 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3777 1380 3841 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3696 2240 3760 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3696 2240 3760 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3696 2154 3760 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3696 2154 3760 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3696 2068 3760 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3696 2068 3760 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3696 1982 3760 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3696 1982 3760 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3696 1896 3760 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3696 1896 3760 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3696 1810 3760 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3696 1810 3760 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3696 1724 3760 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3696 1724 3760 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3696 1638 3760 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3696 1638 3760 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3696 1552 3760 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3696 1552 3760 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3696 1466 3760 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3696 1466 3760 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3696 1380 3760 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3696 1380 3760 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3615 2240 3679 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3615 2240 3679 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3615 2154 3679 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3615 2154 3679 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3615 2068 3679 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3615 2068 3679 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3615 1982 3679 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3615 1982 3679 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3615 1896 3679 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3615 1896 3679 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3615 1810 3679 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3615 1810 3679 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3615 1724 3679 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3615 1724 3679 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3615 1638 3679 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3615 1638 3679 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3615 1552 3679 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3615 1552 3679 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3615 1466 3679 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3615 1466 3679 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3615 1380 3679 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3615 1380 3679 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3534 2240 3598 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3534 2240 3598 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3534 2154 3598 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3534 2154 3598 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3534 2068 3598 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3534 2068 3598 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3534 1982 3598 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3534 1982 3598 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3534 1896 3598 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3534 1896 3598 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3534 1810 3598 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3534 1810 3598 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3534 1724 3598 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3534 1724 3598 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3534 1638 3598 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3534 1638 3598 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3534 1552 3598 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3534 1552 3598 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3534 1466 3598 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3534 1466 3598 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3534 1380 3598 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3534 1380 3598 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3453 2240 3517 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3453 2240 3517 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3453 2154 3517 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3453 2154 3517 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3453 2068 3517 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3453 2068 3517 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3453 1982 3517 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3453 1982 3517 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3453 1896 3517 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3453 1896 3517 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3453 1810 3517 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3453 1810 3517 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3453 1724 3517 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3453 1724 3517 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3453 1638 3517 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3453 1638 3517 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3453 1552 3517 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3453 1552 3517 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3453 1466 3517 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3453 1466 3517 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3453 1380 3517 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3453 1380 3517 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3372 2240 3436 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3372 2240 3436 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3372 2154 3436 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3372 2154 3436 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3372 2068 3436 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3372 2068 3436 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3372 1982 3436 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3372 1982 3436 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3372 1896 3436 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3372 1896 3436 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3372 1810 3436 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3372 1810 3436 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3372 1724 3436 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3372 1724 3436 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3372 1638 3436 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3372 1638 3436 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3372 1552 3436 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3372 1552 3436 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3372 1466 3436 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3372 1466 3436 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3372 1380 3436 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3372 1380 3436 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3291 2240 3355 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3291 2240 3355 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3291 2154 3355 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3291 2154 3355 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3291 2068 3355 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3291 2068 3355 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3291 1982 3355 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3291 1982 3355 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3291 1896 3355 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3291 1896 3355 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3291 1810 3355 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3291 1810 3355 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3291 1724 3355 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3291 1724 3355 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3291 1638 3355 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3291 1638 3355 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3291 1552 3355 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3291 1552 3355 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3291 1466 3355 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3291 1466 3355 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3291 1380 3355 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3291 1380 3355 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3210 2240 3274 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3210 2240 3274 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3210 2154 3274 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3210 2154 3274 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3210 2068 3274 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3210 2068 3274 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3210 1982 3274 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3210 1982 3274 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3210 1896 3274 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3210 1896 3274 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3210 1810 3274 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3210 1810 3274 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3210 1724 3274 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3210 1724 3274 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3210 1638 3274 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3210 1638 3274 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3210 1552 3274 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3210 1552 3274 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3210 1466 3274 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3210 1466 3274 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3210 1380 3274 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3210 1380 3274 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3129 2240 3193 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3129 2240 3193 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3129 2154 3193 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3129 2154 3193 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3129 2068 3193 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3129 2068 3193 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3129 1982 3193 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3129 1982 3193 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3129 1896 3193 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3129 1896 3193 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3129 1810 3193 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3129 1810 3193 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3129 1724 3193 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3129 1724 3193 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3129 1638 3193 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3129 1638 3193 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3129 1552 3193 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3129 1552 3193 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3129 1466 3193 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3129 1466 3193 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3129 1380 3193 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3129 1380 3193 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3048 2240 3112 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3048 2240 3112 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3048 2154 3112 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3048 2154 3112 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3048 2068 3112 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3048 2068 3112 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3048 1982 3112 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3048 1982 3112 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3048 1896 3112 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3048 1896 3112 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3048 1810 3112 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3048 1810 3112 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3048 1724 3112 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3048 1724 3112 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3048 1638 3112 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3048 1638 3112 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3048 1552 3112 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3048 1552 3112 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3048 1466 3112 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3048 1466 3112 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 3048 1380 3112 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 3048 1380 3112 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2967 2240 3031 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2967 2240 3031 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2967 2154 3031 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2967 2154 3031 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2967 2068 3031 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2967 2068 3031 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2967 1982 3031 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2967 1982 3031 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2967 1896 3031 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2967 1896 3031 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2967 1810 3031 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2967 1810 3031 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2967 1724 3031 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2967 1724 3031 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2967 1638 3031 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2967 1638 3031 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2967 1552 3031 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2967 1552 3031 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2967 1466 3031 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2967 1466 3031 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2967 1380 3031 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2967 1380 3031 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2886 2240 2950 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2886 2240 2950 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2886 2154 2950 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2886 2154 2950 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2886 2068 2950 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2886 2068 2950 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2886 1982 2950 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2886 1982 2950 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2886 1896 2950 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2886 1896 2950 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2886 1810 2950 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2886 1810 2950 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2886 1724 2950 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2886 1724 2950 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2886 1638 2950 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2886 1638 2950 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2886 1552 2950 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2886 1552 2950 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2886 1466 2950 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2886 1466 2950 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2886 1380 2950 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2886 1380 2950 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2805 2240 2869 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2805 2240 2869 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2805 2154 2869 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2805 2154 2869 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2805 2068 2869 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2805 2068 2869 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2805 1982 2869 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2805 1982 2869 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2805 1896 2869 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2805 1896 2869 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2805 1810 2869 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2805 1810 2869 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2805 1724 2869 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2805 1724 2869 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2805 1638 2869 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2805 1638 2869 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2805 1552 2869 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2805 1552 2869 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2805 1466 2869 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2805 1466 2869 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2805 1380 2869 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2805 1380 2869 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2724 2240 2788 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2724 2240 2788 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2724 2154 2788 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2724 2154 2788 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2724 2068 2788 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2724 2068 2788 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2724 1982 2788 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2724 1982 2788 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2724 1896 2788 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2724 1896 2788 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2724 1810 2788 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2724 1810 2788 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2724 1724 2788 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2724 1724 2788 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2724 1638 2788 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2724 1638 2788 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2724 1552 2788 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2724 1552 2788 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2724 1466 2788 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2724 1466 2788 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2724 1380 2788 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2724 1380 2788 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2643 2240 2707 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2643 2240 2707 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2643 2154 2707 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2643 2154 2707 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2643 2068 2707 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2643 2068 2707 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2643 1982 2707 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2643 1982 2707 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2643 1896 2707 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2643 1896 2707 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2643 1810 2707 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2643 1810 2707 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2643 1724 2707 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2643 1724 2707 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2643 1638 2707 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2643 1638 2707 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2643 1552 2707 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2643 1552 2707 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2643 1466 2707 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2643 1466 2707 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2643 1380 2707 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2643 1380 2707 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2562 2240 2626 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2562 2240 2626 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2562 2154 2626 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2562 2154 2626 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2562 2068 2626 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2562 2068 2626 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2562 1982 2626 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2562 1982 2626 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2562 1896 2626 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2562 1896 2626 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2562 1810 2626 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2562 1810 2626 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2562 1724 2626 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2562 1724 2626 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2562 1638 2626 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2562 1638 2626 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2562 1552 2626 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2562 1552 2626 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2562 1466 2626 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2562 1466 2626 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2562 1380 2626 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2562 1380 2626 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2481 2240 2545 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2481 2240 2545 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2481 2154 2545 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2481 2154 2545 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2481 2068 2545 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2481 2068 2545 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2481 1982 2545 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2481 1982 2545 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2481 1896 2545 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2481 1896 2545 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2481 1810 2545 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2481 1810 2545 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2481 1724 2545 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2481 1724 2545 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2481 1638 2545 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2481 1638 2545 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2481 1552 2545 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2481 1552 2545 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2481 1466 2545 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2481 1466 2545 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2481 1380 2545 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2481 1380 2545 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2400 2240 2464 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2400 2240 2464 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2400 2154 2464 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2400 2154 2464 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2400 2068 2464 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2400 2068 2464 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2400 1982 2464 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2400 1982 2464 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2400 1896 2464 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2400 1896 2464 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2400 1810 2464 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2400 1810 2464 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2400 1724 2464 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2400 1724 2464 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2400 1638 2464 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2400 1638 2464 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2400 1552 2464 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2400 1552 2464 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2400 1466 2464 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2400 1466 2464 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2400 1380 2464 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2400 1380 2464 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2319 2240 2383 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2319 2240 2383 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2319 2154 2383 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2319 2154 2383 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2319 2068 2383 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2319 2068 2383 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2319 1982 2383 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2319 1982 2383 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2319 1896 2383 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2319 1896 2383 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2319 1810 2383 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2319 1810 2383 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2319 1724 2383 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2319 1724 2383 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2319 1638 2383 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2319 1638 2383 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2319 1552 2383 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2319 1552 2383 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2319 1466 2383 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2319 1466 2383 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2319 1380 2383 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2319 1380 2383 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2238 2240 2302 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2238 2240 2302 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2238 2154 2302 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2238 2154 2302 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2238 2068 2302 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2238 2068 2302 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2238 1982 2302 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2238 1982 2302 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2238 1896 2302 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2238 1896 2302 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2238 1810 2302 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2238 1810 2302 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2238 1724 2302 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2238 1724 2302 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2238 1638 2302 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2238 1638 2302 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2238 1552 2302 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2238 1552 2302 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2238 1466 2302 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2238 1466 2302 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2238 1380 2302 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2238 1380 2302 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2157 2240 2221 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2157 2240 2221 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2157 2154 2221 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2157 2154 2221 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2157 2068 2221 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2157 2068 2221 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2157 1982 2221 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2157 1982 2221 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2157 1896 2221 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2157 1896 2221 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2157 1810 2221 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2157 1810 2221 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2157 1724 2221 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2157 1724 2221 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2157 1638 2221 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2157 1638 2221 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2157 1552 2221 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2157 1552 2221 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2157 1466 2221 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2157 1466 2221 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2157 1380 2221 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2157 1380 2221 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2076 2240 2140 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2076 2240 2140 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2076 2154 2140 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2076 2154 2140 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2076 2068 2140 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2076 2068 2140 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2076 1982 2140 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2076 1982 2140 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2076 1896 2140 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2076 1896 2140 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2076 1810 2140 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2076 1810 2140 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2076 1724 2140 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2076 1724 2140 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2076 1638 2140 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2076 1638 2140 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2076 1552 2140 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2076 1552 2140 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2076 1466 2140 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2076 1466 2140 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 2076 1380 2140 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 2076 1380 2140 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1995 2240 2059 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1995 2240 2059 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1995 2154 2059 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1995 2154 2059 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1995 2068 2059 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1995 2068 2059 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1995 1982 2059 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1995 1982 2059 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1995 1896 2059 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1995 1896 2059 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1995 1810 2059 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1995 1810 2059 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1995 1724 2059 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1995 1724 2059 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1995 1638 2059 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1995 1638 2059 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1995 1552 2059 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1995 1552 2059 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1995 1466 2059 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1995 1466 2059 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1995 1380 2059 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1995 1380 2059 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1914 2240 1978 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1914 2240 1978 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1914 2154 1978 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1914 2154 1978 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1914 2068 1978 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1914 2068 1978 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1914 1982 1978 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1914 1982 1978 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1914 1896 1978 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1914 1896 1978 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1914 1810 1978 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1914 1810 1978 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1914 1724 1978 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1914 1724 1978 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1914 1638 1978 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1914 1638 1978 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1914 1552 1978 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1914 1552 1978 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1914 1466 1978 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1914 1466 1978 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1914 1380 1978 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1914 1380 1978 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1833 2240 1897 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1833 2240 1897 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1833 2154 1897 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1833 2154 1897 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1833 2068 1897 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1833 2068 1897 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1833 1982 1897 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1833 1982 1897 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1833 1896 1897 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1833 1896 1897 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1833 1810 1897 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1833 1810 1897 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1833 1724 1897 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1833 1724 1897 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1833 1638 1897 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1833 1638 1897 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1833 1552 1897 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1833 1552 1897 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1833 1466 1897 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1833 1466 1897 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1833 1380 1897 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1833 1380 1897 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1752 2240 1816 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1752 2240 1816 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1752 2154 1816 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1752 2154 1816 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1752 2068 1816 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1752 2068 1816 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1752 1982 1816 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1752 1982 1816 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1752 1896 1816 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1752 1896 1816 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1752 1810 1816 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1752 1810 1816 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1752 1724 1816 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1752 1724 1816 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1752 1638 1816 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1752 1638 1816 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1752 1552 1816 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1752 1552 1816 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1752 1466 1816 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1752 1466 1816 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1752 1380 1816 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1752 1380 1816 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1671 2240 1735 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1671 2240 1735 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1671 2154 1735 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1671 2154 1735 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1671 2068 1735 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1671 2068 1735 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1671 1982 1735 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1671 1982 1735 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1671 1896 1735 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1671 1896 1735 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1671 1810 1735 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1671 1810 1735 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1671 1724 1735 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1671 1724 1735 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1671 1638 1735 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1671 1638 1735 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1671 1552 1735 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1671 1552 1735 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1671 1466 1735 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1671 1466 1735 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1671 1380 1735 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1671 1380 1735 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1590 2240 1654 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1590 2240 1654 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1590 2154 1654 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1590 2154 1654 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1590 2068 1654 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1590 2068 1654 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1590 1982 1654 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1590 1982 1654 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1590 1896 1654 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1590 1896 1654 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1590 1810 1654 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1590 1810 1654 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1590 1724 1654 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1590 1724 1654 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1590 1638 1654 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1590 1638 1654 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1590 1552 1654 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1590 1552 1654 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1590 1466 1654 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1590 1466 1654 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1590 1380 1654 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1590 1380 1654 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1509 2240 1573 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1509 2240 1573 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1509 2154 1573 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1509 2154 1573 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1509 2068 1573 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1509 2068 1573 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1509 1982 1573 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1509 1982 1573 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1509 1896 1573 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1509 1896 1573 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1509 1810 1573 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1509 1810 1573 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1509 1724 1573 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1509 1724 1573 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1509 1638 1573 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1509 1638 1573 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1509 1552 1573 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1509 1552 1573 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1509 1466 1573 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1509 1466 1573 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1509 1380 1573 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1509 1380 1573 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1428 2240 1492 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1428 2240 1492 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1428 2154 1492 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1428 2154 1492 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1428 2068 1492 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1428 2068 1492 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1428 1982 1492 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1428 1982 1492 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1428 1896 1492 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1428 1896 1492 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1428 1810 1492 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1428 1810 1492 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1428 1724 1492 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1428 1724 1492 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1428 1638 1492 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1428 1638 1492 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1428 1552 1492 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1428 1552 1492 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1428 1466 1492 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1428 1466 1492 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1428 1380 1492 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1428 1380 1492 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1347 2240 1411 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1347 2240 1411 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1347 2154 1411 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1347 2154 1411 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1347 2068 1411 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1347 2068 1411 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1347 1982 1411 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1347 1982 1411 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1347 1896 1411 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1347 1896 1411 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1347 1810 1411 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1347 1810 1411 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1347 1724 1411 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1347 1724 1411 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1347 1638 1411 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1347 1638 1411 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1347 1552 1411 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1347 1552 1411 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1347 1466 1411 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1347 1466 1411 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1347 1380 1411 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1347 1380 1411 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1266 2240 1330 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1266 2240 1330 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1266 2154 1330 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1266 2154 1330 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1266 2068 1330 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1266 2068 1330 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1266 1982 1330 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1266 1982 1330 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1266 1896 1330 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1266 1896 1330 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1266 1810 1330 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1266 1810 1330 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1266 1724 1330 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1266 1724 1330 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1266 1638 1330 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1266 1638 1330 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1266 1552 1330 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1266 1552 1330 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1266 1466 1330 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1266 1466 1330 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1266 1380 1330 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1266 1380 1330 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1185 2240 1249 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1185 2240 1249 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1185 2154 1249 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1185 2154 1249 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1185 2068 1249 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1185 2068 1249 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1185 1982 1249 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1185 1982 1249 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1185 1896 1249 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1185 1896 1249 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1185 1810 1249 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1185 1810 1249 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1185 1724 1249 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1185 1724 1249 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1185 1638 1249 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1185 1638 1249 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1185 1552 1249 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1185 1552 1249 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1185 1466 1249 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1185 1466 1249 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1185 1380 1249 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1185 1380 1249 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1104 2240 1168 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1104 2240 1168 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1104 2154 1168 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1104 2154 1168 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1104 2068 1168 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1104 2068 1168 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1104 1982 1168 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1104 1982 1168 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1104 1896 1168 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1104 1896 1168 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1104 1810 1168 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1104 1810 1168 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1104 1724 1168 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1104 1724 1168 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1104 1638 1168 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1104 1638 1168 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1104 1552 1168 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1104 1552 1168 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1104 1466 1168 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1104 1466 1168 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1104 1380 1168 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1104 1380 1168 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1023 2240 1087 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1023 2240 1087 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1023 2154 1087 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1023 2154 1087 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1023 2068 1087 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1023 2068 1087 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1023 1982 1087 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1023 1982 1087 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1023 1896 1087 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1023 1896 1087 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1023 1810 1087 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1023 1810 1087 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1023 1724 1087 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1023 1724 1087 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1023 1638 1087 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1023 1638 1087 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1023 1552 1087 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1023 1552 1087 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1023 1466 1087 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1023 1466 1087 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 1023 1380 1087 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 1023 1380 1087 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 942 2240 1006 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 942 2240 1006 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 942 2154 1006 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 942 2154 1006 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 942 2068 1006 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 942 2068 1006 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 942 1982 1006 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 942 1982 1006 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 942 1896 1006 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 942 1896 1006 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 942 1810 1006 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 942 1810 1006 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 942 1724 1006 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 942 1724 1006 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 942 1638 1006 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 942 1638 1006 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 942 1552 1006 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 942 1552 1006 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 942 1466 1006 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 942 1466 1006 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 942 1380 1006 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 942 1380 1006 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 861 2240 925 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 861 2240 925 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 861 2154 925 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 861 2154 925 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 861 2068 925 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 861 2068 925 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 861 1982 925 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 861 1982 925 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 861 1896 925 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 861 1896 925 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 861 1810 925 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 861 1810 925 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 861 1724 925 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 861 1724 925 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 861 1638 925 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 861 1638 925 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 861 1552 925 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 861 1552 925 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 861 1466 925 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 861 1466 925 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 861 1380 925 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 861 1380 925 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 780 2240 844 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 780 2240 844 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 780 2154 844 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 780 2154 844 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 780 2068 844 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 780 2068 844 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 780 1982 844 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 780 1982 844 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 780 1896 844 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 780 1896 844 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 780 1810 844 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 780 1810 844 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 780 1724 844 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 780 1724 844 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 780 1638 844 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 780 1638 844 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 780 1552 844 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 780 1552 844 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 780 1466 844 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 780 1466 844 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 780 1380 844 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 780 1380 844 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 699 2240 763 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 699 2240 763 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 699 2154 763 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 699 2154 763 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 699 2068 763 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 699 2068 763 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 699 1982 763 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 699 1982 763 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 699 1896 763 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 699 1896 763 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 699 1810 763 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 699 1810 763 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 699 1724 763 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 699 1724 763 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 699 1638 763 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 699 1638 763 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 699 1552 763 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 699 1552 763 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 699 1466 763 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 699 1466 763 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 699 1380 763 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 699 1380 763 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 618 2240 682 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 618 2240 682 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 618 2154 682 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 618 2154 682 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 618 2068 682 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 618 2068 682 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 618 1982 682 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 618 1982 682 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 618 1896 682 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 618 1896 682 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 618 1810 682 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 618 1810 682 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 618 1724 682 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 618 1724 682 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 618 1638 682 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 618 1638 682 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 618 1552 682 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 618 1552 682 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 618 1466 682 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 618 1466 682 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 618 1380 682 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 618 1380 682 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 536 2240 600 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 536 2240 600 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 536 2154 600 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 536 2154 600 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 536 2068 600 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 536 2068 600 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 536 1982 600 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 536 1982 600 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 536 1896 600 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 536 1896 600 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 536 1810 600 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 536 1810 600 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 536 1724 600 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 536 1724 600 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 536 1638 600 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 536 1638 600 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 536 1552 600 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 536 1552 600 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 536 1466 600 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 536 1466 600 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 536 1380 600 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 536 1380 600 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 454 2240 518 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 454 2240 518 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 454 2154 518 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 454 2154 518 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 454 2068 518 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 454 2068 518 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 454 1982 518 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 454 1982 518 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 454 1896 518 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 454 1896 518 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 454 1810 518 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 454 1810 518 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 454 1724 518 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 454 1724 518 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 454 1638 518 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 454 1638 518 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 454 1552 518 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 454 1552 518 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 454 1466 518 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 454 1466 518 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 454 1380 518 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 454 1380 518 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 372 2240 436 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 372 2240 436 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 372 2154 436 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 372 2154 436 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 372 2068 436 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 372 2068 436 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 372 1982 436 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 372 1982 436 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 372 1896 436 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 372 1896 436 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 372 1810 436 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 372 1810 436 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 372 1724 436 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 372 1724 436 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 372 1638 436 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 372 1638 436 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 372 1552 436 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 372 1552 436 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 372 1466 436 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 372 1466 436 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 372 1380 436 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 372 1380 436 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 290 2240 354 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 290 2240 354 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 290 2154 354 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 290 2154 354 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 290 2068 354 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 290 2068 354 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 290 1982 354 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 290 1982 354 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 290 1896 354 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 290 1896 354 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 290 1810 354 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 290 1810 354 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 290 1724 354 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 290 1724 354 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 290 1638 354 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 290 1638 354 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 290 1552 354 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 290 1552 354 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 290 1466 354 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 290 1466 354 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 290 1380 354 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 290 1380 354 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 254 2240 272 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 208 2240 272 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 254 2154 272 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 208 2154 272 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 254 2068 272 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 208 2068 272 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 254 1982 272 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 208 1982 272 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 254 1896 272 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 208 1896 272 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 254 1810 272 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 208 1810 272 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 254 1724 272 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 208 1724 272 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 254 1638 272 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 208 1638 272 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 254 1552 272 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 208 1552 272 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 254 1466 272 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 208 1466 272 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal4 s 254 1380 272 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 208 1380 272 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 126 2240 190 2304 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 126 2154 190 2218 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 126 2068 190 2132 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 126 1982 190 2046 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 126 1896 190 1960 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 126 1810 190 1874 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 126 1724 190 1788 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 126 1638 190 1702 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 126 1552 190 1616 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 126 1466 190 1530 6 VCCD
port 5 nsew power bidirectional
rlabel metal3 s 126 1380 190 1444 6 VCCD
port 5 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 6 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 6 VDDA
port 6 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 VDDA
port 6 nsew power bidirectional
rlabel metal4 s 0 2587 193 3277 6 VDDA
port 6 nsew power bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 0 11247 254 12137 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal4 s 0 5977 254 6667 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal4 s 0 34757 254 39600 6 VSSIO
port 9 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 10 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 6 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 0 7917 254 8847 6 VSSD
port 10 nsew ground bidirectional
rlabel metal4 s 0 10225 15000 10821 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 0 9273 15000 9869 6 AMUXBUS_B
port 12 nsew signal bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 39600
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 538092
string GDS_START 446284
<< end >>
