magic
tech sky130A
magscale 1 2
timestamp 1651250933
<< nwell >>
rect -84 832 972 1575
<< nmos >>
rect 155 324 185 377
tri 185 324 201 340 sw
rect 155 294 261 324
tri 261 294 291 324 sw
rect 155 193 185 294
tri 185 278 201 294 nw
tri 245 278 261 294 ne
tri 185 193 201 209 sw
tri 245 193 261 209 se
rect 261 193 291 294
tri 155 163 185 193 ne
rect 185 163 261 193
tri 261 163 291 193 nw
rect 599 324 629 377
tri 629 324 645 340 sw
rect 599 294 705 324
tri 705 294 735 324 sw
rect 599 193 629 294
tri 629 278 645 294 nw
tri 689 278 705 294 ne
tri 629 193 645 209 sw
tri 689 193 705 209 se
rect 705 193 735 294
tri 599 163 629 193 ne
rect 629 163 705 193
tri 705 163 735 193 nw
<< pmos >>
rect 163 1050 193 1450
rect 251 1050 281 1450
rect 607 1050 637 1450
rect 695 1050 725 1450
<< ndiff >>
rect 99 361 155 377
rect 99 327 109 361
rect 143 327 155 361
rect 99 289 155 327
rect 185 361 345 377
rect 185 340 303 361
tri 185 324 201 340 ne
rect 201 327 303 340
rect 337 327 345 361
rect 201 324 345 327
tri 261 294 291 324 ne
rect 99 255 109 289
rect 143 255 155 289
rect 99 221 155 255
rect 99 187 109 221
rect 143 187 155 221
tri 185 278 201 294 se
rect 201 278 245 294
tri 245 278 261 294 sw
rect 185 245 261 278
rect 185 211 205 245
rect 239 211 261 245
rect 185 209 261 211
tri 185 193 201 209 ne
rect 201 193 245 209
tri 245 193 261 209 nw
rect 291 289 345 324
rect 291 255 303 289
rect 337 255 345 289
rect 291 221 345 255
rect 99 163 155 187
tri 155 163 185 193 sw
tri 261 163 291 193 se
rect 291 187 303 221
rect 337 187 345 221
rect 291 163 345 187
rect 99 151 345 163
rect 99 117 109 151
rect 143 117 205 151
rect 239 117 303 151
rect 337 117 345 151
rect 99 101 345 117
rect 543 361 599 377
rect 543 327 553 361
rect 587 327 599 361
rect 543 289 599 327
rect 629 361 789 377
rect 629 340 747 361
tri 629 324 645 340 ne
rect 645 327 747 340
rect 781 327 789 361
rect 645 324 789 327
tri 705 294 735 324 ne
rect 543 255 553 289
rect 587 255 599 289
rect 543 221 599 255
rect 543 187 553 221
rect 587 187 599 221
tri 629 278 645 294 se
rect 645 278 689 294
tri 689 278 705 294 sw
rect 629 245 705 278
rect 629 211 649 245
rect 683 211 705 245
rect 629 209 705 211
tri 629 193 645 209 ne
rect 645 193 689 209
tri 689 193 705 209 nw
rect 735 289 789 324
rect 735 255 747 289
rect 781 255 789 289
rect 735 221 789 255
rect 543 163 599 187
tri 599 163 629 193 sw
tri 705 163 735 193 se
rect 735 187 747 221
rect 781 187 789 221
rect 735 163 789 187
rect 543 151 789 163
rect 543 117 553 151
rect 587 117 649 151
rect 683 117 747 151
rect 781 117 789 151
rect 543 101 789 117
<< pdiff >>
rect 107 1412 163 1450
rect 107 1378 117 1412
rect 151 1378 163 1412
rect 107 1344 163 1378
rect 107 1310 117 1344
rect 151 1310 163 1344
rect 107 1276 163 1310
rect 107 1242 117 1276
rect 151 1242 163 1276
rect 107 1208 163 1242
rect 107 1174 117 1208
rect 151 1174 163 1208
rect 107 1139 163 1174
rect 107 1105 117 1139
rect 151 1105 163 1139
rect 107 1050 163 1105
rect 193 1412 251 1450
rect 193 1378 205 1412
rect 239 1378 251 1412
rect 193 1344 251 1378
rect 193 1310 205 1344
rect 239 1310 251 1344
rect 193 1276 251 1310
rect 193 1242 205 1276
rect 239 1242 251 1276
rect 193 1208 251 1242
rect 193 1174 205 1208
rect 239 1174 251 1208
rect 193 1139 251 1174
rect 193 1105 205 1139
rect 239 1105 251 1139
rect 193 1050 251 1105
rect 281 1412 335 1450
rect 281 1378 293 1412
rect 327 1378 335 1412
rect 281 1344 335 1378
rect 281 1310 293 1344
rect 327 1310 335 1344
rect 281 1276 335 1310
rect 281 1242 293 1276
rect 327 1242 335 1276
rect 281 1208 335 1242
rect 281 1174 293 1208
rect 327 1174 335 1208
rect 281 1139 335 1174
rect 281 1105 293 1139
rect 327 1105 335 1139
rect 281 1050 335 1105
rect 551 1412 607 1450
rect 551 1378 561 1412
rect 595 1378 607 1412
rect 551 1344 607 1378
rect 551 1310 561 1344
rect 595 1310 607 1344
rect 551 1276 607 1310
rect 551 1242 561 1276
rect 595 1242 607 1276
rect 551 1208 607 1242
rect 551 1174 561 1208
rect 595 1174 607 1208
rect 551 1139 607 1174
rect 551 1105 561 1139
rect 595 1105 607 1139
rect 551 1050 607 1105
rect 637 1412 695 1450
rect 637 1378 649 1412
rect 683 1378 695 1412
rect 637 1344 695 1378
rect 637 1310 649 1344
rect 683 1310 695 1344
rect 637 1276 695 1310
rect 637 1242 649 1276
rect 683 1242 695 1276
rect 637 1208 695 1242
rect 637 1174 649 1208
rect 683 1174 695 1208
rect 637 1139 695 1174
rect 637 1105 649 1139
rect 683 1105 695 1139
rect 637 1050 695 1105
rect 725 1412 779 1450
rect 725 1378 737 1412
rect 771 1378 779 1412
rect 725 1344 779 1378
rect 725 1310 737 1344
rect 771 1310 779 1344
rect 725 1276 779 1310
rect 725 1242 737 1276
rect 771 1242 779 1276
rect 725 1208 779 1242
rect 725 1174 737 1208
rect 771 1174 779 1208
rect 725 1139 779 1174
rect 725 1105 737 1139
rect 771 1105 779 1139
rect 725 1050 779 1105
<< ndiffc >>
rect 109 327 143 361
rect 303 327 337 361
rect 109 255 143 289
rect 109 187 143 221
rect 205 211 239 245
rect 303 255 337 289
rect 303 187 337 221
rect 109 117 143 151
rect 205 117 239 151
rect 303 117 337 151
rect 553 327 587 361
rect 747 327 781 361
rect 553 255 587 289
rect 553 187 587 221
rect 649 211 683 245
rect 747 255 781 289
rect 747 187 781 221
rect 553 117 587 151
rect 649 117 683 151
rect 747 117 781 151
<< pdiffc >>
rect 117 1378 151 1412
rect 117 1310 151 1344
rect 117 1242 151 1276
rect 117 1174 151 1208
rect 117 1105 151 1139
rect 205 1378 239 1412
rect 205 1310 239 1344
rect 205 1242 239 1276
rect 205 1174 239 1208
rect 205 1105 239 1139
rect 293 1378 327 1412
rect 293 1310 327 1344
rect 293 1242 327 1276
rect 293 1174 327 1208
rect 293 1105 327 1139
rect 561 1378 595 1412
rect 561 1310 595 1344
rect 561 1242 595 1276
rect 561 1174 595 1208
rect 561 1105 595 1139
rect 649 1378 683 1412
rect 649 1310 683 1344
rect 649 1242 683 1276
rect 649 1174 683 1208
rect 649 1105 683 1139
rect 737 1378 771 1412
rect 737 1310 771 1344
rect 737 1242 771 1276
rect 737 1174 771 1208
rect 737 1105 771 1139
<< psubdiff >>
rect -31 546 919 572
rect -31 512 -17 546
rect 17 512 427 546
rect 461 512 871 546
rect 905 512 919 546
rect -31 510 919 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 413 474 475 510
rect -31 368 -17 402
rect 17 368 31 402
rect 413 440 427 474
rect 461 440 475 474
rect 413 402 475 440
rect 857 474 919 510
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 413 368 427 402
rect 461 368 475 402
rect 857 440 871 474
rect 905 440 919 474
rect 857 402 919 440
rect 413 330 475 368
rect 413 296 427 330
rect 461 296 475 330
rect 413 258 475 296
rect 413 224 427 258
rect 461 224 475 258
rect 413 186 475 224
rect 413 152 427 186
rect 461 152 475 186
rect 413 114 475 152
rect -31 47 31 80
rect 413 80 427 114
rect 461 80 475 114
rect 857 368 871 402
rect 905 368 919 402
rect 857 330 919 368
rect 857 296 871 330
rect 905 296 919 330
rect 857 258 919 296
rect 857 224 871 258
rect 905 224 919 258
rect 857 186 919 224
rect 857 152 871 186
rect 905 152 919 186
rect 857 114 919 152
rect 413 47 475 80
rect 857 80 871 114
rect 905 80 919 114
rect 857 47 919 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 649 47
rect 683 13 727 47
rect 761 13 799 47
rect 833 13 919 47
rect -31 11 31 13
rect 413 11 475 13
rect 857 11 919 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 649 1539
rect 683 1505 727 1539
rect 761 1505 799 1539
rect 833 1505 919 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 413 1470 475 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 413 1436 427 1470
rect 461 1436 475 1470
rect 857 1470 919 1505
rect 413 1398 475 1436
rect 413 1364 427 1398
rect 461 1364 475 1398
rect 413 1326 475 1364
rect 413 1292 427 1326
rect 461 1292 475 1326
rect 413 1254 475 1292
rect 413 1220 427 1254
rect 461 1220 475 1254
rect 413 1182 475 1220
rect 413 1148 427 1182
rect 461 1148 475 1182
rect 413 1110 475 1148
rect 413 1076 427 1110
rect 461 1076 475 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 413 1038 475 1076
rect 857 1436 871 1470
rect 905 1436 919 1470
rect 857 1398 919 1436
rect 857 1364 871 1398
rect 905 1364 919 1398
rect 857 1326 919 1364
rect 857 1292 871 1326
rect 905 1292 919 1326
rect 857 1254 919 1292
rect 857 1220 871 1254
rect 905 1220 919 1254
rect 857 1182 919 1220
rect 857 1148 871 1182
rect 905 1148 919 1182
rect 857 1110 919 1148
rect 857 1076 871 1110
rect 905 1076 919 1110
rect 413 1004 427 1038
rect 461 1004 475 1038
rect 413 966 475 1004
rect -31 930 31 932
rect 413 932 427 966
rect 461 932 475 966
rect 857 1038 919 1076
rect 857 1004 871 1038
rect 905 1004 919 1038
rect 857 966 919 1004
rect 413 930 475 932
rect 857 932 871 966
rect 905 932 919 966
rect 857 930 919 932
rect -31 868 919 930
<< psubdiffcont >>
rect -17 512 17 546
rect 427 512 461 546
rect 871 512 905 546
rect -17 440 17 474
rect -17 368 17 402
rect 427 440 461 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 427 368 461 402
rect 871 440 905 474
rect 427 296 461 330
rect 427 224 461 258
rect 427 152 461 186
rect 427 80 461 114
rect 871 368 905 402
rect 871 296 905 330
rect 871 224 905 258
rect 871 152 905 186
rect 871 80 905 114
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
rect 499 13 533 47
rect 571 13 605 47
rect 649 13 683 47
rect 727 13 761 47
rect 799 13 833 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 499 1505 533 1539
rect 571 1505 605 1539
rect 649 1505 683 1539
rect 727 1505 761 1539
rect 799 1505 833 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 427 1436 461 1470
rect 427 1364 461 1398
rect 427 1292 461 1326
rect 427 1220 461 1254
rect 427 1148 461 1182
rect 427 1076 461 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 871 1436 905 1470
rect 871 1364 905 1398
rect 871 1292 905 1326
rect 871 1220 905 1254
rect 871 1148 905 1182
rect 871 1076 905 1110
rect 427 1004 461 1038
rect 427 932 461 966
rect 871 1004 905 1038
rect 871 932 905 966
<< poly >>
rect 163 1450 193 1476
rect 251 1450 281 1476
rect 607 1450 637 1476
rect 695 1450 725 1476
rect 163 1019 193 1050
rect 251 1019 281 1050
rect 121 1003 281 1019
rect 121 969 131 1003
rect 165 989 281 1003
rect 607 1019 637 1050
rect 695 1019 725 1050
rect 165 969 175 989
rect 121 953 175 969
rect 565 1003 725 1019
rect 565 969 575 1003
rect 609 989 725 1003
rect 609 969 619 989
rect 565 953 619 969
rect 121 461 175 477
rect 121 427 131 461
rect 165 441 175 461
rect 165 427 185 441
rect 121 411 185 427
rect 155 377 185 411
rect 565 461 619 477
rect 565 427 575 461
rect 609 441 619 461
rect 609 427 629 441
rect 565 411 629 427
rect 599 377 629 411
<< polycont >>
rect 131 969 165 1003
rect 575 969 609 1003
rect 131 427 165 461
rect 575 427 609 461
<< locali >>
rect -31 1539 919 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 649 1539
rect 683 1505 727 1539
rect 761 1505 799 1539
rect 833 1505 919 1539
rect -31 1492 919 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect 117 1412 151 1492
rect 117 1344 151 1378
rect 117 1276 151 1310
rect 117 1208 151 1242
rect 117 1139 151 1174
rect 117 1083 151 1105
rect 205 1412 239 1450
rect 205 1344 239 1378
rect 205 1276 239 1310
rect 205 1208 239 1242
rect 205 1139 239 1174
rect -31 1038 31 1076
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 131 1003 165 1019
rect 131 683 165 969
rect 205 979 239 1105
rect 293 1412 327 1492
rect 293 1344 327 1378
rect 293 1276 327 1310
rect 293 1208 327 1242
rect 293 1139 327 1174
rect 293 1083 327 1105
rect 413 1470 475 1492
rect 413 1436 427 1470
rect 461 1436 475 1470
rect 413 1398 475 1436
rect 413 1364 427 1398
rect 461 1364 475 1398
rect 413 1326 475 1364
rect 413 1292 427 1326
rect 461 1292 475 1326
rect 413 1254 475 1292
rect 413 1220 427 1254
rect 461 1220 475 1254
rect 413 1182 475 1220
rect 413 1148 427 1182
rect 461 1148 475 1182
rect 413 1110 475 1148
rect 413 1076 427 1110
rect 461 1076 475 1110
rect 561 1412 595 1492
rect 561 1344 595 1378
rect 561 1276 595 1310
rect 561 1208 595 1242
rect 561 1139 595 1174
rect 561 1083 595 1105
rect 649 1412 683 1450
rect 649 1344 683 1378
rect 649 1276 683 1310
rect 649 1208 683 1242
rect 649 1139 683 1174
rect 413 1038 475 1076
rect 413 1004 427 1038
rect 461 1004 475 1038
rect 205 945 313 979
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 131 461 165 649
rect 279 535 313 945
rect 413 966 475 1004
rect 413 932 427 966
rect 461 932 475 966
rect 413 868 475 932
rect 575 1003 609 1019
rect 279 461 313 501
rect 131 411 165 427
rect 205 427 313 461
rect 413 546 475 572
rect 413 512 427 546
rect 461 512 475 546
rect 413 474 475 512
rect 413 440 427 474
rect 461 440 475 474
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect -31 62 31 80
rect 109 361 143 377
rect 109 289 143 327
rect 109 221 143 255
rect 205 245 239 427
rect 413 402 475 440
rect 575 535 609 969
rect 649 979 683 1105
rect 737 1412 771 1492
rect 737 1344 771 1378
rect 737 1276 771 1310
rect 737 1208 771 1242
rect 737 1139 771 1174
rect 737 1083 771 1105
rect 857 1470 919 1492
rect 857 1436 871 1470
rect 905 1436 919 1470
rect 857 1398 919 1436
rect 857 1364 871 1398
rect 905 1364 919 1398
rect 857 1326 919 1364
rect 857 1292 871 1326
rect 905 1292 919 1326
rect 857 1254 919 1292
rect 857 1220 871 1254
rect 905 1220 919 1254
rect 857 1182 919 1220
rect 857 1148 871 1182
rect 905 1148 919 1182
rect 857 1110 919 1148
rect 857 1076 871 1110
rect 905 1076 919 1110
rect 857 1038 919 1076
rect 857 1004 871 1038
rect 905 1004 919 1038
rect 649 945 757 979
rect 575 461 609 501
rect 723 683 757 945
rect 857 966 919 1004
rect 857 932 871 966
rect 905 932 919 966
rect 857 868 919 932
rect 723 461 757 649
rect 575 411 609 427
rect 649 427 757 461
rect 857 546 919 572
rect 857 512 871 546
rect 905 512 919 546
rect 857 474 919 512
rect 857 440 871 474
rect 905 440 919 474
rect 205 195 239 211
rect 303 361 337 377
rect 303 289 337 327
rect 303 221 337 255
rect 109 151 143 187
rect 303 151 337 187
rect 143 117 205 151
rect 239 117 303 151
rect 109 62 143 117
rect 206 62 240 117
rect 303 62 337 117
rect 413 368 427 402
rect 461 368 475 402
rect 413 330 475 368
rect 413 296 427 330
rect 461 296 475 330
rect 413 258 475 296
rect 413 224 427 258
rect 461 224 475 258
rect 413 186 475 224
rect 413 152 427 186
rect 461 152 475 186
rect 413 114 475 152
rect 413 80 427 114
rect 461 80 475 114
rect 413 62 475 80
rect 553 361 587 377
rect 553 289 587 327
rect 553 221 587 255
rect 649 245 683 427
rect 857 402 919 440
rect 649 195 683 211
rect 747 361 781 377
rect 747 289 781 327
rect 747 221 781 255
rect 553 151 587 187
rect 747 151 781 187
rect 587 117 649 151
rect 683 117 747 151
rect 553 62 587 117
rect 650 62 684 117
rect 747 62 781 117
rect 857 368 871 402
rect 905 368 919 402
rect 857 330 919 368
rect 857 296 871 330
rect 905 296 919 330
rect 857 258 919 296
rect 857 224 871 258
rect 905 224 919 258
rect 857 186 919 224
rect 857 152 871 186
rect 905 152 919 186
rect 857 114 919 152
rect 857 80 871 114
rect 905 80 919 114
rect 857 62 919 80
rect -31 47 919 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 649 47
rect 683 13 727 47
rect 761 13 799 47
rect 833 13 919 47
rect -31 0 919 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 205 1505 239 1539
rect 283 1505 317 1539
rect 355 1505 389 1539
rect 499 1505 533 1539
rect 571 1505 605 1539
rect 649 1505 683 1539
rect 727 1505 761 1539
rect 799 1505 833 1539
rect 131 649 165 683
rect 279 501 313 535
rect 575 501 609 535
rect 723 649 757 683
rect 55 13 89 47
rect 127 13 161 47
rect 205 13 239 47
rect 283 13 317 47
rect 355 13 389 47
rect 499 13 533 47
rect 571 13 605 47
rect 649 13 683 47
rect 727 13 761 47
rect 799 13 833 47
<< metal1 >>
rect -31 1539 919 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 205 1539
rect 239 1505 283 1539
rect 317 1505 355 1539
rect 389 1505 499 1539
rect 533 1505 571 1539
rect 605 1505 649 1539
rect 683 1505 727 1539
rect 761 1505 799 1539
rect 833 1505 919 1539
rect -31 1492 919 1505
rect 125 683 171 689
rect 717 683 763 689
rect 95 649 131 683
rect 165 649 177 683
rect 711 649 723 683
rect 757 649 793 683
rect 125 643 171 649
rect 717 643 763 649
rect 273 535 319 541
rect 569 535 615 541
rect 267 501 279 535
rect 313 501 575 535
rect 609 501 621 535
rect 273 495 319 501
rect 569 495 615 501
rect -31 47 919 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 205 47
rect 239 13 283 47
rect 317 13 355 47
rect 389 13 499 47
rect 533 13 571 47
rect 605 13 649 47
rect 683 13 727 47
rect 761 13 799 47
rect 833 13 919 47
rect -31 0 919 13
<< labels >>
rlabel metal1 723 649 757 683 1 Y
port 1 n
rlabel metal1 131 649 165 683 1 A
port 2 n
rlabel metal1 -31 1492 919 1554 1 VDD
port 3 n
rlabel metal1 -31 0 919 62 1 GND
port 4 n
<< end >>
