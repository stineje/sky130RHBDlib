// File: AOI3X1.spi.AOI3X1.pxi
// Created: Tue Oct 15 15:45:23 2024
// 
simulator lang=spectre
x_PM_AOI3X1\%GND ( GND N_GND_c_12_p N_GND_c_27_p N_GND_c_2_p N_GND_c_34_p \
 N_GND_c_53_p N_GND_c_4_p N_GND_c_20_p N_GND_c_65_p N_GND_c_69_p N_GND_c_1_p \
 N_GND_c_3_p N_GND_M0_noxref_d N_GND_M2_noxref_s )  PM_AOI3X1\%GND
x_PM_AOI3X1\%VDD ( VDD N_VDD_c_109_p N_VDD_c_91_p N_VDD_c_92_p N_VDD_c_103_p \
 N_VDD_c_87_n N_VDD_c_88_n N_VDD_c_89_n N_VDD_M4_noxref_s N_VDD_M5_noxref_d \
 N_VDD_M7_noxref_d N_VDD_M8_noxref_d )  PM_AOI3X1\%VDD
x_PM_AOI3X1\%noxref_3 ( N_noxref_3_c_161_n N_noxref_3_c_164_n \
 N_noxref_3_c_184_n N_noxref_3_c_187_n N_noxref_3_c_189_n N_noxref_3_c_165_n \
 N_noxref_3_c_245_p N_noxref_3_c_167_n N_noxref_3_c_169_n N_noxref_3_c_233_p \
 N_noxref_3_c_194_n N_noxref_3_M2_noxref_g N_noxref_3_M8_noxref_g \
 N_noxref_3_M9_noxref_g N_noxref_3_c_172_n N_noxref_3_c_265_p \
 N_noxref_3_c_266_p N_noxref_3_c_174_n N_noxref_3_c_176_n N_noxref_3_c_290_p \
 N_noxref_3_c_254_p N_noxref_3_c_177_n N_noxref_3_c_179_n N_noxref_3_c_201_n \
 N_noxref_3_M1_noxref_d N_noxref_3_M4_noxref_d N_noxref_3_M6_noxref_d )  \
 PM_AOI3X1\%noxref_3
x_PM_AOI3X1\%A ( A A A A A A A N_A_c_304_n N_A_M0_noxref_g N_A_M4_noxref_g \
 N_A_M5_noxref_g N_A_c_305_n N_A_c_307_n N_A_c_308_n N_A_c_309_n N_A_c_310_n \
 N_A_c_311_n N_A_c_312_n N_A_c_314_n N_A_c_321_n )  PM_AOI3X1\%A
x_PM_AOI3X1\%B ( B B B B B B B N_B_c_368_n N_B_c_359_n N_B_M1_noxref_g \
 N_B_M6_noxref_g N_B_M7_noxref_g N_B_c_377_n N_B_c_378_n N_B_c_379_n \
 N_B_c_380_n N_B_c_382_n N_B_c_383_n N_B_c_385_n N_B_c_386_n N_B_c_388_n \
 N_B_c_389_n N_B_c_391_n )  PM_AOI3X1\%B
x_PM_AOI3X1\%noxref_6 ( N_noxref_6_c_447_n N_noxref_6_c_423_n \
 N_noxref_6_c_427_n N_noxref_6_c_431_n N_noxref_6_c_432_n N_noxref_6_c_435_n \
 N_noxref_6_M0_noxref_s )  PM_AOI3X1\%noxref_6
x_PM_AOI3X1\%C ( C C C C C C C N_C_c_486_n N_C_c_474_n N_C_M3_noxref_g \
 N_C_M10_noxref_g N_C_M11_noxref_g N_C_c_476_n N_C_c_498_n N_C_c_501_n \
 N_C_c_514_p N_C_c_478_n N_C_c_479_n N_C_c_480_n N_C_c_505_n N_C_c_506_n \
 N_C_c_508_n N_C_c_509_n )  PM_AOI3X1\%C
x_PM_AOI3X1\%YN ( YN YN YN YN YN YN YN YN N_YN_c_543_n N_YN_c_567_n \
 N_YN_c_560_n N_YN_c_561_n N_YN_c_547_n N_YN_M2_noxref_d N_YN_M3_noxref_d \
 N_YN_M10_noxref_d )  PM_AOI3X1\%YN
x_PM_AOI3X1\%noxref_9 ( N_noxref_9_c_609_n N_noxref_9_c_612_n \
 N_noxref_9_c_613_n N_noxref_9_c_614_n N_noxref_9_M8_noxref_s \
 N_noxref_9_M9_noxref_d N_noxref_9_M11_noxref_d )  PM_AOI3X1\%noxref_9
cc_1 ( N_GND_c_1_p N_VDD_c_87_n ) capacitor c=0.00989031f //x=6.29 //y=0 \
 //x2=6.29 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_88_n ) capacitor c=0.00989031f //x=0.74 //y=0 \
 //x2=0.74 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_89_n ) capacitor c=0.00962895f //x=3.33 //y=0 \
 //x2=3.33 //y2=7.4
cc_4 ( N_GND_c_4_p N_noxref_3_c_161_n ) capacitor c=7.22787e-19 //x=4.425 \
 //y=0.53 //x2=4.325 //y2=2.59
cc_5 ( N_GND_c_3_p N_noxref_3_c_161_n ) capacitor c=0.0435449f //x=3.33 //y=0 \
 //x2=4.325 //y2=2.59
cc_6 ( N_GND_M2_noxref_s N_noxref_3_c_161_n ) capacitor c=0.00494344f //x=3.89 \
 //y=0.365 //x2=4.325 //y2=2.59
cc_7 ( N_GND_c_3_p N_noxref_3_c_164_n ) capacitor c=0.00102529f //x=3.33 //y=0 \
 //x2=2.705 //y2=2.59
cc_8 ( N_GND_c_3_p N_noxref_3_c_165_n ) capacitor c=0.0431271f //x=3.33 //y=0 \
 //x2=2.505 //y2=1.655
cc_9 ( N_GND_M2_noxref_s N_noxref_3_c_165_n ) capacitor c=3.00901e-19 //x=3.89 \
 //y=0.365 //x2=2.505 //y2=1.655
cc_10 ( N_GND_c_2_p N_noxref_3_c_167_n ) capacitor c=0.00101801f //x=0.74 \
 //y=0 //x2=2.59 //y2=2.59
cc_11 ( N_GND_c_3_p N_noxref_3_c_167_n ) capacitor c=5.56859e-19 //x=3.33 \
 //y=0 //x2=2.59 //y2=2.59
cc_12 ( N_GND_c_12_p N_noxref_3_c_169_n ) capacitor c=6.7762e-19 //x=6.29 \
 //y=0 //x2=4.44 //y2=2.08
cc_13 ( N_GND_c_4_p N_noxref_3_c_169_n ) capacitor c=0.00133118f //x=4.425 \
 //y=0.53 //x2=4.44 //y2=2.08
cc_14 ( N_GND_c_3_p N_noxref_3_c_169_n ) capacitor c=0.0147015f //x=3.33 //y=0 \
 //x2=4.44 //y2=2.08
cc_15 ( N_GND_c_4_p N_noxref_3_c_172_n ) capacitor c=0.0122561f //x=4.425 \
 //y=0.53 //x2=4.245 //y2=0.905
cc_16 ( N_GND_M2_noxref_s N_noxref_3_c_172_n ) capacitor c=0.0318086f //x=3.89 \
 //y=0.365 //x2=4.245 //y2=0.905
cc_17 ( N_GND_c_4_p N_noxref_3_c_174_n ) capacitor c=2.1838e-19 //x=4.425 \
 //y=0.53 //x2=4.245 //y2=1.915
cc_18 ( N_GND_c_3_p N_noxref_3_c_174_n ) capacitor c=0.0131707f //x=3.33 //y=0 \
 //x2=4.245 //y2=1.915
cc_19 ( N_GND_M2_noxref_s N_noxref_3_c_176_n ) capacitor c=0.00476335f \
 //x=3.89 //y=0.365 //x2=4.62 //y2=0.75
cc_20 ( N_GND_c_20_p N_noxref_3_c_177_n ) capacitor c=0.0113279f //x=4.91 \
 //y=0.53 //x2=4.775 //y2=0.905
cc_21 ( N_GND_M2_noxref_s N_noxref_3_c_177_n ) capacitor c=0.00514143f \
 //x=3.89 //y=0.365 //x2=4.775 //y2=0.905
cc_22 ( N_GND_M2_noxref_s N_noxref_3_c_179_n ) capacitor c=8.33128e-19 \
 //x=3.89 //y=0.365 //x2=4.775 //y2=1.25
cc_23 ( N_GND_c_2_p N_noxref_3_M1_noxref_d ) capacitor c=8.58106e-19 //x=0.74 \
 //y=0 //x2=1.96 //y2=0.905
cc_24 ( N_GND_c_3_p N_noxref_3_M1_noxref_d ) capacitor c=0.00616547f //x=3.33 \
 //y=0 //x2=1.96 //y2=0.905
cc_25 ( N_GND_M0_noxref_d N_noxref_3_M1_noxref_d ) capacitor c=0.00143464f \
 //x=0.99 //y=0.865 //x2=1.96 //y2=0.905
cc_26 ( N_GND_c_2_p N_A_c_304_n ) capacitor c=0.0180518f //x=0.74 //y=0 \
 //x2=1.11 //y2=2.08
cc_27 ( N_GND_c_27_p N_A_c_305_n ) capacitor c=0.00135046f //x=1.095 //y=0 \
 //x2=0.915 //y2=0.865
cc_28 ( N_GND_M0_noxref_d N_A_c_305_n ) capacitor c=0.00220047f //x=0.99 \
 //y=0.865 //x2=0.915 //y2=0.865
cc_29 ( N_GND_M0_noxref_d N_A_c_307_n ) capacitor c=0.00255985f //x=0.99 \
 //y=0.865 //x2=0.915 //y2=1.21
cc_30 ( N_GND_c_2_p N_A_c_308_n ) capacitor c=0.00264481f //x=0.74 //y=0 \
 //x2=0.915 //y2=1.52
cc_31 ( N_GND_c_2_p N_A_c_309_n ) capacitor c=0.0121947f //x=0.74 //y=0 \
 //x2=0.915 //y2=1.915
cc_32 ( N_GND_M0_noxref_d N_A_c_310_n ) capacitor c=0.0131326f //x=0.99 \
 //y=0.865 //x2=1.29 //y2=0.71
cc_33 ( N_GND_M0_noxref_d N_A_c_311_n ) capacitor c=0.00193127f //x=0.99 \
 //y=0.865 //x2=1.29 //y2=1.365
cc_34 ( N_GND_c_34_p N_A_c_312_n ) capacitor c=0.00130622f //x=3.16 //y=0 \
 //x2=1.445 //y2=0.865
cc_35 ( N_GND_M0_noxref_d N_A_c_312_n ) capacitor c=0.00257848f //x=0.99 \
 //y=0.865 //x2=1.445 //y2=0.865
cc_36 ( N_GND_M0_noxref_d N_A_c_314_n ) capacitor c=0.00255985f //x=0.99 \
 //y=0.865 //x2=1.445 //y2=1.21
cc_37 ( N_GND_c_2_p N_B_c_359_n ) capacitor c=9.2064e-19 //x=0.74 //y=0 \
 //x2=1.85 //y2=2.08
cc_38 ( N_GND_c_3_p N_B_c_359_n ) capacitor c=0.00110071f //x=3.33 //y=0 \
 //x2=1.85 //y2=2.08
cc_39 ( N_GND_c_12_p N_noxref_6_c_423_n ) capacitor c=0.00710948f //x=6.29 \
 //y=0 //x2=1.58 //y2=1.58
cc_40 ( N_GND_c_27_p N_noxref_6_c_423_n ) capacitor c=0.00111428f //x=1.095 \
 //y=0 //x2=1.58 //y2=1.58
cc_41 ( N_GND_c_34_p N_noxref_6_c_423_n ) capacitor c=0.00180846f //x=3.16 \
 //y=0 //x2=1.58 //y2=1.58
cc_42 ( N_GND_M0_noxref_d N_noxref_6_c_423_n ) capacitor c=0.0090983f //x=0.99 \
 //y=0.865 //x2=1.58 //y2=1.58
cc_43 ( N_GND_c_12_p N_noxref_6_c_427_n ) capacitor c=0.00723598f //x=6.29 \
 //y=0 //x2=1.665 //y2=0.615
cc_44 ( N_GND_c_34_p N_noxref_6_c_427_n ) capacitor c=0.0146208f //x=3.16 \
 //y=0 //x2=1.665 //y2=0.615
cc_45 ( N_GND_c_1_p N_noxref_6_c_427_n ) capacitor c=0.00145873f //x=6.29 \
 //y=0 //x2=1.665 //y2=0.615
cc_46 ( N_GND_M0_noxref_d N_noxref_6_c_427_n ) capacitor c=0.033812f //x=0.99 \
 //y=0.865 //x2=1.665 //y2=0.615
cc_47 ( N_GND_c_2_p N_noxref_6_c_431_n ) capacitor c=2.91423e-19 //x=0.74 \
 //y=0 //x2=1.665 //y2=1.495
cc_48 ( N_GND_c_12_p N_noxref_6_c_432_n ) capacitor c=0.0199727f //x=6.29 \
 //y=0 //x2=2.55 //y2=0.53
cc_49 ( N_GND_c_34_p N_noxref_6_c_432_n ) capacitor c=0.0371035f //x=3.16 \
 //y=0 //x2=2.55 //y2=0.53
cc_50 ( N_GND_c_1_p N_noxref_6_c_432_n ) capacitor c=0.002964f //x=6.29 //y=0 \
 //x2=2.55 //y2=0.53
cc_51 ( N_GND_c_12_p N_noxref_6_c_435_n ) capacitor c=0.00719615f //x=6.29 \
 //y=0 //x2=2.635 //y2=0.615
cc_52 ( N_GND_c_34_p N_noxref_6_c_435_n ) capacitor c=0.0144264f //x=3.16 \
 //y=0 //x2=2.635 //y2=0.615
cc_53 ( N_GND_c_53_p N_noxref_6_c_435_n ) capacitor c=9.02073e-19 //x=4.025 \
 //y=0.445 //x2=2.635 //y2=0.615
cc_54 ( N_GND_c_1_p N_noxref_6_c_435_n ) capacitor c=0.00145015f //x=6.29 \
 //y=0 //x2=2.635 //y2=0.615
cc_55 ( N_GND_c_3_p N_noxref_6_c_435_n ) capacitor c=0.0431718f //x=3.33 //y=0 \
 //x2=2.635 //y2=0.615
cc_56 ( N_GND_c_12_p N_noxref_6_M0_noxref_s ) capacitor c=0.00723598f //x=6.29 \
 //y=0 //x2=0.56 //y2=0.365
cc_57 ( N_GND_c_27_p N_noxref_6_M0_noxref_s ) capacitor c=0.0146208f //x=1.095 \
 //y=0 //x2=0.56 //y2=0.365
cc_58 ( N_GND_c_2_p N_noxref_6_M0_noxref_s ) capacitor c=0.0594057f //x=0.74 \
 //y=0 //x2=0.56 //y2=0.365
cc_59 ( N_GND_c_1_p N_noxref_6_M0_noxref_s ) capacitor c=0.00145873f //x=6.29 \
 //y=0 //x2=0.56 //y2=0.365
cc_60 ( N_GND_c_3_p N_noxref_6_M0_noxref_s ) capacitor c=0.00198043f //x=3.33 \
 //y=0 //x2=0.56 //y2=0.365
cc_61 ( N_GND_M0_noxref_d N_noxref_6_M0_noxref_s ) capacitor c=0.0334197f \
 //x=0.99 //y=0.865 //x2=0.56 //y2=0.365
cc_62 ( N_GND_M2_noxref_s N_noxref_6_M0_noxref_s ) capacitor c=9.02073e-19 \
 //x=3.89 //y=0.365 //x2=0.56 //y2=0.365
cc_63 ( N_GND_c_1_p N_C_c_474_n ) capacitor c=9.53263e-19 //x=6.29 //y=0 \
 //x2=5.18 //y2=2.08
cc_64 ( N_GND_c_3_p N_C_c_474_n ) capacitor c=0.00112835f //x=3.33 //y=0 \
 //x2=5.18 //y2=2.08
cc_65 ( N_GND_c_65_p N_C_c_476_n ) capacitor c=0.0109802f //x=5.395 //y=0.53 \
 //x2=5.215 //y2=0.905
cc_66 ( N_GND_M2_noxref_s N_C_c_476_n ) capacitor c=0.00590563f //x=3.89 \
 //y=0.365 //x2=5.215 //y2=0.905
cc_67 ( N_GND_M2_noxref_s N_C_c_478_n ) capacitor c=0.00466751f //x=3.89 \
 //y=0.365 //x2=5.59 //y2=0.75
cc_68 ( N_GND_M2_noxref_s N_C_c_479_n ) capacitor c=0.00316186f //x=3.89 \
 //y=0.365 //x2=5.59 //y2=1.405
cc_69 ( N_GND_c_69_p N_C_c_480_n ) capacitor c=0.0112321f //x=5.88 //y=0.53 \
 //x2=5.745 //y2=0.905
cc_70 ( N_GND_M2_noxref_s N_C_c_480_n ) capacitor c=0.0142835f //x=3.89 \
 //y=0.365 //x2=5.745 //y2=0.905
cc_71 ( N_GND_c_3_p YN ) capacitor c=9.64732e-19 //x=3.33 //y=0 //x2=5.92 \
 //y2=2.22
cc_72 ( N_GND_c_12_p N_YN_c_543_n ) capacitor c=0.00359057f //x=6.29 //y=0 \
 //x2=5.395 //y2=1.655
cc_73 ( N_GND_c_20_p N_YN_c_543_n ) capacitor c=0.00381844f //x=4.91 //y=0.53 \
 //x2=5.395 //y2=1.655
cc_74 ( N_GND_c_65_p N_YN_c_543_n ) capacitor c=0.00323369f //x=5.395 //y=0.53 \
 //x2=5.395 //y2=1.655
cc_75 ( N_GND_M2_noxref_s N_YN_c_543_n ) capacitor c=0.0173679f //x=3.89 \
 //y=0.365 //x2=5.395 //y2=1.655
cc_76 ( N_GND_c_12_p N_YN_c_547_n ) capacitor c=0.00295442f //x=6.29 //y=0 \
 //x2=5.835 //y2=1.655
cc_77 ( N_GND_c_69_p N_YN_c_547_n ) capacitor c=0.0047981f //x=5.88 //y=0.53 \
 //x2=5.835 //y2=1.655
cc_78 ( N_GND_c_1_p N_YN_c_547_n ) capacitor c=0.0471746f //x=6.29 //y=0 \
 //x2=5.835 //y2=1.655
cc_79 ( N_GND_M2_noxref_s N_YN_c_547_n ) capacitor c=0.016186f //x=3.89 \
 //y=0.365 //x2=5.835 //y2=1.655
cc_80 ( N_GND_c_12_p N_YN_M2_noxref_d ) capacitor c=0.00175924f //x=6.29 //y=0 \
 //x2=4.32 //y2=0.905
cc_81 ( N_GND_c_1_p N_YN_M2_noxref_d ) capacitor c=4.88559e-19 //x=6.29 //y=0 \
 //x2=4.32 //y2=0.905
cc_82 ( N_GND_c_3_p N_YN_M2_noxref_d ) capacitor c=0.00416273f //x=3.33 //y=0 \
 //x2=4.32 //y2=0.905
cc_83 ( N_GND_M2_noxref_s N_YN_M2_noxref_d ) capacitor c=0.0769466f //x=3.89 \
 //y=0.365 //x2=4.32 //y2=0.905
cc_84 ( N_GND_c_12_p N_YN_M3_noxref_d ) capacitor c=0.00195394f //x=6.29 //y=0 \
 //x2=5.29 //y2=0.905
cc_85 ( N_GND_c_1_p N_YN_M3_noxref_d ) capacitor c=0.00634044f //x=6.29 //y=0 \
 //x2=5.29 //y2=0.905
cc_86 ( N_GND_M2_noxref_s N_YN_M3_noxref_d ) capacitor c=0.0610175f //x=3.89 \
 //y=0.365 //x2=5.29 //y2=0.905
cc_87 ( N_VDD_c_89_n N_noxref_3_c_161_n ) capacitor c=0.00382812f //x=3.33 \
 //y=7.4 //x2=4.325 //y2=2.59
cc_88 ( N_VDD_c_91_p N_noxref_3_c_184_n ) capacitor c=5.76712e-19 //x=1.585 \
 //y=7.4 //x2=2.025 //y2=5.2
cc_89 ( N_VDD_c_92_p N_noxref_3_c_184_n ) capacitor c=5.76712e-19 //x=2.465 \
 //y=7.4 //x2=2.025 //y2=5.2
cc_90 ( N_VDD_M5_noxref_d N_noxref_3_c_184_n ) capacitor c=0.0132775f \
 //x=1.525 //y=5.02 //x2=2.025 //y2=5.2
cc_91 ( N_VDD_c_88_n N_noxref_3_c_187_n ) capacitor c=0.00989999f //x=0.74 \
 //y=7.4 //x2=1.315 //y2=5.2
cc_92 ( N_VDD_M4_noxref_s N_noxref_3_c_187_n ) capacitor c=0.087833f //x=0.655 \
 //y=5.02 //x2=1.315 //y2=5.2
cc_93 ( N_VDD_c_92_p N_noxref_3_c_189_n ) capacitor c=8.71806e-19 //x=2.465 \
 //y=7.4 //x2=2.505 //y2=5.2
cc_94 ( N_VDD_M7_noxref_d N_noxref_3_c_189_n ) capacitor c=0.0167784f \
 //x=2.405 //y=5.02 //x2=2.505 //y2=5.2
cc_95 ( N_VDD_c_88_n N_noxref_3_c_167_n ) capacitor c=0.00159771f //x=0.74 \
 //y=7.4 //x2=2.59 //y2=2.59
cc_96 ( N_VDD_c_89_n N_noxref_3_c_167_n ) capacitor c=0.0462672f //x=3.33 \
 //y=7.4 //x2=2.59 //y2=2.59
cc_97 ( N_VDD_c_89_n N_noxref_3_c_169_n ) capacitor c=0.0103855f //x=3.33 \
 //y=7.4 //x2=4.44 //y2=2.08
cc_98 ( N_VDD_c_89_n N_noxref_3_c_194_n ) capacitor c=0.00860173f //x=3.33 \
 //y=7.4 //x2=4.285 //y2=4.705
cc_99 ( N_VDD_M8_noxref_d N_noxref_3_c_194_n ) capacitor c=2.85008e-19 \
 //x=4.415 //y=5.025 //x2=4.285 //y2=4.705
cc_100 ( N_VDD_c_103_p N_noxref_3_M8_noxref_g ) capacitor c=0.0067918f \
 //x=4.475 //y=7.4 //x2=4.34 //y2=6.025
cc_101 ( N_VDD_c_89_n N_noxref_3_M8_noxref_g ) capacitor c=0.0105272f //x=3.33 \
 //y=7.4 //x2=4.34 //y2=6.025
cc_102 ( N_VDD_M8_noxref_d N_noxref_3_M8_noxref_g ) capacitor c=0.0156786f \
 //x=4.415 //y=5.025 //x2=4.34 //y2=6.025
cc_103 ( N_VDD_c_87_n N_noxref_3_M9_noxref_g ) capacitor c=0.00678153f \
 //x=6.29 //y=7.4 //x2=4.78 //y2=6.025
cc_104 ( N_VDD_M8_noxref_d N_noxref_3_M9_noxref_g ) capacitor c=0.0183011f \
 //x=4.415 //y=5.025 //x2=4.78 //y2=6.025
cc_105 ( N_VDD_c_89_n N_noxref_3_c_201_n ) capacitor c=0.00890932f //x=3.33 \
 //y=7.4 //x2=4.285 //y2=4.705
cc_106 ( N_VDD_c_109_p N_noxref_3_M4_noxref_d ) capacitor c=0.00719513f \
 //x=6.29 //y=7.4 //x2=1.085 //y2=5.02
cc_107 ( N_VDD_c_91_p N_noxref_3_M4_noxref_d ) capacitor c=0.0138103f \
 //x=1.585 //y=7.4 //x2=1.085 //y2=5.02
cc_108 ( N_VDD_c_87_n N_noxref_3_M4_noxref_d ) capacitor c=0.00135231f \
 //x=6.29 //y=7.4 //x2=1.085 //y2=5.02
cc_109 ( N_VDD_c_89_n N_noxref_3_M4_noxref_d ) capacitor c=6.94454e-19 \
 //x=3.33 //y=7.4 //x2=1.085 //y2=5.02
cc_110 ( N_VDD_M5_noxref_d N_noxref_3_M4_noxref_d ) capacitor c=0.0664752f \
 //x=1.525 //y=5.02 //x2=1.085 //y2=5.02
cc_111 ( N_VDD_c_109_p N_noxref_3_M6_noxref_d ) capacitor c=0.00719513f \
 //x=6.29 //y=7.4 //x2=1.965 //y2=5.02
cc_112 ( N_VDD_c_92_p N_noxref_3_M6_noxref_d ) capacitor c=0.0138379f \
 //x=2.465 //y=7.4 //x2=1.965 //y2=5.02
cc_113 ( N_VDD_c_87_n N_noxref_3_M6_noxref_d ) capacitor c=0.00135231f \
 //x=6.29 //y=7.4 //x2=1.965 //y2=5.02
cc_114 ( N_VDD_c_89_n N_noxref_3_M6_noxref_d ) capacitor c=0.0120541f //x=3.33 \
 //y=7.4 //x2=1.965 //y2=5.02
cc_115 ( N_VDD_M4_noxref_s N_noxref_3_M6_noxref_d ) capacitor c=0.00111971f \
 //x=0.655 //y=5.02 //x2=1.965 //y2=5.02
cc_116 ( N_VDD_M5_noxref_d N_noxref_3_M6_noxref_d ) capacitor c=0.0664752f \
 //x=1.525 //y=5.02 //x2=1.965 //y2=5.02
cc_117 ( N_VDD_M7_noxref_d N_noxref_3_M6_noxref_d ) capacitor c=0.0664752f \
 //x=2.405 //y=5.02 //x2=1.965 //y2=5.02
cc_118 ( N_VDD_c_91_p N_A_c_304_n ) capacitor c=3.97183e-19 //x=1.585 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_119 ( N_VDD_c_88_n N_A_c_304_n ) capacitor c=0.016845f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_120 ( N_VDD_c_91_p N_A_M4_noxref_g ) capacitor c=0.00726866f //x=1.585 \
 //y=7.4 //x2=1.01 //y2=6.02
cc_121 ( N_VDD_M4_noxref_s N_A_M4_noxref_g ) capacitor c=0.054195f //x=0.655 \
 //y=5.02 //x2=1.01 //y2=6.02
cc_122 ( N_VDD_c_91_p N_A_M5_noxref_g ) capacitor c=0.00672952f //x=1.585 \
 //y=7.4 //x2=1.45 //y2=6.02
cc_123 ( N_VDD_M5_noxref_d N_A_M5_noxref_g ) capacitor c=0.015318f //x=1.525 \
 //y=5.02 //x2=1.45 //y2=6.02
cc_124 ( N_VDD_c_88_n N_A_c_321_n ) capacitor c=0.0292267f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=4.7
cc_125 ( N_VDD_c_88_n N_B_c_359_n ) capacitor c=6.61004e-19 //x=0.74 //y=7.4 \
 //x2=1.85 //y2=2.08
cc_126 ( N_VDD_c_89_n N_B_c_359_n ) capacitor c=6.09526e-19 //x=3.33 //y=7.4 \
 //x2=1.85 //y2=2.08
cc_127 ( N_VDD_c_92_p N_B_M6_noxref_g ) capacitor c=0.00673971f //x=2.465 \
 //y=7.4 //x2=1.89 //y2=6.02
cc_128 ( N_VDD_M5_noxref_d N_B_M6_noxref_g ) capacitor c=0.015318f //x=1.525 \
 //y=5.02 //x2=1.89 //y2=6.02
cc_129 ( N_VDD_c_92_p N_B_M7_noxref_g ) capacitor c=0.00672952f //x=2.465 \
 //y=7.4 //x2=2.33 //y2=6.02
cc_130 ( N_VDD_c_89_n N_B_M7_noxref_g ) capacitor c=0.00954586f //x=3.33 \
 //y=7.4 //x2=2.33 //y2=6.02
cc_131 ( N_VDD_M7_noxref_d N_B_M7_noxref_g ) capacitor c=0.0430452f //x=2.405 \
 //y=5.02 //x2=2.33 //y2=6.02
cc_132 ( N_VDD_c_87_n N_C_c_474_n ) capacitor c=6.16704e-19 //x=6.29 //y=7.4 \
 //x2=5.18 //y2=2.08
cc_133 ( N_VDD_c_89_n N_C_c_474_n ) capacitor c=7.02327e-19 //x=3.33 //y=7.4 \
 //x2=5.18 //y2=2.08
cc_134 ( N_VDD_c_87_n N_C_M10_noxref_g ) capacitor c=0.00513565f //x=6.29 \
 //y=7.4 //x2=5.22 //y2=6.025
cc_135 ( N_VDD_c_87_n N_C_M11_noxref_g ) capacitor c=0.0322288f //x=6.29 \
 //y=7.4 //x2=5.66 //y2=6.025
cc_136 ( N_VDD_c_87_n YN ) capacitor c=0.0469841f //x=6.29 //y=7.4 //x2=5.92 \
 //y2=2.22
cc_137 ( N_VDD_c_89_n YN ) capacitor c=0.00155409f //x=3.33 //y=7.4 //x2=5.92 \
 //y2=2.22
cc_138 ( N_VDD_c_87_n N_YN_c_560_n ) capacitor c=9.65117e-19 //x=6.29 //y=7.4 \
 //x2=5.835 //y2=5.21
cc_139 ( N_VDD_c_89_n N_YN_c_561_n ) capacitor c=8.9933e-19 //x=3.33 //y=7.4 \
 //x2=5.525 //y2=5.21
cc_140 ( N_VDD_c_87_n N_YN_M10_noxref_d ) capacitor c=0.00991513f //x=6.29 \
 //y=7.4 //x2=5.295 //y2=5.025
cc_141 ( N_VDD_M8_noxref_d N_YN_M10_noxref_d ) capacitor c=0.00561178f \
 //x=4.415 //y=5.025 //x2=5.295 //y2=5.025
cc_142 ( N_VDD_c_103_p N_noxref_9_c_609_n ) capacitor c=5.81484e-19 //x=4.475 \
 //y=7.4 //x2=4.915 //y2=5.21
cc_143 ( N_VDD_c_87_n N_noxref_9_c_609_n ) capacitor c=0.0034744f //x=6.29 \
 //y=7.4 //x2=4.915 //y2=5.21
cc_144 ( N_VDD_M8_noxref_d N_noxref_9_c_609_n ) capacitor c=0.0132432f \
 //x=4.415 //y=5.025 //x2=4.915 //y2=5.21
cc_145 ( N_VDD_c_89_n N_noxref_9_c_612_n ) capacitor c=0.0669114f //x=3.33 \
 //y=7.4 //x2=4.205 //y2=5.21
cc_146 ( N_VDD_c_87_n N_noxref_9_c_613_n ) capacitor c=0.00358752f //x=6.29 \
 //y=7.4 //x2=5.795 //y2=6.91
cc_147 ( N_VDD_c_109_p N_noxref_9_c_614_n ) capacitor c=0.0370274f //x=6.29 \
 //y=7.4 //x2=5.085 //y2=6.91
cc_148 ( N_VDD_c_87_n N_noxref_9_c_614_n ) capacitor c=0.059856f //x=6.29 \
 //y=7.4 //x2=5.085 //y2=6.91
cc_149 ( N_VDD_c_109_p N_noxref_9_M8_noxref_s ) capacitor c=0.00726388f \
 //x=6.29 //y=7.4 //x2=3.985 //y2=5.025
cc_150 ( N_VDD_c_103_p N_noxref_9_M8_noxref_s ) capacitor c=0.0141117f \
 //x=4.475 //y=7.4 //x2=3.985 //y2=5.025
cc_151 ( N_VDD_c_87_n N_noxref_9_M8_noxref_s ) capacitor c=0.00138926f \
 //x=6.29 //y=7.4 //x2=3.985 //y2=5.025
cc_152 ( N_VDD_M7_noxref_d N_noxref_9_M8_noxref_s ) capacitor c=0.00196306f \
 //x=2.405 //y=5.02 //x2=3.985 //y2=5.025
cc_153 ( N_VDD_M8_noxref_d N_noxref_9_M8_noxref_s ) capacitor c=0.0667021f \
 //x=4.415 //y=5.025 //x2=3.985 //y2=5.025
cc_154 ( N_VDD_c_89_n N_noxref_9_M9_noxref_d ) capacitor c=8.88629e-19 \
 //x=3.33 //y=7.4 //x2=4.855 //y2=5.025
cc_155 ( N_VDD_M8_noxref_d N_noxref_9_M9_noxref_d ) capacitor c=0.0659925f \
 //x=4.415 //y=5.025 //x2=4.855 //y2=5.025
cc_156 ( N_VDD_c_87_n N_noxref_9_M11_noxref_d ) capacitor c=0.0528345f \
 //x=6.29 //y=7.4 //x2=5.735 //y2=5.025
cc_157 ( N_VDD_M8_noxref_d N_noxref_9_M11_noxref_d ) capacitor c=0.00107819f \
 //x=4.415 //y=5.025 //x2=5.735 //y2=5.025
cc_158 ( N_noxref_3_c_187_n N_A_c_304_n ) capacitor c=0.0055959f //x=1.315 \
 //y=5.2 //x2=1.11 //y2=2.08
cc_159 ( N_noxref_3_c_167_n N_A_c_304_n ) capacitor c=0.00407922f //x=2.59 \
 //y=2.59 //x2=1.11 //y2=2.08
cc_160 ( N_noxref_3_c_187_n N_A_M4_noxref_g ) capacitor c=0.0177326f //x=1.315 \
 //y=5.2 //x2=1.01 //y2=6.02
cc_161 ( N_noxref_3_c_184_n N_A_M5_noxref_g ) capacitor c=0.0204115f //x=2.025 \
 //y=5.2 //x2=1.45 //y2=6.02
cc_162 ( N_noxref_3_M4_noxref_d N_A_M5_noxref_g ) capacitor c=0.0173476f \
 //x=1.085 //y=5.02 //x2=1.45 //y2=6.02
cc_163 ( N_noxref_3_c_187_n N_A_c_321_n ) capacitor c=0.00605692f //x=1.315 \
 //y=5.2 //x2=1.11 //y2=4.7
cc_164 ( N_noxref_3_c_184_n N_B_c_368_n ) capacitor c=0.0127867f //x=2.025 \
 //y=5.2 //x2=1.85 //y2=4.535
cc_165 ( N_noxref_3_c_167_n N_B_c_368_n ) capacitor c=0.0101284f //x=2.59 \
 //y=2.59 //x2=1.85 //y2=4.535
cc_166 ( N_noxref_3_c_164_n N_B_c_359_n ) capacitor c=0.00732168f //x=2.705 \
 //y=2.59 //x2=1.85 //y2=2.08
cc_167 ( N_noxref_3_c_167_n N_B_c_359_n ) capacitor c=0.0813981f //x=2.59 \
 //y=2.59 //x2=1.85 //y2=2.08
cc_168 ( N_noxref_3_c_169_n N_B_c_359_n ) capacitor c=9.8819e-19 //x=4.44 \
 //y=2.08 //x2=1.85 //y2=2.08
cc_169 ( N_noxref_3_c_184_n N_B_M6_noxref_g ) capacitor c=0.0166699f //x=2.025 \
 //y=5.2 //x2=1.89 //y2=6.02
cc_170 ( N_noxref_3_M6_noxref_d N_B_M6_noxref_g ) capacitor c=0.0173477f \
 //x=1.965 //y=5.02 //x2=1.89 //y2=6.02
cc_171 ( N_noxref_3_c_189_n N_B_M7_noxref_g ) capacitor c=0.0223814f //x=2.505 \
 //y=5.2 //x2=2.33 //y2=6.02
cc_172 ( N_noxref_3_M6_noxref_d N_B_M7_noxref_g ) capacitor c=0.0179769f \
 //x=1.965 //y=5.02 //x2=2.33 //y2=6.02
cc_173 ( N_noxref_3_M1_noxref_d N_B_c_377_n ) capacitor c=0.00217566f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=0.905
cc_174 ( N_noxref_3_M1_noxref_d N_B_c_378_n ) capacitor c=0.0034598f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=1.25
cc_175 ( N_noxref_3_M1_noxref_d N_B_c_379_n ) capacitor c=0.0065582f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=1.56
cc_176 ( N_noxref_3_c_167_n N_B_c_380_n ) capacitor c=0.0142673f //x=2.59 \
 //y=2.59 //x2=2.255 //y2=4.79
cc_177 ( N_noxref_3_c_233_p N_B_c_380_n ) capacitor c=0.00421574f //x=2.11 \
 //y=5.2 //x2=2.255 //y2=4.79
cc_178 ( N_noxref_3_M1_noxref_d N_B_c_382_n ) capacitor c=0.00241102f //x=1.96 \
 //y=0.905 //x2=2.26 //y2=0.75
cc_179 ( N_noxref_3_c_165_n N_B_c_383_n ) capacitor c=0.00359704f //x=2.505 \
 //y=1.655 //x2=2.26 //y2=1.405
cc_180 ( N_noxref_3_M1_noxref_d N_B_c_383_n ) capacitor c=0.0138845f //x=1.96 \
 //y=0.905 //x2=2.26 //y2=1.405
cc_181 ( N_noxref_3_M1_noxref_d N_B_c_385_n ) capacitor c=0.00132245f //x=1.96 \
 //y=0.905 //x2=2.415 //y2=0.905
cc_182 ( N_noxref_3_c_165_n N_B_c_386_n ) capacitor c=0.00457401f //x=2.505 \
 //y=1.655 //x2=2.415 //y2=1.25
cc_183 ( N_noxref_3_M1_noxref_d N_B_c_386_n ) capacitor c=0.00566463f //x=1.96 \
 //y=0.905 //x2=2.415 //y2=1.25
cc_184 ( N_noxref_3_c_167_n N_B_c_388_n ) capacitor c=0.00877984f //x=2.59 \
 //y=2.59 //x2=1.85 //y2=2.08
cc_185 ( N_noxref_3_c_167_n N_B_c_389_n ) capacitor c=0.00306024f //x=2.59 \
 //y=2.59 //x2=1.85 //y2=1.915
cc_186 ( N_noxref_3_M1_noxref_d N_B_c_389_n ) capacitor c=0.00660593f //x=1.96 \
 //y=0.905 //x2=1.85 //y2=1.915
cc_187 ( N_noxref_3_c_184_n N_B_c_391_n ) capacitor c=0.00399417f //x=2.025 \
 //y=5.2 //x2=1.88 //y2=4.7
cc_188 ( N_noxref_3_c_167_n N_B_c_391_n ) capacitor c=0.00533692f //x=2.59 \
 //y=2.59 //x2=1.88 //y2=4.7
cc_189 ( N_noxref_3_c_245_p N_noxref_6_c_447_n ) capacitor c=3.15806e-19 \
 //x=2.235 //y=1.655 //x2=0.695 //y2=1.495
cc_190 ( N_noxref_3_c_245_p N_noxref_6_c_431_n ) capacitor c=0.0201674f \
 //x=2.235 //y=1.655 //x2=1.665 //y2=1.495
cc_191 ( N_noxref_3_c_165_n N_noxref_6_c_432_n ) capacitor c=0.00468333f \
 //x=2.505 //y=1.655 //x2=2.55 //y2=0.53
cc_192 ( N_noxref_3_M1_noxref_d N_noxref_6_c_432_n ) capacitor c=0.0118355f \
 //x=1.96 //y=0.905 //x2=2.55 //y2=0.53
cc_193 ( N_noxref_3_c_161_n N_noxref_6_M0_noxref_s ) capacitor c=3.03583e-19 \
 //x=4.325 //y=2.59 //x2=0.56 //y2=0.365
cc_194 ( N_noxref_3_c_164_n N_noxref_6_M0_noxref_s ) capacitor c=6.92363e-19 \
 //x=2.705 //y=2.59 //x2=0.56 //y2=0.365
cc_195 ( N_noxref_3_c_165_n N_noxref_6_M0_noxref_s ) capacitor c=0.0129465f \
 //x=2.505 //y=1.655 //x2=0.56 //y2=0.365
cc_196 ( N_noxref_3_M1_noxref_d N_noxref_6_M0_noxref_s ) capacitor \
 c=0.0437911f //x=1.96 //y=0.905 //x2=0.56 //y2=0.365
cc_197 ( N_noxref_3_c_194_n N_C_c_486_n ) capacitor c=0.0467448f //x=4.285 \
 //y=4.705 //x2=5.18 //y2=4.54
cc_198 ( N_noxref_3_c_254_p N_C_c_486_n ) capacitor c=0.00146509f //x=4.705 \
 //y=4.795 //x2=5.18 //y2=4.54
cc_199 ( N_noxref_3_c_201_n N_C_c_486_n ) capacitor c=0.00112871f //x=4.285 \
 //y=4.705 //x2=5.18 //y2=4.54
cc_200 ( N_noxref_3_c_161_n N_C_c_474_n ) capacitor c=0.00732168f //x=4.325 \
 //y=2.59 //x2=5.18 //y2=2.08
cc_201 ( N_noxref_3_c_167_n N_C_c_474_n ) capacitor c=9.8819e-19 //x=2.59 \
 //y=2.59 //x2=5.18 //y2=2.08
cc_202 ( N_noxref_3_c_169_n N_C_c_474_n ) capacitor c=0.0444015f //x=4.44 \
 //y=2.08 //x2=5.18 //y2=2.08
cc_203 ( N_noxref_3_c_174_n N_C_c_474_n ) capacitor c=0.00308814f //x=4.245 \
 //y=1.915 //x2=5.18 //y2=2.08
cc_204 ( N_noxref_3_M8_noxref_g N_C_M10_noxref_g ) capacitor c=0.0100243f \
 //x=4.34 //y=6.025 //x2=5.22 //y2=6.025
cc_205 ( N_noxref_3_M9_noxref_g N_C_M10_noxref_g ) capacitor c=0.107798f \
 //x=4.78 //y=6.025 //x2=5.22 //y2=6.025
cc_206 ( N_noxref_3_M9_noxref_g N_C_M11_noxref_g ) capacitor c=0.0094155f \
 //x=4.78 //y=6.025 //x2=5.66 //y2=6.025
cc_207 ( N_noxref_3_c_172_n N_C_c_476_n ) capacitor c=0.00125788f //x=4.245 \
 //y=0.905 //x2=5.215 //y2=0.905
cc_208 ( N_noxref_3_c_177_n N_C_c_476_n ) capacitor c=0.0126654f //x=4.775 \
 //y=0.905 //x2=5.215 //y2=0.905
cc_209 ( N_noxref_3_c_265_p N_C_c_498_n ) capacitor c=0.00148539f //x=4.245 \
 //y=1.25 //x2=5.215 //y2=1.255
cc_210 ( N_noxref_3_c_266_p N_C_c_498_n ) capacitor c=0.00105591f //x=4.245 \
 //y=1.56 //x2=5.215 //y2=1.255
cc_211 ( N_noxref_3_c_179_n N_C_c_498_n ) capacitor c=0.0126654f //x=4.775 \
 //y=1.25 //x2=5.215 //y2=1.255
cc_212 ( N_noxref_3_c_266_p N_C_c_501_n ) capacitor c=0.00109549f //x=4.245 \
 //y=1.56 //x2=5.215 //y2=1.56
cc_213 ( N_noxref_3_c_179_n N_C_c_501_n ) capacitor c=0.00886999f //x=4.775 \
 //y=1.25 //x2=5.215 //y2=1.56
cc_214 ( N_noxref_3_c_179_n N_C_c_479_n ) capacitor c=0.00123863f //x=4.775 \
 //y=1.25 //x2=5.59 //y2=1.405
cc_215 ( N_noxref_3_c_177_n N_C_c_480_n ) capacitor c=0.00132934f //x=4.775 \
 //y=0.905 //x2=5.745 //y2=0.905
cc_216 ( N_noxref_3_c_179_n N_C_c_505_n ) capacitor c=0.00150734f //x=4.775 \
 //y=1.25 //x2=5.745 //y2=1.255
cc_217 ( N_noxref_3_c_169_n N_C_c_506_n ) capacitor c=0.00307062f //x=4.44 \
 //y=2.08 //x2=5.18 //y2=2.08
cc_218 ( N_noxref_3_c_174_n N_C_c_506_n ) capacitor c=0.0179092f //x=4.245 \
 //y=1.915 //x2=5.18 //y2=2.08
cc_219 ( N_noxref_3_c_174_n N_C_c_508_n ) capacitor c=0.00577193f //x=4.245 \
 //y=1.915 //x2=5.18 //y2=1.915
cc_220 ( N_noxref_3_c_194_n N_C_c_509_n ) capacitor c=0.00336963f //x=4.285 \
 //y=4.705 //x2=5.215 //y2=4.705
cc_221 ( N_noxref_3_c_254_p N_C_c_509_n ) capacitor c=0.020271f //x=4.705 \
 //y=4.795 //x2=5.215 //y2=4.705
cc_222 ( N_noxref_3_c_201_n N_C_c_509_n ) capacitor c=0.00546725f //x=4.285 \
 //y=4.705 //x2=5.215 //y2=4.705
cc_223 ( N_noxref_3_c_167_n YN ) capacitor c=3.55699e-19 //x=2.59 //y=2.59 \
 //x2=5.92 //y2=2.22
cc_224 ( N_noxref_3_c_169_n YN ) capacitor c=0.00392263f //x=4.44 //y=2.08 \
 //x2=5.92 //y2=2.22
cc_225 ( N_noxref_3_c_179_n N_YN_c_543_n ) capacitor c=0.00431513f //x=4.775 \
 //y=1.25 //x2=5.395 //y2=1.655
cc_226 ( N_noxref_3_c_161_n N_YN_c_567_n ) capacitor c=0.0018301f //x=4.325 \
 //y=2.59 //x2=4.595 //y2=1.655
cc_227 ( N_noxref_3_c_169_n N_YN_c_567_n ) capacitor c=0.0107041f //x=4.44 \
 //y=2.08 //x2=4.595 //y2=1.655
cc_228 ( N_noxref_3_c_174_n N_YN_c_567_n ) capacitor c=0.00524371f //x=4.245 \
 //y=1.915 //x2=4.595 //y2=1.655
cc_229 ( N_noxref_3_c_172_n N_YN_M2_noxref_d ) capacitor c=0.0013184f \
 //x=4.245 //y=0.905 //x2=4.32 //y2=0.905
cc_230 ( N_noxref_3_c_265_p N_YN_M2_noxref_d ) capacitor c=0.0034598f \
 //x=4.245 //y=1.25 //x2=4.32 //y2=0.905
cc_231 ( N_noxref_3_c_266_p N_YN_M2_noxref_d ) capacitor c=0.00300148f \
 //x=4.245 //y=1.56 //x2=4.32 //y2=0.905
cc_232 ( N_noxref_3_c_174_n N_YN_M2_noxref_d ) capacitor c=0.00273686f \
 //x=4.245 //y=1.915 //x2=4.32 //y2=0.905
cc_233 ( N_noxref_3_c_176_n N_YN_M2_noxref_d ) capacitor c=0.00241102f \
 //x=4.62 //y=0.75 //x2=4.32 //y2=0.905
cc_234 ( N_noxref_3_c_290_p N_YN_M2_noxref_d ) capacitor c=0.0123304f //x=4.62 \
 //y=1.405 //x2=4.32 //y2=0.905
cc_235 ( N_noxref_3_c_177_n N_YN_M2_noxref_d ) capacitor c=0.00219619f \
 //x=4.775 //y=0.905 //x2=4.32 //y2=0.905
cc_236 ( N_noxref_3_c_179_n N_YN_M2_noxref_d ) capacitor c=0.00603828f \
 //x=4.775 //y=1.25 //x2=4.32 //y2=0.905
cc_237 ( N_noxref_3_c_194_n N_noxref_9_c_609_n ) capacitor c=0.00630079f \
 //x=4.285 //y=4.705 //x2=4.915 //y2=5.21
cc_238 ( N_noxref_3_M8_noxref_g N_noxref_9_c_609_n ) capacitor c=0.0182669f \
 //x=4.34 //y=6.025 //x2=4.915 //y2=5.21
cc_239 ( N_noxref_3_M9_noxref_g N_noxref_9_c_609_n ) capacitor c=0.0204082f \
 //x=4.78 //y=6.025 //x2=4.915 //y2=5.21
cc_240 ( N_noxref_3_c_254_p N_noxref_9_c_609_n ) capacitor c=0.00365818f \
 //x=4.705 //y=4.795 //x2=4.915 //y2=5.21
cc_241 ( N_noxref_3_c_201_n N_noxref_9_c_609_n ) capacitor c=0.0017421f \
 //x=4.285 //y=4.705 //x2=4.915 //y2=5.21
cc_242 ( N_noxref_3_c_189_n N_noxref_9_c_612_n ) capacitor c=2.87761e-19 \
 //x=2.505 //y=5.2 //x2=4.205 //y2=5.21
cc_243 ( N_noxref_3_c_194_n N_noxref_9_c_612_n ) capacitor c=0.0118415f \
 //x=4.285 //y=4.705 //x2=4.205 //y2=5.21
cc_244 ( N_noxref_3_c_201_n N_noxref_9_c_612_n ) capacitor c=0.00613395f \
 //x=4.285 //y=4.705 //x2=4.205 //y2=5.21
cc_245 ( N_noxref_3_M6_noxref_d N_noxref_9_c_612_n ) capacitor c=4.5543e-19 \
 //x=1.965 //y=5.02 //x2=4.205 //y2=5.21
cc_246 ( N_noxref_3_M8_noxref_g N_noxref_9_M8_noxref_s ) capacitor \
 c=0.0473218f //x=4.34 //y=6.025 //x2=3.985 //y2=5.025
cc_247 ( N_noxref_3_M9_noxref_g N_noxref_9_M9_noxref_d ) capacitor \
 c=0.0170604f //x=4.78 //y=6.025 //x2=4.855 //y2=5.025
cc_248 ( N_A_c_304_n N_B_c_368_n ) capacitor c=0.00400249f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=4.535
cc_249 ( N_A_c_321_n N_B_c_368_n ) capacitor c=0.00417994f //x=1.11 //y=4.7 \
 //x2=1.85 //y2=4.535
cc_250 ( N_A_c_304_n N_B_c_359_n ) capacitor c=0.0887263f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=2.08
cc_251 ( N_A_c_309_n N_B_c_359_n ) capacitor c=0.00308814f //x=0.915 //y=1.915 \
 //x2=1.85 //y2=2.08
cc_252 ( N_A_M4_noxref_g N_B_M6_noxref_g ) capacitor c=0.0104611f //x=1.01 \
 //y=6.02 //x2=1.89 //y2=6.02
cc_253 ( N_A_M5_noxref_g N_B_M6_noxref_g ) capacitor c=0.106811f //x=1.45 \
 //y=6.02 //x2=1.89 //y2=6.02
cc_254 ( N_A_M5_noxref_g N_B_M7_noxref_g ) capacitor c=0.0100341f //x=1.45 \
 //y=6.02 //x2=2.33 //y2=6.02
cc_255 ( N_A_c_305_n N_B_c_377_n ) capacitor c=4.86506e-19 //x=0.915 //y=0.865 \
 //x2=1.885 //y2=0.905
cc_256 ( N_A_c_307_n N_B_c_377_n ) capacitor c=0.00152104f //x=0.915 //y=1.21 \
 //x2=1.885 //y2=0.905
cc_257 ( N_A_c_312_n N_B_c_377_n ) capacitor c=0.0151475f //x=1.445 //y=0.865 \
 //x2=1.885 //y2=0.905
cc_258 ( N_A_c_308_n N_B_c_378_n ) capacitor c=0.00109982f //x=0.915 //y=1.52 \
 //x2=1.885 //y2=1.25
cc_259 ( N_A_c_314_n N_B_c_378_n ) capacitor c=0.0111064f //x=1.445 //y=1.21 \
 //x2=1.885 //y2=1.25
cc_260 ( N_A_c_308_n N_B_c_379_n ) capacitor c=9.57794e-19 //x=0.915 //y=1.52 \
 //x2=1.885 //y2=1.56
cc_261 ( N_A_c_309_n N_B_c_379_n ) capacitor c=0.00662747f //x=0.915 //y=1.915 \
 //x2=1.885 //y2=1.56
cc_262 ( N_A_c_314_n N_B_c_379_n ) capacitor c=0.00862358f //x=1.445 //y=1.21 \
 //x2=1.885 //y2=1.56
cc_263 ( N_A_c_312_n N_B_c_385_n ) capacitor c=0.00124821f //x=1.445 //y=0.865 \
 //x2=2.415 //y2=0.905
cc_264 ( N_A_c_314_n N_B_c_386_n ) capacitor c=0.00200715f //x=1.445 //y=1.21 \
 //x2=2.415 //y2=1.25
cc_265 ( N_A_c_304_n N_B_c_388_n ) capacitor c=0.00307062f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=2.08
cc_266 ( N_A_c_309_n N_B_c_388_n ) capacitor c=0.0179092f //x=0.915 //y=1.915 \
 //x2=1.85 //y2=2.08
cc_267 ( N_A_c_304_n N_B_c_391_n ) capacitor c=0.00344981f //x=1.11 //y=2.08 \
 //x2=1.88 //y2=4.7
cc_268 ( N_A_c_321_n N_B_c_391_n ) capacitor c=0.0293367f //x=1.11 //y=4.7 \
 //x2=1.88 //y2=4.7
cc_269 ( N_A_c_309_n N_noxref_6_c_447_n ) capacitor c=0.0034165f //x=0.915 \
 //y=1.915 //x2=0.695 //y2=1.495
cc_270 ( N_A_c_304_n N_noxref_6_c_423_n ) capacitor c=0.0118986f //x=1.11 \
 //y=2.08 //x2=1.58 //y2=1.58
cc_271 ( N_A_c_308_n N_noxref_6_c_423_n ) capacitor c=0.00703567f //x=0.915 \
 //y=1.52 //x2=1.58 //y2=1.58
cc_272 ( N_A_c_309_n N_noxref_6_c_423_n ) capacitor c=0.0216532f //x=0.915 \
 //y=1.915 //x2=1.58 //y2=1.58
cc_273 ( N_A_c_311_n N_noxref_6_c_423_n ) capacitor c=0.00780629f //x=1.29 \
 //y=1.365 //x2=1.58 //y2=1.58
cc_274 ( N_A_c_314_n N_noxref_6_c_423_n ) capacitor c=0.00339872f //x=1.445 \
 //y=1.21 //x2=1.58 //y2=1.58
cc_275 ( N_A_c_309_n N_noxref_6_c_431_n ) capacitor c=6.71402e-19 //x=0.915 \
 //y=1.915 //x2=1.665 //y2=1.495
cc_276 ( N_A_c_305_n N_noxref_6_M0_noxref_s ) capacitor c=0.0326577f //x=0.915 \
 //y=0.865 //x2=0.56 //y2=0.365
cc_277 ( N_A_c_308_n N_noxref_6_M0_noxref_s ) capacitor c=3.48408e-19 \
 //x=0.915 //y=1.52 //x2=0.56 //y2=0.365
cc_278 ( N_A_c_312_n N_noxref_6_M0_noxref_s ) capacitor c=0.0120759f //x=1.445 \
 //y=0.865 //x2=0.56 //y2=0.365
cc_279 ( N_B_c_379_n N_noxref_6_c_431_n ) capacitor c=0.00623646f //x=1.885 \
 //y=1.56 //x2=1.665 //y2=1.495
cc_280 ( N_B_c_388_n N_noxref_6_c_431_n ) capacitor c=0.00172768f //x=1.85 \
 //y=2.08 //x2=1.665 //y2=1.495
cc_281 ( N_B_c_359_n N_noxref_6_c_432_n ) capacitor c=0.00161845f //x=1.85 \
 //y=2.08 //x2=2.55 //y2=0.53
cc_282 ( N_B_c_377_n N_noxref_6_c_432_n ) capacitor c=0.0186143f //x=1.885 \
 //y=0.905 //x2=2.55 //y2=0.53
cc_283 ( N_B_c_385_n N_noxref_6_c_432_n ) capacitor c=0.00656458f //x=2.415 \
 //y=0.905 //x2=2.55 //y2=0.53
cc_284 ( N_B_c_388_n N_noxref_6_c_432_n ) capacitor c=2.1838e-19 //x=1.85 \
 //y=2.08 //x2=2.55 //y2=0.53
cc_285 ( N_B_c_377_n N_noxref_6_M0_noxref_s ) capacitor c=0.00623646f \
 //x=1.885 //y=0.905 //x2=0.56 //y2=0.365
cc_286 ( N_B_c_385_n N_noxref_6_M0_noxref_s ) capacitor c=0.0143002f //x=2.415 \
 //y=0.905 //x2=0.56 //y2=0.365
cc_287 ( N_B_c_386_n N_noxref_6_M0_noxref_s ) capacitor c=0.00290153f \
 //x=2.415 //y=1.25 //x2=0.56 //y2=0.365
cc_288 ( N_C_c_486_n YN ) capacitor c=0.0102183f //x=5.18 //y=4.54 //x2=5.92 \
 //y2=2.22
cc_289 ( N_C_c_474_n YN ) capacitor c=0.0837373f //x=5.18 //y=2.08 //x2=5.92 \
 //y2=2.22
cc_290 ( N_C_c_514_p YN ) capacitor c=0.0144455f //x=5.585 //y=4.795 //x2=5.92 \
 //y2=2.22
cc_291 ( N_C_c_506_n YN ) capacitor c=0.00877984f //x=5.18 //y=2.08 //x2=5.92 \
 //y2=2.22
cc_292 ( N_C_c_508_n YN ) capacitor c=0.00306024f //x=5.18 //y=1.915 //x2=5.92 \
 //y2=2.22
cc_293 ( N_C_c_509_n YN ) capacitor c=0.00537091f //x=5.215 //y=4.705 \
 //x2=5.92 //y2=2.22
cc_294 ( N_C_c_474_n N_YN_c_543_n ) capacitor c=0.0162392f //x=5.18 //y=2.08 \
 //x2=5.395 //y2=1.655
cc_295 ( N_C_c_501_n N_YN_c_543_n ) capacitor c=0.00218915f //x=5.215 //y=1.56 \
 //x2=5.395 //y2=1.655
cc_296 ( N_C_c_506_n N_YN_c_543_n ) capacitor c=0.00633758f //x=5.18 //y=2.08 \
 //x2=5.395 //y2=1.655
cc_297 ( N_C_c_508_n N_YN_c_543_n ) capacitor c=0.0189958f //x=5.18 //y=1.915 \
 //x2=5.395 //y2=1.655
cc_298 ( N_C_M11_noxref_g N_YN_c_560_n ) capacitor c=0.0217751f //x=5.66 \
 //y=6.025 //x2=5.835 //y2=5.21
cc_299 ( N_C_M10_noxref_g N_YN_c_561_n ) capacitor c=0.0132788f //x=5.22 \
 //y=6.025 //x2=5.525 //y2=5.21
cc_300 ( N_C_c_514_p N_YN_c_561_n ) capacitor c=0.00417892f //x=5.585 \
 //y=4.795 //x2=5.525 //y2=5.21
cc_301 ( N_C_c_479_n N_YN_c_547_n ) capacitor c=0.00801563f //x=5.59 //y=1.405 \
 //x2=5.835 //y2=1.655
cc_302 ( N_C_c_501_n N_YN_M2_noxref_d ) capacitor c=0.00148728f //x=5.215 \
 //y=1.56 //x2=4.32 //y2=0.905
cc_303 ( N_C_c_476_n N_YN_M3_noxref_d ) capacitor c=0.00226395f //x=5.215 \
 //y=0.905 //x2=5.29 //y2=0.905
cc_304 ( N_C_c_498_n N_YN_M3_noxref_d ) capacitor c=0.0035101f //x=5.215 \
 //y=1.255 //x2=5.29 //y2=0.905
cc_305 ( N_C_c_501_n N_YN_M3_noxref_d ) capacitor c=0.00546704f //x=5.215 \
 //y=1.56 //x2=5.29 //y2=0.905
cc_306 ( N_C_c_478_n N_YN_M3_noxref_d ) capacitor c=0.00241102f //x=5.59 \
 //y=0.75 //x2=5.29 //y2=0.905
cc_307 ( N_C_c_479_n N_YN_M3_noxref_d ) capacitor c=0.0158021f //x=5.59 \
 //y=1.405 //x2=5.29 //y2=0.905
cc_308 ( N_C_c_480_n N_YN_M3_noxref_d ) capacitor c=0.00132831f //x=5.745 \
 //y=0.905 //x2=5.29 //y2=0.905
cc_309 ( N_C_c_505_n N_YN_M3_noxref_d ) capacitor c=0.0035101f //x=5.745 \
 //y=1.255 //x2=5.29 //y2=0.905
cc_310 ( N_C_c_508_n N_YN_M3_noxref_d ) capacitor c=3.4952e-19 //x=5.18 \
 //y=1.915 //x2=5.29 //y2=0.905
cc_311 ( N_C_M11_noxref_g N_YN_M10_noxref_d ) capacitor c=0.0136385f //x=5.66 \
 //y=6.025 //x2=5.295 //y2=5.025
cc_312 ( N_C_M10_noxref_g N_noxref_9_c_609_n ) capacitor c=0.0170604f //x=5.22 \
 //y=6.025 //x2=4.915 //y2=5.21
cc_313 ( N_C_c_509_n N_noxref_9_c_609_n ) capacitor c=2.3112e-19 //x=5.215 \
 //y=4.705 //x2=4.915 //y2=5.21
cc_314 ( N_C_c_486_n N_noxref_9_c_613_n ) capacitor c=0.00109004f //x=5.18 \
 //y=4.54 //x2=5.795 //y2=6.91
cc_315 ( N_C_M10_noxref_g N_noxref_9_c_613_n ) capacitor c=0.0148484f //x=5.22 \
 //y=6.025 //x2=5.795 //y2=6.91
cc_316 ( N_C_M11_noxref_g N_noxref_9_c_613_n ) capacitor c=0.0163196f //x=5.66 \
 //y=6.025 //x2=5.795 //y2=6.91
cc_317 ( N_C_M11_noxref_g N_noxref_9_M11_noxref_d ) capacitor c=0.0351101f \
 //x=5.66 //y=6.025 //x2=5.735 //y2=5.025
cc_318 ( N_YN_c_561_n N_noxref_9_c_609_n ) capacitor c=0.0348754f //x=5.525 \
 //y=5.21 //x2=4.915 //y2=5.21
cc_319 ( N_YN_c_560_n N_noxref_9_c_613_n ) capacitor c=0.00194034f //x=5.835 \
 //y=5.21 //x2=5.795 //y2=6.91
cc_320 ( N_YN_M10_noxref_d N_noxref_9_c_613_n ) capacitor c=0.0118172f \
 //x=5.295 //y=5.025 //x2=5.795 //y2=6.91
cc_321 ( N_YN_M10_noxref_d N_noxref_9_M8_noxref_s ) capacitor c=0.00107541f \
 //x=5.295 //y=5.025 //x2=3.985 //y2=5.025
cc_322 ( N_YN_M10_noxref_d N_noxref_9_M9_noxref_d ) capacitor c=0.0348754f \
 //x=5.295 //y=5.025 //x2=4.855 //y2=5.025
cc_323 ( N_YN_c_560_n N_noxref_9_M11_noxref_d ) capacitor c=0.0164221f \
 //x=5.835 //y=5.21 //x2=5.735 //y2=5.025
cc_324 ( N_YN_M10_noxref_d N_noxref_9_M11_noxref_d ) capacitor c=0.0458293f \
 //x=5.295 //y=5.025 //x2=5.735 //y2=5.025
