magic
tech sky130A
magscale 1 2
timestamp 1669507611
<< nwell >>
rect -87 786 4083 1550
<< pwell >>
rect -34 -34 4030 544
<< nmos >>
rect 155 297 185 350
tri 185 297 201 313 sw
rect 155 267 261 297
tri 261 267 291 297 sw
rect 155 166 185 267
tri 185 251 201 267 nw
tri 245 251 261 267 ne
tri 185 166 201 182 sw
tri 245 166 261 182 se
rect 261 166 291 267
tri 155 136 185 166 ne
rect 185 136 261 166
tri 261 136 291 166 nw
rect 612 288 642 349
tri 642 288 658 304 sw
rect 806 296 836 349
tri 836 296 852 312 sw
rect 612 258 718 288
tri 718 258 748 288 sw
rect 806 266 912 296
tri 912 266 942 296 sw
rect 612 157 642 258
tri 642 242 658 258 nw
tri 702 242 718 258 ne
tri 642 157 658 173 sw
tri 702 157 718 173 se
rect 718 157 748 258
rect 806 165 836 266
tri 836 250 852 266 nw
tri 896 250 912 266 ne
tri 836 165 852 181 sw
tri 896 165 912 181 se
rect 912 165 942 266
tri 612 127 642 157 ne
rect 642 127 718 157
tri 718 127 748 157 nw
tri 806 135 836 165 ne
rect 836 135 912 165
tri 912 135 942 165 nw
rect 1265 297 1295 350
tri 1295 297 1311 313 sw
rect 1265 267 1371 297
tri 1371 267 1401 297 sw
rect 1265 166 1295 267
tri 1295 251 1311 267 nw
tri 1355 251 1371 267 ne
tri 1295 166 1311 182 sw
tri 1355 166 1371 182 se
rect 1371 166 1401 267
tri 1265 136 1295 166 ne
rect 1295 136 1371 166
tri 1371 136 1401 166 nw
rect 1722 288 1752 349
tri 1752 288 1768 304 sw
rect 1916 296 1946 349
tri 1946 296 1962 312 sw
rect 1722 258 1828 288
tri 1828 258 1858 288 sw
rect 1916 266 2022 296
tri 2022 266 2052 296 sw
rect 1722 157 1752 258
tri 1752 242 1768 258 nw
tri 1812 242 1828 258 ne
tri 1752 157 1768 173 sw
tri 1812 157 1828 173 se
rect 1828 157 1858 258
rect 1916 165 1946 266
tri 1946 250 1962 266 nw
tri 2006 250 2022 266 ne
tri 1946 165 1962 181 sw
tri 2006 165 2022 181 se
rect 2022 165 2052 266
tri 1722 127 1752 157 ne
rect 1752 127 1828 157
tri 1828 127 1858 157 nw
tri 1916 135 1946 165 ne
rect 1946 135 2022 165
tri 2022 135 2052 165 nw
rect 2375 297 2405 350
tri 2405 297 2421 313 sw
rect 2375 267 2481 297
tri 2481 267 2511 297 sw
rect 2375 166 2405 267
tri 2405 251 2421 267 nw
tri 2465 251 2481 267 ne
tri 2405 166 2421 182 sw
tri 2465 166 2481 182 se
rect 2481 166 2511 267
tri 2375 136 2405 166 ne
rect 2405 136 2481 166
tri 2481 136 2511 166 nw
rect 2832 296 2862 349
tri 2862 296 2878 312 sw
rect 3026 296 3056 349
tri 3056 296 3072 312 sw
rect 2832 266 2938 296
tri 2938 266 2968 296 sw
rect 2832 165 2862 266
tri 2862 250 2878 266 nw
tri 2922 250 2938 266 ne
tri 2862 165 2878 181 sw
tri 2922 165 2938 181 se
rect 2938 165 2968 266
rect 3026 266 3132 296
tri 3132 266 3162 296 sw
rect 3026 251 3057 266
tri 3057 251 3072 266 nw
tri 3116 251 3131 266 ne
rect 3131 251 3162 266
tri 2832 135 2862 165 ne
rect 2862 135 2938 165
tri 2938 135 2968 165 nw
rect 3026 165 3056 251
tri 3056 165 3072 181 sw
tri 3116 165 3132 181 se
rect 3132 165 3162 251
tri 3026 135 3056 165 ne
rect 3056 135 3132 165
tri 3132 135 3162 165 nw
rect 3498 296 3528 349
tri 3528 296 3544 312 sw
rect 3692 296 3722 349
tri 3722 296 3738 312 sw
rect 3498 266 3604 296
tri 3604 266 3634 296 sw
rect 3498 165 3528 266
tri 3528 250 3544 266 nw
tri 3588 250 3604 266 ne
tri 3528 165 3544 181 sw
tri 3588 165 3604 181 se
rect 3604 165 3634 266
rect 3692 266 3798 296
tri 3798 266 3828 296 sw
rect 3692 251 3723 266
tri 3723 251 3738 266 nw
tri 3782 251 3797 266 ne
rect 3797 251 3828 266
tri 3498 135 3528 165 ne
rect 3528 135 3604 165
tri 3604 135 3634 165 nw
rect 3692 165 3722 251
tri 3722 165 3738 181 sw
tri 3782 165 3798 181 se
rect 3798 165 3828 251
tri 3692 135 3722 165 ne
rect 3722 135 3798 165
tri 3798 135 3828 165 nw
<< pmos >>
rect 164 1004 194 1404
rect 252 1004 282 1404
rect 631 1004 661 1404
rect 719 1004 749 1404
rect 807 1004 837 1404
rect 895 1004 925 1404
rect 1274 1004 1304 1404
rect 1362 1004 1392 1404
rect 1741 1004 1771 1404
rect 1829 1004 1859 1404
rect 1917 1004 1947 1404
rect 2005 1004 2035 1404
rect 2384 1004 2414 1404
rect 2472 1004 2502 1404
rect 2851 1005 2881 1405
rect 2939 1005 2969 1405
rect 3027 1005 3057 1405
rect 3115 1005 3145 1405
rect 3517 1005 3547 1405
rect 3605 1005 3635 1405
rect 3693 1005 3723 1405
rect 3781 1005 3811 1405
<< ndiff >>
rect 99 334 155 350
rect 99 300 109 334
rect 143 300 155 334
rect 99 262 155 300
rect 185 334 345 350
rect 185 313 303 334
tri 185 297 201 313 ne
rect 201 300 303 313
rect 337 300 345 334
rect 201 297 345 300
tri 261 267 291 297 ne
rect 99 228 109 262
rect 143 228 155 262
rect 99 194 155 228
rect 99 160 109 194
rect 143 160 155 194
tri 185 251 201 267 se
rect 201 251 245 267
tri 245 251 261 267 sw
rect 185 218 261 251
rect 185 184 205 218
rect 239 184 261 218
rect 185 182 261 184
tri 185 166 201 182 ne
rect 201 166 245 182
tri 245 166 261 182 nw
rect 291 262 345 297
rect 291 228 303 262
rect 337 228 345 262
rect 291 194 345 228
rect 99 136 155 160
tri 155 136 185 166 sw
tri 261 136 291 166 se
rect 291 160 303 194
rect 337 160 345 194
rect 291 136 345 160
rect 99 124 345 136
rect 99 90 109 124
rect 143 90 205 124
rect 239 90 303 124
rect 337 90 345 124
rect 99 74 345 90
rect 556 333 612 349
rect 556 299 566 333
rect 600 299 612 333
rect 556 261 612 299
rect 642 333 806 349
rect 642 304 663 333
tri 642 288 658 304 ne
rect 658 299 663 304
rect 697 299 760 333
rect 794 299 806 333
rect 658 288 806 299
rect 836 312 998 349
tri 836 296 852 312 ne
rect 852 296 998 312
rect 556 227 566 261
rect 600 227 612 261
tri 718 258 748 288 ne
rect 748 261 806 288
tri 912 266 942 296 ne
rect 556 193 612 227
rect 556 159 566 193
rect 600 159 612 193
rect 556 127 612 159
tri 642 242 658 258 se
rect 658 242 702 258
tri 702 242 718 258 sw
rect 642 208 718 242
rect 642 174 663 208
rect 697 174 718 208
rect 642 173 718 174
tri 642 157 658 173 ne
rect 658 157 702 173
tri 702 157 718 173 nw
rect 748 227 760 261
rect 794 227 806 261
rect 748 193 806 227
rect 748 159 760 193
rect 794 159 806 193
tri 836 250 852 266 se
rect 852 250 896 266
tri 896 250 912 266 sw
rect 836 217 912 250
rect 836 183 857 217
rect 891 183 912 217
rect 836 181 912 183
tri 836 165 852 181 ne
rect 852 165 896 181
tri 896 165 912 181 nw
rect 942 261 998 296
rect 942 227 954 261
rect 988 227 998 261
rect 942 193 998 227
tri 612 127 642 157 sw
tri 718 127 748 157 se
rect 748 135 806 159
tri 806 135 836 165 sw
tri 912 135 942 165 se
rect 942 159 954 193
rect 988 159 998 193
rect 942 135 998 159
rect 748 127 998 135
rect 556 123 998 127
rect 556 89 566 123
rect 600 89 760 123
rect 794 89 857 123
rect 891 89 954 123
rect 988 89 998 123
rect 556 73 998 89
rect 1209 334 1265 350
rect 1209 300 1219 334
rect 1253 300 1265 334
rect 1209 262 1265 300
rect 1295 334 1455 350
rect 1295 313 1413 334
tri 1295 297 1311 313 ne
rect 1311 300 1413 313
rect 1447 300 1455 334
rect 1311 297 1455 300
tri 1371 267 1401 297 ne
rect 1209 228 1219 262
rect 1253 228 1265 262
rect 1209 194 1265 228
rect 1209 160 1219 194
rect 1253 160 1265 194
tri 1295 251 1311 267 se
rect 1311 251 1355 267
tri 1355 251 1371 267 sw
rect 1295 218 1371 251
rect 1295 184 1315 218
rect 1349 184 1371 218
rect 1295 182 1371 184
tri 1295 166 1311 182 ne
rect 1311 166 1355 182
tri 1355 166 1371 182 nw
rect 1401 262 1455 297
rect 1401 228 1413 262
rect 1447 228 1455 262
rect 1401 194 1455 228
rect 1209 136 1265 160
tri 1265 136 1295 166 sw
tri 1371 136 1401 166 se
rect 1401 160 1413 194
rect 1447 160 1455 194
rect 1401 136 1455 160
rect 1209 124 1455 136
rect 1209 90 1219 124
rect 1253 90 1315 124
rect 1349 90 1413 124
rect 1447 90 1455 124
rect 1209 74 1455 90
rect 1666 333 1722 349
rect 1666 299 1676 333
rect 1710 299 1722 333
rect 1666 261 1722 299
rect 1752 333 1916 349
rect 1752 304 1773 333
tri 1752 288 1768 304 ne
rect 1768 299 1773 304
rect 1807 299 1870 333
rect 1904 299 1916 333
rect 1768 288 1916 299
rect 1946 312 2108 349
tri 1946 296 1962 312 ne
rect 1962 296 2108 312
rect 1666 227 1676 261
rect 1710 227 1722 261
tri 1828 258 1858 288 ne
rect 1858 261 1916 288
tri 2022 266 2052 296 ne
rect 1666 193 1722 227
rect 1666 159 1676 193
rect 1710 159 1722 193
rect 1666 127 1722 159
tri 1752 242 1768 258 se
rect 1768 242 1812 258
tri 1812 242 1828 258 sw
rect 1752 208 1828 242
rect 1752 174 1773 208
rect 1807 174 1828 208
rect 1752 173 1828 174
tri 1752 157 1768 173 ne
rect 1768 157 1812 173
tri 1812 157 1828 173 nw
rect 1858 227 1870 261
rect 1904 227 1916 261
rect 1858 193 1916 227
rect 1858 159 1870 193
rect 1904 159 1916 193
tri 1946 250 1962 266 se
rect 1962 250 2006 266
tri 2006 250 2022 266 sw
rect 1946 217 2022 250
rect 1946 183 1967 217
rect 2001 183 2022 217
rect 1946 181 2022 183
tri 1946 165 1962 181 ne
rect 1962 165 2006 181
tri 2006 165 2022 181 nw
rect 2052 261 2108 296
rect 2052 227 2064 261
rect 2098 227 2108 261
rect 2052 193 2108 227
tri 1722 127 1752 157 sw
tri 1828 127 1858 157 se
rect 1858 135 1916 159
tri 1916 135 1946 165 sw
tri 2022 135 2052 165 se
rect 2052 159 2064 193
rect 2098 159 2108 193
rect 2052 135 2108 159
rect 1858 127 2108 135
rect 1666 123 2108 127
rect 1666 89 1676 123
rect 1710 89 1870 123
rect 1904 89 1967 123
rect 2001 89 2064 123
rect 2098 89 2108 123
rect 1666 73 2108 89
rect 2319 334 2375 350
rect 2319 300 2329 334
rect 2363 300 2375 334
rect 2319 262 2375 300
rect 2405 334 2565 350
rect 2405 313 2523 334
tri 2405 297 2421 313 ne
rect 2421 300 2523 313
rect 2557 300 2565 334
rect 2421 297 2565 300
tri 2481 267 2511 297 ne
rect 2319 228 2329 262
rect 2363 228 2375 262
rect 2319 194 2375 228
rect 2319 160 2329 194
rect 2363 160 2375 194
tri 2405 251 2421 267 se
rect 2421 251 2465 267
tri 2465 251 2481 267 sw
rect 2405 218 2481 251
rect 2405 184 2425 218
rect 2459 184 2481 218
rect 2405 182 2481 184
tri 2405 166 2421 182 ne
rect 2421 166 2465 182
tri 2465 166 2481 182 nw
rect 2511 262 2565 297
rect 2511 228 2523 262
rect 2557 228 2565 262
rect 2511 194 2565 228
rect 2319 136 2375 160
tri 2375 136 2405 166 sw
tri 2481 136 2511 166 se
rect 2511 160 2523 194
rect 2557 160 2565 194
rect 2511 136 2565 160
rect 2319 124 2565 136
rect 2319 90 2329 124
rect 2363 90 2425 124
rect 2459 90 2523 124
rect 2557 90 2565 124
rect 2319 74 2565 90
rect 2776 333 2832 349
rect 2776 299 2786 333
rect 2820 299 2832 333
rect 2776 261 2832 299
rect 2862 312 3026 349
tri 2862 296 2878 312 ne
rect 2878 296 3026 312
rect 3056 312 3218 349
tri 3056 296 3072 312 ne
rect 3072 296 3218 312
tri 2938 266 2968 296 ne
rect 2776 227 2786 261
rect 2820 227 2832 261
rect 2776 193 2832 227
rect 2776 159 2786 193
rect 2820 159 2832 193
tri 2862 250 2878 266 se
rect 2878 250 2922 266
tri 2922 250 2938 266 sw
rect 2862 217 2938 250
rect 2862 183 2883 217
rect 2917 183 2938 217
rect 2862 181 2938 183
tri 2862 165 2878 181 ne
rect 2878 165 2922 181
tri 2922 165 2938 181 nw
rect 2968 261 3026 296
tri 3132 266 3162 296 ne
rect 2968 227 2980 261
rect 3014 227 3026 261
tri 3057 251 3072 266 se
rect 3072 251 3116 266
tri 3116 251 3131 266 sw
rect 3162 261 3218 296
rect 2968 193 3026 227
rect 2776 135 2832 159
tri 2832 135 2862 165 sw
tri 2938 135 2968 165 se
rect 2968 159 2980 193
rect 3014 159 3026 193
rect 3056 217 3132 251
rect 3056 183 3077 217
rect 3111 183 3132 217
rect 3056 181 3132 183
tri 3056 165 3072 181 ne
rect 3072 165 3116 181
tri 3116 165 3132 181 nw
rect 3162 227 3174 261
rect 3208 227 3218 261
rect 3162 193 3218 227
rect 2968 135 3026 159
tri 3026 135 3056 165 sw
tri 3132 135 3162 165 se
rect 3162 159 3174 193
rect 3208 159 3218 193
rect 3162 135 3218 159
rect 2776 123 3218 135
rect 2776 89 2786 123
rect 2820 89 2883 123
rect 2917 89 2980 123
rect 3014 89 3077 123
rect 3111 89 3174 123
rect 3208 89 3218 123
rect 2776 73 3218 89
rect 3442 333 3498 349
rect 3442 299 3452 333
rect 3486 299 3498 333
rect 3442 261 3498 299
rect 3528 312 3692 349
tri 3528 296 3544 312 ne
rect 3544 296 3692 312
rect 3722 312 3884 349
tri 3722 296 3738 312 ne
rect 3738 296 3884 312
tri 3604 266 3634 296 ne
rect 3442 227 3452 261
rect 3486 227 3498 261
rect 3442 193 3498 227
rect 3442 159 3452 193
rect 3486 159 3498 193
tri 3528 250 3544 266 se
rect 3544 250 3588 266
tri 3588 250 3604 266 sw
rect 3528 217 3604 250
rect 3528 183 3549 217
rect 3583 183 3604 217
rect 3528 181 3604 183
tri 3528 165 3544 181 ne
rect 3544 165 3588 181
tri 3588 165 3604 181 nw
rect 3634 261 3692 296
tri 3798 266 3828 296 ne
rect 3634 227 3646 261
rect 3680 227 3692 261
tri 3723 251 3738 266 se
rect 3738 251 3782 266
tri 3782 251 3797 266 sw
rect 3828 261 3884 296
rect 3634 193 3692 227
rect 3442 135 3498 159
tri 3498 135 3528 165 sw
tri 3604 135 3634 165 se
rect 3634 159 3646 193
rect 3680 159 3692 193
rect 3722 217 3798 251
rect 3722 183 3743 217
rect 3777 183 3798 217
rect 3722 181 3798 183
tri 3722 165 3738 181 ne
rect 3738 165 3782 181
tri 3782 165 3798 181 nw
rect 3828 227 3840 261
rect 3874 227 3884 261
rect 3828 193 3884 227
rect 3634 135 3692 159
tri 3692 135 3722 165 sw
tri 3798 135 3828 165 se
rect 3828 159 3840 193
rect 3874 159 3884 193
rect 3828 135 3884 159
rect 3442 123 3884 135
rect 3442 89 3452 123
rect 3486 89 3549 123
rect 3583 89 3646 123
rect 3680 89 3743 123
rect 3777 89 3840 123
rect 3874 89 3884 123
rect 3442 73 3884 89
<< pdiff >>
rect 108 1366 164 1404
rect 108 1332 118 1366
rect 152 1332 164 1366
rect 108 1298 164 1332
rect 108 1264 118 1298
rect 152 1264 164 1298
rect 108 1230 164 1264
rect 108 1196 118 1230
rect 152 1196 164 1230
rect 108 1162 164 1196
rect 108 1128 118 1162
rect 152 1128 164 1162
rect 108 1093 164 1128
rect 108 1059 118 1093
rect 152 1059 164 1093
rect 108 1004 164 1059
rect 194 1366 252 1404
rect 194 1332 206 1366
rect 240 1332 252 1366
rect 194 1298 252 1332
rect 194 1264 206 1298
rect 240 1264 252 1298
rect 194 1230 252 1264
rect 194 1196 206 1230
rect 240 1196 252 1230
rect 194 1162 252 1196
rect 194 1128 206 1162
rect 240 1128 252 1162
rect 194 1093 252 1128
rect 194 1059 206 1093
rect 240 1059 252 1093
rect 194 1004 252 1059
rect 282 1366 336 1404
rect 282 1332 294 1366
rect 328 1332 336 1366
rect 282 1298 336 1332
rect 282 1264 294 1298
rect 328 1264 336 1298
rect 282 1230 336 1264
rect 282 1196 294 1230
rect 328 1196 336 1230
rect 282 1162 336 1196
rect 282 1128 294 1162
rect 328 1128 336 1162
rect 282 1093 336 1128
rect 282 1059 294 1093
rect 328 1059 336 1093
rect 282 1004 336 1059
rect 575 1366 631 1404
rect 575 1332 585 1366
rect 619 1332 631 1366
rect 575 1298 631 1332
rect 575 1264 585 1298
rect 619 1264 631 1298
rect 575 1230 631 1264
rect 575 1196 585 1230
rect 619 1196 631 1230
rect 575 1162 631 1196
rect 575 1128 585 1162
rect 619 1128 631 1162
rect 575 1093 631 1128
rect 575 1059 585 1093
rect 619 1059 631 1093
rect 575 1004 631 1059
rect 661 1366 719 1404
rect 661 1332 673 1366
rect 707 1332 719 1366
rect 661 1298 719 1332
rect 661 1264 673 1298
rect 707 1264 719 1298
rect 661 1230 719 1264
rect 661 1196 673 1230
rect 707 1196 719 1230
rect 661 1162 719 1196
rect 661 1128 673 1162
rect 707 1128 719 1162
rect 661 1093 719 1128
rect 661 1059 673 1093
rect 707 1059 719 1093
rect 661 1004 719 1059
rect 749 1366 807 1404
rect 749 1332 761 1366
rect 795 1332 807 1366
rect 749 1298 807 1332
rect 749 1264 761 1298
rect 795 1264 807 1298
rect 749 1230 807 1264
rect 749 1196 761 1230
rect 795 1196 807 1230
rect 749 1162 807 1196
rect 749 1128 761 1162
rect 795 1128 807 1162
rect 749 1004 807 1128
rect 837 1366 895 1404
rect 837 1332 849 1366
rect 883 1332 895 1366
rect 837 1298 895 1332
rect 837 1264 849 1298
rect 883 1264 895 1298
rect 837 1230 895 1264
rect 837 1196 849 1230
rect 883 1196 895 1230
rect 837 1162 895 1196
rect 837 1128 849 1162
rect 883 1128 895 1162
rect 837 1093 895 1128
rect 837 1059 849 1093
rect 883 1059 895 1093
rect 837 1004 895 1059
rect 925 1366 979 1404
rect 925 1332 937 1366
rect 971 1332 979 1366
rect 925 1298 979 1332
rect 925 1264 937 1298
rect 971 1264 979 1298
rect 925 1230 979 1264
rect 925 1196 937 1230
rect 971 1196 979 1230
rect 925 1162 979 1196
rect 925 1128 937 1162
rect 971 1128 979 1162
rect 925 1004 979 1128
rect 1218 1366 1274 1404
rect 1218 1332 1228 1366
rect 1262 1332 1274 1366
rect 1218 1298 1274 1332
rect 1218 1264 1228 1298
rect 1262 1264 1274 1298
rect 1218 1230 1274 1264
rect 1218 1196 1228 1230
rect 1262 1196 1274 1230
rect 1218 1162 1274 1196
rect 1218 1128 1228 1162
rect 1262 1128 1274 1162
rect 1218 1093 1274 1128
rect 1218 1059 1228 1093
rect 1262 1059 1274 1093
rect 1218 1004 1274 1059
rect 1304 1366 1362 1404
rect 1304 1332 1316 1366
rect 1350 1332 1362 1366
rect 1304 1298 1362 1332
rect 1304 1264 1316 1298
rect 1350 1264 1362 1298
rect 1304 1230 1362 1264
rect 1304 1196 1316 1230
rect 1350 1196 1362 1230
rect 1304 1162 1362 1196
rect 1304 1128 1316 1162
rect 1350 1128 1362 1162
rect 1304 1093 1362 1128
rect 1304 1059 1316 1093
rect 1350 1059 1362 1093
rect 1304 1004 1362 1059
rect 1392 1366 1446 1404
rect 1392 1332 1404 1366
rect 1438 1332 1446 1366
rect 1392 1298 1446 1332
rect 1392 1264 1404 1298
rect 1438 1264 1446 1298
rect 1392 1230 1446 1264
rect 1392 1196 1404 1230
rect 1438 1196 1446 1230
rect 1392 1162 1446 1196
rect 1392 1128 1404 1162
rect 1438 1128 1446 1162
rect 1392 1093 1446 1128
rect 1392 1059 1404 1093
rect 1438 1059 1446 1093
rect 1392 1004 1446 1059
rect 1685 1366 1741 1404
rect 1685 1332 1695 1366
rect 1729 1332 1741 1366
rect 1685 1298 1741 1332
rect 1685 1264 1695 1298
rect 1729 1264 1741 1298
rect 1685 1230 1741 1264
rect 1685 1196 1695 1230
rect 1729 1196 1741 1230
rect 1685 1162 1741 1196
rect 1685 1128 1695 1162
rect 1729 1128 1741 1162
rect 1685 1093 1741 1128
rect 1685 1059 1695 1093
rect 1729 1059 1741 1093
rect 1685 1004 1741 1059
rect 1771 1366 1829 1404
rect 1771 1332 1783 1366
rect 1817 1332 1829 1366
rect 1771 1298 1829 1332
rect 1771 1264 1783 1298
rect 1817 1264 1829 1298
rect 1771 1230 1829 1264
rect 1771 1196 1783 1230
rect 1817 1196 1829 1230
rect 1771 1162 1829 1196
rect 1771 1128 1783 1162
rect 1817 1128 1829 1162
rect 1771 1093 1829 1128
rect 1771 1059 1783 1093
rect 1817 1059 1829 1093
rect 1771 1004 1829 1059
rect 1859 1366 1917 1404
rect 1859 1332 1871 1366
rect 1905 1332 1917 1366
rect 1859 1298 1917 1332
rect 1859 1264 1871 1298
rect 1905 1264 1917 1298
rect 1859 1230 1917 1264
rect 1859 1196 1871 1230
rect 1905 1196 1917 1230
rect 1859 1162 1917 1196
rect 1859 1128 1871 1162
rect 1905 1128 1917 1162
rect 1859 1004 1917 1128
rect 1947 1366 2005 1404
rect 1947 1332 1959 1366
rect 1993 1332 2005 1366
rect 1947 1298 2005 1332
rect 1947 1264 1959 1298
rect 1993 1264 2005 1298
rect 1947 1230 2005 1264
rect 1947 1196 1959 1230
rect 1993 1196 2005 1230
rect 1947 1162 2005 1196
rect 1947 1128 1959 1162
rect 1993 1128 2005 1162
rect 1947 1093 2005 1128
rect 1947 1059 1959 1093
rect 1993 1059 2005 1093
rect 1947 1004 2005 1059
rect 2035 1366 2089 1404
rect 2035 1332 2047 1366
rect 2081 1332 2089 1366
rect 2035 1298 2089 1332
rect 2035 1264 2047 1298
rect 2081 1264 2089 1298
rect 2035 1230 2089 1264
rect 2035 1196 2047 1230
rect 2081 1196 2089 1230
rect 2035 1162 2089 1196
rect 2035 1128 2047 1162
rect 2081 1128 2089 1162
rect 2035 1004 2089 1128
rect 2328 1366 2384 1404
rect 2328 1332 2338 1366
rect 2372 1332 2384 1366
rect 2328 1298 2384 1332
rect 2328 1264 2338 1298
rect 2372 1264 2384 1298
rect 2328 1230 2384 1264
rect 2328 1196 2338 1230
rect 2372 1196 2384 1230
rect 2328 1162 2384 1196
rect 2328 1128 2338 1162
rect 2372 1128 2384 1162
rect 2328 1093 2384 1128
rect 2328 1059 2338 1093
rect 2372 1059 2384 1093
rect 2328 1004 2384 1059
rect 2414 1366 2472 1404
rect 2414 1332 2426 1366
rect 2460 1332 2472 1366
rect 2414 1298 2472 1332
rect 2414 1264 2426 1298
rect 2460 1264 2472 1298
rect 2414 1230 2472 1264
rect 2414 1196 2426 1230
rect 2460 1196 2472 1230
rect 2414 1162 2472 1196
rect 2414 1128 2426 1162
rect 2460 1128 2472 1162
rect 2414 1093 2472 1128
rect 2414 1059 2426 1093
rect 2460 1059 2472 1093
rect 2414 1004 2472 1059
rect 2502 1366 2556 1404
rect 2502 1332 2514 1366
rect 2548 1332 2556 1366
rect 2502 1298 2556 1332
rect 2502 1264 2514 1298
rect 2548 1264 2556 1298
rect 2502 1230 2556 1264
rect 2502 1196 2514 1230
rect 2548 1196 2556 1230
rect 2502 1162 2556 1196
rect 2502 1128 2514 1162
rect 2548 1128 2556 1162
rect 2502 1093 2556 1128
rect 2502 1059 2514 1093
rect 2548 1059 2556 1093
rect 2502 1004 2556 1059
rect 2795 1365 2851 1405
rect 2795 1331 2805 1365
rect 2839 1331 2851 1365
rect 2795 1297 2851 1331
rect 2795 1263 2805 1297
rect 2839 1263 2851 1297
rect 2795 1229 2851 1263
rect 2795 1195 2805 1229
rect 2839 1195 2851 1229
rect 2795 1161 2851 1195
rect 2795 1127 2805 1161
rect 2839 1127 2851 1161
rect 2795 1093 2851 1127
rect 2795 1059 2805 1093
rect 2839 1059 2851 1093
rect 2795 1005 2851 1059
rect 2881 1365 2939 1405
rect 2881 1331 2893 1365
rect 2927 1331 2939 1365
rect 2881 1297 2939 1331
rect 2881 1263 2893 1297
rect 2927 1263 2939 1297
rect 2881 1229 2939 1263
rect 2881 1195 2893 1229
rect 2927 1195 2939 1229
rect 2881 1161 2939 1195
rect 2881 1127 2893 1161
rect 2927 1127 2939 1161
rect 2881 1005 2939 1127
rect 2969 1365 3027 1405
rect 2969 1331 2981 1365
rect 3015 1331 3027 1365
rect 2969 1297 3027 1331
rect 2969 1263 2981 1297
rect 3015 1263 3027 1297
rect 2969 1229 3027 1263
rect 2969 1195 2981 1229
rect 3015 1195 3027 1229
rect 2969 1161 3027 1195
rect 2969 1127 2981 1161
rect 3015 1127 3027 1161
rect 2969 1093 3027 1127
rect 2969 1059 2981 1093
rect 3015 1059 3027 1093
rect 2969 1005 3027 1059
rect 3057 1297 3115 1405
rect 3057 1263 3069 1297
rect 3103 1263 3115 1297
rect 3057 1229 3115 1263
rect 3057 1195 3069 1229
rect 3103 1195 3115 1229
rect 3057 1161 3115 1195
rect 3057 1127 3069 1161
rect 3103 1127 3115 1161
rect 3057 1093 3115 1127
rect 3057 1059 3069 1093
rect 3103 1059 3115 1093
rect 3057 1005 3115 1059
rect 3145 1365 3199 1405
rect 3145 1331 3157 1365
rect 3191 1331 3199 1365
rect 3145 1297 3199 1331
rect 3145 1263 3157 1297
rect 3191 1263 3199 1297
rect 3145 1229 3199 1263
rect 3145 1195 3157 1229
rect 3191 1195 3199 1229
rect 3145 1161 3199 1195
rect 3145 1127 3157 1161
rect 3191 1127 3199 1161
rect 3145 1005 3199 1127
rect 3461 1365 3517 1405
rect 3461 1331 3471 1365
rect 3505 1331 3517 1365
rect 3461 1297 3517 1331
rect 3461 1263 3471 1297
rect 3505 1263 3517 1297
rect 3461 1229 3517 1263
rect 3461 1195 3471 1229
rect 3505 1195 3517 1229
rect 3461 1161 3517 1195
rect 3461 1127 3471 1161
rect 3505 1127 3517 1161
rect 3461 1093 3517 1127
rect 3461 1059 3471 1093
rect 3505 1059 3517 1093
rect 3461 1005 3517 1059
rect 3547 1365 3605 1405
rect 3547 1331 3559 1365
rect 3593 1331 3605 1365
rect 3547 1297 3605 1331
rect 3547 1263 3559 1297
rect 3593 1263 3605 1297
rect 3547 1229 3605 1263
rect 3547 1195 3559 1229
rect 3593 1195 3605 1229
rect 3547 1161 3605 1195
rect 3547 1127 3559 1161
rect 3593 1127 3605 1161
rect 3547 1005 3605 1127
rect 3635 1365 3693 1405
rect 3635 1331 3647 1365
rect 3681 1331 3693 1365
rect 3635 1297 3693 1331
rect 3635 1263 3647 1297
rect 3681 1263 3693 1297
rect 3635 1229 3693 1263
rect 3635 1195 3647 1229
rect 3681 1195 3693 1229
rect 3635 1161 3693 1195
rect 3635 1127 3647 1161
rect 3681 1127 3693 1161
rect 3635 1093 3693 1127
rect 3635 1059 3647 1093
rect 3681 1059 3693 1093
rect 3635 1005 3693 1059
rect 3723 1297 3781 1405
rect 3723 1263 3735 1297
rect 3769 1263 3781 1297
rect 3723 1229 3781 1263
rect 3723 1195 3735 1229
rect 3769 1195 3781 1229
rect 3723 1161 3781 1195
rect 3723 1127 3735 1161
rect 3769 1127 3781 1161
rect 3723 1093 3781 1127
rect 3723 1059 3735 1093
rect 3769 1059 3781 1093
rect 3723 1005 3781 1059
rect 3811 1365 3865 1405
rect 3811 1331 3823 1365
rect 3857 1331 3865 1365
rect 3811 1297 3865 1331
rect 3811 1263 3823 1297
rect 3857 1263 3865 1297
rect 3811 1229 3865 1263
rect 3811 1195 3823 1229
rect 3857 1195 3865 1229
rect 3811 1161 3865 1195
rect 3811 1127 3823 1161
rect 3857 1127 3865 1161
rect 3811 1005 3865 1127
<< ndiffc >>
rect 109 300 143 334
rect 303 300 337 334
rect 109 228 143 262
rect 109 160 143 194
rect 205 184 239 218
rect 303 228 337 262
rect 303 160 337 194
rect 109 90 143 124
rect 205 90 239 124
rect 303 90 337 124
rect 566 299 600 333
rect 663 299 697 333
rect 760 299 794 333
rect 566 227 600 261
rect 566 159 600 193
rect 663 174 697 208
rect 760 227 794 261
rect 760 159 794 193
rect 857 183 891 217
rect 954 227 988 261
rect 954 159 988 193
rect 566 89 600 123
rect 760 89 794 123
rect 857 89 891 123
rect 954 89 988 123
rect 1219 300 1253 334
rect 1413 300 1447 334
rect 1219 228 1253 262
rect 1219 160 1253 194
rect 1315 184 1349 218
rect 1413 228 1447 262
rect 1413 160 1447 194
rect 1219 90 1253 124
rect 1315 90 1349 124
rect 1413 90 1447 124
rect 1676 299 1710 333
rect 1773 299 1807 333
rect 1870 299 1904 333
rect 1676 227 1710 261
rect 1676 159 1710 193
rect 1773 174 1807 208
rect 1870 227 1904 261
rect 1870 159 1904 193
rect 1967 183 2001 217
rect 2064 227 2098 261
rect 2064 159 2098 193
rect 1676 89 1710 123
rect 1870 89 1904 123
rect 1967 89 2001 123
rect 2064 89 2098 123
rect 2329 300 2363 334
rect 2523 300 2557 334
rect 2329 228 2363 262
rect 2329 160 2363 194
rect 2425 184 2459 218
rect 2523 228 2557 262
rect 2523 160 2557 194
rect 2329 90 2363 124
rect 2425 90 2459 124
rect 2523 90 2557 124
rect 2786 299 2820 333
rect 2786 227 2820 261
rect 2786 159 2820 193
rect 2883 183 2917 217
rect 2980 227 3014 261
rect 2980 159 3014 193
rect 3077 183 3111 217
rect 3174 227 3208 261
rect 3174 159 3208 193
rect 2786 89 2820 123
rect 2883 89 2917 123
rect 2980 89 3014 123
rect 3077 89 3111 123
rect 3174 89 3208 123
rect 3452 299 3486 333
rect 3452 227 3486 261
rect 3452 159 3486 193
rect 3549 183 3583 217
rect 3646 227 3680 261
rect 3646 159 3680 193
rect 3743 183 3777 217
rect 3840 227 3874 261
rect 3840 159 3874 193
rect 3452 89 3486 123
rect 3549 89 3583 123
rect 3646 89 3680 123
rect 3743 89 3777 123
rect 3840 89 3874 123
<< pdiffc >>
rect 118 1332 152 1366
rect 118 1264 152 1298
rect 118 1196 152 1230
rect 118 1128 152 1162
rect 118 1059 152 1093
rect 206 1332 240 1366
rect 206 1264 240 1298
rect 206 1196 240 1230
rect 206 1128 240 1162
rect 206 1059 240 1093
rect 294 1332 328 1366
rect 294 1264 328 1298
rect 294 1196 328 1230
rect 294 1128 328 1162
rect 294 1059 328 1093
rect 585 1332 619 1366
rect 585 1264 619 1298
rect 585 1196 619 1230
rect 585 1128 619 1162
rect 585 1059 619 1093
rect 673 1332 707 1366
rect 673 1264 707 1298
rect 673 1196 707 1230
rect 673 1128 707 1162
rect 673 1059 707 1093
rect 761 1332 795 1366
rect 761 1264 795 1298
rect 761 1196 795 1230
rect 761 1128 795 1162
rect 849 1332 883 1366
rect 849 1264 883 1298
rect 849 1196 883 1230
rect 849 1128 883 1162
rect 849 1059 883 1093
rect 937 1332 971 1366
rect 937 1264 971 1298
rect 937 1196 971 1230
rect 937 1128 971 1162
rect 1228 1332 1262 1366
rect 1228 1264 1262 1298
rect 1228 1196 1262 1230
rect 1228 1128 1262 1162
rect 1228 1059 1262 1093
rect 1316 1332 1350 1366
rect 1316 1264 1350 1298
rect 1316 1196 1350 1230
rect 1316 1128 1350 1162
rect 1316 1059 1350 1093
rect 1404 1332 1438 1366
rect 1404 1264 1438 1298
rect 1404 1196 1438 1230
rect 1404 1128 1438 1162
rect 1404 1059 1438 1093
rect 1695 1332 1729 1366
rect 1695 1264 1729 1298
rect 1695 1196 1729 1230
rect 1695 1128 1729 1162
rect 1695 1059 1729 1093
rect 1783 1332 1817 1366
rect 1783 1264 1817 1298
rect 1783 1196 1817 1230
rect 1783 1128 1817 1162
rect 1783 1059 1817 1093
rect 1871 1332 1905 1366
rect 1871 1264 1905 1298
rect 1871 1196 1905 1230
rect 1871 1128 1905 1162
rect 1959 1332 1993 1366
rect 1959 1264 1993 1298
rect 1959 1196 1993 1230
rect 1959 1128 1993 1162
rect 1959 1059 1993 1093
rect 2047 1332 2081 1366
rect 2047 1264 2081 1298
rect 2047 1196 2081 1230
rect 2047 1128 2081 1162
rect 2338 1332 2372 1366
rect 2338 1264 2372 1298
rect 2338 1196 2372 1230
rect 2338 1128 2372 1162
rect 2338 1059 2372 1093
rect 2426 1332 2460 1366
rect 2426 1264 2460 1298
rect 2426 1196 2460 1230
rect 2426 1128 2460 1162
rect 2426 1059 2460 1093
rect 2514 1332 2548 1366
rect 2514 1264 2548 1298
rect 2514 1196 2548 1230
rect 2514 1128 2548 1162
rect 2514 1059 2548 1093
rect 2805 1331 2839 1365
rect 2805 1263 2839 1297
rect 2805 1195 2839 1229
rect 2805 1127 2839 1161
rect 2805 1059 2839 1093
rect 2893 1331 2927 1365
rect 2893 1263 2927 1297
rect 2893 1195 2927 1229
rect 2893 1127 2927 1161
rect 2981 1331 3015 1365
rect 2981 1263 3015 1297
rect 2981 1195 3015 1229
rect 2981 1127 3015 1161
rect 2981 1059 3015 1093
rect 3069 1263 3103 1297
rect 3069 1195 3103 1229
rect 3069 1127 3103 1161
rect 3069 1059 3103 1093
rect 3157 1331 3191 1365
rect 3157 1263 3191 1297
rect 3157 1195 3191 1229
rect 3157 1127 3191 1161
rect 3471 1331 3505 1365
rect 3471 1263 3505 1297
rect 3471 1195 3505 1229
rect 3471 1127 3505 1161
rect 3471 1059 3505 1093
rect 3559 1331 3593 1365
rect 3559 1263 3593 1297
rect 3559 1195 3593 1229
rect 3559 1127 3593 1161
rect 3647 1331 3681 1365
rect 3647 1263 3681 1297
rect 3647 1195 3681 1229
rect 3647 1127 3681 1161
rect 3647 1059 3681 1093
rect 3735 1263 3769 1297
rect 3735 1195 3769 1229
rect 3735 1127 3769 1161
rect 3735 1059 3769 1093
rect 3823 1331 3857 1365
rect 3823 1263 3857 1297
rect 3823 1195 3857 1229
rect 3823 1127 3857 1161
<< psubdiff >>
rect -34 482 4030 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 410 461 478 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 410 427 427 461
rect 461 427 478 461
rect 1076 461 1144 482
rect -34 313 34 353
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 410 313 478 353
rect 1076 427 1093 461
rect 1127 427 1144 461
rect 1520 461 1588 482
rect 1076 387 1144 427
rect 1076 353 1093 387
rect 1127 353 1144 387
rect 1520 427 1537 461
rect 1571 427 1588 461
rect 2186 461 2254 482
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect -34 17 34 57
rect 410 57 427 91
rect 461 57 478 91
rect 1076 313 1144 353
rect 1520 387 1588 427
rect 1520 353 1537 387
rect 1571 353 1588 387
rect 1076 279 1093 313
rect 1127 279 1144 313
rect 1076 239 1144 279
rect 1076 205 1093 239
rect 1127 205 1144 239
rect 1076 165 1144 205
rect 1076 131 1093 165
rect 1127 131 1144 165
rect 1076 91 1144 131
rect 410 17 478 57
rect 1076 57 1093 91
rect 1127 57 1144 91
rect 1520 313 1588 353
rect 2186 427 2203 461
rect 2237 427 2254 461
rect 2630 461 2698 482
rect 2186 387 2254 427
rect 2186 353 2203 387
rect 2237 353 2254 387
rect 2630 427 2647 461
rect 2681 427 2698 461
rect 3296 461 3364 482
rect 1520 279 1537 313
rect 1571 279 1588 313
rect 1520 239 1588 279
rect 1520 205 1537 239
rect 1571 205 1588 239
rect 1520 165 1588 205
rect 1520 131 1537 165
rect 1571 131 1588 165
rect 1520 91 1588 131
rect 1076 17 1144 57
rect 1520 57 1537 91
rect 1571 57 1588 91
rect 2186 313 2254 353
rect 2630 387 2698 427
rect 2630 353 2647 387
rect 2681 353 2698 387
rect 2186 279 2203 313
rect 2237 279 2254 313
rect 2186 239 2254 279
rect 2186 205 2203 239
rect 2237 205 2254 239
rect 2186 165 2254 205
rect 2186 131 2203 165
rect 2237 131 2254 165
rect 2186 91 2254 131
rect 1520 17 1588 57
rect 2186 57 2203 91
rect 2237 57 2254 91
rect 2630 313 2698 353
rect 3296 427 3313 461
rect 3347 427 3364 461
rect 3962 461 4030 482
rect 3296 387 3364 427
rect 3296 353 3313 387
rect 3347 353 3364 387
rect 2630 279 2647 313
rect 2681 279 2698 313
rect 2630 239 2698 279
rect 2630 205 2647 239
rect 2681 205 2698 239
rect 2630 165 2698 205
rect 2630 131 2647 165
rect 2681 131 2698 165
rect 2630 91 2698 131
rect 2186 17 2254 57
rect 2630 57 2647 91
rect 2681 57 2698 91
rect 3296 313 3364 353
rect 3962 427 3979 461
rect 4013 427 4030 461
rect 3962 387 4030 427
rect 3962 353 3979 387
rect 4013 353 4030 387
rect 3296 279 3313 313
rect 3347 279 3364 313
rect 3296 239 3364 279
rect 3296 205 3313 239
rect 3347 205 3364 239
rect 3296 165 3364 205
rect 3296 131 3313 165
rect 3347 131 3364 165
rect 3296 91 3364 131
rect 2630 17 2698 57
rect 3296 57 3313 91
rect 3347 57 3364 91
rect 3962 313 4030 353
rect 3962 279 3979 313
rect 4013 279 4030 313
rect 3962 239 4030 279
rect 3962 205 3979 239
rect 4013 205 4030 239
rect 3962 165 4030 205
rect 3962 131 3979 165
rect 4013 131 4030 165
rect 3962 91 4030 131
rect 3296 17 3364 57
rect 3962 57 3979 91
rect 4013 57 4030 91
rect 3962 17 4030 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 4030 17
rect -34 -34 4030 -17
<< nsubdiff >>
rect -34 1497 4030 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 4030 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 410 1423 478 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 1076 1423 1144 1463
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 410 979 478 1019
rect 1076 1389 1093 1423
rect 1127 1389 1144 1423
rect 1520 1423 1588 1463
rect 1076 1349 1144 1389
rect 1076 1315 1093 1349
rect 1127 1315 1144 1349
rect 1076 1275 1144 1315
rect 1076 1241 1093 1275
rect 1127 1241 1144 1275
rect 1076 1201 1144 1241
rect 1076 1167 1093 1201
rect 1127 1167 1144 1201
rect 1076 1127 1144 1167
rect 1076 1093 1093 1127
rect 1127 1093 1144 1127
rect 1076 1053 1144 1093
rect 1076 1019 1093 1053
rect 1127 1019 1144 1053
rect 410 945 427 979
rect 461 945 478 979
rect -34 871 -17 905
rect 17 884 34 905
rect 410 905 478 945
rect 1076 979 1144 1019
rect 1520 1389 1537 1423
rect 1571 1389 1588 1423
rect 2186 1423 2254 1463
rect 1520 1349 1588 1389
rect 1520 1315 1537 1349
rect 1571 1315 1588 1349
rect 1520 1275 1588 1315
rect 1520 1241 1537 1275
rect 1571 1241 1588 1275
rect 1520 1201 1588 1241
rect 1520 1167 1537 1201
rect 1571 1167 1588 1201
rect 1520 1127 1588 1167
rect 1520 1093 1537 1127
rect 1571 1093 1588 1127
rect 1520 1053 1588 1093
rect 1520 1019 1537 1053
rect 1571 1019 1588 1053
rect 1076 945 1093 979
rect 1127 945 1144 979
rect 410 884 427 905
rect 17 871 427 884
rect 461 884 478 905
rect 1076 905 1144 945
rect 1520 979 1588 1019
rect 2186 1389 2203 1423
rect 2237 1389 2254 1423
rect 2630 1423 2698 1463
rect 2186 1349 2254 1389
rect 2186 1315 2203 1349
rect 2237 1315 2254 1349
rect 2186 1275 2254 1315
rect 2186 1241 2203 1275
rect 2237 1241 2254 1275
rect 2186 1201 2254 1241
rect 2186 1167 2203 1201
rect 2237 1167 2254 1201
rect 2186 1127 2254 1167
rect 2186 1093 2203 1127
rect 2237 1093 2254 1127
rect 2186 1053 2254 1093
rect 2186 1019 2203 1053
rect 2237 1019 2254 1053
rect 1520 945 1537 979
rect 1571 945 1588 979
rect 1076 884 1093 905
rect 461 871 1093 884
rect 1127 884 1144 905
rect 1520 905 1588 945
rect 2186 979 2254 1019
rect 2630 1389 2647 1423
rect 2681 1389 2698 1423
rect 3296 1423 3364 1463
rect 2630 1349 2698 1389
rect 2630 1315 2647 1349
rect 2681 1315 2698 1349
rect 2630 1275 2698 1315
rect 2630 1241 2647 1275
rect 2681 1241 2698 1275
rect 2630 1201 2698 1241
rect 2630 1167 2647 1201
rect 2681 1167 2698 1201
rect 2630 1127 2698 1167
rect 2630 1093 2647 1127
rect 2681 1093 2698 1127
rect 2630 1053 2698 1093
rect 2630 1019 2647 1053
rect 2681 1019 2698 1053
rect 2186 945 2203 979
rect 2237 945 2254 979
rect 1520 884 1537 905
rect 1127 871 1537 884
rect 1571 884 1588 905
rect 2186 905 2254 945
rect 2630 979 2698 1019
rect 3296 1389 3313 1423
rect 3347 1389 3364 1423
rect 3962 1423 4030 1463
rect 3296 1349 3364 1389
rect 3296 1315 3313 1349
rect 3347 1315 3364 1349
rect 3296 1275 3364 1315
rect 3296 1241 3313 1275
rect 3347 1241 3364 1275
rect 3296 1201 3364 1241
rect 3296 1167 3313 1201
rect 3347 1167 3364 1201
rect 3296 1127 3364 1167
rect 3296 1093 3313 1127
rect 3347 1093 3364 1127
rect 3296 1053 3364 1093
rect 3296 1019 3313 1053
rect 3347 1019 3364 1053
rect 2630 945 2647 979
rect 2681 945 2698 979
rect 2186 884 2203 905
rect 1571 871 2203 884
rect 2237 884 2254 905
rect 2630 905 2698 945
rect 3296 979 3364 1019
rect 3962 1389 3979 1423
rect 4013 1389 4030 1423
rect 3962 1349 4030 1389
rect 3962 1315 3979 1349
rect 4013 1315 4030 1349
rect 3962 1275 4030 1315
rect 3962 1241 3979 1275
rect 4013 1241 4030 1275
rect 3962 1201 4030 1241
rect 3962 1167 3979 1201
rect 4013 1167 4030 1201
rect 3962 1127 4030 1167
rect 3962 1093 3979 1127
rect 4013 1093 4030 1127
rect 3962 1053 4030 1093
rect 3962 1019 3979 1053
rect 4013 1019 4030 1053
rect 3296 945 3313 979
rect 3347 945 3364 979
rect 2630 884 2647 905
rect 2237 871 2647 884
rect 2681 884 2698 905
rect 3296 905 3364 945
rect 3962 979 4030 1019
rect 3962 945 3979 979
rect 4013 945 4030 979
rect 3296 884 3313 905
rect 2681 871 3313 884
rect 3347 884 3364 905
rect 3962 905 4030 945
rect 3962 884 3979 905
rect 3347 871 3979 884
rect 4013 871 4030 905
rect -34 822 4030 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 427 427 461 461
rect 427 353 461 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1093 427 1127 461
rect 1093 353 1127 387
rect 1537 427 1571 461
rect 427 279 461 313
rect 427 205 461 239
rect 427 131 461 165
rect 427 57 461 91
rect 1537 353 1571 387
rect 1093 279 1127 313
rect 1093 205 1127 239
rect 1093 131 1127 165
rect 1093 57 1127 91
rect 2203 427 2237 461
rect 2203 353 2237 387
rect 2647 427 2681 461
rect 1537 279 1571 313
rect 1537 205 1571 239
rect 1537 131 1571 165
rect 1537 57 1571 91
rect 2647 353 2681 387
rect 2203 279 2237 313
rect 2203 205 2237 239
rect 2203 131 2237 165
rect 2203 57 2237 91
rect 3313 427 3347 461
rect 3313 353 3347 387
rect 2647 279 2681 313
rect 2647 205 2681 239
rect 2647 131 2681 165
rect 2647 57 2681 91
rect 3979 427 4013 461
rect 3979 353 4013 387
rect 3313 279 3347 313
rect 3313 205 3347 239
rect 3313 131 3347 165
rect 3313 57 3347 91
rect 3979 279 4013 313
rect 3979 205 4013 239
rect 3979 131 4013 165
rect 3979 57 4013 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 427 1389 461 1423
rect 427 1315 461 1349
rect 427 1241 461 1275
rect 427 1167 461 1201
rect 427 1093 461 1127
rect 427 1019 461 1053
rect -17 945 17 979
rect 1093 1389 1127 1423
rect 1093 1315 1127 1349
rect 1093 1241 1127 1275
rect 1093 1167 1127 1201
rect 1093 1093 1127 1127
rect 1093 1019 1127 1053
rect 427 945 461 979
rect -17 871 17 905
rect 1537 1389 1571 1423
rect 1537 1315 1571 1349
rect 1537 1241 1571 1275
rect 1537 1167 1571 1201
rect 1537 1093 1571 1127
rect 1537 1019 1571 1053
rect 1093 945 1127 979
rect 427 871 461 905
rect 2203 1389 2237 1423
rect 2203 1315 2237 1349
rect 2203 1241 2237 1275
rect 2203 1167 2237 1201
rect 2203 1093 2237 1127
rect 2203 1019 2237 1053
rect 1537 945 1571 979
rect 1093 871 1127 905
rect 2647 1389 2681 1423
rect 2647 1315 2681 1349
rect 2647 1241 2681 1275
rect 2647 1167 2681 1201
rect 2647 1093 2681 1127
rect 2647 1019 2681 1053
rect 2203 945 2237 979
rect 1537 871 1571 905
rect 3313 1389 3347 1423
rect 3313 1315 3347 1349
rect 3313 1241 3347 1275
rect 3313 1167 3347 1201
rect 3313 1093 3347 1127
rect 3313 1019 3347 1053
rect 2647 945 2681 979
rect 2203 871 2237 905
rect 3979 1389 4013 1423
rect 3979 1315 4013 1349
rect 3979 1241 4013 1275
rect 3979 1167 4013 1201
rect 3979 1093 4013 1127
rect 3979 1019 4013 1053
rect 3313 945 3347 979
rect 2647 871 2681 905
rect 3979 945 4013 979
rect 3313 871 3347 905
rect 3979 871 4013 905
<< poly >>
rect 164 1404 194 1430
rect 252 1404 282 1430
rect 631 1404 661 1430
rect 719 1404 749 1430
rect 807 1404 837 1430
rect 895 1404 925 1430
rect 164 973 194 1004
rect 252 973 282 1004
rect 121 957 282 973
rect 121 923 131 957
rect 165 943 282 957
rect 1274 1404 1304 1430
rect 1362 1404 1392 1430
rect 165 923 175 943
rect 121 907 175 923
rect 631 973 661 1004
rect 719 973 749 1004
rect 807 973 837 1004
rect 895 973 925 1004
rect 631 957 749 973
rect 631 943 649 957
rect 639 923 649 943
rect 683 943 749 957
rect 793 957 925 973
rect 683 923 693 943
rect 639 907 693 923
rect 793 923 803 957
rect 837 943 925 957
rect 1741 1404 1771 1430
rect 1829 1404 1859 1430
rect 1917 1404 1947 1430
rect 2005 1404 2035 1430
rect 1274 973 1304 1004
rect 1362 973 1392 1004
rect 837 923 847 943
rect 793 907 847 923
rect 1231 957 1392 973
rect 1231 923 1241 957
rect 1275 943 1392 957
rect 2384 1404 2414 1430
rect 2472 1404 2502 1430
rect 1275 923 1285 943
rect 1231 907 1285 923
rect 1741 973 1771 1004
rect 1829 973 1859 1004
rect 1917 973 1947 1004
rect 2005 973 2035 1004
rect 1741 957 1859 973
rect 1741 943 1759 957
rect 1749 923 1759 943
rect 1793 943 1859 957
rect 1903 957 2035 973
rect 1793 923 1803 943
rect 1749 907 1803 923
rect 1903 923 1913 957
rect 1947 943 2035 957
rect 2851 1405 2881 1431
rect 2939 1405 2969 1431
rect 3027 1405 3057 1431
rect 3115 1405 3145 1431
rect 2384 973 2414 1004
rect 2472 973 2502 1004
rect 1947 923 1957 943
rect 1903 907 1957 923
rect 2341 957 2502 973
rect 2341 923 2351 957
rect 2385 943 2502 957
rect 3517 1405 3547 1431
rect 3605 1405 3635 1431
rect 3693 1405 3723 1431
rect 3781 1405 3811 1431
rect 2851 974 2881 1005
rect 2939 974 2969 1005
rect 3027 974 3057 1005
rect 3115 974 3145 1005
rect 2385 923 2395 943
rect 2341 907 2395 923
rect 2828 958 2969 974
rect 2828 924 2838 958
rect 2872 944 2969 958
rect 3014 958 3145 974
rect 2872 924 2882 944
rect 2828 908 2882 924
rect 3014 924 3024 958
rect 3058 944 3145 958
rect 3517 974 3547 1005
rect 3605 974 3635 1005
rect 3693 974 3723 1005
rect 3781 974 3811 1005
rect 3058 924 3068 944
rect 3014 908 3068 924
rect 3494 958 3635 974
rect 3494 924 3504 958
rect 3538 944 3635 958
rect 3680 958 3811 974
rect 3538 924 3548 944
rect 3494 908 3548 924
rect 3680 924 3690 958
rect 3724 944 3811 958
rect 3724 924 3734 944
rect 3680 908 3734 924
rect 121 434 175 450
rect 121 400 131 434
rect 165 413 175 434
rect 165 400 185 413
rect 121 384 185 400
rect 155 350 185 384
rect 639 433 693 449
rect 639 413 649 433
rect 612 399 649 413
rect 683 399 693 433
rect 612 383 693 399
rect 787 433 841 449
rect 787 399 797 433
rect 831 399 841 433
rect 787 383 841 399
rect 612 349 642 383
rect 806 349 836 383
rect 1231 434 1285 450
rect 1231 400 1241 434
rect 1275 413 1285 434
rect 1275 400 1295 413
rect 1231 384 1295 400
rect 1265 350 1295 384
rect 1749 433 1803 449
rect 1749 413 1759 433
rect 1722 399 1759 413
rect 1793 399 1803 433
rect 1722 383 1803 399
rect 1897 433 1951 449
rect 1897 399 1907 433
rect 1941 399 1951 433
rect 1897 383 1951 399
rect 1722 349 1752 383
rect 1916 349 1946 383
rect 2341 434 2395 450
rect 2341 400 2351 434
rect 2385 413 2395 434
rect 2385 400 2405 413
rect 2341 384 2405 400
rect 2375 350 2405 384
rect 2859 433 2913 449
rect 2859 413 2869 433
rect 2832 399 2869 413
rect 2903 399 2913 433
rect 2832 383 2913 399
rect 3007 433 3061 449
rect 3007 399 3017 433
rect 3051 399 3061 433
rect 3007 383 3061 399
rect 3525 433 3579 449
rect 3525 413 3535 433
rect 2832 349 2862 383
rect 3026 349 3056 383
rect 3498 399 3535 413
rect 3569 399 3579 433
rect 3498 383 3579 399
rect 3673 433 3727 449
rect 3673 399 3683 433
rect 3717 399 3727 433
rect 3673 383 3727 399
rect 3498 349 3528 383
rect 3692 349 3722 383
<< polycont >>
rect 131 923 165 957
rect 649 923 683 957
rect 803 923 837 957
rect 1241 923 1275 957
rect 1759 923 1793 957
rect 1913 923 1947 957
rect 2351 923 2385 957
rect 2838 924 2872 958
rect 3024 924 3058 958
rect 3504 924 3538 958
rect 3690 924 3724 958
rect 131 400 165 434
rect 649 399 683 433
rect 797 399 831 433
rect 1241 400 1275 434
rect 1759 399 1793 433
rect 1907 399 1941 433
rect 2351 400 2385 434
rect 2869 399 2903 433
rect 3017 399 3051 433
rect 3535 399 3569 433
rect 3683 399 3717 433
<< locali >>
rect -34 1497 4030 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 4030 1497
rect -34 1446 4030 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 118 1366 152 1446
rect 118 1298 152 1332
rect 118 1230 152 1264
rect 118 1162 152 1196
rect 118 1093 152 1128
rect 118 1037 152 1059
rect 206 1366 240 1404
rect 206 1298 240 1332
rect 206 1230 240 1264
rect 206 1162 240 1196
rect 206 1093 240 1128
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 131 957 165 973
rect 131 831 165 923
rect 206 933 240 1059
rect 294 1366 328 1446
rect 294 1298 328 1332
rect 294 1230 328 1264
rect 294 1162 328 1196
rect 294 1093 328 1128
rect 294 1037 328 1059
rect 410 1423 478 1446
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect 585 1366 619 1446
rect 585 1298 619 1332
rect 585 1230 619 1264
rect 585 1162 619 1196
rect 585 1093 619 1128
rect 585 1027 619 1059
rect 673 1366 707 1404
rect 673 1298 707 1332
rect 673 1230 707 1264
rect 673 1162 707 1196
rect 673 1093 707 1128
rect 761 1366 795 1446
rect 761 1298 795 1332
rect 761 1230 795 1264
rect 761 1162 795 1196
rect 761 1111 795 1128
rect 849 1366 883 1404
rect 849 1298 883 1332
rect 849 1230 883 1264
rect 849 1162 883 1196
rect 673 1057 707 1059
rect 849 1093 883 1128
rect 937 1366 971 1446
rect 937 1298 971 1332
rect 937 1230 971 1264
rect 937 1162 971 1196
rect 937 1111 971 1128
rect 1076 1423 1144 1446
rect 1076 1389 1093 1423
rect 1127 1389 1144 1423
rect 1076 1349 1144 1389
rect 1076 1315 1093 1349
rect 1127 1315 1144 1349
rect 1076 1275 1144 1315
rect 1076 1241 1093 1275
rect 1127 1241 1144 1275
rect 1076 1201 1144 1241
rect 1076 1167 1093 1201
rect 1127 1167 1144 1201
rect 1076 1127 1144 1167
rect 849 1057 883 1059
rect 1076 1093 1093 1127
rect 1127 1093 1144 1127
rect 673 1023 979 1057
rect 410 979 478 1019
rect 410 945 427 979
rect 461 945 478 979
rect 206 899 313 933
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 131 434 165 797
rect 279 757 313 899
rect 410 905 478 945
rect 410 871 427 905
rect 461 871 478 905
rect 410 822 478 871
rect 649 957 683 973
rect 803 957 837 973
rect 279 433 313 723
rect 649 757 683 923
rect 131 384 165 400
rect 205 399 313 433
rect 410 461 478 544
rect 410 427 427 461
rect 461 427 478 461
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect -34 34 34 57
rect 109 334 143 350
rect 109 262 143 300
rect 109 194 143 228
rect 205 218 239 399
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect 649 433 683 723
rect 649 383 683 399
rect 797 923 803 942
rect 797 907 837 923
rect 797 609 831 907
rect 797 433 831 575
rect 797 383 831 399
rect 945 683 979 1023
rect 1076 1053 1144 1093
rect 1076 1019 1093 1053
rect 1127 1019 1144 1053
rect 1228 1366 1262 1446
rect 1228 1298 1262 1332
rect 1228 1230 1262 1264
rect 1228 1162 1262 1196
rect 1228 1093 1262 1128
rect 1228 1037 1262 1059
rect 1316 1366 1350 1404
rect 1316 1298 1350 1332
rect 1316 1230 1350 1264
rect 1316 1162 1350 1196
rect 1316 1093 1350 1128
rect 1076 979 1144 1019
rect 1076 945 1093 979
rect 1127 945 1144 979
rect 1076 905 1144 945
rect 1076 871 1093 905
rect 1127 871 1144 905
rect 1076 822 1144 871
rect 1241 957 1275 973
rect 205 168 239 184
rect 303 334 337 350
rect 303 262 337 300
rect 303 194 337 228
rect 109 124 143 160
rect 303 124 337 160
rect 143 90 205 124
rect 239 90 303 124
rect 109 34 143 90
rect 206 34 240 90
rect 303 34 337 90
rect 410 313 478 353
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect 410 57 427 91
rect 461 57 478 91
rect 566 333 600 349
rect 760 333 794 349
rect 945 348 979 649
rect 1241 683 1275 923
rect 1316 933 1350 1059
rect 1404 1366 1438 1446
rect 1404 1298 1438 1332
rect 1404 1230 1438 1264
rect 1404 1162 1438 1196
rect 1404 1093 1438 1128
rect 1404 1037 1438 1059
rect 1520 1423 1588 1446
rect 1520 1389 1537 1423
rect 1571 1389 1588 1423
rect 1520 1349 1588 1389
rect 1520 1315 1537 1349
rect 1571 1315 1588 1349
rect 1520 1275 1588 1315
rect 1520 1241 1537 1275
rect 1571 1241 1588 1275
rect 1520 1201 1588 1241
rect 1520 1167 1537 1201
rect 1571 1167 1588 1201
rect 1520 1127 1588 1167
rect 1520 1093 1537 1127
rect 1571 1093 1588 1127
rect 1520 1053 1588 1093
rect 1520 1019 1537 1053
rect 1571 1019 1588 1053
rect 1695 1366 1729 1446
rect 1695 1298 1729 1332
rect 1695 1230 1729 1264
rect 1695 1162 1729 1196
rect 1695 1093 1729 1128
rect 1695 1027 1729 1059
rect 1783 1366 1817 1404
rect 1783 1298 1817 1332
rect 1783 1230 1817 1264
rect 1783 1162 1817 1196
rect 1783 1093 1817 1128
rect 1871 1366 1905 1446
rect 1871 1298 1905 1332
rect 1871 1230 1905 1264
rect 1871 1162 1905 1196
rect 1871 1111 1905 1128
rect 1959 1366 1993 1404
rect 1959 1298 1993 1332
rect 1959 1230 1993 1264
rect 1959 1162 1993 1196
rect 1783 1057 1817 1059
rect 1959 1093 1993 1128
rect 2047 1366 2081 1446
rect 2047 1298 2081 1332
rect 2047 1230 2081 1264
rect 2047 1162 2081 1196
rect 2047 1111 2081 1128
rect 2186 1423 2254 1446
rect 2186 1389 2203 1423
rect 2237 1389 2254 1423
rect 2186 1349 2254 1389
rect 2186 1315 2203 1349
rect 2237 1315 2254 1349
rect 2186 1275 2254 1315
rect 2186 1241 2203 1275
rect 2237 1241 2254 1275
rect 2186 1201 2254 1241
rect 2186 1167 2203 1201
rect 2237 1167 2254 1201
rect 2186 1127 2254 1167
rect 1959 1057 1993 1059
rect 2186 1093 2203 1127
rect 2237 1093 2254 1127
rect 1783 1023 2089 1057
rect 1520 979 1588 1019
rect 1520 945 1537 979
rect 1571 945 1588 979
rect 1316 899 1423 933
rect 600 299 663 333
rect 697 299 760 333
rect 566 261 600 299
rect 566 193 600 227
rect 760 261 794 299
rect 566 123 600 159
rect 566 73 600 89
rect 663 208 697 224
rect 410 34 478 57
rect 663 34 697 174
rect 760 193 794 227
rect 857 314 979 348
rect 1076 461 1144 544
rect 1076 427 1093 461
rect 1127 427 1144 461
rect 1076 387 1144 427
rect 1076 353 1093 387
rect 1127 353 1144 387
rect 1241 434 1275 649
rect 1389 757 1423 899
rect 1520 905 1588 945
rect 1520 871 1537 905
rect 1571 871 1588 905
rect 1520 822 1588 871
rect 1759 957 1793 973
rect 1913 957 1947 973
rect 1389 433 1423 723
rect 1759 609 1793 923
rect 1241 384 1275 400
rect 1315 399 1423 433
rect 1520 461 1588 544
rect 1520 427 1537 461
rect 1571 427 1588 461
rect 857 217 891 314
rect 1076 313 1144 353
rect 1076 279 1093 313
rect 1127 279 1144 313
rect 857 167 891 183
rect 954 261 988 277
rect 954 193 988 227
rect 760 123 794 159
rect 954 123 988 159
rect 794 89 857 123
rect 891 89 954 123
rect 760 73 794 89
rect 954 73 988 89
rect 1076 239 1144 279
rect 1076 205 1093 239
rect 1127 205 1144 239
rect 1076 165 1144 205
rect 1076 131 1093 165
rect 1127 131 1144 165
rect 1076 91 1144 131
rect 1076 57 1093 91
rect 1127 57 1144 91
rect 1076 34 1144 57
rect 1219 334 1253 350
rect 1219 262 1253 300
rect 1219 194 1253 228
rect 1315 218 1349 399
rect 1520 387 1588 427
rect 1520 353 1537 387
rect 1571 353 1588 387
rect 1759 433 1793 575
rect 1759 383 1793 399
rect 1907 923 1913 942
rect 1907 907 1947 923
rect 1907 831 1941 907
rect 1907 433 1941 797
rect 1907 383 1941 399
rect 2055 683 2089 1023
rect 2186 1053 2254 1093
rect 2186 1019 2203 1053
rect 2237 1019 2254 1053
rect 2338 1366 2372 1446
rect 2338 1298 2372 1332
rect 2338 1230 2372 1264
rect 2338 1162 2372 1196
rect 2338 1093 2372 1128
rect 2338 1037 2372 1059
rect 2426 1366 2460 1404
rect 2426 1298 2460 1332
rect 2426 1230 2460 1264
rect 2426 1162 2460 1196
rect 2426 1093 2460 1128
rect 2186 979 2254 1019
rect 2186 945 2203 979
rect 2237 945 2254 979
rect 2186 905 2254 945
rect 2186 871 2203 905
rect 2237 871 2254 905
rect 2186 822 2254 871
rect 2351 957 2385 973
rect 1315 168 1349 184
rect 1413 334 1447 350
rect 1413 262 1447 300
rect 1413 194 1447 228
rect 1219 124 1253 160
rect 1413 124 1447 160
rect 1253 90 1315 124
rect 1349 90 1413 124
rect 1219 34 1253 90
rect 1316 34 1350 90
rect 1413 34 1447 90
rect 1520 313 1588 353
rect 1520 279 1537 313
rect 1571 279 1588 313
rect 1520 239 1588 279
rect 1520 205 1537 239
rect 1571 205 1588 239
rect 1520 165 1588 205
rect 1520 131 1537 165
rect 1571 131 1588 165
rect 1520 91 1588 131
rect 1520 57 1537 91
rect 1571 57 1588 91
rect 1676 333 1710 349
rect 1870 333 1904 349
rect 2055 348 2089 649
rect 2351 683 2385 923
rect 2426 933 2460 1059
rect 2514 1366 2548 1446
rect 2514 1298 2548 1332
rect 2514 1230 2548 1264
rect 2514 1162 2548 1196
rect 2514 1093 2548 1128
rect 2514 1037 2548 1059
rect 2630 1423 2698 1446
rect 2630 1389 2647 1423
rect 2681 1389 2698 1423
rect 2630 1349 2698 1389
rect 2630 1315 2647 1349
rect 2681 1315 2698 1349
rect 2630 1275 2698 1315
rect 2630 1241 2647 1275
rect 2681 1241 2698 1275
rect 2630 1201 2698 1241
rect 2630 1167 2647 1201
rect 2681 1167 2698 1201
rect 2630 1127 2698 1167
rect 2630 1093 2647 1127
rect 2681 1093 2698 1127
rect 2630 1053 2698 1093
rect 2630 1019 2647 1053
rect 2681 1019 2698 1053
rect 2805 1365 2839 1405
rect 2805 1297 2839 1331
rect 2805 1229 2839 1263
rect 2805 1161 2839 1195
rect 2805 1093 2839 1127
rect 2893 1365 2927 1446
rect 3296 1423 3364 1446
rect 2893 1297 2927 1331
rect 2893 1229 2927 1263
rect 2893 1161 2927 1195
rect 2893 1111 2927 1127
rect 2981 1365 3191 1399
rect 2981 1297 3015 1331
rect 2981 1229 3015 1263
rect 2981 1161 3015 1195
rect 2981 1093 3015 1127
rect 2805 1025 3015 1059
rect 3069 1297 3103 1313
rect 3069 1229 3103 1263
rect 3069 1161 3103 1195
rect 3069 1093 3103 1127
rect 3157 1297 3191 1331
rect 3157 1229 3191 1263
rect 3157 1161 3191 1195
rect 3157 1111 3191 1127
rect 3296 1389 3313 1423
rect 3347 1389 3364 1423
rect 3296 1349 3364 1389
rect 3296 1315 3313 1349
rect 3347 1315 3364 1349
rect 3296 1275 3364 1315
rect 3296 1241 3313 1275
rect 3347 1241 3364 1275
rect 3296 1201 3364 1241
rect 3296 1167 3313 1201
rect 3347 1167 3364 1201
rect 3296 1127 3364 1167
rect 3296 1093 3313 1127
rect 3347 1093 3364 1127
rect 3069 1025 3199 1059
rect 2630 979 2698 1019
rect 2630 945 2647 979
rect 2681 945 2698 979
rect 2426 899 2533 933
rect 1710 299 1773 333
rect 1807 299 1870 333
rect 1676 261 1710 299
rect 1676 193 1710 227
rect 1870 261 1904 299
rect 1676 123 1710 159
rect 1676 73 1710 89
rect 1773 208 1807 224
rect 1520 34 1588 57
rect 1773 34 1807 174
rect 1870 193 1904 227
rect 1967 314 2089 348
rect 2186 461 2254 544
rect 2186 427 2203 461
rect 2237 427 2254 461
rect 2186 387 2254 427
rect 2186 353 2203 387
rect 2237 353 2254 387
rect 2351 434 2385 649
rect 2499 831 2533 899
rect 2630 905 2698 945
rect 2838 958 2872 974
rect 3024 958 3058 974
rect 2872 924 2903 942
rect 2838 908 2903 924
rect 2630 871 2647 905
rect 2681 871 2698 905
rect 2630 822 2698 871
rect 2499 433 2533 797
rect 2869 757 2903 908
rect 2351 384 2385 400
rect 2425 399 2533 433
rect 2630 461 2698 544
rect 2630 427 2647 461
rect 2681 427 2698 461
rect 1967 217 2001 314
rect 2186 313 2254 353
rect 2186 279 2203 313
rect 2237 279 2254 313
rect 1967 167 2001 183
rect 2064 261 2098 277
rect 2064 193 2098 227
rect 1870 123 1904 159
rect 2064 123 2098 159
rect 1904 89 1967 123
rect 2001 89 2064 123
rect 1870 73 1904 89
rect 2064 73 2098 89
rect 2186 239 2254 279
rect 2186 205 2203 239
rect 2237 205 2254 239
rect 2186 165 2254 205
rect 2186 131 2203 165
rect 2237 131 2254 165
rect 2186 91 2254 131
rect 2186 57 2203 91
rect 2237 57 2254 91
rect 2186 34 2254 57
rect 2329 334 2363 350
rect 2329 262 2363 300
rect 2329 194 2363 228
rect 2425 218 2459 399
rect 2630 387 2698 427
rect 2630 353 2647 387
rect 2681 353 2698 387
rect 2869 433 2903 723
rect 2869 383 2903 399
rect 3017 924 3024 942
rect 3017 908 3058 924
rect 3017 757 3051 908
rect 3017 433 3051 723
rect 3017 383 3051 399
rect 3165 683 3199 1025
rect 3296 1053 3364 1093
rect 3296 1019 3313 1053
rect 3347 1019 3364 1053
rect 3471 1365 3505 1405
rect 3471 1297 3505 1331
rect 3471 1229 3505 1263
rect 3471 1161 3505 1195
rect 3471 1093 3505 1127
rect 3559 1365 3593 1446
rect 3962 1423 4030 1446
rect 3559 1297 3593 1331
rect 3559 1229 3593 1263
rect 3559 1161 3593 1195
rect 3559 1111 3593 1127
rect 3647 1365 3857 1399
rect 3647 1297 3681 1331
rect 3647 1229 3681 1263
rect 3647 1161 3681 1195
rect 3647 1093 3681 1127
rect 3471 1025 3681 1059
rect 3735 1297 3769 1313
rect 3735 1229 3769 1263
rect 3735 1161 3769 1195
rect 3735 1093 3769 1127
rect 3823 1297 3857 1331
rect 3823 1229 3857 1263
rect 3823 1161 3857 1195
rect 3823 1111 3857 1127
rect 3962 1389 3979 1423
rect 4013 1389 4030 1423
rect 3962 1349 4030 1389
rect 3962 1315 3979 1349
rect 4013 1315 4030 1349
rect 3962 1275 4030 1315
rect 3962 1241 3979 1275
rect 4013 1241 4030 1275
rect 3962 1201 4030 1241
rect 3962 1167 3979 1201
rect 4013 1167 4030 1201
rect 3962 1127 4030 1167
rect 3962 1093 3979 1127
rect 4013 1093 4030 1127
rect 3735 1025 3865 1059
rect 3296 979 3364 1019
rect 3296 945 3313 979
rect 3347 945 3364 979
rect 3296 905 3364 945
rect 3504 958 3538 974
rect 3690 958 3724 974
rect 3538 924 3569 942
rect 3504 908 3569 924
rect 3296 871 3313 905
rect 3347 871 3364 905
rect 3296 822 3364 871
rect 2425 168 2459 184
rect 2523 334 2557 350
rect 2523 262 2557 300
rect 2523 194 2557 228
rect 2329 124 2363 160
rect 2523 124 2557 160
rect 2363 90 2425 124
rect 2459 90 2523 124
rect 2329 34 2363 90
rect 2426 34 2460 90
rect 2523 34 2557 90
rect 2630 313 2698 353
rect 2630 279 2647 313
rect 2681 279 2698 313
rect 2630 239 2698 279
rect 2630 205 2647 239
rect 2681 205 2698 239
rect 2630 165 2698 205
rect 2630 131 2647 165
rect 2681 131 2698 165
rect 2630 91 2698 131
rect 2630 57 2647 91
rect 2681 57 2698 91
rect 2630 34 2698 57
rect 2786 333 2820 349
rect 3165 348 3199 649
rect 3535 683 3569 908
rect 2786 261 2820 299
rect 2786 193 2820 227
rect 2883 314 3199 348
rect 3296 461 3364 544
rect 3296 427 3313 461
rect 3347 427 3364 461
rect 3296 387 3364 427
rect 3296 353 3313 387
rect 3347 353 3364 387
rect 3535 433 3569 649
rect 3535 383 3569 399
rect 3683 924 3690 942
rect 3683 908 3724 924
rect 3683 831 3717 908
rect 3683 433 3717 797
rect 3683 383 3717 399
rect 3831 757 3865 1025
rect 3962 1053 4030 1093
rect 3962 1019 3979 1053
rect 4013 1019 4030 1053
rect 3962 979 4030 1019
rect 3962 945 3979 979
rect 4013 945 4030 979
rect 3962 905 4030 945
rect 3962 871 3979 905
rect 4013 871 4030 905
rect 3962 822 4030 871
rect 2883 217 2917 314
rect 2883 167 2917 183
rect 2980 261 3014 278
rect 2980 193 3014 227
rect 2786 123 2820 159
rect 3077 217 3111 314
rect 3296 313 3364 353
rect 3296 279 3313 313
rect 3347 279 3364 313
rect 3077 167 3111 183
rect 3174 261 3208 278
rect 3174 193 3208 227
rect 2980 123 3014 159
rect 3174 123 3208 159
rect 2820 89 2883 123
rect 2917 89 2980 123
rect 3014 89 3077 123
rect 3111 89 3174 123
rect 2786 34 2820 89
rect 2883 34 2917 89
rect 2980 34 3014 89
rect 3077 34 3111 89
rect 3174 34 3208 89
rect 3296 239 3364 279
rect 3296 205 3313 239
rect 3347 205 3364 239
rect 3296 165 3364 205
rect 3296 131 3313 165
rect 3347 131 3364 165
rect 3296 91 3364 131
rect 3296 57 3313 91
rect 3347 57 3364 91
rect 3296 34 3364 57
rect 3452 333 3486 349
rect 3831 348 3865 723
rect 3452 261 3486 299
rect 3452 193 3486 227
rect 3549 314 3865 348
rect 3962 461 4030 544
rect 3962 427 3979 461
rect 4013 427 4030 461
rect 3962 387 4030 427
rect 3962 353 3979 387
rect 4013 353 4030 387
rect 3549 217 3583 314
rect 3549 167 3583 183
rect 3646 261 3680 278
rect 3646 193 3680 227
rect 3452 123 3486 159
rect 3743 217 3777 314
rect 3962 313 4030 353
rect 3962 279 3979 313
rect 4013 279 4030 313
rect 3743 167 3777 183
rect 3840 261 3874 278
rect 3840 193 3874 227
rect 3646 123 3680 159
rect 3840 123 3874 159
rect 3486 89 3549 123
rect 3583 89 3646 123
rect 3680 89 3743 123
rect 3777 89 3840 123
rect 3452 34 3486 89
rect 3549 34 3583 89
rect 3646 34 3680 89
rect 3743 34 3777 89
rect 3840 34 3874 89
rect 3962 239 4030 279
rect 3962 205 3979 239
rect 4013 205 4030 239
rect 3962 165 4030 205
rect 3962 131 3979 165
rect 4013 131 4030 165
rect 3962 91 4030 131
rect 3962 57 3979 91
rect 4013 57 4030 91
rect 3962 34 4030 57
rect -34 17 4030 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 4030 17
rect -34 -34 4030 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 131 797 165 831
rect 279 723 313 757
rect 649 723 683 757
rect 797 575 831 609
rect 945 649 979 683
rect 1241 649 1275 683
rect 1389 723 1423 757
rect 1759 575 1793 609
rect 1907 797 1941 831
rect 2055 649 2089 683
rect 2351 649 2385 683
rect 2499 797 2533 831
rect 2869 723 2903 757
rect 3017 723 3051 757
rect 3165 649 3199 683
rect 3535 649 3569 683
rect 3683 797 3717 831
rect 3831 723 3865 757
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
<< metal1 >>
rect -34 1497 4030 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 4030 1497
rect -34 1446 4030 1463
rect 125 831 171 837
rect 1901 831 1947 837
rect 2493 831 2539 837
rect 3677 831 3723 837
rect 119 797 131 831
rect 165 797 1907 831
rect 1941 797 1953 831
rect 2487 797 2499 831
rect 2533 797 3683 831
rect 3717 797 3729 831
rect 125 791 171 797
rect 1901 791 1947 797
rect 2493 791 2539 797
rect 3677 791 3723 797
rect 273 757 319 763
rect 643 757 689 763
rect 1383 757 1429 763
rect 2863 757 2909 763
rect 3011 757 3057 763
rect 3825 757 3871 763
rect 267 723 279 757
rect 313 723 649 757
rect 683 723 695 757
rect 1377 723 1389 757
rect 1423 723 2869 757
rect 2903 723 2915 757
rect 3005 723 3017 757
rect 3051 723 3831 757
rect 3865 723 3877 757
rect 273 717 319 723
rect 643 717 689 723
rect 1383 717 1429 723
rect 2863 717 2909 723
rect 3011 717 3057 723
rect 3825 717 3871 723
rect 939 683 985 689
rect 1235 683 1281 689
rect 2049 683 2095 689
rect 2345 683 2391 689
rect 3159 683 3205 689
rect 3529 683 3575 689
rect 933 649 945 683
rect 979 649 1241 683
rect 1275 649 1287 683
rect 2043 649 2055 683
rect 2089 649 2351 683
rect 2385 649 2397 683
rect 3153 649 3165 683
rect 3199 649 3535 683
rect 3569 649 3581 683
rect 939 643 985 649
rect 1235 643 1281 649
rect 2049 643 2095 649
rect 2345 643 2391 649
rect 3159 643 3205 649
rect 3529 643 3575 649
rect 791 609 837 615
rect 1753 609 1799 615
rect 785 575 797 609
rect 831 575 1759 609
rect 1793 575 1805 609
rect 791 569 837 575
rect 1753 569 1799 575
rect -34 17 4030 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 4030 17
rect -34 -34 4030 -17
<< labels >>
rlabel metal1 3165 649 3199 683 1 Q
port 1 n
rlabel metal1 3165 575 3199 609 1 Q
port 2 n
rlabel metal1 3165 501 3199 535 1 Q
port 3 n
rlabel metal1 3165 427 3199 461 1 Q
port 4 n
rlabel metal1 3165 871 3199 905 1 Q
port 5 n
rlabel metal1 3535 427 3569 461 1 Q
port 6 n
rlabel metal1 3535 501 3569 535 1 Q
port 7 n
rlabel metal1 3535 575 3569 609 1 Q
port 8 n
rlabel metal1 3535 649 3569 683 1 Q
port 9 n
rlabel metal1 3535 871 3569 905 1 Q
port 10 n
rlabel metal1 131 797 165 831 1 D
port 11 n
rlabel metal1 131 871 165 905 1 D
port 12 n
rlabel metal1 131 723 165 757 1 D
port 13 n
rlabel metal1 131 649 165 683 1 D
port 14 n
rlabel metal1 131 575 165 609 1 D
port 15 n
rlabel metal1 131 501 165 535 1 D
port 16 n
rlabel metal1 131 427 165 461 1 D
port 17 n
rlabel metal1 1907 427 1941 461 1 D
port 18 n
rlabel metal1 1907 501 1941 535 1 D
port 19 n
rlabel metal1 1907 575 1941 609 1 D
port 20 n
rlabel metal1 1907 649 1941 683 1 D
port 21 n
rlabel metal1 1907 797 1941 831 1 D
port 22 n
rlabel metal1 1907 871 1941 905 1 D
port 23 n
rlabel metal1 797 575 831 609 1 GATE
port 24 n
rlabel metal1 797 501 831 535 1 GATE
port 25 n
rlabel metal1 797 649 831 683 1 GATE
port 26 n
rlabel metal1 797 723 831 757 1 GATE
port 27 n
rlabel metal1 797 871 831 905 1 GATE
port 28 n
rlabel metal1 1759 501 1793 535 1 GATE
port 29 n
rlabel metal1 1759 575 1793 609 1 GATE
port 30 n
rlabel metal1 1759 649 1793 683 1 GATE
port 31 n
rlabel metal1 1759 871 1793 905 1 GATE
port 32 n
rlabel metal1 -34 1446 4030 1514 1 VPWR
port 33 n
rlabel metal1 -34 -34 4030 34 1 VGND
port 34 n
rlabel nwell 57 1463 91 1497 1 VPB
port 35 n
rlabel pwell 57 -17 91 17 1 VNB
port 36 n
<< end >>
