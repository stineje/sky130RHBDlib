* SPICE3 file created from AOI3X1.ext - technology: sky130A

.subckt AOI3X1 YN A B C VDD GND
X0 YN a_217_1004 GND GND nshort w=3 l=0.15
X1 VDD B a_217_1004 VDD pshort w=2 l=0.15 M=2
X2 GND A a_112_73 GND nshort w=3 l=0.15
X3 a_797_1005 C YN VDD pshort w=2 l=0.15 M=2
X4 a_217_1004 A VDD VDD pshort w=2 l=0.15 M=2
X5 a_217_1004 B a_112_73 GND nshort w=3 l=0.15
X6 YN C GND GND nshort w=3 l=0.15
X7 a_797_1005 a_217_1004 VDD VDD pshort w=2 l=0.15 M=2
C0 VDD GND 3.54fF
.ends
