magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect 419 4416 9008 4522
rect 9038 3851 9109 4552
<< pwell >>
rect 417 3446 8713 3532
<< psubdiff >>
rect 443 3472 519 3506
rect 553 3472 587 3506
rect 621 3472 655 3506
rect 689 3472 723 3506
rect 757 3472 791 3506
rect 825 3472 859 3506
rect 893 3472 927 3506
rect 961 3472 995 3506
rect 1029 3472 1063 3506
rect 1097 3472 1131 3506
rect 1165 3472 1199 3506
rect 1233 3472 1267 3506
rect 1301 3472 1335 3506
rect 1369 3472 1403 3506
rect 1437 3472 1471 3506
rect 1505 3472 1539 3506
rect 1573 3472 1607 3506
rect 1641 3472 1675 3506
rect 1709 3472 1743 3506
rect 1777 3472 1811 3506
rect 1845 3472 1879 3506
rect 1913 3472 1947 3506
rect 1981 3472 2015 3506
rect 2049 3472 2083 3506
rect 2117 3472 2151 3506
rect 2185 3472 2219 3506
rect 2253 3472 2287 3506
rect 2321 3472 2355 3506
rect 2389 3472 2423 3506
rect 2457 3472 2491 3506
<< nsubdiff >>
rect 429 4452 479 4486
rect 513 4452 547 4486
rect 581 4452 615 4486
rect 649 4452 683 4486
rect 717 4452 751 4486
rect 785 4452 819 4486
rect 853 4452 887 4486
rect 921 4452 955 4486
rect 989 4452 1023 4486
rect 1057 4452 1091 4486
rect 1125 4452 1159 4486
rect 1193 4452 1227 4486
rect 1261 4452 1295 4486
rect 1329 4452 1363 4486
rect 1397 4452 1431 4486
rect 1465 4452 1499 4486
rect 1533 4452 1567 4486
rect 1601 4452 1635 4486
rect 1669 4452 1703 4486
rect 1737 4452 1771 4486
rect 1805 4452 1839 4486
rect 1873 4452 1907 4486
rect 1941 4452 1975 4486
rect 2009 4452 2043 4486
rect 2077 4452 2111 4486
rect 2145 4452 2179 4486
rect 2213 4452 2247 4486
rect 2281 4452 2315 4486
rect 2349 4452 2383 4486
rect 2417 4452 2451 4486
rect 2485 4452 2505 4486
<< mvpsubdiff >>
rect 2525 3472 2559 3506
rect 2593 3472 2627 3506
rect 2661 3472 2695 3506
rect 2729 3472 2763 3506
rect 2797 3472 2831 3506
rect 2865 3472 2899 3506
rect 2933 3472 2967 3506
rect 3001 3472 3035 3506
rect 3069 3472 3103 3506
rect 3137 3472 3171 3506
rect 3205 3472 3239 3506
rect 3273 3472 3307 3506
rect 3341 3472 3375 3506
rect 3409 3472 3443 3506
rect 3477 3472 3511 3506
rect 3545 3472 3579 3506
rect 3613 3472 3647 3506
rect 3681 3472 3715 3506
rect 3749 3472 3783 3506
rect 3817 3472 3851 3506
rect 3885 3472 3919 3506
rect 3953 3472 3987 3506
rect 4021 3472 4055 3506
rect 4089 3472 4123 3506
rect 4157 3472 4191 3506
rect 4225 3472 4259 3506
rect 4293 3472 4327 3506
rect 4361 3472 4395 3506
rect 4429 3472 4463 3506
rect 4497 3472 4531 3506
rect 4565 3472 4599 3506
rect 4633 3472 4667 3506
rect 4701 3472 4735 3506
rect 4769 3472 4803 3506
rect 4837 3472 4871 3506
rect 4905 3472 4939 3506
rect 4973 3472 5007 3506
rect 5041 3472 5075 3506
rect 5109 3472 5143 3506
rect 5177 3472 5211 3506
rect 5245 3472 5279 3506
rect 5313 3472 5347 3506
rect 5381 3472 5415 3506
rect 5449 3472 5483 3506
rect 5517 3472 5551 3506
rect 5585 3472 5619 3506
rect 5653 3472 5687 3506
rect 5721 3472 5755 3506
rect 5789 3472 5823 3506
rect 5857 3472 5891 3506
rect 5925 3472 5959 3506
rect 5993 3472 6027 3506
rect 6061 3472 6095 3506
rect 6129 3472 6163 3506
rect 6197 3472 6231 3506
rect 6265 3472 6299 3506
rect 6333 3472 6367 3506
rect 6401 3472 6435 3506
rect 6469 3472 6503 3506
rect 6537 3472 6571 3506
rect 6605 3472 6639 3506
rect 6673 3472 6707 3506
rect 6741 3472 6775 3506
rect 6809 3472 6843 3506
rect 6877 3472 6911 3506
rect 6945 3472 6979 3506
rect 7013 3472 7047 3506
rect 7081 3472 7115 3506
rect 7149 3472 7183 3506
rect 7217 3472 7251 3506
rect 7285 3472 7319 3506
rect 7353 3472 7387 3506
rect 7421 3472 7455 3506
rect 7489 3472 7523 3506
rect 7557 3472 7591 3506
rect 7625 3472 7659 3506
rect 7693 3472 7727 3506
rect 7761 3472 7795 3506
rect 7829 3472 7863 3506
rect 7897 3472 7931 3506
rect 7965 3472 7999 3506
rect 8033 3472 8067 3506
rect 8101 3472 8135 3506
rect 8169 3472 8203 3506
rect 8237 3472 8271 3506
rect 8305 3472 8339 3506
rect 8373 3472 8407 3506
rect 8441 3472 8475 3506
rect 8509 3472 8543 3506
rect 8577 3472 8611 3506
rect 8645 3472 8687 3506
<< mvnsubdiff >>
rect 2505 4452 2519 4486
rect 2553 4452 2587 4486
rect 2621 4452 2655 4486
rect 2689 4452 2723 4486
rect 2757 4452 2791 4486
rect 2825 4452 2859 4486
rect 2893 4452 2927 4486
rect 2961 4452 2995 4486
rect 3029 4452 3063 4486
rect 3097 4452 3131 4486
rect 3165 4452 3199 4486
rect 3233 4452 3267 4486
rect 3301 4452 3335 4486
rect 3369 4452 3403 4486
rect 3437 4452 3471 4486
rect 3505 4452 3539 4486
rect 3573 4452 3607 4486
rect 3641 4452 3675 4486
rect 3709 4452 3743 4486
rect 3777 4452 3811 4486
rect 3845 4452 3879 4486
rect 3913 4452 3947 4486
rect 3981 4452 4015 4486
rect 4049 4452 4083 4486
rect 4117 4452 4151 4486
rect 4185 4452 4219 4486
rect 4253 4452 4287 4486
rect 4321 4452 4355 4486
rect 4389 4452 4423 4486
rect 4457 4452 4491 4486
rect 4525 4452 4559 4486
rect 4593 4452 4627 4486
rect 4661 4452 4695 4486
rect 4729 4452 4763 4486
rect 4797 4452 4831 4486
rect 4865 4452 4899 4486
rect 4933 4452 4967 4486
rect 5001 4452 5035 4486
rect 5069 4452 5103 4486
rect 5137 4452 5171 4486
rect 5205 4452 5239 4486
rect 5273 4452 5307 4486
rect 5341 4452 5375 4486
rect 5409 4452 5443 4486
rect 5477 4452 5511 4486
rect 5545 4452 5579 4486
rect 5613 4452 5647 4486
rect 5681 4452 5715 4486
rect 5749 4452 5783 4486
rect 5817 4452 5851 4486
rect 5885 4452 5919 4486
rect 5953 4452 5987 4486
rect 6021 4452 6055 4486
rect 6089 4452 6123 4486
rect 6157 4452 6191 4486
rect 6225 4452 6259 4486
rect 6293 4452 6327 4486
rect 6361 4452 6395 4486
rect 6429 4452 6463 4486
rect 6497 4452 6531 4486
rect 6565 4452 6599 4486
rect 6633 4452 6667 4486
rect 6701 4452 6735 4486
rect 6769 4452 6803 4486
rect 6837 4452 6871 4486
rect 6905 4452 6939 4486
rect 6973 4452 7007 4486
rect 7041 4452 7075 4486
rect 7109 4452 7143 4486
rect 7177 4452 7211 4486
rect 7245 4452 7279 4486
rect 7313 4452 7347 4486
rect 7381 4452 7415 4486
rect 7449 4452 7483 4486
rect 7517 4452 7551 4486
rect 7585 4452 7619 4486
rect 7653 4452 7687 4486
rect 7721 4452 7755 4486
rect 7789 4452 7823 4486
rect 7857 4452 7891 4486
rect 7925 4452 7959 4486
rect 7993 4452 8027 4486
rect 8061 4452 8095 4486
rect 8129 4452 8163 4486
rect 8197 4452 8231 4486
rect 8265 4452 8299 4486
rect 8333 4452 8367 4486
rect 8401 4452 8435 4486
rect 8469 4452 8503 4486
rect 8537 4452 8571 4486
rect 8605 4452 8639 4486
rect 8673 4452 8707 4486
rect 8741 4452 8775 4486
rect 8809 4452 8843 4486
rect 8877 4452 8911 4486
rect 8945 4452 8972 4486
<< psubdiffcont >>
rect 519 3472 553 3506
rect 587 3472 621 3506
rect 655 3472 689 3506
rect 723 3472 757 3506
rect 791 3472 825 3506
rect 859 3472 893 3506
rect 927 3472 961 3506
rect 995 3472 1029 3506
rect 1063 3472 1097 3506
rect 1131 3472 1165 3506
rect 1199 3472 1233 3506
rect 1267 3472 1301 3506
rect 1335 3472 1369 3506
rect 1403 3472 1437 3506
rect 1471 3472 1505 3506
rect 1539 3472 1573 3506
rect 1607 3472 1641 3506
rect 1675 3472 1709 3506
rect 1743 3472 1777 3506
rect 1811 3472 1845 3506
rect 1879 3472 1913 3506
rect 1947 3472 1981 3506
rect 2015 3472 2049 3506
rect 2083 3472 2117 3506
rect 2151 3472 2185 3506
rect 2219 3472 2253 3506
rect 2287 3472 2321 3506
rect 2355 3472 2389 3506
rect 2423 3472 2457 3506
rect 2491 3472 2505 3506
<< nsubdiffcont >>
rect 479 4452 513 4486
rect 547 4452 581 4486
rect 615 4452 649 4486
rect 683 4452 717 4486
rect 751 4452 785 4486
rect 819 4452 853 4486
rect 887 4452 921 4486
rect 955 4452 989 4486
rect 1023 4452 1057 4486
rect 1091 4452 1125 4486
rect 1159 4452 1193 4486
rect 1227 4452 1261 4486
rect 1295 4452 1329 4486
rect 1363 4452 1397 4486
rect 1431 4452 1465 4486
rect 1499 4452 1533 4486
rect 1567 4452 1601 4486
rect 1635 4452 1669 4486
rect 1703 4452 1737 4486
rect 1771 4452 1805 4486
rect 1839 4452 1873 4486
rect 1907 4452 1941 4486
rect 1975 4452 2009 4486
rect 2043 4452 2077 4486
rect 2111 4452 2145 4486
rect 2179 4452 2213 4486
rect 2247 4452 2281 4486
rect 2315 4452 2349 4486
rect 2383 4452 2417 4486
rect 2451 4452 2485 4486
<< mvpsubdiffcont >>
rect 2505 3472 2525 3506
rect 2559 3472 2593 3506
rect 2627 3472 2661 3506
rect 2695 3472 2729 3506
rect 2763 3472 2797 3506
rect 2831 3472 2865 3506
rect 2899 3472 2933 3506
rect 2967 3472 3001 3506
rect 3035 3472 3069 3506
rect 3103 3472 3137 3506
rect 3171 3472 3205 3506
rect 3239 3472 3273 3506
rect 3307 3472 3341 3506
rect 3375 3472 3409 3506
rect 3443 3472 3477 3506
rect 3511 3472 3545 3506
rect 3579 3472 3613 3506
rect 3647 3472 3681 3506
rect 3715 3472 3749 3506
rect 3783 3472 3817 3506
rect 3851 3472 3885 3506
rect 3919 3472 3953 3506
rect 3987 3472 4021 3506
rect 4055 3472 4089 3506
rect 4123 3472 4157 3506
rect 4191 3472 4225 3506
rect 4259 3472 4293 3506
rect 4327 3472 4361 3506
rect 4395 3472 4429 3506
rect 4463 3472 4497 3506
rect 4531 3472 4565 3506
rect 4599 3472 4633 3506
rect 4667 3472 4701 3506
rect 4735 3472 4769 3506
rect 4803 3472 4837 3506
rect 4871 3472 4905 3506
rect 4939 3472 4973 3506
rect 5007 3472 5041 3506
rect 5075 3472 5109 3506
rect 5143 3472 5177 3506
rect 5211 3472 5245 3506
rect 5279 3472 5313 3506
rect 5347 3472 5381 3506
rect 5415 3472 5449 3506
rect 5483 3472 5517 3506
rect 5551 3472 5585 3506
rect 5619 3472 5653 3506
rect 5687 3472 5721 3506
rect 5755 3472 5789 3506
rect 5823 3472 5857 3506
rect 5891 3472 5925 3506
rect 5959 3472 5993 3506
rect 6027 3472 6061 3506
rect 6095 3472 6129 3506
rect 6163 3472 6197 3506
rect 6231 3472 6265 3506
rect 6299 3472 6333 3506
rect 6367 3472 6401 3506
rect 6435 3472 6469 3506
rect 6503 3472 6537 3506
rect 6571 3472 6605 3506
rect 6639 3472 6673 3506
rect 6707 3472 6741 3506
rect 6775 3472 6809 3506
rect 6843 3472 6877 3506
rect 6911 3472 6945 3506
rect 6979 3472 7013 3506
rect 7047 3472 7081 3506
rect 7115 3472 7149 3506
rect 7183 3472 7217 3506
rect 7251 3472 7285 3506
rect 7319 3472 7353 3506
rect 7387 3472 7421 3506
rect 7455 3472 7489 3506
rect 7523 3472 7557 3506
rect 7591 3472 7625 3506
rect 7659 3472 7693 3506
rect 7727 3472 7761 3506
rect 7795 3472 7829 3506
rect 7863 3472 7897 3506
rect 7931 3472 7965 3506
rect 7999 3472 8033 3506
rect 8067 3472 8101 3506
rect 8135 3472 8169 3506
rect 8203 3472 8237 3506
rect 8271 3472 8305 3506
rect 8339 3472 8373 3506
rect 8407 3472 8441 3506
rect 8475 3472 8509 3506
rect 8543 3472 8577 3506
rect 8611 3472 8645 3506
<< mvnsubdiffcont >>
rect 2519 4452 2553 4486
rect 2587 4452 2621 4486
rect 2655 4452 2689 4486
rect 2723 4452 2757 4486
rect 2791 4452 2825 4486
rect 2859 4452 2893 4486
rect 2927 4452 2961 4486
rect 2995 4452 3029 4486
rect 3063 4452 3097 4486
rect 3131 4452 3165 4486
rect 3199 4452 3233 4486
rect 3267 4452 3301 4486
rect 3335 4452 3369 4486
rect 3403 4452 3437 4486
rect 3471 4452 3505 4486
rect 3539 4452 3573 4486
rect 3607 4452 3641 4486
rect 3675 4452 3709 4486
rect 3743 4452 3777 4486
rect 3811 4452 3845 4486
rect 3879 4452 3913 4486
rect 3947 4452 3981 4486
rect 4015 4452 4049 4486
rect 4083 4452 4117 4486
rect 4151 4452 4185 4486
rect 4219 4452 4253 4486
rect 4287 4452 4321 4486
rect 4355 4452 4389 4486
rect 4423 4452 4457 4486
rect 4491 4452 4525 4486
rect 4559 4452 4593 4486
rect 4627 4452 4661 4486
rect 4695 4452 4729 4486
rect 4763 4452 4797 4486
rect 4831 4452 4865 4486
rect 4899 4452 4933 4486
rect 4967 4452 5001 4486
rect 5035 4452 5069 4486
rect 5103 4452 5137 4486
rect 5171 4452 5205 4486
rect 5239 4452 5273 4486
rect 5307 4452 5341 4486
rect 5375 4452 5409 4486
rect 5443 4452 5477 4486
rect 5511 4452 5545 4486
rect 5579 4452 5613 4486
rect 5647 4452 5681 4486
rect 5715 4452 5749 4486
rect 5783 4452 5817 4486
rect 5851 4452 5885 4486
rect 5919 4452 5953 4486
rect 5987 4452 6021 4486
rect 6055 4452 6089 4486
rect 6123 4452 6157 4486
rect 6191 4452 6225 4486
rect 6259 4452 6293 4486
rect 6327 4452 6361 4486
rect 6395 4452 6429 4486
rect 6463 4452 6497 4486
rect 6531 4452 6565 4486
rect 6599 4452 6633 4486
rect 6667 4452 6701 4486
rect 6735 4452 6769 4486
rect 6803 4452 6837 4486
rect 6871 4452 6905 4486
rect 6939 4452 6973 4486
rect 7007 4452 7041 4486
rect 7075 4452 7109 4486
rect 7143 4452 7177 4486
rect 7211 4452 7245 4486
rect 7279 4452 7313 4486
rect 7347 4452 7381 4486
rect 7415 4452 7449 4486
rect 7483 4452 7517 4486
rect 7551 4452 7585 4486
rect 7619 4452 7653 4486
rect 7687 4452 7721 4486
rect 7755 4452 7789 4486
rect 7823 4452 7857 4486
rect 7891 4452 7925 4486
rect 7959 4452 7993 4486
rect 8027 4452 8061 4486
rect 8095 4452 8129 4486
rect 8163 4452 8197 4486
rect 8231 4452 8265 4486
rect 8299 4452 8333 4486
rect 8367 4452 8401 4486
rect 8435 4452 8469 4486
rect 8503 4452 8537 4486
rect 8571 4452 8605 4486
rect 8639 4452 8673 4486
rect 8707 4452 8741 4486
rect 8775 4452 8809 4486
rect 8843 4452 8877 4486
rect 8911 4452 8945 4486
<< locali >>
rect 429 4452 467 4486
rect 513 4452 539 4486
rect 581 4452 611 4486
rect 649 4452 683 4486
rect 717 4452 751 4486
rect 789 4452 819 4486
rect 861 4452 887 4486
rect 933 4452 955 4486
rect 1005 4452 1023 4486
rect 1077 4452 1091 4486
rect 1149 4452 1159 4486
rect 1221 4452 1227 4486
rect 1293 4452 1295 4486
rect 1329 4452 1331 4486
rect 1397 4452 1403 4486
rect 1465 4452 1475 4486
rect 1533 4452 1547 4486
rect 1601 4452 1619 4486
rect 1669 4452 1691 4486
rect 1737 4452 1763 4486
rect 1805 4452 1835 4486
rect 1873 4452 1907 4486
rect 1941 4452 1975 4486
rect 2013 4452 2043 4486
rect 2085 4452 2111 4486
rect 2157 4452 2179 4486
rect 2229 4452 2247 4486
rect 2301 4452 2315 4486
rect 2373 4452 2383 4486
rect 2445 4452 2451 4486
rect 2517 4452 2519 4486
rect 2553 4452 2555 4486
rect 2621 4452 2627 4486
rect 2689 4452 2699 4486
rect 2757 4452 2771 4486
rect 2825 4452 2843 4486
rect 2893 4452 2915 4486
rect 2961 4452 2987 4486
rect 3029 4452 3059 4486
rect 3097 4452 3131 4486
rect 3165 4452 3199 4486
rect 3237 4452 3267 4486
rect 3309 4452 3335 4486
rect 3381 4452 3403 4486
rect 3453 4452 3471 4486
rect 3525 4452 3539 4486
rect 3597 4452 3607 4486
rect 3669 4452 3675 4486
rect 3741 4452 3743 4486
rect 3777 4452 3779 4486
rect 3845 4452 3851 4486
rect 3913 4452 3923 4486
rect 3981 4452 3995 4486
rect 4049 4452 4067 4486
rect 4117 4452 4139 4486
rect 4185 4452 4211 4486
rect 4253 4452 4283 4486
rect 4321 4452 4355 4486
rect 4389 4452 4423 4486
rect 4461 4452 4491 4486
rect 4533 4452 4559 4486
rect 4605 4452 4627 4486
rect 4677 4452 4695 4486
rect 4749 4452 4763 4486
rect 4821 4452 4831 4486
rect 4893 4452 4899 4486
rect 4965 4452 4967 4486
rect 5001 4452 5003 4486
rect 5069 4452 5075 4486
rect 5137 4452 5147 4486
rect 5205 4452 5219 4486
rect 5273 4452 5291 4486
rect 5341 4452 5363 4486
rect 5409 4452 5435 4486
rect 5477 4452 5507 4486
rect 5545 4452 5579 4486
rect 5613 4452 5647 4486
rect 5685 4452 5715 4486
rect 5757 4452 5783 4486
rect 5829 4452 5851 4486
rect 5901 4452 5919 4486
rect 5973 4452 5987 4486
rect 6045 4452 6055 4486
rect 6117 4452 6123 4486
rect 6189 4452 6191 4486
rect 6225 4452 6227 4486
rect 6293 4452 6299 4486
rect 6361 4452 6371 4486
rect 6429 4452 6443 4486
rect 6497 4452 6515 4486
rect 6565 4452 6587 4486
rect 6633 4452 6659 4486
rect 6701 4452 6731 4486
rect 6769 4452 6803 4486
rect 6837 4452 6871 4486
rect 6909 4452 6939 4486
rect 6981 4452 7007 4486
rect 7053 4452 7075 4486
rect 7125 4452 7143 4486
rect 7197 4452 7211 4486
rect 7269 4452 7279 4486
rect 7341 4452 7347 4486
rect 7413 4452 7415 4486
rect 7449 4452 7451 4486
rect 7517 4452 7523 4486
rect 7585 4452 7595 4486
rect 7653 4452 7667 4486
rect 7721 4452 7739 4486
rect 7789 4452 7811 4486
rect 7857 4452 7883 4486
rect 7925 4452 7955 4486
rect 7993 4452 8027 4486
rect 8061 4452 8095 4486
rect 8133 4452 8163 4486
rect 8205 4452 8231 4486
rect 8277 4452 8299 4486
rect 8349 4452 8367 4486
rect 8421 4452 8435 4486
rect 8493 4452 8503 4486
rect 8565 4452 8571 4486
rect 8637 4452 8639 4486
rect 8673 4452 8675 4486
rect 8741 4452 8747 4486
rect 8809 4452 8819 4486
rect 8877 4452 8891 4486
rect 8945 4452 8972 4486
rect 8998 4230 9064 4242
rect 2625 4126 2659 4164
rect 8998 4196 9014 4230
rect 9048 4196 9064 4230
rect 3417 4121 3455 4155
rect 7293 4074 7359 4156
rect 7293 4040 7308 4074
rect 7342 4040 7359 4074
rect 7293 4002 7359 4040
rect 8650 4149 8716 4161
rect 8650 4115 8666 4149
rect 8700 4115 8716 4149
rect 8650 4077 8716 4115
rect 8650 4043 8666 4077
rect 8700 4043 8716 4077
rect 7293 3968 7308 4002
rect 7342 3968 7359 4002
rect 2696 3862 2889 3885
rect 2923 3862 2943 3885
rect 2696 3824 2943 3862
rect 2696 3790 2889 3824
rect 2923 3790 2943 3824
rect 2696 3768 2943 3790
rect 3061 3805 3095 3843
rect 3154 3768 3351 3870
rect 3488 3869 3653 3870
rect 3500 3835 3538 3869
rect 3572 3835 3653 3869
rect 3488 3768 3653 3835
rect 7222 3859 7256 3897
rect 7293 3870 7359 3968
rect 8474 3992 8540 4019
rect 8474 3958 8486 3992
rect 8520 3958 8540 3992
rect 8474 3920 8540 3958
rect 8226 3864 8260 3920
rect 8474 3886 8486 3920
rect 8520 3886 8540 3920
rect 8226 3792 8260 3830
rect 2588 3709 2626 3743
rect 3154 3726 3232 3768
rect 8474 3870 8540 3886
rect 8650 3870 8716 4043
rect 8998 4158 9064 4196
rect 8998 4124 9014 4158
rect 9048 4124 9064 4158
rect 8312 3800 8346 3838
rect 8998 3870 9064 4124
rect 8754 3800 8788 3838
rect 8893 3768 9064 3870
rect 2978 3589 3232 3726
rect 443 3472 507 3506
rect 553 3472 579 3506
rect 621 3472 651 3506
rect 689 3472 723 3506
rect 757 3472 791 3506
rect 829 3472 859 3506
rect 901 3472 927 3506
rect 973 3472 995 3506
rect 1045 3472 1063 3506
rect 1117 3472 1131 3506
rect 1189 3472 1199 3506
rect 1261 3472 1267 3506
rect 1333 3472 1335 3506
rect 1369 3472 1371 3506
rect 1437 3472 1443 3506
rect 1505 3472 1515 3506
rect 1573 3472 1587 3506
rect 1641 3472 1659 3506
rect 1709 3472 1731 3506
rect 1777 3472 1803 3506
rect 1845 3472 1875 3506
rect 1913 3472 1947 3506
rect 1981 3472 2015 3506
rect 2053 3472 2083 3506
rect 2125 3472 2151 3506
rect 2197 3472 2219 3506
rect 2269 3472 2287 3506
rect 2341 3472 2355 3506
rect 2413 3472 2423 3506
rect 2485 3472 2491 3506
rect 2557 3472 2559 3506
rect 2593 3472 2595 3506
rect 2661 3472 2667 3506
rect 2729 3472 2739 3506
rect 2797 3472 2811 3506
rect 2865 3472 2883 3506
rect 2933 3472 2955 3506
rect 3001 3472 3027 3506
rect 3069 3472 3099 3506
rect 3137 3472 3171 3506
rect 3205 3472 3239 3506
rect 3277 3472 3307 3506
rect 3349 3472 3375 3506
rect 3421 3472 3443 3506
rect 3493 3472 3511 3506
rect 3565 3472 3579 3506
rect 3637 3472 3647 3506
rect 3709 3472 3715 3506
rect 3781 3472 3783 3506
rect 3817 3472 3819 3506
rect 3885 3472 3891 3506
rect 3953 3472 3963 3506
rect 4021 3472 4035 3506
rect 4089 3472 4107 3506
rect 4157 3472 4179 3506
rect 4225 3472 4251 3506
rect 4293 3472 4323 3506
rect 4361 3472 4395 3506
rect 4429 3472 4463 3506
rect 4501 3472 4531 3506
rect 4573 3472 4599 3506
rect 4645 3472 4667 3506
rect 4717 3472 4735 3506
rect 4789 3472 4803 3506
rect 4861 3472 4871 3506
rect 4933 3472 4939 3506
rect 5005 3472 5007 3506
rect 5041 3472 5043 3506
rect 5109 3472 5115 3506
rect 5177 3472 5187 3506
rect 5245 3472 5259 3506
rect 5313 3472 5331 3506
rect 5381 3472 5403 3506
rect 5449 3472 5475 3506
rect 5517 3472 5547 3506
rect 5585 3472 5619 3506
rect 5653 3472 5687 3506
rect 5725 3472 5755 3506
rect 5797 3472 5823 3506
rect 5869 3472 5891 3506
rect 5941 3472 5959 3506
rect 6013 3472 6027 3506
rect 6085 3472 6095 3506
rect 6157 3472 6163 3506
rect 6229 3472 6231 3506
rect 6265 3472 6267 3506
rect 6333 3472 6339 3506
rect 6401 3472 6411 3506
rect 6469 3472 6483 3506
rect 6537 3472 6555 3506
rect 6605 3472 6627 3506
rect 6673 3472 6699 3506
rect 6741 3472 6771 3506
rect 6809 3472 6843 3506
rect 6877 3472 6911 3506
rect 6949 3472 6979 3506
rect 7021 3472 7047 3506
rect 7093 3472 7115 3506
rect 7165 3472 7183 3506
rect 7237 3472 7251 3506
rect 7309 3472 7319 3506
rect 7381 3472 7387 3506
rect 7453 3472 7455 3506
rect 7489 3472 7491 3506
rect 7557 3472 7563 3506
rect 7625 3472 7635 3506
rect 7693 3472 7707 3506
rect 7761 3472 7779 3506
rect 7829 3472 7851 3506
rect 7897 3472 7923 3506
rect 7965 3472 7995 3506
rect 8033 3472 8067 3506
rect 8101 3472 8135 3506
rect 8173 3472 8203 3506
rect 8245 3472 8271 3506
rect 8317 3472 8339 3506
rect 8389 3472 8407 3506
rect 8461 3472 8475 3506
rect 8533 3472 8543 3506
rect 8605 3472 8611 3506
rect 8645 3472 8687 3506
<< viali >>
rect 467 4452 479 4486
rect 479 4452 501 4486
rect 539 4452 547 4486
rect 547 4452 573 4486
rect 611 4452 615 4486
rect 615 4452 645 4486
rect 683 4452 717 4486
rect 755 4452 785 4486
rect 785 4452 789 4486
rect 827 4452 853 4486
rect 853 4452 861 4486
rect 899 4452 921 4486
rect 921 4452 933 4486
rect 971 4452 989 4486
rect 989 4452 1005 4486
rect 1043 4452 1057 4486
rect 1057 4452 1077 4486
rect 1115 4452 1125 4486
rect 1125 4452 1149 4486
rect 1187 4452 1193 4486
rect 1193 4452 1221 4486
rect 1259 4452 1261 4486
rect 1261 4452 1293 4486
rect 1331 4452 1363 4486
rect 1363 4452 1365 4486
rect 1403 4452 1431 4486
rect 1431 4452 1437 4486
rect 1475 4452 1499 4486
rect 1499 4452 1509 4486
rect 1547 4452 1567 4486
rect 1567 4452 1581 4486
rect 1619 4452 1635 4486
rect 1635 4452 1653 4486
rect 1691 4452 1703 4486
rect 1703 4452 1725 4486
rect 1763 4452 1771 4486
rect 1771 4452 1797 4486
rect 1835 4452 1839 4486
rect 1839 4452 1869 4486
rect 1907 4452 1941 4486
rect 1979 4452 2009 4486
rect 2009 4452 2013 4486
rect 2051 4452 2077 4486
rect 2077 4452 2085 4486
rect 2123 4452 2145 4486
rect 2145 4452 2157 4486
rect 2195 4452 2213 4486
rect 2213 4452 2229 4486
rect 2267 4452 2281 4486
rect 2281 4452 2301 4486
rect 2339 4452 2349 4486
rect 2349 4452 2373 4486
rect 2411 4452 2417 4486
rect 2417 4452 2445 4486
rect 2483 4452 2485 4486
rect 2485 4452 2517 4486
rect 2555 4452 2587 4486
rect 2587 4452 2589 4486
rect 2627 4452 2655 4486
rect 2655 4452 2661 4486
rect 2699 4452 2723 4486
rect 2723 4452 2733 4486
rect 2771 4452 2791 4486
rect 2791 4452 2805 4486
rect 2843 4452 2859 4486
rect 2859 4452 2877 4486
rect 2915 4452 2927 4486
rect 2927 4452 2949 4486
rect 2987 4452 2995 4486
rect 2995 4452 3021 4486
rect 3059 4452 3063 4486
rect 3063 4452 3093 4486
rect 3131 4452 3165 4486
rect 3203 4452 3233 4486
rect 3233 4452 3237 4486
rect 3275 4452 3301 4486
rect 3301 4452 3309 4486
rect 3347 4452 3369 4486
rect 3369 4452 3381 4486
rect 3419 4452 3437 4486
rect 3437 4452 3453 4486
rect 3491 4452 3505 4486
rect 3505 4452 3525 4486
rect 3563 4452 3573 4486
rect 3573 4452 3597 4486
rect 3635 4452 3641 4486
rect 3641 4452 3669 4486
rect 3707 4452 3709 4486
rect 3709 4452 3741 4486
rect 3779 4452 3811 4486
rect 3811 4452 3813 4486
rect 3851 4452 3879 4486
rect 3879 4452 3885 4486
rect 3923 4452 3947 4486
rect 3947 4452 3957 4486
rect 3995 4452 4015 4486
rect 4015 4452 4029 4486
rect 4067 4452 4083 4486
rect 4083 4452 4101 4486
rect 4139 4452 4151 4486
rect 4151 4452 4173 4486
rect 4211 4452 4219 4486
rect 4219 4452 4245 4486
rect 4283 4452 4287 4486
rect 4287 4452 4317 4486
rect 4355 4452 4389 4486
rect 4427 4452 4457 4486
rect 4457 4452 4461 4486
rect 4499 4452 4525 4486
rect 4525 4452 4533 4486
rect 4571 4452 4593 4486
rect 4593 4452 4605 4486
rect 4643 4452 4661 4486
rect 4661 4452 4677 4486
rect 4715 4452 4729 4486
rect 4729 4452 4749 4486
rect 4787 4452 4797 4486
rect 4797 4452 4821 4486
rect 4859 4452 4865 4486
rect 4865 4452 4893 4486
rect 4931 4452 4933 4486
rect 4933 4452 4965 4486
rect 5003 4452 5035 4486
rect 5035 4452 5037 4486
rect 5075 4452 5103 4486
rect 5103 4452 5109 4486
rect 5147 4452 5171 4486
rect 5171 4452 5181 4486
rect 5219 4452 5239 4486
rect 5239 4452 5253 4486
rect 5291 4452 5307 4486
rect 5307 4452 5325 4486
rect 5363 4452 5375 4486
rect 5375 4452 5397 4486
rect 5435 4452 5443 4486
rect 5443 4452 5469 4486
rect 5507 4452 5511 4486
rect 5511 4452 5541 4486
rect 5579 4452 5613 4486
rect 5651 4452 5681 4486
rect 5681 4452 5685 4486
rect 5723 4452 5749 4486
rect 5749 4452 5757 4486
rect 5795 4452 5817 4486
rect 5817 4452 5829 4486
rect 5867 4452 5885 4486
rect 5885 4452 5901 4486
rect 5939 4452 5953 4486
rect 5953 4452 5973 4486
rect 6011 4452 6021 4486
rect 6021 4452 6045 4486
rect 6083 4452 6089 4486
rect 6089 4452 6117 4486
rect 6155 4452 6157 4486
rect 6157 4452 6189 4486
rect 6227 4452 6259 4486
rect 6259 4452 6261 4486
rect 6299 4452 6327 4486
rect 6327 4452 6333 4486
rect 6371 4452 6395 4486
rect 6395 4452 6405 4486
rect 6443 4452 6463 4486
rect 6463 4452 6477 4486
rect 6515 4452 6531 4486
rect 6531 4452 6549 4486
rect 6587 4452 6599 4486
rect 6599 4452 6621 4486
rect 6659 4452 6667 4486
rect 6667 4452 6693 4486
rect 6731 4452 6735 4486
rect 6735 4452 6765 4486
rect 6803 4452 6837 4486
rect 6875 4452 6905 4486
rect 6905 4452 6909 4486
rect 6947 4452 6973 4486
rect 6973 4452 6981 4486
rect 7019 4452 7041 4486
rect 7041 4452 7053 4486
rect 7091 4452 7109 4486
rect 7109 4452 7125 4486
rect 7163 4452 7177 4486
rect 7177 4452 7197 4486
rect 7235 4452 7245 4486
rect 7245 4452 7269 4486
rect 7307 4452 7313 4486
rect 7313 4452 7341 4486
rect 7379 4452 7381 4486
rect 7381 4452 7413 4486
rect 7451 4452 7483 4486
rect 7483 4452 7485 4486
rect 7523 4452 7551 4486
rect 7551 4452 7557 4486
rect 7595 4452 7619 4486
rect 7619 4452 7629 4486
rect 7667 4452 7687 4486
rect 7687 4452 7701 4486
rect 7739 4452 7755 4486
rect 7755 4452 7773 4486
rect 7811 4452 7823 4486
rect 7823 4452 7845 4486
rect 7883 4452 7891 4486
rect 7891 4452 7917 4486
rect 7955 4452 7959 4486
rect 7959 4452 7989 4486
rect 8027 4452 8061 4486
rect 8099 4452 8129 4486
rect 8129 4452 8133 4486
rect 8171 4452 8197 4486
rect 8197 4452 8205 4486
rect 8243 4452 8265 4486
rect 8265 4452 8277 4486
rect 8315 4452 8333 4486
rect 8333 4452 8349 4486
rect 8387 4452 8401 4486
rect 8401 4452 8421 4486
rect 8459 4452 8469 4486
rect 8469 4452 8493 4486
rect 8531 4452 8537 4486
rect 8537 4452 8565 4486
rect 8603 4452 8605 4486
rect 8605 4452 8637 4486
rect 8675 4452 8707 4486
rect 8707 4452 8709 4486
rect 8747 4452 8775 4486
rect 8775 4452 8781 4486
rect 8819 4452 8843 4486
rect 8843 4452 8853 4486
rect 8891 4452 8911 4486
rect 8911 4452 8925 4486
rect 2625 4164 2659 4198
rect 9014 4196 9048 4230
rect 2625 4092 2659 4126
rect 3383 4121 3417 4155
rect 3455 4121 3489 4155
rect 7308 4040 7342 4074
rect 8666 4115 8700 4149
rect 8666 4043 8700 4077
rect 7308 3968 7342 4002
rect 7222 3897 7256 3931
rect 2889 3862 2923 3896
rect 2889 3790 2923 3824
rect 3061 3843 3095 3877
rect 3061 3771 3095 3805
rect 3466 3835 3500 3869
rect 3538 3835 3572 3869
rect 8486 3958 8520 3992
rect 7222 3825 7256 3859
rect 8486 3886 8520 3920
rect 8226 3830 8260 3864
rect 2554 3709 2588 3743
rect 2626 3709 2660 3743
rect 8226 3758 8260 3792
rect 8312 3838 8346 3872
rect 9014 4124 9048 4158
rect 8312 3766 8346 3800
rect 8754 3838 8788 3872
rect 8754 3766 8788 3800
rect 507 3472 519 3506
rect 519 3472 541 3506
rect 579 3472 587 3506
rect 587 3472 613 3506
rect 651 3472 655 3506
rect 655 3472 685 3506
rect 723 3472 757 3506
rect 795 3472 825 3506
rect 825 3472 829 3506
rect 867 3472 893 3506
rect 893 3472 901 3506
rect 939 3472 961 3506
rect 961 3472 973 3506
rect 1011 3472 1029 3506
rect 1029 3472 1045 3506
rect 1083 3472 1097 3506
rect 1097 3472 1117 3506
rect 1155 3472 1165 3506
rect 1165 3472 1189 3506
rect 1227 3472 1233 3506
rect 1233 3472 1261 3506
rect 1299 3472 1301 3506
rect 1301 3472 1333 3506
rect 1371 3472 1403 3506
rect 1403 3472 1405 3506
rect 1443 3472 1471 3506
rect 1471 3472 1477 3506
rect 1515 3472 1539 3506
rect 1539 3472 1549 3506
rect 1587 3472 1607 3506
rect 1607 3472 1621 3506
rect 1659 3472 1675 3506
rect 1675 3472 1693 3506
rect 1731 3472 1743 3506
rect 1743 3472 1765 3506
rect 1803 3472 1811 3506
rect 1811 3472 1837 3506
rect 1875 3472 1879 3506
rect 1879 3472 1909 3506
rect 1947 3472 1981 3506
rect 2019 3472 2049 3506
rect 2049 3472 2053 3506
rect 2091 3472 2117 3506
rect 2117 3472 2125 3506
rect 2163 3472 2185 3506
rect 2185 3472 2197 3506
rect 2235 3472 2253 3506
rect 2253 3472 2269 3506
rect 2307 3472 2321 3506
rect 2321 3472 2341 3506
rect 2379 3472 2389 3506
rect 2389 3472 2413 3506
rect 2451 3472 2457 3506
rect 2457 3472 2485 3506
rect 2523 3472 2525 3506
rect 2525 3472 2557 3506
rect 2595 3472 2627 3506
rect 2627 3472 2629 3506
rect 2667 3472 2695 3506
rect 2695 3472 2701 3506
rect 2739 3472 2763 3506
rect 2763 3472 2773 3506
rect 2811 3472 2831 3506
rect 2831 3472 2845 3506
rect 2883 3472 2899 3506
rect 2899 3472 2917 3506
rect 2955 3472 2967 3506
rect 2967 3472 2989 3506
rect 3027 3472 3035 3506
rect 3035 3472 3061 3506
rect 3099 3472 3103 3506
rect 3103 3472 3133 3506
rect 3171 3472 3205 3506
rect 3243 3472 3273 3506
rect 3273 3472 3277 3506
rect 3315 3472 3341 3506
rect 3341 3472 3349 3506
rect 3387 3472 3409 3506
rect 3409 3472 3421 3506
rect 3459 3472 3477 3506
rect 3477 3472 3493 3506
rect 3531 3472 3545 3506
rect 3545 3472 3565 3506
rect 3603 3472 3613 3506
rect 3613 3472 3637 3506
rect 3675 3472 3681 3506
rect 3681 3472 3709 3506
rect 3747 3472 3749 3506
rect 3749 3472 3781 3506
rect 3819 3472 3851 3506
rect 3851 3472 3853 3506
rect 3891 3472 3919 3506
rect 3919 3472 3925 3506
rect 3963 3472 3987 3506
rect 3987 3472 3997 3506
rect 4035 3472 4055 3506
rect 4055 3472 4069 3506
rect 4107 3472 4123 3506
rect 4123 3472 4141 3506
rect 4179 3472 4191 3506
rect 4191 3472 4213 3506
rect 4251 3472 4259 3506
rect 4259 3472 4285 3506
rect 4323 3472 4327 3506
rect 4327 3472 4357 3506
rect 4395 3472 4429 3506
rect 4467 3472 4497 3506
rect 4497 3472 4501 3506
rect 4539 3472 4565 3506
rect 4565 3472 4573 3506
rect 4611 3472 4633 3506
rect 4633 3472 4645 3506
rect 4683 3472 4701 3506
rect 4701 3472 4717 3506
rect 4755 3472 4769 3506
rect 4769 3472 4789 3506
rect 4827 3472 4837 3506
rect 4837 3472 4861 3506
rect 4899 3472 4905 3506
rect 4905 3472 4933 3506
rect 4971 3472 4973 3506
rect 4973 3472 5005 3506
rect 5043 3472 5075 3506
rect 5075 3472 5077 3506
rect 5115 3472 5143 3506
rect 5143 3472 5149 3506
rect 5187 3472 5211 3506
rect 5211 3472 5221 3506
rect 5259 3472 5279 3506
rect 5279 3472 5293 3506
rect 5331 3472 5347 3506
rect 5347 3472 5365 3506
rect 5403 3472 5415 3506
rect 5415 3472 5437 3506
rect 5475 3472 5483 3506
rect 5483 3472 5509 3506
rect 5547 3472 5551 3506
rect 5551 3472 5581 3506
rect 5619 3472 5653 3506
rect 5691 3472 5721 3506
rect 5721 3472 5725 3506
rect 5763 3472 5789 3506
rect 5789 3472 5797 3506
rect 5835 3472 5857 3506
rect 5857 3472 5869 3506
rect 5907 3472 5925 3506
rect 5925 3472 5941 3506
rect 5979 3472 5993 3506
rect 5993 3472 6013 3506
rect 6051 3472 6061 3506
rect 6061 3472 6085 3506
rect 6123 3472 6129 3506
rect 6129 3472 6157 3506
rect 6195 3472 6197 3506
rect 6197 3472 6229 3506
rect 6267 3472 6299 3506
rect 6299 3472 6301 3506
rect 6339 3472 6367 3506
rect 6367 3472 6373 3506
rect 6411 3472 6435 3506
rect 6435 3472 6445 3506
rect 6483 3472 6503 3506
rect 6503 3472 6517 3506
rect 6555 3472 6571 3506
rect 6571 3472 6589 3506
rect 6627 3472 6639 3506
rect 6639 3472 6661 3506
rect 6699 3472 6707 3506
rect 6707 3472 6733 3506
rect 6771 3472 6775 3506
rect 6775 3472 6805 3506
rect 6843 3472 6877 3506
rect 6915 3472 6945 3506
rect 6945 3472 6949 3506
rect 6987 3472 7013 3506
rect 7013 3472 7021 3506
rect 7059 3472 7081 3506
rect 7081 3472 7093 3506
rect 7131 3472 7149 3506
rect 7149 3472 7165 3506
rect 7203 3472 7217 3506
rect 7217 3472 7237 3506
rect 7275 3472 7285 3506
rect 7285 3472 7309 3506
rect 7347 3472 7353 3506
rect 7353 3472 7381 3506
rect 7419 3472 7421 3506
rect 7421 3472 7453 3506
rect 7491 3472 7523 3506
rect 7523 3472 7525 3506
rect 7563 3472 7591 3506
rect 7591 3472 7597 3506
rect 7635 3472 7659 3506
rect 7659 3472 7669 3506
rect 7707 3472 7727 3506
rect 7727 3472 7741 3506
rect 7779 3472 7795 3506
rect 7795 3472 7813 3506
rect 7851 3472 7863 3506
rect 7863 3472 7885 3506
rect 7923 3472 7931 3506
rect 7931 3472 7957 3506
rect 7995 3472 7999 3506
rect 7999 3472 8029 3506
rect 8067 3472 8101 3506
rect 8139 3472 8169 3506
rect 8169 3472 8173 3506
rect 8211 3472 8237 3506
rect 8237 3472 8245 3506
rect 8283 3472 8305 3506
rect 8305 3472 8317 3506
rect 8355 3472 8373 3506
rect 8373 3472 8389 3506
rect 8427 3472 8441 3506
rect 8441 3472 8461 3506
rect 8499 3472 8509 3506
rect 8509 3472 8533 3506
rect 8571 3472 8577 3506
rect 8577 3472 8605 3506
<< metal1 >>
rect 455 4486 8972 4498
rect 455 4452 467 4486
rect 501 4452 539 4486
rect 573 4452 611 4486
rect 645 4452 683 4486
rect 717 4452 755 4486
rect 789 4452 827 4486
rect 861 4452 899 4486
rect 933 4452 971 4486
rect 1005 4452 1043 4486
rect 1077 4452 1115 4486
rect 1149 4452 1187 4486
rect 1221 4452 1259 4486
rect 1293 4452 1331 4486
rect 1365 4452 1403 4486
rect 1437 4452 1475 4486
rect 1509 4452 1547 4486
rect 1581 4452 1619 4486
rect 1653 4452 1691 4486
rect 1725 4452 1763 4486
rect 1797 4452 1835 4486
rect 1869 4452 1907 4486
rect 1941 4452 1979 4486
rect 2013 4452 2051 4486
rect 2085 4452 2123 4486
rect 2157 4452 2195 4486
rect 2229 4452 2267 4486
rect 2301 4452 2339 4486
rect 2373 4452 2411 4486
rect 2445 4452 2483 4486
rect 2517 4452 2555 4486
rect 2589 4452 2627 4486
rect 2661 4452 2699 4486
rect 2733 4452 2771 4486
rect 2805 4452 2843 4486
rect 2877 4452 2915 4486
rect 2949 4452 2987 4486
rect 3021 4452 3059 4486
rect 3093 4452 3131 4486
rect 3165 4452 3203 4486
rect 3237 4452 3275 4486
rect 3309 4452 3347 4486
rect 3381 4452 3419 4486
rect 3453 4452 3491 4486
rect 3525 4452 3563 4486
rect 3597 4452 3635 4486
rect 3669 4452 3707 4486
rect 3741 4452 3779 4486
rect 3813 4452 3851 4486
rect 3885 4452 3923 4486
rect 3957 4452 3995 4486
rect 4029 4452 4067 4486
rect 4101 4452 4139 4486
rect 4173 4452 4211 4486
rect 4245 4452 4283 4486
rect 4317 4452 4355 4486
rect 4389 4452 4427 4486
rect 4461 4452 4499 4486
rect 4533 4452 4571 4486
rect 4605 4452 4643 4486
rect 4677 4452 4715 4486
rect 4749 4452 4787 4486
rect 4821 4452 4859 4486
rect 4893 4452 4931 4486
rect 4965 4452 5003 4486
rect 5037 4452 5075 4486
rect 5109 4452 5147 4486
rect 5181 4452 5219 4486
rect 5253 4452 5291 4486
rect 5325 4452 5363 4486
rect 5397 4452 5435 4486
rect 5469 4452 5507 4486
rect 5541 4452 5579 4486
rect 5613 4452 5651 4486
rect 5685 4452 5723 4486
rect 5757 4452 5795 4486
rect 5829 4452 5867 4486
rect 5901 4452 5939 4486
rect 5973 4452 6011 4486
rect 6045 4452 6083 4486
rect 6117 4452 6155 4486
rect 6189 4452 6227 4486
rect 6261 4452 6299 4486
rect 6333 4452 6371 4486
rect 6405 4452 6443 4486
rect 6477 4452 6515 4486
rect 6549 4452 6587 4486
rect 6621 4452 6659 4486
rect 6693 4452 6731 4486
rect 6765 4452 6803 4486
rect 6837 4452 6875 4486
rect 6909 4452 6947 4486
rect 6981 4452 7019 4486
rect 7053 4452 7091 4486
rect 7125 4452 7163 4486
rect 7197 4452 7235 4486
rect 7269 4452 7307 4486
rect 7341 4452 7379 4486
rect 7413 4452 7451 4486
rect 7485 4452 7523 4486
rect 7557 4452 7595 4486
rect 7629 4452 7667 4486
rect 7701 4452 7739 4486
rect 7773 4452 7811 4486
rect 7845 4452 7883 4486
rect 7917 4452 7955 4486
rect 7989 4452 8027 4486
rect 8061 4452 8099 4486
rect 8133 4452 8171 4486
rect 8205 4452 8243 4486
rect 8277 4452 8315 4486
rect 8349 4452 8387 4486
rect 8421 4452 8459 4486
rect 8493 4452 8531 4486
rect 8565 4452 8603 4486
rect 8637 4452 8675 4486
rect 8709 4452 8747 4486
rect 8781 4452 8819 4486
rect 8853 4452 8891 4486
rect 8925 4452 8972 4486
rect 455 4440 8972 4452
rect 2709 4335 2832 4438
rect 3200 4296 3266 4440
rect 3501 4295 3566 4440
rect 7145 4296 7209 4440
rect 8149 4295 8214 4440
rect 8976 4295 9041 4498
rect 2619 4198 2665 4210
rect 3684 4201 5050 4253
rect 5102 4201 5114 4253
rect 5166 4201 5172 4253
rect 2619 4164 2625 4198
rect 2659 4167 2665 4198
rect 5874 4196 5880 4248
rect 5932 4196 5944 4248
rect 5996 4242 6002 4248
tri 6002 4242 6008 4248 sw
rect 5996 4230 9054 4242
rect 5996 4196 9014 4230
rect 9048 4196 9054 4230
tri 2665 4167 2694 4196 sw
tri 8974 4167 9003 4196 ne
rect 9003 4167 9054 4196
rect 2659 4164 2694 4167
rect 2619 4161 2694 4164
tri 2694 4161 2700 4167 sw
tri 4791 4161 4797 4167 se
rect 4797 4161 4803 4167
rect 2619 4158 2700 4161
tri 2700 4158 2703 4161 sw
rect 2619 4155 2703 4158
tri 2703 4155 2706 4158 sw
rect 3371 4155 4803 4161
rect 2619 4126 2706 4155
rect 2619 4092 2625 4126
rect 2659 4121 2706 4126
tri 2706 4121 2740 4155 sw
rect 3371 4121 3383 4155
rect 3417 4121 3455 4155
rect 3489 4121 4803 4155
rect 2659 4115 2740 4121
tri 2740 4115 2746 4121 sw
rect 3371 4115 4803 4121
rect 4855 4115 4867 4167
rect 4919 4161 4925 4167
tri 4925 4161 4931 4167 sw
tri 9003 4162 9008 4167 ne
rect 4919 4149 8706 4161
rect 4919 4115 8666 4149
rect 8700 4115 8706 4149
rect 2659 4092 2746 4115
rect 2619 4086 2746 4092
tri 2746 4086 2775 4115 sw
tri 8626 4086 8655 4115 ne
rect 8655 4086 8706 4115
rect 9008 4158 9054 4167
rect 9008 4124 9014 4158
rect 9048 4124 9054 4158
rect 9008 4112 9054 4124
rect 2619 4080 7348 4086
tri 8655 4081 8660 4086 ne
tri 2684 4077 2687 4080 ne
rect 2687 4077 7348 4080
tri 2687 4074 2690 4077 ne
rect 2690 4074 7348 4077
tri 2690 4058 2706 4074 ne
rect 2706 4058 7308 4074
tri 7268 4040 7286 4058 ne
rect 7286 4040 7308 4058
rect 7342 4040 7348 4074
tri 7286 4024 7302 4040 ne
rect 7302 4002 7348 4040
rect 8660 4077 8706 4086
rect 8660 4043 8666 4077
rect 8700 4043 8706 4077
rect 8660 4031 8706 4043
rect 7302 3968 7308 4002
rect 7342 3968 7348 4002
tri 8475 3992 8480 3997 se
rect 8480 3992 8526 4004
tri 3553 3961 3559 3967 sw
tri 5658 3961 5664 3967 se
tri 5792 3961 5798 3967 sw
rect 3552 3915 3701 3961
rect 3703 3915 3707 3961
rect 4188 3915 4352 3961
rect 5597 3915 5608 3961
rect 5613 3915 5806 3961
rect 5811 3915 5854 3961
rect 7302 3956 7348 3968
tri 8444 3961 8475 3992 se
rect 8475 3961 8486 3992
rect 8008 3958 8486 3961
rect 8520 3958 8526 3992
rect 7216 3931 7262 3943
tri 4272 3908 4279 3915 ne
rect 4279 3908 4352 3915
rect 2883 3896 2929 3908
tri 4279 3897 4290 3908 ne
rect 4290 3897 4352 3908
tri 4352 3897 4364 3909 sw
rect 7216 3897 7222 3931
rect 7256 3915 7262 3931
rect 8008 3920 8526 3958
tri 7262 3915 7266 3919 sw
rect 8008 3915 8486 3920
rect 7256 3897 7266 3915
rect 2883 3862 2889 3896
rect 2923 3862 2929 3896
tri 4290 3889 4298 3897 ne
rect 4298 3889 4364 3897
rect 2883 3842 2929 3862
rect 2456 3824 2929 3842
rect 2456 3790 2889 3824
rect 2923 3790 2929 3824
rect 2456 3778 2929 3790
rect 3055 3877 3101 3889
tri 4298 3886 4301 3889 ne
rect 4301 3886 4364 3889
tri 4364 3886 4375 3897 sw
rect 7216 3886 7266 3897
tri 7266 3886 7295 3915 sw
tri 8444 3886 8473 3915 ne
rect 8473 3886 8486 3915
rect 8520 3886 8526 3920
tri 4301 3882 4305 3886 ne
rect 4305 3882 4375 3886
tri 4186 3881 4187 3882 se
tri 4305 3881 4306 3882 ne
rect 3055 3843 3061 3877
rect 3095 3843 3101 3877
tri 4180 3875 4186 3881 se
rect 4186 3875 4187 3881
rect 4306 3875 4375 3882
tri 4375 3875 4386 3886 sw
rect 7216 3884 7295 3886
tri 7295 3884 7297 3886 sw
tri 8473 3884 8475 3886 ne
rect 8475 3884 8526 3886
rect 7216 3876 7297 3884
tri 7297 3876 7305 3884 sw
rect 7216 3875 7305 3876
tri 7305 3875 7306 3876 sw
rect 3055 3805 3101 3843
rect 3454 3869 3602 3875
rect 3454 3835 3466 3869
rect 3500 3835 3538 3869
rect 3572 3835 3602 3869
rect 3454 3829 3602 3835
rect 5700 3829 5714 3875
rect 7216 3859 7527 3875
rect 7216 3825 7222 3859
rect 7256 3829 7527 3859
rect 8217 3870 8269 3876
rect 7256 3825 7262 3829
rect 7216 3813 7262 3825
tri 7262 3813 7278 3829 nw
rect 2446 3771 2453 3778
tri 2453 3771 2460 3778 nw
rect 3055 3771 3061 3805
rect 3095 3771 3101 3805
rect 2446 3770 2452 3771
tri 2452 3770 2453 3771 nw
rect 3055 3759 3101 3771
rect 8217 3804 8269 3818
tri 3355 3749 3361 3755 se
rect 3361 3749 3968 3755
rect 2542 3746 2672 3749
tri 2672 3746 2675 3749 sw
tri 3352 3746 3355 3749 se
rect 3355 3746 3968 3749
rect 2542 3743 2675 3746
rect 2542 3709 2554 3743
rect 2588 3709 2626 3743
rect 2660 3731 2675 3743
tri 2675 3731 2690 3746 sw
tri 3337 3731 3352 3746 se
rect 3352 3731 3968 3746
rect 2660 3709 3968 3731
rect 2542 3703 3968 3709
rect 4020 3703 4032 3755
rect 4084 3703 4090 3755
rect 8306 3874 8352 3884
tri 8475 3879 8480 3884 ne
tri 8352 3874 8354 3876 sw
rect 8480 3874 8526 3884
tri 8746 3874 8748 3876 se
rect 8748 3874 8794 3884
rect 8306 3872 8354 3874
tri 8354 3872 8356 3874 sw
tri 8744 3872 8746 3874 se
rect 8746 3872 8794 3874
rect 8306 3838 8312 3872
rect 8346 3842 8356 3872
tri 8356 3842 8386 3872 sw
tri 8714 3842 8744 3872 se
rect 8744 3842 8754 3872
rect 8346 3838 8754 3842
rect 8788 3838 8794 3872
rect 8306 3800 8794 3838
rect 8306 3766 8312 3800
rect 8346 3796 8754 3800
rect 8346 3766 8356 3796
tri 8356 3766 8386 3796 nw
tri 8714 3766 8744 3796 ne
rect 8744 3766 8754 3796
rect 8788 3766 8794 3800
rect 8306 3754 8352 3766
tri 8352 3762 8356 3766 nw
tri 8744 3762 8748 3766 ne
rect 8748 3754 8794 3766
rect 8217 3746 8269 3752
rect 2754 3518 2929 3557
rect 3200 3518 3230 3675
rect 3542 3518 3545 3675
rect 7145 3518 7168 3674
rect 8149 3518 8214 3675
rect 495 3506 8687 3518
rect 495 3472 507 3506
rect 541 3472 579 3506
rect 613 3472 651 3506
rect 685 3472 723 3506
rect 757 3472 795 3506
rect 829 3472 867 3506
rect 901 3472 939 3506
rect 973 3472 1011 3506
rect 1045 3472 1083 3506
rect 1117 3472 1155 3506
rect 1189 3472 1227 3506
rect 1261 3472 1299 3506
rect 1333 3472 1371 3506
rect 1405 3472 1443 3506
rect 1477 3472 1515 3506
rect 1549 3472 1587 3506
rect 1621 3472 1659 3506
rect 1693 3472 1731 3506
rect 1765 3472 1803 3506
rect 1837 3472 1875 3506
rect 1909 3472 1947 3506
rect 1981 3472 2019 3506
rect 2053 3472 2091 3506
rect 2125 3472 2163 3506
rect 2197 3472 2235 3506
rect 2269 3472 2307 3506
rect 2341 3472 2379 3506
rect 2413 3472 2451 3506
rect 2485 3472 2523 3506
rect 2557 3472 2595 3506
rect 2629 3472 2667 3506
rect 2701 3472 2739 3506
rect 2773 3472 2811 3506
rect 2845 3472 2883 3506
rect 2917 3472 2955 3506
rect 2989 3472 3027 3506
rect 3061 3472 3099 3506
rect 3133 3472 3171 3506
rect 3205 3472 3243 3506
rect 3277 3472 3315 3506
rect 3349 3472 3387 3506
rect 3421 3472 3459 3506
rect 3493 3472 3531 3506
rect 3565 3472 3603 3506
rect 3637 3472 3675 3506
rect 3709 3472 3747 3506
rect 3781 3472 3819 3506
rect 3853 3472 3891 3506
rect 3925 3472 3963 3506
rect 3997 3472 4035 3506
rect 4069 3472 4107 3506
rect 4141 3472 4179 3506
rect 4213 3472 4251 3506
rect 4285 3472 4323 3506
rect 4357 3472 4395 3506
rect 4429 3472 4467 3506
rect 4501 3472 4539 3506
rect 4573 3472 4611 3506
rect 4645 3472 4683 3506
rect 4717 3472 4755 3506
rect 4789 3472 4827 3506
rect 4861 3472 4899 3506
rect 4933 3472 4971 3506
rect 5005 3472 5043 3506
rect 5077 3472 5115 3506
rect 5149 3472 5187 3506
rect 5221 3472 5259 3506
rect 5293 3472 5331 3506
rect 5365 3472 5403 3506
rect 5437 3472 5475 3506
rect 5509 3472 5547 3506
rect 5581 3472 5619 3506
rect 5653 3472 5691 3506
rect 5725 3472 5763 3506
rect 5797 3472 5835 3506
rect 5869 3472 5907 3506
rect 5941 3472 5979 3506
rect 6013 3472 6051 3506
rect 6085 3472 6123 3506
rect 6157 3472 6195 3506
rect 6229 3472 6267 3506
rect 6301 3472 6339 3506
rect 6373 3472 6411 3506
rect 6445 3472 6483 3506
rect 6517 3472 6555 3506
rect 6589 3472 6627 3506
rect 6661 3472 6699 3506
rect 6733 3472 6771 3506
rect 6805 3472 6843 3506
rect 6877 3472 6915 3506
rect 6949 3472 6987 3506
rect 7021 3472 7059 3506
rect 7093 3472 7131 3506
rect 7165 3472 7203 3506
rect 7237 3472 7275 3506
rect 7309 3472 7347 3506
rect 7381 3472 7419 3506
rect 7453 3472 7491 3506
rect 7525 3472 7563 3506
rect 7597 3472 7635 3506
rect 7669 3472 7707 3506
rect 7741 3472 7779 3506
rect 7813 3472 7851 3506
rect 7885 3472 7923 3506
rect 7957 3472 7995 3506
rect 8029 3472 8067 3506
rect 8101 3472 8139 3506
rect 8173 3472 8211 3506
rect 8245 3472 8283 3506
rect 8317 3472 8355 3506
rect 8389 3472 8427 3506
rect 8461 3472 8499 3506
rect 8533 3472 8571 3506
rect 8605 3472 8687 3506
rect 495 3460 8687 3472
rect 8976 3460 9000 3675
rect 5044 3215 5050 3267
rect 5102 3215 5114 3267
rect 5166 3215 5172 3267
rect 4118 2623 4170 2629
tri 4082 2553 4118 2589 se
rect 4671 2610 4723 2616
rect 4118 2559 4170 2571
tri 4170 2553 4200 2583 sw
tri 5797 2586 5803 2592 se
rect 4118 2501 4170 2507
rect 4671 2540 4723 2558
rect 5803 2540 5809 2592
rect 5861 2540 5873 2592
rect 5925 2540 5931 2592
tri 5931 2586 5937 2592 sw
rect 4671 2482 4723 2488
tri 4097 1871 4131 1905 ne
rect 4131 1810 4183 1905
tri 4183 1871 4217 1905 nw
tri 4322 1607 4331 1616 se
rect 4331 1607 4377 1648
rect 4088 1601 4140 1607
tri 4300 1585 4322 1607 se
rect 4322 1596 4377 1607
rect 4322 1585 4336 1596
tri 4140 1555 4170 1585 sw
tri 4270 1555 4300 1585 se
rect 4300 1555 4336 1585
tri 4336 1555 4377 1596 nw
rect 4140 1549 4290 1555
rect 4088 1537 4290 1549
rect 4140 1509 4290 1537
tri 4290 1509 4336 1555 nw
rect 4088 1479 4140 1485
tri 4140 1479 4170 1509 nw
rect 4824 1247 5182 1360
<< rmetal1 >>
rect 3701 3915 3703 3961
rect 5608 3915 5613 3961
rect 5806 3915 5811 3961
<< via1 >>
rect 5050 4201 5102 4253
rect 5114 4201 5166 4253
rect 5880 4196 5932 4248
rect 5944 4196 5996 4248
rect 4803 4115 4855 4167
rect 4867 4115 4919 4167
rect 8217 3864 8269 3870
rect 8217 3830 8226 3864
rect 8226 3830 8260 3864
rect 8260 3830 8269 3864
rect 8217 3818 8269 3830
rect 8217 3792 8269 3804
rect 8217 3758 8226 3792
rect 8226 3758 8260 3792
rect 8260 3758 8269 3792
rect 3968 3703 4020 3755
rect 4032 3703 4084 3755
rect 8217 3752 8269 3758
rect 5050 3215 5102 3267
rect 5114 3215 5166 3267
rect 4118 2571 4170 2623
rect 4118 2507 4170 2559
rect 4671 2558 4723 2610
rect 5809 2540 5861 2592
rect 5873 2540 5925 2592
rect 4671 2488 4723 2540
rect 4088 1549 4140 1601
rect 4088 1485 4140 1537
<< metal2 >>
tri 3556 4196 3561 4201 ne
rect 3561 4196 3614 4201
tri 3561 4182 3575 4196 ne
rect 3575 4182 3614 4196
rect 3665 4196 3679 4201
tri 3679 4196 3684 4201 nw
rect 3665 4183 3666 4196
tri 3666 4183 3679 4196 nw
tri 3665 4182 3666 4183 nw
tri 3575 4167 3590 4182 ne
rect 3590 4167 3614 4182
tri 3590 4143 3614 4167 ne
rect 4110 4025 4162 4213
rect 5044 4201 5050 4253
rect 5102 4201 5114 4253
rect 5166 4201 5172 4253
tri 5044 4196 5049 4201 ne
rect 5049 4196 5156 4201
tri 5156 4196 5161 4201 nw
rect 5874 4196 5880 4248
rect 5932 4196 5944 4248
rect 5996 4196 6002 4248
tri 5049 4170 5075 4196 ne
rect 5075 4183 5143 4196
tri 5143 4183 5156 4196 nw
tri 5875 4183 5888 4196 ne
rect 5888 4183 5962 4196
rect 4797 4115 4803 4167
rect 4855 4115 4867 4167
rect 4919 4115 4925 4167
tri 4162 4025 4170 4033 sw
rect 4110 4011 4170 4025
tri 4110 4003 4118 4011 ne
rect 3962 3703 3968 3755
rect 4020 3703 4032 3755
rect 4084 3703 4090 3755
tri 3983 3648 4038 3703 ne
rect 4038 2399 4090 3703
rect 4118 2623 4170 4011
tri 4787 3818 4797 3828 se
rect 4797 3818 4851 4115
tri 4851 4081 4885 4115 nw
tri 4773 3804 4787 3818 se
rect 4787 3804 4851 3818
tri 4744 3775 4773 3804 se
rect 4773 3775 4851 3804
rect 4744 3723 4851 3775
rect 4118 2559 4170 2571
rect 4118 2501 4170 2507
tri 4671 2773 4744 2846 se
rect 4744 2824 4796 3723
tri 4796 3668 4851 3723 nw
tri 5044 3267 5075 3298 se
rect 5075 3267 5127 4183
tri 5127 4167 5143 4183 nw
tri 5888 4167 5904 4183 ne
rect 5904 4167 5962 4183
tri 5904 4161 5910 4167 ne
tri 5127 3267 5161 3301 sw
rect 5044 3215 5050 3267
rect 5102 3215 5114 3267
rect 5166 3215 5172 3267
rect 4744 2773 4745 2824
tri 4745 2773 4796 2824 nw
tri 5844 2857 5910 2923 se
rect 5910 2901 5962 4167
tri 5962 4161 5997 4196 nw
rect 8217 3870 8269 3876
rect 8217 3804 8269 3818
rect 8217 3746 8269 3752
rect 5910 2857 5918 2901
tri 5918 2857 5962 2901 nw
rect 4671 2610 4723 2773
tri 4723 2751 4745 2773 nw
tri 5809 2592 5844 2627 se
rect 5844 2592 5896 2857
tri 5896 2835 5918 2857 nw
tri 5896 2592 5931 2627 sw
rect 4671 2540 4723 2558
rect 5803 2540 5809 2592
rect 5861 2540 5873 2592
rect 5925 2540 5931 2592
rect 4671 2482 4723 2488
tri 4038 2371 4066 2399 ne
rect 4066 2371 4090 2399
tri 4090 2371 4140 2421 sw
tri 4066 2349 4088 2371 ne
rect 4088 1601 4140 2371
rect 4088 1537 4140 1549
rect 4088 1479 4140 1485
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1645210163
transform -1 0 2910 0 1 3436
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1645210163
transform -1 0 7506 0 1 3436
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_2
timestamp 1645210163
transform 1 0 3204 0 1 3436
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x4  sky130_fd_io__hvsbt_inv_x4_0
timestamp 1645210163
transform 1 0 7324 0 1 3436
box -42 24 913 1116
use sky130_fd_io__hvsbt_inv_x4  sky130_fd_io__hvsbt_inv_x4_1
timestamp 1645210163
transform 1 0 3504 0 1 3436
box -42 24 913 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1645210163
transform 1 0 8504 0 1 3436
box 0 24 534 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_1
timestamp 1645210163
transform -1 0 8686 0 1 3436
box 0 24 534 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1645210163
transform 1 0 2728 0 1 3436
box -42 24 569 1116
use sky130_fd_io__hvsbt_inv_x8  sky130_fd_io__hvsbt_inv_x8_0
timestamp 1645210163
transform 1 0 5616 0 1 3436
box -42 24 1632 1116
use sky130_fd_io__com_ctl_ls  sky130_fd_io__com_ctl_ls_0
timestamp 1645210163
transform -1 0 6098 0 -1 3226
box -71 10 2077 2019
use sky130_fd_io__hvsbt_inv_x8v2  sky130_fd_io__hvsbt_inv_x8v2_0
timestamp 1645210163
transform 1 0 4208 0 1 3436
box -42 24 1632 1116
<< labels >>
flabel metal2 s 4128 4183 4156 4207 3 FreeSans 520 0 0 0 HLD_OVR
port 1 nsew
flabel metal1 s 5581 2998 5581 2998 0 FreeSans 440 0 0 0 VCC_IO
port 2 nsew
flabel metal1 s 2709 4335 2832 4438 3 FreeSans 520 0 0 0 VCC_IO
port 2 nsew
flabel metal1 s 2754 3479 2929 3557 3 FreeSans 520 0 0 0 VGND
port 3 nsew
flabel metal1 s 5639 3921 5793 3954 3 FreeSans 520 0 0 0 HLD_I_H_N
port 4 nsew
flabel metal1 s 8026 3927 8091 3951 3 FreeSans 520 0 0 0 OD_I_H
port 5 nsew
flabel metal1 s 5725 1995 5725 1995 0 FreeSans 440 0 0 0 VGND
port 3 nsew
flabel metal1 s 5699 2830 5699 2830 0 FreeSans 440 0 0 0 VPWR
port 6 nsew
flabel metal1 s 4824 1247 5182 1360 3 FreeSans 520 0 0 0 VPWR
port 6 nsew
flabel metal1 s 3552 3915 3606 3961 3 FreeSans 520 0 0 0 HLD_I_H
port 7 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 8052828
string GDS_START 8008754
<< end >>
