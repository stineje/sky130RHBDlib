magic
tech sky130A
magscale 1 2
timestamp 1648064704
<< metal1 >>
rect 867 649 1057 683
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 1110 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 814 0 -1 666
box -53 -33 29 33
use nand3x1_pcell  nand3x1_pcell_0
timestamp 1648064657
transform 1 0 0 0 1 0
box -84 0 1046 1575
use invx1_pcell  invx1_pcell_0
timestamp 1648064504
transform 1 0 962 0 1 0
box -84 0 528 1575
<< end >>
