magic
tech sky130A
magscale 1 2
timestamp 1669564290
<< nwell >>
rect -87 786 4379 1550
<< pwell >>
rect -34 -34 4326 544
<< nmos >>
rect 147 290 177 351
tri 177 290 193 306 sw
rect 447 290 477 351
rect 147 260 253 290
tri 253 260 283 290 sw
rect 147 159 177 260
tri 177 244 193 260 nw
tri 237 244 253 260 ne
tri 177 159 193 175 sw
tri 237 159 253 175 se
rect 253 159 283 260
tri 342 260 372 290 se
rect 372 260 477 290
rect 342 166 372 260
tri 372 244 388 260 nw
tri 431 244 447 260 ne
tri 372 166 388 182 sw
tri 431 166 447 182 se
rect 447 166 477 260
tri 147 129 177 159 ne
rect 177 129 253 159
tri 253 129 283 159 nw
tri 342 136 372 166 ne
rect 372 136 447 166
tri 447 136 477 166 nw
rect 649 298 679 351
tri 679 298 695 314 sw
rect 649 268 755 298
tri 755 268 785 298 sw
rect 649 167 679 268
tri 679 252 695 268 nw
tri 739 252 755 268 ne
tri 679 167 695 183 sw
tri 739 167 755 183 se
rect 755 167 785 268
tri 649 137 679 167 ne
rect 679 137 755 167
tri 755 137 785 167 nw
rect 1130 288 1160 349
tri 1160 288 1176 304 sw
rect 1324 296 1354 349
tri 1354 296 1370 312 sw
rect 1130 258 1236 288
tri 1236 258 1266 288 sw
rect 1324 266 1430 296
tri 1430 266 1460 296 sw
rect 1130 157 1160 258
tri 1160 242 1176 258 nw
tri 1220 242 1236 258 ne
tri 1160 157 1176 173 sw
tri 1220 157 1236 173 se
rect 1236 157 1266 258
rect 1324 165 1354 266
tri 1354 250 1370 266 nw
tri 1414 250 1430 266 ne
tri 1354 165 1370 181 sw
tri 1414 165 1430 181 se
rect 1430 165 1460 266
tri 1130 127 1160 157 ne
rect 1160 127 1236 157
tri 1236 127 1266 157 nw
tri 1324 135 1354 165 ne
rect 1354 135 1430 165
tri 1430 135 1460 165 nw
rect 1796 288 1826 349
tri 1826 288 1842 304 sw
rect 1990 296 2020 349
tri 2020 296 2036 312 sw
rect 1796 258 1902 288
tri 1902 258 1932 288 sw
rect 1990 266 2096 296
tri 2096 266 2126 296 sw
rect 1796 157 1826 258
tri 1826 242 1842 258 nw
tri 1886 242 1902 258 ne
tri 1826 157 1842 173 sw
tri 1886 157 1902 173 se
rect 1902 157 1932 258
rect 1990 165 2020 266
tri 2020 250 2036 266 nw
tri 2080 250 2096 266 ne
tri 2020 165 2036 181 sw
tri 2080 165 2096 181 se
rect 2096 165 2126 266
tri 1796 127 1826 157 ne
rect 1826 127 1902 157
tri 1902 127 1932 157 nw
tri 1990 135 2020 165 ne
rect 2020 135 2096 165
tri 2096 135 2126 165 nw
rect 2462 288 2492 349
tri 2492 288 2508 304 sw
rect 2656 296 2686 349
tri 2686 296 2702 312 sw
rect 2462 258 2568 288
tri 2568 258 2598 288 sw
rect 2656 266 2762 296
tri 2762 266 2792 296 sw
rect 2462 157 2492 258
tri 2492 242 2508 258 nw
tri 2552 242 2568 258 ne
tri 2492 157 2508 173 sw
tri 2552 157 2568 173 se
rect 2568 157 2598 258
rect 2656 165 2686 266
tri 2686 250 2702 266 nw
tri 2746 250 2762 266 ne
tri 2686 165 2702 181 sw
tri 2746 165 2762 181 se
rect 2762 165 2792 266
tri 2462 127 2492 157 ne
rect 2492 127 2568 157
tri 2568 127 2598 157 nw
tri 2656 135 2686 165 ne
rect 2686 135 2762 165
tri 2762 135 2792 165 nw
rect 3128 288 3158 349
tri 3158 288 3174 304 sw
rect 3322 296 3352 349
tri 3352 296 3368 312 sw
rect 3128 258 3234 288
tri 3234 258 3264 288 sw
rect 3322 266 3428 296
tri 3428 266 3458 296 sw
rect 3128 157 3158 258
tri 3158 242 3174 258 nw
tri 3218 242 3234 258 ne
tri 3158 157 3174 173 sw
tri 3218 157 3234 173 se
rect 3234 157 3264 258
rect 3322 165 3352 266
tri 3352 250 3368 266 nw
tri 3412 250 3428 266 ne
tri 3352 165 3368 181 sw
tri 3412 165 3428 181 se
rect 3428 165 3458 266
tri 3128 127 3158 157 ne
rect 3158 127 3234 157
tri 3234 127 3264 157 nw
tri 3322 135 3352 165 ne
rect 3352 135 3428 165
tri 3428 135 3458 165 nw
rect 3794 288 3824 349
tri 3824 288 3840 304 sw
rect 3988 296 4018 349
tri 4018 296 4034 312 sw
rect 3794 258 3900 288
tri 3900 258 3930 288 sw
rect 3988 266 4094 296
tri 4094 266 4124 296 sw
rect 3794 157 3824 258
tri 3824 242 3840 258 nw
tri 3884 242 3900 258 ne
tri 3824 157 3840 173 sw
tri 3884 157 3900 173 se
rect 3900 157 3930 258
rect 3988 165 4018 266
tri 4018 250 4034 266 nw
tri 4078 250 4094 266 ne
tri 4018 165 4034 181 sw
tri 4078 165 4094 181 se
rect 4094 165 4124 266
tri 3794 127 3824 157 ne
rect 3824 127 3900 157
tri 3900 127 3930 157 nw
tri 3988 135 4018 165 ne
rect 4018 135 4094 165
tri 4094 135 4124 165 nw
<< pmos >>
rect 247 1004 277 1404
rect 335 1004 365 1404
rect 423 1004 453 1404
rect 511 1004 541 1404
rect 599 1004 629 1404
rect 687 1004 717 1404
rect 1149 1004 1179 1404
rect 1237 1004 1267 1404
rect 1325 1004 1355 1404
rect 1413 1004 1443 1404
rect 1815 1004 1845 1404
rect 1903 1004 1933 1404
rect 1991 1004 2021 1404
rect 2079 1004 2109 1404
rect 2481 1004 2511 1404
rect 2569 1004 2599 1404
rect 2657 1004 2687 1404
rect 2745 1004 2775 1404
rect 3147 1004 3177 1404
rect 3235 1004 3265 1404
rect 3323 1004 3353 1404
rect 3411 1004 3441 1404
rect 3813 1004 3843 1404
rect 3901 1004 3931 1404
rect 3989 1004 4019 1404
rect 4077 1004 4107 1404
<< ndiff >>
rect 91 335 147 351
rect 91 301 101 335
rect 135 301 147 335
rect 91 263 147 301
rect 177 335 447 351
rect 177 306 198 335
tri 177 290 193 306 ne
rect 193 301 198 306
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 447 335
rect 193 290 447 301
rect 477 335 533 351
rect 477 301 489 335
rect 523 301 533 335
rect 91 229 101 263
rect 135 229 147 263
tri 253 260 283 290 ne
rect 283 263 342 290
rect 91 195 147 229
rect 91 161 101 195
rect 135 161 147 195
rect 91 129 147 161
tri 177 244 193 260 se
rect 193 244 237 260
tri 237 244 253 260 sw
rect 177 210 253 244
rect 177 176 198 210
rect 232 176 253 210
rect 177 175 253 176
tri 177 159 193 175 ne
rect 193 159 237 175
tri 237 159 253 175 nw
rect 283 229 295 263
rect 329 229 342 263
tri 342 260 372 290 nw
rect 283 195 342 229
rect 283 161 295 195
rect 329 161 342 195
tri 372 244 388 260 se
rect 388 244 431 260
tri 431 244 447 260 sw
rect 372 216 447 244
rect 372 182 393 216
rect 427 182 447 216
tri 372 166 388 182 ne
rect 388 166 431 182
tri 431 166 447 182 nw
tri 147 129 177 159 sw
tri 253 129 283 159 se
rect 283 136 342 161
tri 342 136 372 166 sw
tri 447 136 477 166 se
rect 477 136 533 301
rect 283 129 533 136
rect 91 125 533 129
rect 91 91 101 125
rect 135 91 295 125
rect 329 91 392 125
rect 426 91 489 125
rect 523 91 533 125
rect 91 75 533 91
rect 593 335 649 351
rect 593 301 603 335
rect 637 301 649 335
rect 593 263 649 301
rect 679 314 841 351
tri 679 298 695 314 ne
rect 695 298 841 314
tri 755 268 785 298 ne
rect 593 229 603 263
rect 637 229 649 263
rect 593 195 649 229
rect 593 161 603 195
rect 637 161 649 195
tri 679 252 695 268 se
rect 695 252 739 268
tri 739 252 755 268 sw
rect 679 219 755 252
rect 679 185 700 219
rect 734 185 755 219
rect 679 183 755 185
tri 679 167 695 183 ne
rect 695 167 739 183
tri 739 167 755 183 nw
rect 785 263 841 298
rect 785 229 797 263
rect 831 229 841 263
rect 785 195 841 229
rect 593 137 649 161
tri 649 137 679 167 sw
tri 755 137 785 167 se
rect 785 161 797 195
rect 831 161 841 195
rect 785 137 841 161
rect 593 125 841 137
rect 593 91 603 125
rect 637 91 700 125
rect 734 91 797 125
rect 831 91 841 125
rect 593 75 841 91
rect 1074 333 1130 349
rect 1074 299 1084 333
rect 1118 299 1130 333
rect 1074 261 1130 299
rect 1160 333 1324 349
rect 1160 304 1181 333
tri 1160 288 1176 304 ne
rect 1176 299 1181 304
rect 1215 299 1278 333
rect 1312 299 1324 333
rect 1176 288 1324 299
rect 1354 312 1516 349
tri 1354 296 1370 312 ne
rect 1370 296 1516 312
rect 1074 227 1084 261
rect 1118 227 1130 261
tri 1236 258 1266 288 ne
rect 1266 261 1324 288
tri 1430 266 1460 296 ne
rect 1074 193 1130 227
rect 1074 159 1084 193
rect 1118 159 1130 193
rect 1074 127 1130 159
tri 1160 242 1176 258 se
rect 1176 242 1220 258
tri 1220 242 1236 258 sw
rect 1160 208 1236 242
rect 1160 174 1181 208
rect 1215 174 1236 208
rect 1160 173 1236 174
tri 1160 157 1176 173 ne
rect 1176 157 1220 173
tri 1220 157 1236 173 nw
rect 1266 227 1278 261
rect 1312 227 1324 261
rect 1266 193 1324 227
rect 1266 159 1278 193
rect 1312 159 1324 193
tri 1354 250 1370 266 se
rect 1370 250 1414 266
tri 1414 250 1430 266 sw
rect 1354 217 1430 250
rect 1354 183 1375 217
rect 1409 183 1430 217
rect 1354 181 1430 183
tri 1354 165 1370 181 ne
rect 1370 165 1414 181
tri 1414 165 1430 181 nw
rect 1460 261 1516 296
rect 1460 227 1472 261
rect 1506 227 1516 261
rect 1460 193 1516 227
tri 1130 127 1160 157 sw
tri 1236 127 1266 157 se
rect 1266 135 1324 159
tri 1324 135 1354 165 sw
tri 1430 135 1460 165 se
rect 1460 159 1472 193
rect 1506 159 1516 193
rect 1460 135 1516 159
rect 1266 127 1516 135
rect 1074 123 1516 127
rect 1074 89 1084 123
rect 1118 89 1278 123
rect 1312 89 1375 123
rect 1409 89 1472 123
rect 1506 89 1516 123
rect 1074 73 1516 89
rect 1740 333 1796 349
rect 1740 299 1750 333
rect 1784 299 1796 333
rect 1740 261 1796 299
rect 1826 333 1990 349
rect 1826 304 1847 333
tri 1826 288 1842 304 ne
rect 1842 299 1847 304
rect 1881 299 1944 333
rect 1978 299 1990 333
rect 1842 288 1990 299
rect 2020 312 2182 349
tri 2020 296 2036 312 ne
rect 2036 296 2182 312
rect 1740 227 1750 261
rect 1784 227 1796 261
tri 1902 258 1932 288 ne
rect 1932 261 1990 288
tri 2096 266 2126 296 ne
rect 1740 193 1796 227
rect 1740 159 1750 193
rect 1784 159 1796 193
rect 1740 127 1796 159
tri 1826 242 1842 258 se
rect 1842 242 1886 258
tri 1886 242 1902 258 sw
rect 1826 208 1902 242
rect 1826 174 1847 208
rect 1881 174 1902 208
rect 1826 173 1902 174
tri 1826 157 1842 173 ne
rect 1842 157 1886 173
tri 1886 157 1902 173 nw
rect 1932 227 1944 261
rect 1978 227 1990 261
rect 1932 193 1990 227
rect 1932 159 1944 193
rect 1978 159 1990 193
tri 2020 250 2036 266 se
rect 2036 250 2080 266
tri 2080 250 2096 266 sw
rect 2020 217 2096 250
rect 2020 183 2041 217
rect 2075 183 2096 217
rect 2020 181 2096 183
tri 2020 165 2036 181 ne
rect 2036 165 2080 181
tri 2080 165 2096 181 nw
rect 2126 261 2182 296
rect 2126 227 2138 261
rect 2172 227 2182 261
rect 2126 193 2182 227
tri 1796 127 1826 157 sw
tri 1902 127 1932 157 se
rect 1932 135 1990 159
tri 1990 135 2020 165 sw
tri 2096 135 2126 165 se
rect 2126 159 2138 193
rect 2172 159 2182 193
rect 2126 135 2182 159
rect 1932 127 2182 135
rect 1740 123 2182 127
rect 1740 89 1750 123
rect 1784 89 1944 123
rect 1978 89 2041 123
rect 2075 89 2138 123
rect 2172 89 2182 123
rect 1740 73 2182 89
rect 2406 333 2462 349
rect 2406 299 2416 333
rect 2450 299 2462 333
rect 2406 261 2462 299
rect 2492 333 2656 349
rect 2492 304 2513 333
tri 2492 288 2508 304 ne
rect 2508 299 2513 304
rect 2547 299 2610 333
rect 2644 299 2656 333
rect 2508 288 2656 299
rect 2686 312 2848 349
tri 2686 296 2702 312 ne
rect 2702 296 2848 312
rect 2406 227 2416 261
rect 2450 227 2462 261
tri 2568 258 2598 288 ne
rect 2598 261 2656 288
tri 2762 266 2792 296 ne
rect 2406 193 2462 227
rect 2406 159 2416 193
rect 2450 159 2462 193
rect 2406 127 2462 159
tri 2492 242 2508 258 se
rect 2508 242 2552 258
tri 2552 242 2568 258 sw
rect 2492 208 2568 242
rect 2492 174 2513 208
rect 2547 174 2568 208
rect 2492 173 2568 174
tri 2492 157 2508 173 ne
rect 2508 157 2552 173
tri 2552 157 2568 173 nw
rect 2598 227 2610 261
rect 2644 227 2656 261
rect 2598 193 2656 227
rect 2598 159 2610 193
rect 2644 159 2656 193
tri 2686 250 2702 266 se
rect 2702 250 2746 266
tri 2746 250 2762 266 sw
rect 2686 217 2762 250
rect 2686 183 2707 217
rect 2741 183 2762 217
rect 2686 181 2762 183
tri 2686 165 2702 181 ne
rect 2702 165 2746 181
tri 2746 165 2762 181 nw
rect 2792 261 2848 296
rect 2792 227 2804 261
rect 2838 227 2848 261
rect 2792 193 2848 227
tri 2462 127 2492 157 sw
tri 2568 127 2598 157 se
rect 2598 135 2656 159
tri 2656 135 2686 165 sw
tri 2762 135 2792 165 se
rect 2792 159 2804 193
rect 2838 159 2848 193
rect 2792 135 2848 159
rect 2598 127 2848 135
rect 2406 123 2848 127
rect 2406 89 2416 123
rect 2450 89 2610 123
rect 2644 89 2707 123
rect 2741 89 2804 123
rect 2838 89 2848 123
rect 2406 73 2848 89
rect 3072 333 3128 349
rect 3072 299 3082 333
rect 3116 299 3128 333
rect 3072 261 3128 299
rect 3158 333 3322 349
rect 3158 304 3179 333
tri 3158 288 3174 304 ne
rect 3174 299 3179 304
rect 3213 299 3276 333
rect 3310 299 3322 333
rect 3174 288 3322 299
rect 3352 312 3514 349
tri 3352 296 3368 312 ne
rect 3368 296 3514 312
rect 3072 227 3082 261
rect 3116 227 3128 261
tri 3234 258 3264 288 ne
rect 3264 261 3322 288
tri 3428 266 3458 296 ne
rect 3072 193 3128 227
rect 3072 159 3082 193
rect 3116 159 3128 193
rect 3072 127 3128 159
tri 3158 242 3174 258 se
rect 3174 242 3218 258
tri 3218 242 3234 258 sw
rect 3158 208 3234 242
rect 3158 174 3179 208
rect 3213 174 3234 208
rect 3158 173 3234 174
tri 3158 157 3174 173 ne
rect 3174 157 3218 173
tri 3218 157 3234 173 nw
rect 3264 227 3276 261
rect 3310 227 3322 261
rect 3264 193 3322 227
rect 3264 159 3276 193
rect 3310 159 3322 193
tri 3352 250 3368 266 se
rect 3368 250 3412 266
tri 3412 250 3428 266 sw
rect 3352 217 3428 250
rect 3352 183 3373 217
rect 3407 183 3428 217
rect 3352 181 3428 183
tri 3352 165 3368 181 ne
rect 3368 165 3412 181
tri 3412 165 3428 181 nw
rect 3458 261 3514 296
rect 3458 227 3470 261
rect 3504 227 3514 261
rect 3458 193 3514 227
tri 3128 127 3158 157 sw
tri 3234 127 3264 157 se
rect 3264 135 3322 159
tri 3322 135 3352 165 sw
tri 3428 135 3458 165 se
rect 3458 159 3470 193
rect 3504 159 3514 193
rect 3458 135 3514 159
rect 3264 127 3514 135
rect 3072 123 3514 127
rect 3072 89 3082 123
rect 3116 89 3276 123
rect 3310 89 3373 123
rect 3407 89 3470 123
rect 3504 89 3514 123
rect 3072 73 3514 89
rect 3738 333 3794 349
rect 3738 299 3748 333
rect 3782 299 3794 333
rect 3738 261 3794 299
rect 3824 333 3988 349
rect 3824 304 3845 333
tri 3824 288 3840 304 ne
rect 3840 299 3845 304
rect 3879 299 3942 333
rect 3976 299 3988 333
rect 3840 288 3988 299
rect 4018 312 4180 349
tri 4018 296 4034 312 ne
rect 4034 296 4180 312
rect 3738 227 3748 261
rect 3782 227 3794 261
tri 3900 258 3930 288 ne
rect 3930 261 3988 288
tri 4094 266 4124 296 ne
rect 3738 193 3794 227
rect 3738 159 3748 193
rect 3782 159 3794 193
rect 3738 127 3794 159
tri 3824 242 3840 258 se
rect 3840 242 3884 258
tri 3884 242 3900 258 sw
rect 3824 208 3900 242
rect 3824 174 3845 208
rect 3879 174 3900 208
rect 3824 173 3900 174
tri 3824 157 3840 173 ne
rect 3840 157 3884 173
tri 3884 157 3900 173 nw
rect 3930 227 3942 261
rect 3976 227 3988 261
rect 3930 193 3988 227
rect 3930 159 3942 193
rect 3976 159 3988 193
tri 4018 250 4034 266 se
rect 4034 250 4078 266
tri 4078 250 4094 266 sw
rect 4018 217 4094 250
rect 4018 183 4039 217
rect 4073 183 4094 217
rect 4018 181 4094 183
tri 4018 165 4034 181 ne
rect 4034 165 4078 181
tri 4078 165 4094 181 nw
rect 4124 261 4180 296
rect 4124 227 4136 261
rect 4170 227 4180 261
rect 4124 193 4180 227
tri 3794 127 3824 157 sw
tri 3900 127 3930 157 se
rect 3930 135 3988 159
tri 3988 135 4018 165 sw
tri 4094 135 4124 165 se
rect 4124 159 4136 193
rect 4170 159 4180 193
rect 4124 135 4180 159
rect 3930 127 4180 135
rect 3738 123 4180 127
rect 3738 89 3748 123
rect 3782 89 3942 123
rect 3976 89 4039 123
rect 4073 89 4136 123
rect 4170 89 4180 123
rect 3738 73 4180 89
<< pdiff >>
rect 191 1366 247 1404
rect 191 1332 201 1366
rect 235 1332 247 1366
rect 191 1298 247 1332
rect 191 1264 201 1298
rect 235 1264 247 1298
rect 191 1230 247 1264
rect 191 1196 201 1230
rect 235 1196 247 1230
rect 191 1162 247 1196
rect 191 1128 201 1162
rect 235 1128 247 1162
rect 191 1093 247 1128
rect 191 1059 201 1093
rect 235 1059 247 1093
rect 191 1004 247 1059
rect 277 1366 335 1404
rect 277 1332 289 1366
rect 323 1332 335 1366
rect 277 1298 335 1332
rect 277 1264 289 1298
rect 323 1264 335 1298
rect 277 1230 335 1264
rect 277 1196 289 1230
rect 323 1196 335 1230
rect 277 1162 335 1196
rect 277 1128 289 1162
rect 323 1128 335 1162
rect 277 1093 335 1128
rect 277 1059 289 1093
rect 323 1059 335 1093
rect 277 1004 335 1059
rect 365 1366 423 1404
rect 365 1332 377 1366
rect 411 1332 423 1366
rect 365 1298 423 1332
rect 365 1264 377 1298
rect 411 1264 423 1298
rect 365 1230 423 1264
rect 365 1196 377 1230
rect 411 1196 423 1230
rect 365 1162 423 1196
rect 365 1128 377 1162
rect 411 1128 423 1162
rect 365 1004 423 1128
rect 453 1366 511 1404
rect 453 1332 465 1366
rect 499 1332 511 1366
rect 453 1298 511 1332
rect 453 1264 465 1298
rect 499 1264 511 1298
rect 453 1230 511 1264
rect 453 1196 465 1230
rect 499 1196 511 1230
rect 453 1162 511 1196
rect 453 1128 465 1162
rect 499 1128 511 1162
rect 453 1093 511 1128
rect 453 1059 465 1093
rect 499 1059 511 1093
rect 453 1004 511 1059
rect 541 1366 599 1404
rect 541 1332 553 1366
rect 587 1332 599 1366
rect 541 1298 599 1332
rect 541 1264 553 1298
rect 587 1264 599 1298
rect 541 1230 599 1264
rect 541 1196 553 1230
rect 587 1196 599 1230
rect 541 1162 599 1196
rect 541 1128 553 1162
rect 587 1128 599 1162
rect 541 1004 599 1128
rect 629 1366 687 1404
rect 629 1332 641 1366
rect 675 1332 687 1366
rect 629 1298 687 1332
rect 629 1264 641 1298
rect 675 1264 687 1298
rect 629 1230 687 1264
rect 629 1196 641 1230
rect 675 1196 687 1230
rect 629 1162 687 1196
rect 629 1128 641 1162
rect 675 1128 687 1162
rect 629 1093 687 1128
rect 629 1059 641 1093
rect 675 1059 687 1093
rect 629 1004 687 1059
rect 717 1366 771 1404
rect 717 1332 729 1366
rect 763 1332 771 1366
rect 717 1298 771 1332
rect 717 1264 729 1298
rect 763 1264 771 1298
rect 717 1230 771 1264
rect 717 1196 729 1230
rect 763 1196 771 1230
rect 717 1162 771 1196
rect 717 1128 729 1162
rect 763 1128 771 1162
rect 717 1004 771 1128
rect 1093 1366 1149 1404
rect 1093 1332 1103 1366
rect 1137 1332 1149 1366
rect 1093 1298 1149 1332
rect 1093 1264 1103 1298
rect 1137 1264 1149 1298
rect 1093 1230 1149 1264
rect 1093 1196 1103 1230
rect 1137 1196 1149 1230
rect 1093 1162 1149 1196
rect 1093 1128 1103 1162
rect 1137 1128 1149 1162
rect 1093 1093 1149 1128
rect 1093 1059 1103 1093
rect 1137 1059 1149 1093
rect 1093 1004 1149 1059
rect 1179 1366 1237 1404
rect 1179 1332 1191 1366
rect 1225 1332 1237 1366
rect 1179 1298 1237 1332
rect 1179 1264 1191 1298
rect 1225 1264 1237 1298
rect 1179 1230 1237 1264
rect 1179 1196 1191 1230
rect 1225 1196 1237 1230
rect 1179 1162 1237 1196
rect 1179 1128 1191 1162
rect 1225 1128 1237 1162
rect 1179 1093 1237 1128
rect 1179 1059 1191 1093
rect 1225 1059 1237 1093
rect 1179 1004 1237 1059
rect 1267 1366 1325 1404
rect 1267 1332 1279 1366
rect 1313 1332 1325 1366
rect 1267 1298 1325 1332
rect 1267 1264 1279 1298
rect 1313 1264 1325 1298
rect 1267 1230 1325 1264
rect 1267 1196 1279 1230
rect 1313 1196 1325 1230
rect 1267 1162 1325 1196
rect 1267 1128 1279 1162
rect 1313 1128 1325 1162
rect 1267 1004 1325 1128
rect 1355 1366 1413 1404
rect 1355 1332 1367 1366
rect 1401 1332 1413 1366
rect 1355 1298 1413 1332
rect 1355 1264 1367 1298
rect 1401 1264 1413 1298
rect 1355 1230 1413 1264
rect 1355 1196 1367 1230
rect 1401 1196 1413 1230
rect 1355 1162 1413 1196
rect 1355 1128 1367 1162
rect 1401 1128 1413 1162
rect 1355 1093 1413 1128
rect 1355 1059 1367 1093
rect 1401 1059 1413 1093
rect 1355 1004 1413 1059
rect 1443 1366 1497 1404
rect 1443 1332 1455 1366
rect 1489 1332 1497 1366
rect 1443 1298 1497 1332
rect 1443 1264 1455 1298
rect 1489 1264 1497 1298
rect 1443 1230 1497 1264
rect 1443 1196 1455 1230
rect 1489 1196 1497 1230
rect 1443 1162 1497 1196
rect 1443 1128 1455 1162
rect 1489 1128 1497 1162
rect 1443 1004 1497 1128
rect 1759 1366 1815 1404
rect 1759 1332 1769 1366
rect 1803 1332 1815 1366
rect 1759 1298 1815 1332
rect 1759 1264 1769 1298
rect 1803 1264 1815 1298
rect 1759 1230 1815 1264
rect 1759 1196 1769 1230
rect 1803 1196 1815 1230
rect 1759 1162 1815 1196
rect 1759 1128 1769 1162
rect 1803 1128 1815 1162
rect 1759 1093 1815 1128
rect 1759 1059 1769 1093
rect 1803 1059 1815 1093
rect 1759 1004 1815 1059
rect 1845 1366 1903 1404
rect 1845 1332 1857 1366
rect 1891 1332 1903 1366
rect 1845 1298 1903 1332
rect 1845 1264 1857 1298
rect 1891 1264 1903 1298
rect 1845 1230 1903 1264
rect 1845 1196 1857 1230
rect 1891 1196 1903 1230
rect 1845 1162 1903 1196
rect 1845 1128 1857 1162
rect 1891 1128 1903 1162
rect 1845 1093 1903 1128
rect 1845 1059 1857 1093
rect 1891 1059 1903 1093
rect 1845 1004 1903 1059
rect 1933 1366 1991 1404
rect 1933 1332 1945 1366
rect 1979 1332 1991 1366
rect 1933 1298 1991 1332
rect 1933 1264 1945 1298
rect 1979 1264 1991 1298
rect 1933 1230 1991 1264
rect 1933 1196 1945 1230
rect 1979 1196 1991 1230
rect 1933 1162 1991 1196
rect 1933 1128 1945 1162
rect 1979 1128 1991 1162
rect 1933 1004 1991 1128
rect 2021 1366 2079 1404
rect 2021 1332 2033 1366
rect 2067 1332 2079 1366
rect 2021 1298 2079 1332
rect 2021 1264 2033 1298
rect 2067 1264 2079 1298
rect 2021 1230 2079 1264
rect 2021 1196 2033 1230
rect 2067 1196 2079 1230
rect 2021 1162 2079 1196
rect 2021 1128 2033 1162
rect 2067 1128 2079 1162
rect 2021 1093 2079 1128
rect 2021 1059 2033 1093
rect 2067 1059 2079 1093
rect 2021 1004 2079 1059
rect 2109 1366 2163 1404
rect 2109 1332 2121 1366
rect 2155 1332 2163 1366
rect 2109 1298 2163 1332
rect 2109 1264 2121 1298
rect 2155 1264 2163 1298
rect 2109 1230 2163 1264
rect 2109 1196 2121 1230
rect 2155 1196 2163 1230
rect 2109 1162 2163 1196
rect 2109 1128 2121 1162
rect 2155 1128 2163 1162
rect 2109 1004 2163 1128
rect 2425 1366 2481 1404
rect 2425 1332 2435 1366
rect 2469 1332 2481 1366
rect 2425 1298 2481 1332
rect 2425 1264 2435 1298
rect 2469 1264 2481 1298
rect 2425 1230 2481 1264
rect 2425 1196 2435 1230
rect 2469 1196 2481 1230
rect 2425 1162 2481 1196
rect 2425 1128 2435 1162
rect 2469 1128 2481 1162
rect 2425 1093 2481 1128
rect 2425 1059 2435 1093
rect 2469 1059 2481 1093
rect 2425 1004 2481 1059
rect 2511 1366 2569 1404
rect 2511 1332 2523 1366
rect 2557 1332 2569 1366
rect 2511 1298 2569 1332
rect 2511 1264 2523 1298
rect 2557 1264 2569 1298
rect 2511 1230 2569 1264
rect 2511 1196 2523 1230
rect 2557 1196 2569 1230
rect 2511 1162 2569 1196
rect 2511 1128 2523 1162
rect 2557 1128 2569 1162
rect 2511 1093 2569 1128
rect 2511 1059 2523 1093
rect 2557 1059 2569 1093
rect 2511 1004 2569 1059
rect 2599 1366 2657 1404
rect 2599 1332 2611 1366
rect 2645 1332 2657 1366
rect 2599 1298 2657 1332
rect 2599 1264 2611 1298
rect 2645 1264 2657 1298
rect 2599 1230 2657 1264
rect 2599 1196 2611 1230
rect 2645 1196 2657 1230
rect 2599 1162 2657 1196
rect 2599 1128 2611 1162
rect 2645 1128 2657 1162
rect 2599 1004 2657 1128
rect 2687 1366 2745 1404
rect 2687 1332 2699 1366
rect 2733 1332 2745 1366
rect 2687 1298 2745 1332
rect 2687 1264 2699 1298
rect 2733 1264 2745 1298
rect 2687 1230 2745 1264
rect 2687 1196 2699 1230
rect 2733 1196 2745 1230
rect 2687 1162 2745 1196
rect 2687 1128 2699 1162
rect 2733 1128 2745 1162
rect 2687 1093 2745 1128
rect 2687 1059 2699 1093
rect 2733 1059 2745 1093
rect 2687 1004 2745 1059
rect 2775 1366 2829 1404
rect 2775 1332 2787 1366
rect 2821 1332 2829 1366
rect 2775 1298 2829 1332
rect 2775 1264 2787 1298
rect 2821 1264 2829 1298
rect 2775 1230 2829 1264
rect 2775 1196 2787 1230
rect 2821 1196 2829 1230
rect 2775 1162 2829 1196
rect 2775 1128 2787 1162
rect 2821 1128 2829 1162
rect 2775 1004 2829 1128
rect 3091 1366 3147 1404
rect 3091 1332 3101 1366
rect 3135 1332 3147 1366
rect 3091 1298 3147 1332
rect 3091 1264 3101 1298
rect 3135 1264 3147 1298
rect 3091 1230 3147 1264
rect 3091 1196 3101 1230
rect 3135 1196 3147 1230
rect 3091 1162 3147 1196
rect 3091 1128 3101 1162
rect 3135 1128 3147 1162
rect 3091 1093 3147 1128
rect 3091 1059 3101 1093
rect 3135 1059 3147 1093
rect 3091 1004 3147 1059
rect 3177 1366 3235 1404
rect 3177 1332 3189 1366
rect 3223 1332 3235 1366
rect 3177 1298 3235 1332
rect 3177 1264 3189 1298
rect 3223 1264 3235 1298
rect 3177 1230 3235 1264
rect 3177 1196 3189 1230
rect 3223 1196 3235 1230
rect 3177 1162 3235 1196
rect 3177 1128 3189 1162
rect 3223 1128 3235 1162
rect 3177 1093 3235 1128
rect 3177 1059 3189 1093
rect 3223 1059 3235 1093
rect 3177 1004 3235 1059
rect 3265 1366 3323 1404
rect 3265 1332 3277 1366
rect 3311 1332 3323 1366
rect 3265 1298 3323 1332
rect 3265 1264 3277 1298
rect 3311 1264 3323 1298
rect 3265 1230 3323 1264
rect 3265 1196 3277 1230
rect 3311 1196 3323 1230
rect 3265 1162 3323 1196
rect 3265 1128 3277 1162
rect 3311 1128 3323 1162
rect 3265 1004 3323 1128
rect 3353 1366 3411 1404
rect 3353 1332 3365 1366
rect 3399 1332 3411 1366
rect 3353 1298 3411 1332
rect 3353 1264 3365 1298
rect 3399 1264 3411 1298
rect 3353 1230 3411 1264
rect 3353 1196 3365 1230
rect 3399 1196 3411 1230
rect 3353 1162 3411 1196
rect 3353 1128 3365 1162
rect 3399 1128 3411 1162
rect 3353 1093 3411 1128
rect 3353 1059 3365 1093
rect 3399 1059 3411 1093
rect 3353 1004 3411 1059
rect 3441 1366 3495 1404
rect 3441 1332 3453 1366
rect 3487 1332 3495 1366
rect 3441 1298 3495 1332
rect 3441 1264 3453 1298
rect 3487 1264 3495 1298
rect 3441 1230 3495 1264
rect 3441 1196 3453 1230
rect 3487 1196 3495 1230
rect 3441 1162 3495 1196
rect 3441 1128 3453 1162
rect 3487 1128 3495 1162
rect 3441 1004 3495 1128
rect 3757 1366 3813 1404
rect 3757 1332 3767 1366
rect 3801 1332 3813 1366
rect 3757 1298 3813 1332
rect 3757 1264 3767 1298
rect 3801 1264 3813 1298
rect 3757 1230 3813 1264
rect 3757 1196 3767 1230
rect 3801 1196 3813 1230
rect 3757 1162 3813 1196
rect 3757 1128 3767 1162
rect 3801 1128 3813 1162
rect 3757 1093 3813 1128
rect 3757 1059 3767 1093
rect 3801 1059 3813 1093
rect 3757 1004 3813 1059
rect 3843 1366 3901 1404
rect 3843 1332 3855 1366
rect 3889 1332 3901 1366
rect 3843 1298 3901 1332
rect 3843 1264 3855 1298
rect 3889 1264 3901 1298
rect 3843 1230 3901 1264
rect 3843 1196 3855 1230
rect 3889 1196 3901 1230
rect 3843 1162 3901 1196
rect 3843 1128 3855 1162
rect 3889 1128 3901 1162
rect 3843 1093 3901 1128
rect 3843 1059 3855 1093
rect 3889 1059 3901 1093
rect 3843 1004 3901 1059
rect 3931 1366 3989 1404
rect 3931 1332 3943 1366
rect 3977 1332 3989 1366
rect 3931 1298 3989 1332
rect 3931 1264 3943 1298
rect 3977 1264 3989 1298
rect 3931 1230 3989 1264
rect 3931 1196 3943 1230
rect 3977 1196 3989 1230
rect 3931 1162 3989 1196
rect 3931 1128 3943 1162
rect 3977 1128 3989 1162
rect 3931 1004 3989 1128
rect 4019 1366 4077 1404
rect 4019 1332 4031 1366
rect 4065 1332 4077 1366
rect 4019 1298 4077 1332
rect 4019 1264 4031 1298
rect 4065 1264 4077 1298
rect 4019 1230 4077 1264
rect 4019 1196 4031 1230
rect 4065 1196 4077 1230
rect 4019 1162 4077 1196
rect 4019 1128 4031 1162
rect 4065 1128 4077 1162
rect 4019 1093 4077 1128
rect 4019 1059 4031 1093
rect 4065 1059 4077 1093
rect 4019 1004 4077 1059
rect 4107 1366 4161 1404
rect 4107 1332 4119 1366
rect 4153 1332 4161 1366
rect 4107 1298 4161 1332
rect 4107 1264 4119 1298
rect 4153 1264 4161 1298
rect 4107 1230 4161 1264
rect 4107 1196 4119 1230
rect 4153 1196 4161 1230
rect 4107 1162 4161 1196
rect 4107 1128 4119 1162
rect 4153 1128 4161 1162
rect 4107 1004 4161 1128
<< ndiffc >>
rect 101 301 135 335
rect 198 301 232 335
rect 295 301 329 335
rect 392 301 426 335
rect 489 301 523 335
rect 101 229 135 263
rect 101 161 135 195
rect 198 176 232 210
rect 295 229 329 263
rect 295 161 329 195
rect 393 182 427 216
rect 101 91 135 125
rect 295 91 329 125
rect 392 91 426 125
rect 489 91 523 125
rect 603 301 637 335
rect 603 229 637 263
rect 603 161 637 195
rect 700 185 734 219
rect 797 229 831 263
rect 797 161 831 195
rect 603 91 637 125
rect 700 91 734 125
rect 797 91 831 125
rect 1084 299 1118 333
rect 1181 299 1215 333
rect 1278 299 1312 333
rect 1084 227 1118 261
rect 1084 159 1118 193
rect 1181 174 1215 208
rect 1278 227 1312 261
rect 1278 159 1312 193
rect 1375 183 1409 217
rect 1472 227 1506 261
rect 1472 159 1506 193
rect 1084 89 1118 123
rect 1278 89 1312 123
rect 1375 89 1409 123
rect 1472 89 1506 123
rect 1750 299 1784 333
rect 1847 299 1881 333
rect 1944 299 1978 333
rect 1750 227 1784 261
rect 1750 159 1784 193
rect 1847 174 1881 208
rect 1944 227 1978 261
rect 1944 159 1978 193
rect 2041 183 2075 217
rect 2138 227 2172 261
rect 2138 159 2172 193
rect 1750 89 1784 123
rect 1944 89 1978 123
rect 2041 89 2075 123
rect 2138 89 2172 123
rect 2416 299 2450 333
rect 2513 299 2547 333
rect 2610 299 2644 333
rect 2416 227 2450 261
rect 2416 159 2450 193
rect 2513 174 2547 208
rect 2610 227 2644 261
rect 2610 159 2644 193
rect 2707 183 2741 217
rect 2804 227 2838 261
rect 2804 159 2838 193
rect 2416 89 2450 123
rect 2610 89 2644 123
rect 2707 89 2741 123
rect 2804 89 2838 123
rect 3082 299 3116 333
rect 3179 299 3213 333
rect 3276 299 3310 333
rect 3082 227 3116 261
rect 3082 159 3116 193
rect 3179 174 3213 208
rect 3276 227 3310 261
rect 3276 159 3310 193
rect 3373 183 3407 217
rect 3470 227 3504 261
rect 3470 159 3504 193
rect 3082 89 3116 123
rect 3276 89 3310 123
rect 3373 89 3407 123
rect 3470 89 3504 123
rect 3748 299 3782 333
rect 3845 299 3879 333
rect 3942 299 3976 333
rect 3748 227 3782 261
rect 3748 159 3782 193
rect 3845 174 3879 208
rect 3942 227 3976 261
rect 3942 159 3976 193
rect 4039 183 4073 217
rect 4136 227 4170 261
rect 4136 159 4170 193
rect 3748 89 3782 123
rect 3942 89 3976 123
rect 4039 89 4073 123
rect 4136 89 4170 123
<< pdiffc >>
rect 201 1332 235 1366
rect 201 1264 235 1298
rect 201 1196 235 1230
rect 201 1128 235 1162
rect 201 1059 235 1093
rect 289 1332 323 1366
rect 289 1264 323 1298
rect 289 1196 323 1230
rect 289 1128 323 1162
rect 289 1059 323 1093
rect 377 1332 411 1366
rect 377 1264 411 1298
rect 377 1196 411 1230
rect 377 1128 411 1162
rect 465 1332 499 1366
rect 465 1264 499 1298
rect 465 1196 499 1230
rect 465 1128 499 1162
rect 465 1059 499 1093
rect 553 1332 587 1366
rect 553 1264 587 1298
rect 553 1196 587 1230
rect 553 1128 587 1162
rect 641 1332 675 1366
rect 641 1264 675 1298
rect 641 1196 675 1230
rect 641 1128 675 1162
rect 641 1059 675 1093
rect 729 1332 763 1366
rect 729 1264 763 1298
rect 729 1196 763 1230
rect 729 1128 763 1162
rect 1103 1332 1137 1366
rect 1103 1264 1137 1298
rect 1103 1196 1137 1230
rect 1103 1128 1137 1162
rect 1103 1059 1137 1093
rect 1191 1332 1225 1366
rect 1191 1264 1225 1298
rect 1191 1196 1225 1230
rect 1191 1128 1225 1162
rect 1191 1059 1225 1093
rect 1279 1332 1313 1366
rect 1279 1264 1313 1298
rect 1279 1196 1313 1230
rect 1279 1128 1313 1162
rect 1367 1332 1401 1366
rect 1367 1264 1401 1298
rect 1367 1196 1401 1230
rect 1367 1128 1401 1162
rect 1367 1059 1401 1093
rect 1455 1332 1489 1366
rect 1455 1264 1489 1298
rect 1455 1196 1489 1230
rect 1455 1128 1489 1162
rect 1769 1332 1803 1366
rect 1769 1264 1803 1298
rect 1769 1196 1803 1230
rect 1769 1128 1803 1162
rect 1769 1059 1803 1093
rect 1857 1332 1891 1366
rect 1857 1264 1891 1298
rect 1857 1196 1891 1230
rect 1857 1128 1891 1162
rect 1857 1059 1891 1093
rect 1945 1332 1979 1366
rect 1945 1264 1979 1298
rect 1945 1196 1979 1230
rect 1945 1128 1979 1162
rect 2033 1332 2067 1366
rect 2033 1264 2067 1298
rect 2033 1196 2067 1230
rect 2033 1128 2067 1162
rect 2033 1059 2067 1093
rect 2121 1332 2155 1366
rect 2121 1264 2155 1298
rect 2121 1196 2155 1230
rect 2121 1128 2155 1162
rect 2435 1332 2469 1366
rect 2435 1264 2469 1298
rect 2435 1196 2469 1230
rect 2435 1128 2469 1162
rect 2435 1059 2469 1093
rect 2523 1332 2557 1366
rect 2523 1264 2557 1298
rect 2523 1196 2557 1230
rect 2523 1128 2557 1162
rect 2523 1059 2557 1093
rect 2611 1332 2645 1366
rect 2611 1264 2645 1298
rect 2611 1196 2645 1230
rect 2611 1128 2645 1162
rect 2699 1332 2733 1366
rect 2699 1264 2733 1298
rect 2699 1196 2733 1230
rect 2699 1128 2733 1162
rect 2699 1059 2733 1093
rect 2787 1332 2821 1366
rect 2787 1264 2821 1298
rect 2787 1196 2821 1230
rect 2787 1128 2821 1162
rect 3101 1332 3135 1366
rect 3101 1264 3135 1298
rect 3101 1196 3135 1230
rect 3101 1128 3135 1162
rect 3101 1059 3135 1093
rect 3189 1332 3223 1366
rect 3189 1264 3223 1298
rect 3189 1196 3223 1230
rect 3189 1128 3223 1162
rect 3189 1059 3223 1093
rect 3277 1332 3311 1366
rect 3277 1264 3311 1298
rect 3277 1196 3311 1230
rect 3277 1128 3311 1162
rect 3365 1332 3399 1366
rect 3365 1264 3399 1298
rect 3365 1196 3399 1230
rect 3365 1128 3399 1162
rect 3365 1059 3399 1093
rect 3453 1332 3487 1366
rect 3453 1264 3487 1298
rect 3453 1196 3487 1230
rect 3453 1128 3487 1162
rect 3767 1332 3801 1366
rect 3767 1264 3801 1298
rect 3767 1196 3801 1230
rect 3767 1128 3801 1162
rect 3767 1059 3801 1093
rect 3855 1332 3889 1366
rect 3855 1264 3889 1298
rect 3855 1196 3889 1230
rect 3855 1128 3889 1162
rect 3855 1059 3889 1093
rect 3943 1332 3977 1366
rect 3943 1264 3977 1298
rect 3943 1196 3977 1230
rect 3943 1128 3977 1162
rect 4031 1332 4065 1366
rect 4031 1264 4065 1298
rect 4031 1196 4065 1230
rect 4031 1128 4065 1162
rect 4031 1059 4065 1093
rect 4119 1332 4153 1366
rect 4119 1264 4153 1298
rect 4119 1196 4153 1230
rect 4119 1128 4153 1162
<< psubdiff >>
rect -34 482 4326 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 928 461 996 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 928 427 945 461
rect 979 427 996 461
rect 1594 461 1662 482
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 928 313 996 353
rect 1594 427 1611 461
rect 1645 427 1662 461
rect 2260 461 2328 482
rect 1594 387 1662 427
rect 1594 353 1611 387
rect 1645 353 1662 387
rect 928 279 945 313
rect 979 279 996 313
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect -34 17 34 57
rect 928 57 945 91
rect 979 57 996 91
rect 1594 313 1662 353
rect 2260 427 2277 461
rect 2311 427 2328 461
rect 2926 461 2994 482
rect 2260 387 2328 427
rect 2260 353 2277 387
rect 2311 353 2328 387
rect 1594 279 1611 313
rect 1645 279 1662 313
rect 1594 239 1662 279
rect 1594 205 1611 239
rect 1645 205 1662 239
rect 1594 165 1662 205
rect 1594 131 1611 165
rect 1645 131 1662 165
rect 1594 91 1662 131
rect 928 17 996 57
rect 1594 57 1611 91
rect 1645 57 1662 91
rect 2260 313 2328 353
rect 2926 427 2943 461
rect 2977 427 2994 461
rect 3592 461 3660 482
rect 2926 387 2994 427
rect 2926 353 2943 387
rect 2977 353 2994 387
rect 2260 279 2277 313
rect 2311 279 2328 313
rect 2260 239 2328 279
rect 2260 205 2277 239
rect 2311 205 2328 239
rect 2260 165 2328 205
rect 2260 131 2277 165
rect 2311 131 2328 165
rect 2260 91 2328 131
rect 1594 17 1662 57
rect 2260 57 2277 91
rect 2311 57 2328 91
rect 2926 313 2994 353
rect 3592 427 3609 461
rect 3643 427 3660 461
rect 4258 461 4326 482
rect 3592 387 3660 427
rect 3592 353 3609 387
rect 3643 353 3660 387
rect 2926 279 2943 313
rect 2977 279 2994 313
rect 2926 239 2994 279
rect 2926 205 2943 239
rect 2977 205 2994 239
rect 2926 165 2994 205
rect 2926 131 2943 165
rect 2977 131 2994 165
rect 2926 91 2994 131
rect 2260 17 2328 57
rect 2926 57 2943 91
rect 2977 57 2994 91
rect 3592 313 3660 353
rect 4258 427 4275 461
rect 4309 427 4326 461
rect 4258 387 4326 427
rect 4258 353 4275 387
rect 4309 353 4326 387
rect 3592 279 3609 313
rect 3643 279 3660 313
rect 3592 239 3660 279
rect 3592 205 3609 239
rect 3643 205 3660 239
rect 3592 165 3660 205
rect 3592 131 3609 165
rect 3643 131 3660 165
rect 3592 91 3660 131
rect 2926 17 2994 57
rect 3592 57 3609 91
rect 3643 57 3660 91
rect 4258 313 4326 353
rect 4258 279 4275 313
rect 4309 279 4326 313
rect 4258 239 4326 279
rect 4258 205 4275 239
rect 4309 205 4326 239
rect 4258 165 4326 205
rect 4258 131 4275 165
rect 4309 131 4326 165
rect 4258 91 4326 131
rect 3592 17 3660 57
rect 4258 57 4275 91
rect 4309 57 4326 91
rect 4258 17 4326 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4326 17
rect -34 -34 4326 -17
<< nsubdiff >>
rect -34 1497 4326 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4326 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 928 1423 996 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 1594 1423 1662 1463
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect 928 1019 945 1053
rect 979 1019 996 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 928 979 996 1019
rect 1594 1389 1611 1423
rect 1645 1389 1662 1423
rect 2260 1423 2328 1463
rect 1594 1349 1662 1389
rect 1594 1315 1611 1349
rect 1645 1315 1662 1349
rect 1594 1275 1662 1315
rect 1594 1241 1611 1275
rect 1645 1241 1662 1275
rect 1594 1201 1662 1241
rect 1594 1167 1611 1201
rect 1645 1167 1662 1201
rect 1594 1127 1662 1167
rect 1594 1093 1611 1127
rect 1645 1093 1662 1127
rect 1594 1053 1662 1093
rect 1594 1019 1611 1053
rect 1645 1019 1662 1053
rect 928 945 945 979
rect 979 945 996 979
rect -34 871 -17 905
rect 17 884 34 905
rect 928 905 996 945
rect 1594 979 1662 1019
rect 2260 1389 2277 1423
rect 2311 1389 2328 1423
rect 2926 1423 2994 1463
rect 2260 1349 2328 1389
rect 2260 1315 2277 1349
rect 2311 1315 2328 1349
rect 2260 1275 2328 1315
rect 2260 1241 2277 1275
rect 2311 1241 2328 1275
rect 2260 1201 2328 1241
rect 2260 1167 2277 1201
rect 2311 1167 2328 1201
rect 2260 1127 2328 1167
rect 2260 1093 2277 1127
rect 2311 1093 2328 1127
rect 2260 1053 2328 1093
rect 2260 1019 2277 1053
rect 2311 1019 2328 1053
rect 1594 945 1611 979
rect 1645 945 1662 979
rect 928 884 945 905
rect 17 871 945 884
rect 979 884 996 905
rect 1594 905 1662 945
rect 2260 979 2328 1019
rect 2926 1389 2943 1423
rect 2977 1389 2994 1423
rect 3592 1423 3660 1463
rect 2926 1349 2994 1389
rect 2926 1315 2943 1349
rect 2977 1315 2994 1349
rect 2926 1275 2994 1315
rect 2926 1241 2943 1275
rect 2977 1241 2994 1275
rect 2926 1201 2994 1241
rect 2926 1167 2943 1201
rect 2977 1167 2994 1201
rect 2926 1127 2994 1167
rect 2926 1093 2943 1127
rect 2977 1093 2994 1127
rect 2926 1053 2994 1093
rect 2926 1019 2943 1053
rect 2977 1019 2994 1053
rect 2260 945 2277 979
rect 2311 945 2328 979
rect 1594 884 1611 905
rect 979 871 1611 884
rect 1645 884 1662 905
rect 2260 905 2328 945
rect 2926 979 2994 1019
rect 3592 1389 3609 1423
rect 3643 1389 3660 1423
rect 4258 1423 4326 1463
rect 3592 1349 3660 1389
rect 3592 1315 3609 1349
rect 3643 1315 3660 1349
rect 3592 1275 3660 1315
rect 3592 1241 3609 1275
rect 3643 1241 3660 1275
rect 3592 1201 3660 1241
rect 3592 1167 3609 1201
rect 3643 1167 3660 1201
rect 3592 1127 3660 1167
rect 3592 1093 3609 1127
rect 3643 1093 3660 1127
rect 3592 1053 3660 1093
rect 3592 1019 3609 1053
rect 3643 1019 3660 1053
rect 2926 945 2943 979
rect 2977 945 2994 979
rect 2260 884 2277 905
rect 1645 871 2277 884
rect 2311 884 2328 905
rect 2926 905 2994 945
rect 3592 979 3660 1019
rect 4258 1389 4275 1423
rect 4309 1389 4326 1423
rect 4258 1349 4326 1389
rect 4258 1315 4275 1349
rect 4309 1315 4326 1349
rect 4258 1275 4326 1315
rect 4258 1241 4275 1275
rect 4309 1241 4326 1275
rect 4258 1201 4326 1241
rect 4258 1167 4275 1201
rect 4309 1167 4326 1201
rect 4258 1127 4326 1167
rect 4258 1093 4275 1127
rect 4309 1093 4326 1127
rect 4258 1053 4326 1093
rect 4258 1019 4275 1053
rect 4309 1019 4326 1053
rect 3592 945 3609 979
rect 3643 945 3660 979
rect 2926 884 2943 905
rect 2311 871 2943 884
rect 2977 884 2994 905
rect 3592 905 3660 945
rect 4258 979 4326 1019
rect 4258 945 4275 979
rect 4309 945 4326 979
rect 3592 884 3609 905
rect 2977 871 3609 884
rect 3643 884 3660 905
rect 4258 905 4326 945
rect 4258 884 4275 905
rect 3643 871 4275 884
rect 4309 871 4326 905
rect -34 822 4326 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 945 427 979 461
rect 945 353 979 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1611 427 1645 461
rect 1611 353 1645 387
rect 945 279 979 313
rect 945 205 979 239
rect 945 131 979 165
rect 945 57 979 91
rect 2277 427 2311 461
rect 2277 353 2311 387
rect 1611 279 1645 313
rect 1611 205 1645 239
rect 1611 131 1645 165
rect 1611 57 1645 91
rect 2943 427 2977 461
rect 2943 353 2977 387
rect 2277 279 2311 313
rect 2277 205 2311 239
rect 2277 131 2311 165
rect 2277 57 2311 91
rect 3609 427 3643 461
rect 3609 353 3643 387
rect 2943 279 2977 313
rect 2943 205 2977 239
rect 2943 131 2977 165
rect 2943 57 2977 91
rect 4275 427 4309 461
rect 4275 353 4309 387
rect 3609 279 3643 313
rect 3609 205 3643 239
rect 3609 131 3643 165
rect 3609 57 3643 91
rect 4275 279 4309 313
rect 4275 205 4309 239
rect 4275 131 4309 165
rect 4275 57 4309 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 945 1389 979 1423
rect 945 1315 979 1349
rect 945 1241 979 1275
rect 945 1167 979 1201
rect 945 1093 979 1127
rect 945 1019 979 1053
rect -17 945 17 979
rect 1611 1389 1645 1423
rect 1611 1315 1645 1349
rect 1611 1241 1645 1275
rect 1611 1167 1645 1201
rect 1611 1093 1645 1127
rect 1611 1019 1645 1053
rect 945 945 979 979
rect -17 871 17 905
rect 2277 1389 2311 1423
rect 2277 1315 2311 1349
rect 2277 1241 2311 1275
rect 2277 1167 2311 1201
rect 2277 1093 2311 1127
rect 2277 1019 2311 1053
rect 1611 945 1645 979
rect 945 871 979 905
rect 2943 1389 2977 1423
rect 2943 1315 2977 1349
rect 2943 1241 2977 1275
rect 2943 1167 2977 1201
rect 2943 1093 2977 1127
rect 2943 1019 2977 1053
rect 2277 945 2311 979
rect 1611 871 1645 905
rect 3609 1389 3643 1423
rect 3609 1315 3643 1349
rect 3609 1241 3643 1275
rect 3609 1167 3643 1201
rect 3609 1093 3643 1127
rect 3609 1019 3643 1053
rect 2943 945 2977 979
rect 2277 871 2311 905
rect 4275 1389 4309 1423
rect 4275 1315 4309 1349
rect 4275 1241 4309 1275
rect 4275 1167 4309 1201
rect 4275 1093 4309 1127
rect 4275 1019 4309 1053
rect 3609 945 3643 979
rect 2943 871 2977 905
rect 4275 945 4309 979
rect 3609 871 3643 905
rect 4275 871 4309 905
<< poly >>
rect 247 1404 277 1430
rect 335 1404 365 1430
rect 423 1404 453 1430
rect 511 1404 541 1430
rect 599 1404 629 1430
rect 687 1404 717 1430
rect 1149 1404 1179 1430
rect 1237 1404 1267 1430
rect 1325 1404 1355 1430
rect 1413 1404 1443 1430
rect 247 973 277 1004
rect 335 973 365 1004
rect 423 973 453 1004
rect 511 973 541 1004
rect 195 957 365 973
rect 195 923 205 957
rect 239 943 365 957
rect 417 957 541 973
rect 239 923 249 943
rect 195 907 249 923
rect 417 923 427 957
rect 461 943 541 957
rect 599 973 629 1004
rect 687 973 717 1004
rect 599 957 717 973
rect 599 943 649 957
rect 461 923 471 943
rect 417 907 471 923
rect 639 923 649 943
rect 683 943 717 957
rect 1815 1404 1845 1430
rect 1903 1404 1933 1430
rect 1991 1404 2021 1430
rect 2079 1404 2109 1430
rect 683 923 693 943
rect 639 907 693 923
rect 1149 973 1179 1004
rect 1237 973 1267 1004
rect 1325 973 1355 1004
rect 1413 973 1443 1004
rect 1149 957 1267 973
rect 1149 943 1167 957
rect 1157 923 1167 943
rect 1201 943 1267 957
rect 1311 957 1443 973
rect 1201 923 1211 943
rect 1157 907 1211 923
rect 1311 923 1321 957
rect 1355 943 1443 957
rect 2481 1404 2511 1430
rect 2569 1404 2599 1430
rect 2657 1404 2687 1430
rect 2745 1404 2775 1430
rect 1355 923 1365 943
rect 1311 907 1365 923
rect 1815 973 1845 1004
rect 1903 973 1933 1004
rect 1991 973 2021 1004
rect 2079 973 2109 1004
rect 1815 957 1933 973
rect 1815 943 1833 957
rect 1823 923 1833 943
rect 1867 943 1933 957
rect 1977 957 2109 973
rect 1867 923 1877 943
rect 1823 907 1877 923
rect 1977 923 1987 957
rect 2021 943 2109 957
rect 3147 1404 3177 1430
rect 3235 1404 3265 1430
rect 3323 1404 3353 1430
rect 3411 1404 3441 1430
rect 2021 923 2031 943
rect 1977 907 2031 923
rect 2481 973 2511 1004
rect 2569 973 2599 1004
rect 2657 973 2687 1004
rect 2745 973 2775 1004
rect 2481 957 2599 973
rect 2481 943 2499 957
rect 2489 923 2499 943
rect 2533 943 2599 957
rect 2643 957 2775 973
rect 2533 923 2543 943
rect 2489 907 2543 923
rect 2643 923 2653 957
rect 2687 943 2775 957
rect 3813 1404 3843 1430
rect 3901 1404 3931 1430
rect 3989 1404 4019 1430
rect 4077 1404 4107 1430
rect 2687 923 2697 943
rect 2643 907 2697 923
rect 3147 973 3177 1004
rect 3235 973 3265 1004
rect 3323 973 3353 1004
rect 3411 973 3441 1004
rect 3147 957 3265 973
rect 3147 943 3165 957
rect 3155 923 3165 943
rect 3199 943 3265 957
rect 3309 957 3441 973
rect 3199 923 3209 943
rect 3155 907 3209 923
rect 3309 923 3319 957
rect 3353 943 3441 957
rect 3353 923 3363 943
rect 3309 907 3363 923
rect 3813 973 3843 1004
rect 3901 973 3931 1004
rect 3989 973 4019 1004
rect 4077 973 4107 1004
rect 3813 957 3931 973
rect 3813 943 3831 957
rect 3821 923 3831 943
rect 3865 943 3931 957
rect 3975 957 4107 973
rect 3865 923 3875 943
rect 3821 907 3875 923
rect 3975 923 3985 957
rect 4019 943 4107 957
rect 4019 923 4029 943
rect 3975 907 4029 923
rect 195 433 249 449
rect 195 413 205 433
rect 147 399 205 413
rect 239 399 249 433
rect 147 383 249 399
rect 417 433 471 449
rect 417 399 427 433
rect 461 413 471 433
rect 639 433 693 449
rect 461 399 477 413
rect 417 383 477 399
rect 639 399 649 433
rect 683 399 693 433
rect 639 383 693 399
rect 1157 433 1211 449
rect 1157 413 1167 433
rect 147 351 177 383
rect 447 351 477 383
rect 649 351 679 383
rect 1130 399 1167 413
rect 1201 399 1211 433
rect 1130 383 1211 399
rect 1305 433 1359 449
rect 1305 399 1315 433
rect 1349 399 1359 433
rect 1305 383 1359 399
rect 1823 433 1877 449
rect 1823 413 1833 433
rect 1130 349 1160 383
rect 1324 349 1354 383
rect 1796 399 1833 413
rect 1867 399 1877 433
rect 1796 383 1877 399
rect 1971 433 2025 449
rect 1971 399 1981 433
rect 2015 399 2025 433
rect 1971 383 2025 399
rect 2489 433 2543 449
rect 2489 413 2499 433
rect 1796 349 1826 383
rect 1990 349 2020 383
rect 2462 399 2499 413
rect 2533 399 2543 433
rect 2462 383 2543 399
rect 2637 433 2691 449
rect 2637 399 2647 433
rect 2681 399 2691 433
rect 2637 383 2691 399
rect 3155 433 3209 449
rect 3155 413 3165 433
rect 2462 349 2492 383
rect 2656 349 2686 383
rect 3128 399 3165 413
rect 3199 399 3209 433
rect 3128 383 3209 399
rect 3303 433 3357 449
rect 3303 399 3313 433
rect 3347 399 3357 433
rect 3303 383 3357 399
rect 3821 433 3875 449
rect 3821 413 3831 433
rect 3128 349 3158 383
rect 3322 349 3352 383
rect 3794 399 3831 413
rect 3865 399 3875 433
rect 3794 383 3875 399
rect 3969 433 4023 449
rect 3969 399 3979 433
rect 4013 399 4023 433
rect 3969 383 4023 399
rect 3794 349 3824 383
rect 3988 349 4018 383
<< polycont >>
rect 205 923 239 957
rect 427 923 461 957
rect 649 923 683 957
rect 1167 923 1201 957
rect 1321 923 1355 957
rect 1833 923 1867 957
rect 1987 923 2021 957
rect 2499 923 2533 957
rect 2653 923 2687 957
rect 3165 923 3199 957
rect 3319 923 3353 957
rect 3831 923 3865 957
rect 3985 923 4019 957
rect 205 399 239 433
rect 427 399 461 433
rect 649 399 683 433
rect 1167 399 1201 433
rect 1315 399 1349 433
rect 1833 399 1867 433
rect 1981 399 2015 433
rect 2499 399 2533 433
rect 2647 399 2681 433
rect 3165 399 3199 433
rect 3313 399 3347 433
rect 3831 399 3865 433
rect 3979 399 4013 433
<< locali >>
rect -34 1497 4326 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4326 1497
rect -34 1446 4326 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 201 1366 235 1446
rect 201 1298 235 1332
rect 201 1230 235 1264
rect 201 1162 235 1196
rect 201 1093 235 1128
rect 201 1043 235 1059
rect 289 1366 323 1404
rect 289 1298 323 1332
rect 289 1230 323 1264
rect 289 1162 323 1196
rect 289 1093 323 1128
rect 377 1366 411 1446
rect 377 1298 411 1332
rect 377 1230 411 1264
rect 377 1162 411 1196
rect 377 1111 411 1128
rect 465 1366 499 1404
rect 465 1298 499 1332
rect 465 1230 499 1264
rect 465 1162 499 1196
rect 289 1048 323 1059
rect 465 1093 499 1128
rect 553 1366 587 1446
rect 553 1298 587 1332
rect 553 1230 587 1264
rect 553 1162 587 1196
rect 553 1111 587 1128
rect 641 1366 675 1404
rect 641 1298 675 1332
rect 641 1230 675 1264
rect 641 1162 675 1196
rect 465 1048 499 1059
rect 641 1093 675 1128
rect 729 1366 763 1446
rect 729 1298 763 1332
rect 729 1230 763 1264
rect 729 1162 763 1196
rect 729 1111 763 1128
rect 928 1423 996 1446
rect 928 1389 945 1423
rect 979 1389 996 1423
rect 928 1349 996 1389
rect 928 1315 945 1349
rect 979 1315 996 1349
rect 928 1275 996 1315
rect 928 1241 945 1275
rect 979 1241 996 1275
rect 928 1201 996 1241
rect 928 1167 945 1201
rect 979 1167 996 1201
rect 928 1127 996 1167
rect 641 1048 675 1059
rect 928 1093 945 1127
rect 979 1093 996 1127
rect 928 1053 996 1093
rect -34 979 34 1019
rect 289 1014 831 1048
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect 205 831 239 923
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 797
rect 205 383 239 399
rect 427 957 461 973
rect 427 905 461 923
rect 427 433 461 871
rect 427 383 461 399
rect 649 957 683 973
rect 649 683 683 923
rect 649 433 683 649
rect 649 383 683 399
rect 797 757 831 1014
rect 928 1019 945 1053
rect 979 1019 996 1053
rect 1103 1366 1137 1446
rect 1103 1298 1137 1332
rect 1103 1230 1137 1264
rect 1103 1162 1137 1196
rect 1103 1093 1137 1128
rect 1103 1027 1137 1059
rect 1191 1366 1225 1404
rect 1191 1298 1225 1332
rect 1191 1230 1225 1264
rect 1191 1162 1225 1196
rect 1191 1093 1225 1128
rect 1279 1366 1313 1446
rect 1279 1298 1313 1332
rect 1279 1230 1313 1264
rect 1279 1162 1313 1196
rect 1279 1111 1313 1128
rect 1367 1366 1401 1404
rect 1367 1298 1401 1332
rect 1367 1230 1401 1264
rect 1367 1162 1401 1196
rect 1191 1057 1225 1059
rect 1367 1093 1401 1128
rect 1455 1366 1489 1446
rect 1455 1298 1489 1332
rect 1455 1230 1489 1264
rect 1455 1162 1489 1196
rect 1455 1111 1489 1128
rect 1594 1423 1662 1446
rect 1594 1389 1611 1423
rect 1645 1389 1662 1423
rect 1594 1349 1662 1389
rect 1594 1315 1611 1349
rect 1645 1315 1662 1349
rect 1594 1275 1662 1315
rect 1594 1241 1611 1275
rect 1645 1241 1662 1275
rect 1594 1201 1662 1241
rect 1594 1167 1611 1201
rect 1645 1167 1662 1201
rect 1594 1127 1662 1167
rect 1367 1057 1401 1059
rect 1594 1093 1611 1127
rect 1645 1093 1662 1127
rect 1191 1023 1497 1057
rect 928 979 996 1019
rect 928 945 945 979
rect 979 945 996 979
rect 928 905 996 945
rect 928 871 945 905
rect 979 871 996 905
rect 928 822 996 871
rect 1167 957 1201 973
rect 1321 957 1355 973
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 101 335 135 351
rect 295 335 329 351
rect 489 335 523 351
rect 135 301 198 335
rect 232 301 295 335
rect 329 301 392 335
rect 426 301 489 335
rect 101 263 135 301
rect 101 195 135 229
rect 295 263 329 301
rect 489 285 523 301
rect 603 335 637 351
rect 797 350 831 723
rect 1167 757 1201 923
rect 603 263 637 301
rect 101 125 135 161
rect 101 75 135 91
rect 198 210 232 226
rect -34 34 34 57
rect 198 34 232 176
rect 295 195 329 229
rect 393 216 427 232
rect 603 216 637 229
rect 427 195 637 216
rect 427 182 603 195
rect 393 166 427 182
rect 295 125 329 161
rect 700 316 831 350
rect 928 461 996 544
rect 928 427 945 461
rect 979 427 996 461
rect 928 387 996 427
rect 928 353 945 387
rect 979 353 996 387
rect 1167 433 1201 723
rect 1167 383 1201 399
rect 1315 923 1321 942
rect 1315 907 1355 923
rect 1315 433 1349 907
rect 1315 383 1349 399
rect 1463 683 1497 1023
rect 1594 1053 1662 1093
rect 1594 1019 1611 1053
rect 1645 1019 1662 1053
rect 1769 1366 1803 1446
rect 1769 1298 1803 1332
rect 1769 1230 1803 1264
rect 1769 1162 1803 1196
rect 1769 1093 1803 1128
rect 1769 1027 1803 1059
rect 1857 1366 1891 1404
rect 1857 1298 1891 1332
rect 1857 1230 1891 1264
rect 1857 1162 1891 1196
rect 1857 1093 1891 1128
rect 1945 1366 1979 1446
rect 1945 1298 1979 1332
rect 1945 1230 1979 1264
rect 1945 1162 1979 1196
rect 1945 1111 1979 1128
rect 2033 1366 2067 1404
rect 2033 1298 2067 1332
rect 2033 1230 2067 1264
rect 2033 1162 2067 1196
rect 1857 1057 1891 1059
rect 2033 1093 2067 1128
rect 2121 1366 2155 1446
rect 2121 1298 2155 1332
rect 2121 1230 2155 1264
rect 2121 1162 2155 1196
rect 2121 1111 2155 1128
rect 2260 1423 2328 1446
rect 2260 1389 2277 1423
rect 2311 1389 2328 1423
rect 2260 1349 2328 1389
rect 2260 1315 2277 1349
rect 2311 1315 2328 1349
rect 2260 1275 2328 1315
rect 2260 1241 2277 1275
rect 2311 1241 2328 1275
rect 2260 1201 2328 1241
rect 2260 1167 2277 1201
rect 2311 1167 2328 1201
rect 2260 1127 2328 1167
rect 2033 1057 2067 1059
rect 2260 1093 2277 1127
rect 2311 1093 2328 1127
rect 1857 1023 2163 1057
rect 1594 979 1662 1019
rect 1594 945 1611 979
rect 1645 945 1662 979
rect 1594 905 1662 945
rect 1594 871 1611 905
rect 1645 871 1662 905
rect 1594 822 1662 871
rect 1833 957 1867 973
rect 1987 957 2021 973
rect 700 219 734 316
rect 928 313 996 353
rect 928 279 945 313
rect 979 279 996 313
rect 700 169 734 185
rect 797 263 831 279
rect 797 195 831 229
rect 489 125 523 141
rect 329 91 392 125
rect 426 91 489 125
rect 295 75 329 91
rect 489 75 523 91
rect 603 125 637 161
rect 797 125 831 161
rect 637 91 700 125
rect 734 91 797 125
rect 603 75 637 91
rect 797 75 831 91
rect 928 239 996 279
rect 928 205 945 239
rect 979 205 996 239
rect 928 165 996 205
rect 928 131 945 165
rect 979 131 996 165
rect 928 91 996 131
rect 928 57 945 91
rect 979 57 996 91
rect 1084 333 1118 349
rect 1278 333 1312 349
rect 1463 348 1497 649
rect 1833 683 1867 923
rect 1118 299 1181 333
rect 1215 299 1278 333
rect 1084 261 1118 299
rect 1084 193 1118 227
rect 1278 261 1312 299
rect 1084 123 1118 159
rect 1084 73 1118 89
rect 1181 208 1215 224
rect 928 34 996 57
rect 1181 34 1215 174
rect 1278 193 1312 227
rect 1375 314 1497 348
rect 1594 461 1662 544
rect 1594 427 1611 461
rect 1645 427 1662 461
rect 1594 387 1662 427
rect 1594 353 1611 387
rect 1645 353 1662 387
rect 1833 433 1867 649
rect 1833 383 1867 399
rect 1981 923 1987 942
rect 1981 907 2021 923
rect 1981 831 2015 907
rect 1981 433 2015 797
rect 1981 383 2015 399
rect 2129 683 2163 1023
rect 2260 1053 2328 1093
rect 2260 1019 2277 1053
rect 2311 1019 2328 1053
rect 2435 1366 2469 1446
rect 2435 1298 2469 1332
rect 2435 1230 2469 1264
rect 2435 1162 2469 1196
rect 2435 1093 2469 1128
rect 2435 1027 2469 1059
rect 2523 1366 2557 1404
rect 2523 1298 2557 1332
rect 2523 1230 2557 1264
rect 2523 1162 2557 1196
rect 2523 1093 2557 1128
rect 2611 1366 2645 1446
rect 2611 1298 2645 1332
rect 2611 1230 2645 1264
rect 2611 1162 2645 1196
rect 2611 1111 2645 1128
rect 2699 1366 2733 1404
rect 2699 1298 2733 1332
rect 2699 1230 2733 1264
rect 2699 1162 2733 1196
rect 2523 1057 2557 1059
rect 2699 1093 2733 1128
rect 2787 1366 2821 1446
rect 2787 1298 2821 1332
rect 2787 1230 2821 1264
rect 2787 1162 2821 1196
rect 2787 1111 2821 1128
rect 2926 1423 2994 1446
rect 2926 1389 2943 1423
rect 2977 1389 2994 1423
rect 2926 1349 2994 1389
rect 2926 1315 2943 1349
rect 2977 1315 2994 1349
rect 2926 1275 2994 1315
rect 2926 1241 2943 1275
rect 2977 1241 2994 1275
rect 2926 1201 2994 1241
rect 2926 1167 2943 1201
rect 2977 1167 2994 1201
rect 2926 1127 2994 1167
rect 2699 1057 2733 1059
rect 2926 1093 2943 1127
rect 2977 1093 2994 1127
rect 2523 1023 2829 1057
rect 2260 979 2328 1019
rect 2260 945 2277 979
rect 2311 945 2328 979
rect 2260 905 2328 945
rect 2260 871 2277 905
rect 2311 871 2328 905
rect 2260 822 2328 871
rect 2499 957 2533 973
rect 2653 957 2687 973
rect 1375 217 1409 314
rect 1594 313 1662 353
rect 1594 279 1611 313
rect 1645 279 1662 313
rect 1375 167 1409 183
rect 1472 261 1506 277
rect 1472 193 1506 227
rect 1278 123 1312 159
rect 1472 123 1506 159
rect 1312 89 1375 123
rect 1409 89 1472 123
rect 1278 73 1312 89
rect 1472 73 1506 89
rect 1594 239 1662 279
rect 1594 205 1611 239
rect 1645 205 1662 239
rect 1594 165 1662 205
rect 1594 131 1611 165
rect 1645 131 1662 165
rect 1594 91 1662 131
rect 1594 57 1611 91
rect 1645 57 1662 91
rect 1750 333 1784 349
rect 1944 333 1978 349
rect 2129 348 2163 649
rect 2499 683 2533 923
rect 1784 299 1847 333
rect 1881 299 1944 333
rect 1750 261 1784 299
rect 1750 193 1784 227
rect 1944 261 1978 299
rect 1750 123 1784 159
rect 1750 73 1784 89
rect 1847 208 1881 224
rect 1594 34 1662 57
rect 1847 34 1881 174
rect 1944 193 1978 227
rect 2041 314 2163 348
rect 2260 461 2328 544
rect 2260 427 2277 461
rect 2311 427 2328 461
rect 2260 387 2328 427
rect 2260 353 2277 387
rect 2311 353 2328 387
rect 2499 433 2533 649
rect 2499 383 2533 399
rect 2647 923 2653 942
rect 2647 907 2687 923
rect 2647 905 2681 907
rect 2647 433 2681 871
rect 2647 383 2681 399
rect 2795 831 2829 1023
rect 2926 1053 2994 1093
rect 2926 1019 2943 1053
rect 2977 1019 2994 1053
rect 3101 1366 3135 1446
rect 3101 1298 3135 1332
rect 3101 1230 3135 1264
rect 3101 1162 3135 1196
rect 3101 1093 3135 1128
rect 3101 1027 3135 1059
rect 3189 1366 3223 1404
rect 3189 1298 3223 1332
rect 3189 1230 3223 1264
rect 3189 1162 3223 1196
rect 3189 1093 3223 1128
rect 3277 1366 3311 1446
rect 3277 1298 3311 1332
rect 3277 1230 3311 1264
rect 3277 1162 3311 1196
rect 3277 1111 3311 1128
rect 3365 1366 3399 1404
rect 3365 1298 3399 1332
rect 3365 1230 3399 1264
rect 3365 1162 3399 1196
rect 3189 1057 3223 1059
rect 3365 1093 3399 1128
rect 3453 1366 3487 1446
rect 3453 1298 3487 1332
rect 3453 1230 3487 1264
rect 3453 1162 3487 1196
rect 3453 1111 3487 1128
rect 3592 1423 3660 1446
rect 3592 1389 3609 1423
rect 3643 1389 3660 1423
rect 3592 1349 3660 1389
rect 3592 1315 3609 1349
rect 3643 1315 3660 1349
rect 3592 1275 3660 1315
rect 3592 1241 3609 1275
rect 3643 1241 3660 1275
rect 3592 1201 3660 1241
rect 3592 1167 3609 1201
rect 3643 1167 3660 1201
rect 3592 1127 3660 1167
rect 3365 1057 3399 1059
rect 3592 1093 3609 1127
rect 3643 1093 3660 1127
rect 3189 1023 3495 1057
rect 2926 979 2994 1019
rect 2926 945 2943 979
rect 2977 945 2994 979
rect 2926 905 2994 945
rect 2926 871 2943 905
rect 2977 871 2994 905
rect 2926 822 2994 871
rect 3165 957 3199 973
rect 3319 957 3353 973
rect 2041 217 2075 314
rect 2260 313 2328 353
rect 2260 279 2277 313
rect 2311 279 2328 313
rect 2041 167 2075 183
rect 2138 261 2172 277
rect 2138 193 2172 227
rect 1944 123 1978 159
rect 2138 123 2172 159
rect 1978 89 2041 123
rect 2075 89 2138 123
rect 1944 73 1978 89
rect 2138 73 2172 89
rect 2260 239 2328 279
rect 2260 205 2277 239
rect 2311 205 2328 239
rect 2260 165 2328 205
rect 2260 131 2277 165
rect 2311 131 2328 165
rect 2260 91 2328 131
rect 2260 57 2277 91
rect 2311 57 2328 91
rect 2416 333 2450 349
rect 2610 333 2644 349
rect 2795 348 2829 797
rect 3165 757 3199 923
rect 2450 299 2513 333
rect 2547 299 2610 333
rect 2416 261 2450 299
rect 2416 193 2450 227
rect 2610 261 2644 299
rect 2416 123 2450 159
rect 2416 73 2450 89
rect 2513 208 2547 224
rect 2260 34 2328 57
rect 2513 34 2547 174
rect 2610 193 2644 227
rect 2707 314 2829 348
rect 2926 461 2994 544
rect 2926 427 2943 461
rect 2977 427 2994 461
rect 2926 387 2994 427
rect 2926 353 2943 387
rect 2977 353 2994 387
rect 3165 433 3199 723
rect 3165 383 3199 399
rect 3313 923 3319 942
rect 3313 907 3353 923
rect 3313 757 3347 907
rect 3313 433 3347 723
rect 3313 383 3347 399
rect 3461 683 3495 1023
rect 3592 1053 3660 1093
rect 3592 1019 3609 1053
rect 3643 1019 3660 1053
rect 3767 1366 3801 1446
rect 3767 1298 3801 1332
rect 3767 1230 3801 1264
rect 3767 1162 3801 1196
rect 3767 1093 3801 1128
rect 3767 1027 3801 1059
rect 3855 1366 3889 1404
rect 3855 1298 3889 1332
rect 3855 1230 3889 1264
rect 3855 1162 3889 1196
rect 3855 1093 3889 1128
rect 3943 1366 3977 1446
rect 3943 1298 3977 1332
rect 3943 1230 3977 1264
rect 3943 1162 3977 1196
rect 3943 1111 3977 1128
rect 4031 1366 4065 1404
rect 4031 1298 4065 1332
rect 4031 1230 4065 1264
rect 4031 1162 4065 1196
rect 3855 1057 3889 1059
rect 4031 1093 4065 1128
rect 4119 1366 4153 1446
rect 4119 1298 4153 1332
rect 4119 1230 4153 1264
rect 4119 1162 4153 1196
rect 4119 1111 4153 1128
rect 4258 1423 4326 1446
rect 4258 1389 4275 1423
rect 4309 1389 4326 1423
rect 4258 1349 4326 1389
rect 4258 1315 4275 1349
rect 4309 1315 4326 1349
rect 4258 1275 4326 1315
rect 4258 1241 4275 1275
rect 4309 1241 4326 1275
rect 4258 1201 4326 1241
rect 4258 1167 4275 1201
rect 4309 1167 4326 1201
rect 4258 1127 4326 1167
rect 4031 1057 4065 1059
rect 4258 1093 4275 1127
rect 4309 1093 4326 1127
rect 3855 1023 4161 1057
rect 3592 979 3660 1019
rect 3592 945 3609 979
rect 3643 945 3660 979
rect 3592 905 3660 945
rect 3592 871 3609 905
rect 3643 871 3660 905
rect 3592 822 3660 871
rect 3831 957 3865 973
rect 3985 957 4019 973
rect 2707 217 2741 314
rect 2926 313 2994 353
rect 2926 279 2943 313
rect 2977 279 2994 313
rect 2707 167 2741 183
rect 2804 261 2838 277
rect 2804 193 2838 227
rect 2610 123 2644 159
rect 2804 123 2838 159
rect 2644 89 2707 123
rect 2741 89 2804 123
rect 2610 73 2644 89
rect 2804 73 2838 89
rect 2926 239 2994 279
rect 2926 205 2943 239
rect 2977 205 2994 239
rect 2926 165 2994 205
rect 2926 131 2943 165
rect 2977 131 2994 165
rect 2926 91 2994 131
rect 2926 57 2943 91
rect 2977 57 2994 91
rect 3082 333 3116 349
rect 3276 333 3310 349
rect 3461 348 3495 649
rect 3831 683 3865 923
rect 3116 299 3179 333
rect 3213 299 3276 333
rect 3082 261 3116 299
rect 3082 193 3116 227
rect 3276 261 3310 299
rect 3082 123 3116 159
rect 3082 73 3116 89
rect 3179 208 3213 224
rect 2926 34 2994 57
rect 3179 34 3213 174
rect 3276 193 3310 227
rect 3373 314 3495 348
rect 3592 461 3660 544
rect 3592 427 3609 461
rect 3643 427 3660 461
rect 3592 387 3660 427
rect 3592 353 3609 387
rect 3643 353 3660 387
rect 3831 433 3865 649
rect 3831 383 3865 399
rect 3979 923 3985 942
rect 3979 907 4019 923
rect 3979 831 4013 907
rect 3979 433 4013 797
rect 3979 383 4013 399
rect 4127 757 4161 1023
rect 4258 1053 4326 1093
rect 4258 1019 4275 1053
rect 4309 1019 4326 1053
rect 4258 979 4326 1019
rect 4258 945 4275 979
rect 4309 945 4326 979
rect 4258 905 4326 945
rect 4258 871 4275 905
rect 4309 871 4326 905
rect 4258 822 4326 871
rect 3373 217 3407 314
rect 3592 313 3660 353
rect 3592 279 3609 313
rect 3643 279 3660 313
rect 3373 167 3407 183
rect 3470 261 3504 277
rect 3470 193 3504 227
rect 3276 123 3310 159
rect 3470 123 3504 159
rect 3310 89 3373 123
rect 3407 89 3470 123
rect 3276 73 3310 89
rect 3470 73 3504 89
rect 3592 239 3660 279
rect 3592 205 3609 239
rect 3643 205 3660 239
rect 3592 165 3660 205
rect 3592 131 3609 165
rect 3643 131 3660 165
rect 3592 91 3660 131
rect 3592 57 3609 91
rect 3643 57 3660 91
rect 3748 333 3782 349
rect 3942 333 3976 349
rect 4127 348 4161 723
rect 3782 299 3845 333
rect 3879 299 3942 333
rect 3748 261 3782 299
rect 3748 193 3782 227
rect 3942 261 3976 299
rect 3748 123 3782 159
rect 3748 73 3782 89
rect 3845 208 3879 224
rect 3592 34 3660 57
rect 3845 34 3879 174
rect 3942 193 3976 227
rect 4039 314 4161 348
rect 4258 461 4326 544
rect 4258 427 4275 461
rect 4309 427 4326 461
rect 4258 387 4326 427
rect 4258 353 4275 387
rect 4309 353 4326 387
rect 4039 217 4073 314
rect 4258 313 4326 353
rect 4258 279 4275 313
rect 4309 279 4326 313
rect 4039 167 4073 183
rect 4136 261 4170 277
rect 4136 193 4170 227
rect 3942 123 3976 159
rect 4136 123 4170 159
rect 3976 89 4039 123
rect 4073 89 4136 123
rect 3942 73 3976 89
rect 4136 73 4170 89
rect 4258 239 4326 279
rect 4258 205 4275 239
rect 4309 205 4326 239
rect 4258 165 4326 205
rect 4258 131 4275 165
rect 4309 131 4326 165
rect 4258 91 4326 131
rect 4258 57 4275 91
rect 4309 57 4326 91
rect 4258 34 4326 57
rect -34 17 4326 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4326 17
rect -34 -34 4326 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2573 1463 2607 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3239 1463 3273 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3905 1463 3939 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 205 797 239 831
rect 427 871 461 905
rect 649 649 683 683
rect 797 723 831 757
rect 1167 723 1201 757
rect 1463 649 1497 683
rect 1833 649 1867 683
rect 1981 797 2015 831
rect 2129 649 2163 683
rect 2499 649 2533 683
rect 2647 871 2681 905
rect 2795 797 2829 831
rect 3165 723 3199 757
rect 3313 723 3347 757
rect 3461 649 3495 683
rect 3831 649 3865 683
rect 3979 797 4013 831
rect 4127 723 4161 757
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2573 -17 2607 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3239 -17 3273 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3905 -17 3939 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
<< metal1 >>
rect -34 1497 4326 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2573 1497
rect 2607 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3239 1497
rect 3273 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3905 1497
rect 3939 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4326 1497
rect -34 1445 4326 1463
rect 421 905 467 911
rect 2641 905 2687 911
rect 415 871 427 905
rect 461 871 2647 905
rect 2681 871 2693 905
rect 421 865 467 871
rect 2641 865 2687 871
rect 199 831 245 837
rect 1975 831 2021 837
rect 2789 831 2835 837
rect 3973 831 4019 837
rect 193 797 205 831
rect 239 797 1981 831
rect 2015 797 2795 831
rect 2829 797 3979 831
rect 4013 797 4025 831
rect 199 791 245 797
rect 1975 791 2021 797
rect 2789 791 2835 797
rect 3973 791 4019 797
rect 791 757 837 763
rect 1161 757 1207 763
rect 3159 757 3205 763
rect 3307 757 3353 763
rect 4121 757 4167 763
rect 785 723 797 757
rect 831 723 1167 757
rect 1201 723 3165 757
rect 3199 723 3211 757
rect 3301 723 3313 757
rect 3347 723 4127 757
rect 4161 723 4173 757
rect 791 717 837 723
rect 1161 717 1207 723
rect 3159 717 3205 723
rect 3307 717 3353 723
rect 4121 717 4167 723
rect 643 683 689 689
rect 1457 683 1503 689
rect 1827 683 1873 689
rect 2123 683 2169 689
rect 2493 683 2539 689
rect 3455 683 3501 689
rect 3825 683 3871 689
rect 637 649 649 683
rect 683 649 1463 683
rect 1497 649 1833 683
rect 1867 649 1879 683
rect 2117 649 2129 683
rect 2163 649 2499 683
rect 2533 649 2545 683
rect 3449 649 3461 683
rect 3495 649 3831 683
rect 3865 649 3877 683
rect 643 643 689 649
rect 1457 643 1503 649
rect 1827 643 1873 649
rect 2123 643 2169 649
rect 2493 643 2539 649
rect 3455 643 3501 649
rect 3825 643 3871 649
rect -34 17 4326 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2573 17
rect 2607 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3239 17
rect 3273 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3905 17
rect 3939 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4326 17
rect -34 -34 4326 -17
<< labels >>
rlabel metal1 4127 723 4161 757 1 Q
port 1 n
rlabel metal1 4127 797 4161 831 1 Q
port 2 n
rlabel metal1 4127 871 4161 905 1 Q
port 3 n
rlabel metal1 4127 945 4161 979 1 Q
port 4 n
rlabel metal1 4127 649 4161 683 1 Q
port 5 n
rlabel metal1 4127 575 4161 609 1 Q
port 6 n
rlabel metal1 4127 501 4161 535 1 Q
port 7 n
rlabel metal1 4127 427 4161 461 1 Q
port 8 n
rlabel metal1 3313 871 3347 905 1 Q
port 9 n
rlabel metal1 3313 723 3347 757 1 Q
port 10 n
rlabel metal1 3313 649 3347 683 1 Q
port 11 n
rlabel metal1 3313 575 3347 609 1 Q
port 12 n
rlabel metal1 3313 501 3347 535 1 Q
port 13 n
rlabel metal1 3313 427 3347 461 1 Q
port 14 n
rlabel metal1 3831 649 3865 683 1 QN
port 15 n
rlabel metal1 3831 871 3865 905 1 QN
port 16 n
rlabel metal1 3831 575 3865 609 1 QN
port 17 n
rlabel metal1 3831 501 3865 535 1 QN
port 18 n
rlabel metal1 3831 427 3865 461 1 QN
port 19 n
rlabel metal1 3461 427 3495 461 1 QN
port 20 n
rlabel metal1 3461 501 3495 535 1 QN
port 21 n
rlabel metal1 3461 575 3495 609 1 QN
port 22 n
rlabel metal1 3461 649 3495 683 1 QN
port 23 n
rlabel metal1 3461 871 3495 905 1 QN
port 24 n
rlabel metal1 3461 945 3495 979 1 QN
port 25 n
rlabel metal1 1315 575 1349 609 1 D
port 26 n
rlabel metal1 1315 501 1349 535 1 D
port 27 n
rlabel metal1 1315 427 1349 461 1 D
port 28 n
rlabel metal1 427 871 461 905 1 CLK
port 29 n
rlabel metal1 427 723 461 757 1 CLK
port 30 n
rlabel metal1 427 649 461 683 1 CLK
port 31 n
rlabel metal1 427 575 461 609 1 CLK
port 32 n
rlabel metal1 427 501 461 535 1 CLK
port 33 n
rlabel metal1 427 427 461 461 1 CLK
port 34 n
rlabel metal1 2647 427 2681 461 1 CLK
port 35 n
rlabel metal1 2647 501 2681 535 1 CLK
port 36 n
rlabel metal1 2647 575 2681 609 1 CLK
port 37 n
rlabel metal1 2647 649 2681 683 1 CLK
port 38 n
rlabel metal1 2647 871 2681 905 1 CLK
port 39 n
rlabel metal1 -34 1445 4326 1514 1 VPWR
port 40 n
rlabel metal1 -34 -34 4326 34 1 VGND
port 41 n
rlabel nwell 57 1463 91 1497 1 VPB
port 42 n
rlabel pwell 57 -17 91 17 1 VNB
port 43 n
<< end >>
