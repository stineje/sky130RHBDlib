`timescale 1ns/1ps

module tb ();

  logic a, b;
  

  always
  begin

  end


  initial
  begin


    $stop;
  end


endmodule
