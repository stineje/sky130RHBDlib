* SPICE3 file created from NAND2X1.ext - technology: sky130A

.subckt NAND2X1 Y A B VDD VSS
X0 VDD A Y VDD sky130_fd_pr__pfet_01v8 ad=0.00168 pd=1.368 as=0.00116 ps=9.16 w=2 l=0.15 M=2
X1 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X2 VSS A a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0 ps=0 w=3 l=0.15
X3 Y B a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0 ps=0 w=3 l=0.15
.ends
