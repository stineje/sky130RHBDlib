* SPICE3 file created from AND3X1.ext - technology: sky130A

.subckt AND3X1 Y A B C VDD GND
X0 VDD B a_277_1004 VDD pshort w=2 l=0.15 M=2
X1 GND A a_91_75 GND nshort w=3 l=0.15
X2 VDD C a_277_1004 VDD pshort w=2 l=0.15 M=2
X3 a_372_182 B a_91_75 GND nshort w=3 l=0.15
X4 a_277_1004 A VDD VDD pshort w=2 l=0.15 M=2
X5 VDD a_277_1004 Y VDD pshort w=2 l=0.15 M=2
X6 Y a_277_1004 GND GND nshort w=3 l=0.15
X7 a_277_1004 C a_372_182 GND nshort w=3 l=0.15
C0 VDD GND 3.71fF
.ends
