// File: FA.spi.pex
// Created: Tue Oct 15 15:48:52 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_FA\%GND ( 1 65 77 81 84 89 95 101 107 115 123 126 131 135 143 149 \
 157 161 164 169 173 181 189 197 205 208 213 217 220 225 229 237 245 248 253 \
 257 260 265 271 277 283 288 293 297 305 309 317 321 329 333 341 347 355 359 \
 370 373 384 387 389 401 413 415 417 429 431 443 446 458 478 490 491 492 493 \
 494 495 496 497 498 499 500 501 502 503 )
c557 ( 503 0 ) capacitor c=0.0600324f //x=37.125 //y=0.37
c558 ( 502 0 ) capacitor c=0.0699409f //x=33.86 //y=0.365
c559 ( 501 0 ) capacitor c=0.0572693f //x=31.575 //y=0.37
c560 ( 500 0 ) capacitor c=0.0207059f //x=28.74 //y=0.865
c561 ( 499 0 ) capacitor c=0.0562168f //x=26.025 //y=0.37
c562 ( 498 0 ) capacitor c=0.0207059f //x=23.19 //y=0.865
c563 ( 497 0 ) capacitor c=0.0561333f //x=20.475 //y=0.37
c564 ( 496 0 ) capacitor c=0.0209533f //x=17.64 //y=0.87
c565 ( 495 0 ) capacitor c=0.0209533f //x=14.31 //y=0.87
c566 ( 494 0 ) capacitor c=0.0561333f //x=11.595 //y=0.37
c567 ( 493 0 ) capacitor c=0.0561333f //x=9.375 //y=0.37
c568 ( 492 0 ) capacitor c=0.0209533f //x=6.54 //y=0.87
c569 ( 491 0 ) capacitor c=0.0209533f //x=3.21 //y=0.87
c570 ( 490 0 ) capacitor c=0.0582156f //x=0.495 //y=0.37
c571 ( 478 0 ) capacitor c=0.0992376f //x=36.63 //y=0
c572 ( 458 0 ) capacitor c=0.102761f //x=33.3 //y=0
c573 ( 446 0 ) capacitor c=0.0997852f //x=31.08 //y=0
c574 ( 445 0 ) capacitor c=0.00440095f //x=28.86 //y=0
c575 ( 443 0 ) capacitor c=0.100398f //x=27.75 //y=0
c576 ( 431 0 ) capacitor c=0.100609f //x=25.53 //y=0
c577 ( 430 0 ) capacitor c=0.00440095f //x=23.38 //y=0
c578 ( 429 0 ) capacitor c=0.0986577f //x=22.2 //y=0
c579 ( 417 0 ) capacitor c=0.100431f //x=19.98 //y=0
c580 ( 416 0 ) capacitor c=0.0044012f //x=17.83 //y=0
c581 ( 415 0 ) capacitor c=0.103425f //x=16.65 //y=0
c582 ( 414 0 ) capacitor c=0.0044012f //x=14.5 //y=0
c583 ( 413 0 ) capacitor c=0.0998974f //x=13.32 //y=0
c584 ( 401 0 ) capacitor c=0.0921731f //x=11.1 //y=0
c585 ( 389 0 ) capacitor c=0.101392f //x=8.88 //y=0
c586 ( 388 0 ) capacitor c=0.0044012f //x=6.73 //y=0
c587 ( 387 0 ) capacitor c=0.10347f //x=5.55 //y=0
c588 ( 386 0 ) capacitor c=0.0044012f //x=3.33 //y=0
c589 ( 384 0 ) capacitor c=0.100929f //x=2.22 //y=0
c590 ( 373 0 ) capacitor c=0.192382f //x=0.63 //y=0
c591 ( 370 0 ) capacitor c=0.198211f //x=38.48 //y=0
c592 ( 368 0 ) capacitor c=0.0360689f //x=38.315 //y=0
c593 ( 362 0 ) capacitor c=0.00587411f //x=38.23 //y=0.45
c594 ( 359 0 ) capacitor c=0.00542558f //x=38.145 //y=0.535
c595 ( 358 0 ) capacitor c=0.00479856f //x=37.745 //y=0.45
c596 ( 355 0 ) capacitor c=0.0068422f //x=37.66 //y=0.535
c597 ( 350 0 ) capacitor c=0.00592191f //x=37.26 //y=0.45
c598 ( 347 0 ) capacitor c=0.0164879f //x=37.175 //y=0
c599 ( 342 0 ) capacitor c=0.0660122f //x=36.02 //y=0
c600 ( 341 0 ) capacitor c=0.0195795f //x=36.46 //y=0
c601 ( 336 0 ) capacitor c=0.00609805f //x=35.935 //y=0.445
c602 ( 333 0 ) capacitor c=0.00508468f //x=35.85 //y=0.53
c603 ( 332 0 ) capacitor c=0.00468234f //x=35.45 //y=0.445
c604 ( 329 0 ) capacitor c=0.00551137f //x=35.365 //y=0.53
c605 ( 324 0 ) capacitor c=0.00468234f //x=34.965 //y=0.445
c606 ( 321 0 ) capacitor c=0.00533847f //x=34.88 //y=0.53
c607 ( 320 0 ) capacitor c=0.00468234f //x=34.48 //y=0.445
c608 ( 317 0 ) capacitor c=0.00625032f //x=34.395 //y=0.53
c609 ( 312 0 ) capacitor c=0.00609805f //x=33.995 //y=0.445
c610 ( 309 0 ) capacitor c=0.0195795f //x=33.91 //y=0
c611 ( 306 0 ) capacitor c=0.0360881f //x=32.765 //y=0
c612 ( 305 0 ) capacitor c=0.0160123f //x=33.13 //y=0
c613 ( 300 0 ) capacitor c=0.00583665f //x=32.68 //y=0.45
c614 ( 297 0 ) capacitor c=0.00531808f //x=32.595 //y=0.535
c615 ( 296 0 ) capacitor c=0.00479856f //x=32.195 //y=0.45
c616 ( 293 0 ) capacitor c=0.006266f //x=32.11 //y=0.535
c617 ( 288 0 ) capacitor c=0.00588377f //x=31.71 //y=0.45
c618 ( 283 0 ) capacitor c=0.0164879f //x=31.625 //y=0
c619 ( 277 0 ) capacitor c=0.0718128f //x=30.91 //y=0
c620 ( 271 0 ) capacitor c=0.038871f //x=28.845 //y=0
c621 ( 266 0 ) capacitor c=0.0360821f //x=27.215 //y=0
c622 ( 265 0 ) capacitor c=0.0160123f //x=27.58 //y=0
c623 ( 260 0 ) capacitor c=0.00583665f //x=27.13 //y=0.45
c624 ( 257 0 ) capacitor c=0.0051464f //x=27.045 //y=0.535
c625 ( 256 0 ) capacitor c=0.00479856f //x=26.645 //y=0.45
c626 ( 253 0 ) capacitor c=0.00591695f //x=26.56 //y=0.535
c627 ( 248 0 ) capacitor c=0.00588377f //x=26.16 //y=0.45
c628 ( 245 0 ) capacitor c=0.0164879f //x=26.075 //y=0
c629 ( 237 0 ) capacitor c=0.071756f //x=25.36 //y=0
c630 ( 229 0 ) capacitor c=0.038871f //x=23.295 //y=0
c631 ( 226 0 ) capacitor c=0.0360821f //x=21.655 //y=0
c632 ( 225 0 ) capacitor c=0.0164879f //x=22.03 //y=0
c633 ( 220 0 ) capacitor c=0.00588377f //x=21.57 //y=0.45
c634 ( 217 0 ) capacitor c=0.00591695f //x=21.485 //y=0.535
c635 ( 216 0 ) capacitor c=0.00479856f //x=21.085 //y=0.45
c636 ( 213 0 ) capacitor c=0.0051464f //x=21 //y=0.535
c637 ( 208 0 ) capacitor c=0.00587411f //x=20.6 //y=0.45
c638 ( 205 0 ) capacitor c=0.0160123f //x=20.515 //y=0
c639 ( 197 0 ) capacitor c=0.0719474f //x=19.81 //y=0
c640 ( 189 0 ) capacitor c=0.0388897f //x=17.745 //y=0
c641 ( 181 0 ) capacitor c=0.0719474f //x=16.48 //y=0
c642 ( 173 0 ) capacitor c=0.0388897f //x=14.415 //y=0
c643 ( 170 0 ) capacitor c=0.0360821f //x=12.785 //y=0
c644 ( 169 0 ) capacitor c=0.0160123f //x=13.15 //y=0
c645 ( 164 0 ) capacitor c=0.00587411f //x=12.7 //y=0.45
c646 ( 161 0 ) capacitor c=0.0051464f //x=12.615 //y=0.535
c647 ( 160 0 ) capacitor c=0.00479856f //x=12.215 //y=0.45
c648 ( 157 0 ) capacitor c=0.00591695f //x=12.13 //y=0.535
c649 ( 152 0 ) capacitor c=0.00592191f //x=11.73 //y=0.45
c650 ( 149 0 ) capacitor c=0.0164879f //x=11.645 //y=0
c651 ( 144 0 ) capacitor c=0.0360821f //x=10.555 //y=0
c652 ( 143 0 ) capacitor c=0.0164879f //x=10.93 //y=0
c653 ( 138 0 ) capacitor c=0.00592191f //x=10.47 //y=0.45
c654 ( 135 0 ) capacitor c=0.00591695f //x=10.385 //y=0.535
c655 ( 134 0 ) capacitor c=0.00479856f //x=9.985 //y=0.45
c656 ( 131 0 ) capacitor c=0.0051464f //x=9.9 //y=0.535
c657 ( 126 0 ) capacitor c=0.00587411f //x=9.5 //y=0.45
c658 ( 123 0 ) capacitor c=0.0160123f //x=9.415 //y=0
c659 ( 115 0 ) capacitor c=0.0719474f //x=8.71 //y=0
c660 ( 107 0 ) capacitor c=0.0388897f //x=6.645 //y=0
c661 ( 101 0 ) capacitor c=0.0719474f //x=5.38 //y=0
c662 ( 95 0 ) capacitor c=0.0389232f //x=3.315 //y=0
c663 ( 90 0 ) capacitor c=0.0360673f //x=1.685 //y=0
c664 ( 89 0 ) capacitor c=0.0160123f //x=2.05 //y=0
c665 ( 84 0 ) capacitor c=0.00587411f //x=1.6 //y=0.45
c666 ( 81 0 ) capacitor c=0.00534353f //x=1.515 //y=0.535
c667 ( 80 0 ) capacitor c=0.00479856f //x=1.115 //y=0.45
c668 ( 77 0 ) capacitor c=0.00707849f //x=1.03 //y=0.535
c669 ( 72 0 ) capacitor c=0.00592191f //x=0.63 //y=0.45
c670 ( 65 0 ) capacitor c=1.233f //x=38.48 //y=0
r671 (  482 483 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=37.745 //y=0 //x2=38.23 //y2=0
r672 (  481 482 ) resistor r=0.179272 //w=0.357 //l=0.005 //layer=li \
 //thickness=0.1 //x=37.74 //y=0 //x2=37.745 //y2=0
r673 (  479 481 ) resistor r=17.2101 //w=0.357 //l=0.48 //layer=li \
 //thickness=0.1 //x=37.26 //y=0 //x2=37.74 //y2=0
r674 (  466 467 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=35.45 //y=0 //x2=35.935 //y2=0
r675 (  465 466 ) resistor r=10.7563 //w=0.357 //l=0.3 //layer=li \
 //thickness=0.1 //x=35.15 //y=0 //x2=35.45 //y2=0
r676 (  463 465 ) resistor r=6.63305 //w=0.357 //l=0.185 //layer=li \
 //thickness=0.1 //x=34.965 //y=0 //x2=35.15 //y2=0
r677 (  462 463 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=34.48 //y=0 //x2=34.965 //y2=0
r678 (  461 462 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=34.04 //y=0 //x2=34.48 //y2=0
r679 (  459 461 ) resistor r=1.61345 //w=0.357 //l=0.045 //layer=li \
 //thickness=0.1 //x=33.995 //y=0 //x2=34.04 //y2=0
r680 (  450 451 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=32.56 //y=0 //x2=32.68 //y2=0
r681 (  448 450 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=32.195 //y=0 //x2=32.56 //y2=0
r682 (  447 448 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=31.71 //y=0 //x2=32.195 //y2=0
r683 (  435 436 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.645 //y=0 //x2=27.13 //y2=0
r684 (  434 435 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=26.27 //y=0 //x2=26.645 //y2=0
r685 (  432 434 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=26.16 //y=0 //x2=26.27 //y2=0
r686 (  421 422 ) resistor r=17.2101 //w=0.357 //l=0.48 //layer=li \
 //thickness=0.1 //x=21.09 //y=0 //x2=21.57 //y2=0
r687 (  419 421 ) resistor r=0.179272 //w=0.357 //l=0.005 //layer=li \
 //thickness=0.1 //x=21.085 //y=0 //x2=21.09 //y2=0
r688 (  418 419 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.6 //y=0 //x2=21.085 //y2=0
r689 (  405 406 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.215 //y=0 //x2=12.7 //y2=0
r690 (  404 405 ) resistor r=0.179272 //w=0.357 //l=0.005 //layer=li \
 //thickness=0.1 //x=12.21 //y=0 //x2=12.215 //y2=0
r691 (  402 404 ) resistor r=17.2101 //w=0.357 //l=0.48 //layer=li \
 //thickness=0.1 //x=11.73 //y=0 //x2=12.21 //y2=0
r692 (  393 394 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=9.985 //y=0 //x2=10.47 //y2=0
r693 (  392 393 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=9.62 //y=0 //x2=9.985 //y2=0
r694 (  390 392 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=9.5 //y=0 //x2=9.62 //y2=0
r695 (  376 377 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.115 //y=0 //x2=1.6 //y2=0
r696 (  375 376 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.115 //y2=0
r697 (  373 375 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=0.63 //y=0 //x2=0.74 //y2=0
r698 (  368 483 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.315 //y=0 //x2=38.23 //y2=0
r699 (  368 370 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=38.315 //y=0 //x2=38.48 //y2=0
r700 (  363 503 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.23 //y=0.62 //x2=38.23 //y2=0.535
r701 (  363 503 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=38.23 //y=0.62 //x2=38.23 //y2=1.225
r702 (  362 503 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.23 //y=0.45 //x2=38.23 //y2=0.535
r703 (  361 483 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.23 //y=0.17 //x2=38.23 //y2=0
r704 (  361 362 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=38.23 //y=0.17 //x2=38.23 //y2=0.45
r705 (  360 503 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.83 //y=0.535 //x2=37.745 //y2=0.535
r706 (  359 503 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.145 //y=0.535 //x2=38.23 //y2=0.535
r707 (  359 360 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=38.145 //y=0.535 //x2=37.83 //y2=0.535
r708 (  358 503 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.745 //y=0.45 //x2=37.745 //y2=0.535
r709 (  357 482 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.745 //y=0.17 //x2=37.745 //y2=0
r710 (  357 358 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=37.745 //y=0.17 //x2=37.745 //y2=0.45
r711 (  356 503 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.345 //y=0.535 //x2=37.26 //y2=0.535
r712 (  355 503 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.66 //y=0.535 //x2=37.745 //y2=0.535
r713 (  355 356 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=37.66 //y=0.535 //x2=37.345 //y2=0.535
r714 (  351 503 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.26 //y=0.62 //x2=37.26 //y2=0.535
r715 (  351 503 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=37.26 //y=0.62 //x2=37.26 //y2=1.225
r716 (  350 503 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.26 //y=0.45 //x2=37.26 //y2=0.535
r717 (  349 479 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.26 //y=0.17 //x2=37.26 //y2=0
r718 (  349 350 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=37.26 //y=0.17 //x2=37.26 //y2=0.45
r719 (  348 478 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.8 //y=0 //x2=36.63 //y2=0
r720 (  347 479 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.175 //y=0 //x2=37.26 //y2=0
r721 (  347 348 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=37.175 //y=0 //x2=36.8 //y2=0
r722 (  342 467 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.02 //y=0 //x2=35.935 //y2=0
r723 (  342 344 ) resistor r=8.60504 //w=0.357 //l=0.24 //layer=li \
 //thickness=0.1 //x=36.02 //y=0 //x2=36.26 //y2=0
r724 (  341 478 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.46 //y=0 //x2=36.63 //y2=0
r725 (  341 344 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=36.46 //y=0 //x2=36.26 //y2=0
r726 (  337 502 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.935 //y=0.615 //x2=35.935 //y2=0.53
r727 (  337 502 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=35.935 //y=0.615 //x2=35.935 //y2=0.88
r728 (  336 502 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.935 //y=0.445 //x2=35.935 //y2=0.53
r729 (  335 467 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=35.935 //y=0.17 //x2=35.935 //y2=0
r730 (  335 336 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=35.935 //y=0.17 //x2=35.935 //y2=0.445
r731 (  334 502 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.535 //y=0.53 //x2=35.45 //y2=0.53
r732 (  333 502 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.85 //y=0.53 //x2=35.935 //y2=0.53
r733 (  333 334 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=35.85 //y=0.53 //x2=35.535 //y2=0.53
r734 (  332 502 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.45 //y=0.445 //x2=35.45 //y2=0.53
r735 (  331 466 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=35.45 //y=0.17 //x2=35.45 //y2=0
r736 (  331 332 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=35.45 //y=0.17 //x2=35.45 //y2=0.445
r737 (  330 502 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=35.05 //y=0.53 //x2=34.965 //y2=0.53
r738 (  329 502 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.365 //y=0.53 //x2=35.45 //y2=0.53
r739 (  329 330 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=35.365 //y=0.53 //x2=35.05 //y2=0.53
r740 (  325 502 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=34.965 //y=0.615 //x2=34.965 //y2=0.53
r741 (  325 502 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=34.965 //y=0.615 //x2=34.965 //y2=0.88
r742 (  324 502 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=34.965 //y=0.445 //x2=34.965 //y2=0.53
r743 (  323 463 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=34.965 //y=0.17 //x2=34.965 //y2=0
r744 (  323 324 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=34.965 //y=0.17 //x2=34.965 //y2=0.445
r745 (  322 502 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.565 //y=0.53 //x2=34.48 //y2=0.53
r746 (  321 502 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=34.88 //y=0.53 //x2=34.965 //y2=0.53
r747 (  321 322 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=34.88 //y=0.53 //x2=34.565 //y2=0.53
r748 (  320 502 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.48 //y=0.445 //x2=34.48 //y2=0.53
r749 (  319 462 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=34.48 //y=0.17 //x2=34.48 //y2=0
r750 (  319 320 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=34.48 //y=0.17 //x2=34.48 //y2=0.445
r751 (  318 502 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.08 //y=0.53 //x2=33.995 //y2=0.53
r752 (  317 502 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.395 //y=0.53 //x2=34.48 //y2=0.53
r753 (  317 318 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=34.395 //y=0.53 //x2=34.08 //y2=0.53
r754 (  313 502 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.995 //y=0.615 //x2=33.995 //y2=0.53
r755 (  313 502 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=33.995 //y=0.615 //x2=33.995 //y2=1.22
r756 (  312 502 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.995 //y=0.445 //x2=33.995 //y2=0.53
r757 (  311 459 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.995 //y=0.17 //x2=33.995 //y2=0
r758 (  311 312 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=33.995 //y=0.17 //x2=33.995 //y2=0.445
r759 (  310 458 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.47 //y=0 //x2=33.3 //y2=0
r760 (  309 459 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.91 //y=0 //x2=33.995 //y2=0
r761 (  309 310 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=33.91 //y=0 //x2=33.47 //y2=0
r762 (  306 451 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.765 //y=0 //x2=32.68 //y2=0
r763 (  305 458 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.13 //y=0 //x2=33.3 //y2=0
r764 (  305 306 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=33.13 //y=0 //x2=32.765 //y2=0
r765 (  301 501 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.68 //y=0.62 //x2=32.68 //y2=0.535
r766 (  301 501 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=32.68 //y=0.62 //x2=32.68 //y2=1.225
r767 (  300 501 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.68 //y=0.45 //x2=32.68 //y2=0.535
r768 (  299 451 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.68 //y=0.17 //x2=32.68 //y2=0
r769 (  299 300 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=32.68 //y=0.17 //x2=32.68 //y2=0.45
r770 (  298 501 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.28 //y=0.535 //x2=32.195 //y2=0.535
r771 (  297 501 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.595 //y=0.535 //x2=32.68 //y2=0.535
r772 (  297 298 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=32.595 //y=0.535 //x2=32.28 //y2=0.535
r773 (  296 501 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.195 //y=0.45 //x2=32.195 //y2=0.535
r774 (  295 448 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.195 //y=0.17 //x2=32.195 //y2=0
r775 (  295 296 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=32.195 //y=0.17 //x2=32.195 //y2=0.45
r776 (  294 501 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.795 //y=0.535 //x2=31.71 //y2=0.535
r777 (  293 501 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.11 //y=0.535 //x2=32.195 //y2=0.535
r778 (  293 294 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=32.11 //y=0.535 //x2=31.795 //y2=0.535
r779 (  289 501 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.71 //y=0.62 //x2=31.71 //y2=0.535
r780 (  289 501 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=31.71 //y=0.62 //x2=31.71 //y2=1.225
r781 (  288 501 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.71 //y=0.45 //x2=31.71 //y2=0.535
r782 (  287 447 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=31.71 //y=0.17 //x2=31.71 //y2=0
r783 (  287 288 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=31.71 //y=0.17 //x2=31.71 //y2=0.45
r784 (  284 446 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=31.25 //y=0 //x2=31.08 //y2=0
r785 (  284 286 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=31.25 //y=0 //x2=31.45 //y2=0
r786 (  283 447 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.625 //y=0 //x2=31.71 //y2=0
r787 (  283 286 ) resistor r=6.27451 //w=0.357 //l=0.175 //layer=li \
 //thickness=0.1 //x=31.625 //y=0 //x2=31.45 //y2=0
r788 (  278 445 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.015 //y=0 //x2=28.93 //y2=0
r789 (  278 280 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=29.015 //y=0 //x2=29.97 //y2=0
r790 (  277 446 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.91 //y=0 //x2=31.08 //y2=0
r791 (  277 280 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=30.91 //y=0 //x2=29.97 //y2=0
r792 (  273 445 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=28.93 //y=0.17 //x2=28.93 //y2=0
r793 (  273 500 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=28.93 //y=0.17 //x2=28.93 //y2=0.955
r794 (  272 443 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.92 //y=0 //x2=27.75 //y2=0
r795 (  271 445 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.845 //y=0 //x2=28.93 //y2=0
r796 (  271 272 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=28.845 //y=0 //x2=27.92 //y2=0
r797 (  266 436 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.215 //y=0 //x2=27.13 //y2=0
r798 (  266 268 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=27.215 //y=0 //x2=27.38 //y2=0
r799 (  265 443 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.58 //y=0 //x2=27.75 //y2=0
r800 (  265 268 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=27.58 //y=0 //x2=27.38 //y2=0
r801 (  261 499 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.13 //y=0.62 //x2=27.13 //y2=0.535
r802 (  261 499 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=27.13 //y=0.62 //x2=27.13 //y2=1.225
r803 (  260 499 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.13 //y=0.45 //x2=27.13 //y2=0.535
r804 (  259 436 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.13 //y=0.17 //x2=27.13 //y2=0
r805 (  259 260 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=27.13 //y=0.17 //x2=27.13 //y2=0.45
r806 (  258 499 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.73 //y=0.535 //x2=26.645 //y2=0.535
r807 (  257 499 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.045 //y=0.535 //x2=27.13 //y2=0.535
r808 (  257 258 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=27.045 //y=0.535 //x2=26.73 //y2=0.535
r809 (  256 499 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.645 //y=0.45 //x2=26.645 //y2=0.535
r810 (  255 435 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.645 //y=0.17 //x2=26.645 //y2=0
r811 (  255 256 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=26.645 //y=0.17 //x2=26.645 //y2=0.45
r812 (  254 499 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.245 //y=0.535 //x2=26.16 //y2=0.535
r813 (  253 499 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.56 //y=0.535 //x2=26.645 //y2=0.535
r814 (  253 254 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=26.56 //y=0.535 //x2=26.245 //y2=0.535
r815 (  249 499 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.16 //y=0.62 //x2=26.16 //y2=0.535
r816 (  249 499 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=26.16 //y=0.62 //x2=26.16 //y2=1.225
r817 (  248 499 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.16 //y=0.45 //x2=26.16 //y2=0.535
r818 (  247 432 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.16 //y=0.17 //x2=26.16 //y2=0
r819 (  247 248 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=26.16 //y=0.17 //x2=26.16 //y2=0.45
r820 (  246 431 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.7 //y=0 //x2=25.53 //y2=0
r821 (  245 432 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.075 //y=0 //x2=26.16 //y2=0
r822 (  245 246 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=26.075 //y=0 //x2=25.7 //y2=0
r823 (  240 242 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=23.68 //y=0 //x2=24.79 //y2=0
r824 (  238 430 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.465 //y=0 //x2=23.38 //y2=0
r825 (  238 240 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=23.465 //y=0 //x2=23.68 //y2=0
r826 (  237 431 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.36 //y=0 //x2=25.53 //y2=0
r827 (  237 242 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=25.36 //y=0 //x2=24.79 //y2=0
r828 (  233 430 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.38 //y=0.17 //x2=23.38 //y2=0
r829 (  233 498 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=23.38 //y=0.17 //x2=23.38 //y2=0.955
r830 (  230 429 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.37 //y=0 //x2=22.2 //y2=0
r831 (  230 232 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=22.37 //y=0 //x2=22.57 //y2=0
r832 (  229 430 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.295 //y=0 //x2=23.38 //y2=0
r833 (  229 232 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=23.295 //y=0 //x2=22.57 //y2=0
r834 (  226 422 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.655 //y=0 //x2=21.57 //y2=0
r835 (  225 429 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.03 //y=0 //x2=22.2 //y2=0
r836 (  225 226 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=22.03 //y=0 //x2=21.655 //y2=0
r837 (  221 497 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.57 //y=0.62 //x2=21.57 //y2=0.535
r838 (  221 497 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=21.57 //y=0.62 //x2=21.57 //y2=1.225
r839 (  220 497 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.57 //y=0.45 //x2=21.57 //y2=0.535
r840 (  219 422 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.57 //y=0.17 //x2=21.57 //y2=0
r841 (  219 220 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=21.57 //y=0.17 //x2=21.57 //y2=0.45
r842 (  218 497 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.17 //y=0.535 //x2=21.085 //y2=0.535
r843 (  217 497 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.485 //y=0.535 //x2=21.57 //y2=0.535
r844 (  217 218 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=21.485 //y=0.535 //x2=21.17 //y2=0.535
r845 (  216 497 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.085 //y=0.45 //x2=21.085 //y2=0.535
r846 (  215 419 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.085 //y=0.17 //x2=21.085 //y2=0
r847 (  215 216 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=21.085 //y=0.17 //x2=21.085 //y2=0.45
r848 (  214 497 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.685 //y=0.535 //x2=20.6 //y2=0.535
r849 (  213 497 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21 //y=0.535 //x2=21.085 //y2=0.535
r850 (  213 214 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=21 //y=0.535 //x2=20.685 //y2=0.535
r851 (  209 497 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.6 //y=0.62 //x2=20.6 //y2=0.535
r852 (  209 497 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=20.6 //y=0.62 //x2=20.6 //y2=1.225
r853 (  208 497 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.6 //y=0.45 //x2=20.6 //y2=0.535
r854 (  207 418 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.6 //y=0.17 //x2=20.6 //y2=0
r855 (  207 208 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=20.6 //y=0.17 //x2=20.6 //y2=0.45
r856 (  206 417 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.15 //y=0 //x2=19.98 //y2=0
r857 (  205 418 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.515 //y=0 //x2=20.6 //y2=0
r858 (  205 206 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=20.515 //y=0 //x2=20.15 //y2=0
r859 (  200 202 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=18.5 //y=0 //x2=19.61 //y2=0
r860 (  198 416 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.915 //y=0 //x2=17.83 //y2=0
r861 (  198 200 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=17.915 //y=0 //x2=18.5 //y2=0
r862 (  197 417 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.81 //y=0 //x2=19.98 //y2=0
r863 (  197 202 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=19.81 //y=0 //x2=19.61 //y2=0
r864 (  193 416 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.83 //y=0.17 //x2=17.83 //y2=0
r865 (  193 496 ) resistor r=54.0749 //w=0.187 //l=0.79 //layer=li \
 //thickness=0.1 //x=17.83 //y=0.17 //x2=17.83 //y2=0.96
r866 (  190 415 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.82 //y=0 //x2=16.65 //y2=0
r867 (  190 192 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=16.82 //y=0 //x2=17.39 //y2=0
r868 (  189 416 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.745 //y=0 //x2=17.83 //y2=0
r869 (  189 192 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=17.745 //y=0 //x2=17.39 //y2=0
r870 (  184 186 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=14.8 //y=0 //x2=15.91 //y2=0
r871 (  182 414 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.585 //y=0 //x2=14.5 //y2=0
r872 (  182 184 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=14.585 //y=0 //x2=14.8 //y2=0
r873 (  181 415 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.48 //y=0 //x2=16.65 //y2=0
r874 (  181 186 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=16.48 //y=0 //x2=15.91 //y2=0
r875 (  177 414 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.5 //y=0.17 //x2=14.5 //y2=0
r876 (  177 495 ) resistor r=54.0749 //w=0.187 //l=0.79 //layer=li \
 //thickness=0.1 //x=14.5 //y=0.17 //x2=14.5 //y2=0.96
r877 (  174 413 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.49 //y=0 //x2=13.32 //y2=0
r878 (  174 176 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=13.49 //y=0 //x2=13.69 //y2=0
r879 (  173 414 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.415 //y=0 //x2=14.5 //y2=0
r880 (  173 176 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=14.415 //y=0 //x2=13.69 //y2=0
r881 (  170 406 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.785 //y=0 //x2=12.7 //y2=0
r882 (  169 413 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.15 //y=0 //x2=13.32 //y2=0
r883 (  169 170 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=13.15 //y=0 //x2=12.785 //y2=0
r884 (  165 494 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.7 //y=0.62 //x2=12.7 //y2=0.535
r885 (  165 494 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=12.7 //y=0.62 //x2=12.7 //y2=1.225
r886 (  164 494 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.7 //y=0.45 //x2=12.7 //y2=0.535
r887 (  163 406 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.7 //y=0.17 //x2=12.7 //y2=0
r888 (  163 164 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=12.7 //y=0.17 //x2=12.7 //y2=0.45
r889 (  162 494 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.3 //y=0.535 //x2=12.215 //y2=0.535
r890 (  161 494 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.615 //y=0.535 //x2=12.7 //y2=0.535
r891 (  161 162 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=12.615 //y=0.535 //x2=12.3 //y2=0.535
r892 (  160 494 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.215 //y=0.45 //x2=12.215 //y2=0.535
r893 (  159 405 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.215 //y=0.17 //x2=12.215 //y2=0
r894 (  159 160 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=12.215 //y=0.17 //x2=12.215 //y2=0.45
r895 (  158 494 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.815 //y=0.535 //x2=11.73 //y2=0.535
r896 (  157 494 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.13 //y=0.535 //x2=12.215 //y2=0.535
r897 (  157 158 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=12.13 //y=0.535 //x2=11.815 //y2=0.535
r898 (  153 494 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.73 //y=0.62 //x2=11.73 //y2=0.535
r899 (  153 494 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=11.73 //y=0.62 //x2=11.73 //y2=1.225
r900 (  152 494 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.73 //y=0.45 //x2=11.73 //y2=0.535
r901 (  151 402 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.73 //y=0.17 //x2=11.73 //y2=0
r902 (  151 152 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=11.73 //y=0.17 //x2=11.73 //y2=0.45
r903 (  150 401 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.27 //y=0 //x2=11.1 //y2=0
r904 (  149 402 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.645 //y=0 //x2=11.73 //y2=0
r905 (  149 150 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=11.645 //y=0 //x2=11.27 //y2=0
r906 (  144 394 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.555 //y=0 //x2=10.47 //y2=0
r907 (  144 146 ) resistor r=6.27451 //w=0.357 //l=0.175 //layer=li \
 //thickness=0.1 //x=10.555 //y=0 //x2=10.73 //y2=0
r908 (  143 401 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.93 //y=0 //x2=11.1 //y2=0
r909 (  143 146 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=10.93 //y=0 //x2=10.73 //y2=0
r910 (  139 493 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.47 //y=0.62 //x2=10.47 //y2=0.535
r911 (  139 493 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=10.47 //y=0.62 //x2=10.47 //y2=1.225
r912 (  138 493 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.47 //y=0.45 //x2=10.47 //y2=0.535
r913 (  137 394 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.47 //y=0.17 //x2=10.47 //y2=0
r914 (  137 138 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=10.47 //y=0.17 //x2=10.47 //y2=0.45
r915 (  136 493 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.07 //y=0.535 //x2=9.985 //y2=0.535
r916 (  135 493 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.385 //y=0.535 //x2=10.47 //y2=0.535
r917 (  135 136 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=10.385 //y=0.535 //x2=10.07 //y2=0.535
r918 (  134 493 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.985 //y=0.45 //x2=9.985 //y2=0.535
r919 (  133 393 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.985 //y=0.17 //x2=9.985 //y2=0
r920 (  133 134 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=9.985 //y=0.17 //x2=9.985 //y2=0.45
r921 (  132 493 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.585 //y=0.535 //x2=9.5 //y2=0.535
r922 (  131 493 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.9 //y=0.535 //x2=9.985 //y2=0.535
r923 (  131 132 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=9.9 //y=0.535 //x2=9.585 //y2=0.535
r924 (  127 493 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.5 //y=0.62 //x2=9.5 //y2=0.535
r925 (  127 493 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=9.5 //y=0.62 //x2=9.5 //y2=1.225
r926 (  126 493 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.5 //y=0.45 //x2=9.5 //y2=0.535
r927 (  125 390 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.5 //y=0.17 //x2=9.5 //y2=0
r928 (  125 126 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=9.5 //y=0.17 //x2=9.5 //y2=0.45
r929 (  124 389 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.05 //y=0 //x2=8.88 //y2=0
r930 (  123 390 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.415 //y=0 //x2=9.5 //y2=0
r931 (  123 124 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=9.415 //y=0 //x2=9.05 //y2=0
r932 (  118 120 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=7.03 //y=0 //x2=8.14 //y2=0
r933 (  116 388 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.815 //y=0 //x2=6.73 //y2=0
r934 (  116 118 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=6.815 //y=0 //x2=7.03 //y2=0
r935 (  115 389 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.71 //y=0 //x2=8.88 //y2=0
r936 (  115 120 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=8.71 //y=0 //x2=8.14 //y2=0
r937 (  111 388 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.73 //y=0.17 //x2=6.73 //y2=0
r938 (  111 492 ) resistor r=54.0749 //w=0.187 //l=0.79 //layer=li \
 //thickness=0.1 //x=6.73 //y=0.17 //x2=6.73 //y2=0.96
r939 (  108 387 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.72 //y=0 //x2=5.55 //y2=0
r940 (  108 110 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=5.72 //y=0 //x2=5.92 //y2=0
r941 (  107 388 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.645 //y=0 //x2=6.73 //y2=0
r942 (  107 110 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=6.645 //y=0 //x2=5.92 //y2=0
r943 (  102 386 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.485 //y=0 //x2=3.4 //y2=0
r944 (  102 104 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=3.485 //y=0 //x2=4.44 //y2=0
r945 (  101 387 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.38 //y=0 //x2=5.55 //y2=0
r946 (  101 104 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=5.38 //y=0 //x2=4.44 //y2=0
r947 (  97 386 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.4 //y=0.17 //x2=3.4 //y2=0
r948 (  97 491 ) resistor r=54.0749 //w=0.187 //l=0.79 //layer=li \
 //thickness=0.1 //x=3.4 //y=0.17 //x2=3.4 //y2=0.96
r949 (  96 384 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.39 //y=0 //x2=2.22 //y2=0
r950 (  95 386 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.315 //y=0 //x2=3.4 //y2=0
r951 (  95 96 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=3.315 //y=0 //x2=2.39 //y2=0
r952 (  90 377 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.685 //y=0 //x2=1.6 //y2=0
r953 (  90 92 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=1.685 //y=0 //x2=1.85 //y2=0
r954 (  89 384 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.05 //y=0 //x2=2.22 //y2=0
r955 (  89 92 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=2.05 //y=0 //x2=1.85 //y2=0
r956 (  85 490 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=0.535
r957 (  85 490 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=1.225
r958 (  84 490 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.45 //x2=1.6 //y2=0.535
r959 (  83 377 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0
r960 (  83 84 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0.45
r961 (  82 490 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.2 //y=0.535 //x2=1.115 //y2=0.535
r962 (  81 490 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.6 //y2=0.535
r963 (  81 82 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.2 //y2=0.535
r964 (  80 490 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.45 //x2=1.115 //y2=0.535
r965 (  79 376 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0
r966 (  79 80 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0.45
r967 (  78 490 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.715 //y=0.535 //x2=0.63 //y2=0.535
r968 (  77 490 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=1.115 //y2=0.535
r969 (  77 78 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=0.715 //y2=0.535
r970 (  73 490 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=0.535
r971 (  73 490 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=1.225
r972 (  72 490 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.45 //x2=0.63 //y2=0.535
r973 (  71 373 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0
r974 (  71 72 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0.45
r975 (  65 370 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=38.48 //y=0 //x2=38.48 //y2=0
r976 (  63 481 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37.74 //y=0 //x2=37.74 //y2=0
r977 (  63 65 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=37.74 //y=0 //x2=38.48 //y2=0
r978 (  61 344 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=36.26 //y=0 //x2=36.26 //y2=0
r979 (  61 63 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=36.26 //y=0 //x2=37.74 //y2=0
r980 (  59 465 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.15 //y=0 //x2=35.15 //y2=0
r981 (  59 61 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=35.15 //y=0 //x2=36.26 //y2=0
r982 (  57 461 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.04 //y=0 //x2=34.04 //y2=0
r983 (  57 59 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=34.04 //y=0 //x2=35.15 //y2=0
r984 (  55 450 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.56 //y=0 //x2=32.56 //y2=0
r985 (  55 57 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=32.56 //y=0 //x2=34.04 //y2=0
r986 (  53 286 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.45 //y=0 //x2=31.45 //y2=0
r987 (  53 55 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.45 //y=0 //x2=32.56 //y2=0
r988 (  51 280 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=29.97 //y=0 //x2=29.97 //y2=0
r989 (  51 53 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=29.97 //y=0 //x2=31.45 //y2=0
r990 (  49 445 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.86 //y=0 //x2=28.86 //y2=0
r991 (  49 51 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=28.86 //y=0 //x2=29.97 //y2=0
r992 (  47 268 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.38 //y=0 //x2=27.38 //y2=0
r993 (  47 49 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=27.38 //y=0 //x2=28.86 //y2=0
r994 (  45 434 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=26.27 //y=0 //x2=26.27 //y2=0
r995 (  45 47 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=26.27 //y=0 //x2=27.38 //y2=0
r996 (  43 242 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=0 //x2=24.79 //y2=0
r997 (  43 45 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=0 //x2=26.27 //y2=0
r998 (  41 240 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=0 //x2=23.68 //y2=0
r999 (  41 43 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=23.68 //y=0 //x2=24.79 //y2=0
r1000 (  39 232 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.57 //y=0 //x2=22.57 //y2=0
r1001 (  39 41 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.57 //y=0 //x2=23.68 //y2=0
r1002 (  37 421 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=0 //x2=21.09 //y2=0
r1003 (  37 39 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=0 //x2=22.57 //y2=0
r1004 (  35 202 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.61 //y=0 //x2=19.61 //y2=0
r1005 (  35 37 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=19.61 //y=0 //x2=21.09 //y2=0
r1006 (  32 200 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=0 //x2=18.5 //y2=0
r1007 (  30 192 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=0 //x2=17.39 //y2=0
r1008 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=0 //x2=18.5 //y2=0
r1009 (  28 186 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.91 //y=0 //x2=15.91 //y2=0
r1010 (  28 30 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=15.91 //y=0 //x2=17.39 //y2=0
r1011 (  26 184 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.8 //y=0 //x2=14.8 //y2=0
r1012 (  26 28 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.8 //y=0 //x2=15.91 //y2=0
r1013 (  24 176 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=0 //x2=13.69 //y2=0
r1014 (  24 26 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=13.69 //y=0 //x2=14.8 //y2=0
r1015 (  22 404 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.21 //y=0 //x2=12.21 //y2=0
r1016 (  22 24 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.21 //y=0 //x2=13.69 //y2=0
r1017 (  20 146 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.73 //y=0 //x2=10.73 //y2=0
r1018 (  20 22 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=0 //x2=12.21 //y2=0
r1019 (  18 392 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.62 //y=0 //x2=9.62 //y2=0
r1020 (  18 20 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.62 //y=0 //x2=10.73 //y2=0
r1021 (  16 120 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.14 //y=0 //x2=8.14 //y2=0
r1022 (  16 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.14 //y=0 //x2=9.62 //y2=0
r1023 (  14 118 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=0 //x2=7.03 //y2=0
r1024 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=0 //x2=8.14 //y2=0
r1025 (  12 110 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.92 //y=0 //x2=5.92 //y2=0
r1026 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.92 //y=0 //x2=7.03 //y2=0
r1027 (  10 104 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r1028 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.92 //y2=0
r1029 (  8 386 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=3.33 //y=0 //x2=3.33 //y2=0
r1030 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=0 //x2=4.44 //y2=0
r1031 (  6 92 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r1032 (  6 8 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=3.33 //y2=0
r1033 (  3 375 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r1034 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r1035 (  1 35 ) resistor r=0.0768272 //w=0.301 //l=0.185 //layer=m1 \
 //thickness=0.36 //x=19.425 //y=0 //x2=19.61 //y2=0
r1036 (  1 32 ) resistor r=0.384136 //w=0.301 //l=0.925 //layer=m1 \
 //thickness=0.36 //x=19.425 //y=0 //x2=18.5 //y2=0
ends PM_FA\%GND

subckt PM_FA\%VDD ( 1 65 77 85 91 99 105 113 121 129 137 143 151 161 165 173 \
 181 189 197 205 215 219 229 239 247 251 259 267 273 281 291 315 327 337 353 \
 366 370 372 374 376 380 383 385 387 390 395 399 403 407 409 412 413 414 415 \
 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433 434 \
 435 436 )
c530 ( 436 0 ) capacitor c=0.0451925f //x=38.04 //y=5.02
c531 ( 435 0 ) capacitor c=0.0423715f //x=37.17 //y=5.02
c532 ( 434 0 ) capacitor c=0.0256052f //x=34.385 //y=5.025
c533 ( 433 0 ) capacitor c=0.0436617f //x=32.49 //y=5.02
c534 ( 432 0 ) capacitor c=0.042362f //x=31.62 //y=5.02
c535 ( 431 0 ) capacitor c=0.0382536f //x=30.155 //y=5.02
c536 ( 430 0 ) capacitor c=0.024222f //x=29.275 //y=5.02
c537 ( 429 0 ) capacitor c=0.0488152f //x=28.405 //y=5.02
c538 ( 428 0 ) capacitor c=0.0428352f //x=26.94 //y=5.02
c539 ( 427 0 ) capacitor c=0.0420515f //x=26.07 //y=5.02
c540 ( 426 0 ) capacitor c=0.0379601f //x=24.605 //y=5.02
c541 ( 425 0 ) capacitor c=0.0239037f //x=23.725 //y=5.02
c542 ( 424 0 ) capacitor c=0.0488145f //x=22.855 //y=5.02
c543 ( 423 0 ) capacitor c=0.0418661f //x=21.38 //y=5.02
c544 ( 422 0 ) capacitor c=0.0431307f //x=20.52 //y=5.02
c545 ( 421 0 ) capacitor c=0.0265379f //x=17.735 //y=5.02
c546 ( 420 0 ) capacitor c=0.026371f //x=14.405 //y=5.02
c547 ( 419 0 ) capacitor c=0.0428352f //x=12.51 //y=5.02
c548 ( 418 0 ) capacitor c=0.0418661f //x=11.64 //y=5.02
c549 ( 417 0 ) capacitor c=0.0418242f //x=10.28 //y=5.02
c550 ( 416 0 ) capacitor c=0.0433633f //x=9.42 //y=5.02
c551 ( 415 0 ) capacitor c=0.0266033f //x=6.635 //y=5.02
c552 ( 414 0 ) capacitor c=0.0265296f //x=3.305 //y=5.02
c553 ( 413 0 ) capacitor c=0.0432963f //x=1.41 //y=5.02
c554 ( 412 0 ) capacitor c=0.0421443f //x=0.54 //y=5.02
c555 ( 411 0 ) capacitor c=0.00591168f //x=38.185 //y=7.4
c556 ( 410 0 ) capacitor c=0.00591168f //x=37.305 //y=7.4
c557 ( 409 0 ) capacitor c=0.109776f //x=36.63 //y=7.4
c558 ( 408 0 ) capacitor c=0.00591168f //x=34.53 //y=7.4
c559 ( 407 0 ) capacitor c=0.112698f //x=33.3 //y=7.4
c560 ( 406 0 ) capacitor c=0.00591168f //x=32.56 //y=7.4
c561 ( 404 0 ) capacitor c=0.00591168f //x=31.755 //y=7.4
c562 ( 403 0 ) capacitor c=0.110461f //x=31.08 //y=7.4
c563 ( 402 0 ) capacitor c=0.00591168f //x=30.3 //y=7.4
c564 ( 401 0 ) capacitor c=0.00591168f //x=29.42 //y=7.4
c565 ( 400 0 ) capacitor c=0.00591168f //x=28.54 //y=7.4
c566 ( 399 0 ) capacitor c=0.117626f //x=27.75 //y=7.4
c567 ( 398 0 ) capacitor c=0.00591168f //x=27.085 //y=7.4
c568 ( 397 0 ) capacitor c=0.00591168f //x=26.27 //y=7.4
c569 ( 395 0 ) capacitor c=0.111282f //x=25.53 //y=7.4
c570 ( 394 0 ) capacitor c=0.00591168f //x=24.79 //y=7.4
c571 ( 392 0 ) capacitor c=0.00591168f //x=23.87 //y=7.4
c572 ( 391 0 ) capacitor c=0.00591168f //x=22.99 //y=7.4
c573 ( 390 0 ) capacitor c=0.115106f //x=22.2 //y=7.4
c574 ( 389 0 ) capacitor c=0.00591168f //x=21.525 //y=7.4
c575 ( 388 0 ) capacitor c=0.00591168f //x=20.645 //y=7.4
c576 ( 387 0 ) capacitor c=0.106476f //x=19.98 //y=7.4
c577 ( 386 0 ) capacitor c=0.00591168f //x=17.88 //y=7.4
c578 ( 385 0 ) capacitor c=0.112325f //x=16.65 //y=7.4
c579 ( 384 0 ) capacitor c=0.00591168f //x=14.55 //y=7.4
c580 ( 383 0 ) capacitor c=0.112188f //x=13.32 //y=7.4
c581 ( 382 0 ) capacitor c=0.00591168f //x=12.655 //y=7.4
c582 ( 381 0 ) capacitor c=0.00591168f //x=11.775 //y=7.4
c583 ( 380 0 ) capacitor c=0.105409f //x=11.1 //y=7.4
c584 ( 379 0 ) capacitor c=0.00591168f //x=10.425 //y=7.4
c585 ( 378 0 ) capacitor c=0.00591168f //x=9.62 //y=7.4
c586 ( 376 0 ) capacitor c=0.105229f //x=8.88 //y=7.4
c587 ( 375 0 ) capacitor c=0.00591168f //x=6.78 //y=7.4
c588 ( 374 0 ) capacitor c=0.111763f //x=5.55 //y=7.4
c589 ( 373 0 ) capacitor c=0.00591168f //x=3.45 //y=7.4
c590 ( 372 0 ) capacitor c=0.111559f //x=2.22 //y=7.4
c591 ( 371 0 ) capacitor c=0.00591168f //x=1.555 //y=7.4
c592 ( 370 0 ) capacitor c=0.232987f //x=0.74 //y=7.4
c593 ( 366 0 ) capacitor c=0.228884f //x=38.48 //y=7.4
c594 ( 353 0 ) capacitor c=0.0287207f //x=38.1 //y=7.4
c595 ( 345 0 ) capacitor c=0.0216067f //x=37.22 //y=7.4
c596 ( 337 0 ) capacitor c=0.0778183f //x=36.46 //y=7.4
c597 ( 327 0 ) capacitor c=0.0465804f //x=34.445 //y=7.4
c598 ( 323 0 ) capacitor c=0.0210379f //x=33.13 //y=7.4
c599 ( 315 0 ) capacitor c=0.0287207f //x=32.55 //y=7.4
c600 ( 305 0 ) capacitor c=0.0216067f //x=31.67 //y=7.4
c601 ( 301 0 ) capacitor c=0.0275781f //x=30.91 //y=7.4
c602 ( 291 0 ) capacitor c=0.0285035f //x=30.215 //y=7.4
c603 ( 281 0 ) capacitor c=0.0291677f //x=29.335 //y=7.4
c604 ( 273 0 ) capacitor c=0.0240981f //x=28.455 //y=7.4
c605 ( 267 0 ) capacitor c=0.0181526f //x=27.58 //y=7.4
c606 ( 259 0 ) capacitor c=0.0288667f //x=27 //y=7.4
c607 ( 251 0 ) capacitor c=0.0186283f //x=26.12 //y=7.4
c608 ( 247 0 ) capacitor c=0.0236224f //x=25.36 //y=7.4
c609 ( 239 0 ) capacitor c=0.0288042f //x=24.665 //y=7.4
c610 ( 229 0 ) capacitor c=0.02888f //x=23.785 //y=7.4
c611 ( 219 0 ) capacitor c=0.0240981f //x=22.905 //y=7.4
c612 ( 215 0 ) capacitor c=0.0186283f //x=22.03 //y=7.4
c613 ( 205 0 ) capacitor c=0.0288667f //x=21.44 //y=7.4
c614 ( 197 0 ) capacitor c=0.0181526f //x=20.56 //y=7.4
c615 ( 189 0 ) capacitor c=0.0746972f //x=19.81 //y=7.4
c616 ( 181 0 ) capacitor c=0.0428451f //x=17.795 //y=7.4
c617 ( 173 0 ) capacitor c=0.0746972f //x=16.48 //y=7.4
c618 ( 165 0 ) capacitor c=0.0428451f //x=14.465 //y=7.4
c619 ( 161 0 ) capacitor c=0.0181526f //x=13.15 //y=7.4
c620 ( 151 0 ) capacitor c=0.0288667f //x=12.57 //y=7.4
c621 ( 143 0 ) capacitor c=0.0186283f //x=11.69 //y=7.4
c622 ( 137 0 ) capacitor c=0.0186283f //x=10.93 //y=7.4
c623 ( 129 0 ) capacitor c=0.0290039f //x=10.34 //y=7.4
c624 ( 121 0 ) capacitor c=0.0181526f //x=9.46 //y=7.4
c625 ( 113 0 ) capacitor c=0.0747638f //x=8.71 //y=7.4
c626 ( 105 0 ) capacitor c=0.042882f //x=6.695 //y=7.4
c627 ( 99 0 ) capacitor c=0.074629f //x=5.38 //y=7.4
c628 ( 91 0 ) capacitor c=0.042884f //x=3.365 //y=7.4
c629 ( 85 0 ) capacitor c=0.0181526f //x=2.05 //y=7.4
c630 ( 77 0 ) capacitor c=0.0291066f //x=1.47 //y=7.4
c631 ( 65 0 ) capacitor c=1.2943f //x=38.48 //y=7.4
r632 (  364 411 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.27 //y=7.4 //x2=38.185 //y2=7.4
r633 (  364 366 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=38.27 //y=7.4 //x2=38.48 //y2=7.4
r634 (  357 411 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.185 //y=7.23 //x2=38.185 //y2=7.4
r635 (  357 436 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=38.185 //y=7.23 //x2=38.185 //y2=6.405
r636 (  354 410 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.39 //y=7.4 //x2=37.305 //y2=7.4
r637 (  354 356 ) resistor r=12.549 //w=0.357 //l=0.35 //layer=li \
 //thickness=0.1 //x=37.39 //y=7.4 //x2=37.74 //y2=7.4
r638 (  353 411 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.1 //y=7.4 //x2=38.185 //y2=7.4
r639 (  353 356 ) resistor r=12.9076 //w=0.357 //l=0.36 //layer=li \
 //thickness=0.1 //x=38.1 //y=7.4 //x2=37.74 //y2=7.4
r640 (  347 410 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.305 //y=7.23 //x2=37.305 //y2=7.4
r641 (  347 435 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=37.305 //y=7.23 //x2=37.305 //y2=6.405
r642 (  346 409 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.8 //y=7.4 //x2=36.63 //y2=7.4
r643 (  345 410 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.22 //y=7.4 //x2=37.305 //y2=7.4
r644 (  345 346 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=37.22 //y=7.4 //x2=36.8 //y2=7.4
r645 (  340 342 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=35.15 //y=7.4 //x2=36.26 //y2=7.4
r646 (  338 408 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.615 //y=7.4 //x2=34.53 //y2=7.4
r647 (  338 340 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=34.615 //y=7.4 //x2=35.15 //y2=7.4
r648 (  337 409 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.46 //y=7.4 //x2=36.63 //y2=7.4
r649 (  337 342 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=36.46 //y=7.4 //x2=36.26 //y2=7.4
r650 (  331 408 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=34.53 //y=7.23 //x2=34.53 //y2=7.4
r651 (  331 434 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=34.53 //y=7.23 //x2=34.53 //y2=6.74
r652 (  328 407 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.47 //y=7.4 //x2=33.3 //y2=7.4
r653 (  328 330 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=33.47 //y=7.4 //x2=34.04 //y2=7.4
r654 (  327 408 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.445 //y=7.4 //x2=34.53 //y2=7.4
r655 (  327 330 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=34.445 //y=7.4 //x2=34.04 //y2=7.4
r656 (  324 406 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.72 //y=7.4 //x2=32.635 //y2=7.4
r657 (  323 407 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.13 //y=7.4 //x2=33.3 //y2=7.4
r658 (  323 324 ) resistor r=14.7003 //w=0.357 //l=0.41 //layer=li \
 //thickness=0.1 //x=33.13 //y=7.4 //x2=32.72 //y2=7.4
r659 (  317 406 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.635 //y=7.23 //x2=32.635 //y2=7.4
r660 (  317 433 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=32.635 //y=7.23 //x2=32.635 //y2=6.405
r661 (  316 404 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.84 //y=7.4 //x2=31.755 //y2=7.4
r662 (  315 406 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.55 //y=7.4 //x2=32.635 //y2=7.4
r663 (  315 316 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=32.55 //y=7.4 //x2=31.84 //y2=7.4
r664 (  309 404 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=31.755 //y=7.23 //x2=31.755 //y2=7.4
r665 (  309 432 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=31.755 //y=7.23 //x2=31.755 //y2=6.405
r666 (  306 403 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=31.25 //y=7.4 //x2=31.08 //y2=7.4
r667 (  306 308 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=31.25 //y=7.4 //x2=31.45 //y2=7.4
r668 (  305 404 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.67 //y=7.4 //x2=31.755 //y2=7.4
r669 (  305 308 ) resistor r=7.88796 //w=0.357 //l=0.22 //layer=li \
 //thickness=0.1 //x=31.67 //y=7.4 //x2=31.45 //y2=7.4
r670 (  302 402 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.385 //y=7.4 //x2=30.3 //y2=7.4
r671 (  301 403 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.91 //y=7.4 //x2=31.08 //y2=7.4
r672 (  301 302 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=30.91 //y=7.4 //x2=30.385 //y2=7.4
r673 (  295 402 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.3 //y=7.23 //x2=30.3 //y2=7.4
r674 (  295 431 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=30.3 //y=7.23 //x2=30.3 //y2=6.745
r675 (  292 401 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.505 //y=7.4 //x2=29.42 //y2=7.4
r676 (  292 294 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=29.505 //y=7.4 //x2=29.97 //y2=7.4
r677 (  291 402 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.215 //y=7.4 //x2=30.3 //y2=7.4
r678 (  291 294 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=30.215 //y=7.4 //x2=29.97 //y2=7.4
r679 (  285 401 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.42 //y=7.23 //x2=29.42 //y2=7.4
r680 (  285 430 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=29.42 //y=7.23 //x2=29.42 //y2=6.745
r681 (  282 400 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.625 //y=7.4 //x2=28.54 //y2=7.4
r682 (  282 284 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=28.625 //y=7.4 //x2=28.86 //y2=7.4
r683 (  281 401 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.335 //y=7.4 //x2=29.42 //y2=7.4
r684 (  281 284 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=29.335 //y=7.4 //x2=28.86 //y2=7.4
r685 (  275 400 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=28.54 //y=7.23 //x2=28.54 //y2=7.4
r686 (  275 429 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=28.54 //y=7.23 //x2=28.54 //y2=6.405
r687 (  274 399 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.92 //y=7.4 //x2=27.75 //y2=7.4
r688 (  273 400 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.455 //y=7.4 //x2=28.54 //y2=7.4
r689 (  273 274 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=28.455 //y=7.4 //x2=27.92 //y2=7.4
r690 (  268 398 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.17 //y=7.4 //x2=27.085 //y2=7.4
r691 (  268 270 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=27.17 //y=7.4 //x2=27.38 //y2=7.4
r692 (  267 399 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.58 //y=7.4 //x2=27.75 //y2=7.4
r693 (  267 270 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=27.58 //y=7.4 //x2=27.38 //y2=7.4
r694 (  261 398 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.085 //y=7.23 //x2=27.085 //y2=7.4
r695 (  261 428 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=27.085 //y=7.23 //x2=27.085 //y2=6.405
r696 (  260 397 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.29 //y=7.4 //x2=26.205 //y2=7.4
r697 (  259 398 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27 //y=7.4 //x2=27.085 //y2=7.4
r698 (  259 260 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=27 //y=7.4 //x2=26.29 //y2=7.4
r699 (  253 397 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.205 //y=7.23 //x2=26.205 //y2=7.4
r700 (  253 427 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=26.205 //y=7.23 //x2=26.205 //y2=6.405
r701 (  252 395 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.7 //y=7.4 //x2=25.53 //y2=7.4
r702 (  251 397 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.12 //y=7.4 //x2=26.205 //y2=7.4
r703 (  251 252 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=26.12 //y=7.4 //x2=25.7 //y2=7.4
r704 (  248 394 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.835 //y=7.4 //x2=24.75 //y2=7.4
r705 (  247 395 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.36 //y=7.4 //x2=25.53 //y2=7.4
r706 (  247 248 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=25.36 //y=7.4 //x2=24.835 //y2=7.4
r707 (  241 394 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.75 //y=7.23 //x2=24.75 //y2=7.4
r708 (  241 426 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=24.75 //y=7.23 //x2=24.75 //y2=6.745
r709 (  240 392 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.955 //y=7.4 //x2=23.87 //y2=7.4
r710 (  239 394 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.665 //y=7.4 //x2=24.75 //y2=7.4
r711 (  239 240 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=24.665 //y=7.4 //x2=23.955 //y2=7.4
r712 (  233 392 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.87 //y=7.23 //x2=23.87 //y2=7.4
r713 (  233 425 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=23.87 //y=7.23 //x2=23.87 //y2=6.745
r714 (  230 391 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.075 //y=7.4 //x2=22.99 //y2=7.4
r715 (  230 232 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=23.075 //y=7.4 //x2=23.68 //y2=7.4
r716 (  229 392 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.785 //y=7.4 //x2=23.87 //y2=7.4
r717 (  229 232 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=23.785 //y=7.4 //x2=23.68 //y2=7.4
r718 (  223 391 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.99 //y=7.23 //x2=22.99 //y2=7.4
r719 (  223 424 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=22.99 //y=7.23 //x2=22.99 //y2=6.405
r720 (  220 390 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.37 //y=7.4 //x2=22.2 //y2=7.4
r721 (  220 222 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=22.37 //y=7.4 //x2=22.57 //y2=7.4
r722 (  219 391 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.905 //y=7.4 //x2=22.99 //y2=7.4
r723 (  219 222 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=22.905 //y=7.4 //x2=22.57 //y2=7.4
r724 (  216 389 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.61 //y=7.4 //x2=21.525 //y2=7.4
r725 (  215 390 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.03 //y=7.4 //x2=22.2 //y2=7.4
r726 (  215 216 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=22.03 //y=7.4 //x2=21.61 //y2=7.4
r727 (  209 389 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.525 //y=7.23 //x2=21.525 //y2=7.4
r728 (  209 423 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=21.525 //y=7.23 //x2=21.525 //y2=6.405
r729 (  206 388 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.73 //y=7.4 //x2=20.645 //y2=7.4
r730 (  206 208 ) resistor r=12.9076 //w=0.357 //l=0.36 //layer=li \
 //thickness=0.1 //x=20.73 //y=7.4 //x2=21.09 //y2=7.4
r731 (  205 389 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.44 //y=7.4 //x2=21.525 //y2=7.4
r732 (  205 208 ) resistor r=12.549 //w=0.357 //l=0.35 //layer=li \
 //thickness=0.1 //x=21.44 //y=7.4 //x2=21.09 //y2=7.4
r733 (  199 388 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.645 //y=7.23 //x2=20.645 //y2=7.4
r734 (  199 422 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=20.645 //y=7.23 //x2=20.645 //y2=6.405
r735 (  198 387 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.15 //y=7.4 //x2=19.98 //y2=7.4
r736 (  197 388 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.56 //y=7.4 //x2=20.645 //y2=7.4
r737 (  197 198 ) resistor r=14.7003 //w=0.357 //l=0.41 //layer=li \
 //thickness=0.1 //x=20.56 //y=7.4 //x2=20.15 //y2=7.4
r738 (  192 194 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=18.5 //y=7.4 //x2=19.61 //y2=7.4
r739 (  190 386 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.965 //y=7.4 //x2=17.88 //y2=7.4
r740 (  190 192 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=17.965 //y=7.4 //x2=18.5 //y2=7.4
r741 (  189 387 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.81 //y=7.4 //x2=19.98 //y2=7.4
r742 (  189 194 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=19.81 //y=7.4 //x2=19.61 //y2=7.4
r743 (  185 386 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.88 //y=7.23 //x2=17.88 //y2=7.4
r744 (  185 421 ) resistor r=80.4278 //w=0.187 //l=1.175 //layer=li \
 //thickness=0.1 //x=17.88 //y=7.23 //x2=17.88 //y2=6.055
r745 (  182 385 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.82 //y=7.4 //x2=16.65 //y2=7.4
r746 (  182 184 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=16.82 //y=7.4 //x2=17.39 //y2=7.4
r747 (  181 386 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.795 //y=7.4 //x2=17.88 //y2=7.4
r748 (  181 184 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=17.795 //y=7.4 //x2=17.39 //y2=7.4
r749 (  176 178 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=14.8 //y=7.4 //x2=15.91 //y2=7.4
r750 (  174 384 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.635 //y=7.4 //x2=14.55 //y2=7.4
r751 (  174 176 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=14.635 //y=7.4 //x2=14.8 //y2=7.4
r752 (  173 385 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.48 //y=7.4 //x2=16.65 //y2=7.4
r753 (  173 178 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=16.48 //y=7.4 //x2=15.91 //y2=7.4
r754 (  169 384 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.55 //y=7.23 //x2=14.55 //y2=7.4
r755 (  169 420 ) resistor r=80.4278 //w=0.187 //l=1.175 //layer=li \
 //thickness=0.1 //x=14.55 //y=7.23 //x2=14.55 //y2=6.055
r756 (  166 383 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.49 //y=7.4 //x2=13.32 //y2=7.4
r757 (  166 168 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=13.49 //y=7.4 //x2=13.69 //y2=7.4
r758 (  165 384 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.465 //y=7.4 //x2=14.55 //y2=7.4
r759 (  165 168 ) resistor r=27.7871 //w=0.357 //l=0.775 //layer=li \
 //thickness=0.1 //x=14.465 //y=7.4 //x2=13.69 //y2=7.4
r760 (  162 382 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.74 //y=7.4 //x2=12.655 //y2=7.4
r761 (  161 383 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.15 //y=7.4 //x2=13.32 //y2=7.4
r762 (  161 162 ) resistor r=14.7003 //w=0.357 //l=0.41 //layer=li \
 //thickness=0.1 //x=13.15 //y=7.4 //x2=12.74 //y2=7.4
r763 (  155 382 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.655 //y=7.23 //x2=12.655 //y2=7.4
r764 (  155 419 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=12.655 //y=7.23 //x2=12.655 //y2=6.405
r765 (  152 381 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.86 //y=7.4 //x2=11.775 //y2=7.4
r766 (  152 154 ) resistor r=12.549 //w=0.357 //l=0.35 //layer=li \
 //thickness=0.1 //x=11.86 //y=7.4 //x2=12.21 //y2=7.4
r767 (  151 382 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.57 //y=7.4 //x2=12.655 //y2=7.4
r768 (  151 154 ) resistor r=12.9076 //w=0.357 //l=0.36 //layer=li \
 //thickness=0.1 //x=12.57 //y=7.4 //x2=12.21 //y2=7.4
r769 (  145 381 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.775 //y=7.23 //x2=11.775 //y2=7.4
r770 (  145 418 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=11.775 //y=7.23 //x2=11.775 //y2=6.405
r771 (  144 380 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.27 //y=7.4 //x2=11.1 //y2=7.4
r772 (  143 381 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.69 //y=7.4 //x2=11.775 //y2=7.4
r773 (  143 144 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=11.69 //y=7.4 //x2=11.27 //y2=7.4
r774 (  138 379 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.51 //y=7.4 //x2=10.425 //y2=7.4
r775 (  138 140 ) resistor r=7.88796 //w=0.357 //l=0.22 //layer=li \
 //thickness=0.1 //x=10.51 //y=7.4 //x2=10.73 //y2=7.4
r776 (  137 380 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.93 //y=7.4 //x2=11.1 //y2=7.4
r777 (  137 140 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=10.93 //y=7.4 //x2=10.73 //y2=7.4
r778 (  131 379 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.425 //y=7.23 //x2=10.425 //y2=7.4
r779 (  131 417 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=10.425 //y=7.23 //x2=10.425 //y2=6.405
r780 (  130 378 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.63 //y=7.4 //x2=9.545 //y2=7.4
r781 (  129 379 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.34 //y=7.4 //x2=10.425 //y2=7.4
r782 (  129 130 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.34 //y=7.4 //x2=9.63 //y2=7.4
r783 (  123 378 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.545 //y=7.23 //x2=9.545 //y2=7.4
r784 (  123 416 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=9.545 //y=7.23 //x2=9.545 //y2=6.405
r785 (  122 376 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.05 //y=7.4 //x2=8.88 //y2=7.4
r786 (  121 378 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.46 //y=7.4 //x2=9.545 //y2=7.4
r787 (  121 122 ) resistor r=14.7003 //w=0.357 //l=0.41 //layer=li \
 //thickness=0.1 //x=9.46 //y=7.4 //x2=9.05 //y2=7.4
r788 (  116 118 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=7.03 //y=7.4 //x2=8.14 //y2=7.4
r789 (  114 375 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.865 //y=7.4 //x2=6.78 //y2=7.4
r790 (  114 116 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=6.865 //y=7.4 //x2=7.03 //y2=7.4
r791 (  113 376 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.71 //y=7.4 //x2=8.88 //y2=7.4
r792 (  113 118 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=8.71 //y=7.4 //x2=8.14 //y2=7.4
r793 (  109 375 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=7.4
r794 (  109 415 ) resistor r=80.4278 //w=0.187 //l=1.175 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=6.055
r795 (  106 374 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.72 //y=7.4 //x2=5.55 //y2=7.4
r796 (  106 108 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=5.72 //y=7.4 //x2=5.92 //y2=7.4
r797 (  105 375 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.78 //y2=7.4
r798 (  105 108 ) resistor r=27.7871 //w=0.357 //l=0.775 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=5.92 //y2=7.4
r799 (  100 373 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.535 //y=7.4 //x2=3.45 //y2=7.4
r800 (  100 102 ) resistor r=32.4482 //w=0.357 //l=0.905 //layer=li \
 //thickness=0.1 //x=3.535 //y=7.4 //x2=4.44 //y2=7.4
r801 (  99 374 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.38 //y=7.4 //x2=5.55 //y2=7.4
r802 (  99 102 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=5.38 //y=7.4 //x2=4.44 //y2=7.4
r803 (  95 373 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.45 //y=7.23 //x2=3.45 //y2=7.4
r804 (  95 414 ) resistor r=80.4278 //w=0.187 //l=1.175 //layer=li \
 //thickness=0.1 //x=3.45 //y=7.23 //x2=3.45 //y2=6.055
r805 (  92 372 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.39 //y=7.4 //x2=2.22 //y2=7.4
r806 (  92 94 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=2.39 //y=7.4 //x2=3.33 //y2=7.4
r807 (  91 373 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.365 //y=7.4 //x2=3.45 //y2=7.4
r808 (  91 94 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=3.365 //y=7.4 //x2=3.33 //y2=7.4
r809 (  86 371 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.64 //y=7.4 //x2=1.555 //y2=7.4
r810 (  86 88 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=1.64 //y=7.4 //x2=1.85 //y2=7.4
r811 (  85 372 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.05 //y=7.4 //x2=2.22 //y2=7.4
r812 (  85 88 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=2.05 //y=7.4 //x2=1.85 //y2=7.4
r813 (  79 371 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=7.4
r814 (  79 413 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=6.405
r815 (  78 370 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.76 //y=7.4 //x2=0.675 //y2=7.4
r816 (  77 371 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=1.555 //y2=7.4
r817 (  77 78 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=0.76 //y2=7.4
r818 (  71 370 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=7.4
r819 (  71 412 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=6.405
r820 (  65 366 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=38.48 //y=7.4 //x2=38.48 //y2=7.4
r821 (  63 356 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37.74 //y=7.4 //x2=37.74 //y2=7.4
r822 (  63 65 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=37.74 //y=7.4 //x2=38.48 //y2=7.4
r823 (  61 342 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=36.26 //y=7.4 //x2=36.26 //y2=7.4
r824 (  61 63 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=36.26 //y=7.4 //x2=37.74 //y2=7.4
r825 (  59 340 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.15 //y=7.4 //x2=35.15 //y2=7.4
r826 (  59 61 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=35.15 //y=7.4 //x2=36.26 //y2=7.4
r827 (  57 330 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.04 //y=7.4 //x2=34.04 //y2=7.4
r828 (  57 59 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=34.04 //y=7.4 //x2=35.15 //y2=7.4
r829 (  55 406 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.56 //y=7.4 //x2=32.56 //y2=7.4
r830 (  55 57 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=32.56 //y=7.4 //x2=34.04 //y2=7.4
r831 (  53 308 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.45 //y=7.4 //x2=31.45 //y2=7.4
r832 (  53 55 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.45 //y=7.4 //x2=32.56 //y2=7.4
r833 (  51 294 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=29.97 //y=7.4 //x2=29.97 //y2=7.4
r834 (  51 53 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=29.97 //y=7.4 //x2=31.45 //y2=7.4
r835 (  49 284 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.86 //y=7.4 //x2=28.86 //y2=7.4
r836 (  49 51 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=28.86 //y=7.4 //x2=29.97 //y2=7.4
r837 (  47 270 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.38 //y=7.4 //x2=27.38 //y2=7.4
r838 (  47 49 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=27.38 //y=7.4 //x2=28.86 //y2=7.4
r839 (  45 397 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=26.27 //y=7.4 //x2=26.27 //y2=7.4
r840 (  45 47 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=26.27 //y=7.4 //x2=27.38 //y2=7.4
r841 (  43 394 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=7.4 //x2=24.79 //y2=7.4
r842 (  43 45 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=7.4 //x2=26.27 //y2=7.4
r843 (  41 232 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=7.4 //x2=23.68 //y2=7.4
r844 (  41 43 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=23.68 //y=7.4 //x2=24.79 //y2=7.4
r845 (  39 222 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.57 //y=7.4 //x2=22.57 //y2=7.4
r846 (  39 41 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.57 //y=7.4 //x2=23.68 //y2=7.4
r847 (  37 208 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=7.4 //x2=21.09 //y2=7.4
r848 (  37 39 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=7.4 //x2=22.57 //y2=7.4
r849 (  35 194 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.61 //y=7.4 //x2=19.61 //y2=7.4
r850 (  35 37 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=19.61 //y=7.4 //x2=21.09 //y2=7.4
r851 (  32 192 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=7.4 //x2=18.5 //y2=7.4
r852 (  30 184 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=7.4 //x2=17.39 //y2=7.4
r853 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=7.4 //x2=18.5 //y2=7.4
r854 (  28 178 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.91 //y=7.4 //x2=15.91 //y2=7.4
r855 (  28 30 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=15.91 //y=7.4 //x2=17.39 //y2=7.4
r856 (  26 176 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.8 //y=7.4 //x2=14.8 //y2=7.4
r857 (  26 28 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.8 //y=7.4 //x2=15.91 //y2=7.4
r858 (  24 168 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=7.4 //x2=13.69 //y2=7.4
r859 (  24 26 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=13.69 //y=7.4 //x2=14.8 //y2=7.4
r860 (  22 154 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.21 //y=7.4 //x2=12.21 //y2=7.4
r861 (  22 24 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.21 //y=7.4 //x2=13.69 //y2=7.4
r862 (  20 140 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.73 //y=7.4 //x2=10.73 //y2=7.4
r863 (  20 22 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=7.4 //x2=12.21 //y2=7.4
r864 (  18 378 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.62 //y=7.4 //x2=9.62 //y2=7.4
r865 (  18 20 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.62 //y=7.4 //x2=10.73 //y2=7.4
r866 (  16 118 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.14 //y=7.4 //x2=8.14 //y2=7.4
r867 (  16 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.14 //y=7.4 //x2=9.62 //y2=7.4
r868 (  14 116 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=7.4 //x2=7.03 //y2=7.4
r869 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=7.4 //x2=8.14 //y2=7.4
r870 (  12 108 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.92 //y=7.4 //x2=5.92 //y2=7.4
r871 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.92 //y=7.4 //x2=7.03 //y2=7.4
r872 (  10 102 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r873 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.92 //y2=7.4
r874 (  8 94 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=3.33 //y=7.4 //x2=3.33 //y2=7.4
r875 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=7.4 //x2=4.44 //y2=7.4
r876 (  6 88 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r877 (  6 8 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=3.33 //y2=7.4
r878 (  3 370 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r879 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r880 (  1 35 ) resistor r=0.0768272 //w=0.301 //l=0.185 //layer=m1 \
 //thickness=0.36 //x=19.425 //y=7.4 //x2=19.61 //y2=7.4
r881 (  1 32 ) resistor r=0.384136 //w=0.301 //l=0.925 //layer=m1 \
 //thickness=0.36 //x=19.425 //y=7.4 //x2=18.5 //y2=7.4
ends PM_FA\%VDD

subckt PM_FA\%A ( 1 2 4 5 6 8 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 \
 33 34 36 59 73 74 75 76 77 78 79 80 81 82 83 84 85 89 90 91 93 99 100 101 102 \
 103 104 108 110 113 114 118 119 120 125 127 129 135 136 138 152 156 157 160 )
c377 ( 160 0 ) capacitor c=0.0347334f //x=29.63 //y=4.7
c378 ( 157 0 ) capacitor c=0.0273722f //x=29.6 //y=1.915
c379 ( 156 0 ) capacitor c=0.0405821f //x=29.6 //y=2.08
c380 ( 152 0 ) capacitor c=0.0661295f //x=3.33 //y=4.7
c381 ( 138 0 ) capacitor c=0.0537799f //x=0.74 //y=2.085
c382 ( 136 0 ) capacitor c=0.0429696f //x=30.165 //y=1.25
c383 ( 135 0 ) capacitor c=0.0192208f //x=30.165 //y=0.905
c384 ( 129 0 ) capacitor c=0.0158629f //x=30.01 //y=1.405
c385 ( 127 0 ) capacitor c=0.0157803f //x=30.01 //y=0.75
c386 ( 125 0 ) capacitor c=0.0367015f //x=30.005 //y=4.79
c387 ( 120 0 ) capacitor c=0.0205163f //x=29.635 //y=1.56
c388 ( 119 0 ) capacitor c=0.0168481f //x=29.635 //y=1.25
c389 ( 118 0 ) capacitor c=0.0174142f //x=29.635 //y=0.905
c390 ( 114 0 ) capacitor c=0.0318948f //x=3.665 //y=1.215
c391 ( 113 0 ) capacitor c=0.0186029f //x=3.665 //y=0.87
c392 ( 110 0 ) capacitor c=0.0141798f //x=3.51 //y=1.37
c393 ( 108 0 ) capacitor c=0.0149852f //x=3.51 //y=0.715
c394 ( 104 0 ) capacitor c=0.0809667f //x=3.135 //y=1.92
c395 ( 103 0 ) capacitor c=0.0229153f //x=3.135 //y=1.525
c396 ( 102 0 ) capacitor c=0.0234352f //x=3.135 //y=1.215
c397 ( 101 0 ) capacitor c=0.0197989f //x=3.135 //y=0.87
c398 ( 100 0 ) capacitor c=0.0435629f //x=1.38 //y=1.255
c399 ( 99 0 ) capacitor c=0.0200386f //x=1.38 //y=0.91
c400 ( 93 0 ) capacitor c=0.0152946f //x=1.225 //y=1.41
c401 ( 91 0 ) capacitor c=0.0157804f //x=1.225 //y=0.755
c402 ( 90 0 ) capacitor c=0.048995f //x=0.97 //y=4.79
c403 ( 89 0 ) capacitor c=0.0303096f //x=1.26 //y=4.79
c404 ( 85 0 ) capacitor c=0.0290017f //x=0.85 //y=1.92
c405 ( 84 0 ) capacitor c=0.0250027f //x=0.85 //y=1.565
c406 ( 83 0 ) capacitor c=0.0234316f //x=0.85 //y=1.255
c407 ( 82 0 ) capacitor c=0.0200596f //x=0.85 //y=0.91
c408 ( 81 0 ) capacitor c=0.15358f //x=30.08 //y=6.02
c409 ( 80 0 ) capacitor c=0.110184f //x=29.64 //y=6.02
c410 ( 79 0 ) capacitor c=0.110797f //x=3.67 //y=6.02
c411 ( 78 0 ) capacitor c=0.154322f //x=3.23 //y=6.02
c412 ( 77 0 ) capacitor c=0.154218f //x=1.335 //y=6.02
c413 ( 76 0 ) capacitor c=0.154243f //x=0.895 //y=6.02
c414 ( 59 0 ) capacitor c=0.00415003f //x=29.6 //y=4.535
c415 ( 36 0 ) capacitor c=0.110862f //x=0.74 //y=2.085
c416 ( 34 0 ) capacitor c=0.00913498f //x=29.6 //y=2.22
c417 ( 33 0 ) capacitor c=0.0103502f //x=3.33 //y=2.22
c418 ( 28 0 ) capacitor c=0.0719211f //x=29.6 //y=2.59
c419 ( 23 0 ) capacitor c=0.101802f //x=3.33 //y=2.96
c420 ( 8 0 ) capacitor c=0.0133532f //x=29.6 //y=2.105
c421 ( 6 0 ) capacitor c=0.0050701f //x=3.415 //y=1.85
c422 ( 5 0 ) capacitor c=0.487085f //x=29.515 //y=1.85
c423 ( 4 0 ) capacitor c=0.0229105f //x=3.33 //y=2.105
c424 ( 2 0 ) capacitor c=0.0144527f //x=0.855 //y=4.07
c425 ( 1 0 ) capacitor c=0.0967174f //x=3.215 //y=4.07
r426 (  162 163 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=29.63 //y=4.79 //x2=29.63 //y2=4.865
r427 (  160 162 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=29.63 //y=4.7 //x2=29.63 //y2=4.79
r428 (  156 157 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=29.6 //y=2.08 //x2=29.6 //y2=1.915
r429 (  150 152 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=3.23 //y=4.7 //x2=3.33 //y2=4.7
r430 (  138 139 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=0.74 //y=2.085 //x2=0.85 //y2=2.085
r431 (  136 167 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.165 //y=1.25 //x2=30.125 //y2=1.405
r432 (  135 166 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.165 //y=0.905 //x2=30.125 //y2=0.75
r433 (  135 136 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=30.165 //y=0.905 //x2=30.165 //y2=1.25
r434 (  130 165 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.79 //y=1.405 //x2=29.675 //y2=1.405
r435 (  129 167 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.01 //y=1.405 //x2=30.125 //y2=1.405
r436 (  128 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.79 //y=0.75 //x2=29.675 //y2=0.75
r437 (  127 166 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=30.01 //y=0.75 //x2=30.125 //y2=0.75
r438 (  127 128 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=30.01 //y=0.75 //x2=29.79 //y2=0.75
r439 (  126 162 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=29.765 //y=4.79 //x2=29.63 //y2=4.79
r440 (  125 132 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=30.005 //y=4.79 //x2=30.08 //y2=4.865
r441 (  125 126 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=30.005 //y=4.79 //x2=29.765 //y2=4.79
r442 (  120 165 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.635 //y=1.56 //x2=29.675 //y2=1.405
r443 (  120 157 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=29.635 //y=1.56 //x2=29.635 //y2=1.915
r444 (  119 165 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.635 //y=1.25 //x2=29.675 //y2=1.405
r445 (  118 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.635 //y=0.905 //x2=29.675 //y2=0.75
r446 (  118 119 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=29.635 //y=0.905 //x2=29.635 //y2=1.25
r447 (  115 152 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=3.67 //y=4.865 //x2=3.33 //y2=4.7
r448 (  114 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.665 //y=1.215 //x2=3.625 //y2=1.37
r449 (  113 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.665 //y=0.87 //x2=3.625 //y2=0.715
r450 (  113 114 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.665 //y=0.87 //x2=3.665 //y2=1.215
r451 (  111 149 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.29 //y=1.37 //x2=3.175 //y2=1.37
r452 (  110 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.51 //y=1.37 //x2=3.625 //y2=1.37
r453 (  109 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.29 //y=0.715 //x2=3.175 //y2=0.715
r454 (  108 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.51 //y=0.715 //x2=3.625 //y2=0.715
r455 (  108 109 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.51 //y=0.715 //x2=3.29 //y2=0.715
r456 (  105 150 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.23 //y=4.865 //x2=3.23 //y2=4.7
r457 (  104 147 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.92 //x2=3.33 //y2=2.085
r458 (  103 149 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.525 //x2=3.175 //y2=1.37
r459 (  103 104 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.525 //x2=3.135 //y2=1.92
r460 (  102 149 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.135 //y=1.215 //x2=3.175 //y2=1.37
r461 (  101 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.135 //y=0.87 //x2=3.175 //y2=0.715
r462 (  101 102 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.135 //y=0.87 //x2=3.135 //y2=1.215
r463 (  100 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=1.255 //x2=1.34 //y2=1.41
r464 (  99 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.34 //y2=0.755
r465 (  99 100 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.38 //y2=1.255
r466 (  94 143 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=1.41 //x2=0.89 //y2=1.41
r467 (  93 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=1.41 //x2=1.34 //y2=1.41
r468 (  92 142 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=0.755 //x2=0.89 //y2=0.755
r469 (  91 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.34 //y2=0.755
r470 (  91 92 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.005 //y2=0.755
r471 (  89 96 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=1.335 //y2=4.865
r472 (  89 90 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=0.97 //y2=4.79
r473 (  86 90 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.97 //y2=4.79
r474 (  86 141 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.74 //y2=4.7
r475 (  85 139 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.92 //x2=0.85 //y2=2.085
r476 (  84 143 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.89 //y2=1.41
r477 (  84 85 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.85 //y2=1.92
r478 (  83 143 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.255 //x2=0.89 //y2=1.41
r479 (  82 142 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.89 //y2=0.755
r480 (  82 83 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.85 //y2=1.255
r481 (  81 132 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=30.08 //y=6.02 //x2=30.08 //y2=4.865
r482 (  80 163 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=29.64 //y=6.02 //x2=29.64 //y2=4.865
r483 (  79 115 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.67 //y=6.02 //x2=3.67 //y2=4.865
r484 (  78 105 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.23 //y=6.02 //x2=3.23 //y2=4.865
r485 (  77 96 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.335 //y=6.02 //x2=1.335 //y2=4.865
r486 (  76 86 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=0.895 //y=6.02 //x2=0.895 //y2=4.865
r487 (  75 129 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=29.9 //y=1.405 //x2=30.01 //y2=1.405
r488 (  75 130 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=29.9 //y=1.405 //x2=29.79 //y2=1.405
r489 (  74 110 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.4 //y=1.37 //x2=3.51 //y2=1.37
r490 (  74 111 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.4 //y=1.37 //x2=3.29 //y2=1.37
r491 (  73 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.225 //y2=1.41
r492 (  73 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.005 //y2=1.41
r493 (  69 160 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=29.63 //y=4.7 //x2=29.63 //y2=4.7
r494 (  59 69 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=29.6 //y=4.535 //x2=29.615 //y2=4.7
r495 (  56 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r496 (  46 141 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=4.7 //x2=0.74 //y2=4.7
r497 (  36 138 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=2.085 //x2=0.74 //y2=2.085
r498 (  34 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=29.6 //y=2.08 //x2=29.6 //y2=2.08
r499 (  34 58 ) resistor r=3.9234 //w=0.284 //l=0.195 //layer=li \
 //thickness=0.1 //x=29.6 //y=2.11 //x2=29.6 //y2=2.305
r500 (  33 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.085 //x2=3.33 //y2=2.085
r501 (  33 48 ) resistor r=3.85819 //w=0.281 //l=0.193 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.112 //x2=3.33 //y2=2.305
r502 (  32 59 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=29.6 //y=4.44 //x2=29.6 //y2=4.535
r503 (  31 32 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=29.6 //y=4.07 //x2=29.6 //y2=4.44
r504 (  30 31 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=29.6 //y=3.7 //x2=29.6 //y2=4.07
r505 (  29 30 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=29.6 //y=3.33 //x2=29.6 //y2=3.7
r506 (  28 29 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=29.6 //y=2.59 //x2=29.6 //y2=3.33
r507 (  28 58 ) resistor r=19.508 //w=0.187 //l=0.285 //layer=li \
 //thickness=0.1 //x=29.6 //y=2.59 //x2=29.6 //y2=2.305
r508 (  27 56 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=3.33 //y=4.44 //x2=3.33 //y2=4.7
r509 (  26 27 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=4.07 //x2=3.33 //y2=4.44
r510 (  25 26 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=3.7 //x2=3.33 //y2=4.07
r511 (  24 25 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=3.33 //x2=3.33 //y2=3.7
r512 (  23 24 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.96 //x2=3.33 //y2=3.33
r513 (  23 48 ) resistor r=44.8342 //w=0.187 //l=0.655 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.96 //x2=3.33 //y2=2.305
r514 (  22 46 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=0.74 //y=4.44 //x2=0.74 //y2=4.7
r515 (  21 22 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=4.07 //x2=0.74 //y2=4.44
r516 (  20 21 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=3.7 //x2=0.74 //y2=4.07
r517 (  19 20 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=3.33 //x2=0.74 //y2=3.7
r518 (  18 19 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=2.96 //x2=0.74 //y2=3.33
r519 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=2.59 //x2=0.74 //y2=2.96
r520 (  17 36 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=0.74 //y=2.59 //x2=0.74 //y2=2.085
r521 (  16 34 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=29.6 //y=2.22 //x2=29.6 //y2=2.22
r522 (  14 26 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=4.07 //x2=3.33 //y2=4.07
r523 (  12 33 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=2.22 //x2=3.33 //y2=2.22
r524 (  10 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=0.74 //y=4.07 //x2=0.74 //y2=4.07
r525 (  8 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=29.6 //y=2.105 //x2=29.6 //y2=2.22
r526 (  7 8 ) resistor r=0.162214 //w=0.131 //l=0.17 //layer=m1 \
 //thickness=0.36 //x=29.6 //y=1.935 //x2=29.6 //y2=2.105
r527 (  5 7 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=29.515 //y=1.85 //x2=29.6 //y2=1.935
r528 (  5 6 ) resistor r=24.9046 //w=0.131 //l=26.1 //layer=m1 \
 //thickness=0.36 //x=29.515 //y=1.85 //x2=3.415 //y2=1.85
r529 (  4 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=2.105 //x2=3.33 //y2=2.22
r530 (  3 6 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=1.935 //x2=3.415 //y2=1.85
r531 (  3 4 ) resistor r=0.162214 //w=0.131 //l=0.17 //layer=m1 \
 //thickness=0.36 //x=3.33 //y=1.935 //x2=3.33 //y2=2.105
r532 (  2 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=0.855 //y=4.07 //x2=0.74 //y2=4.07
r533 (  1 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.215 //y=4.07 //x2=3.33 //y2=4.07
r534 (  1 2 ) resistor r=2.25191 //w=0.131 //l=2.36 //layer=m1 \
 //thickness=0.36 //x=3.215 //y=4.07 //x2=0.855 //y2=4.07
ends PM_FA\%A

subckt PM_FA\%noxref_4 ( 1 2 17 18 19 20 24 26 33 34 35 36 37 38 39 43 45 51 \
 52 60 62 64 )
c161 ( 64 0 ) capacitor c=0.0288629f //x=0.97 //y=5.02
c162 ( 62 0 ) capacitor c=0.0170302f //x=0.925 //y=0.91
c163 ( 60 0 ) capacitor c=0.058481f //x=7.77 //y=4.7
c164 ( 52 0 ) capacitor c=0.0417768f //x=7.965 //y=1.255
c165 ( 51 0 ) capacitor c=0.01899f //x=7.965 //y=0.91
c166 ( 45 0 ) capacitor c=0.0124204f //x=7.81 //y=1.41
c167 ( 43 0 ) capacitor c=0.0157803f //x=7.81 //y=0.755
c168 ( 39 0 ) capacitor c=0.0889632f //x=7.435 //y=1.92
c169 ( 38 0 ) capacitor c=0.0194674f //x=7.435 //y=1.565
c170 ( 37 0 ) capacitor c=0.0168481f //x=7.435 //y=1.255
c171 ( 36 0 ) capacitor c=0.0173364f //x=7.435 //y=0.91
c172 ( 35 0 ) capacitor c=0.153255f //x=7.88 //y=6.02
c173 ( 34 0 ) capacitor c=0.110227f //x=7.44 //y=6.02
c174 ( 26 0 ) capacitor c=0.0735823f //x=7.77 //y=2.085
c175 ( 24 0 ) capacitor c=0.0865771f //x=1.48 //y=2.59
c176 ( 20 0 ) capacitor c=0.00417404f //x=1.2 //y=4.58
c177 ( 19 0 ) capacitor c=0.0118896f //x=1.395 //y=4.58
c178 ( 18 0 ) capacitor c=0.00621372f //x=1.195 //y=2.08
c179 ( 17 0 ) capacitor c=0.0132255f //x=1.395 //y=2.08
c180 ( 2 0 ) capacitor c=0.0163395f //x=1.595 //y=2.59
c181 ( 1 0 ) capacitor c=0.155274f //x=7.655 //y=2.59
r182 (  60 61 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.77 //y=4.7 //x2=7.88 //y2=4.7
r183 (  52 58 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.965 //y=1.255 //x2=7.925 //y2=1.41
r184 (  51 57 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.965 //y=0.91 //x2=7.925 //y2=0.755
r185 (  51 52 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.965 //y=0.91 //x2=7.965 //y2=1.255
r186 (  48 61 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=7.88 //y=4.865 //x2=7.88 //y2=4.7
r187 (  46 54 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.59 //y=1.41 //x2=7.475 //y2=1.41
r188 (  45 58 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.81 //y=1.41 //x2=7.925 //y2=1.41
r189 (  44 53 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.59 //y=0.755 //x2=7.475 //y2=0.755
r190 (  43 57 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.81 //y=0.755 //x2=7.925 //y2=0.755
r191 (  43 44 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.81 //y=0.755 //x2=7.59 //y2=0.755
r192 (  40 60 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=7.44 //y=4.865 //x2=7.77 //y2=4.7
r193 (  39 56 ) resistor r=67.2792 //w=0.24 //l=0.438891 //layer=ply \
 //thickness=0.18 //x=7.435 //y=1.92 //x2=7.77 //y2=2.16
r194 (  38 54 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.435 //y=1.565 //x2=7.475 //y2=1.41
r195 (  38 39 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=7.435 //y=1.565 //x2=7.435 //y2=1.92
r196 (  37 54 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.435 //y=1.255 //x2=7.475 //y2=1.41
r197 (  36 53 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.435 //y=0.91 //x2=7.475 //y2=0.755
r198 (  36 37 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.435 //y=0.91 //x2=7.435 //y2=1.255
r199 (  35 48 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.88 //y=6.02 //x2=7.88 //y2=4.865
r200 (  34 40 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.44 //y=6.02 //x2=7.44 //y2=4.865
r201 (  33 45 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.7 //y=1.41 //x2=7.81 //y2=1.41
r202 (  33 46 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.7 //y=1.41 //x2=7.59 //y2=1.41
r203 (  31 60 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.77 //y=4.7 //x2=7.77 //y2=4.7
r204 (  29 31 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=7.77 //y=2.59 //x2=7.77 //y2=4.7
r205 (  26 56 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.77 //y=2.085 //x2=7.77 //y2=2.085
r206 (  26 29 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=7.77 //y=2.085 //x2=7.77 //y2=2.59
r207 (  22 24 ) resistor r=130.396 //w=0.187 //l=1.905 //layer=li \
 //thickness=0.1 //x=1.48 //y=4.495 //x2=1.48 //y2=2.59
r208 (  21 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.48 //y=2.165 //x2=1.48 //y2=2.59
r209 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.48 //y2=4.495
r210 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.2 //y2=4.58
r211 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.48 //y2=2.165
r212 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.195 //y2=2.08
r213 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.2 //y2=4.58
r214 (  11 64 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.115 //y2=5.725
r215 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.195 //y2=2.08
r216 (  7 62 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.11 //y2=1.005
r217 (  6 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.77 //y=2.59 //x2=7.77 //y2=2.59
r218 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.48 //y=2.59 //x2=1.48 //y2=2.59
r219 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.595 //y=2.59 //x2=1.48 //y2=2.59
r220 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.655 //y=2.59 //x2=7.77 //y2=2.59
r221 (  1 2 ) resistor r=5.78244 //w=0.131 //l=6.06 //layer=m1 \
 //thickness=0.36 //x=7.655 //y=2.59 //x2=1.595 //y2=2.59
ends PM_FA\%noxref_4

subckt PM_FA\%noxref_5 ( 1 2 3 4 14 20 28 31 32 33 34 45 46 47 54 55 56 57 58 \
 60 63 64 66 74 76 )
c175 ( 76 0 ) capacitor c=0.0284262f //x=9.84 //y=5.02
c176 ( 74 0 ) capacitor c=0.0170943f //x=9.795 //y=0.91
c177 ( 66 0 ) capacitor c=0.0636249f //x=4.44 //y=4.7
c178 ( 64 0 ) capacitor c=0.0318948f //x=6.995 //y=1.215
c179 ( 63 0 ) capacitor c=0.0186029f //x=6.995 //y=0.87
c180 ( 60 0 ) capacitor c=0.0141798f //x=6.84 //y=1.37
c181 ( 58 0 ) capacitor c=0.0149852f //x=6.84 //y=0.715
c182 ( 57 0 ) capacitor c=0.0827875f //x=6.465 //y=1.92
c183 ( 56 0 ) capacitor c=0.0229212f //x=6.465 //y=1.525
c184 ( 55 0 ) capacitor c=0.0234352f //x=6.465 //y=1.215
c185 ( 54 0 ) capacitor c=0.0197989f //x=6.465 //y=0.87
c186 ( 47 0 ) capacitor c=0.153255f //x=4.55 //y=6.02
c187 ( 46 0 ) capacitor c=0.110227f //x=4.11 //y=6.02
c188 ( 34 0 ) capacitor c=0.00670488f //x=9.705 //y=4.58
c189 ( 33 0 ) capacitor c=0.0136086f //x=9.9 //y=4.58
c190 ( 32 0 ) capacitor c=0.00507261f //x=9.705 //y=2.08
c191 ( 31 0 ) capacitor c=0.0124351f //x=9.905 //y=2.08
c192 ( 28 0 ) capacitor c=0.0754874f //x=9.62 //y=3.33
c193 ( 20 0 ) capacitor c=0.0548742f //x=6.66 //y=2.085
c194 ( 14 0 ) capacitor c=0.024985f //x=4.44 //y=4.07
c195 ( 4 0 ) capacitor c=0.0126928f //x=6.775 //y=3.33
c196 ( 3 0 ) capacitor c=0.0521532f //x=9.505 //y=3.33
c197 ( 2 0 ) capacitor c=0.01091f //x=4.555 //y=4.07
c198 ( 1 0 ) capacitor c=0.10314f //x=9.505 //y=4.07
r199 (  66 67 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.44 //y=4.7 //x2=4.55 //y2=4.7
r200 (  64 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.995 //y=1.215 //x2=6.955 //y2=1.37
r201 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.995 //y=0.87 //x2=6.955 //y2=0.715
r202 (  63 64 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.995 //y=0.87 //x2=6.995 //y2=1.215
r203 (  61 71 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.62 //y=1.37 //x2=6.505 //y2=1.37
r204 (  60 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.84 //y=1.37 //x2=6.955 //y2=1.37
r205 (  59 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.62 //y=0.715 //x2=6.505 //y2=0.715
r206 (  58 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.84 //y=0.715 //x2=6.955 //y2=0.715
r207 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=6.84 //y=0.715 //x2=6.62 //y2=0.715
r208 (  57 69 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=6.465 //y=1.92 //x2=6.66 //y2=2.085
r209 (  56 71 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.465 //y=1.525 //x2=6.505 //y2=1.37
r210 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=6.465 //y=1.525 //x2=6.465 //y2=1.92
r211 (  55 71 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.465 //y=1.215 //x2=6.505 //y2=1.37
r212 (  54 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.465 //y=0.87 //x2=6.505 //y2=0.715
r213 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.465 //y=0.87 //x2=6.465 //y2=1.215
r214 (  51 67 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=4.55 //y=4.865 //x2=4.55 //y2=4.7
r215 (  48 66 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=4.11 //y=4.865 //x2=4.44 //y2=4.7
r216 (  47 51 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.55 //y=6.02 //x2=4.55 //y2=4.865
r217 (  46 48 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.11 //y=6.02 //x2=4.11 //y2=4.865
r218 (  45 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.73 //y=1.37 //x2=6.84 //y2=1.37
r219 (  45 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.73 //y=1.37 //x2=6.62 //y2=1.37
r220 (  41 74 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=9.99 //y=1.995 //x2=9.99 //y2=1.005
r221 (  35 76 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=9.985 //y=4.665 //x2=9.985 //y2=5.725
r222 (  33 35 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.9 //y=4.58 //x2=9.985 //y2=4.665
r223 (  33 34 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=9.9 //y=4.58 //x2=9.705 //y2=4.58
r224 (  31 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.905 //y=2.08 //x2=9.99 //y2=1.995
r225 (  31 32 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=9.905 //y=2.08 //x2=9.705 //y2=2.08
r226 (  28 30 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=9.62 //y=3.33 //x2=9.62 //y2=4.07
r227 (  26 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.62 //y=4.495 //x2=9.705 //y2=4.58
r228 (  26 30 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=9.62 //y=4.495 //x2=9.62 //y2=4.07
r229 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.62 //y=2.165 //x2=9.705 //y2=2.08
r230 (  25 28 ) resistor r=79.7433 //w=0.187 //l=1.165 //layer=li \
 //thickness=0.1 //x=9.62 //y=2.165 //x2=9.62 //y2=3.33
r231 (  20 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=2.085 //x2=6.66 //y2=2.085
r232 (  20 23 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=6.66 //y=2.085 //x2=6.66 //y2=3.33
r233 (  17 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=4.7 //x2=4.44 //y2=4.7
r234 (  14 17 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=4.44 //y=4.07 //x2=4.44 //y2=4.7
r235 (  12 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.62 //y=4.07 //x2=9.62 //y2=4.07
r236 (  10 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.62 //y=3.33 //x2=9.62 //y2=3.33
r237 (  8 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.66 //y=3.33 //x2=6.66 //y2=3.33
r238 (  6 14 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.44 //y=4.07 //x2=4.44 //y2=4.07
r239 (  4 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.775 //y=3.33 //x2=6.66 //y2=3.33
r240 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.505 //y=3.33 //x2=9.62 //y2=3.33
r241 (  3 4 ) resistor r=2.60496 //w=0.131 //l=2.73 //layer=m1 \
 //thickness=0.36 //x=9.505 //y=3.33 //x2=6.775 //y2=3.33
r242 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.555 //y=4.07 //x2=4.44 //y2=4.07
r243 (  1 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.505 //y=4.07 //x2=9.62 //y2=4.07
r244 (  1 2 ) resistor r=4.72328 //w=0.131 //l=4.95 //layer=m1 \
 //thickness=0.36 //x=9.505 //y=4.07 //x2=4.555 //y2=4.07
ends PM_FA\%noxref_5

subckt PM_FA\%B ( 1 2 3 4 5 6 18 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 \
 36 49 65 75 76 77 78 79 80 81 82 83 84 85 86 87 88 90 93 94 101 102 106 107 \
 108 110 113 116 117 118 119 120 121 122 123 127 129 132 133 145 150 161 )
c381 ( 161 0 ) capacitor c=0.0627475f //x=28.86 //y=4.7
c382 ( 150 0 ) capacitor c=0.0513056f //x=10.25 //y=2.085
c383 ( 145 0 ) capacitor c=0.0606915f //x=6.66 //y=4.7
c384 ( 133 0 ) capacitor c=0.0318948f //x=29.195 //y=1.21
c385 ( 132 0 ) capacitor c=0.0187384f //x=29.195 //y=0.865
c386 ( 129 0 ) capacitor c=0.0141798f //x=29.04 //y=1.365
c387 ( 127 0 ) capacitor c=0.0149844f //x=29.04 //y=0.71
c388 ( 123 0 ) capacitor c=0.0811005f //x=28.665 //y=1.915
c389 ( 122 0 ) capacitor c=0.0229212f //x=28.665 //y=1.52
c390 ( 121 0 ) capacitor c=0.0234352f //x=28.665 //y=1.21
c391 ( 120 0 ) capacitor c=0.0199343f //x=28.665 //y=0.865
c392 ( 119 0 ) capacitor c=0.0293214f //x=10.25 //y=1.92
c393 ( 118 0 ) capacitor c=0.0250171f //x=10.25 //y=1.565
c394 ( 117 0 ) capacitor c=0.0234316f //x=10.25 //y=1.255
c395 ( 116 0 ) capacitor c=0.0199789f //x=10.25 //y=0.91
c396 ( 113 0 ) capacitor c=0.0488408f //x=10.205 //y=4.865
c397 ( 110 0 ) capacitor c=0.0148979f //x=10.095 //y=1.41
c398 ( 108 0 ) capacitor c=0.0157804f //x=10.095 //y=0.755
c399 ( 107 0 ) capacitor c=0.0129718f //x=9.84 //y=4.79
c400 ( 106 0 ) capacitor c=0.0172687f //x=10.13 //y=4.79
c401 ( 102 0 ) capacitor c=0.0435512f //x=9.72 //y=1.255
c402 ( 101 0 ) capacitor c=0.0199346f //x=9.72 //y=0.91
c403 ( 94 0 ) capacitor c=0.0417768f //x=4.635 //y=1.255
c404 ( 93 0 ) capacitor c=0.01899f //x=4.635 //y=0.91
c405 ( 90 0 ) capacitor c=0.0124204f //x=4.48 //y=1.41
c406 ( 88 0 ) capacitor c=0.0157803f //x=4.48 //y=0.755
c407 ( 87 0 ) capacitor c=0.0889343f //x=4.105 //y=1.92
c408 ( 86 0 ) capacitor c=0.0194674f //x=4.105 //y=1.565
c409 ( 85 0 ) capacitor c=0.0168481f //x=4.105 //y=1.255
c410 ( 84 0 ) capacitor c=0.0173364f //x=4.105 //y=0.91
c411 ( 83 0 ) capacitor c=0.110274f //x=29.2 //y=6.02
c412 ( 82 0 ) capacitor c=0.154186f //x=28.76 //y=6.02
c413 ( 81 0 ) capacitor c=0.1536f //x=10.205 //y=6.02
c414 ( 80 0 ) capacitor c=0.154218f //x=9.765 //y=6.02
c415 ( 79 0 ) capacitor c=0.110797f //x=7 //y=6.02
c416 ( 78 0 ) capacitor c=0.154322f //x=6.56 //y=6.02
c417 ( 65 0 ) capacitor c=0.0938005f //x=28.86 //y=2.08
c418 ( 49 0 ) capacitor c=0.0850502f //x=10.36 //y=2.085
c419 ( 36 0 ) capacitor c=0.029964f //x=4.44 //y=2.085
c420 ( 34 0 ) capacitor c=0.00995663f //x=28.86 //y=4.81
c421 ( 22 0 ) capacitor c=0.0150587f //x=6.66 //y=4.44
c422 ( 18 0 ) capacitor c=0.0148475f //x=28.86 //y=4.63
c423 ( 6 0 ) capacitor c=0.0111878f //x=10.475 //y=4.81
c424 ( 5 0 ) capacitor c=0.430557f //x=28.745 //y=4.81
c425 ( 4 0 ) capacitor c=0.015004f //x=6.775 //y=4.44
c426 ( 3 0 ) capacitor c=0.0883217f //x=10.245 //y=4.44
c427 ( 2 0 ) capacitor c=0.0154186f //x=4.555 //y=2.96
c428 ( 1 0 ) capacitor c=0.113504f //x=10.245 //y=2.96
r429 (  159 161 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=28.76 //y=4.7 //x2=28.86 //y2=4.7
r430 (  150 152 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.25 //y=2.085 //x2=10.36 //y2=2.085
r431 (  143 145 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=6.56 //y=4.7 //x2=6.66 //y2=4.7
r432 (  134 161 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=29.2 //y=4.865 //x2=28.86 //y2=4.7
r433 (  133 163 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.195 //y=1.21 //x2=29.155 //y2=1.365
r434 (  132 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.195 //y=0.865 //x2=29.155 //y2=0.71
r435 (  132 133 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=29.195 //y=0.865 //x2=29.195 //y2=1.21
r436 (  130 158 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.82 //y=1.365 //x2=28.705 //y2=1.365
r437 (  129 163 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.04 //y=1.365 //x2=29.155 //y2=1.365
r438 (  128 157 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.82 //y=0.71 //x2=28.705 //y2=0.71
r439 (  127 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.04 //y=0.71 //x2=29.155 //y2=0.71
r440 (  127 128 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=29.04 //y=0.71 //x2=28.82 //y2=0.71
r441 (  124 159 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=28.76 //y=4.865 //x2=28.76 //y2=4.7
r442 (  123 156 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=28.665 //y=1.915 //x2=28.86 //y2=2.08
r443 (  122 158 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.665 //y=1.52 //x2=28.705 //y2=1.365
r444 (  122 123 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=28.665 //y=1.52 //x2=28.665 //y2=1.915
r445 (  121 158 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.665 //y=1.21 //x2=28.705 //y2=1.365
r446 (  120 157 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.665 //y=0.865 //x2=28.705 //y2=0.71
r447 (  120 121 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=28.665 //y=0.865 //x2=28.665 //y2=1.21
r448 (  119 150 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=10.25 //y=1.92 //x2=10.25 //y2=2.085
r449 (  118 149 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.25 //y=1.565 //x2=10.21 //y2=1.41
r450 (  118 119 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=10.25 //y=1.565 //x2=10.25 //y2=1.92
r451 (  117 149 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.25 //y=1.255 //x2=10.21 //y2=1.41
r452 (  116 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.25 //y=0.91 //x2=10.21 //y2=0.755
r453 (  116 117 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.25 //y=0.91 //x2=10.25 //y2=1.255
r454 (  113 154 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=10.205 //y=4.865 //x2=10.36 //y2=4.7
r455 (  111 147 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.875 //y=1.41 //x2=9.76 //y2=1.41
r456 (  110 149 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.095 //y=1.41 //x2=10.21 //y2=1.41
r457 (  109 146 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.875 //y=0.755 //x2=9.76 //y2=0.755
r458 (  108 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.095 //y=0.755 //x2=10.21 //y2=0.755
r459 (  108 109 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.095 //y=0.755 //x2=9.875 //y2=0.755
r460 (  106 113 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.13 //y=4.79 //x2=10.205 //y2=4.865
r461 (  106 107 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=10.13 //y=4.79 //x2=9.84 //y2=4.79
r462 (  103 107 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=9.765 //y=4.865 //x2=9.84 //y2=4.79
r463 (  102 147 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.72 //y=1.255 //x2=9.76 //y2=1.41
r464 (  101 146 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.72 //y=0.91 //x2=9.76 //y2=0.755
r465 (  101 102 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.72 //y=0.91 //x2=9.72 //y2=1.255
r466 (  98 145 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=7 //y=4.865 //x2=6.66 //y2=4.7
r467 (  95 143 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.56 //y=4.865 //x2=6.56 //y2=4.7
r468 (  94 142 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.635 //y=1.255 //x2=4.595 //y2=1.41
r469 (  93 141 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.635 //y=0.91 //x2=4.595 //y2=0.755
r470 (  93 94 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.635 //y=0.91 //x2=4.635 //y2=1.255
r471 (  91 138 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.26 //y=1.41 //x2=4.145 //y2=1.41
r472 (  90 142 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.48 //y=1.41 //x2=4.595 //y2=1.41
r473 (  89 137 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.26 //y=0.755 //x2=4.145 //y2=0.755
r474 (  88 141 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.48 //y=0.755 //x2=4.595 //y2=0.755
r475 (  88 89 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.48 //y=0.755 //x2=4.26 //y2=0.755
r476 (  87 140 ) resistor r=67.2792 //w=0.24 //l=0.438891 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.92 //x2=4.44 //y2=2.16
r477 (  86 138 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.565 //x2=4.145 //y2=1.41
r478 (  86 87 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.565 //x2=4.105 //y2=1.92
r479 (  85 138 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.105 //y=1.255 //x2=4.145 //y2=1.41
r480 (  84 137 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.105 //y=0.91 //x2=4.145 //y2=0.755
r481 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.105 //y=0.91 //x2=4.105 //y2=1.255
r482 (  83 134 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=29.2 //y=6.02 //x2=29.2 //y2=4.865
r483 (  82 124 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=28.76 //y=6.02 //x2=28.76 //y2=4.865
r484 (  81 113 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.205 //y=6.02 //x2=10.205 //y2=4.865
r485 (  80 103 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.765 //y=6.02 //x2=9.765 //y2=4.865
r486 (  79 98 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7 //y=6.02 //x2=7 //y2=4.865
r487 (  78 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.56 //y=6.02 //x2=6.56 //y2=4.865
r488 (  77 129 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=28.93 //y=1.365 //x2=29.04 //y2=1.365
r489 (  77 130 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=28.93 //y=1.365 //x2=28.82 //y2=1.365
r490 (  76 110 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.985 //y=1.41 //x2=10.095 //y2=1.41
r491 (  76 111 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.985 //y=1.41 //x2=9.875 //y2=1.41
r492 (  75 90 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.37 //y=1.41 //x2=4.48 //y2=1.41
r493 (  75 91 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.37 //y=1.41 //x2=4.26 //y2=1.41
r494 (  65 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=28.86 //y=2.08 //x2=28.86 //y2=2.08
r495 (  59 154 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.36 //y=4.7 //x2=10.36 //y2=4.7
r496 (  49 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.36 //y=2.085 //x2=10.36 //y2=2.085
r497 (  46 145 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=4.7 //x2=6.66 //y2=4.7
r498 (  36 140 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=2.085 //x2=4.44 //y2=2.085
r499 (  34 161 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=28.86 //y=4.7 //x2=28.86 //y2=4.7
r500 (  34 63 ) resistor r=3.4525 //w=0.263 //l=0.175 //layer=li \
 //thickness=0.1 //x=28.86 //y=4.72 //x2=28.86 //y2=4.545
r501 (  33 63 ) resistor r=7.18717 //w=0.187 //l=0.105 //layer=li \
 //thickness=0.1 //x=28.86 //y=4.44 //x2=28.86 //y2=4.545
r502 (  32 33 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=28.86 //y=4.07 //x2=28.86 //y2=4.44
r503 (  31 32 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=28.86 //y=3.7 //x2=28.86 //y2=4.07
r504 (  30 31 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=28.86 //y=3.33 //x2=28.86 //y2=3.7
r505 (  29 30 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=28.86 //y=2.59 //x2=28.86 //y2=3.33
r506 (  29 65 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=28.86 //y=2.59 //x2=28.86 //y2=2.08
r507 (  28 59 ) resistor r=7.52941 //w=0.187 //l=0.11 //layer=li \
 //thickness=0.1 //x=10.36 //y=4.81 //x2=10.36 //y2=4.7
r508 (  27 59 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=10.36 //y=4.44 //x2=10.36 //y2=4.7
r509 (  26 27 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=10.36 //y=4.07 //x2=10.36 //y2=4.44
r510 (  25 26 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=10.36 //y=3.33 //x2=10.36 //y2=4.07
r511 (  24 25 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.96 //x2=10.36 //y2=3.33
r512 (  23 24 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.59 //x2=10.36 //y2=2.96
r513 (  23 49 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.59 //x2=10.36 //y2=2.085
r514 (  22 46 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=6.66 //y=4.44 //x2=6.66 //y2=4.7
r515 (  20 21 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.22 //x2=4.44 //y2=2.96
r516 (  20 36 ) resistor r=9.24064 //w=0.187 //l=0.135 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.22 //x2=4.44 //y2=2.085
r517 (  18 34 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=28.86 //y=4.63 //x2=28.86 //y2=4.63
r518 (  18 19 ) resistor r=0.104651 //w=0.215 //l=0.18 //layer=m1 \
 //thickness=0.36 //x=28.86 //y=4.63 //x2=28.86 //y2=4.81
r519 (  16 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.36 //y=4.44 //x2=10.36 //y2=4.44
r520 (  14 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.36 //y=2.96 //x2=10.36 //y2=2.96
r521 (  12 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.36 //y=4.81 //x2=10.36 //y2=4.81
r522 (  10 22 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.66 //y=4.44 //x2=6.66 //y2=4.44
r523 (  8 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.44 //y=2.96 //x2=4.44 //y2=2.96
r524 (  6 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.475 //y=4.81 //x2=10.36 //y2=4.81
r525 (  5 19 ) resistor r=0.0216707 //w=0.215 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=28.745 //y=4.81 //x2=28.86 //y2=4.81
r526 (  5 6 ) resistor r=17.4332 //w=0.131 //l=18.27 //layer=m1 \
 //thickness=0.36 //x=28.745 //y=4.81 //x2=10.475 //y2=4.81
r527 (  4 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.775 //y=4.44 //x2=6.66 //y2=4.44
r528 (  3 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.245 //y=4.44 //x2=10.36 //y2=4.44
r529 (  3 4 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=10.245 //y=4.44 //x2=6.775 //y2=4.44
r530 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.555 //y=2.96 //x2=4.44 //y2=2.96
r531 (  1 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.245 //y=2.96 //x2=10.36 //y2=2.96
r532 (  1 2 ) resistor r=5.42939 //w=0.131 //l=5.69 //layer=m1 \
 //thickness=0.36 //x=10.245 //y=2.96 //x2=4.555 //y2=2.96
ends PM_FA\%B

subckt PM_FA\%noxref_7 ( 1 2 3 4 5 6 7 8 33 34 35 36 40 51 52 53 54 58 60 72 \
 79 81 87 88 89 90 91 92 93 94 95 96 97 98 99 103 104 105 107 113 114 115 116 \
 117 118 122 124 127 128 132 133 134 139 141 143 149 150 152 166 170 171 174 \
 182 183 186 187 )
c420 ( 187 0 ) capacitor c=0.0159588f //x=7.515 //y=5.02
c421 ( 186 0 ) capacitor c=0.0159588f //x=4.185 //y=5.02
c422 ( 183 0 ) capacitor c=0.00827922f //x=7.51 //y=0.91
c423 ( 182 0 ) capacitor c=0.00846882f //x=4.18 //y=0.91
c424 ( 174 0 ) capacitor c=0.0347773f //x=24.08 //y=4.7
c425 ( 171 0 ) capacitor c=0.0270331f //x=24.05 //y=1.915
c426 ( 170 0 ) capacitor c=0.0423789f //x=24.05 //y=2.08
c427 ( 166 0 ) capacitor c=0.06601f //x=14.43 //y=4.7
c428 ( 152 0 ) capacitor c=0.0505038f //x=11.84 //y=2.085
c429 ( 150 0 ) capacitor c=0.0429696f //x=24.615 //y=1.25
c430 ( 149 0 ) capacitor c=0.0190738f //x=24.615 //y=0.905
c431 ( 143 0 ) capacitor c=0.0148572f //x=24.46 //y=1.405
c432 ( 141 0 ) capacitor c=0.0157803f //x=24.46 //y=0.75
c433 ( 139 0 ) capacitor c=0.037277f //x=24.455 //y=4.79
c434 ( 134 0 ) capacitor c=0.0205163f //x=24.085 //y=1.56
c435 ( 133 0 ) capacitor c=0.0168481f //x=24.085 //y=1.25
c436 ( 132 0 ) capacitor c=0.0174142f //x=24.085 //y=0.905
c437 ( 128 0 ) capacitor c=0.0318948f //x=14.765 //y=1.215
c438 ( 127 0 ) capacitor c=0.0186029f //x=14.765 //y=0.87
c439 ( 124 0 ) capacitor c=0.0141798f //x=14.61 //y=1.37
c440 ( 122 0 ) capacitor c=0.0149852f //x=14.61 //y=0.715
c441 ( 118 0 ) capacitor c=0.0823795f //x=14.235 //y=1.92
c442 ( 117 0 ) capacitor c=0.0229212f //x=14.235 //y=1.525
c443 ( 116 0 ) capacitor c=0.0234352f //x=14.235 //y=1.215
c444 ( 115 0 ) capacitor c=0.0197989f //x=14.235 //y=0.87
c445 ( 114 0 ) capacitor c=0.0435629f //x=12.48 //y=1.255
c446 ( 113 0 ) capacitor c=0.0199463f //x=12.48 //y=0.91
c447 ( 107 0 ) capacitor c=0.0148979f //x=12.325 //y=1.41
c448 ( 105 0 ) capacitor c=0.0157804f //x=12.325 //y=0.755
c449 ( 104 0 ) capacitor c=0.049215f //x=12.07 //y=4.79
c450 ( 103 0 ) capacitor c=0.030248f //x=12.36 //y=4.79
c451 ( 99 0 ) capacitor c=0.0293214f //x=11.95 //y=1.92
c452 ( 98 0 ) capacitor c=0.0250027f //x=11.95 //y=1.565
c453 ( 97 0 ) capacitor c=0.0234316f //x=11.95 //y=1.255
c454 ( 96 0 ) capacitor c=0.0199673f //x=11.95 //y=0.91
c455 ( 95 0 ) capacitor c=0.15358f //x=24.53 //y=6.02
c456 ( 94 0 ) capacitor c=0.110117f //x=24.09 //y=6.02
c457 ( 93 0 ) capacitor c=0.110632f //x=14.77 //y=6.02
c458 ( 92 0 ) capacitor c=0.154209f //x=14.33 //y=6.02
c459 ( 91 0 ) capacitor c=0.154131f //x=12.435 //y=6.02
c460 ( 90 0 ) capacitor c=0.154154f //x=11.995 //y=6.02
c461 ( 81 0 ) capacitor c=0.0762812f //x=24.05 //y=2.08
c462 ( 79 0 ) capacitor c=0.00307329f //x=24.05 //y=4.535
c463 ( 72 0 ) capacitor c=0.104556f //x=14.43 //y=2.085
c464 ( 60 0 ) capacitor c=0.0826372f //x=11.84 //y=2.085
c465 ( 58 0 ) capacitor c=0.0885032f //x=8.14 //y=3.7
c466 ( 54 0 ) capacitor c=0.0016874f //x=7.785 //y=1.655
c467 ( 53 0 ) capacitor c=0.014358f //x=8.055 //y=1.655
c468 ( 52 0 ) capacitor c=0.00235465f //x=7.745 //y=5.205
c469 ( 51 0 ) capacitor c=0.0121398f //x=8.055 //y=5.205
c470 ( 40 0 ) capacitor c=0.104613f //x=4.81 //y=3.7
c471 ( 36 0 ) capacitor c=0.0016874f //x=4.455 //y=1.655
c472 ( 35 0 ) capacitor c=0.014358f //x=4.725 //y=1.655
c473 ( 34 0 ) capacitor c=0.0027221f //x=4.415 //y=5.205
c474 ( 33 0 ) capacitor c=0.0121701f //x=4.725 //y=5.205
c475 ( 8 0 ) capacitor c=0.00719749f //x=11.955 //y=4.07
c476 ( 7 0 ) capacitor c=0.0689485f //x=14.315 //y=4.07
c477 ( 6 0 ) capacitor c=0.0140175f //x=11.955 //y=2.22
c478 ( 5 0 ) capacitor c=0.201199f //x=23.935 //y=2.22
c479 ( 4 0 ) capacitor c=0.00275131f //x=8.255 //y=3.7
c480 ( 3 0 ) capacitor c=0.0880917f //x=11.725 //y=3.7
c481 ( 2 0 ) capacitor c=0.0134265f //x=4.925 //y=3.7
c482 ( 1 0 ) capacitor c=0.0544718f //x=8.025 //y=3.7
r483 (  176 177 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=24.08 //y=4.79 //x2=24.08 //y2=4.865
r484 (  174 176 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=24.08 //y=4.7 //x2=24.08 //y2=4.79
r485 (  170 171 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=24.05 //y=2.08 //x2=24.05 //y2=1.915
r486 (  164 166 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=14.33 //y=4.7 //x2=14.43 //y2=4.7
r487 (  152 153 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.84 //y=2.085 //x2=11.95 //y2=2.085
r488 (  150 181 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.615 //y=1.25 //x2=24.575 //y2=1.405
r489 (  149 180 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.615 //y=0.905 //x2=24.575 //y2=0.75
r490 (  149 150 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.615 //y=0.905 //x2=24.615 //y2=1.25
r491 (  144 179 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.24 //y=1.405 //x2=24.125 //y2=1.405
r492 (  143 181 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.46 //y=1.405 //x2=24.575 //y2=1.405
r493 (  142 178 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.24 //y=0.75 //x2=24.125 //y2=0.75
r494 (  141 180 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.46 //y=0.75 //x2=24.575 //y2=0.75
r495 (  141 142 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=24.46 //y=0.75 //x2=24.24 //y2=0.75
r496 (  140 176 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=24.215 //y=4.79 //x2=24.08 //y2=4.79
r497 (  139 146 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=24.455 //y=4.79 //x2=24.53 //y2=4.865
r498 (  139 140 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=24.455 //y=4.79 //x2=24.215 //y2=4.79
r499 (  134 179 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.085 //y=1.56 //x2=24.125 //y2=1.405
r500 (  134 171 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=24.085 //y=1.56 //x2=24.085 //y2=1.915
r501 (  133 179 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.085 //y=1.25 //x2=24.125 //y2=1.405
r502 (  132 178 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.085 //y=0.905 //x2=24.125 //y2=0.75
r503 (  132 133 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.085 //y=0.905 //x2=24.085 //y2=1.25
r504 (  129 166 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=14.77 //y=4.865 //x2=14.43 //y2=4.7
r505 (  128 168 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.765 //y=1.215 //x2=14.725 //y2=1.37
r506 (  127 167 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.765 //y=0.87 //x2=14.725 //y2=0.715
r507 (  127 128 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.765 //y=0.87 //x2=14.765 //y2=1.215
r508 (  125 163 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.39 //y=1.37 //x2=14.275 //y2=1.37
r509 (  124 168 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.61 //y=1.37 //x2=14.725 //y2=1.37
r510 (  123 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.39 //y=0.715 //x2=14.275 //y2=0.715
r511 (  122 167 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.61 //y=0.715 //x2=14.725 //y2=0.715
r512 (  122 123 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=14.61 //y=0.715 //x2=14.39 //y2=0.715
r513 (  119 164 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=14.33 //y=4.865 //x2=14.33 //y2=4.7
r514 (  118 161 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=14.235 //y=1.92 //x2=14.43 //y2=2.085
r515 (  117 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.235 //y=1.525 //x2=14.275 //y2=1.37
r516 (  117 118 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=14.235 //y=1.525 //x2=14.235 //y2=1.92
r517 (  116 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.235 //y=1.215 //x2=14.275 //y2=1.37
r518 (  115 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.235 //y=0.87 //x2=14.275 //y2=0.715
r519 (  115 116 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.235 //y=0.87 //x2=14.235 //y2=1.215
r520 (  114 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.48 //y=1.255 //x2=12.44 //y2=1.41
r521 (  113 158 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.48 //y=0.91 //x2=12.44 //y2=0.755
r522 (  113 114 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.48 //y=0.91 //x2=12.48 //y2=1.255
r523 (  108 157 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.105 //y=1.41 //x2=11.99 //y2=1.41
r524 (  107 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.325 //y=1.41 //x2=12.44 //y2=1.41
r525 (  106 156 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.105 //y=0.755 //x2=11.99 //y2=0.755
r526 (  105 158 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=12.325 //y=0.755 //x2=12.44 //y2=0.755
r527 (  105 106 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=12.325 //y=0.755 //x2=12.105 //y2=0.755
r528 (  103 110 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=12.36 //y=4.79 //x2=12.435 //y2=4.865
r529 (  103 104 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=12.36 //y=4.79 //x2=12.07 //y2=4.79
r530 (  100 104 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=11.995 //y=4.865 //x2=12.07 //y2=4.79
r531 (  100 155 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=11.995 //y=4.865 //x2=11.84 //y2=4.7
r532 (  99 153 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=11.95 //y=1.92 //x2=11.95 //y2=2.085
r533 (  98 157 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.95 //y=1.565 //x2=11.99 //y2=1.41
r534 (  98 99 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=11.95 //y=1.565 //x2=11.95 //y2=1.92
r535 (  97 157 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.95 //y=1.255 //x2=11.99 //y2=1.41
r536 (  96 156 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.95 //y=0.91 //x2=11.99 //y2=0.755
r537 (  96 97 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.95 //y=0.91 //x2=11.95 //y2=1.255
r538 (  95 146 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=24.53 //y=6.02 //x2=24.53 //y2=4.865
r539 (  94 177 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=24.09 //y=6.02 //x2=24.09 //y2=4.865
r540 (  93 129 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.77 //y=6.02 //x2=14.77 //y2=4.865
r541 (  92 119 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.33 //y=6.02 //x2=14.33 //y2=4.865
r542 (  91 110 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.435 //y=6.02 //x2=12.435 //y2=4.865
r543 (  90 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.995 //y=6.02 //x2=11.995 //y2=4.865
r544 (  89 143 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=24.35 //y=1.405 //x2=24.46 //y2=1.405
r545 (  89 144 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=24.35 //y=1.405 //x2=24.24 //y2=1.405
r546 (  88 124 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.5 //y=1.37 //x2=14.61 //y2=1.37
r547 (  88 125 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.5 //y=1.37 //x2=14.39 //y2=1.37
r548 (  87 107 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.215 //y=1.41 //x2=12.325 //y2=1.41
r549 (  87 108 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=12.215 //y=1.41 //x2=12.105 //y2=1.41
r550 (  86 174 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=24.08 //y=4.7 //x2=24.08 //y2=4.7
r551 (  81 170 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=24.05 //y=2.08 //x2=24.05 //y2=2.08
r552 (  81 84 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=24.05 //y=2.08 //x2=24.05 //y2=2.22
r553 (  79 86 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=24.05 //y=4.535 //x2=24.065 //y2=4.7
r554 (  79 84 ) resistor r=158.46 //w=0.187 //l=2.315 //layer=li \
 //thickness=0.1 //x=24.05 //y=4.535 //x2=24.05 //y2=2.22
r555 (  77 166 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.43 //y=4.7 //x2=14.43 //y2=4.7
r556 (  75 77 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=14.43 //y=4.07 //x2=14.43 //y2=4.7
r557 (  72 161 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.43 //y=2.085 //x2=14.43 //y2=2.085
r558 (  72 75 ) resistor r=135.872 //w=0.187 //l=1.985 //layer=li \
 //thickness=0.1 //x=14.43 //y=2.085 //x2=14.43 //y2=4.07
r559 (  69 155 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=4.7 //x2=11.84 //y2=4.7
r560 (  67 69 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=11.84 //y=4.07 //x2=11.84 //y2=4.7
r561 (  65 67 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=11.84 //y=3.7 //x2=11.84 //y2=4.07
r562 (  63 65 ) resistor r=101.305 //w=0.187 //l=1.48 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.22 //x2=11.84 //y2=3.7
r563 (  60 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=2.085 //x2=11.84 //y2=2.085
r564 (  60 63 ) resistor r=9.24064 //w=0.187 //l=0.135 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.085 //x2=11.84 //y2=2.22
r565 (  56 58 ) resistor r=97.1979 //w=0.187 //l=1.42 //layer=li \
 //thickness=0.1 //x=8.14 //y=5.12 //x2=8.14 //y2=3.7
r566 (  55 58 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=8.14 //y=1.74 //x2=8.14 //y2=3.7
r567 (  53 55 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.055 //y=1.655 //x2=8.14 //y2=1.74
r568 (  53 54 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=8.055 //y=1.655 //x2=7.785 //y2=1.655
r569 (  51 56 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.055 //y=5.205 //x2=8.14 //y2=5.12
r570 (  51 52 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=8.055 //y=5.205 //x2=7.745 //y2=5.205
r571 (  47 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.7 //y=1.57 //x2=7.785 //y2=1.655
r572 (  47 183 ) resistor r=38.6738 //w=0.187 //l=0.565 //layer=li \
 //thickness=0.1 //x=7.7 //y=1.57 //x2=7.7 //y2=1.005
r573 (  41 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.66 //y=5.29 //x2=7.745 //y2=5.205
r574 (  41 187 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=7.66 //y=5.29 //x2=7.66 //y2=5.715
r575 (  38 40 ) resistor r=97.1979 //w=0.187 //l=1.42 //layer=li \
 //thickness=0.1 //x=4.81 //y=5.12 //x2=4.81 //y2=3.7
r576 (  37 40 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=4.81 //y=1.74 //x2=4.81 //y2=3.7
r577 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=1.655 //x2=4.81 //y2=1.74
r578 (  35 36 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=4.725 //y=1.655 //x2=4.455 //y2=1.655
r579 (  33 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=5.205 //x2=4.81 //y2=5.12
r580 (  33 34 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=4.725 //y=5.205 //x2=4.415 //y2=5.205
r581 (  29 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.37 //y=1.57 //x2=4.455 //y2=1.655
r582 (  29 182 ) resistor r=38.6738 //w=0.187 //l=0.565 //layer=li \
 //thickness=0.1 //x=4.37 //y=1.57 //x2=4.37 //y2=1.005
r583 (  23 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.33 //y=5.29 //x2=4.415 //y2=5.205
r584 (  23 186 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=4.33 //y=5.29 //x2=4.33 //y2=5.715
r585 (  22 84 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=24.05 //y=2.22 //x2=24.05 //y2=2.22
r586 (  20 75 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.43 //y=4.07 //x2=14.43 //y2=4.07
r587 (  18 65 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.84 //y=3.7 //x2=11.84 //y2=3.7
r588 (  16 67 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.84 //y=4.07 //x2=11.84 //y2=4.07
r589 (  14 63 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.84 //y=2.22 //x2=11.84 //y2=2.22
r590 (  12 58 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.14 //y=3.7 //x2=8.14 //y2=3.7
r591 (  10 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.81 //y=3.7 //x2=4.81 //y2=3.7
r592 (  8 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.955 //y=4.07 //x2=11.84 //y2=4.07
r593 (  7 20 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=14.315 //y=4.07 //x2=14.43 //y2=4.07
r594 (  7 8 ) resistor r=2.25191 //w=0.131 //l=2.36 //layer=m1 \
 //thickness=0.36 //x=14.315 //y=4.07 //x2=11.955 //y2=4.07
r595 (  6 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.955 //y=2.22 //x2=11.84 //y2=2.22
r596 (  5 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.935 //y=2.22 //x2=24.05 //y2=2.22
r597 (  5 6 ) resistor r=11.4313 //w=0.131 //l=11.98 //layer=m1 \
 //thickness=0.36 //x=23.935 //y=2.22 //x2=11.955 //y2=2.22
r598 (  4 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.255 //y=3.7 //x2=8.14 //y2=3.7
r599 (  3 18 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.725 //y=3.7 //x2=11.84 //y2=3.7
r600 (  3 4 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=11.725 //y=3.7 //x2=8.255 //y2=3.7
r601 (  2 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.925 //y=3.7 //x2=4.81 //y2=3.7
r602 (  1 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.025 //y=3.7 //x2=8.14 //y2=3.7
r603 (  1 2 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=8.025 //y=3.7 //x2=4.925 //y2=3.7
ends PM_FA\%noxref_7

subckt PM_FA\%noxref_8 ( 1 2 17 18 19 20 24 26 33 34 35 36 37 38 39 43 45 51 \
 52 60 62 64 )
c163 ( 64 0 ) capacitor c=0.0280624f //x=12.07 //y=5.02
c164 ( 62 0 ) capacitor c=0.0170084f //x=12.025 //y=0.91
c165 ( 60 0 ) capacitor c=0.0588976f //x=18.87 //y=4.7
c166 ( 52 0 ) capacitor c=0.0417768f //x=19.065 //y=1.255
c167 ( 51 0 ) capacitor c=0.01899f //x=19.065 //y=0.91
c168 ( 45 0 ) capacitor c=0.0124204f //x=18.91 //y=1.41
c169 ( 43 0 ) capacitor c=0.0157803f //x=18.91 //y=0.755
c170 ( 39 0 ) capacitor c=0.0889138f //x=18.535 //y=1.92
c171 ( 38 0 ) capacitor c=0.0194674f //x=18.535 //y=1.565
c172 ( 37 0 ) capacitor c=0.0168481f //x=18.535 //y=1.255
c173 ( 36 0 ) capacitor c=0.0173364f //x=18.535 //y=0.91
c174 ( 35 0 ) capacitor c=0.153256f //x=18.98 //y=6.02
c175 ( 34 0 ) capacitor c=0.110062f //x=18.54 //y=6.02
c176 ( 26 0 ) capacitor c=0.0699117f //x=18.87 //y=2.085
c177 ( 24 0 ) capacitor c=0.0843781f //x=12.58 //y=2.59
c178 ( 20 0 ) capacitor c=0.00413007f //x=12.3 //y=4.58
c179 ( 19 0 ) capacitor c=0.0103938f //x=12.495 //y=4.58
c180 ( 18 0 ) capacitor c=0.00476658f //x=12.295 //y=2.08
c181 ( 17 0 ) capacitor c=0.0155174f //x=12.495 //y=2.08
c182 ( 2 0 ) capacitor c=0.0146857f //x=12.695 //y=2.59
c183 ( 1 0 ) capacitor c=0.121614f //x=18.755 //y=2.59
r184 (  60 61 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.87 //y=4.7 //x2=18.98 //y2=4.7
r185 (  52 58 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.065 //y=1.255 //x2=19.025 //y2=1.41
r186 (  51 57 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.065 //y=0.91 //x2=19.025 //y2=0.755
r187 (  51 52 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=19.065 //y=0.91 //x2=19.065 //y2=1.255
r188 (  48 61 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=18.98 //y=4.865 //x2=18.98 //y2=4.7
r189 (  46 54 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.69 //y=1.41 //x2=18.575 //y2=1.41
r190 (  45 58 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.91 //y=1.41 //x2=19.025 //y2=1.41
r191 (  44 53 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.69 //y=0.755 //x2=18.575 //y2=0.755
r192 (  43 57 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.91 //y=0.755 //x2=19.025 //y2=0.755
r193 (  43 44 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=18.91 //y=0.755 //x2=18.69 //y2=0.755
r194 (  40 60 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=18.54 //y=4.865 //x2=18.87 //y2=4.7
r195 (  39 56 ) resistor r=67.2792 //w=0.24 //l=0.438891 //layer=ply \
 //thickness=0.18 //x=18.535 //y=1.92 //x2=18.87 //y2=2.16
r196 (  38 54 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.535 //y=1.565 //x2=18.575 //y2=1.41
r197 (  38 39 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=18.535 //y=1.565 //x2=18.535 //y2=1.92
r198 (  37 54 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.535 //y=1.255 //x2=18.575 //y2=1.41
r199 (  36 53 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.535 //y=0.91 //x2=18.575 //y2=0.755
r200 (  36 37 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.535 //y=0.91 //x2=18.535 //y2=1.255
r201 (  35 48 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.98 //y=6.02 //x2=18.98 //y2=4.865
r202 (  34 40 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.54 //y=6.02 //x2=18.54 //y2=4.865
r203 (  33 45 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.8 //y=1.41 //x2=18.91 //y2=1.41
r204 (  33 46 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.8 //y=1.41 //x2=18.69 //y2=1.41
r205 (  31 60 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.87 //y=4.7 //x2=18.87 //y2=4.7
r206 (  29 31 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=18.87 //y=2.59 //x2=18.87 //y2=4.7
r207 (  26 56 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.87 //y=2.085 //x2=18.87 //y2=2.085
r208 (  26 29 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=18.87 //y=2.085 //x2=18.87 //y2=2.59
r209 (  22 24 ) resistor r=130.396 //w=0.187 //l=1.905 //layer=li \
 //thickness=0.1 //x=12.58 //y=4.495 //x2=12.58 //y2=2.59
r210 (  21 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=12.58 //y=2.165 //x2=12.58 //y2=2.59
r211 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.495 //y=4.58 //x2=12.58 //y2=4.495
r212 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=12.495 //y=4.58 //x2=12.3 //y2=4.58
r213 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.495 //y=2.08 //x2=12.58 //y2=2.165
r214 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.495 //y=2.08 //x2=12.295 //y2=2.08
r215 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.215 //y=4.665 //x2=12.3 //y2=4.58
r216 (  11 64 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=12.215 //y=4.665 //x2=12.215 //y2=5.725
r217 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.21 //y=1.995 //x2=12.295 //y2=2.08
r218 (  7 62 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=12.21 //y=1.995 //x2=12.21 //y2=1.005
r219 (  6 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.87 //y=2.59 //x2=18.87 //y2=2.59
r220 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.58 //y=2.59 //x2=12.58 //y2=2.59
r221 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.695 //y=2.59 //x2=12.58 //y2=2.59
r222 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.755 //y=2.59 //x2=18.87 //y2=2.59
r223 (  1 2 ) resistor r=5.78244 //w=0.131 //l=6.06 //layer=m1 \
 //thickness=0.36 //x=18.755 //y=2.59 //x2=12.695 //y2=2.59
ends PM_FA\%noxref_8

subckt PM_FA\%SUM ( 1 2 7 8 9 10 11 22 23 24 25 42 43 44 45 51 52 55 56 )
c148 ( 56 0 ) capacitor c=0.0159588f //x=18.615 //y=5.02
c149 ( 55 0 ) capacitor c=0.0159588f //x=15.285 //y=5.02
c150 ( 52 0 ) capacitor c=0.00827922f //x=18.61 //y=0.91
c151 ( 51 0 ) capacitor c=0.00846882f //x=15.28 //y=0.91
c152 ( 45 0 ) capacitor c=0.0016874f //x=18.885 //y=1.655
c153 ( 44 0 ) capacitor c=0.014358f //x=19.155 //y=1.655
c154 ( 43 0 ) capacitor c=0.00222879f //x=18.845 //y=5.205
c155 ( 42 0 ) capacitor c=0.011934f //x=19.155 //y=5.205
c156 ( 25 0 ) capacitor c=0.0016874f //x=15.555 //y=1.655
c157 ( 24 0 ) capacitor c=0.014358f //x=15.825 //y=1.655
c158 ( 23 0 ) capacitor c=0.00222879f //x=15.515 //y=5.205
c159 ( 22 0 ) capacitor c=0.0117456f //x=15.825 //y=5.205
c160 ( 10 0 ) capacitor c=0.0870285f //x=19.24 //y=2.59
c161 ( 7 0 ) capacitor c=0.103261f //x=15.91 //y=3.33
c162 ( 2 0 ) capacitor c=0.0103701f //x=16.025 //y=3.7
c163 ( 1 0 ) capacitor c=0.0661877f //x=19.125 //y=3.7
r164 (  44 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=19.155 //y=1.655 //x2=19.24 //y2=1.74
r165 (  44 45 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=19.155 //y=1.655 //x2=18.885 //y2=1.655
r166 (  42 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=19.155 //y=5.205 //x2=19.24 //y2=5.12
r167 (  42 43 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=19.155 //y=5.205 //x2=18.845 //y2=5.205
r168 (  38 45 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.8 //y=1.57 //x2=18.885 //y2=1.655
r169 (  38 52 ) resistor r=38.6738 //w=0.187 //l=0.565 //layer=li \
 //thickness=0.1 //x=18.8 //y=1.57 //x2=18.8 //y2=1.005
r170 (  32 43 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.76 //y=5.29 //x2=18.845 //y2=5.205
r171 (  32 56 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=18.76 //y=5.29 //x2=18.76 //y2=5.715
r172 (  24 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.825 //y=1.655 //x2=15.91 //y2=1.74
r173 (  24 25 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=15.825 //y=1.655 //x2=15.555 //y2=1.655
r174 (  22 27 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.825 //y=5.205 //x2=15.91 //y2=5.12
r175 (  22 23 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=15.825 //y=5.205 //x2=15.515 //y2=5.205
r176 (  18 25 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.47 //y=1.57 //x2=15.555 //y2=1.655
r177 (  18 51 ) resistor r=38.6738 //w=0.187 //l=0.565 //layer=li \
 //thickness=0.1 //x=15.47 //y=1.57 //x2=15.47 //y2=1.005
r178 (  12 23 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.43 //y=5.29 //x2=15.515 //y2=5.205
r179 (  12 55 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=15.43 //y=5.29 //x2=15.43 //y2=5.715
r180 (  11 47 ) resistor r=97.1979 //w=0.187 //l=1.42 //layer=li \
 //thickness=0.1 //x=19.24 //y=3.7 //x2=19.24 //y2=5.12
r181 (  10 11 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=19.24 //y=2.59 //x2=19.24 //y2=3.7
r182 (  10 46 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=19.24 //y=2.59 //x2=19.24 //y2=1.74
r183 (  9 27 ) resistor r=46.5455 //w=0.187 //l=0.68 //layer=li \
 //thickness=0.1 //x=15.91 //y=4.44 //x2=15.91 //y2=5.12
r184 (  8 9 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li //thickness=0.1 \
 //x=15.91 //y=3.7 //x2=15.91 //y2=4.44
r185 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=15.91 //y=3.33 //x2=15.91 //y2=3.7
r186 (  7 26 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=15.91 //y=3.33 //x2=15.91 //y2=1.74
r187 (  6 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=19.24 //y=3.7 //x2=19.24 //y2=3.7
r188 (  4 8 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.91 //y=3.7 //x2=15.91 //y2=3.7
r189 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.025 //y=3.7 //x2=15.91 //y2=3.7
r190 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=19.125 //y=3.7 //x2=19.24 //y2=3.7
r191 (  1 2 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=19.125 //y=3.7 //x2=16.025 //y2=3.7
ends PM_FA\%SUM

subckt PM_FA\%noxref_10 ( 1 2 3 4 14 20 28 31 32 33 34 45 46 47 54 55 56 57 58 \
 60 63 64 66 74 76 )
c172 ( 76 0 ) capacitor c=0.0279647f //x=20.94 //y=5.02
c173 ( 74 0 ) capacitor c=0.0170596f //x=20.895 //y=0.91
c174 ( 66 0 ) capacitor c=0.0640415f //x=15.54 //y=4.7
c175 ( 64 0 ) capacitor c=0.0318948f //x=18.095 //y=1.215
c176 ( 63 0 ) capacitor c=0.0186029f //x=18.095 //y=0.87
c177 ( 60 0 ) capacitor c=0.0141798f //x=17.94 //y=1.37
c178 ( 58 0 ) capacitor c=0.0149852f //x=17.94 //y=0.715
c179 ( 57 0 ) capacitor c=0.0823795f //x=17.565 //y=1.92
c180 ( 56 0 ) capacitor c=0.0229212f //x=17.565 //y=1.525
c181 ( 55 0 ) capacitor c=0.0234352f //x=17.565 //y=1.215
c182 ( 54 0 ) capacitor c=0.0197989f //x=17.565 //y=0.87
c183 ( 47 0 ) capacitor c=0.153256f //x=15.65 //y=6.02
c184 ( 46 0 ) capacitor c=0.110062f //x=15.21 //y=6.02
c185 ( 34 0 ) capacitor c=0.00614759f //x=20.805 //y=4.58
c186 ( 33 0 ) capacitor c=0.0137356f //x=21 //y=4.58
c187 ( 32 0 ) capacitor c=0.00618684f //x=20.805 //y=2.08
c188 ( 31 0 ) capacitor c=0.0139695f //x=21.005 //y=2.08
c189 ( 28 0 ) capacitor c=0.0765759f //x=20.72 //y=3.33
c190 ( 20 0 ) capacitor c=0.0523393f //x=17.76 //y=2.085
c191 ( 14 0 ) capacitor c=0.0234413f //x=15.54 //y=4.07
c192 ( 4 0 ) capacitor c=0.0126928f //x=17.875 //y=3.33
c193 ( 3 0 ) capacitor c=0.0515075f //x=20.605 //y=3.33
c194 ( 2 0 ) capacitor c=0.00869386f //x=15.655 //y=4.07
c195 ( 1 0 ) capacitor c=0.0895659f //x=20.605 //y=4.07
r196 (  66 67 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.54 //y=4.7 //x2=15.65 //y2=4.7
r197 (  64 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.095 //y=1.215 //x2=18.055 //y2=1.37
r198 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.095 //y=0.87 //x2=18.055 //y2=0.715
r199 (  63 64 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.095 //y=0.87 //x2=18.095 //y2=1.215
r200 (  61 71 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.72 //y=1.37 //x2=17.605 //y2=1.37
r201 (  60 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.94 //y=1.37 //x2=18.055 //y2=1.37
r202 (  59 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.72 //y=0.715 //x2=17.605 //y2=0.715
r203 (  58 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.94 //y=0.715 //x2=18.055 //y2=0.715
r204 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=17.94 //y=0.715 //x2=17.72 //y2=0.715
r205 (  57 69 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=17.565 //y=1.92 //x2=17.76 //y2=2.085
r206 (  56 71 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.565 //y=1.525 //x2=17.605 //y2=1.37
r207 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=17.565 //y=1.525 //x2=17.565 //y2=1.92
r208 (  55 71 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.565 //y=1.215 //x2=17.605 //y2=1.37
r209 (  54 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.565 //y=0.87 //x2=17.605 //y2=0.715
r210 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.565 //y=0.87 //x2=17.565 //y2=1.215
r211 (  51 67 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=15.65 //y=4.865 //x2=15.65 //y2=4.7
r212 (  48 66 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=15.21 //y=4.865 //x2=15.54 //y2=4.7
r213 (  47 51 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.65 //y=6.02 //x2=15.65 //y2=4.865
r214 (  46 48 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.21 //y=6.02 //x2=15.21 //y2=4.865
r215 (  45 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.83 //y=1.37 //x2=17.94 //y2=1.37
r216 (  45 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.83 //y=1.37 //x2=17.72 //y2=1.37
r217 (  41 74 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=21.09 //y=1.995 //x2=21.09 //y2=1.005
r218 (  35 76 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=21.085 //y=4.665 //x2=21.085 //y2=5.725
r219 (  33 35 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21 //y=4.58 //x2=21.085 //y2=4.665
r220 (  33 34 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=21 //y=4.58 //x2=20.805 //y2=4.58
r221 (  31 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.005 //y=2.08 //x2=21.09 //y2=1.995
r222 (  31 32 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=21.005 //y=2.08 //x2=20.805 //y2=2.08
r223 (  28 30 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=20.72 //y=3.33 //x2=20.72 //y2=4.07
r224 (  26 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.72 //y=4.495 //x2=20.805 //y2=4.58
r225 (  26 30 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=20.72 //y=4.495 //x2=20.72 //y2=4.07
r226 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.72 //y=2.165 //x2=20.805 //y2=2.08
r227 (  25 28 ) resistor r=79.7433 //w=0.187 //l=1.165 //layer=li \
 //thickness=0.1 //x=20.72 //y=2.165 //x2=20.72 //y2=3.33
r228 (  20 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.76 //y=2.085 //x2=17.76 //y2=2.085
r229 (  20 23 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.085 //x2=17.76 //y2=3.33
r230 (  17 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.54 //y=4.7 //x2=15.54 //y2=4.7
r231 (  14 17 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=15.54 //y=4.07 //x2=15.54 //y2=4.7
r232 (  12 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=20.72 //y=4.07 //x2=20.72 //y2=4.07
r233 (  10 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=20.72 //y=3.33 //x2=20.72 //y2=3.33
r234 (  8 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.76 //y=3.33 //x2=17.76 //y2=3.33
r235 (  6 14 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.54 //y=4.07 //x2=15.54 //y2=4.07
r236 (  4 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.875 //y=3.33 //x2=17.76 //y2=3.33
r237 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=3.33 //x2=20.72 //y2=3.33
r238 (  3 4 ) resistor r=2.60496 //w=0.131 //l=2.73 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=3.33 //x2=17.875 //y2=3.33
r239 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.655 //y=4.07 //x2=15.54 //y2=4.07
r240 (  1 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=4.07 //x2=20.72 //y2=4.07
r241 (  1 2 ) resistor r=4.72328 //w=0.131 //l=4.95 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=4.07 //x2=15.655 //y2=4.07
ends PM_FA\%noxref_10

subckt PM_FA\%CIN ( 1 2 3 4 5 6 17 18 19 20 21 22 23 24 25 26 27 28 29 30 32 \
 44 58 70 71 72 73 74 75 76 77 78 79 80 81 82 83 85 88 89 96 97 101 102 103 \
 105 108 111 112 113 114 115 116 117 118 122 124 127 128 140 145 156 )
c251 ( 156 0 ) capacitor c=0.064035f //x=23.31 //y=4.7
c252 ( 145 0 ) capacitor c=0.0503242f //x=21.35 //y=2.085
c253 ( 140 0 ) capacitor c=0.0605721f //x=17.76 //y=4.7
c254 ( 128 0 ) capacitor c=0.0318948f //x=23.645 //y=1.21
c255 ( 127 0 ) capacitor c=0.0187384f //x=23.645 //y=0.865
c256 ( 124 0 ) capacitor c=0.0141798f //x=23.49 //y=1.365
c257 ( 122 0 ) capacitor c=0.0149844f //x=23.49 //y=0.71
c258 ( 118 0 ) capacitor c=0.0804766f //x=23.115 //y=1.915
c259 ( 117 0 ) capacitor c=0.0229212f //x=23.115 //y=1.52
c260 ( 116 0 ) capacitor c=0.0234352f //x=23.115 //y=1.21
c261 ( 115 0 ) capacitor c=0.0199343f //x=23.115 //y=0.865
c262 ( 114 0 ) capacitor c=0.0293214f //x=21.35 //y=1.92
c263 ( 113 0 ) capacitor c=0.0250171f //x=21.35 //y=1.565
c264 ( 112 0 ) capacitor c=0.0234316f //x=21.35 //y=1.255
c265 ( 111 0 ) capacitor c=0.0199789f //x=21.35 //y=0.91
c266 ( 108 0 ) capacitor c=0.0490825f //x=21.305 //y=4.865
c267 ( 105 0 ) capacitor c=0.0148979f //x=21.195 //y=1.41
c268 ( 103 0 ) capacitor c=0.0157804f //x=21.195 //y=0.755
c269 ( 102 0 ) capacitor c=0.0129101f //x=20.94 //y=4.79
c270 ( 101 0 ) capacitor c=0.0173472f //x=21.23 //y=4.79
c271 ( 97 0 ) capacitor c=0.0435512f //x=20.82 //y=1.255
c272 ( 96 0 ) capacitor c=0.0199346f //x=20.82 //y=0.91
c273 ( 89 0 ) capacitor c=0.0417768f //x=15.735 //y=1.255
c274 ( 88 0 ) capacitor c=0.01899f //x=15.735 //y=0.91
c275 ( 85 0 ) capacitor c=0.0124204f //x=15.58 //y=1.41
c276 ( 83 0 ) capacitor c=0.0157803f //x=15.58 //y=0.755
c277 ( 82 0 ) capacitor c=0.0889138f //x=15.205 //y=1.92
c278 ( 81 0 ) capacitor c=0.0194674f //x=15.205 //y=1.565
c279 ( 80 0 ) capacitor c=0.0168481f //x=15.205 //y=1.255
c280 ( 79 0 ) capacitor c=0.0173364f //x=15.205 //y=0.91
c281 ( 78 0 ) capacitor c=0.11011f //x=23.65 //y=6.02
c282 ( 77 0 ) capacitor c=0.154192f //x=23.21 //y=6.02
c283 ( 76 0 ) capacitor c=0.154154f //x=21.305 //y=6.02
c284 ( 75 0 ) capacitor c=0.154131f //x=20.865 //y=6.02
c285 ( 74 0 ) capacitor c=0.110632f //x=18.1 //y=6.02
c286 ( 73 0 ) capacitor c=0.154209f //x=17.66 //y=6.02
c287 ( 58 0 ) capacitor c=0.0957711f //x=23.31 //y=2.08
c288 ( 44 0 ) capacitor c=0.0865219f //x=21.46 //y=2.085
c289 ( 32 0 ) capacitor c=0.0283262f //x=15.54 //y=2.085
c290 ( 18 0 ) capacitor c=0.0131564f //x=17.76 //y=4.44
c291 ( 6 0 ) capacitor c=0.0027479f //x=21.575 //y=4.44
c292 ( 5 0 ) capacitor c=0.0578447f //x=23.195 //y=4.44
c293 ( 4 0 ) capacitor c=0.0125654f //x=17.875 //y=4.44
c294 ( 3 0 ) capacitor c=0.0440536f //x=21.345 //y=4.44
c295 ( 2 0 ) capacitor c=0.0154186f //x=15.655 //y=2.96
c296 ( 1 0 ) capacitor c=0.110748f //x=21.345 //y=2.96
r297 (  154 156 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=23.21 //y=4.7 //x2=23.31 //y2=4.7
r298 (  145 147 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=21.35 //y=2.085 //x2=21.46 //y2=2.085
r299 (  138 140 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=17.66 //y=4.7 //x2=17.76 //y2=4.7
r300 (  129 156 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=23.65 //y=4.865 //x2=23.31 //y2=4.7
r301 (  128 158 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.645 //y=1.21 //x2=23.605 //y2=1.365
r302 (  127 157 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.645 //y=0.865 //x2=23.605 //y2=0.71
r303 (  127 128 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=23.645 //y=0.865 //x2=23.645 //y2=1.21
r304 (  125 153 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.27 //y=1.365 //x2=23.155 //y2=1.365
r305 (  124 158 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.49 //y=1.365 //x2=23.605 //y2=1.365
r306 (  123 152 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.27 //y=0.71 //x2=23.155 //y2=0.71
r307 (  122 157 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.49 //y=0.71 //x2=23.605 //y2=0.71
r308 (  122 123 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=23.49 //y=0.71 //x2=23.27 //y2=0.71
r309 (  119 154 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=23.21 //y=4.865 //x2=23.21 //y2=4.7
r310 (  118 151 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=23.115 //y=1.915 //x2=23.31 //y2=2.08
r311 (  117 153 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.115 //y=1.52 //x2=23.155 //y2=1.365
r312 (  117 118 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=23.115 //y=1.52 //x2=23.115 //y2=1.915
r313 (  116 153 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.115 //y=1.21 //x2=23.155 //y2=1.365
r314 (  115 152 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.115 //y=0.865 //x2=23.155 //y2=0.71
r315 (  115 116 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=23.115 //y=0.865 //x2=23.115 //y2=1.21
r316 (  114 145 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=21.35 //y=1.92 //x2=21.35 //y2=2.085
r317 (  113 144 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.35 //y=1.565 //x2=21.31 //y2=1.41
r318 (  113 114 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=21.35 //y=1.565 //x2=21.35 //y2=1.92
r319 (  112 144 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.35 //y=1.255 //x2=21.31 //y2=1.41
r320 (  111 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.35 //y=0.91 //x2=21.31 //y2=0.755
r321 (  111 112 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=21.35 //y=0.91 //x2=21.35 //y2=1.255
r322 (  108 149 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=21.305 //y=4.865 //x2=21.46 //y2=4.7
r323 (  106 142 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.975 //y=1.41 //x2=20.86 //y2=1.41
r324 (  105 144 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.195 //y=1.41 //x2=21.31 //y2=1.41
r325 (  104 141 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.975 //y=0.755 //x2=20.86 //y2=0.755
r326 (  103 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.195 //y=0.755 //x2=21.31 //y2=0.755
r327 (  103 104 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=21.195 //y=0.755 //x2=20.975 //y2=0.755
r328 (  101 108 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=21.23 //y=4.79 //x2=21.305 //y2=4.865
r329 (  101 102 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=21.23 //y=4.79 //x2=20.94 //y2=4.79
r330 (  98 102 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.865 //y=4.865 //x2=20.94 //y2=4.79
r331 (  97 142 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.82 //y=1.255 //x2=20.86 //y2=1.41
r332 (  96 141 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.82 //y=0.91 //x2=20.86 //y2=0.755
r333 (  96 97 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.82 //y=0.91 //x2=20.82 //y2=1.255
r334 (  93 140 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=18.1 //y=4.865 //x2=17.76 //y2=4.7
r335 (  90 138 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=17.66 //y=4.865 //x2=17.66 //y2=4.7
r336 (  89 137 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.735 //y=1.255 //x2=15.695 //y2=1.41
r337 (  88 136 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.735 //y=0.91 //x2=15.695 //y2=0.755
r338 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.735 //y=0.91 //x2=15.735 //y2=1.255
r339 (  86 133 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.36 //y=1.41 //x2=15.245 //y2=1.41
r340 (  85 137 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.58 //y=1.41 //x2=15.695 //y2=1.41
r341 (  84 132 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.36 //y=0.755 //x2=15.245 //y2=0.755
r342 (  83 136 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.58 //y=0.755 //x2=15.695 //y2=0.755
r343 (  83 84 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=15.58 //y=0.755 //x2=15.36 //y2=0.755
r344 (  82 135 ) resistor r=67.2792 //w=0.24 //l=0.438891 //layer=ply \
 //thickness=0.18 //x=15.205 //y=1.92 //x2=15.54 //y2=2.16
r345 (  81 133 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.205 //y=1.565 //x2=15.245 //y2=1.41
r346 (  81 82 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=15.205 //y=1.565 //x2=15.205 //y2=1.92
r347 (  80 133 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.205 //y=1.255 //x2=15.245 //y2=1.41
r348 (  79 132 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.205 //y=0.91 //x2=15.245 //y2=0.755
r349 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.205 //y=0.91 //x2=15.205 //y2=1.255
r350 (  78 129 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=23.65 //y=6.02 //x2=23.65 //y2=4.865
r351 (  77 119 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=23.21 //y=6.02 //x2=23.21 //y2=4.865
r352 (  76 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.305 //y=6.02 //x2=21.305 //y2=4.865
r353 (  75 98 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.865 //y=6.02 //x2=20.865 //y2=4.865
r354 (  74 93 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.1 //y=6.02 //x2=18.1 //y2=4.865
r355 (  73 90 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.66 //y=6.02 //x2=17.66 //y2=4.865
r356 (  72 124 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.38 //y=1.365 //x2=23.49 //y2=1.365
r357 (  72 125 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.38 //y=1.365 //x2=23.27 //y2=1.365
r358 (  71 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=21.085 //y=1.41 //x2=21.195 //y2=1.41
r359 (  71 106 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=21.085 //y=1.41 //x2=20.975 //y2=1.41
r360 (  70 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.47 //y=1.41 //x2=15.58 //y2=1.41
r361 (  70 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.47 //y=1.41 //x2=15.36 //y2=1.41
r362 (  68 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=23.31 //y=4.7 //x2=23.31 //y2=4.7
r363 (  58 151 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=23.31 //y=2.08 //x2=23.31 //y2=2.08
r364 (  55 149 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.46 //y=4.7 //x2=21.46 //y2=4.7
r365 (  44 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.46 //y=2.085 //x2=21.46 //y2=2.085
r366 (  41 140 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.76 //y=4.7 //x2=17.76 //y2=4.7
r367 (  32 135 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.54 //y=2.085 //x2=15.54 //y2=2.085
r368 (  30 68 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=23.31 //y=4.44 //x2=23.31 //y2=4.7
r369 (  29 30 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.31 //y=4.07 //x2=23.31 //y2=4.44
r370 (  28 29 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.31 //y=3.7 //x2=23.31 //y2=4.07
r371 (  27 28 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.31 //y=3.33 //x2=23.31 //y2=3.7
r372 (  26 27 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.31 //y=2.96 //x2=23.31 //y2=3.33
r373 (  25 26 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.31 //y=2.59 //x2=23.31 //y2=2.96
r374 (  25 58 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=23.31 //y=2.59 //x2=23.31 //y2=2.08
r375 (  24 55 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=21.46 //y=4.44 //x2=21.46 //y2=4.7
r376 (  23 24 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.46 //y=4.07 //x2=21.46 //y2=4.44
r377 (  22 23 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.46 //y=3.7 //x2=21.46 //y2=4.07
r378 (  21 22 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.46 //y=3.33 //x2=21.46 //y2=3.7
r379 (  20 21 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.96 //x2=21.46 //y2=3.33
r380 (  19 20 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.59 //x2=21.46 //y2=2.96
r381 (  19 44 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.59 //x2=21.46 //y2=2.085
r382 (  18 41 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=17.76 //y=4.44 //x2=17.76 //y2=4.7
r383 (  17 32 ) resistor r=59.893 //w=0.187 //l=0.875 //layer=li \
 //thickness=0.1 //x=15.54 //y=2.96 //x2=15.54 //y2=2.085
r384 (  16 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=23.31 //y=4.44 //x2=23.31 //y2=4.44
r385 (  14 20 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.46 //y=2.96 //x2=21.46 //y2=2.96
r386 (  12 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.46 //y=4.44 //x2=21.46 //y2=4.44
r387 (  10 18 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.76 //y=4.44 //x2=17.76 //y2=4.44
r388 (  8 17 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.54 //y=2.96 //x2=15.54 //y2=2.96
r389 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.575 //y=4.44 //x2=21.46 //y2=4.44
r390 (  5 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.195 //y=4.44 //x2=23.31 //y2=4.44
r391 (  5 6 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=23.195 //y=4.44 //x2=21.575 //y2=4.44
r392 (  4 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.875 //y=4.44 //x2=17.76 //y2=4.44
r393 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=4.44 //x2=21.46 //y2=4.44
r394 (  3 4 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=4.44 //x2=17.875 //y2=4.44
r395 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.655 //y=2.96 //x2=15.54 //y2=2.96
r396 (  1 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=2.96 //x2=21.46 //y2=2.96
r397 (  1 2 ) resistor r=5.42939 //w=0.131 //l=5.69 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=2.96 //x2=15.655 //y2=2.96
ends PM_FA\%CIN

subckt PM_FA\%noxref_12 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 48 52 \
 53 54 56 62 63 65 73 75 76 )
c139 ( 76 0 ) capacitor c=0.0220291f //x=24.165 //y=5.02
c140 ( 75 0 ) capacitor c=0.0217503f //x=23.285 //y=5.02
c141 ( 73 0 ) capacitor c=0.0084702f //x=24.16 //y=0.905
c142 ( 65 0 ) capacitor c=0.0530483f //x=26.27 //y=2.085
c143 ( 63 0 ) capacitor c=0.0435629f //x=26.91 //y=1.255
c144 ( 62 0 ) capacitor c=0.0199463f //x=26.91 //y=0.91
c145 ( 56 0 ) capacitor c=0.0148979f //x=26.755 //y=1.41
c146 ( 54 0 ) capacitor c=0.0157804f //x=26.755 //y=0.755
c147 ( 53 0 ) capacitor c=0.0527191f //x=26.5 //y=4.79
c148 ( 52 0 ) capacitor c=0.0322367f //x=26.79 //y=4.79
c149 ( 48 0 ) capacitor c=0.0293214f //x=26.38 //y=1.92
c150 ( 47 0 ) capacitor c=0.0250027f //x=26.38 //y=1.565
c151 ( 46 0 ) capacitor c=0.0234316f //x=26.38 //y=1.255
c152 ( 45 0 ) capacitor c=0.0199673f //x=26.38 //y=0.91
c153 ( 44 0 ) capacitor c=0.154131f //x=26.865 //y=6.02
c154 ( 43 0 ) capacitor c=0.154154f //x=26.425 //y=6.02
c155 ( 41 0 ) capacitor c=0.00194742f //x=24.31 //y=5.2
c156 ( 34 0 ) capacitor c=0.088828f //x=26.27 //y=2.085
c157 ( 32 0 ) capacitor c=0.110774f //x=24.79 //y=3.33
c158 ( 28 0 ) capacitor c=0.00384212f //x=24.435 //y=1.655
c159 ( 27 0 ) capacitor c=0.0158293f //x=24.705 //y=1.655
c160 ( 25 0 ) capacitor c=0.013629f //x=24.705 //y=5.2
c161 ( 14 0 ) capacitor c=0.00238935f //x=23.515 //y=5.2
c162 ( 13 0 ) capacitor c=0.0136432f //x=24.225 //y=5.2
c163 ( 2 0 ) capacitor c=0.0111187f //x=24.905 //y=3.33
c164 ( 1 0 ) capacitor c=0.0546065f //x=26.155 //y=3.33
r165 (  65 66 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=26.27 //y=2.085 //x2=26.38 //y2=2.085
r166 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.91 //y=1.255 //x2=26.87 //y2=1.41
r167 (  62 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.91 //y=0.91 //x2=26.87 //y2=0.755
r168 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=26.91 //y=0.91 //x2=26.91 //y2=1.255
r169 (  57 70 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.535 //y=1.41 //x2=26.42 //y2=1.41
r170 (  56 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.755 //y=1.41 //x2=26.87 //y2=1.41
r171 (  55 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.535 //y=0.755 //x2=26.42 //y2=0.755
r172 (  54 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.755 //y=0.755 //x2=26.87 //y2=0.755
r173 (  54 55 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=26.755 //y=0.755 //x2=26.535 //y2=0.755
r174 (  52 59 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=26.79 //y=4.79 //x2=26.865 //y2=4.865
r175 (  52 53 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=26.79 //y=4.79 //x2=26.5 //y2=4.79
r176 (  49 53 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=26.425 //y=4.865 //x2=26.5 //y2=4.79
r177 (  49 68 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=26.425 //y=4.865 //x2=26.27 //y2=4.7
r178 (  48 66 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=26.38 //y=1.92 //x2=26.38 //y2=2.085
r179 (  47 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.38 //y=1.565 //x2=26.42 //y2=1.41
r180 (  47 48 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=26.38 //y=1.565 //x2=26.38 //y2=1.92
r181 (  46 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.38 //y=1.255 //x2=26.42 //y2=1.41
r182 (  45 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.38 //y=0.91 //x2=26.42 //y2=0.755
r183 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=26.38 //y=0.91 //x2=26.38 //y2=1.255
r184 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.865 //y=6.02 //x2=26.865 //y2=4.865
r185 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.425 //y=6.02 //x2=26.425 //y2=4.865
r186 (  42 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=26.645 //y=1.41 //x2=26.755 //y2=1.41
r187 (  42 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=26.645 //y=1.41 //x2=26.535 //y2=1.41
r188 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.27 //y=4.7 //x2=26.27 //y2=4.7
r189 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=26.27 //y=3.33 //x2=26.27 //y2=4.7
r190 (  34 65 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.27 //y=2.085 //x2=26.27 //y2=2.085
r191 (  34 37 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.085 //x2=26.27 //y2=3.33
r192 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=24.79 //y=5.115 //x2=24.79 //y2=3.33
r193 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=24.79 //y=1.74 //x2=24.79 //y2=3.33
r194 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=24.705 //y=1.655 //x2=24.79 //y2=1.74
r195 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=24.705 //y=1.655 //x2=24.435 //y2=1.655
r196 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.395 //y=5.2 //x2=24.31 //y2=5.2
r197 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=24.705 //y=5.2 //x2=24.79 //y2=5.115
r198 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=24.705 //y=5.2 //x2=24.395 //y2=5.2
r199 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=24.35 //y=1.57 //x2=24.435 //y2=1.655
r200 (  21 73 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.35 //y=1.57 //x2=24.35 //y2=1
r201 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.31 //y=5.285 //x2=24.31 //y2=5.2
r202 (  15 76 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=24.31 //y=5.285 //x2=24.31 //y2=5.725
r203 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.225 //y=5.2 //x2=24.31 //y2=5.2
r204 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=24.225 //y=5.2 //x2=23.515 //y2=5.2
r205 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.43 //y=5.285 //x2=23.515 //y2=5.2
r206 (  7 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=23.43 //y=5.285 //x2=23.43 //y2=5.725
r207 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=26.27 //y=3.33 //x2=26.27 //y2=3.33
r208 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=24.79 //y=3.33 //x2=24.79 //y2=3.33
r209 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=24.905 //y=3.33 //x2=24.79 //y2=3.33
r210 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=26.155 //y=3.33 //x2=26.27 //y2=3.33
r211 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=26.155 //y=3.33 //x2=24.905 //y2=3.33
ends PM_FA\%noxref_12

subckt PM_FA\%noxref_13 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 48 52 \
 53 54 56 62 63 65 73 75 76 )
c142 ( 76 0 ) capacitor c=0.0220291f //x=29.715 //y=5.02
c143 ( 75 0 ) capacitor c=0.0217503f //x=28.835 //y=5.02
c144 ( 73 0 ) capacitor c=0.0084702f //x=29.71 //y=0.905
c145 ( 65 0 ) capacitor c=0.0511458f //x=31.82 //y=2.085
c146 ( 63 0 ) capacitor c=0.0435629f //x=32.46 //y=1.255
c147 ( 62 0 ) capacitor c=0.0200386f //x=32.46 //y=0.91
c148 ( 56 0 ) capacitor c=0.0152946f //x=32.305 //y=1.41
c149 ( 54 0 ) capacitor c=0.0157804f //x=32.305 //y=0.755
c150 ( 53 0 ) capacitor c=0.0524991f //x=32.05 //y=4.79
c151 ( 52 0 ) capacitor c=0.0323689f //x=32.34 //y=4.79
c152 ( 48 0 ) capacitor c=0.0290017f //x=31.93 //y=1.92
c153 ( 47 0 ) capacitor c=0.0250027f //x=31.93 //y=1.565
c154 ( 46 0 ) capacitor c=0.0234316f //x=31.93 //y=1.255
c155 ( 45 0 ) capacitor c=0.0200596f //x=31.93 //y=0.91
c156 ( 44 0 ) capacitor c=0.154218f //x=32.415 //y=6.02
c157 ( 43 0 ) capacitor c=0.154243f //x=31.975 //y=6.02
c158 ( 41 0 ) capacitor c=0.00279371f //x=29.86 //y=5.2
c159 ( 34 0 ) capacitor c=0.0918279f //x=31.82 //y=2.085
c160 ( 32 0 ) capacitor c=0.10823f //x=30.34 //y=3.33
c161 ( 28 0 ) capacitor c=0.00468667f //x=29.985 //y=1.655
c162 ( 27 0 ) capacitor c=0.0131863f //x=30.255 //y=1.655
c163 ( 25 0 ) capacitor c=0.0148609f //x=30.255 //y=5.2
c164 ( 14 0 ) capacitor c=0.0022661f //x=29.065 //y=5.2
c165 ( 13 0 ) capacitor c=0.0169929f //x=29.775 //y=5.2
c166 ( 2 0 ) capacitor c=0.0113927f //x=30.455 //y=3.33
c167 ( 1 0 ) capacitor c=0.0516026f //x=31.705 //y=3.33
r168 (  65 66 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=31.82 //y=2.085 //x2=31.93 //y2=2.085
r169 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.46 //y=1.255 //x2=32.42 //y2=1.41
r170 (  62 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.46 //y=0.91 //x2=32.42 //y2=0.755
r171 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=32.46 //y=0.91 //x2=32.46 //y2=1.255
r172 (  57 70 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.085 //y=1.41 //x2=31.97 //y2=1.41
r173 (  56 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.305 //y=1.41 //x2=32.42 //y2=1.41
r174 (  55 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.085 //y=0.755 //x2=31.97 //y2=0.755
r175 (  54 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.305 //y=0.755 //x2=32.42 //y2=0.755
r176 (  54 55 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=32.305 //y=0.755 //x2=32.085 //y2=0.755
r177 (  52 59 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=32.34 //y=4.79 //x2=32.415 //y2=4.865
r178 (  52 53 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=32.34 //y=4.79 //x2=32.05 //y2=4.79
r179 (  49 53 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=31.975 //y=4.865 //x2=32.05 //y2=4.79
r180 (  49 68 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=31.975 //y=4.865 //x2=31.82 //y2=4.7
r181 (  48 66 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=31.93 //y=1.92 //x2=31.93 //y2=2.085
r182 (  47 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.93 //y=1.565 //x2=31.97 //y2=1.41
r183 (  47 48 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=31.93 //y=1.565 //x2=31.93 //y2=1.92
r184 (  46 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.93 //y=1.255 //x2=31.97 //y2=1.41
r185 (  45 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.93 //y=0.91 //x2=31.97 //y2=0.755
r186 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=31.93 //y=0.91 //x2=31.93 //y2=1.255
r187 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=32.415 //y=6.02 //x2=32.415 //y2=4.865
r188 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=31.975 //y=6.02 //x2=31.975 //y2=4.865
r189 (  42 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=32.195 //y=1.41 //x2=32.305 //y2=1.41
r190 (  42 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=32.195 //y=1.41 //x2=32.085 //y2=1.41
r191 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.82 //y=4.7 //x2=31.82 //y2=4.7
r192 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=31.82 //y=3.33 //x2=31.82 //y2=4.7
r193 (  34 65 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.82 //y=2.085 //x2=31.82 //y2=2.085
r194 (  34 37 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=31.82 //y=2.085 //x2=31.82 //y2=3.33
r195 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=30.34 //y=5.115 //x2=30.34 //y2=3.33
r196 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=30.34 //y=1.74 //x2=30.34 //y2=3.33
r197 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=30.255 //y=1.655 //x2=30.34 //y2=1.74
r198 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=30.255 //y=1.655 //x2=29.985 //y2=1.655
r199 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.945 //y=5.2 //x2=29.86 //y2=5.2
r200 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=30.255 //y=5.2 //x2=30.34 //y2=5.115
r201 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=30.255 //y=5.2 //x2=29.945 //y2=5.2
r202 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=29.9 //y=1.57 //x2=29.985 //y2=1.655
r203 (  21 73 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=29.9 //y=1.57 //x2=29.9 //y2=1
r204 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.86 //y=5.285 //x2=29.86 //y2=5.2
r205 (  15 76 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=29.86 //y=5.285 //x2=29.86 //y2=5.725
r206 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.775 //y=5.2 //x2=29.86 //y2=5.2
r207 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=29.775 //y=5.2 //x2=29.065 //y2=5.2
r208 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=28.98 //y=5.285 //x2=29.065 //y2=5.2
r209 (  7 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=28.98 //y=5.285 //x2=28.98 //y2=5.725
r210 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=31.82 //y=3.33 //x2=31.82 //y2=3.33
r211 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=30.34 //y=3.33 //x2=30.34 //y2=3.33
r212 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=30.455 //y=3.33 //x2=30.34 //y2=3.33
r213 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.705 //y=3.33 //x2=31.82 //y2=3.33
r214 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=31.705 //y=3.33 //x2=30.455 //y2=3.33
ends PM_FA\%noxref_13

subckt PM_FA\%noxref_14 ( 1 2 17 18 19 20 24 27 32 34 35 36 37 38 39 40 44 46 \
 49 51 52 57 67 69 )
c165 ( 69 0 ) capacitor c=0.0279852f //x=26.5 //y=5.02
c166 ( 67 0 ) capacitor c=0.016967f //x=26.455 //y=0.91
c167 ( 57 0 ) capacitor c=0.0422106f //x=34.255 //y=4.705
c168 ( 52 0 ) capacitor c=0.0321911f //x=34.745 //y=1.25
c169 ( 51 0 ) capacitor c=0.0185201f //x=34.745 //y=0.905
c170 ( 49 0 ) capacitor c=0.0344254f //x=34.675 //y=4.795
c171 ( 46 0 ) capacitor c=0.0133656f //x=34.59 //y=1.405
c172 ( 44 0 ) capacitor c=0.0157804f //x=34.59 //y=0.75
c173 ( 40 0 ) capacitor c=0.0788505f //x=34.215 //y=1.915
c174 ( 39 0 ) capacitor c=0.022867f //x=34.215 //y=1.56
c175 ( 38 0 ) capacitor c=0.0234318f //x=34.215 //y=1.25
c176 ( 37 0 ) capacitor c=0.0192004f //x=34.215 //y=0.905
c177 ( 36 0 ) capacitor c=0.110795f //x=34.75 //y=6.025
c178 ( 35 0 ) capacitor c=0.153847f //x=34.31 //y=6.025
c179 ( 32 0 ) capacitor c=0.00993392f //x=34.255 //y=4.705
c180 ( 27 0 ) capacitor c=0.0921769f //x=34.41 //y=2.08
c181 ( 24 0 ) capacitor c=0.0882674f //x=27.01 //y=2.96
c182 ( 20 0 ) capacitor c=0.00573423f //x=26.73 //y=4.58
c183 ( 19 0 ) capacitor c=0.0118959f //x=26.925 //y=4.58
c184 ( 18 0 ) capacitor c=0.00630489f //x=26.725 //y=2.08
c185 ( 17 0 ) capacitor c=0.012513f //x=26.925 //y=2.08
c186 ( 2 0 ) capacitor c=0.0155528f //x=27.125 //y=2.96
c187 ( 1 0 ) capacitor c=0.23241f //x=34.295 //y=2.96
r188 (  59 60 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=34.255 //y=4.795 //x2=34.255 //y2=4.87
r189 (  57 59 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=34.255 //y=4.705 //x2=34.255 //y2=4.795
r190 (  52 66 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.745 //y=1.25 //x2=34.705 //y2=1.405
r191 (  51 65 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.745 //y=0.905 //x2=34.705 //y2=0.75
r192 (  51 52 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=34.745 //y=0.905 //x2=34.745 //y2=1.25
r193 (  50 59 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=34.39 //y=4.795 //x2=34.255 //y2=4.795
r194 (  49 53 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=34.675 //y=4.795 //x2=34.75 //y2=4.87
r195 (  49 50 ) resistor r=146.138 //w=0.094 //l=0.285 //layer=ply \
 //thickness=0.18 //x=34.675 //y=4.795 //x2=34.39 //y2=4.795
r196 (  47 64 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.37 //y=1.405 //x2=34.255 //y2=1.405
r197 (  46 66 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.59 //y=1.405 //x2=34.705 //y2=1.405
r198 (  45 63 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.37 //y=0.75 //x2=34.255 //y2=0.75
r199 (  44 65 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.59 //y=0.75 //x2=34.705 //y2=0.75
r200 (  44 45 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=34.59 //y=0.75 //x2=34.37 //y2=0.75
r201 (  40 62 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=34.215 //y=1.915 //x2=34.41 //y2=2.08
r202 (  39 64 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.215 //y=1.56 //x2=34.255 //y2=1.405
r203 (  39 40 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=34.215 //y=1.56 //x2=34.215 //y2=1.915
r204 (  38 64 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.215 //y=1.25 //x2=34.255 //y2=1.405
r205 (  37 63 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.215 //y=0.905 //x2=34.255 //y2=0.75
r206 (  37 38 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=34.215 //y=0.905 //x2=34.215 //y2=1.25
r207 (  36 53 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=34.75 //y=6.025 //x2=34.75 //y2=4.87
r208 (  35 60 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=34.31 //y=6.025 //x2=34.31 //y2=4.87
r209 (  34 46 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=34.48 //y=1.405 //x2=34.59 //y2=1.405
r210 (  34 47 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=34.48 //y=1.405 //x2=34.37 //y2=1.405
r211 (  32 57 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.255 //y=4.705 //x2=34.255 //y2=4.705
r212 (  32 33 ) resistor r=7.81102 //w=0.254 //l=0.155 //layer=li \
 //thickness=0.1 //x=34.255 //y=4.705 //x2=34.41 //y2=4.705
r213 (  27 62 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.41 //y=2.08 //x2=34.41 //y2=2.08
r214 (  27 30 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=34.41 //y=2.08 //x2=34.41 //y2=2.96
r215 (  25 33 ) resistor r=3.23951 //w=0.254 //l=0.165 //layer=li \
 //thickness=0.1 //x=34.41 //y=4.54 //x2=34.41 //y2=4.705
r216 (  25 30 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=34.41 //y=4.54 //x2=34.41 //y2=2.96
r217 (  22 24 ) resistor r=105.07 //w=0.187 //l=1.535 //layer=li \
 //thickness=0.1 //x=27.01 //y=4.495 //x2=27.01 //y2=2.96
r218 (  21 24 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=27.01 //y=2.165 //x2=27.01 //y2=2.96
r219 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=26.925 //y=4.58 //x2=27.01 //y2=4.495
r220 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=26.925 //y=4.58 //x2=26.73 //y2=4.58
r221 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=26.925 //y=2.08 //x2=27.01 //y2=2.165
r222 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=26.925 //y=2.08 //x2=26.725 //y2=2.08
r223 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=26.645 //y=4.665 //x2=26.73 //y2=4.58
r224 (  11 69 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=26.645 //y=4.665 //x2=26.645 //y2=5.725
r225 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=26.64 //y=1.995 //x2=26.725 //y2=2.08
r226 (  7 67 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=26.64 //y=1.995 //x2=26.64 //y2=1.005
r227 (  6 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=34.41 //y=2.96 //x2=34.41 //y2=2.96
r228 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=27.01 //y=2.96 //x2=27.01 //y2=2.96
r229 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=27.125 //y=2.96 //x2=27.01 //y2=2.96
r230 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.295 //y=2.96 //x2=34.41 //y2=2.96
r231 (  1 2 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=34.295 //y=2.96 //x2=27.125 //y2=2.96
ends PM_FA\%noxref_14

subckt PM_FA\%noxref_15 ( 1 2 17 18 19 20 24 25 27 33 34 35 36 37 38 43 45 47 \
 53 54 56 57 60 68 70 )
c137 ( 70 0 ) capacitor c=0.0288456f //x=32.05 //y=5.02
c138 ( 68 0 ) capacitor c=0.0172738f //x=32.005 //y=0.91
c139 ( 60 0 ) capacitor c=0.0369822f //x=35.185 //y=4.705
c140 ( 57 0 ) capacitor c=0.0279572f //x=35.15 //y=1.915
c141 ( 56 0 ) capacitor c=0.0413537f //x=35.15 //y=2.08
c142 ( 54 0 ) capacitor c=0.0237734f //x=35.715 //y=1.255
c143 ( 53 0 ) capacitor c=0.0191782f //x=35.715 //y=0.905
c144 ( 47 0 ) capacitor c=0.0346941f //x=35.56 //y=1.405
c145 ( 45 0 ) capacitor c=0.0157803f //x=35.56 //y=0.75
c146 ( 43 0 ) capacitor c=0.0360787f //x=35.555 //y=4.795
c147 ( 38 0 ) capacitor c=0.0199921f //x=35.185 //y=1.56
c148 ( 37 0 ) capacitor c=0.0169608f //x=35.185 //y=1.255
c149 ( 36 0 ) capacitor c=0.0185462f //x=35.185 //y=0.905
c150 ( 35 0 ) capacitor c=0.15325f //x=35.63 //y=6.025
c151 ( 34 0 ) capacitor c=0.110232f //x=35.19 //y=6.025
c152 ( 27 0 ) capacitor c=0.0785323f //x=35.15 //y=2.08
c153 ( 25 0 ) capacitor c=0.00515516f //x=35.15 //y=4.54
c154 ( 24 0 ) capacitor c=0.0863121f //x=32.56 //y=3.33
c155 ( 20 0 ) capacitor c=0.00558395f //x=32.28 //y=4.58
c156 ( 19 0 ) capacitor c=0.0134399f //x=32.475 //y=4.58
c157 ( 18 0 ) capacitor c=0.00547024f //x=32.275 //y=2.08
c158 ( 17 0 ) capacitor c=0.013178f //x=32.475 //y=2.08
c159 ( 2 0 ) capacitor c=0.00731142f //x=32.675 //y=3.33
c160 ( 1 0 ) capacitor c=0.091903f //x=35.035 //y=3.33
r161 (  62 63 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=35.185 //y=4.795 //x2=35.185 //y2=4.87
r162 (  60 62 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=35.185 //y=4.705 //x2=35.185 //y2=4.795
r163 (  56 57 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=35.15 //y=2.08 //x2=35.15 //y2=1.915
r164 (  54 67 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=35.715 //y=1.255 //x2=35.715 //y2=1.367
r165 (  53 66 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.715 //y=0.905 //x2=35.675 //y2=0.75
r166 (  53 54 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=35.715 //y=0.905 //x2=35.715 //y2=1.255
r167 (  48 65 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.34 //y=1.405 //x2=35.225 //y2=1.405
r168 (  47 67 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=35.56 //y=1.405 //x2=35.715 //y2=1.367
r169 (  46 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.34 //y=0.75 //x2=35.225 //y2=0.75
r170 (  45 66 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=35.56 //y=0.75 //x2=35.675 //y2=0.75
r171 (  45 46 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=35.56 //y=0.75 //x2=35.34 //y2=0.75
r172 (  44 62 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=35.32 //y=4.795 //x2=35.185 //y2=4.795
r173 (  43 50 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=35.555 //y=4.795 //x2=35.63 //y2=4.87
r174 (  43 44 ) resistor r=120.5 //w=0.094 //l=0.235 //layer=ply \
 //thickness=0.18 //x=35.555 //y=4.795 //x2=35.32 //y2=4.795
r175 (  38 65 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.185 //y=1.56 //x2=35.225 //y2=1.405
r176 (  38 57 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=35.185 //y=1.56 //x2=35.185 //y2=1.915
r177 (  37 65 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=35.185 //y=1.255 //x2=35.225 //y2=1.405
r178 (  36 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.185 //y=0.905 //x2=35.225 //y2=0.75
r179 (  36 37 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=35.185 //y=0.905 //x2=35.185 //y2=1.255
r180 (  35 50 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=35.63 //y=6.025 //x2=35.63 //y2=4.87
r181 (  34 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=35.19 //y=6.025 //x2=35.19 //y2=4.87
r182 (  33 47 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=35.45 //y=1.405 //x2=35.56 //y2=1.405
r183 (  33 48 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=35.45 //y=1.405 //x2=35.34 //y2=1.405
r184 (  32 60 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=35.185 //y=4.705 //x2=35.185 //y2=4.705
r185 (  27 56 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=35.15 //y=2.08 //x2=35.15 //y2=2.08
r186 (  27 30 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=35.15 //y=2.08 //x2=35.15 //y2=3.33
r187 (  25 32 ) resistor r=11.332 //w=0.189 //l=0.173292 //layer=li \
 //thickness=0.1 //x=35.15 //y=4.54 //x2=35.167 //y2=4.705
r188 (  25 30 ) resistor r=82.8235 //w=0.187 //l=1.21 //layer=li \
 //thickness=0.1 //x=35.15 //y=4.54 //x2=35.15 //y2=3.33
r189 (  22 24 ) resistor r=79.7433 //w=0.187 //l=1.165 //layer=li \
 //thickness=0.1 //x=32.56 //y=4.495 //x2=32.56 //y2=3.33
r190 (  21 24 ) resistor r=79.7433 //w=0.187 //l=1.165 //layer=li \
 //thickness=0.1 //x=32.56 //y=2.165 //x2=32.56 //y2=3.33
r191 (  19 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.475 //y=4.58 //x2=32.56 //y2=4.495
r192 (  19 20 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=32.475 //y=4.58 //x2=32.28 //y2=4.58
r193 (  17 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.475 //y=2.08 //x2=32.56 //y2=2.165
r194 (  17 18 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li \
 //thickness=0.1 //x=32.475 //y=2.08 //x2=32.275 //y2=2.08
r195 (  11 20 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.195 //y=4.665 //x2=32.28 //y2=4.58
r196 (  11 70 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=32.195 //y=4.665 //x2=32.195 //y2=5.725
r197 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.19 //y=1.995 //x2=32.275 //y2=2.08
r198 (  7 68 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li \
 //thickness=0.1 //x=32.19 //y=1.995 //x2=32.19 //y2=1.005
r199 (  6 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=35.15 //y=3.33 //x2=35.15 //y2=3.33
r200 (  4 24 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=32.56 //y=3.33 //x2=32.56 //y2=3.33
r201 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=32.675 //y=3.33 //x2=32.56 //y2=3.33
r202 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=35.035 //y=3.33 //x2=35.15 //y2=3.33
r203 (  1 2 ) resistor r=2.25191 //w=0.131 //l=2.36 //layer=m1 \
 //thickness=0.36 //x=35.035 //y=3.33 //x2=32.675 //y2=3.33
ends PM_FA\%noxref_15

subckt PM_FA\%noxref_16 ( 1 2 11 12 23 24 25 30 32 40 41 42 43 44 45 46 50 51 \
 52 54 60 61 63 71 72 75 )
c140 ( 75 0 ) capacitor c=0.0159573f //x=35.265 //y=5.025
c141 ( 72 0 ) capacitor c=0.00905936f //x=35.26 //y=0.905
c142 ( 71 0 ) capacitor c=0.007684f //x=34.29 //y=0.905
c143 ( 63 0 ) capacitor c=0.0528806f //x=37.37 //y=2.085
c144 ( 61 0 ) capacitor c=0.0435629f //x=38.01 //y=1.255
c145 ( 60 0 ) capacitor c=0.0200386f //x=38.01 //y=0.91
c146 ( 54 0 ) capacitor c=0.0152946f //x=37.855 //y=1.41
c147 ( 52 0 ) capacitor c=0.0157804f //x=37.855 //y=0.755
c148 ( 51 0 ) capacitor c=0.0524991f //x=37.6 //y=4.79
c149 ( 50 0 ) capacitor c=0.0322983f //x=37.89 //y=4.79
c150 ( 46 0 ) capacitor c=0.0290017f //x=37.48 //y=1.92
c151 ( 45 0 ) capacitor c=0.0250027f //x=37.48 //y=1.565
c152 ( 44 0 ) capacitor c=0.0234316f //x=37.48 //y=1.255
c153 ( 43 0 ) capacitor c=0.0200596f //x=37.48 //y=0.91
c154 ( 42 0 ) capacitor c=0.154218f //x=37.965 //y=6.02
c155 ( 41 0 ) capacitor c=0.154243f //x=37.525 //y=6.02
c156 ( 39 0 ) capacitor c=0.00710337f //x=35.45 //y=1.655
c157 ( 32 0 ) capacitor c=0.0944545f //x=37.37 //y=2.085
c158 ( 30 0 ) capacitor c=0.112585f //x=35.89 //y=3.33
c159 ( 25 0 ) capacitor c=0.0162468f //x=35.805 //y=1.655
c160 ( 24 0 ) capacitor c=0.00499395f //x=35.495 //y=5.21
c161 ( 23 0 ) capacitor c=0.0155365f //x=35.805 //y=5.21
c162 ( 12 0 ) capacitor c=0.00210564f //x=34.565 //y=1.655
c163 ( 11 0 ) capacitor c=0.0217261f //x=35.365 //y=1.655
c164 ( 2 0 ) capacitor c=0.00861659f //x=36.005 //y=3.33
c165 ( 1 0 ) capacitor c=0.0802319f //x=37.255 //y=3.33
r166 (  63 64 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=37.37 //y=2.085 //x2=37.48 //y2=2.085
r167 (  61 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.01 //y=1.255 //x2=37.97 //y2=1.41
r168 (  60 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.01 //y=0.91 //x2=37.97 //y2=0.755
r169 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=38.01 //y=0.91 //x2=38.01 //y2=1.255
r170 (  55 68 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.635 //y=1.41 //x2=37.52 //y2=1.41
r171 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.855 //y=1.41 //x2=37.97 //y2=1.41
r172 (  53 67 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.635 //y=0.755 //x2=37.52 //y2=0.755
r173 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.855 //y=0.755 //x2=37.97 //y2=0.755
r174 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=37.855 //y=0.755 //x2=37.635 //y2=0.755
r175 (  50 57 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=37.89 //y=4.79 //x2=37.965 //y2=4.865
r176 (  50 51 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=37.89 //y=4.79 //x2=37.6 //y2=4.79
r177 (  47 51 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=37.525 //y=4.865 //x2=37.6 //y2=4.79
r178 (  47 66 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=37.525 //y=4.865 //x2=37.37 //y2=4.7
r179 (  46 64 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=37.48 //y=1.92 //x2=37.48 //y2=2.085
r180 (  45 68 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.48 //y=1.565 //x2=37.52 //y2=1.41
r181 (  45 46 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=37.48 //y=1.565 //x2=37.48 //y2=1.92
r182 (  44 68 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.48 //y=1.255 //x2=37.52 //y2=1.41
r183 (  43 67 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.48 //y=0.91 //x2=37.52 //y2=0.755
r184 (  43 44 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=37.48 //y=0.91 //x2=37.48 //y2=1.255
r185 (  42 57 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=37.965 //y=6.02 //x2=37.965 //y2=4.865
r186 (  41 47 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=37.525 //y=6.02 //x2=37.525 //y2=4.865
r187 (  40 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=37.745 //y=1.41 //x2=37.855 //y2=1.41
r188 (  40 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=37.745 //y=1.41 //x2=37.635 //y2=1.41
r189 (  37 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=37.37 //y=4.7 //x2=37.37 //y2=4.7
r190 (  35 37 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=37.37 //y=3.33 //x2=37.37 //y2=4.7
r191 (  32 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=37.37 //y=2.085 //x2=37.37 //y2=2.085
r192 (  32 35 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=37.37 //y=2.085 //x2=37.37 //y2=3.33
r193 (  28 30 ) resistor r=122.866 //w=0.187 //l=1.795 //layer=li \
 //thickness=0.1 //x=35.89 //y=5.125 //x2=35.89 //y2=3.33
r194 (  27 30 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=35.89 //y=1.74 //x2=35.89 //y2=3.33
r195 (  26 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.535 //y=1.655 //x2=35.45 //y2=1.655
r196 (  25 27 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=35.805 //y=1.655 //x2=35.89 //y2=1.74
r197 (  25 26 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=35.805 //y=1.655 //x2=35.535 //y2=1.655
r198 (  23 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=35.805 //y=5.21 //x2=35.89 //y2=5.125
r199 (  23 24 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=35.805 //y=5.21 //x2=35.495 //y2=5.21
r200 (  19 39 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.45 //y=1.57 //x2=35.45 //y2=1.655
r201 (  19 72 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=35.45 //y=1.57 //x2=35.45 //y2=1
r202 (  13 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=35.41 //y=5.295 //x2=35.495 //y2=5.21
r203 (  13 75 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=35.41 //y=5.295 //x2=35.41 //y2=5.72
r204 (  11 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.365 //y=1.655 //x2=35.45 //y2=1.655
r205 (  11 12 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li \
 //thickness=0.1 //x=35.365 //y=1.655 //x2=34.565 //y2=1.655
r206 (  7 12 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=34.48 //y=1.57 //x2=34.565 //y2=1.655
r207 (  7 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=34.48 //y=1.57 //x2=34.48 //y2=1
r208 (  6 35 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=37.37 //y=3.33 //x2=37.37 //y2=3.33
r209 (  4 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=35.89 //y=3.33 //x2=35.89 //y2=3.33
r210 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=36.005 //y=3.33 //x2=35.89 //y2=3.33
r211 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=37.255 //y=3.33 //x2=37.37 //y2=3.33
r212 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=37.255 //y=3.33 //x2=36.005 //y2=3.33
ends PM_FA\%noxref_16

subckt PM_FA\%noxref_17 ( 7 8 15 16 23 24 25 )
c39 ( 25 0 ) capacitor c=0.0306618f //x=4.625 //y=5.02
c40 ( 24 0 ) capacitor c=0.0185379f //x=3.745 //y=5.02
c41 ( 23 0 ) capacitor c=0.0384176f //x=2.875 //y=5.02
c42 ( 16 0 ) capacitor c=0.00194711f //x=3.975 //y=6.905
c43 ( 15 0 ) capacitor c=0.014216f //x=4.685 //y=6.905
c44 ( 8 0 ) capacitor c=0.00644339f //x=3.095 //y=5.205
c45 ( 7 0 ) capacitor c=0.0207865f //x=3.805 //y=5.205
r46 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.77 //y=6.82 //x2=4.77 //y2=6.735
r47 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.685 //y=6.905 //x2=4.77 //y2=6.82
r48 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=4.685 //y=6.905 //x2=3.975 //y2=6.905
r49 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.89 //y=6.82 //x2=3.975 //y2=6.905
r50 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=3.89 //y=6.82 //x2=3.89 //y2=6.395
r51 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=3.89 //y=5.29 //x2=3.89 //y2=5.715
r52 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.805 //y=5.205 //x2=3.89 //y2=5.29
r53 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=3.805 //y=5.205 //x2=3.095 //y2=5.205
r54 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.01 //y=5.29 //x2=3.095 //y2=5.205
r55 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=3.01 //y=5.29 //x2=3.01 //y2=5.715
ends PM_FA\%noxref_17

subckt PM_FA\%noxref_18 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0629093f //x=2.78 //y=0.37
c52 ( 17 0 ) capacitor c=0.00723243f //x=4.855 //y=0.62
c53 ( 13 0 ) capacitor c=0.0149083f //x=4.77 //y=0.535
c54 ( 10 0 ) capacitor c=0.00604817f //x=3.885 //y=1.5
c55 ( 9 0 ) capacitor c=0.00677124f //x=3.885 //y=0.62
c56 ( 5 0 ) capacitor c=0.0230272f //x=3.8 //y=1.585
c57 ( 1 0 ) capacitor c=0.0076549f //x=2.915 //y=1.5
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.855 //y=0.62 //x2=4.855 //y2=0.495
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.855 //y=0.62 //x2=4.855 //y2=0.885
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.97 //y=0.535 //x2=3.885 //y2=0.495
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.97 //y=0.535 //x2=4.37 //y2=0.535
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.77 //y=0.535 //x2=4.855 //y2=0.495
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.77 //y=0.535 //x2=4.37 //y2=0.535
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=3.885 //y=1.5 //x2=3.885 //y2=1.625
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=3.885 //y=1.5 //x2=3.885 //y2=0.885
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.885 //y=0.62 //x2=3.885 //y2=0.495
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.885 //y=0.62 //x2=3.885 //y2=0.885
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3 //y=1.585 //x2=2.915 //y2=1.625
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3 //y=1.585 //x2=3.4 //y2=1.585
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.8 //y=1.585 //x2=3.885 //y2=1.625
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.8 //y=1.585 //x2=3.4 //y2=1.585
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=2.915 //y=1.5 //x2=2.915 //y2=1.625
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.915 //y=1.5 //x2=2.915 //y2=0.885
ends PM_FA\%noxref_18

subckt PM_FA\%noxref_19 ( 7 8 15 16 23 24 25 )
c41 ( 25 0 ) capacitor c=0.0305804f //x=7.955 //y=5.02
c42 ( 24 0 ) capacitor c=0.0185379f //x=7.075 //y=5.02
c43 ( 23 0 ) capacitor c=0.0384176f //x=6.205 //y=5.02
c44 ( 16 0 ) capacitor c=0.00194711f //x=7.305 //y=6.905
c45 ( 15 0 ) capacitor c=0.0133643f //x=8.015 //y=6.905
c46 ( 8 0 ) capacitor c=0.00631451f //x=6.425 //y=5.205
c47 ( 7 0 ) capacitor c=0.0183784f //x=7.135 //y=5.205
r48 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.1 //y=6.82 //x2=8.1 //y2=6.735
r49 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.015 //y=6.905 //x2=8.1 //y2=6.82
r50 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.015 //y=6.905 //x2=7.305 //y2=6.905
r51 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.22 //y=6.82 //x2=7.305 //y2=6.905
r52 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=7.22 //y=6.82 //x2=7.22 //y2=6.395
r53 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.29 //x2=7.22 //y2=5.715
r54 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.205 //x2=7.22 //y2=5.29
r55 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=7.135 //y=5.205 //x2=6.425 //y2=5.205
r56 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.29 //x2=6.425 //y2=5.205
r57 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.29 //x2=6.34 //y2=5.715
ends PM_FA\%noxref_19

subckt PM_FA\%noxref_20 ( 1 5 9 10 13 17 29 )
c50 ( 29 0 ) capacitor c=0.0630989f //x=6.11 //y=0.37
c51 ( 17 0 ) capacitor c=0.00723243f //x=8.185 //y=0.62
c52 ( 13 0 ) capacitor c=0.0149083f //x=8.1 //y=0.535
c53 ( 10 0 ) capacitor c=0.00604817f //x=7.215 //y=1.5
c54 ( 9 0 ) capacitor c=0.00677124f //x=7.215 //y=0.62
c55 ( 5 0 ) capacitor c=0.0245898f //x=7.13 //y=1.585
c56 ( 1 0 ) capacitor c=0.0071362f //x=6.245 //y=1.5
r57 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=8.185 //y=0.62 //x2=8.185 //y2=0.495
r58 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=8.185 //y=0.62 //x2=8.185 //y2=0.885
r59 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.3 //y=0.535 //x2=7.215 //y2=0.495
r60 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.3 //y=0.535 //x2=7.7 //y2=0.535
r61 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.1 //y=0.535 //x2=8.185 //y2=0.495
r62 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.1 //y=0.535 //x2=7.7 //y2=0.535
r63 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=7.215 //y=1.5 //x2=7.215 //y2=1.625
r64 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=7.215 //y=1.5 //x2=7.215 //y2=0.885
r65 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=7.215 //y=0.62 //x2=7.215 //y2=0.495
r66 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=7.215 //y=0.62 //x2=7.215 //y2=0.885
r67 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.33 //y=1.585 //x2=6.245 //y2=1.625
r68 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.33 //y=1.585 //x2=6.73 //y2=1.585
r69 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.13 //y=1.585 //x2=7.215 //y2=1.625
r70 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.13 //y=1.585 //x2=6.73 //y2=1.585
r71 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.245 //y=1.5 //x2=6.245 //y2=1.625
r72 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.245 //y=1.5 //x2=6.245 //y2=0.885
ends PM_FA\%noxref_20

subckt PM_FA\%noxref_21 ( 7 8 15 16 23 24 25 )
c37 ( 25 0 ) capacitor c=0.0304741f //x=15.725 //y=5.02
c38 ( 24 0 ) capacitor c=0.0185379f //x=14.845 //y=5.02
c39 ( 23 0 ) capacitor c=0.0384176f //x=13.975 //y=5.02
c40 ( 16 0 ) capacitor c=0.00194711f //x=15.075 //y=6.905
c41 ( 15 0 ) capacitor c=0.0133605f //x=15.785 //y=6.905
c42 ( 8 0 ) capacitor c=0.00580995f //x=14.195 //y=5.205
c43 ( 7 0 ) capacitor c=0.0174896f //x=14.905 //y=5.205
r44 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.87 //y=6.82 //x2=15.87 //y2=6.735
r45 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.785 //y=6.905 //x2=15.87 //y2=6.82
r46 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=15.785 //y=6.905 //x2=15.075 //y2=6.905
r47 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.99 //y=6.82 //x2=15.075 //y2=6.905
r48 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=14.99 //y=6.82 //x2=14.99 //y2=6.395
r49 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=14.99 //y=5.29 //x2=14.99 //y2=5.715
r50 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.905 //y=5.205 //x2=14.99 //y2=5.29
r51 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=14.905 //y=5.205 //x2=14.195 //y2=5.205
r52 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.11 //y=5.29 //x2=14.195 //y2=5.205
r53 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=14.11 //y=5.29 //x2=14.11 //y2=5.715
ends PM_FA\%noxref_21

subckt PM_FA\%noxref_22 ( 1 5 9 10 13 17 29 )
c49 ( 29 0 ) capacitor c=0.0629093f //x=13.88 //y=0.37
c50 ( 17 0 ) capacitor c=0.00723243f //x=15.955 //y=0.62
c51 ( 13 0 ) capacitor c=0.0149083f //x=15.87 //y=0.535
c52 ( 10 0 ) capacitor c=0.00604817f //x=14.985 //y=1.5
c53 ( 9 0 ) capacitor c=0.00677124f //x=14.985 //y=0.62
c54 ( 5 0 ) capacitor c=0.0245898f //x=14.9 //y=1.585
c55 ( 1 0 ) capacitor c=0.0071362f //x=14.015 //y=1.5
r56 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=15.955 //y=0.62 //x2=15.955 //y2=0.495
r57 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=15.955 //y=0.62 //x2=15.955 //y2=0.885
r58 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.07 //y=0.535 //x2=14.985 //y2=0.495
r59 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.07 //y=0.535 //x2=15.47 //y2=0.535
r60 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.87 //y=0.535 //x2=15.955 //y2=0.495
r61 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.87 //y=0.535 //x2=15.47 //y2=0.535
r62 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=14.985 //y=1.5 //x2=14.985 //y2=1.625
r63 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=14.985 //y=1.5 //x2=14.985 //y2=0.885
r64 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=14.985 //y=0.62 //x2=14.985 //y2=0.495
r65 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=14.985 //y=0.62 //x2=14.985 //y2=0.885
r66 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.1 //y=1.585 //x2=14.015 //y2=1.625
r67 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.1 //y=1.585 //x2=14.5 //y2=1.585
r68 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.9 //y=1.585 //x2=14.985 //y2=1.625
r69 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.9 //y=1.585 //x2=14.5 //y2=1.585
r70 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=14.015 //y=1.5 //x2=14.015 //y2=1.625
r71 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=14.015 //y=1.5 //x2=14.015 //y2=0.885
ends PM_FA\%noxref_22

subckt PM_FA\%noxref_23 ( 7 8 15 16 23 24 25 )
c39 ( 25 0 ) capacitor c=0.0304741f //x=19.055 //y=5.02
c40 ( 24 0 ) capacitor c=0.0185379f //x=18.175 //y=5.02
c41 ( 23 0 ) capacitor c=0.0384176f //x=17.305 //y=5.02
c42 ( 16 0 ) capacitor c=0.00194711f //x=18.405 //y=6.905
c43 ( 15 0 ) capacitor c=0.0131936f //x=19.115 //y=6.905
c44 ( 8 0 ) capacitor c=0.00568107f //x=17.525 //y=5.205
c45 ( 7 0 ) capacitor c=0.0174896f //x=18.235 //y=5.205
r46 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.2 //y=6.82 //x2=19.2 //y2=6.735
r47 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=19.115 //y=6.905 //x2=19.2 //y2=6.82
r48 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=19.115 //y=6.905 //x2=18.405 //y2=6.905
r49 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.32 //y=6.82 //x2=18.405 //y2=6.905
r50 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=18.32 //y=6.82 //x2=18.32 //y2=6.395
r51 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=18.32 //y=5.29 //x2=18.32 //y2=5.715
r52 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.235 //y=5.205 //x2=18.32 //y2=5.29
r53 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=18.235 //y=5.205 //x2=17.525 //y2=5.205
r54 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.44 //y=5.29 //x2=17.525 //y2=5.205
r55 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=17.44 //y=5.29 //x2=17.44 //y2=5.715
ends PM_FA\%noxref_23

subckt PM_FA\%noxref_24 ( 1 5 9 10 13 17 29 )
c50 ( 29 0 ) capacitor c=0.0630989f //x=17.21 //y=0.37
c51 ( 17 0 ) capacitor c=0.00723243f //x=19.285 //y=0.62
c52 ( 13 0 ) capacitor c=0.0149083f //x=19.2 //y=0.535
c53 ( 10 0 ) capacitor c=0.00604817f //x=18.315 //y=1.5
c54 ( 9 0 ) capacitor c=0.00677124f //x=18.315 //y=0.62
c55 ( 5 0 ) capacitor c=0.0245898f //x=18.23 //y=1.585
c56 ( 1 0 ) capacitor c=0.0071362f //x=17.345 //y=1.5
r57 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=19.285 //y=0.62 //x2=19.285 //y2=0.495
r58 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=19.285 //y=0.62 //x2=19.285 //y2=0.885
r59 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.4 //y=0.535 //x2=18.315 //y2=0.495
r60 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.4 //y=0.535 //x2=18.8 //y2=0.535
r61 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.2 //y=0.535 //x2=19.285 //y2=0.495
r62 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.2 //y=0.535 //x2=18.8 //y2=0.535
r63 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=18.315 //y=1.5 //x2=18.315 //y2=1.625
r64 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=18.315 //y=1.5 //x2=18.315 //y2=0.885
r65 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=18.315 //y=0.62 //x2=18.315 //y2=0.495
r66 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=18.315 //y=0.62 //x2=18.315 //y2=0.885
r67 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.43 //y=1.585 //x2=17.345 //y2=1.625
r68 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.43 //y=1.585 //x2=17.83 //y2=1.585
r69 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.23 //y=1.585 //x2=18.315 //y2=1.625
r70 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.23 //y=1.585 //x2=17.83 //y2=1.585
r71 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=17.345 //y=1.5 //x2=17.345 //y2=1.625
r72 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=17.345 //y=1.5 //x2=17.345 //y2=0.885
ends PM_FA\%noxref_24

subckt PM_FA\%noxref_25 ( 1 5 9 10 13 17 29 )
c53 ( 29 0 ) capacitor c=0.0626874f //x=22.76 //y=0.365
c54 ( 17 0 ) capacitor c=0.00722223f //x=24.835 //y=0.615
c55 ( 13 0 ) capacitor c=0.0143165f //x=24.75 //y=0.53
c56 ( 10 0 ) capacitor c=0.00565173f //x=23.865 //y=1.495
c57 ( 9 0 ) capacitor c=0.006761f //x=23.865 //y=0.615
c58 ( 5 0 ) capacitor c=0.0245809f //x=23.78 //y=1.58
c59 ( 1 0 ) capacitor c=0.0071365f //x=22.895 //y=1.495
r60 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=24.835 //y=0.615 //x2=24.835 //y2=0.49
r61 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=24.835 //y=0.615 //x2=24.835 //y2=0.88
r62 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.95 //y=0.53 //x2=23.865 //y2=0.49
r63 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.95 //y=0.53 //x2=24.35 //y2=0.53
r64 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=24.75 //y=0.53 //x2=24.835 //y2=0.49
r65 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=24.75 //y=0.53 //x2=24.35 //y2=0.53
r66 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=23.865 //y=1.495 //x2=23.865 //y2=1.62
r67 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=23.865 //y=1.495 //x2=23.865 //y2=0.88
r68 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=23.865 //y=0.615 //x2=23.865 //y2=0.49
r69 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=23.865 //y=0.615 //x2=23.865 //y2=0.88
r70 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=22.98 //y=1.58 //x2=22.895 //y2=1.62
r71 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.98 //y=1.58 //x2=23.38 //y2=1.58
r72 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.78 //y=1.58 //x2=23.865 //y2=1.62
r73 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.78 //y=1.58 //x2=23.38 //y2=1.58
r74 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=22.895 //y=1.495 //x2=22.895 //y2=1.62
r75 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=22.895 //y=1.495 //x2=22.895 //y2=0.88
ends PM_FA\%noxref_25

subckt PM_FA\%noxref_26 ( 1 5 9 10 13 17 29 )
c57 ( 29 0 ) capacitor c=0.0631306f //x=28.31 //y=0.365
c58 ( 17 0 ) capacitor c=0.00722223f //x=30.385 //y=0.615
c59 ( 13 0 ) capacitor c=0.0143072f //x=30.3 //y=0.53
c60 ( 10 0 ) capacitor c=0.00519634f //x=29.415 //y=1.495
c61 ( 9 0 ) capacitor c=0.006761f //x=29.415 //y=0.615
c62 ( 5 0 ) capacitor c=0.0243504f //x=29.33 //y=1.58
c63 ( 1 0 ) capacitor c=0.0071365f //x=28.445 //y=1.495
r64 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=30.385 //y=0.615 //x2=30.385 //y2=0.49
r65 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=30.385 //y=0.615 //x2=30.385 //y2=0.88
r66 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=29.5 //y=0.53 //x2=29.415 //y2=0.49
r67 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=29.5 //y=0.53 //x2=29.9 //y2=0.53
r68 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=30.3 //y=0.53 //x2=30.385 //y2=0.49
r69 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.3 //y=0.53 //x2=29.9 //y2=0.53
r70 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=29.415 //y=1.495 //x2=29.415 //y2=1.62
r71 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=29.415 //y=1.495 //x2=29.415 //y2=0.88
r72 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=29.415 //y=0.615 //x2=29.415 //y2=0.49
r73 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=29.415 //y=0.615 //x2=29.415 //y2=0.88
r74 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=28.53 //y=1.58 //x2=28.445 //y2=1.62
r75 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=28.53 //y=1.58 //x2=28.93 //y2=1.58
r76 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=29.33 //y=1.58 //x2=29.415 //y2=1.62
r77 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=29.33 //y=1.58 //x2=28.93 //y2=1.58
r78 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=28.445 //y=1.495 //x2=28.445 //y2=1.62
r79 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=28.445 //y=1.495 //x2=28.445 //y2=0.88
ends PM_FA\%noxref_26

subckt PM_FA\%noxref_27 ( 7 8 15 16 23 24 25 )
c42 ( 25 0 ) capacitor c=0.030764f //x=35.705 //y=5.025
c43 ( 24 0 ) capacitor c=0.0185379f //x=34.825 //y=5.025
c44 ( 23 0 ) capacitor c=0.0409962f //x=33.955 //y=5.025
c45 ( 16 0 ) capacitor c=0.00193672f //x=35.055 //y=6.91
c46 ( 15 0 ) capacitor c=0.01354f //x=35.765 //y=6.91
c47 ( 8 0 ) capacitor c=0.0062284f //x=34.175 //y=5.21
c48 ( 7 0 ) capacitor c=0.0182952f //x=34.885 //y=5.21
r49 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.85 //y=6.825 //x2=35.85 //y2=6.74
r50 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=35.765 //y=6.91 //x2=35.85 //y2=6.825
r51 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=35.765 //y=6.91 //x2=35.055 //y2=6.91
r52 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=34.97 //y=6.825 //x2=35.055 //y2=6.91
r53 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=34.97 //y=6.825 //x2=34.97 //y2=6.4
r54 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=34.97 //y=5.295 //x2=34.97 //y2=5.72
r55 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=34.885 //y=5.21 //x2=34.97 //y2=5.295
r56 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=34.885 //y=5.21 //x2=34.175 //y2=5.21
r57 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=34.09 //y=5.295 //x2=34.175 //y2=5.21
r58 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=34.09 //y=5.295 //x2=34.09 //y2=5.72
ends PM_FA\%noxref_27

subckt PM_FA\%COUT ( 1 2 3 4 5 6 7 18 19 20 21 31 33 )
c44 ( 33 0 ) capacitor c=0.028734f //x=37.6 //y=5.02
c45 ( 31 0 ) capacitor c=0.0173218f //x=37.555 //y=0.91
c46 ( 21 0 ) capacitor c=0.00575887f //x=37.83 //y=4.58
c47 ( 20 0 ) capacitor c=0.0136889f //x=38.025 //y=4.58
c48 ( 19 0 ) capacitor c=0.00636159f //x=37.825 //y=2.08
c49 ( 18 0 ) capacitor c=0.0140707f //x=38.025 //y=2.08
c50 ( 1 0 ) capacitor c=0.105613f //x=38.11 //y=2.22
r51 (  20 23 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=38.025 //y=4.58 //x2=38.11 //y2=4.495
r52 (  20 21 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=38.025 //y=4.58 //x2=37.83 //y2=4.58
r53 (  18 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=38.025 //y=2.08 //x2=38.11 //y2=2.165
r54 (  18 19 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=38.025 //y=2.08 //x2=37.825 //y2=2.08
r55 (  12 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=37.745 //y=4.665 //x2=37.83 //y2=4.58
r56 (  12 33 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=37.745 //y=4.665 //x2=37.745 //y2=5.725
r57 (  8 19 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=37.74 //y=1.995 //x2=37.825 //y2=2.08
r58 (  8 31 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=37.74 //y=1.995 //x2=37.74 //y2=1.005
r59 (  7 23 ) resistor r=3.76471 //w=0.187 //l=0.055 //layer=li \
 //thickness=0.1 //x=38.11 //y=4.44 //x2=38.11 //y2=4.495
r60 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=38.11 //y=4.07 //x2=38.11 //y2=4.44
r61 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=38.11 //y=3.7 //x2=38.11 //y2=4.07
r62 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=38.11 //y=3.33 //x2=38.11 //y2=3.7
r63 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=38.11 //y=2.96 //x2=38.11 //y2=3.33
r64 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=38.11 //y=2.59 //x2=38.11 //y2=2.96
r65 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=38.11 //y=2.22 //x2=38.11 //y2=2.59
r66 (  1 22 ) resistor r=3.76471 //w=0.187 //l=0.055 //layer=li \
 //thickness=0.1 //x=38.11 //y=2.22 //x2=38.11 //y2=2.165
ends PM_FA\%COUT

