magic
tech sky130A
magscale 1 2
timestamp 1652327672
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 205 871 239 905
rect 353 871 387 905
rect 501 871 535 905
rect 205 797 239 831
rect 353 797 387 831
rect 501 797 535 831
rect 205 723 239 757
rect 353 723 387 757
rect 501 723 535 757
rect 205 649 239 683
rect 353 649 387 683
rect 501 649 535 683
rect 205 575 239 609
rect 353 575 387 609
rect 501 575 535 609
rect 205 501 239 535
rect 353 501 387 535
rect 501 501 535 535
rect 205 427 239 461
rect 353 427 387 461
rect 501 427 535 461
<< metal1 >>
rect -34 1446 700 1514
rect -34 -34 700 34
use nor2x1_pcell  nor2x1_pcell_0 pcells
timestamp 1652323563
transform 1 0 0 0 1 0
box -87 -34 753 1550
<< labels >>
rlabel locali 501 427 535 461 1 Y
port 1 nsew signal output
rlabel locali 501 501 535 535 1 Y
port 1 nsew signal output
rlabel locali 501 575 535 609 1 Y
port 1 nsew signal output
rlabel locali 501 649 535 683 1 Y
port 1 nsew signal output
rlabel locali 501 723 535 757 1 Y
port 1 nsew signal output
rlabel locali 501 797 535 831 1 Y
port 1 nsew signal output
rlabel locali 501 871 535 905 1 Y
port 1 nsew signal output
rlabel locali 205 427 239 461 1 A
port 2 nsew signal input
rlabel locali 205 501 239 535 1 A
port 2 nsew signal input
rlabel locali 205 575 239 609 1 A
port 2 nsew signal input
rlabel locali 205 649 239 683 1 A
port 2 nsew signal input
rlabel locali 205 723 239 757 1 A
port 2 nsew signal input
rlabel locali 205 797 239 831 1 A
port 2 nsew signal input
rlabel locali 205 871 239 905 1 A
port 2 nsew signal input
rlabel locali 353 427 387 461 1 B
port 3 nsew signal input
rlabel locali 353 501 387 535 1 B
port 3 nsew signal input
rlabel locali 353 575 387 609 1 B
port 3 nsew signal input
rlabel locali 353 649 387 683 1 B
port 3 nsew signal input
rlabel locali 353 723 387 757 1 B
port 3 nsew signal input
rlabel locali 353 797 387 831 1 B
port 3 nsew signal input
rlabel locali 353 871 387 905 1 B
port 3 nsew signal input
rlabel metal1 -34 1446 700 1514 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 -34 -34 700 34 1 GND
port 5 nsew power bidirectional abutment


<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 666 1480
string LEFsymmetry X Y R90
<< end >>
