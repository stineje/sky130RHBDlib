* SPICE3 file created from AOI3X1.ext - technology: sky130A

.subckt AOI3X1 YN A B C VPB VNB
M1000 VNB a_168_157# a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=2.1157p pd=14.51u as=0p ps=0u
M1001 VPB.t3 a_168_157# a_217_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPB.t5 a_217_1004.t5 a_797_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t1 a_343_383# a_217_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_797_1005.t1 a_1009_383# a_864_181.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_217_1004.t4 a_168_157# VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_217_1004.t2 a_343_383# VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_797_1005.t2 a_217_1004.t6 VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_864_181.t1 a_1009_383# a_797_1005.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 a_168_157# VPB 0.08fF
C1 a_168_157# a_343_383# 0.26fF
C2 VPB a_1009_383# 0.07fF
C3 VPB a_343_383# 0.07fF
R0 a_217_1004.n4 a_217_1004.t6 486.819
R1 a_217_1004.n4 a_217_1004.t5 384.527
R2 a_217_1004.n6 a_217_1004.n3 215.652
R3 a_217_1004.n5 a_217_1004.t7 207.443
R4 a_217_1004.n5 a_217_1004.n4 169.7
R5 a_217_1004.n6 a_217_1004.n5 153.315
R6 a_217_1004.n8 a_217_1004.n6 140.981
R7 a_217_1004.n3 a_217_1004.n2 76.002
R8 a_217_1004.n8 a_217_1004.n7 30
R9 a_217_1004.n9 a_217_1004.n0 24.383
R10 a_217_1004.n9 a_217_1004.n8 23.684
R11 a_217_1004.n1 a_217_1004.t1 14.282
R12 a_217_1004.n1 a_217_1004.t2 14.282
R13 a_217_1004.n2 a_217_1004.t3 14.282
R14 a_217_1004.n2 a_217_1004.t4 14.282
R15 a_217_1004.n3 a_217_1004.n1 12.85
R16 VPB VPB.n137 126.832
R17 VPB.n115 VPB.n113 94.117
R18 VPB.n121 VPB.n120 76
R19 VPB.n130 VPB.n129 76
R20 VPB.n75 VPB.n74 61.764
R21 VPB.n91 VPB.t2 55.106
R22 VPB.n109 VPB.t1 55.106
R23 VPB.n106 VPB.n105 48.952
R24 VPB.n63 VPB.n62 44.502
R25 VPB.n93 VPB.n92 44.502
R26 VPB.n61 VPB.n22 41.183
R27 VPB.n100 VPB.n90 40.824
R28 VPB.n134 VPB.n130 20.452
R29 VPB.n46 VPB.n43 20.452
R30 VPB.n102 VPB.n101 17.801
R31 VPB.n90 VPB.t0 14.282
R32 VPB.n90 VPB.t3 14.282
R33 VPB.n22 VPB.t4 14.282
R34 VPB.n22 VPB.t5 14.282
R35 VPB.n46 VPB.n45 13.653
R36 VPB.n45 VPB.n44 13.653
R37 VPB.n50 VPB.n49 13.653
R38 VPB.n49 VPB.n48 13.653
R39 VPB.n53 VPB.n52 13.653
R40 VPB.n52 VPB.n51 13.653
R41 VPB.n56 VPB.n55 13.653
R42 VPB.n55 VPB.n54 13.653
R43 VPB.n60 VPB.n59 13.653
R44 VPB.n59 VPB.n58 13.653
R45 VPB.n65 VPB.n64 13.653
R46 VPB.n64 VPB.n63 13.653
R47 VPB.n68 VPB.n67 13.653
R48 VPB.n67 VPB.n66 13.653
R49 VPB.n120 VPB.n119 13.653
R50 VPB.n119 VPB.n118 13.653
R51 VPB.n116 VPB.n115 13.653
R52 VPB.n115 VPB.n114 13.653
R53 VPB.n112 VPB.n111 13.653
R54 VPB.n111 VPB.n110 13.653
R55 VPB.n108 VPB.n107 13.653
R56 VPB.n107 VPB.n106 13.653
R57 VPB.n104 VPB.n103 13.653
R58 VPB.n103 VPB.n102 13.653
R59 VPB.n99 VPB.n98 13.653
R60 VPB.n98 VPB.n97 13.653
R61 VPB.n95 VPB.n94 13.653
R62 VPB.n94 VPB.n93 13.653
R63 VPB.n16 VPB.n15 13.653
R64 VPB.n15 VPB.n14 13.653
R65 VPB.n130 VPB.n0 13.653
R66 VPB VPB.n0 13.653
R67 VPB.n58 VPB.n57 13.35
R68 VPB.n97 VPB.n96 13.35
R69 VPB.n134 VPB.n133 13.276
R70 VPB.n133 VPB.n131 13.276
R71 VPB.n89 VPB.n71 13.276
R72 VPB.n71 VPB.n69 13.276
R73 VPB.n53 VPB.n50 13.276
R74 VPB.n56 VPB.n53 13.276
R75 VPB.n60 VPB.n56 13.276
R76 VPB.n68 VPB.n65 13.276
R77 VPB.n120 VPB.n68 13.276
R78 VPB.n120 VPB.n117 13.276
R79 VPB.n117 VPB.n116 13.276
R80 VPB.n116 VPB.n112 13.276
R81 VPB.n108 VPB.n104 13.276
R82 VPB.n99 VPB.n95 13.276
R83 VPB.n130 VPB.n16 13.276
R84 VPB.n43 VPB.n25 13.276
R85 VPB.n25 VPB.n23 13.276
R86 VPB.n30 VPB.n28 12.796
R87 VPB.n30 VPB.n29 12.564
R88 VPB.n39 VPB.n38 12.198
R89 VPB.n36 VPB.n35 12.198
R90 VPB.n36 VPB.n33 12.198
R91 VPB.n109 VPB.n108 11.841
R92 VPB.n95 VPB.n91 11.482
R93 VPB.n61 VPB.n60 8.97
R94 VPB.n43 VPB.n42 7.5
R95 VPB.n28 VPB.n27 7.5
R96 VPB.n35 VPB.n34 7.5
R97 VPB.n33 VPB.n32 7.5
R98 VPB.n25 VPB.n24 7.5
R99 VPB.n40 VPB.n26 7.5
R100 VPB.n71 VPB.n70 7.5
R101 VPB.n84 VPB.n83 7.5
R102 VPB.n78 VPB.n77 7.5
R103 VPB.n80 VPB.n79 7.5
R104 VPB.n73 VPB.n72 7.5
R105 VPB.n89 VPB.n88 7.5
R106 VPB.n133 VPB.n132 7.5
R107 VPB.n12 VPB.n11 7.5
R108 VPB.n6 VPB.n5 7.5
R109 VPB.n8 VPB.n7 7.5
R110 VPB.n2 VPB.n1 7.5
R111 VPB.n135 VPB.n134 7.5
R112 VPB.n117 VPB.n89 7.176
R113 VPB.n100 VPB.n99 6.817
R114 VPB.n85 VPB.n82 6.729
R115 VPB.n81 VPB.n78 6.729
R116 VPB.n76 VPB.n73 6.729
R117 VPB.n13 VPB.n10 6.729
R118 VPB.n9 VPB.n6 6.729
R119 VPB.n4 VPB.n2 6.729
R120 VPB.n76 VPB.n75 6.728
R121 VPB.n81 VPB.n80 6.728
R122 VPB.n85 VPB.n84 6.728
R123 VPB.n88 VPB.n87 6.728
R124 VPB.n4 VPB.n3 6.728
R125 VPB.n9 VPB.n8 6.728
R126 VPB.n13 VPB.n12 6.728
R127 VPB.n136 VPB.n135 6.728
R128 VPB.n104 VPB.n100 6.458
R129 VPB.n42 VPB.n41 6.398
R130 VPB.n47 VPB.n46 6.112
R131 VPB.n50 VPB.n47 6.101
R132 VPB.n65 VPB.n61 4.305
R133 VPB.n91 VPB.n16 1.794
R134 VPB.n112 VPB.n109 1.435
R135 VPB.n40 VPB.n31 1.402
R136 VPB.n40 VPB.n36 1.402
R137 VPB.n40 VPB.n37 1.402
R138 VPB.n40 VPB.n39 1.402
R139 VPB.n41 VPB.n40 0.735
R140 VPB.n40 VPB.n30 0.735
R141 VPB.n86 VPB.n85 0.387
R142 VPB.n86 VPB.n81 0.387
R143 VPB.n86 VPB.n76 0.387
R144 VPB.n87 VPB.n86 0.387
R145 VPB.n137 VPB.n13 0.387
R146 VPB.n137 VPB.n9 0.387
R147 VPB.n137 VPB.n4 0.387
R148 VPB.n137 VPB.n136 0.387
R149 VPB.n129 VPB 0.198
R150 VPB.n18 VPB.n17 0.136
R151 VPB.n19 VPB.n18 0.136
R152 VPB.n20 VPB.n19 0.136
R153 VPB.n21 VPB.n20 0.136
R154 VPB.n121 VPB.n21 0.136
R155 VPB VPB.n121 0.136
R156 VPB.n122 VPB 0.136
R157 VPB.n123 VPB.n122 0.136
R158 VPB.n124 VPB.n123 0.136
R159 VPB.n125 VPB.n124 0.136
R160 VPB.n126 VPB.n125 0.136
R161 VPB.n127 VPB.n126 0.136
R162 VPB.n128 VPB.n127 0.136
R163 VPB.n129 VPB.n128 0.136
R164 a_797_1005.n0 a_797_1005.t1 101.66
R165 a_797_1005.n0 a_797_1005.t3 101.66
R166 a_797_1005.n0 a_797_1005.t0 14.294
R167 a_797_1005.t2 a_797_1005.n0 14.282
R168 a_112_73.t0 a_112_73.n1 93.333
R169 a_112_73.n4 a_112_73.n2 55.07
R170 a_112_73.t0 a_112_73.n0 8.137
R171 a_112_73.n4 a_112_73.n3 4.619
R172 a_112_73.t0 a_112_73.n4 0.071
R173 VNB VNB.n138 300.778
R174 VNB.n85 VNB.n84 199.897
R175 VNB.n110 VNB.n108 154.509
R176 VNB.n61 VNB.n60 121.366
R177 VNB.n95 VNB.n91 84.842
R178 VNB.n125 VNB.n124 76
R179 VNB.n116 VNB.n115 76
R180 VNB.n14 VNB.t2 39.412
R181 VNB.n55 VNB.n54 36.937
R182 VNB.n56 VNB.n55 36.937
R183 VNB.n62 VNB.n61 36.937
R184 VNB.n93 VNB.n92 36.678
R185 VNB.n68 VNB.n67 27.855
R186 VNB.n44 VNB.n41 20.452
R187 VNB.n126 VNB.n125 20.452
R188 VNB.n65 VNB.n17 19.735
R189 VNB.n59 VNB.n21 19.735
R190 VNB.n52 VNB.n23 19.735
R191 VNB.n45 VNB.n26 19.735
R192 VNB.n74 VNB.n15 19.735
R193 VNB.n14 VNB.n13 17.185
R194 VNB.n25 VNB.n24 17.006
R195 VNB.n69 VNB.n68 16.721
R196 VNB.n20 VNB.t0 13.654
R197 VNB.n20 VNB.n19 13.654
R198 VNB.n48 VNB.n47 13.653
R199 VNB.n47 VNB.n46 13.653
R200 VNB.n51 VNB.n50 13.653
R201 VNB.n50 VNB.n49 13.653
R202 VNB.n58 VNB.n57 13.653
R203 VNB.n57 VNB.n56 13.653
R204 VNB.n64 VNB.n63 13.653
R205 VNB.n63 VNB.n62 13.653
R206 VNB.n70 VNB.n69 13.653
R207 VNB.n73 VNB.n72 13.653
R208 VNB.n72 VNB.n71 13.653
R209 VNB.n115 VNB.n114 13.653
R210 VNB.n114 VNB.n113 13.653
R211 VNB.n111 VNB.n110 13.653
R212 VNB.n110 VNB.n109 13.653
R213 VNB.n107 VNB.n106 13.653
R214 VNB.n106 VNB.n105 13.653
R215 VNB.n104 VNB.n103 13.653
R216 VNB.n103 VNB.n102 13.653
R217 VNB.n101 VNB.n100 13.653
R218 VNB.n100 VNB.n99 13.653
R219 VNB.n98 VNB.n97 13.653
R220 VNB.n97 VNB.n96 13.653
R221 VNB.n94 VNB.n93 13.653
R222 VNB.n6 VNB.n5 13.653
R223 VNB.n5 VNB.n4 13.653
R224 VNB.n125 VNB.n0 13.653
R225 VNB VNB.n0 13.653
R226 VNB.n44 VNB.n43 13.653
R227 VNB.n43 VNB.n42 13.653
R228 VNB.n133 VNB.n130 13.577
R229 VNB.n29 VNB.n27 13.276
R230 VNB.n41 VNB.n29 13.276
R231 VNB.n77 VNB.n75 13.276
R232 VNB.n90 VNB.n77 13.276
R233 VNB.n51 VNB.n48 13.276
R234 VNB.n73 VNB.n70 13.276
R235 VNB.n115 VNB.n112 13.276
R236 VNB.n112 VNB.n111 13.276
R237 VNB.n111 VNB.n107 13.276
R238 VNB.n107 VNB.n104 13.276
R239 VNB.n104 VNB.n101 13.276
R240 VNB.n101 VNB.n98 13.276
R241 VNB.n94 VNB.n6 13.276
R242 VNB.n125 VNB.n6 13.276
R243 VNB.n3 VNB.n1 13.276
R244 VNB.n126 VNB.n3 13.276
R245 VNB.n45 VNB.n44 11.661
R246 VNB.n115 VNB.n74 11.661
R247 VNB.n58 VNB.n52 10.764
R248 VNB.n65 VNB.n64 10.764
R249 VNB.n98 VNB.n95 10.764
R250 VNB.n23 VNB.n22 7.5
R251 VNB.n17 VNB.n16 7.5
R252 VNB.n135 VNB.n134 7.5
R253 VNB.n83 VNB.n82 7.5
R254 VNB.n79 VNB.n78 7.5
R255 VNB.n77 VNB.n76 7.5
R256 VNB.n90 VNB.n89 7.5
R257 VNB.n127 VNB.n126 7.5
R258 VNB.n3 VNB.n2 7.5
R259 VNB.n132 VNB.n131 7.5
R260 VNB.n35 VNB.n34 7.5
R261 VNB.n31 VNB.n30 7.5
R262 VNB.n29 VNB.n28 7.5
R263 VNB.n41 VNB.n40 7.5
R264 VNB.n112 VNB.n90 7.176
R265 VNB.t0 VNB.n18 7.04
R266 VNB.n137 VNB.n135 7.011
R267 VNB.n86 VNB.n83 7.011
R268 VNB.n81 VNB.n79 7.011
R269 VNB.n37 VNB.n35 7.011
R270 VNB.n33 VNB.n31 7.011
R271 VNB.n89 VNB.n88 7.01
R272 VNB.n81 VNB.n80 7.01
R273 VNB.n86 VNB.n85 7.01
R274 VNB.n40 VNB.n39 7.01
R275 VNB.n33 VNB.n32 7.01
R276 VNB.n37 VNB.n36 7.01
R277 VNB.n137 VNB.n136 7.01
R278 VNB.n133 VNB.n132 6.788
R279 VNB.n128 VNB.n127 6.788
R280 VNB.n59 VNB.n58 6.638
R281 VNB.n64 VNB.n59 6.638
R282 VNB.n26 VNB.n25 6.323
R283 VNB.n15 VNB.n14 6.139
R284 VNB.n21 VNB.n20 5.774
R285 VNB.n54 VNB.n53 5.276
R286 VNB.n52 VNB.n51 2.511
R287 VNB.n70 VNB.n65 2.511
R288 VNB.n95 VNB.n94 2.511
R289 VNB.n68 VNB.n66 1.99
R290 VNB.n48 VNB.n45 1.614
R291 VNB.n74 VNB.n73 1.614
R292 VNB.n138 VNB.n129 0.921
R293 VNB.n138 VNB.n133 0.476
R294 VNB.n138 VNB.n128 0.475
R295 VNB.n87 VNB.n81 0.246
R296 VNB.n88 VNB.n87 0.246
R297 VNB.n87 VNB.n86 0.246
R298 VNB.n38 VNB.n33 0.246
R299 VNB.n39 VNB.n38 0.246
R300 VNB.n38 VNB.n37 0.246
R301 VNB.n138 VNB.n137 0.246
R302 VNB.n124 VNB 0.198
R303 VNB.n8 VNB.n7 0.136
R304 VNB.n9 VNB.n8 0.136
R305 VNB.n10 VNB.n9 0.136
R306 VNB.n11 VNB.n10 0.136
R307 VNB.n12 VNB.n11 0.136
R308 VNB.n116 VNB.n12 0.136
R309 VNB VNB.n116 0.136
R310 VNB.n117 VNB 0.136
R311 VNB.n118 VNB.n117 0.136
R312 VNB.n119 VNB.n118 0.136
R313 VNB.n120 VNB.n119 0.136
R314 VNB.n121 VNB.n120 0.136
R315 VNB.n122 VNB.n121 0.136
R316 VNB.n123 VNB.n122 0.136
R317 VNB.n124 VNB.n123 0.136
R318 a_864_181.n4 a_864_181.n0 321.065
R319 a_864_181.n4 a_864_181.n3 133.539
R320 a_864_181.n6 a_864_181.n4 55.263
R321 a_864_181.n3 a_864_181.n2 22.578
R322 a_864_181.n6 a_864_181.n5 15.001
R323 a_864_181.n0 a_864_181.t2 14.282
R324 a_864_181.n0 a_864_181.t1 14.282
R325 a_864_181.n7 a_864_181.n6 12.632
R326 a_864_181.n3 a_864_181.n1 8.58
C4 VPB VNB 6.16fF
C5 a_864_181.n0 VNB 0.85fF
C6 a_864_181.n1 VNB 0.04fF
C7 a_864_181.n2 VNB 0.05fF
C8 a_864_181.n3 VNB 0.19fF
C9 a_864_181.n4 VNB 0.62fF
C10 a_864_181.n5 VNB 0.08fF
C11 a_864_181.n6 VNB 0.08fF
C12 a_864_181.n7 VNB 0.05fF
C13 a_112_73.n0 VNB 0.05fF
C14 a_112_73.n1 VNB 0.02fF
C15 a_112_73.n2 VNB 0.12fF
C16 a_112_73.n3 VNB 0.04fF
C17 a_112_73.n4 VNB 0.16fF
C18 a_797_1005.n0 VNB 0.52fF
C19 VPB.n0 VNB 0.03fF
C20 VPB.n1 VNB 0.03fF
C21 VPB.n2 VNB 0.02fF
C22 VPB.n3 VNB 0.13fF
C23 VPB.n5 VNB 0.02fF
C24 VPB.n6 VNB 0.02fF
C25 VPB.n7 VNB 0.02fF
C26 VPB.n8 VNB 0.02fF
C27 VPB.n10 VNB 0.02fF
C28 VPB.n11 VNB 0.02fF
C29 VPB.n12 VNB 0.02fF
C30 VPB.n14 VNB 0.23fF
C31 VPB.n15 VNB 0.02fF
C32 VPB.n16 VNB 0.01fF
C33 VPB.n17 VNB 0.09fF
C34 VPB.n18 VNB 0.02fF
C35 VPB.n19 VNB 0.02fF
C36 VPB.n20 VNB 0.02fF
C37 VPB.n21 VNB 0.02fF
C38 VPB.n22 VNB 0.10fF
C39 VPB.n23 VNB 0.02fF
C40 VPB.n24 VNB 0.02fF
C41 VPB.n25 VNB 0.02fF
C42 VPB.n26 VNB 0.13fF
C43 VPB.n27 VNB 0.03fF
C44 VPB.n28 VNB 0.02fF
C45 VPB.n29 VNB 0.04fF
C46 VPB.n30 VNB 0.01fF
C47 VPB.n32 VNB 0.02fF
C48 VPB.n33 VNB 0.02fF
C49 VPB.n34 VNB 0.02fF
C50 VPB.n35 VNB 0.02fF
C51 VPB.n38 VNB 0.02fF
C52 VPB.n40 VNB 0.44fF
C53 VPB.n42 VNB 0.03fF
C54 VPB.n43 VNB 0.04fF
C55 VPB.n44 VNB 0.26fF
C56 VPB.n45 VNB 0.03fF
C57 VPB.n46 VNB 0.03fF
C58 VPB.n47 VNB 0.00fF
C59 VPB.n48 VNB 0.26fF
C60 VPB.n49 VNB 0.02fF
C61 VPB.n50 VNB 0.02fF
C62 VPB.n51 VNB 0.26fF
C63 VPB.n52 VNB 0.02fF
C64 VPB.n53 VNB 0.02fF
C65 VPB.n54 VNB 0.26fF
C66 VPB.n55 VNB 0.02fF
C67 VPB.n56 VNB 0.02fF
C68 VPB.n57 VNB 0.13fF
C69 VPB.n58 VNB 0.14fF
C70 VPB.n59 VNB 0.02fF
C71 VPB.n60 VNB 0.02fF
C72 VPB.n61 VNB 0.02fF
C73 VPB.n62 VNB 0.13fF
C74 VPB.n63 VNB 0.15fF
C75 VPB.n64 VNB 0.02fF
C76 VPB.n65 VNB 0.02fF
C77 VPB.n66 VNB 0.23fF
C78 VPB.n67 VNB 0.02fF
C79 VPB.n68 VNB 0.02fF
C80 VPB.n69 VNB 0.02fF
C81 VPB.n70 VNB 0.02fF
C82 VPB.n71 VNB 0.02fF
C83 VPB.n72 VNB 0.03fF
C84 VPB.n73 VNB 0.02fF
C85 VPB.n74 VNB 0.20fF
C86 VPB.n75 VNB 0.04fF
C87 VPB.n77 VNB 0.02fF
C88 VPB.n78 VNB 0.02fF
C89 VPB.n79 VNB 0.02fF
C90 VPB.n80 VNB 0.02fF
C91 VPB.n82 VNB 0.02fF
C92 VPB.n83 VNB 0.02fF
C93 VPB.n84 VNB 0.02fF
C94 VPB.n86 VNB 0.26fF
C95 VPB.n88 VNB 0.02fF
C96 VPB.n89 VNB 0.02fF
C97 VPB.n90 VNB 0.10fF
C98 VPB.n91 VNB 0.06fF
C99 VPB.n92 VNB 0.13fF
C100 VPB.n93 VNB 0.15fF
C101 VPB.n94 VNB 0.02fF
C102 VPB.n95 VNB 0.02fF
C103 VPB.n96 VNB 0.13fF
C104 VPB.n97 VNB 0.14fF
C105 VPB.n98 VNB 0.02fF
C106 VPB.n99 VNB 0.02fF
C107 VPB.n100 VNB 0.02fF
C108 VPB.n101 VNB 0.13fF
C109 VPB.n102 VNB 0.14fF
C110 VPB.n103 VNB 0.02fF
C111 VPB.n104 VNB 0.02fF
C112 VPB.n105 VNB 0.13fF
C113 VPB.n106 VNB 0.15fF
C114 VPB.n107 VNB 0.02fF
C115 VPB.n108 VNB 0.02fF
C116 VPB.n109 VNB 0.05fF
C117 VPB.n110 VNB 0.22fF
C118 VPB.n111 VNB 0.02fF
C119 VPB.n112 VNB 0.01fF
C120 VPB.n113 VNB 0.03fF
C121 VPB.n114 VNB 0.26fF
C122 VPB.n115 VNB 0.01fF
C123 VPB.n116 VNB 0.02fF
C124 VPB.n117 VNB 0.03fF
C125 VPB.n118 VNB 0.26fF
C126 VPB.n119 VNB 0.01fF
C127 VPB.n120 VNB 0.02fF
C128 VPB.n121 VNB 0.02fF
C129 VPB.n122 VNB 0.02fF
C130 VPB.n123 VNB 0.02fF
C131 VPB.n124 VNB 0.02fF
C132 VPB.n125 VNB 0.02fF
C133 VPB.n126 VNB 0.02fF
C134 VPB.n127 VNB 0.02fF
C135 VPB.n128 VNB 0.02fF
C136 VPB.n129 VNB 0.03fF
C137 VPB.n130 VNB 0.03fF
C138 VPB.n131 VNB 0.02fF
C139 VPB.n132 VNB 0.02fF
C140 VPB.n133 VNB 0.02fF
C141 VPB.n134 VNB 0.04fF
C142 VPB.n135 VNB 0.03fF
C143 VPB.n137 VNB 0.41fF
C144 a_217_1004.n0 VNB 0.03fF
C145 a_217_1004.n1 VNB 0.43fF
C146 a_217_1004.n2 VNB 0.51fF
C147 a_217_1004.n3 VNB 0.31fF
C148 a_217_1004.n4 VNB 0.35fF
C149 a_217_1004.t7 VNB 0.38fF
C150 a_217_1004.n5 VNB 0.45fF
C151 a_217_1004.n6 VNB 0.48fF
C152 a_217_1004.n7 VNB 0.03fF
C153 a_217_1004.n8 VNB 0.17fF
C154 a_217_1004.n9 VNB 0.04fF
.ends
