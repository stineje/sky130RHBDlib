* SPICE3 file created from AOA4X1.ext - technology: sky130A

.subckt AOA4X1 Y A B C D VDD GND
X0 a_864_181 a_217_1004 GND GND nshort w=3 l=0.15
X1 VDD B a_217_1004 VDD pshort w=2 l=0.15 M=2
X2 GND A a_112_73 GND nshort w=3 l=0.15
X3 GND a_864_181 a_1444_73 GND nshort w=3 l=0.15
X4 VDD a_864_181 a_1549_1004 VDD pshort w=2 l=0.15 M=2
X5 a_1549_1004 D a_1444_73 GND nshort w=3 l=0.15
X6 VDD a_1549_1004 Y VDD pshort w=2 l=0.15 M=2
X7 a_797_1005 C a_864_181 VDD pshort w=2 l=0.15 M=2
X8 a_217_1004 A VDD VDD pshort w=2 l=0.15 M=2
X9 a_217_1004 B a_112_73 GND nshort w=3 l=0.15
X10 VDD D a_1549_1004 VDD pshort w=2 l=0.15 M=2
X11 a_864_181 C GND GND nshort w=3 l=0.15
X12 a_797_1005 a_217_1004 VDD VDD pshort w=2 l=0.15 M=2
X13 Y a_1549_1004 GND GND nshort w=3 l=0.15
C0 VDD GND 6.16fF
.ends
