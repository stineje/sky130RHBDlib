* SPICE3 file created from AND2X1.ext - technology: sky130A

.subckt AND2X1 Y A B VPB VNB
X0 VPB a_343_383# a_217_1004# VPB sky130_fd_pr__pfet_01v8 ad=2.78e+12p pd=2.278e+07u as=0p ps=0u w=2e+06u l=150000u M=2
X1 VNB a_168_157# a_112_73# VNB sky130_fd_pr__nfet_01v8 ad=1.3199e+12p pd=9.67e+06u as=0p ps=0u w=3e+06u l=150000u
X2 a_851_182# a_217_1004# VNB VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X3 VPB a_217_1004# a_851_182# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X4 a_217_1004# a_168_157# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X5 a_217_1004# a_343_383# a_112_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
.ends
