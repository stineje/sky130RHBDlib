* SPICE3 file created from DFFSNRNQX1.ext - technology: sky130A

.subckt DFFSNRNQX1 Q D CLK SN RN VDD GND
M1000 VDD.t32 a_2201_1050.t7 a_1561_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 Q.t1 SN.t0 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t6 D.t0 a_277_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 GND D.t1 a_91_103.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1004 a_599_989.t1 CLK.t1 VDD.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VDD.t5 a_277_1050.t7 a_2201_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VDD.t13 CLK.t2 a_1561_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VDD.t9 RN.t0 a_277_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_599_989.t6 a_1561_989.t7 VDD.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VDD.t2 RN.t1 a_1561_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VDD.t17 SN.t1 a_2201_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_4125_1050.t1 a_599_989.t8 VDD.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_4125_1050.t6 Q.t7 VDD.t33 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1561_989.t2 CLK.t3 VDD.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t0 a_599_989.t9 a_277_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 GND a_277_1050.t9 a_2015_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1016 VDD.t29 a_1561_989.t8 a_2201_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_4125_1050.t3 RN.t2 VDD.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_1561_989.t12 a_5182_210.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1019 a_1561_989.t5 a_2201_1050.t8 VDD.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 VDD.t21 a_4125_1050.t8 Q.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_277_1050.t5 D.t2 VDD.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 GND a_2201_1050.t9 a_2977_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1023 VDD.t35 a_277_1050.t8 a_599_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 GND a_277_1050.t10 a_1053_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1025 VDD.t26 a_1561_989.t11 a_599_989.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VDD.t23 SN.t2 Q.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_277_1050.t4 RN.t5 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 GND a_599_989.t11 a_3939_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1029 VDD.t10 CLK.t4 a_599_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1561_989.t4 RN.t6 VDD.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 VDD.t30 a_1561_989.t13 Q.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_599_989.t2 a_277_1050.t11 VDD.t34 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_2201_1050.t0 SN.t3 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 VDD.t14 RN.t7 a_4125_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_277_1050.t2 a_599_989.t10 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 GND a_4125_1050.t7 a_4901_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_2201_1050.t4 a_277_1050.t12 VDD.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_2201_1050.t6 a_1561_989.t14 VDD.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 VDD.t24 a_599_989.t12 a_4125_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 VDD.t4 Q.t9 a_4125_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 Q.t2 a_4125_1050.t9 VDD.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 Q.t5 a_1561_989.t15 VDD.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 D RN 0.18fF
C1 CLK SN 0.48fF
C2 VDD CLK 0.10fF
C3 SN Q 0.39fF
C4 VDD SN 0.10fF
C5 RN CLK 0.73fF
C6 VDD Q 1.83fF
C7 RN SN 0.37fF
C8 VDD D 0.08fF
C9 RN Q 0.18fF
C10 VDD RN 2.04fF
R0 CLK.n2 CLK.t4 479.223
R1 CLK.n0 CLK.t2 479.223
R2 CLK.n2 CLK.t1 375.52
R3 CLK.n0 CLK.t3 375.52
R4 CLK.n3 CLK.t5 215.154
R5 CLK.n1 CLK.t0 215.154
R6 CLK.n3 CLK.n2 122.323
R7 CLK.n1 CLK.n0 122.323
R8 CLK.n4 CLK.n1 83.028
R9 CLK.n4 CLK.n3 76
R10 CLK.n4 CLK 0.046
R11 a_2977_103.t0 a_2977_103.n0 117.777
R12 a_2977_103.n2 a_2977_103.n1 55.228
R13 a_2977_103.n4 a_2977_103.n3 9.111
R14 a_2977_103.n8 a_2977_103.n6 7.859
R15 a_2977_103.t0 a_2977_103.n2 4.04
R16 a_2977_103.t0 a_2977_103.n8 3.034
R17 a_2977_103.n6 a_2977_103.n4 1.964
R18 a_2977_103.n6 a_2977_103.n5 1.964
R19 a_2977_103.n8 a_2977_103.n7 0.443
R20 a_3258_210.n12 a_3258_210.n5 96.467
R21 a_3258_210.t0 a_3258_210.n1 46.91
R22 a_3258_210.n9 a_3258_210.n7 34.805
R23 a_3258_210.n9 a_3258_210.n8 32.622
R24 a_3258_210.t0 a_3258_210.n12 32.417
R25 a_3258_210.n5 a_3258_210.n4 22.349
R26 a_3258_210.n11 a_3258_210.n9 19.017
R27 a_3258_210.n1 a_3258_210.n0 17.006
R28 a_3258_210.n5 a_3258_210.n3 8.443
R29 a_3258_210.t0 a_3258_210.n2 8.137
R30 a_3258_210.n7 a_3258_210.n6 7.5
R31 a_3258_210.n11 a_3258_210.n10 7.5
R32 a_3258_210.n12 a_3258_210.n11 1.435
R33 a_4125_1050.n5 a_4125_1050.t8 512.525
R34 a_4125_1050.n5 a_4125_1050.t9 371.139
R35 a_4125_1050.n6 a_4125_1050.t7 261.115
R36 a_4125_1050.n7 a_4125_1050.n4 197.352
R37 a_4125_1050.n9 a_4125_1050.n7 193.073
R38 a_4125_1050.n6 a_4125_1050.n5 189.266
R39 a_4125_1050.n7 a_4125_1050.n6 153.315
R40 a_4125_1050.n3 a_4125_1050.n2 79.232
R41 a_4125_1050.n4 a_4125_1050.n3 63.152
R42 a_4125_1050.n4 a_4125_1050.n0 16.08
R43 a_4125_1050.n3 a_4125_1050.n1 16.08
R44 a_4125_1050.n9 a_4125_1050.n8 15.218
R45 a_4125_1050.n0 a_4125_1050.t0 14.282
R46 a_4125_1050.n0 a_4125_1050.t6 14.282
R47 a_4125_1050.n1 a_4125_1050.t2 14.282
R48 a_4125_1050.n1 a_4125_1050.t3 14.282
R49 a_4125_1050.n2 a_4125_1050.t4 14.282
R50 a_4125_1050.n2 a_4125_1050.t1 14.282
R51 a_4125_1050.n10 a_4125_1050.n9 12.014
R52 a_4901_103.t0 a_4901_103.n0 117.777
R53 a_4901_103.n2 a_4901_103.n1 55.228
R54 a_4901_103.n4 a_4901_103.n3 9.111
R55 a_4901_103.t0 a_4901_103.n2 4.04
R56 a_4901_103.n8 a_4901_103.n7 2.455
R57 a_4901_103.n6 a_4901_103.n4 1.964
R58 a_4901_103.n6 a_4901_103.n5 1.964
R59 a_4901_103.n8 a_4901_103.n6 0.636
R60 a_4901_103.t0 a_4901_103.n8 0.246
R61 GND.n38 GND.n36 219.745
R62 GND.n161 GND.n160 219.745
R63 GND.n203 GND.n201 219.745
R64 GND.n241 GND.n239 219.745
R65 GND.n80 GND.n79 219.745
R66 GND.n27 GND.n26 85.559
R67 GND.n69 GND.n68 85.559
R68 GND.n111 GND.n110 85.559
R69 GND.n212 GND.n211 85.559
R70 GND.n170 GND.n169 85.559
R71 GND.n128 GND.n127 85.559
R72 GND.n38 GND.n37 85.529
R73 GND.n161 GND.n159 85.529
R74 GND.n203 GND.n202 85.529
R75 GND.n241 GND.n240 85.529
R76 GND.n80 GND.n78 85.529
R77 GND.n122 GND.n121 76
R78 GND.n12 GND.n11 76
R79 GND.n15 GND.n14 76
R80 GND.n18 GND.n17 76
R81 GND.n21 GND.n20 76
R82 GND.n24 GND.n23 76
R83 GND.n29 GND.n28 76
R84 GND.n32 GND.n31 76
R85 GND.n35 GND.n34 76
R86 GND.n42 GND.n41 76
R87 GND.n45 GND.n44 76
R88 GND.n48 GND.n47 76
R89 GND.n51 GND.n50 76
R90 GND.n54 GND.n53 76
R91 GND.n57 GND.n56 76
R92 GND.n60 GND.n59 76
R93 GND.n63 GND.n62 76
R94 GND.n66 GND.n65 76
R95 GND.n71 GND.n70 76
R96 GND.n74 GND.n73 76
R97 GND.n77 GND.n76 76
R98 GND.n84 GND.n83 76
R99 GND.n87 GND.n86 76
R100 GND.n90 GND.n89 76
R101 GND.n93 GND.n92 76
R102 GND.n96 GND.n95 76
R103 GND.n99 GND.n98 76
R104 GND.n102 GND.n101 76
R105 GND.n105 GND.n104 76
R106 GND.n108 GND.n107 76
R107 GND.n113 GND.n112 76
R108 GND.n116 GND.n115 76
R109 GND.n119 GND.n118 76
R110 GND.n245 GND.n244 76
R111 GND.n238 GND.n237 76
R112 GND.n235 GND.n234 76
R113 GND.n232 GND.n231 76
R114 GND.n229 GND.n228 76
R115 GND.n226 GND.n225 76
R116 GND.n223 GND.n222 76
R117 GND.n220 GND.n219 76
R118 GND.n217 GND.n216 76
R119 GND.n214 GND.n213 76
R120 GND.n209 GND.n208 76
R121 GND.n206 GND.n205 76
R122 GND.n199 GND.n198 76
R123 GND.n196 GND.n195 76
R124 GND.n193 GND.n192 76
R125 GND.n190 GND.n189 76
R126 GND.n187 GND.n186 76
R127 GND.n184 GND.n183 76
R128 GND.n181 GND.n180 76
R129 GND.n178 GND.n177 76
R130 GND.n175 GND.n174 76
R131 GND.n172 GND.n171 76
R132 GND.n167 GND.n166 76
R133 GND.n164 GND.n163 76
R134 GND.n157 GND.n156 76
R135 GND.n154 GND.n153 76
R136 GND.n151 GND.n150 76
R137 GND.n148 GND.n147 76
R138 GND.n145 GND.n144 76
R139 GND.n142 GND.n141 76
R140 GND.n139 GND.n138 76
R141 GND.n136 GND.n135 76
R142 GND.n133 GND.n132 76
R143 GND.n130 GND.n129 76
R144 GND.n125 GND.n124 76
R145 GND.n8 GND.n7 34.942
R146 GND.n6 GND.n5 14.167
R147 GND.n5 GND.n4 14.167
R148 GND.n41 GND.n39 14.167
R149 GND.n83 GND.n81 14.167
R150 GND.n244 GND.n242 14.167
R151 GND.n205 GND.n204 14.167
R152 GND.n163 GND.n162 14.167
R153 GND.n124 GND.n123 13.653
R154 GND.n129 GND.n126 13.653
R155 GND.n132 GND.n131 13.653
R156 GND.n135 GND.n134 13.653
R157 GND.n138 GND.n137 13.653
R158 GND.n141 GND.n140 13.653
R159 GND.n144 GND.n143 13.653
R160 GND.n147 GND.n146 13.653
R161 GND.n150 GND.n149 13.653
R162 GND.n153 GND.n152 13.653
R163 GND.n156 GND.n155 13.653
R164 GND.n163 GND.n158 13.653
R165 GND.n166 GND.n165 13.653
R166 GND.n171 GND.n168 13.653
R167 GND.n174 GND.n173 13.653
R168 GND.n177 GND.n176 13.653
R169 GND.n180 GND.n179 13.653
R170 GND.n183 GND.n182 13.653
R171 GND.n186 GND.n185 13.653
R172 GND.n189 GND.n188 13.653
R173 GND.n192 GND.n191 13.653
R174 GND.n195 GND.n194 13.653
R175 GND.n198 GND.n197 13.653
R176 GND.n205 GND.n200 13.653
R177 GND.n208 GND.n207 13.653
R178 GND.n213 GND.n210 13.653
R179 GND.n216 GND.n215 13.653
R180 GND.n219 GND.n218 13.653
R181 GND.n222 GND.n221 13.653
R182 GND.n225 GND.n224 13.653
R183 GND.n228 GND.n227 13.653
R184 GND.n231 GND.n230 13.653
R185 GND.n234 GND.n233 13.653
R186 GND.n237 GND.n236 13.653
R187 GND.n244 GND.n243 13.653
R188 GND.n118 GND.n117 13.653
R189 GND.n115 GND.n114 13.653
R190 GND.n112 GND.n109 13.653
R191 GND.n107 GND.n106 13.653
R192 GND.n104 GND.n103 13.653
R193 GND.n101 GND.n100 13.653
R194 GND.n98 GND.n97 13.653
R195 GND.n95 GND.n94 13.653
R196 GND.n92 GND.n91 13.653
R197 GND.n89 GND.n88 13.653
R198 GND.n86 GND.n85 13.653
R199 GND.n83 GND.n82 13.653
R200 GND.n76 GND.n75 13.653
R201 GND.n73 GND.n72 13.653
R202 GND.n70 GND.n67 13.653
R203 GND.n65 GND.n64 13.653
R204 GND.n62 GND.n61 13.653
R205 GND.n59 GND.n58 13.653
R206 GND.n56 GND.n55 13.653
R207 GND.n53 GND.n52 13.653
R208 GND.n50 GND.n49 13.653
R209 GND.n47 GND.n46 13.653
R210 GND.n44 GND.n43 13.653
R211 GND.n41 GND.n40 13.653
R212 GND.n34 GND.n33 13.653
R213 GND.n31 GND.n30 13.653
R214 GND.n28 GND.n25 13.653
R215 GND.n23 GND.n22 13.653
R216 GND.n20 GND.n19 13.653
R217 GND.n17 GND.n16 13.653
R218 GND.n14 GND.n13 13.653
R219 GND.n11 GND.n10 13.653
R220 GND.n4 GND.n3 13.653
R221 GND.n5 GND.n2 13.653
R222 GND.n6 GND.n1 13.653
R223 GND.n39 GND.n38 7.312
R224 GND.n162 GND.n161 7.312
R225 GND.n204 GND.n203 7.312
R226 GND.n242 GND.n241 7.312
R227 GND.n81 GND.n80 7.312
R228 GND.n7 GND.n0 7.083
R229 GND.n7 GND.n6 6.474
R230 GND.n121 GND.n120 0.596
R231 GND.n42 GND.n35 0.29
R232 GND.n84 GND.n77 0.29
R233 GND.n206 GND.n199 0.29
R234 GND.n164 GND.n157 0.29
R235 GND.n122 GND 0.207
R236 GND.n18 GND.n15 0.197
R237 GND.n60 GND.n57 0.197
R238 GND.n102 GND.n99 0.197
R239 GND.n226 GND.n223 0.197
R240 GND.n184 GND.n181 0.197
R241 GND.n142 GND.n139 0.197
R242 GND.n28 GND.n27 0.196
R243 GND.n70 GND.n69 0.196
R244 GND.n112 GND.n111 0.196
R245 GND.n213 GND.n212 0.196
R246 GND.n171 GND.n170 0.196
R247 GND.n129 GND.n128 0.196
R248 GND.n9 GND.n8 0.145
R249 GND.n12 GND.n9 0.145
R250 GND.n15 GND.n12 0.145
R251 GND.n21 GND.n18 0.145
R252 GND.n24 GND.n21 0.145
R253 GND.n29 GND.n24 0.145
R254 GND.n32 GND.n29 0.145
R255 GND.n35 GND.n32 0.145
R256 GND.n45 GND.n42 0.145
R257 GND.n48 GND.n45 0.145
R258 GND.n51 GND.n48 0.145
R259 GND.n54 GND.n51 0.145
R260 GND.n57 GND.n54 0.145
R261 GND.n63 GND.n60 0.145
R262 GND.n66 GND.n63 0.145
R263 GND.n71 GND.n66 0.145
R264 GND.n74 GND.n71 0.145
R265 GND.n77 GND.n74 0.145
R266 GND.n87 GND.n84 0.145
R267 GND.n90 GND.n87 0.145
R268 GND.n93 GND.n90 0.145
R269 GND.n96 GND.n93 0.145
R270 GND.n99 GND.n96 0.145
R271 GND.n105 GND.n102 0.145
R272 GND.n108 GND.n105 0.145
R273 GND.n113 GND.n108 0.145
R274 GND.n116 GND.n113 0.145
R275 GND.n119 GND.n116 0.145
R276 GND GND.n119 0.145
R277 GND GND.n245 0.145
R278 GND.n245 GND.n238 0.145
R279 GND.n238 GND.n235 0.145
R280 GND.n235 GND.n232 0.145
R281 GND.n232 GND.n229 0.145
R282 GND.n229 GND.n226 0.145
R283 GND.n223 GND.n220 0.145
R284 GND.n220 GND.n217 0.145
R285 GND.n217 GND.n214 0.145
R286 GND.n214 GND.n209 0.145
R287 GND.n209 GND.n206 0.145
R288 GND.n199 GND.n196 0.145
R289 GND.n196 GND.n193 0.145
R290 GND.n193 GND.n190 0.145
R291 GND.n190 GND.n187 0.145
R292 GND.n187 GND.n184 0.145
R293 GND.n181 GND.n178 0.145
R294 GND.n178 GND.n175 0.145
R295 GND.n175 GND.n172 0.145
R296 GND.n172 GND.n167 0.145
R297 GND.n167 GND.n164 0.145
R298 GND.n157 GND.n154 0.145
R299 GND.n154 GND.n151 0.145
R300 GND.n151 GND.n148 0.145
R301 GND.n148 GND.n145 0.145
R302 GND.n145 GND.n142 0.145
R303 GND.n139 GND.n136 0.145
R304 GND.n136 GND.n133 0.145
R305 GND.n133 GND.n130 0.145
R306 GND.n130 GND.n125 0.145
R307 GND.n125 GND.n122 0.145
R308 a_2201_1050.n5 a_2201_1050.t7 512.525
R309 a_2201_1050.n5 a_2201_1050.t8 371.139
R310 a_2201_1050.n6 a_2201_1050.t9 234.562
R311 a_2201_1050.n7 a_2201_1050.n4 223.905
R312 a_2201_1050.n6 a_2201_1050.n5 215.819
R313 a_2201_1050.n9 a_2201_1050.n7 166.52
R314 a_2201_1050.n7 a_2201_1050.n6 153.315
R315 a_2201_1050.n3 a_2201_1050.n2 79.232
R316 a_2201_1050.n4 a_2201_1050.n3 63.152
R317 a_2201_1050.n4 a_2201_1050.n0 16.08
R318 a_2201_1050.n3 a_2201_1050.n1 16.08
R319 a_2201_1050.n9 a_2201_1050.n8 15.218
R320 a_2201_1050.n0 a_2201_1050.t5 14.282
R321 a_2201_1050.n0 a_2201_1050.t6 14.282
R322 a_2201_1050.n1 a_2201_1050.t3 14.282
R323 a_2201_1050.n1 a_2201_1050.t0 14.282
R324 a_2201_1050.n2 a_2201_1050.t1 14.282
R325 a_2201_1050.n2 a_2201_1050.t4 14.282
R326 a_2201_1050.n10 a_2201_1050.n9 12.014
R327 a_1561_989.n7 a_1561_989.t14 454.685
R328 a_1561_989.n9 a_1561_989.t7 454.685
R329 a_1561_989.n5 a_1561_989.t15 454.685
R330 a_1561_989.n7 a_1561_989.t8 428.979
R331 a_1561_989.n9 a_1561_989.t11 428.979
R332 a_1561_989.n5 a_1561_989.t13 428.979
R333 a_1561_989.n8 a_1561_989.t9 264.512
R334 a_1561_989.n6 a_1561_989.t12 264.512
R335 a_1561_989.n10 a_1561_989.t10 264.173
R336 a_1561_989.n15 a_1561_989.n13 246.179
R337 a_1561_989.n13 a_1561_989.n4 144.246
R338 a_1561_989.n12 a_1561_989.n6 82.484
R339 a_1561_989.n11 a_1561_989.n10 79.495
R340 a_1561_989.n3 a_1561_989.n2 79.232
R341 a_1561_989.n11 a_1561_989.n8 76
R342 a_1561_989.n13 a_1561_989.n12 76
R343 a_1561_989.n8 a_1561_989.n7 71.894
R344 a_1561_989.n6 a_1561_989.n5 71.894
R345 a_1561_989.n10 a_1561_989.n9 71.555
R346 a_1561_989.n4 a_1561_989.n3 63.152
R347 a_1561_989.n4 a_1561_989.n0 16.08
R348 a_1561_989.n3 a_1561_989.n1 16.08
R349 a_1561_989.n15 a_1561_989.n14 15.218
R350 a_1561_989.n0 a_1561_989.t0 14.282
R351 a_1561_989.n0 a_1561_989.t4 14.282
R352 a_1561_989.n1 a_1561_989.t3 14.282
R353 a_1561_989.n1 a_1561_989.t2 14.282
R354 a_1561_989.n2 a_1561_989.t6 14.282
R355 a_1561_989.n2 a_1561_989.t5 14.282
R356 a_1561_989.n16 a_1561_989.n15 12.014
R357 a_1561_989.n12 a_1561_989.n11 4.035
R358 VDD.n344 VDD.n342 144.705
R359 VDD.n502 VDD.n500 144.705
R360 VDD.n425 VDD.n423 144.705
R361 VDD.n184 VDD.n182 144.705
R362 VDD.n103 VDD.n101 144.705
R363 VDD.n43 VDD.n42 76
R364 VDD.n48 VDD.n47 76
R365 VDD.n53 VDD.n52 76
R366 VDD.n60 VDD.n59 76
R367 VDD.n65 VDD.n64 76
R368 VDD.n70 VDD.n69 76
R369 VDD.n74 VDD.n73 76
R370 VDD.n78 VDD.n77 76
R371 VDD.n105 VDD.n104 76
R372 VDD.n109 VDD.n108 76
R373 VDD.n113 VDD.n112 76
R374 VDD.n118 VDD.n117 76
R375 VDD.n125 VDD.n124 76
R376 VDD.n130 VDD.n129 76
R377 VDD.n135 VDD.n134 76
R378 VDD.n142 VDD.n141 76
R379 VDD.n147 VDD.n146 76
R380 VDD.n152 VDD.n151 76
R381 VDD.n156 VDD.n155 76
R382 VDD.n160 VDD.n159 76
R383 VDD.n186 VDD.n185 76
R384 VDD.n190 VDD.n189 76
R385 VDD.n194 VDD.n193 76
R386 VDD.n199 VDD.n198 76
R387 VDD.n206 VDD.n205 76
R388 VDD.n211 VDD.n210 76
R389 VDD.n216 VDD.n215 76
R390 VDD.n223 VDD.n222 76
R391 VDD.n228 VDD.n227 76
R392 VDD.n233 VDD.n232 76
R393 VDD.n237 VDD.n236 76
R394 VDD.n241 VDD.n240 76
R395 VDD.n504 VDD.n503 76
R396 VDD.n478 VDD.n477 76
R397 VDD.n474 VDD.n473 76
R398 VDD.n470 VDD.n469 76
R399 VDD.n465 VDD.n464 76
R400 VDD.n458 VDD.n457 76
R401 VDD.n453 VDD.n452 76
R402 VDD.n448 VDD.n447 76
R403 VDD.n441 VDD.n440 76
R404 VDD.n436 VDD.n435 76
R405 VDD.n431 VDD.n430 76
R406 VDD.n427 VDD.n426 76
R407 VDD.n401 VDD.n400 76
R408 VDD.n397 VDD.n396 76
R409 VDD.n393 VDD.n392 76
R410 VDD.n389 VDD.n388 76
R411 VDD.n384 VDD.n383 76
R412 VDD.n377 VDD.n376 76
R413 VDD.n372 VDD.n371 76
R414 VDD.n367 VDD.n366 76
R415 VDD.n360 VDD.n359 76
R416 VDD.n355 VDD.n354 76
R417 VDD.n350 VDD.n349 76
R418 VDD.n346 VDD.n345 76
R419 VDD.n319 VDD.n318 76
R420 VDD.n315 VDD.n314 76
R421 VDD.n311 VDD.n310 76
R422 VDD.n307 VDD.n306 76
R423 VDD.n302 VDD.n301 76
R424 VDD.n295 VDD.n294 76
R425 VDD.n290 VDD.n289 76
R426 VDD.n285 VDD.n284 76
R427 VDD.n278 VDD.n277 76
R428 VDD.n273 VDD.n272 76
R429 VDD.n268 VDD.n267 76
R430 VDD.n264 VDD.n263 76
R431 VDD.n27 VDD.n26 64.064
R432 VDD.n115 VDD.n114 64.064
R433 VDD.n196 VDD.n195 64.064
R434 VDD.n467 VDD.n466 64.064
R435 VDD.n386 VDD.n385 64.064
R436 VDD.n304 VDD.n303 64.064
R437 VDD.n62 VDD.n61 59.488
R438 VDD.n144 VDD.n143 59.488
R439 VDD.n225 VDD.n224 59.488
R440 VDD.n438 VDD.n437 59.488
R441 VDD.n357 VDD.n356 59.488
R442 VDD.n275 VDD.n274 59.488
R443 VDD.n269 VDD.t20 55.106
R444 VDD.n351 VDD.t34 55.106
R445 VDD.n432 VDD.t19 55.106
R446 VDD.n229 VDD.t31 55.106
R447 VDD.n148 VDD.t7 55.106
R448 VDD.n66 VDD.t22 55.106
R449 VDD.n310 VDD.t0 55.106
R450 VDD.n392 VDD.t26 55.106
R451 VDD.n473 VDD.t29 55.106
R452 VDD.n193 VDD.t2 55.106
R453 VDD.n112 VDD.t4 55.106
R454 VDD.n30 VDD.t30 55.106
R455 VDD.n280 VDD.n279 40.824
R456 VDD.n300 VDD.n299 40.824
R457 VDD.n362 VDD.n361 40.824
R458 VDD.n382 VDD.n381 40.824
R459 VDD.n443 VDD.n442 40.824
R460 VDD.n463 VDD.n462 40.824
R461 VDD.n218 VDD.n217 40.824
R462 VDD.n204 VDD.n203 40.824
R463 VDD.n137 VDD.n136 40.824
R464 VDD.n123 VDD.n122 40.824
R465 VDD.n55 VDD.n54 40.824
R466 VDD.n41 VDD.n40 40.824
R467 VDD.n406 VDD.n405 36.774
R468 VDD.n483 VDD.n482 36.774
R469 VDD.n165 VDD.n164 36.774
R470 VDD.n83 VDD.n82 36.774
R471 VDD.n335 VDD.n334 36.774
R472 VDD.n35 VDD.n34 34.942
R473 VDD.n38 VDD.n37 27.456
R474 VDD.n120 VDD.n119 27.456
R475 VDD.n201 VDD.n200 27.456
R476 VDD.n460 VDD.n459 27.456
R477 VDD.n379 VDD.n378 27.456
R478 VDD.n297 VDD.n296 27.456
R479 VDD.n57 VDD.n56 22.88
R480 VDD.n139 VDD.n138 22.88
R481 VDD.n220 VDD.n219 22.88
R482 VDD.n445 VDD.n444 22.88
R483 VDD.n364 VDD.n363 22.88
R484 VDD.n282 VDD.n281 22.88
R485 VDD.n263 VDD.n260 21.841
R486 VDD.n23 VDD.n20 21.841
R487 VDD.n279 VDD.t18 14.282
R488 VDD.n279 VDD.t6 14.282
R489 VDD.n299 VDD.t3 14.282
R490 VDD.n299 VDD.t9 14.282
R491 VDD.n361 VDD.t11 14.282
R492 VDD.n361 VDD.t35 14.282
R493 VDD.n381 VDD.t25 14.282
R494 VDD.n381 VDD.t10 14.282
R495 VDD.n442 VDD.t1 14.282
R496 VDD.n442 VDD.t5 14.282
R497 VDD.n462 VDD.t28 14.282
R498 VDD.n462 VDD.t17 14.282
R499 VDD.n217 VDD.t12 14.282
R500 VDD.n217 VDD.t32 14.282
R501 VDD.n203 VDD.t15 14.282
R502 VDD.n203 VDD.t13 14.282
R503 VDD.n136 VDD.t16 14.282
R504 VDD.n136 VDD.t24 14.282
R505 VDD.n122 VDD.t33 14.282
R506 VDD.n122 VDD.t14 14.282
R507 VDD.n54 VDD.t8 14.282
R508 VDD.n54 VDD.t21 14.282
R509 VDD.n40 VDD.t27 14.282
R510 VDD.n40 VDD.t23 14.282
R511 VDD.n260 VDD.n243 14.167
R512 VDD.n243 VDD.n242 14.167
R513 VDD.n421 VDD.n403 14.167
R514 VDD.n403 VDD.n402 14.167
R515 VDD.n498 VDD.n480 14.167
R516 VDD.n480 VDD.n479 14.167
R517 VDD.n180 VDD.n162 14.167
R518 VDD.n162 VDD.n161 14.167
R519 VDD.n99 VDD.n80 14.167
R520 VDD.n80 VDD.n79 14.167
R521 VDD.n340 VDD.n321 14.167
R522 VDD.n321 VDD.n320 14.167
R523 VDD.n20 VDD.n19 14.167
R524 VDD.n19 VDD.n17 14.167
R525 VDD.n33 VDD.n30 14.167
R526 VDD.n30 VDD.n29 14.167
R527 VDD.n104 VDD.n100 14.167
R528 VDD.n185 VDD.n181 14.167
R529 VDD.n503 VDD.n499 14.167
R530 VDD.n426 VDD.n422 14.167
R531 VDD.n345 VDD.n341 14.167
R532 VDD.n50 VDD.n49 13.728
R533 VDD.n132 VDD.n131 13.728
R534 VDD.n213 VDD.n212 13.728
R535 VDD.n450 VDD.n449 13.728
R536 VDD.n369 VDD.n368 13.728
R537 VDD.n287 VDD.n286 13.728
R538 VDD.n23 VDD.n22 13.653
R539 VDD.n22 VDD.n21 13.653
R540 VDD.n33 VDD.n32 13.653
R541 VDD.n32 VDD.n31 13.653
R542 VDD.n30 VDD.n25 13.653
R543 VDD.n25 VDD.n24 13.653
R544 VDD.n29 VDD.n28 13.653
R545 VDD.n28 VDD.n27 13.653
R546 VDD.n42 VDD.n39 13.653
R547 VDD.n39 VDD.n38 13.653
R548 VDD.n47 VDD.n46 13.653
R549 VDD.n46 VDD.n45 13.653
R550 VDD.n52 VDD.n51 13.653
R551 VDD.n51 VDD.n50 13.653
R552 VDD.n59 VDD.n58 13.653
R553 VDD.n58 VDD.n57 13.653
R554 VDD.n64 VDD.n63 13.653
R555 VDD.n63 VDD.n62 13.653
R556 VDD.n69 VDD.n68 13.653
R557 VDD.n68 VDD.n67 13.653
R558 VDD.n73 VDD.n72 13.653
R559 VDD.n72 VDD.n71 13.653
R560 VDD.n77 VDD.n76 13.653
R561 VDD.n76 VDD.n75 13.653
R562 VDD.n104 VDD.n103 13.653
R563 VDD.n103 VDD.n102 13.653
R564 VDD.n108 VDD.n107 13.653
R565 VDD.n107 VDD.n106 13.653
R566 VDD.n112 VDD.n111 13.653
R567 VDD.n111 VDD.n110 13.653
R568 VDD.n117 VDD.n116 13.653
R569 VDD.n116 VDD.n115 13.653
R570 VDD.n124 VDD.n121 13.653
R571 VDD.n121 VDD.n120 13.653
R572 VDD.n129 VDD.n128 13.653
R573 VDD.n128 VDD.n127 13.653
R574 VDD.n134 VDD.n133 13.653
R575 VDD.n133 VDD.n132 13.653
R576 VDD.n141 VDD.n140 13.653
R577 VDD.n140 VDD.n139 13.653
R578 VDD.n146 VDD.n145 13.653
R579 VDD.n145 VDD.n144 13.653
R580 VDD.n151 VDD.n150 13.653
R581 VDD.n150 VDD.n149 13.653
R582 VDD.n155 VDD.n154 13.653
R583 VDD.n154 VDD.n153 13.653
R584 VDD.n159 VDD.n158 13.653
R585 VDD.n158 VDD.n157 13.653
R586 VDD.n185 VDD.n184 13.653
R587 VDD.n184 VDD.n183 13.653
R588 VDD.n189 VDD.n188 13.653
R589 VDD.n188 VDD.n187 13.653
R590 VDD.n193 VDD.n192 13.653
R591 VDD.n192 VDD.n191 13.653
R592 VDD.n198 VDD.n197 13.653
R593 VDD.n197 VDD.n196 13.653
R594 VDD.n205 VDD.n202 13.653
R595 VDD.n202 VDD.n201 13.653
R596 VDD.n210 VDD.n209 13.653
R597 VDD.n209 VDD.n208 13.653
R598 VDD.n215 VDD.n214 13.653
R599 VDD.n214 VDD.n213 13.653
R600 VDD.n222 VDD.n221 13.653
R601 VDD.n221 VDD.n220 13.653
R602 VDD.n227 VDD.n226 13.653
R603 VDD.n226 VDD.n225 13.653
R604 VDD.n232 VDD.n231 13.653
R605 VDD.n231 VDD.n230 13.653
R606 VDD.n236 VDD.n235 13.653
R607 VDD.n235 VDD.n234 13.653
R608 VDD.n240 VDD.n239 13.653
R609 VDD.n239 VDD.n238 13.653
R610 VDD.n503 VDD.n502 13.653
R611 VDD.n502 VDD.n501 13.653
R612 VDD.n477 VDD.n476 13.653
R613 VDD.n476 VDD.n475 13.653
R614 VDD.n473 VDD.n472 13.653
R615 VDD.n472 VDD.n471 13.653
R616 VDD.n469 VDD.n468 13.653
R617 VDD.n468 VDD.n467 13.653
R618 VDD.n464 VDD.n461 13.653
R619 VDD.n461 VDD.n460 13.653
R620 VDD.n457 VDD.n456 13.653
R621 VDD.n456 VDD.n455 13.653
R622 VDD.n452 VDD.n451 13.653
R623 VDD.n451 VDD.n450 13.653
R624 VDD.n447 VDD.n446 13.653
R625 VDD.n446 VDD.n445 13.653
R626 VDD.n440 VDD.n439 13.653
R627 VDD.n439 VDD.n438 13.653
R628 VDD.n435 VDD.n434 13.653
R629 VDD.n434 VDD.n433 13.653
R630 VDD.n430 VDD.n429 13.653
R631 VDD.n429 VDD.n428 13.653
R632 VDD.n426 VDD.n425 13.653
R633 VDD.n425 VDD.n424 13.653
R634 VDD.n400 VDD.n399 13.653
R635 VDD.n399 VDD.n398 13.653
R636 VDD.n396 VDD.n395 13.653
R637 VDD.n395 VDD.n394 13.653
R638 VDD.n392 VDD.n391 13.653
R639 VDD.n391 VDD.n390 13.653
R640 VDD.n388 VDD.n387 13.653
R641 VDD.n387 VDD.n386 13.653
R642 VDD.n383 VDD.n380 13.653
R643 VDD.n380 VDD.n379 13.653
R644 VDD.n376 VDD.n375 13.653
R645 VDD.n375 VDD.n374 13.653
R646 VDD.n371 VDD.n370 13.653
R647 VDD.n370 VDD.n369 13.653
R648 VDD.n366 VDD.n365 13.653
R649 VDD.n365 VDD.n364 13.653
R650 VDD.n359 VDD.n358 13.653
R651 VDD.n358 VDD.n357 13.653
R652 VDD.n354 VDD.n353 13.653
R653 VDD.n353 VDD.n352 13.653
R654 VDD.n349 VDD.n348 13.653
R655 VDD.n348 VDD.n347 13.653
R656 VDD.n345 VDD.n344 13.653
R657 VDD.n344 VDD.n343 13.653
R658 VDD.n318 VDD.n317 13.653
R659 VDD.n317 VDD.n316 13.653
R660 VDD.n314 VDD.n313 13.653
R661 VDD.n313 VDD.n312 13.653
R662 VDD.n310 VDD.n309 13.653
R663 VDD.n309 VDD.n308 13.653
R664 VDD.n306 VDD.n305 13.653
R665 VDD.n305 VDD.n304 13.653
R666 VDD.n301 VDD.n298 13.653
R667 VDD.n298 VDD.n297 13.653
R668 VDD.n294 VDD.n293 13.653
R669 VDD.n293 VDD.n292 13.653
R670 VDD.n289 VDD.n288 13.653
R671 VDD.n288 VDD.n287 13.653
R672 VDD.n284 VDD.n283 13.653
R673 VDD.n283 VDD.n282 13.653
R674 VDD.n277 VDD.n276 13.653
R675 VDD.n276 VDD.n275 13.653
R676 VDD.n272 VDD.n271 13.653
R677 VDD.n271 VDD.n270 13.653
R678 VDD.n267 VDD.n266 13.653
R679 VDD.n266 VDD.n265 13.653
R680 VDD.n263 VDD.n262 13.653
R681 VDD.n262 VDD.n261 13.653
R682 VDD.n4 VDD.n2 12.915
R683 VDD.n4 VDD.n3 12.66
R684 VDD.n10 VDD.n9 12.343
R685 VDD.n12 VDD.n11 12.343
R686 VDD.n10 VDD.n7 12.343
R687 VDD.n45 VDD.n44 9.152
R688 VDD.n127 VDD.n126 9.152
R689 VDD.n208 VDD.n207 9.152
R690 VDD.n455 VDD.n454 9.152
R691 VDD.n374 VDD.n373 9.152
R692 VDD.n292 VDD.n291 9.152
R693 VDD.n422 VDD.n421 7.674
R694 VDD.n499 VDD.n498 7.674
R695 VDD.n181 VDD.n180 7.674
R696 VDD.n100 VDD.n99 7.674
R697 VDD.n341 VDD.n340 7.674
R698 VDD.n94 VDD.n93 7.5
R699 VDD.n88 VDD.n87 7.5
R700 VDD.n90 VDD.n89 7.5
R701 VDD.n85 VDD.n84 7.5
R702 VDD.n99 VDD.n98 7.5
R703 VDD.n175 VDD.n174 7.5
R704 VDD.n169 VDD.n168 7.5
R705 VDD.n171 VDD.n170 7.5
R706 VDD.n177 VDD.n167 7.5
R707 VDD.n177 VDD.n165 7.5
R708 VDD.n180 VDD.n179 7.5
R709 VDD.n493 VDD.n492 7.5
R710 VDD.n487 VDD.n486 7.5
R711 VDD.n489 VDD.n488 7.5
R712 VDD.n495 VDD.n485 7.5
R713 VDD.n495 VDD.n483 7.5
R714 VDD.n498 VDD.n497 7.5
R715 VDD.n416 VDD.n415 7.5
R716 VDD.n410 VDD.n409 7.5
R717 VDD.n412 VDD.n411 7.5
R718 VDD.n418 VDD.n408 7.5
R719 VDD.n418 VDD.n406 7.5
R720 VDD.n421 VDD.n420 7.5
R721 VDD.n325 VDD.n324 7.5
R722 VDD.n328 VDD.n327 7.5
R723 VDD.n330 VDD.n329 7.5
R724 VDD.n333 VDD.n332 7.5
R725 VDD.n340 VDD.n339 7.5
R726 VDD.n255 VDD.n254 7.5
R727 VDD.n249 VDD.n248 7.5
R728 VDD.n251 VDD.n250 7.5
R729 VDD.n257 VDD.n247 7.5
R730 VDD.n257 VDD.n245 7.5
R731 VDD.n260 VDD.n259 7.5
R732 VDD.n20 VDD.n16 7.5
R733 VDD.n2 VDD.n1 7.5
R734 VDD.n9 VDD.n8 7.5
R735 VDD.n7 VDD.n6 7.5
R736 VDD.n19 VDD.n18 7.5
R737 VDD.n14 VDD.n0 7.5
R738 VDD.n86 VDD.n83 6.772
R739 VDD.n97 VDD.n81 6.772
R740 VDD.n95 VDD.n92 6.772
R741 VDD.n91 VDD.n88 6.772
R742 VDD.n178 VDD.n163 6.772
R743 VDD.n176 VDD.n173 6.772
R744 VDD.n172 VDD.n169 6.772
R745 VDD.n496 VDD.n481 6.772
R746 VDD.n494 VDD.n491 6.772
R747 VDD.n490 VDD.n487 6.772
R748 VDD.n419 VDD.n404 6.772
R749 VDD.n417 VDD.n414 6.772
R750 VDD.n413 VDD.n410 6.772
R751 VDD.n258 VDD.n244 6.772
R752 VDD.n256 VDD.n253 6.772
R753 VDD.n252 VDD.n249 6.772
R754 VDD.n86 VDD.n85 6.772
R755 VDD.n91 VDD.n90 6.772
R756 VDD.n95 VDD.n94 6.772
R757 VDD.n98 VDD.n97 6.772
R758 VDD.n172 VDD.n171 6.772
R759 VDD.n176 VDD.n175 6.772
R760 VDD.n179 VDD.n178 6.772
R761 VDD.n490 VDD.n489 6.772
R762 VDD.n494 VDD.n493 6.772
R763 VDD.n497 VDD.n496 6.772
R764 VDD.n413 VDD.n412 6.772
R765 VDD.n417 VDD.n416 6.772
R766 VDD.n420 VDD.n419 6.772
R767 VDD.n252 VDD.n251 6.772
R768 VDD.n256 VDD.n255 6.772
R769 VDD.n259 VDD.n258 6.772
R770 VDD.n339 VDD.n338 6.772
R771 VDD.n326 VDD.n323 6.772
R772 VDD.n331 VDD.n328 6.772
R773 VDD.n336 VDD.n333 6.772
R774 VDD.n336 VDD.n335 6.772
R775 VDD.n331 VDD.n330 6.772
R776 VDD.n326 VDD.n325 6.772
R777 VDD.n338 VDD.n322 6.772
R778 VDD.n59 VDD.n55 6.69
R779 VDD.n141 VDD.n137 6.69
R780 VDD.n222 VDD.n218 6.69
R781 VDD.n447 VDD.n443 6.69
R782 VDD.n366 VDD.n362 6.69
R783 VDD.n284 VDD.n280 6.69
R784 VDD.n34 VDD.n23 6.487
R785 VDD.n34 VDD.n33 6.475
R786 VDD.n16 VDD.n15 6.458
R787 VDD.n42 VDD.n41 6.296
R788 VDD.n124 VDD.n123 6.296
R789 VDD.n205 VDD.n204 6.296
R790 VDD.n464 VDD.n463 6.296
R791 VDD.n383 VDD.n382 6.296
R792 VDD.n301 VDD.n300 6.296
R793 VDD.n167 VDD.n166 6.202
R794 VDD.n485 VDD.n484 6.202
R795 VDD.n408 VDD.n407 6.202
R796 VDD.n247 VDD.n246 6.202
R797 VDD.n14 VDD.n5 1.329
R798 VDD.n14 VDD.n10 1.329
R799 VDD.n14 VDD.n12 1.329
R800 VDD.n14 VDD.n13 1.329
R801 VDD.n15 VDD.n14 0.696
R802 VDD.n14 VDD.n4 0.696
R803 VDD.n69 VDD.n66 0.393
R804 VDD.n151 VDD.n148 0.393
R805 VDD.n232 VDD.n229 0.393
R806 VDD.n435 VDD.n432 0.393
R807 VDD.n354 VDD.n351 0.393
R808 VDD.n272 VDD.n269 0.393
R809 VDD.n96 VDD.n95 0.365
R810 VDD.n96 VDD.n91 0.365
R811 VDD.n96 VDD.n86 0.365
R812 VDD.n97 VDD.n96 0.365
R813 VDD.n177 VDD.n176 0.365
R814 VDD.n177 VDD.n172 0.365
R815 VDD.n178 VDD.n177 0.365
R816 VDD.n495 VDD.n494 0.365
R817 VDD.n495 VDD.n490 0.365
R818 VDD.n496 VDD.n495 0.365
R819 VDD.n418 VDD.n417 0.365
R820 VDD.n418 VDD.n413 0.365
R821 VDD.n419 VDD.n418 0.365
R822 VDD.n257 VDD.n256 0.365
R823 VDD.n257 VDD.n252 0.365
R824 VDD.n258 VDD.n257 0.365
R825 VDD.n337 VDD.n336 0.365
R826 VDD.n337 VDD.n331 0.365
R827 VDD.n337 VDD.n326 0.365
R828 VDD.n338 VDD.n337 0.365
R829 VDD.n105 VDD.n78 0.29
R830 VDD.n186 VDD.n160 0.29
R831 VDD.n427 VDD.n401 0.29
R832 VDD.n346 VDD.n319 0.29
R833 VDD.n264 VDD 0.207
R834 VDD.n53 VDD.n48 0.197
R835 VDD.n135 VDD.n130 0.197
R836 VDD.n216 VDD.n211 0.197
R837 VDD.n458 VDD.n453 0.197
R838 VDD.n377 VDD.n372 0.197
R839 VDD.n295 VDD.n290 0.197
R840 VDD.n36 VDD.n35 0.145
R841 VDD.n43 VDD.n36 0.145
R842 VDD.n48 VDD.n43 0.145
R843 VDD.n60 VDD.n53 0.145
R844 VDD.n65 VDD.n60 0.145
R845 VDD.n70 VDD.n65 0.145
R846 VDD.n74 VDD.n70 0.145
R847 VDD.n78 VDD.n74 0.145
R848 VDD.n109 VDD.n105 0.145
R849 VDD.n113 VDD.n109 0.145
R850 VDD.n118 VDD.n113 0.145
R851 VDD.n125 VDD.n118 0.145
R852 VDD.n130 VDD.n125 0.145
R853 VDD.n142 VDD.n135 0.145
R854 VDD.n147 VDD.n142 0.145
R855 VDD.n152 VDD.n147 0.145
R856 VDD.n156 VDD.n152 0.145
R857 VDD.n160 VDD.n156 0.145
R858 VDD.n190 VDD.n186 0.145
R859 VDD.n194 VDD.n190 0.145
R860 VDD.n199 VDD.n194 0.145
R861 VDD.n206 VDD.n199 0.145
R862 VDD.n211 VDD.n206 0.145
R863 VDD.n223 VDD.n216 0.145
R864 VDD.n228 VDD.n223 0.145
R865 VDD.n233 VDD.n228 0.145
R866 VDD.n237 VDD.n233 0.145
R867 VDD.n241 VDD.n237 0.145
R868 VDD VDD.n241 0.145
R869 VDD VDD.n504 0.145
R870 VDD.n504 VDD.n478 0.145
R871 VDD.n478 VDD.n474 0.145
R872 VDD.n474 VDD.n470 0.145
R873 VDD.n470 VDD.n465 0.145
R874 VDD.n465 VDD.n458 0.145
R875 VDD.n453 VDD.n448 0.145
R876 VDD.n448 VDD.n441 0.145
R877 VDD.n441 VDD.n436 0.145
R878 VDD.n436 VDD.n431 0.145
R879 VDD.n431 VDD.n427 0.145
R880 VDD.n401 VDD.n397 0.145
R881 VDD.n397 VDD.n393 0.145
R882 VDD.n393 VDD.n389 0.145
R883 VDD.n389 VDD.n384 0.145
R884 VDD.n384 VDD.n377 0.145
R885 VDD.n372 VDD.n367 0.145
R886 VDD.n367 VDD.n360 0.145
R887 VDD.n360 VDD.n355 0.145
R888 VDD.n355 VDD.n350 0.145
R889 VDD.n350 VDD.n346 0.145
R890 VDD.n319 VDD.n315 0.145
R891 VDD.n315 VDD.n311 0.145
R892 VDD.n311 VDD.n307 0.145
R893 VDD.n307 VDD.n302 0.145
R894 VDD.n302 VDD.n295 0.145
R895 VDD.n290 VDD.n285 0.145
R896 VDD.n285 VDD.n278 0.145
R897 VDD.n278 VDD.n273 0.145
R898 VDD.n273 VDD.n268 0.145
R899 VDD.n268 VDD.n264 0.145
R900 SN.n2 SN.t1 479.223
R901 SN.n0 SN.t2 479.223
R902 SN.n2 SN.t3 375.52
R903 SN.n0 SN.t0 375.52
R904 SN.n1 SN.n0 175.429
R905 SN.n3 SN.n2 175.07
R906 SN.n3 SN.t4 162.407
R907 SN.n1 SN.t5 162.048
R908 SN.n4 SN.n1 86.561
R909 SN.n4 SN.n3 76
R910 SN.n4 SN 0.046
R911 Q.n10 Q.t7 454.685
R912 Q.n10 Q.t9 428.979
R913 Q.n11 Q.t8 237.959
R914 Q.n9 Q.n8 213.104
R915 Q.n9 Q.n4 170.799
R916 Q.n11 Q.n10 98.447
R917 Q Q.n11 79.989
R918 Q.n3 Q.n2 79.232
R919 Q.n12 Q.n9 76
R920 Q.n4 Q.n3 63.152
R921 Q.n8 Q.n7 30
R922 Q.n6 Q.n5 24.383
R923 Q.n8 Q.n6 23.684
R924 Q.n4 Q.n0 16.08
R925 Q.n3 Q.n1 16.08
R926 Q.n0 Q.t6 14.282
R927 Q.n0 Q.t5 14.282
R928 Q.n1 Q.t0 14.282
R929 Q.n1 Q.t1 14.282
R930 Q.n2 Q.t3 14.282
R931 Q.n2 Q.t2 14.282
R932 Q.n12 Q 0.046
R933 D.n0 D.t0 512.525
R934 D.n0 D.t2 371.139
R935 D.n1 D.t1 234.562
R936 D.n1 D.n0 215.819
R937 D.n2 D.n1 76
R938 D.n2 D 0.046
R939 a_277_1050.n4 a_277_1050.t8 512.525
R940 a_277_1050.n2 a_277_1050.t7 512.525
R941 a_277_1050.n4 a_277_1050.t11 371.139
R942 a_277_1050.n2 a_277_1050.t12 371.139
R943 a_277_1050.n5 a_277_1050.t10 234.921
R944 a_277_1050.n3 a_277_1050.t9 234.921
R945 a_277_1050.n9 a_277_1050.n8 223.546
R946 a_277_1050.n5 a_277_1050.n4 215.46
R947 a_277_1050.n3 a_277_1050.n2 215.46
R948 a_277_1050.n8 a_277_1050.n7 182.096
R949 a_277_1050.n6 a_277_1050.n3 79.491
R950 a_277_1050.n11 a_277_1050.n10 79.231
R951 a_277_1050.n8 a_277_1050.n6 77.315
R952 a_277_1050.n6 a_277_1050.n5 76
R953 a_277_1050.n10 a_277_1050.n9 63.152
R954 a_277_1050.n9 a_277_1050.n1 16.08
R955 a_277_1050.n10 a_277_1050.n0 16.08
R956 a_277_1050.n1 a_277_1050.t0 14.282
R957 a_277_1050.n1 a_277_1050.t2 14.282
R958 a_277_1050.n0 a_277_1050.t3 14.282
R959 a_277_1050.n0 a_277_1050.t4 14.282
R960 a_277_1050.t6 a_277_1050.n11 14.282
R961 a_277_1050.n11 a_277_1050.t5 14.282
R962 a_599_989.n1 a_599_989.t12 512.525
R963 a_599_989.n3 a_599_989.t10 454.685
R964 a_599_989.n3 a_599_989.t9 428.979
R965 a_599_989.n1 a_599_989.t8 371.139
R966 a_599_989.n2 a_599_989.t11 287.668
R967 a_599_989.n4 a_599_989.t7 237.959
R968 a_599_989.n10 a_599_989.n9 213.104
R969 a_599_989.n11 a_599_989.n10 170.799
R970 a_599_989.n2 a_599_989.n1 162.713
R971 a_599_989.n4 a_599_989.n3 98.447
R972 a_599_989.n5 a_599_989.n2 84.388
R973 a_599_989.n5 a_599_989.n4 80.035
R974 a_599_989.n13 a_599_989.n12 79.232
R975 a_599_989.n10 a_599_989.n5 76
R976 a_599_989.n13 a_599_989.n11 63.152
R977 a_599_989.n9 a_599_989.n8 30
R978 a_599_989.n7 a_599_989.n6 24.383
R979 a_599_989.n9 a_599_989.n7 23.684
R980 a_599_989.n11 a_599_989.n0 16.08
R981 a_599_989.n14 a_599_989.n13 16.078
R982 a_599_989.n0 a_599_989.t5 14.282
R983 a_599_989.n0 a_599_989.t6 14.282
R984 a_599_989.n12 a_599_989.t3 14.282
R985 a_599_989.n12 a_599_989.t2 14.282
R986 a_599_989.n14 a_599_989.t0 14.282
R987 a_599_989.t1 a_599_989.n14 14.282
R988 a_372_210.n10 a_372_210.n8 82.852
R989 a_372_210.n11 a_372_210.n0 49.6
R990 a_372_210.n7 a_372_210.n6 32.833
R991 a_372_210.n8 a_372_210.t1 32.416
R992 a_372_210.n10 a_372_210.n9 27.2
R993 a_372_210.n3 a_372_210.n2 23.284
R994 a_372_210.n11 a_372_210.n10 22.4
R995 a_372_210.n7 a_372_210.n4 19.017
R996 a_372_210.n6 a_372_210.n5 13.494
R997 a_372_210.t1 a_372_210.n1 7.04
R998 a_372_210.t1 a_372_210.n3 5.727
R999 a_372_210.n8 a_372_210.n7 1.435
R1000 RN.n5 RN.t0 479.223
R1001 RN.n0 RN.t7 479.223
R1002 RN.n2 RN.t6 454.685
R1003 RN.n2 RN.t1 428.979
R1004 RN.n5 RN.t5 375.52
R1005 RN.n0 RN.t2 375.52
R1006 RN.n6 RN.t3 294.813
R1007 RN.n1 RN.t8 294.813
R1008 RN.n3 RN.t4 291.065
R1009 RN.n4 RN.n1 78.675
R1010 RN.n4 RN.n3 76
R1011 RN.n7 RN.n6 76
R1012 RN.n3 RN.n2 45.341
R1013 RN.n6 RN.n5 42.664
R1014 RN.n1 RN.n0 42.664
R1015 RN.n7 RN.n4 11.381
R1016 RN.n7 RN 0.046
R1017 a_91_103.n5 a_91_103.n4 19.724
R1018 a_91_103.t0 a_91_103.n3 11.595
R1019 a_91_103.t0 a_91_103.n5 9.207
R1020 a_91_103.n2 a_91_103.n1 2.455
R1021 a_91_103.n2 a_91_103.n0 1.32
R1022 a_91_103.t0 a_91_103.n2 0.246
R1023 a_2296_210.n10 a_2296_210.n8 82.852
R1024 a_2296_210.n7 a_2296_210.n6 32.833
R1025 a_2296_210.n8 a_2296_210.t1 32.416
R1026 a_2296_210.n10 a_2296_210.n9 27.2
R1027 a_2296_210.n11 a_2296_210.n0 23.498
R1028 a_2296_210.n3 a_2296_210.n2 23.284
R1029 a_2296_210.n11 a_2296_210.n10 22.4
R1030 a_2296_210.n7 a_2296_210.n4 19.017
R1031 a_2296_210.n6 a_2296_210.n5 13.494
R1032 a_2296_210.t1 a_2296_210.n1 7.04
R1033 a_2296_210.t1 a_2296_210.n3 5.727
R1034 a_2296_210.n8 a_2296_210.n7 1.435
R1035 a_4220_210.n9 a_4220_210.n7 82.852
R1036 a_4220_210.n3 a_4220_210.n1 44.628
R1037 a_4220_210.t0 a_4220_210.n9 32.417
R1038 a_4220_210.n7 a_4220_210.n6 27.2
R1039 a_4220_210.n5 a_4220_210.n4 23.498
R1040 a_4220_210.n3 a_4220_210.n2 23.284
R1041 a_4220_210.n7 a_4220_210.n5 22.4
R1042 a_4220_210.t0 a_4220_210.n11 20.241
R1043 a_4220_210.n11 a_4220_210.n10 13.494
R1044 a_4220_210.t0 a_4220_210.n0 8.137
R1045 a_4220_210.t0 a_4220_210.n3 5.727
R1046 a_4220_210.n9 a_4220_210.n8 1.435
R1047 a_1334_210.n10 a_1334_210.n8 82.852
R1048 a_1334_210.n7 a_1334_210.n6 32.833
R1049 a_1334_210.n8 a_1334_210.t1 32.416
R1050 a_1334_210.n10 a_1334_210.n9 27.2
R1051 a_1334_210.n11 a_1334_210.n0 23.498
R1052 a_1334_210.n3 a_1334_210.n2 23.284
R1053 a_1334_210.n11 a_1334_210.n10 22.4
R1054 a_1334_210.n7 a_1334_210.n4 19.017
R1055 a_1334_210.n6 a_1334_210.n5 13.494
R1056 a_1334_210.t1 a_1334_210.n1 7.04
R1057 a_1334_210.t1 a_1334_210.n3 5.727
R1058 a_1334_210.n8 a_1334_210.n7 1.435
R1059 a_2015_103.n1 a_2015_103.n0 25.576
R1060 a_2015_103.n3 a_2015_103.n2 9.111
R1061 a_2015_103.n7 a_2015_103.n6 2.455
R1062 a_2015_103.n5 a_2015_103.n3 1.964
R1063 a_2015_103.n5 a_2015_103.n4 1.964
R1064 a_2015_103.t0 a_2015_103.n1 1.871
R1065 a_2015_103.n7 a_2015_103.n5 0.636
R1066 a_2015_103.t0 a_2015_103.n7 0.246
R1067 a_5182_210.n10 a_5182_210.n8 82.852
R1068 a_5182_210.n11 a_5182_210.n0 49.6
R1069 a_5182_210.n7 a_5182_210.n6 32.833
R1070 a_5182_210.n8 a_5182_210.t1 32.416
R1071 a_5182_210.n10 a_5182_210.n9 27.2
R1072 a_5182_210.n3 a_5182_210.n2 23.284
R1073 a_5182_210.n11 a_5182_210.n10 22.4
R1074 a_5182_210.n7 a_5182_210.n4 19.017
R1075 a_5182_210.n6 a_5182_210.n5 13.494
R1076 a_5182_210.t1 a_5182_210.n1 7.04
R1077 a_5182_210.t1 a_5182_210.n3 5.727
R1078 a_5182_210.n8 a_5182_210.n7 1.435
R1079 a_1053_103.n1 a_1053_103.n0 25.576
R1080 a_1053_103.n3 a_1053_103.n2 9.111
R1081 a_1053_103.n7 a_1053_103.n6 2.455
R1082 a_1053_103.n5 a_1053_103.n3 1.964
R1083 a_1053_103.n5 a_1053_103.n4 1.964
R1084 a_1053_103.t0 a_1053_103.n1 1.871
R1085 a_1053_103.n7 a_1053_103.n5 0.636
R1086 a_1053_103.t0 a_1053_103.n7 0.246
R1087 a_3939_103.n5 a_3939_103.n4 19.724
R1088 a_3939_103.t0 a_3939_103.n3 11.595
R1089 a_3939_103.t0 a_3939_103.n5 9.207
R1090 a_3939_103.n2 a_3939_103.n1 2.455
R1091 a_3939_103.n2 a_3939_103.n0 1.32
R1092 a_3939_103.t0 a_3939_103.n2 0.246
C11 SN GND 2.29fF
C12 RN GND 1.35fF
C13 VDD GND 21.17fF
C14 a_3939_103.n0 GND 0.10fF
C15 a_3939_103.n1 GND 0.04fF
C16 a_3939_103.n2 GND 0.03fF
C17 a_3939_103.n3 GND 0.07fF
C18 a_3939_103.n4 GND 0.08fF
C19 a_3939_103.n5 GND 0.06fF
C20 a_1053_103.n0 GND 0.09fF
C21 a_1053_103.n1 GND 0.10fF
C22 a_1053_103.n2 GND 0.05fF
C23 a_1053_103.n3 GND 0.03fF
C24 a_1053_103.n4 GND 0.04fF
C25 a_1053_103.n5 GND 0.03fF
C26 a_1053_103.n6 GND 0.04fF
C27 a_5182_210.n0 GND 0.02fF
C28 a_5182_210.n1 GND 0.09fF
C29 a_5182_210.n2 GND 0.13fF
C30 a_5182_210.n3 GND 0.11fF
C31 a_5182_210.n4 GND 0.09fF
C32 a_5182_210.n5 GND 0.05fF
C33 a_5182_210.n6 GND 0.01fF
C34 a_5182_210.n7 GND 0.03fF
C35 a_5182_210.n8 GND 0.11fF
C36 a_5182_210.n9 GND 0.02fF
C37 a_5182_210.n10 GND 0.05fF
C38 a_5182_210.n11 GND 0.02fF
C39 a_2015_103.n0 GND 0.09fF
C40 a_2015_103.n1 GND 0.10fF
C41 a_2015_103.n2 GND 0.05fF
C42 a_2015_103.n3 GND 0.03fF
C43 a_2015_103.n4 GND 0.04fF
C44 a_2015_103.n5 GND 0.03fF
C45 a_2015_103.n6 GND 0.04fF
C46 a_1334_210.n0 GND 0.02fF
C47 a_1334_210.n1 GND 0.09fF
C48 a_1334_210.n2 GND 0.13fF
C49 a_1334_210.n3 GND 0.11fF
C50 a_1334_210.t1 GND 0.30fF
C51 a_1334_210.n4 GND 0.09fF
C52 a_1334_210.n5 GND 0.06fF
C53 a_1334_210.n6 GND 0.01fF
C54 a_1334_210.n7 GND 0.03fF
C55 a_1334_210.n8 GND 0.11fF
C56 a_1334_210.n9 GND 0.02fF
C57 a_1334_210.n10 GND 0.05fF
C58 a_1334_210.n11 GND 0.03fF
C59 a_4220_210.n0 GND 0.07fF
C60 a_4220_210.n1 GND 0.09fF
C61 a_4220_210.n2 GND 0.13fF
C62 a_4220_210.n3 GND 0.11fF
C63 a_4220_210.n4 GND 0.02fF
C64 a_4220_210.n5 GND 0.03fF
C65 a_4220_210.n6 GND 0.02fF
C66 a_4220_210.n7 GND 0.05fF
C67 a_4220_210.n8 GND 0.03fF
C68 a_4220_210.n9 GND 0.11fF
C69 a_4220_210.n10 GND 0.06fF
C70 a_4220_210.n11 GND 0.01fF
C71 a_4220_210.t0 GND 0.33fF
C72 a_2296_210.n0 GND 0.02fF
C73 a_2296_210.n1 GND 0.09fF
C74 a_2296_210.n2 GND 0.13fF
C75 a_2296_210.n3 GND 0.11fF
C76 a_2296_210.t1 GND 0.30fF
C77 a_2296_210.n4 GND 0.09fF
C78 a_2296_210.n5 GND 0.06fF
C79 a_2296_210.n6 GND 0.01fF
C80 a_2296_210.n7 GND 0.03fF
C81 a_2296_210.n8 GND 0.11fF
C82 a_2296_210.n9 GND 0.02fF
C83 a_2296_210.n10 GND 0.05fF
C84 a_2296_210.n11 GND 0.03fF
C85 a_91_103.n0 GND 0.10fF
C86 a_91_103.n1 GND 0.04fF
C87 a_91_103.n2 GND 0.03fF
C88 a_91_103.n3 GND 0.06fF
C89 a_91_103.n4 GND 0.08fF
C90 a_91_103.n5 GND 0.06fF
C91 RN.n0 GND 0.44fF
C92 RN.t8 GND 0.77fF
C93 RN.n1 GND 0.51fF
C94 RN.n2 GND 0.42fF
C95 RN.t4 GND 0.78fF
C96 RN.n3 GND 0.50fF
C97 RN.n4 GND 2.53fF
C98 RN.n5 GND 0.44fF
C99 RN.t3 GND 0.77fF
C100 RN.n6 GND 0.50fF
C101 RN.n7 GND 1.71fF
C102 a_372_210.n0 GND 0.02fF
C103 a_372_210.n1 GND 0.09fF
C104 a_372_210.n2 GND 0.13fF
C105 a_372_210.n3 GND 0.11fF
C106 a_372_210.t1 GND 0.30fF
C107 a_372_210.n4 GND 0.09fF
C108 a_372_210.n5 GND 0.06fF
C109 a_372_210.n6 GND 0.01fF
C110 a_372_210.n7 GND 0.03fF
C111 a_372_210.n8 GND 0.11fF
C112 a_372_210.n9 GND 0.02fF
C113 a_372_210.n10 GND 0.05fF
C114 a_372_210.n11 GND 0.02fF
C115 a_599_989.n0 GND 0.78fF
C116 a_599_989.n1 GND 0.49fF
C117 a_599_989.n2 GND 0.83fF
C118 a_599_989.n3 GND 0.54fF
C119 a_599_989.t7 GND 0.77fF
C120 a_599_989.n4 GND 0.57fF
C121 a_599_989.n5 GND 3.94fF
C122 a_599_989.n6 GND 0.06fF
C123 a_599_989.n7 GND 0.08fF
C124 a_599_989.n8 GND 0.05fF
C125 a_599_989.n9 GND 0.44fF
C126 a_599_989.n10 GND 0.65fF
C127 a_599_989.n11 GND 0.44fF
C128 a_599_989.n12 GND 0.91fF
C129 a_599_989.n13 GND 0.29fF
C130 a_599_989.n14 GND 0.78fF
C131 a_277_1050.n0 GND 0.49fF
C132 a_277_1050.n1 GND 0.49fF
C133 a_277_1050.n2 GND 0.36fF
C134 a_277_1050.n3 GND 0.44fF
C135 a_277_1050.n4 GND 0.36fF
C136 a_277_1050.n5 GND 0.43fF
C137 a_277_1050.n6 GND 1.03fF
C138 a_277_1050.n7 GND 0.31fF
C139 a_277_1050.n8 GND 0.44fF
C140 a_277_1050.n9 GND 0.33fF
C141 a_277_1050.n10 GND 0.18fF
C142 a_277_1050.n11 GND 0.57fF
C143 Q.n0 GND 0.54fF
C144 Q.n1 GND 0.54fF
C145 Q.n2 GND 0.63fF
C146 Q.n3 GND 0.20fF
C147 Q.n4 GND 0.31fF
C148 Q.n5 GND 0.04fF
C149 Q.n6 GND 0.05fF
C150 Q.n7 GND 0.03fF
C151 Q.n8 GND 0.30fF
C152 Q.n9 GND 0.45fF
C153 Q.n10 GND 0.38fF
C154 Q.t8 GND 0.54fF
C155 Q.n11 GND 0.39fF
C156 Q.n12 GND 0.03fF
C157 SN.n0 GND 0.54fF
C158 SN.t5 GND 0.49fF
C159 SN.n1 GND 0.57fF
C160 SN.n2 GND 0.54fF
C161 SN.t4 GND 0.49fF
C162 SN.n3 GND 0.40fF
C163 SN.n4 GND 2.52fF
C164 VDD.n0 GND 0.19fF
C165 VDD.n1 GND 0.02fF
C166 VDD.n2 GND 0.02fF
C167 VDD.n3 GND 0.04fF
C168 VDD.n4 GND 0.01fF
C169 VDD.n6 GND 0.02fF
C170 VDD.n7 GND 0.02fF
C171 VDD.n8 GND 0.02fF
C172 VDD.n9 GND 0.02fF
C173 VDD.n11 GND 0.02fF
C174 VDD.n14 GND 0.44fF
C175 VDD.n16 GND 0.03fF
C176 VDD.n17 GND 0.02fF
C177 VDD.n18 GND 0.02fF
C178 VDD.n19 GND 0.02fF
C179 VDD.n20 GND 0.03fF
C180 VDD.n21 GND 0.26fF
C181 VDD.n22 GND 0.02fF
C182 VDD.n23 GND 0.03fF
C183 VDD.n24 GND 0.21fF
C184 VDD.n25 GND 0.01fF
C185 VDD.n26 GND 0.13fF
C186 VDD.n27 GND 0.16fF
C187 VDD.n28 GND 0.01fF
C188 VDD.n29 GND 0.02fF
C189 VDD.n30 GND 0.06fF
C190 VDD.n31 GND 0.26fF
C191 VDD.n32 GND 0.01fF
C192 VDD.n33 GND 0.02fF
C193 VDD.n34 GND 0.00fF
C194 VDD.n35 GND 0.09fF
C195 VDD.n36 GND 0.02fF
C196 VDD.n37 GND 0.13fF
C197 VDD.n38 GND 0.15fF
C198 VDD.n39 GND 0.01fF
C199 VDD.n40 GND 0.10fF
C200 VDD.n41 GND 0.02fF
C201 VDD.n42 GND 0.02fF
C202 VDD.n43 GND 0.02fF
C203 VDD.n44 GND 0.17fF
C204 VDD.n45 GND 0.14fF
C205 VDD.n46 GND 0.01fF
C206 VDD.n47 GND 0.02fF
C207 VDD.n48 GND 0.03fF
C208 VDD.n49 GND 0.17fF
C209 VDD.n50 GND 0.14fF
C210 VDD.n51 GND 0.01fF
C211 VDD.n52 GND 0.02fF
C212 VDD.n53 GND 0.03fF
C213 VDD.n54 GND 0.10fF
C214 VDD.n55 GND 0.02fF
C215 VDD.n56 GND 0.13fF
C216 VDD.n57 GND 0.15fF
C217 VDD.n58 GND 0.01fF
C218 VDD.n59 GND 0.02fF
C219 VDD.n60 GND 0.02fF
C220 VDD.n61 GND 0.13fF
C221 VDD.n62 GND 0.16fF
C222 VDD.n63 GND 0.01fF
C223 VDD.n64 GND 0.02fF
C224 VDD.n65 GND 0.02fF
C225 VDD.n66 GND 0.06fF
C226 VDD.n67 GND 0.22fF
C227 VDD.n68 GND 0.01fF
C228 VDD.n69 GND 0.01fF
C229 VDD.n70 GND 0.02fF
C230 VDD.n71 GND 0.26fF
C231 VDD.n72 GND 0.01fF
C232 VDD.n73 GND 0.02fF
C233 VDD.n74 GND 0.02fF
C234 VDD.n75 GND 0.26fF
C235 VDD.n76 GND 0.01fF
C236 VDD.n77 GND 0.02fF
C237 VDD.n78 GND 0.03fF
C238 VDD.n79 GND 0.02fF
C239 VDD.n80 GND 0.02fF
C240 VDD.n81 GND 0.02fF
C241 VDD.n82 GND 0.30fF
C242 VDD.n83 GND 0.04fF
C243 VDD.n84 GND 0.03fF
C244 VDD.n85 GND 0.02fF
C245 VDD.n87 GND 0.02fF
C246 VDD.n88 GND 0.02fF
C247 VDD.n89 GND 0.02fF
C248 VDD.n90 GND 0.02fF
C249 VDD.n92 GND 0.02fF
C250 VDD.n93 GND 0.02fF
C251 VDD.n94 GND 0.02fF
C252 VDD.n96 GND 0.26fF
C253 VDD.n98 GND 0.02fF
C254 VDD.n99 GND 0.02fF
C255 VDD.n100 GND 0.03fF
C256 VDD.n101 GND 0.02fF
C257 VDD.n102 GND 0.26fF
C258 VDD.n103 GND 0.01fF
C259 VDD.n104 GND 0.02fF
C260 VDD.n105 GND 0.03fF
C261 VDD.n106 GND 0.26fF
C262 VDD.n107 GND 0.01fF
C263 VDD.n108 GND 0.02fF
C264 VDD.n109 GND 0.02fF
C265 VDD.n110 GND 0.21fF
C266 VDD.n111 GND 0.01fF
C267 VDD.n112 GND 0.06fF
C268 VDD.n113 GND 0.02fF
C269 VDD.n114 GND 0.13fF
C270 VDD.n115 GND 0.16fF
C271 VDD.n116 GND 0.01fF
C272 VDD.n117 GND 0.02fF
C273 VDD.n118 GND 0.02fF
C274 VDD.n119 GND 0.13fF
C275 VDD.n120 GND 0.15fF
C276 VDD.n121 GND 0.01fF
C277 VDD.n122 GND 0.10fF
C278 VDD.n123 GND 0.02fF
C279 VDD.n124 GND 0.02fF
C280 VDD.n125 GND 0.02fF
C281 VDD.n126 GND 0.17fF
C282 VDD.n127 GND 0.14fF
C283 VDD.n128 GND 0.01fF
C284 VDD.n129 GND 0.02fF
C285 VDD.n130 GND 0.03fF
C286 VDD.n131 GND 0.17fF
C287 VDD.n132 GND 0.14fF
C288 VDD.n133 GND 0.01fF
C289 VDD.n134 GND 0.02fF
C290 VDD.n135 GND 0.03fF
C291 VDD.n136 GND 0.10fF
C292 VDD.n137 GND 0.02fF
C293 VDD.n138 GND 0.13fF
C294 VDD.n139 GND 0.15fF
C295 VDD.n140 GND 0.01fF
C296 VDD.n141 GND 0.02fF
C297 VDD.n142 GND 0.02fF
C298 VDD.n143 GND 0.13fF
C299 VDD.n144 GND 0.16fF
C300 VDD.n145 GND 0.01fF
C301 VDD.n146 GND 0.02fF
C302 VDD.n147 GND 0.02fF
C303 VDD.n148 GND 0.06fF
C304 VDD.n149 GND 0.22fF
C305 VDD.n150 GND 0.01fF
C306 VDD.n151 GND 0.01fF
C307 VDD.n152 GND 0.02fF
C308 VDD.n153 GND 0.26fF
C309 VDD.n154 GND 0.01fF
C310 VDD.n155 GND 0.02fF
C311 VDD.n156 GND 0.02fF
C312 VDD.n157 GND 0.26fF
C313 VDD.n158 GND 0.01fF
C314 VDD.n159 GND 0.02fF
C315 VDD.n160 GND 0.03fF
C316 VDD.n161 GND 0.02fF
C317 VDD.n162 GND 0.02fF
C318 VDD.n163 GND 0.02fF
C319 VDD.n164 GND 0.30fF
C320 VDD.n165 GND 0.04fF
C321 VDD.n166 GND 0.03fF
C322 VDD.n167 GND 0.02fF
C323 VDD.n168 GND 0.02fF
C324 VDD.n169 GND 0.02fF
C325 VDD.n170 GND 0.02fF
C326 VDD.n171 GND 0.02fF
C327 VDD.n173 GND 0.02fF
C328 VDD.n174 GND 0.02fF
C329 VDD.n175 GND 0.02fF
C330 VDD.n177 GND 0.26fF
C331 VDD.n179 GND 0.02fF
C332 VDD.n180 GND 0.02fF
C333 VDD.n181 GND 0.03fF
C334 VDD.n182 GND 0.02fF
C335 VDD.n183 GND 0.26fF
C336 VDD.n184 GND 0.01fF
C337 VDD.n185 GND 0.02fF
C338 VDD.n186 GND 0.03fF
C339 VDD.n187 GND 0.26fF
C340 VDD.n188 GND 0.01fF
C341 VDD.n189 GND 0.02fF
C342 VDD.n190 GND 0.02fF
C343 VDD.n191 GND 0.21fF
C344 VDD.n192 GND 0.01fF
C345 VDD.n193 GND 0.06fF
C346 VDD.n194 GND 0.02fF
C347 VDD.n195 GND 0.13fF
C348 VDD.n196 GND 0.16fF
C349 VDD.n197 GND 0.01fF
C350 VDD.n198 GND 0.02fF
C351 VDD.n199 GND 0.02fF
C352 VDD.n200 GND 0.13fF
C353 VDD.n201 GND 0.15fF
C354 VDD.n202 GND 0.01fF
C355 VDD.n203 GND 0.10fF
C356 VDD.n204 GND 0.02fF
C357 VDD.n205 GND 0.02fF
C358 VDD.n206 GND 0.02fF
C359 VDD.n207 GND 0.17fF
C360 VDD.n208 GND 0.14fF
C361 VDD.n209 GND 0.01fF
C362 VDD.n210 GND 0.02fF
C363 VDD.n211 GND 0.03fF
C364 VDD.n212 GND 0.17fF
C365 VDD.n213 GND 0.14fF
C366 VDD.n214 GND 0.01fF
C367 VDD.n215 GND 0.02fF
C368 VDD.n216 GND 0.03fF
C369 VDD.n217 GND 0.10fF
C370 VDD.n218 GND 0.02fF
C371 VDD.n219 GND 0.13fF
C372 VDD.n220 GND 0.15fF
C373 VDD.n221 GND 0.01fF
C374 VDD.n222 GND 0.02fF
C375 VDD.n223 GND 0.02fF
C376 VDD.n224 GND 0.13fF
C377 VDD.n225 GND 0.16fF
C378 VDD.n226 GND 0.01fF
C379 VDD.n227 GND 0.02fF
C380 VDD.n228 GND 0.02fF
C381 VDD.n229 GND 0.06fF
C382 VDD.n230 GND 0.22fF
C383 VDD.n231 GND 0.01fF
C384 VDD.n232 GND 0.01fF
C385 VDD.n233 GND 0.02fF
C386 VDD.n234 GND 0.26fF
C387 VDD.n235 GND 0.01fF
C388 VDD.n236 GND 0.02fF
C389 VDD.n237 GND 0.02fF
C390 VDD.n238 GND 0.26fF
C391 VDD.n239 GND 0.01fF
C392 VDD.n240 GND 0.02fF
C393 VDD.n241 GND 0.02fF
C394 VDD.n242 GND 0.02fF
C395 VDD.n243 GND 0.02fF
C396 VDD.n244 GND 0.02fF
C397 VDD.n245 GND 0.19fF
C398 VDD.n246 GND 0.03fF
C399 VDD.n247 GND 0.02fF
C400 VDD.n248 GND 0.02fF
C401 VDD.n249 GND 0.02fF
C402 VDD.n250 GND 0.02fF
C403 VDD.n251 GND 0.02fF
C404 VDD.n253 GND 0.02fF
C405 VDD.n254 GND 0.02fF
C406 VDD.n255 GND 0.02fF
C407 VDD.n257 GND 0.44fF
C408 VDD.n259 GND 0.03fF
C409 VDD.n260 GND 0.03fF
C410 VDD.n261 GND 0.26fF
C411 VDD.n262 GND 0.02fF
C412 VDD.n263 GND 0.03fF
C413 VDD.n264 GND 0.03fF
C414 VDD.n265 GND 0.26fF
C415 VDD.n266 GND 0.01fF
C416 VDD.n267 GND 0.02fF
C417 VDD.n268 GND 0.02fF
C418 VDD.n269 GND 0.06fF
C419 VDD.n270 GND 0.22fF
C420 VDD.n271 GND 0.01fF
C421 VDD.n272 GND 0.01fF
C422 VDD.n273 GND 0.02fF
C423 VDD.n274 GND 0.13fF
C424 VDD.n275 GND 0.16fF
C425 VDD.n276 GND 0.01fF
C426 VDD.n277 GND 0.02fF
C427 VDD.n278 GND 0.02fF
C428 VDD.n279 GND 0.10fF
C429 VDD.n280 GND 0.02fF
C430 VDD.n281 GND 0.13fF
C431 VDD.n282 GND 0.15fF
C432 VDD.n283 GND 0.01fF
C433 VDD.n284 GND 0.02fF
C434 VDD.n285 GND 0.02fF
C435 VDD.n286 GND 0.17fF
C436 VDD.n287 GND 0.14fF
C437 VDD.n288 GND 0.01fF
C438 VDD.n289 GND 0.02fF
C439 VDD.n290 GND 0.03fF
C440 VDD.n291 GND 0.17fF
C441 VDD.n292 GND 0.14fF
C442 VDD.n293 GND 0.01fF
C443 VDD.n294 GND 0.02fF
C444 VDD.n295 GND 0.03fF
C445 VDD.n296 GND 0.13fF
C446 VDD.n297 GND 0.15fF
C447 VDD.n298 GND 0.01fF
C448 VDD.n299 GND 0.10fF
C449 VDD.n300 GND 0.02fF
C450 VDD.n301 GND 0.02fF
C451 VDD.n302 GND 0.02fF
C452 VDD.n303 GND 0.13fF
C453 VDD.n304 GND 0.16fF
C454 VDD.n305 GND 0.01fF
C455 VDD.n306 GND 0.02fF
C456 VDD.n307 GND 0.02fF
C457 VDD.n308 GND 0.21fF
C458 VDD.n309 GND 0.01fF
C459 VDD.n310 GND 0.06fF
C460 VDD.n311 GND 0.02fF
C461 VDD.n312 GND 0.26fF
C462 VDD.n313 GND 0.01fF
C463 VDD.n314 GND 0.02fF
C464 VDD.n315 GND 0.02fF
C465 VDD.n316 GND 0.26fF
C466 VDD.n317 GND 0.01fF
C467 VDD.n318 GND 0.02fF
C468 VDD.n319 GND 0.03fF
C469 VDD.n320 GND 0.02fF
C470 VDD.n321 GND 0.02fF
C471 VDD.n322 GND 0.02fF
C472 VDD.n323 GND 0.02fF
C473 VDD.n324 GND 0.02fF
C474 VDD.n325 GND 0.02fF
C475 VDD.n327 GND 0.02fF
C476 VDD.n328 GND 0.02fF
C477 VDD.n329 GND 0.02fF
C478 VDD.n330 GND 0.02fF
C479 VDD.n332 GND 0.03fF
C480 VDD.n333 GND 0.02fF
C481 VDD.n334 GND 0.30fF
C482 VDD.n335 GND 0.04fF
C483 VDD.n337 GND 0.26fF
C484 VDD.n339 GND 0.02fF
C485 VDD.n340 GND 0.02fF
C486 VDD.n341 GND 0.03fF
C487 VDD.n342 GND 0.02fF
C488 VDD.n343 GND 0.26fF
C489 VDD.n344 GND 0.01fF
C490 VDD.n345 GND 0.02fF
C491 VDD.n346 GND 0.03fF
C492 VDD.n347 GND 0.26fF
C493 VDD.n348 GND 0.01fF
C494 VDD.n349 GND 0.02fF
C495 VDD.n350 GND 0.02fF
C496 VDD.n351 GND 0.06fF
C497 VDD.n352 GND 0.22fF
C498 VDD.n353 GND 0.01fF
C499 VDD.n354 GND 0.01fF
C500 VDD.n355 GND 0.02fF
C501 VDD.n356 GND 0.13fF
C502 VDD.n357 GND 0.16fF
C503 VDD.n358 GND 0.01fF
C504 VDD.n359 GND 0.02fF
C505 VDD.n360 GND 0.02fF
C506 VDD.n361 GND 0.10fF
C507 VDD.n362 GND 0.02fF
C508 VDD.n363 GND 0.13fF
C509 VDD.n364 GND 0.15fF
C510 VDD.n365 GND 0.01fF
C511 VDD.n366 GND 0.02fF
C512 VDD.n367 GND 0.02fF
C513 VDD.n368 GND 0.17fF
C514 VDD.n369 GND 0.14fF
C515 VDD.n370 GND 0.01fF
C516 VDD.n371 GND 0.02fF
C517 VDD.n372 GND 0.03fF
C518 VDD.n373 GND 0.17fF
C519 VDD.n374 GND 0.14fF
C520 VDD.n375 GND 0.01fF
C521 VDD.n376 GND 0.02fF
C522 VDD.n377 GND 0.03fF
C523 VDD.n378 GND 0.13fF
C524 VDD.n379 GND 0.15fF
C525 VDD.n380 GND 0.01fF
C526 VDD.n381 GND 0.10fF
C527 VDD.n382 GND 0.02fF
C528 VDD.n383 GND 0.02fF
C529 VDD.n384 GND 0.02fF
C530 VDD.n385 GND 0.13fF
C531 VDD.n386 GND 0.16fF
C532 VDD.n387 GND 0.01fF
C533 VDD.n388 GND 0.02fF
C534 VDD.n389 GND 0.02fF
C535 VDD.n390 GND 0.21fF
C536 VDD.n391 GND 0.01fF
C537 VDD.n392 GND 0.06fF
C538 VDD.n393 GND 0.02fF
C539 VDD.n394 GND 0.26fF
C540 VDD.n395 GND 0.01fF
C541 VDD.n396 GND 0.02fF
C542 VDD.n397 GND 0.02fF
C543 VDD.n398 GND 0.26fF
C544 VDD.n399 GND 0.01fF
C545 VDD.n400 GND 0.02fF
C546 VDD.n401 GND 0.03fF
C547 VDD.n402 GND 0.02fF
C548 VDD.n403 GND 0.02fF
C549 VDD.n404 GND 0.02fF
C550 VDD.n405 GND 0.30fF
C551 VDD.n406 GND 0.04fF
C552 VDD.n407 GND 0.03fF
C553 VDD.n408 GND 0.02fF
C554 VDD.n409 GND 0.02fF
C555 VDD.n410 GND 0.02fF
C556 VDD.n411 GND 0.02fF
C557 VDD.n412 GND 0.02fF
C558 VDD.n414 GND 0.02fF
C559 VDD.n415 GND 0.02fF
C560 VDD.n416 GND 0.02fF
C561 VDD.n418 GND 0.26fF
C562 VDD.n420 GND 0.02fF
C563 VDD.n421 GND 0.02fF
C564 VDD.n422 GND 0.03fF
C565 VDD.n423 GND 0.02fF
C566 VDD.n424 GND 0.26fF
C567 VDD.n425 GND 0.01fF
C568 VDD.n426 GND 0.02fF
C569 VDD.n427 GND 0.03fF
C570 VDD.n428 GND 0.26fF
C571 VDD.n429 GND 0.01fF
C572 VDD.n430 GND 0.02fF
C573 VDD.n431 GND 0.02fF
C574 VDD.n432 GND 0.06fF
C575 VDD.n433 GND 0.22fF
C576 VDD.n434 GND 0.01fF
C577 VDD.n435 GND 0.01fF
C578 VDD.n436 GND 0.02fF
C579 VDD.n437 GND 0.13fF
C580 VDD.n438 GND 0.16fF
C581 VDD.n439 GND 0.01fF
C582 VDD.n440 GND 0.02fF
C583 VDD.n441 GND 0.02fF
C584 VDD.n442 GND 0.10fF
C585 VDD.n443 GND 0.02fF
C586 VDD.n444 GND 0.13fF
C587 VDD.n445 GND 0.15fF
C588 VDD.n446 GND 0.01fF
C589 VDD.n447 GND 0.02fF
C590 VDD.n448 GND 0.02fF
C591 VDD.n449 GND 0.17fF
C592 VDD.n450 GND 0.14fF
C593 VDD.n451 GND 0.01fF
C594 VDD.n452 GND 0.02fF
C595 VDD.n453 GND 0.03fF
C596 VDD.n454 GND 0.17fF
C597 VDD.n455 GND 0.14fF
C598 VDD.n456 GND 0.01fF
C599 VDD.n457 GND 0.02fF
C600 VDD.n458 GND 0.03fF
C601 VDD.n459 GND 0.13fF
C602 VDD.n460 GND 0.15fF
C603 VDD.n461 GND 0.01fF
C604 VDD.n462 GND 0.10fF
C605 VDD.n463 GND 0.02fF
C606 VDD.n464 GND 0.02fF
C607 VDD.n465 GND 0.02fF
C608 VDD.n466 GND 0.13fF
C609 VDD.n467 GND 0.16fF
C610 VDD.n468 GND 0.01fF
C611 VDD.n469 GND 0.02fF
C612 VDD.n470 GND 0.02fF
C613 VDD.n471 GND 0.21fF
C614 VDD.n472 GND 0.01fF
C615 VDD.n473 GND 0.06fF
C616 VDD.n474 GND 0.02fF
C617 VDD.n475 GND 0.26fF
C618 VDD.n476 GND 0.01fF
C619 VDD.n477 GND 0.02fF
C620 VDD.n478 GND 0.02fF
C621 VDD.n479 GND 0.02fF
C622 VDD.n480 GND 0.02fF
C623 VDD.n481 GND 0.02fF
C624 VDD.n482 GND 0.30fF
C625 VDD.n483 GND 0.04fF
C626 VDD.n484 GND 0.03fF
C627 VDD.n485 GND 0.02fF
C628 VDD.n486 GND 0.02fF
C629 VDD.n487 GND 0.02fF
C630 VDD.n488 GND 0.02fF
C631 VDD.n489 GND 0.02fF
C632 VDD.n491 GND 0.02fF
C633 VDD.n492 GND 0.02fF
C634 VDD.n493 GND 0.02fF
C635 VDD.n495 GND 0.26fF
C636 VDD.n497 GND 0.02fF
C637 VDD.n498 GND 0.02fF
C638 VDD.n499 GND 0.03fF
C639 VDD.n500 GND 0.02fF
C640 VDD.n501 GND 0.26fF
C641 VDD.n502 GND 0.01fF
C642 VDD.n503 GND 0.02fF
C643 VDD.n504 GND 0.02fF
C644 a_1561_989.n0 GND 0.76fF
C645 a_1561_989.n1 GND 0.76fF
C646 a_1561_989.n2 GND 0.89fF
C647 a_1561_989.n3 GND 0.28fF
C648 a_1561_989.n4 GND 0.39fF
C649 a_1561_989.n5 GND 0.49fF
C650 a_1561_989.n6 GND 0.61fF
C651 a_1561_989.n7 GND 0.49fF
C652 a_1561_989.t9 GND 0.79fF
C653 a_1561_989.n8 GND 0.52fF
C654 a_1561_989.n9 GND 0.49fF
C655 a_1561_989.t10 GND 0.79fF
C656 a_1561_989.n10 GND 0.55fF
C657 a_1561_989.n11 GND 1.78fF
C658 a_1561_989.n12 GND 2.66fF
C659 a_1561_989.n13 GND 0.65fF
C660 a_1561_989.n14 GND 0.12fF
C661 a_1561_989.n15 GND 0.46fF
C662 a_1561_989.n16 GND 0.06fF
C663 a_2201_1050.n0 GND 0.52fF
C664 a_2201_1050.n1 GND 0.52fF
C665 a_2201_1050.n2 GND 0.62fF
C666 a_2201_1050.n3 GND 0.19fF
C667 a_2201_1050.n4 GND 0.36fF
C668 a_2201_1050.n5 GND 0.39fF
C669 a_2201_1050.n6 GND 0.63fF
C670 a_2201_1050.n7 GND 0.62fF
C671 a_2201_1050.n8 GND 0.08fF
C672 a_2201_1050.n9 GND 0.22fF
C673 a_2201_1050.n10 GND 0.04fF
C674 a_4901_103.n0 GND 0.03fF
C675 a_4901_103.n1 GND 0.10fF
C676 a_4901_103.n2 GND 0.10fF
C677 a_4901_103.n3 GND 0.05fF
C678 a_4901_103.n4 GND 0.03fF
C679 a_4901_103.n5 GND 0.04fF
C680 a_4901_103.n6 GND 0.03fF
C681 a_4901_103.n7 GND 0.04fF
C682 a_4125_1050.n0 GND 0.47fF
C683 a_4125_1050.n1 GND 0.47fF
C684 a_4125_1050.n2 GND 0.55fF
C685 a_4125_1050.n3 GND 0.17fF
C686 a_4125_1050.n4 GND 0.29fF
C687 a_4125_1050.n5 GND 0.32fF
C688 a_4125_1050.n6 GND 0.57fF
C689 a_4125_1050.n7 GND 0.55fF
C690 a_4125_1050.n8 GND 0.07fF
C691 a_4125_1050.n9 GND 0.23fF
C692 a_4125_1050.n10 GND 0.04fF
C693 a_3258_210.n0 GND 0.07fF
C694 a_3258_210.n1 GND 0.13fF
C695 a_3258_210.n2 GND 0.07fF
C696 a_3258_210.n3 GND 0.02fF
C697 a_3258_210.n4 GND 0.03fF
C698 a_3258_210.n5 GND 0.06fF
C699 a_3258_210.n6 GND 0.05fF
C700 a_3258_210.n7 GND 0.06fF
C701 a_3258_210.n8 GND 0.07fF
C702 a_3258_210.n9 GND 0.07fF
C703 a_3258_210.n10 GND 0.03fF
C704 a_3258_210.n11 GND 0.01fF
C705 a_3258_210.n12 GND 0.12fF
C706 a_3258_210.t0 GND 0.28fF
C707 a_2977_103.n0 GND 0.03fF
C708 a_2977_103.n1 GND 0.10fF
C709 a_2977_103.n2 GND 0.10fF
C710 a_2977_103.n3 GND 0.05fF
C711 a_2977_103.n4 GND 0.03fF
C712 a_2977_103.n5 GND 0.04fF
C713 a_2977_103.n6 GND 0.11fF
C714 a_2977_103.n7 GND 0.04fF
.ends
