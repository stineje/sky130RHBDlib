* SPICE3 file created from NAND3X1.ext - technology: sky130A

.subckt NAND3X1 Y A B C VPB VNB
M1000 VPB.t3 a_147_159# a_277_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VPB.t5 a_342_166# a_277_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VNB a_147_159# a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1003 VPB.t1 a_599_943# a_277_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_277_1004.t3 a_147_159# VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_277_1004.t5 a_342_166# VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_277_1004.t0 a_599_943# VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 a_147_159# VPB 0.08fF
C1 a_342_166# VPB 0.05fF
C2 a_147_159# a_599_943# 0.02fF
C3 a_342_166# a_599_943# 0.18fF
C4 VPB a_599_943# 0.06fF
C5 a_342_166# a_147_159# 0.18fF
R0 a_277_1004.n7 a_277_1004.n5 377.444
R1 a_277_1004.n4 a_277_1004.n3 79.232
R2 a_277_1004.n5 a_277_1004.n4 63.152
R3 a_277_1004.n7 a_277_1004.n6 30
R4 a_277_1004.n8 a_277_1004.n0 24.383
R5 a_277_1004.n8 a_277_1004.n7 23.684
R6 a_277_1004.n5 a_277_1004.n1 16.08
R7 a_277_1004.n4 a_277_1004.n2 16.08
R8 a_277_1004.n1 a_277_1004.t2 14.282
R9 a_277_1004.n1 a_277_1004.t0 14.282
R10 a_277_1004.n2 a_277_1004.t6 14.282
R11 a_277_1004.n2 a_277_1004.t5 14.282
R12 a_277_1004.n3 a_277_1004.t4 14.282
R13 a_277_1004.n3 a_277_1004.t3 14.282
R14 VPB VPB.n98 126.832
R15 VPB.n54 VPB.n53 80.104
R16 VPB.n84 VPB.n83 76
R17 VPB.n91 VPB.n90 76
R18 VPB.n68 VPB.n67 75.654
R19 VPB.n63 VPB.t2 55.106
R20 VPB.n49 VPB.t1 55.106
R21 VPB.n58 VPB.n57 48.952
R22 VPB.n72 VPB.n71 44.502
R23 VPB.n75 VPB.n62 40.824
R24 VPB.n61 VPB.n20 40.824
R25 VPB.n95 VPB.n91 20.452
R26 VPB.n44 VPB.n41 20.452
R27 VPB.n81 VPB.n80 17.801
R28 VPB.n62 VPB.t4 14.282
R29 VPB.n62 VPB.t3 14.282
R30 VPB.n20 VPB.t0 14.282
R31 VPB.n20 VPB.t5 14.282
R32 VPB.n44 VPB.n43 13.653
R33 VPB.n43 VPB.n42 13.653
R34 VPB.n48 VPB.n47 13.653
R35 VPB.n47 VPB.n46 13.653
R36 VPB.n52 VPB.n51 13.653
R37 VPB.n51 VPB.n50 13.653
R38 VPB.n56 VPB.n55 13.653
R39 VPB.n55 VPB.n54 13.653
R40 VPB.n60 VPB.n59 13.653
R41 VPB.n59 VPB.n58 13.653
R42 VPB.n83 VPB.n82 13.653
R43 VPB.n82 VPB.n81 13.653
R44 VPB.n79 VPB.n78 13.653
R45 VPB.n78 VPB.n77 13.653
R46 VPB.n74 VPB.n73 13.653
R47 VPB.n73 VPB.n72 13.653
R48 VPB.n70 VPB.n69 13.653
R49 VPB.n69 VPB.n68 13.653
R50 VPB.n66 VPB.n65 13.653
R51 VPB.n65 VPB.n64 13.653
R52 VPB.n16 VPB.n15 13.653
R53 VPB.n15 VPB.n14 13.653
R54 VPB.n91 VPB.n0 13.653
R55 VPB VPB.n0 13.653
R56 VPB.n77 VPB.n76 13.35
R57 VPB.n95 VPB.n94 13.276
R58 VPB.n94 VPB.n92 13.276
R59 VPB.n56 VPB.n52 13.276
R60 VPB.n60 VPB.n56 13.276
R61 VPB.n83 VPB.n79 13.276
R62 VPB.n74 VPB.n70 13.276
R63 VPB.n70 VPB.n66 13.276
R64 VPB.n91 VPB.n16 13.276
R65 VPB.n41 VPB.n23 13.276
R66 VPB.n23 VPB.n21 13.276
R67 VPB.n28 VPB.n26 12.796
R68 VPB.n28 VPB.n27 12.564
R69 VPB.n63 VPB.n16 12.558
R70 VPB.n49 VPB.n48 12.2
R71 VPB.n37 VPB.n36 12.198
R72 VPB.n34 VPB.n33 12.198
R73 VPB.n31 VPB.n30 12.198
R74 VPB.n83 VPB.n61 9.329
R75 VPB.n79 VPB.n75 8.97
R76 VPB.n41 VPB.n40 7.5
R77 VPB.n26 VPB.n25 7.5
R78 VPB.n30 VPB.n29 7.5
R79 VPB.n33 VPB.n32 7.5
R80 VPB.n23 VPB.n22 7.5
R81 VPB.n38 VPB.n24 7.5
R82 VPB.n94 VPB.n93 7.5
R83 VPB.n12 VPB.n11 7.5
R84 VPB.n6 VPB.n5 7.5
R85 VPB.n8 VPB.n7 7.5
R86 VPB.n2 VPB.n1 7.5
R87 VPB.n96 VPB.n95 7.5
R88 VPB.n13 VPB.n10 6.729
R89 VPB.n9 VPB.n6 6.729
R90 VPB.n4 VPB.n2 6.729
R91 VPB.n4 VPB.n3 6.728
R92 VPB.n9 VPB.n8 6.728
R93 VPB.n13 VPB.n12 6.728
R94 VPB.n97 VPB.n96 6.728
R95 VPB.n40 VPB.n39 6.398
R96 VPB.n45 VPB.n44 6.112
R97 VPB.n48 VPB.n45 6.101
R98 VPB.n75 VPB.n74 4.305
R99 VPB.n61 VPB.n60 3.947
R100 VPB.n38 VPB.n31 1.402
R101 VPB.n38 VPB.n34 1.402
R102 VPB.n38 VPB.n35 1.402
R103 VPB.n38 VPB.n37 1.402
R104 VPB.n52 VPB.n49 1.076
R105 VPB.n39 VPB.n38 0.735
R106 VPB.n38 VPB.n28 0.735
R107 VPB.n66 VPB.n63 0.717
R108 VPB.n98 VPB.n13 0.387
R109 VPB.n98 VPB.n9 0.387
R110 VPB.n98 VPB.n4 0.387
R111 VPB.n98 VPB.n97 0.387
R112 VPB.n90 VPB 0.198
R113 VPB.n18 VPB.n17 0.136
R114 VPB.n19 VPB.n18 0.136
R115 VPB.n84 VPB.n19 0.136
R116 VPB.n86 VPB.n85 0.136
R117 VPB.n87 VPB.n86 0.136
R118 VPB.n88 VPB.n87 0.136
R119 VPB.n89 VPB.n88 0.136
R120 VPB.n90 VPB.n89 0.136
R121 VPB VPB.n84 0.068
R122 VPB.n85 VPB 0.068
R123 a_91_75.t0 a_91_75.n3 117.777
R124 a_91_75.n6 a_91_75.n5 45.444
R125 a_91_75.t0 a_91_75.n6 21.213
R126 a_91_75.t0 a_91_75.n4 11.595
R127 a_91_75.n2 a_91_75.n0 8.543
R128 a_91_75.t0 a_91_75.n2 3.034
R129 a_91_75.n2 a_91_75.n1 0.443
R130 a_372_182.n8 a_372_182.n6 96.467
R131 a_372_182.n3 a_372_182.n1 44.628
R132 a_372_182.t0 a_372_182.n8 32.417
R133 a_372_182.n3 a_372_182.n2 23.284
R134 a_372_182.n6 a_372_182.n5 22.349
R135 a_372_182.t0 a_372_182.n10 20.241
R136 a_372_182.n10 a_372_182.n9 13.494
R137 a_372_182.n6 a_372_182.n4 8.443
R138 a_372_182.t0 a_372_182.n0 8.137
R139 a_372_182.t0 a_372_182.n3 5.727
R140 a_372_182.n8 a_372_182.n7 1.435
R141 VNB VNB.n78 300.778
R142 VNB.n42 VNB.n41 85.559
R143 VNB.n65 VNB.n64 76
R144 VNB.n58 VNB.n57 76
R145 VNB.n44 VNB.n43 41.971
R146 VNB.n27 VNB.n24 20.452
R147 VNB.n66 VNB.n65 20.452
R148 VNB.n31 VNB.n30 13.653
R149 VNB.n30 VNB.n29 13.653
R150 VNB.n34 VNB.n33 13.653
R151 VNB.n33 VNB.n32 13.653
R152 VNB.n37 VNB.n36 13.653
R153 VNB.n36 VNB.n35 13.653
R154 VNB.n40 VNB.n39 13.653
R155 VNB.n39 VNB.n38 13.653
R156 VNB.n57 VNB.n56 13.653
R157 VNB.n56 VNB.n55 13.653
R158 VNB.n54 VNB.n53 13.653
R159 VNB.n53 VNB.n52 13.653
R160 VNB.n51 VNB.n50 13.653
R161 VNB.n50 VNB.n49 13.653
R162 VNB.n48 VNB.n47 13.653
R163 VNB.n47 VNB.n46 13.653
R164 VNB.n45 VNB.n44 13.653
R165 VNB.n6 VNB.n5 13.653
R166 VNB.n5 VNB.n4 13.653
R167 VNB.n65 VNB.n0 13.653
R168 VNB VNB.n0 13.653
R169 VNB.n27 VNB.n26 13.653
R170 VNB.n26 VNB.n25 13.653
R171 VNB.n73 VNB.n70 13.577
R172 VNB.n12 VNB.n10 13.276
R173 VNB.n24 VNB.n12 13.276
R174 VNB.n34 VNB.n31 13.276
R175 VNB.n37 VNB.n34 13.276
R176 VNB.n40 VNB.n37 13.276
R177 VNB.n57 VNB.n40 13.276
R178 VNB.n57 VNB.n54 13.276
R179 VNB.n54 VNB.n51 13.276
R180 VNB.n51 VNB.n48 13.276
R181 VNB.n48 VNB.n45 13.276
R182 VNB.n65 VNB.n6 13.276
R183 VNB.n3 VNB.n1 13.276
R184 VNB.n66 VNB.n3 13.276
R185 VNB.n42 VNB.n6 12.02
R186 VNB.n75 VNB.n74 7.5
R187 VNB.n67 VNB.n66 7.5
R188 VNB.n3 VNB.n2 7.5
R189 VNB.n72 VNB.n71 7.5
R190 VNB.n18 VNB.n17 7.5
R191 VNB.n14 VNB.n13 7.5
R192 VNB.n12 VNB.n11 7.5
R193 VNB.n24 VNB.n23 7.5
R194 VNB.n77 VNB.n75 7.011
R195 VNB.n20 VNB.n18 7.011
R196 VNB.n16 VNB.n14 7.011
R197 VNB.n23 VNB.n22 7.01
R198 VNB.n16 VNB.n15 7.01
R199 VNB.n20 VNB.n19 7.01
R200 VNB.n77 VNB.n76 7.01
R201 VNB.n73 VNB.n72 6.788
R202 VNB.n68 VNB.n67 6.788
R203 VNB.n28 VNB.n27 6.111
R204 VNB.n31 VNB.n28 6.1
R205 VNB.n45 VNB.n42 1.255
R206 VNB.n78 VNB.n69 0.921
R207 VNB.n78 VNB.n73 0.476
R208 VNB.n78 VNB.n68 0.475
R209 VNB.n21 VNB.n16 0.246
R210 VNB.n22 VNB.n21 0.246
R211 VNB.n21 VNB.n20 0.246
R212 VNB.n78 VNB.n77 0.246
R213 VNB.n64 VNB 0.198
R214 VNB.n8 VNB.n7 0.136
R215 VNB.n9 VNB.n8 0.136
R216 VNB.n58 VNB.n9 0.136
R217 VNB.n60 VNB.n59 0.136
R218 VNB.n61 VNB.n60 0.136
R219 VNB.n62 VNB.n61 0.136
R220 VNB.n63 VNB.n62 0.136
R221 VNB.n64 VNB.n63 0.136
R222 VNB VNB.n58 0.068
R223 VNB.n59 VNB 0.068
C6 VPB VNB 4.63fF
C7 a_372_182.n0 VNB 0.07fF
C8 a_372_182.n1 VNB 0.09fF
C9 a_372_182.n2 VNB 0.13fF
C10 a_372_182.n3 VNB 0.11fF
C11 a_372_182.n4 VNB 0.02fF
C12 a_372_182.n5 VNB 0.03fF
C13 a_372_182.n6 VNB 0.06fF
C14 a_372_182.n7 VNB 0.03fF
C15 a_372_182.n8 VNB 0.12fF
C16 a_372_182.n9 VNB 0.05fF
C17 a_372_182.n10 VNB 0.01fF
C18 a_372_182.t0 VNB 0.32fF
C19 a_91_75.n0 VNB 0.19fF
C20 a_91_75.n1 VNB 0.04fF
C21 a_91_75.n2 VNB 0.01fF
C22 a_91_75.n3 VNB 0.03fF
C23 a_91_75.n4 VNB 0.05fF
C24 a_91_75.n5 VNB 0.08fF
C25 a_91_75.n6 VNB 0.07fF
C26 VPB.n0 VNB 0.03fF
C27 VPB.n1 VNB 0.03fF
C28 VPB.n2 VNB 0.02fF
C29 VPB.n3 VNB 0.17fF
C30 VPB.n5 VNB 0.02fF
C31 VPB.n6 VNB 0.02fF
C32 VPB.n7 VNB 0.02fF
C33 VPB.n8 VNB 0.02fF
C34 VPB.n10 VNB 0.02fF
C35 VPB.n11 VNB 0.02fF
C36 VPB.n12 VNB 0.02fF
C37 VPB.n14 VNB 0.25fF
C38 VPB.n15 VNB 0.02fF
C39 VPB.n16 VNB 0.02fF
C40 VPB.n17 VNB 0.09fF
C41 VPB.n18 VNB 0.02fF
C42 VPB.n19 VNB 0.02fF
C43 VPB.n20 VNB 0.09fF
C44 VPB.n21 VNB 0.02fF
C45 VPB.n22 VNB 0.02fF
C46 VPB.n23 VNB 0.02fF
C47 VPB.n24 VNB 0.17fF
C48 VPB.n25 VNB 0.02fF
C49 VPB.n26 VNB 0.02fF
C50 VPB.n27 VNB 0.04fF
C51 VPB.n28 VNB 0.01fF
C52 VPB.n29 VNB 0.02fF
C53 VPB.n30 VNB 0.02fF
C54 VPB.n32 VNB 0.02fF
C55 VPB.n33 VNB 0.02fF
C56 VPB.n36 VNB 0.02fF
C57 VPB.n38 VNB 0.42fF
C58 VPB.n40 VNB 0.03fF
C59 VPB.n41 VNB 0.03fF
C60 VPB.n42 VNB 0.25fF
C61 VPB.n43 VNB 0.03fF
C62 VPB.n44 VNB 0.03fF
C63 VPB.n45 VNB 0.00fF
C64 VPB.n46 VNB 0.25fF
C65 VPB.n47 VNB 0.02fF
C66 VPB.n48 VNB 0.02fF
C67 VPB.n49 VNB 0.05fF
C68 VPB.n50 VNB 0.19fF
C69 VPB.n51 VNB 0.02fF
C70 VPB.n52 VNB 0.01fF
C71 VPB.n53 VNB 0.12fF
C72 VPB.n54 VNB 0.15fF
C73 VPB.n55 VNB 0.02fF
C74 VPB.n56 VNB 0.02fF
C75 VPB.n57 VNB 0.12fF
C76 VPB.n58 VNB 0.15fF
C77 VPB.n59 VNB 0.02fF
C78 VPB.n60 VNB 0.01fF
C79 VPB.n61 VNB 0.02fF
C80 VPB.n62 VNB 0.09fF
C81 VPB.n63 VNB 0.05fF
C82 VPB.n64 VNB 0.19fF
C83 VPB.n65 VNB 0.02fF
C84 VPB.n66 VNB 0.01fF
C85 VPB.n67 VNB 0.12fF
C86 VPB.n68 VNB 0.15fF
C87 VPB.n69 VNB 0.02fF
C88 VPB.n70 VNB 0.02fF
C89 VPB.n71 VNB 0.12fF
C90 VPB.n72 VNB 0.15fF
C91 VPB.n73 VNB 0.02fF
C92 VPB.n74 VNB 0.01fF
C93 VPB.n75 VNB 0.02fF
C94 VPB.n76 VNB 0.12fF
C95 VPB.n77 VNB 0.13fF
C96 VPB.n78 VNB 0.02fF
C97 VPB.n79 VNB 0.02fF
C98 VPB.n80 VNB 0.12fF
C99 VPB.n81 VNB 0.14fF
C100 VPB.n82 VNB 0.02fF
C101 VPB.n83 VNB 0.02fF
C102 VPB.n84 VNB 0.02fF
C103 VPB.n85 VNB 0.02fF
C104 VPB.n86 VNB 0.02fF
C105 VPB.n87 VNB 0.02fF
C106 VPB.n88 VNB 0.02fF
C107 VPB.n89 VNB 0.02fF
C108 VPB.n90 VNB 0.03fF
C109 VPB.n91 VNB 0.03fF
C110 VPB.n92 VNB 0.02fF
C111 VPB.n93 VNB 0.02fF
C112 VPB.n94 VNB 0.02fF
C113 VPB.n95 VNB 0.03fF
C114 VPB.n96 VNB 0.03fF
C115 VPB.n98 VNB 0.39fF
C116 a_277_1004.n0 VNB 0.03fF
C117 a_277_1004.n1 VNB 0.42fF
C118 a_277_1004.n2 VNB 0.42fF
C119 a_277_1004.n3 VNB 0.49fF
C120 a_277_1004.n4 VNB 0.15fF
C121 a_277_1004.n5 VNB 0.43fF
C122 a_277_1004.n6 VNB 0.03fF
C123 a_277_1004.n7 VNB 0.38fF
C124 a_277_1004.n8 VNB 0.04fF
.ends
