// File: DFFQX1.spi.DFFQX1.pxi
// Created: Tue Oct 15 15:46:01 2024
// 
simulator lang=spectre
x_PM_DFFQX1\%GND ( GND N_GND_c_8_p N_GND_c_117_p N_GND_c_1_p N_GND_c_9_p \
 N_GND_c_10_p N_GND_c_11_p N_GND_c_16_p N_GND_c_30_p N_GND_c_38_p N_GND_c_51_p \
 N_GND_c_75_p N_GND_c_82_p N_GND_c_88_p N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p \
 N_GND_c_5_p N_GND_c_6_p N_GND_c_7_p N_GND_M0_noxref_d N_GND_M3_noxref_d \
 N_GND_M5_noxref_d N_GND_M7_noxref_d N_GND_M9_noxref_d N_GND_M11_noxref_d )  \
 PM_DFFQX1\%GND
x_PM_DFFQX1\%VDD ( VDD N_VDD_c_272_p N_VDD_c_264_n N_VDD_c_372_p N_VDD_c_361_p \
 N_VDD_c_287_p N_VDD_c_339_p N_VDD_c_340_p N_VDD_c_273_p N_VDD_c_274_p \
 N_VDD_c_342_p N_VDD_c_343_p N_VDD_c_285_p N_VDD_c_309_p N_VDD_c_345_p \
 N_VDD_c_346_p N_VDD_c_320_p N_VDD_c_365_p N_VDD_c_458_p N_VDD_c_459_p \
 N_VDD_c_390_p N_VDD_c_419_p N_VDD_c_461_p N_VDD_c_462_p N_VDD_c_430_p \
 N_VDD_c_500_p N_VDD_c_265_n N_VDD_c_266_n N_VDD_c_267_n N_VDD_c_268_n \
 N_VDD_c_269_n N_VDD_c_270_n N_VDD_M13_noxref_s N_VDD_M14_noxref_d \
 N_VDD_M16_noxref_d N_VDD_M18_noxref_d N_VDD_M19_noxref_s N_VDD_M20_noxref_d \
 N_VDD_M22_noxref_d N_VDD_M23_noxref_s N_VDD_M24_noxref_d N_VDD_M26_noxref_d \
 N_VDD_M27_noxref_s N_VDD_M28_noxref_d N_VDD_M30_noxref_d N_VDD_M31_noxref_s \
 N_VDD_M32_noxref_d N_VDD_M34_noxref_d N_VDD_M35_noxref_s N_VDD_M36_noxref_d \
 N_VDD_M38_noxref_d )  PM_DFFQX1\%VDD
x_PM_DFFQX1\%noxref_3 ( N_noxref_3_c_555_n N_noxref_3_c_560_n \
 N_noxref_3_c_561_n N_noxref_3_c_565_n N_noxref_3_c_566_n N_noxref_3_c_584_n \
 N_noxref_3_c_588_n N_noxref_3_c_590_n N_noxref_3_c_567_n N_noxref_3_c_764_p \
 N_noxref_3_c_568_n N_noxref_3_c_569_n N_noxref_3_c_751_p \
 N_noxref_3_M2_noxref_g N_noxref_3_M5_noxref_g N_noxref_3_M17_noxref_g \
 N_noxref_3_M18_noxref_g N_noxref_3_M23_noxref_g N_noxref_3_M24_noxref_g \
 N_noxref_3_c_644_p N_noxref_3_c_645_p N_noxref_3_c_646_p N_noxref_3_c_688_p \
 N_noxref_3_c_665_p N_noxref_3_c_690_p N_noxref_3_c_666_p N_noxref_3_c_570_n \
 N_noxref_3_c_572_n N_noxref_3_c_573_n N_noxref_3_c_574_n N_noxref_3_c_575_n \
 N_noxref_3_c_576_n N_noxref_3_c_577_n N_noxref_3_c_579_n N_noxref_3_c_639_p \
 N_noxref_3_c_649_p N_noxref_3_c_634_p N_noxref_3_c_607_n \
 N_noxref_3_M4_noxref_d N_noxref_3_M19_noxref_d N_noxref_3_M21_noxref_d )  \
 PM_DFFQX1\%noxref_3
x_PM_DFFQX1\%noxref_4 ( N_noxref_4_c_787_n N_noxref_4_c_791_n \
 N_noxref_4_c_808_n N_noxref_4_c_812_n N_noxref_4_c_814_n N_noxref_4_c_792_n \
 N_noxref_4_c_877_p N_noxref_4_c_793_n N_noxref_4_c_794_n N_noxref_4_c_904_p \
 N_noxref_4_M7_noxref_g N_noxref_4_M27_noxref_g N_noxref_4_M28_noxref_g \
 N_noxref_4_c_795_n N_noxref_4_c_797_n N_noxref_4_c_798_n N_noxref_4_c_799_n \
 N_noxref_4_c_800_n N_noxref_4_c_801_n N_noxref_4_c_802_n N_noxref_4_c_804_n \
 N_noxref_4_c_827_n N_noxref_4_M6_noxref_d N_noxref_4_M23_noxref_d \
 N_noxref_4_M25_noxref_d )  PM_DFFQX1\%noxref_4
x_PM_DFFQX1\%CLK ( N_CLK_c_940_n N_CLK_c_958_n CLK CLK CLK CLK CLK \
 N_CLK_c_937_n N_CLK_c_1003_n N_CLK_c_938_n N_CLK_M1_noxref_g \
 N_CLK_M8_noxref_g N_CLK_M15_noxref_g N_CLK_M16_noxref_g N_CLK_M29_noxref_g \
 N_CLK_M30_noxref_g N_CLK_c_1083_p N_CLK_c_1085_p N_CLK_c_1117_p \
 N_CLK_c_1124_p N_CLK_c_989_n N_CLK_c_990_n N_CLK_c_991_n N_CLK_c_992_n \
 N_CLK_c_995_n N_CLK_c_1012_n N_CLK_c_1015_n N_CLK_c_1017_n N_CLK_c_1053_p \
 N_CLK_c_1102_p N_CLK_c_1070_p N_CLK_c_1020_n N_CLK_c_1021_n N_CLK_c_996_n \
 N_CLK_c_1022_n N_CLK_c_1077_p N_CLK_c_1024_n )  PM_DFFQX1\%CLK
x_PM_DFFQX1\%noxref_6 ( N_noxref_6_c_1215_n N_noxref_6_c_1216_n \
 N_noxref_6_c_1142_n N_noxref_6_c_1223_n N_noxref_6_c_1169_n \
 N_noxref_6_c_1173_n N_noxref_6_c_1175_n N_noxref_6_c_1179_n \
 N_noxref_6_c_1144_n N_noxref_6_c_1229_n N_noxref_6_c_1183_n \
 N_noxref_6_c_1145_n N_noxref_6_c_1146_n N_noxref_6_c_1277_n \
 N_noxref_6_c_1241_n N_noxref_6_M3_noxref_g N_noxref_6_M9_noxref_g \
 N_noxref_6_M19_noxref_g N_noxref_6_M20_noxref_g N_noxref_6_M31_noxref_g \
 N_noxref_6_M32_noxref_g N_noxref_6_c_1147_n N_noxref_6_c_1149_n \
 N_noxref_6_c_1150_n N_noxref_6_c_1151_n N_noxref_6_c_1152_n \
 N_noxref_6_c_1153_n N_noxref_6_c_1154_n N_noxref_6_c_1156_n \
 N_noxref_6_c_1157_n N_noxref_6_c_1159_n N_noxref_6_c_1160_n \
 N_noxref_6_c_1161_n N_noxref_6_c_1162_n N_noxref_6_c_1163_n \
 N_noxref_6_c_1164_n N_noxref_6_c_1166_n N_noxref_6_c_1198_n \
 N_noxref_6_c_1199_n N_noxref_6_M2_noxref_d N_noxref_6_M13_noxref_d \
 N_noxref_6_M15_noxref_d N_noxref_6_M17_noxref_d )  PM_DFFQX1\%noxref_6
x_PM_DFFQX1\%noxref_7 ( N_noxref_7_c_1395_n N_noxref_7_c_1399_n \
 N_noxref_7_c_1416_n N_noxref_7_c_1420_n N_noxref_7_c_1422_n \
 N_noxref_7_c_1400_n N_noxref_7_c_1486_p N_noxref_7_c_1401_n \
 N_noxref_7_c_1402_n N_noxref_7_c_1509_p N_noxref_7_M11_noxref_g \
 N_noxref_7_M35_noxref_g N_noxref_7_M36_noxref_g N_noxref_7_c_1403_n \
 N_noxref_7_c_1405_n N_noxref_7_c_1406_n N_noxref_7_c_1407_n \
 N_noxref_7_c_1408_n N_noxref_7_c_1409_n N_noxref_7_c_1410_n \
 N_noxref_7_c_1412_n N_noxref_7_c_1435_n N_noxref_7_M10_noxref_d \
 N_noxref_7_M31_noxref_d N_noxref_7_M33_noxref_d )  PM_DFFQX1\%noxref_7
x_PM_DFFQX1\%noxref_8 ( N_noxref_8_c_1542_n N_noxref_8_c_1543_n \
 N_noxref_8_c_1572_n N_noxref_8_c_1642_n N_noxref_8_c_1544_n \
 N_noxref_8_c_1586_n N_noxref_8_c_1545_n N_noxref_8_c_1644_n \
 N_noxref_8_c_1546_n N_noxref_8_c_1594_n N_noxref_8_c_1598_n \
 N_noxref_8_c_1600_n N_noxref_8_c_1548_n N_noxref_8_c_1782_n \
 N_noxref_8_c_1549_n N_noxref_8_c_1797_n N_noxref_8_c_1550_n \
 N_noxref_8_c_1737_n N_noxref_8_M0_noxref_g N_noxref_8_M6_noxref_g \
 N_noxref_8_M12_noxref_g N_noxref_8_M13_noxref_g N_noxref_8_M14_noxref_g \
 N_noxref_8_M25_noxref_g N_noxref_8_M26_noxref_g N_noxref_8_M37_noxref_g \
 N_noxref_8_M38_noxref_g N_noxref_8_c_1552_n N_noxref_8_c_1554_n \
 N_noxref_8_c_1555_n N_noxref_8_c_1556_n N_noxref_8_c_1557_n \
 N_noxref_8_c_1558_n N_noxref_8_c_1559_n N_noxref_8_c_1561_n \
 N_noxref_8_c_1751_n N_noxref_8_c_1622_n N_noxref_8_c_1653_n \
 N_noxref_8_c_1656_n N_noxref_8_c_1658_n N_noxref_8_c_1690_n \
 N_noxref_8_c_1692_n N_noxref_8_c_1693_n N_noxref_8_c_1661_n \
 N_noxref_8_c_1662_n N_noxref_8_c_1806_n N_noxref_8_c_1809_n \
 N_noxref_8_c_1811_n N_noxref_8_c_1822_p N_noxref_8_c_1849_p \
 N_noxref_8_c_1841_p N_noxref_8_c_1814_n N_noxref_8_c_1815_n \
 N_noxref_8_c_1663_n N_noxref_8_c_1699_n N_noxref_8_c_1665_n \
 N_noxref_8_c_1816_n N_noxref_8_c_1830_p N_noxref_8_c_1818_n \
 N_noxref_8_M8_noxref_d N_noxref_8_M27_noxref_d N_noxref_8_M29_noxref_d )  \
 PM_DFFQX1\%noxref_8
x_PM_DFFQX1\%Q ( N_Q_c_1900_n N_Q_c_1901_n Q Q Q Q Q Q Q Q N_Q_c_1941_n \
 N_Q_c_1903_n N_Q_c_1915_n N_Q_c_1919_n N_Q_c_1921_n N_Q_c_1905_n N_Q_c_2048_p \
 N_Q_c_2024_n N_Q_M10_noxref_g N_Q_M33_noxref_g N_Q_M34_noxref_g N_Q_c_1949_n \
 N_Q_c_1952_n N_Q_c_1954_n N_Q_c_1987_n N_Q_c_1989_n N_Q_c_1990_n N_Q_c_1957_n \
 N_Q_c_1958_n N_Q_c_1959_n N_Q_c_1996_n N_Q_c_1961_n N_Q_M12_noxref_d \
 N_Q_M35_noxref_d N_Q_M37_noxref_d )  PM_DFFQX1\%Q
x_PM_DFFQX1\%noxref_10 ( N_noxref_10_c_2083_n N_noxref_10_c_2058_n \
 N_noxref_10_c_2062_n N_noxref_10_c_2065_n N_noxref_10_c_2076_n \
 N_noxref_10_M0_noxref_s )  PM_DFFQX1\%noxref_10
x_PM_DFFQX1\%noxref_11 ( N_noxref_11_c_2105_n N_noxref_11_c_2107_n \
 N_noxref_11_c_2110_n N_noxref_11_c_2113_n N_noxref_11_c_2124_n \
 N_noxref_11_M1_noxref_d N_noxref_11_M2_noxref_s )  PM_DFFQX1\%noxref_11
x_PM_DFFQX1\%D ( D D D N_D_c_2167_n N_D_c_2158_n N_D_M4_noxref_g \
 N_D_M21_noxref_g N_D_M22_noxref_g N_D_c_2177_n N_D_c_2178_n N_D_c_2179_n \
 N_D_c_2180_n N_D_c_2182_n N_D_c_2183_n N_D_c_2185_n N_D_c_2186_n N_D_c_2188_n \
 N_D_c_2189_n N_D_c_2191_n )  PM_DFFQX1\%D
x_PM_DFFQX1\%noxref_13 ( N_noxref_13_c_2250_n N_noxref_13_c_2231_n \
 N_noxref_13_c_2235_n N_noxref_13_c_2238_n N_noxref_13_c_2239_n \
 N_noxref_13_c_2242_n N_noxref_13_M3_noxref_s )  PM_DFFQX1\%noxref_13
x_PM_DFFQX1\%noxref_14 ( N_noxref_14_c_2302_n N_noxref_14_c_2283_n \
 N_noxref_14_c_2287_n N_noxref_14_c_2290_n N_noxref_14_c_2291_n \
 N_noxref_14_c_2294_n N_noxref_14_M5_noxref_s )  PM_DFFQX1\%noxref_14
x_PM_DFFQX1\%noxref_15 ( N_noxref_15_c_2355_n N_noxref_15_c_2336_n \
 N_noxref_15_c_2340_n N_noxref_15_c_2343_n N_noxref_15_c_2344_n \
 N_noxref_15_c_2347_n N_noxref_15_M7_noxref_s )  PM_DFFQX1\%noxref_15
x_PM_DFFQX1\%noxref_16 ( N_noxref_16_c_2408_n N_noxref_16_c_2389_n \
 N_noxref_16_c_2393_n N_noxref_16_c_2396_n N_noxref_16_c_2397_n \
 N_noxref_16_c_2400_n N_noxref_16_M9_noxref_s )  PM_DFFQX1\%noxref_16
x_PM_DFFQX1\%noxref_17 ( N_noxref_17_c_2460_n N_noxref_17_c_2443_n \
 N_noxref_17_c_2447_n N_noxref_17_c_2450_n N_noxref_17_c_2451_n \
 N_noxref_17_c_2453_n N_noxref_17_M11_noxref_s )  PM_DFFQX1\%noxref_17
cc_1 ( N_GND_c_1_p N_VDD_c_264_n ) capacitor c=0.00989031f //x=0.74 //y=0 \
 //x2=0.74 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_265_n ) capacitor c=0.00989031f //x=21.09 //y=0 \
 //x2=21.09 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_266_n ) capacitor c=0.00500587f //x=4.81 //y=0 \
 //x2=4.81 //y2=7.4
cc_4 ( N_GND_c_4_p N_VDD_c_267_n ) capacitor c=0.00500587f //x=8.14 //y=0 \
 //x2=8.14 //y2=7.4
cc_5 ( N_GND_c_5_p N_VDD_c_268_n ) capacitor c=0.00500587f //x=11.47 //y=0 \
 //x2=11.47 //y2=7.4
cc_6 ( N_GND_c_6_p N_VDD_c_269_n ) capacitor c=0.00524516f //x=14.8 //y=0 \
 //x2=14.8 //y2=7.4
cc_7 ( N_GND_c_7_p N_VDD_c_270_n ) capacitor c=0.00500587f //x=18.13 //y=0 \
 //x2=18.13 //y2=7.4
cc_8 ( N_GND_c_8_p N_noxref_3_c_555_n ) capacitor c=0.0264756f //x=21.09 //y=0 \
 //x2=7.285 //y2=3.33
cc_9 ( N_GND_c_9_p N_noxref_3_c_555_n ) capacitor c=0.00174514f //x=4.64 //y=0 \
 //x2=7.285 //y2=3.33
cc_10 ( N_GND_c_10_p N_noxref_3_c_555_n ) capacitor c=0.00192599f //x=5.905 \
 //y=0 //x2=7.285 //y2=3.33
cc_11 ( N_GND_c_11_p N_noxref_3_c_555_n ) capacitor c=5.39691e-19 //x=7.97 \
 //y=0 //x2=7.285 //y2=3.33
cc_12 ( N_GND_c_3_p N_noxref_3_c_555_n ) capacitor c=0.00820844f //x=4.81 \
 //y=0 //x2=7.285 //y2=3.33
cc_13 ( N_GND_c_8_p N_noxref_3_c_560_n ) capacitor c=0.00172266f //x=21.09 \
 //y=0 //x2=3.445 //y2=3.33
cc_14 ( N_GND_c_8_p N_noxref_3_c_561_n ) capacitor c=0.0143714f //x=21.09 \
 //y=0 //x2=9.135 //y2=3.33
cc_15 ( N_GND_c_11_p N_noxref_3_c_561_n ) capacitor c=0.00157139f //x=7.97 \
 //y=0 //x2=9.135 //y2=3.33
cc_16 ( N_GND_c_16_p N_noxref_3_c_561_n ) capacitor c=0.00189853f //x=9.235 \
 //y=0 //x2=9.135 //y2=3.33
cc_17 ( N_GND_c_4_p N_noxref_3_c_561_n ) capacitor c=0.00820844f //x=8.14 \
 //y=0 //x2=9.135 //y2=3.33
cc_18 ( N_GND_c_8_p N_noxref_3_c_565_n ) capacitor c=0.00153258f //x=21.09 \
 //y=0 //x2=7.515 //y2=3.33
cc_19 ( N_GND_c_3_p N_noxref_3_c_566_n ) capacitor c=9.53263e-19 //x=4.81 \
 //y=0 //x2=3.33 //y2=2.08
cc_20 ( N_GND_c_4_p N_noxref_3_c_567_n ) capacitor c=0.0462817f //x=8.14 //y=0 \
 //x2=7.315 //y2=1.655
cc_21 ( N_GND_c_3_p N_noxref_3_c_568_n ) capacitor c=9.64732e-19 //x=4.81 \
 //y=0 //x2=7.4 //y2=3.33
cc_22 ( N_GND_c_4_p N_noxref_3_c_569_n ) capacitor c=0.0179404f //x=8.14 //y=0 \
 //x2=9.25 //y2=2.08
cc_23 ( N_GND_c_16_p N_noxref_3_c_570_n ) capacitor c=0.00135046f //x=9.235 \
 //y=0 //x2=9.055 //y2=0.865
cc_24 ( N_GND_M5_noxref_d N_noxref_3_c_570_n ) capacitor c=0.00220047f \
 //x=9.13 //y=0.865 //x2=9.055 //y2=0.865
cc_25 ( N_GND_M5_noxref_d N_noxref_3_c_572_n ) capacitor c=0.00255985f \
 //x=9.13 //y=0.865 //x2=9.055 //y2=1.21
cc_26 ( N_GND_c_4_p N_noxref_3_c_573_n ) capacitor c=0.0018059f //x=8.14 //y=0 \
 //x2=9.055 //y2=1.52
cc_27 ( N_GND_c_4_p N_noxref_3_c_574_n ) capacitor c=0.0114883f //x=8.14 //y=0 \
 //x2=9.055 //y2=1.915
cc_28 ( N_GND_M5_noxref_d N_noxref_3_c_575_n ) capacitor c=0.0131326f //x=9.13 \
 //y=0.865 //x2=9.43 //y2=0.71
cc_29 ( N_GND_M5_noxref_d N_noxref_3_c_576_n ) capacitor c=0.00193127f \
 //x=9.13 //y=0.865 //x2=9.43 //y2=1.365
cc_30 ( N_GND_c_30_p N_noxref_3_c_577_n ) capacitor c=0.00130622f //x=11.3 \
 //y=0 //x2=9.585 //y2=0.865
cc_31 ( N_GND_M5_noxref_d N_noxref_3_c_577_n ) capacitor c=0.00257848f \
 //x=9.13 //y=0.865 //x2=9.585 //y2=0.865
cc_32 ( N_GND_M5_noxref_d N_noxref_3_c_579_n ) capacitor c=0.00255985f \
 //x=9.13 //y=0.865 //x2=9.585 //y2=1.21
cc_33 ( N_GND_c_3_p N_noxref_3_M4_noxref_d ) capacitor c=8.58106e-19 //x=4.81 \
 //y=0 //x2=6.77 //y2=0.905
cc_34 ( N_GND_c_4_p N_noxref_3_M4_noxref_d ) capacitor c=0.00616547f //x=8.14 \
 //y=0 //x2=6.77 //y2=0.905
cc_35 ( N_GND_M3_noxref_d N_noxref_3_M4_noxref_d ) capacitor c=0.00143464f \
 //x=5.8 //y=0.865 //x2=6.77 //y2=0.905
cc_36 ( N_GND_c_8_p N_noxref_4_c_787_n ) capacitor c=0.0143714f //x=21.09 \
 //y=0 //x2=12.465 //y2=3.33
cc_37 ( N_GND_c_30_p N_noxref_4_c_787_n ) capacitor c=0.00157139f //x=11.3 \
 //y=0 //x2=12.465 //y2=3.33
cc_38 ( N_GND_c_38_p N_noxref_4_c_787_n ) capacitor c=0.00189853f //x=12.565 \
 //y=0 //x2=12.465 //y2=3.33
cc_39 ( N_GND_c_5_p N_noxref_4_c_787_n ) capacitor c=0.00820844f //x=11.47 \
 //y=0 //x2=12.465 //y2=3.33
cc_40 ( N_GND_c_8_p N_noxref_4_c_791_n ) capacitor c=0.00174211f //x=21.09 \
 //y=0 //x2=10.845 //y2=3.33
cc_41 ( N_GND_c_5_p N_noxref_4_c_792_n ) capacitor c=0.0462817f //x=11.47 \
 //y=0 //x2=10.645 //y2=1.655
cc_42 ( N_GND_c_4_p N_noxref_4_c_793_n ) capacitor c=9.64732e-19 //x=8.14 \
 //y=0 //x2=10.73 //y2=3.33
cc_43 ( N_GND_c_5_p N_noxref_4_c_794_n ) capacitor c=0.0179404f //x=11.47 \
 //y=0 //x2=12.58 //y2=2.08
cc_44 ( N_GND_c_38_p N_noxref_4_c_795_n ) capacitor c=0.00135046f //x=12.565 \
 //y=0 //x2=12.385 //y2=0.865
cc_45 ( N_GND_M7_noxref_d N_noxref_4_c_795_n ) capacitor c=0.00220047f \
 //x=12.46 //y=0.865 //x2=12.385 //y2=0.865
cc_46 ( N_GND_M7_noxref_d N_noxref_4_c_797_n ) capacitor c=0.00255985f \
 //x=12.46 //y=0.865 //x2=12.385 //y2=1.21
cc_47 ( N_GND_c_5_p N_noxref_4_c_798_n ) capacitor c=0.0018059f //x=11.47 \
 //y=0 //x2=12.385 //y2=1.52
cc_48 ( N_GND_c_5_p N_noxref_4_c_799_n ) capacitor c=0.0114883f //x=11.47 \
 //y=0 //x2=12.385 //y2=1.915
cc_49 ( N_GND_M7_noxref_d N_noxref_4_c_800_n ) capacitor c=0.0131326f \
 //x=12.46 //y=0.865 //x2=12.76 //y2=0.71
cc_50 ( N_GND_M7_noxref_d N_noxref_4_c_801_n ) capacitor c=0.00193127f \
 //x=12.46 //y=0.865 //x2=12.76 //y2=1.365
cc_51 ( N_GND_c_51_p N_noxref_4_c_802_n ) capacitor c=0.00130622f //x=14.63 \
 //y=0 //x2=12.915 //y2=0.865
cc_52 ( N_GND_M7_noxref_d N_noxref_4_c_802_n ) capacitor c=0.00257848f \
 //x=12.46 //y=0.865 //x2=12.915 //y2=0.865
cc_53 ( N_GND_M7_noxref_d N_noxref_4_c_804_n ) capacitor c=0.00255985f \
 //x=12.46 //y=0.865 //x2=12.915 //y2=1.21
cc_54 ( N_GND_c_4_p N_noxref_4_M6_noxref_d ) capacitor c=8.58106e-19 //x=8.14 \
 //y=0 //x2=10.1 //y2=0.905
cc_55 ( N_GND_c_5_p N_noxref_4_M6_noxref_d ) capacitor c=0.00616547f //x=11.47 \
 //y=0 //x2=10.1 //y2=0.905
cc_56 ( N_GND_M5_noxref_d N_noxref_4_M6_noxref_d ) capacitor c=0.00143464f \
 //x=9.13 //y=0.865 //x2=10.1 //y2=0.905
cc_57 ( N_GND_c_1_p N_CLK_c_937_n ) capacitor c=7.64246e-19 //x=0.74 //y=0 \
 //x2=2.22 //y2=2.08
cc_58 ( N_GND_c_5_p N_CLK_c_938_n ) capacitor c=9.2064e-19 //x=11.47 //y=0 \
 //x2=13.32 //y2=2.08
cc_59 ( N_GND_c_6_p N_CLK_c_938_n ) capacitor c=9.53263e-19 //x=14.8 //y=0 \
 //x2=13.32 //y2=2.08
cc_60 ( N_GND_c_8_p N_noxref_6_c_1142_n ) capacitor c=0.046817f //x=21.09 \
 //y=0 //x2=15.795 //y2=3.7
cc_61 ( N_GND_c_6_p N_noxref_6_c_1142_n ) capacitor c=0.00533016f //x=14.8 \
 //y=0 //x2=15.795 //y2=3.7
cc_62 ( N_GND_c_3_p N_noxref_6_c_1144_n ) capacitor c=0.0459932f //x=4.81 \
 //y=0 //x2=3.985 //y2=1.665
cc_63 ( N_GND_c_3_p N_noxref_6_c_1145_n ) capacitor c=0.0179404f //x=4.81 \
 //y=0 //x2=5.92 //y2=2.08
cc_64 ( N_GND_c_6_p N_noxref_6_c_1146_n ) capacitor c=0.0179404f //x=14.8 \
 //y=0 //x2=15.91 //y2=2.08
cc_65 ( N_GND_c_10_p N_noxref_6_c_1147_n ) capacitor c=0.00135046f //x=5.905 \
 //y=0 //x2=5.725 //y2=0.865
cc_66 ( N_GND_M3_noxref_d N_noxref_6_c_1147_n ) capacitor c=0.00220047f \
 //x=5.8 //y=0.865 //x2=5.725 //y2=0.865
cc_67 ( N_GND_M3_noxref_d N_noxref_6_c_1149_n ) capacitor c=0.00255985f \
 //x=5.8 //y=0.865 //x2=5.725 //y2=1.21
cc_68 ( N_GND_c_3_p N_noxref_6_c_1150_n ) capacitor c=0.00189421f //x=4.81 \
 //y=0 //x2=5.725 //y2=1.52
cc_69 ( N_GND_c_3_p N_noxref_6_c_1151_n ) capacitor c=0.0114883f //x=4.81 \
 //y=0 //x2=5.725 //y2=1.915
cc_70 ( N_GND_M3_noxref_d N_noxref_6_c_1152_n ) capacitor c=0.0131326f //x=5.8 \
 //y=0.865 //x2=6.1 //y2=0.71
cc_71 ( N_GND_M3_noxref_d N_noxref_6_c_1153_n ) capacitor c=0.00193127f \
 //x=5.8 //y=0.865 //x2=6.1 //y2=1.365
cc_72 ( N_GND_c_11_p N_noxref_6_c_1154_n ) capacitor c=0.00130622f //x=7.97 \
 //y=0 //x2=6.255 //y2=0.865
cc_73 ( N_GND_M3_noxref_d N_noxref_6_c_1154_n ) capacitor c=0.00257848f \
 //x=5.8 //y=0.865 //x2=6.255 //y2=0.865
cc_74 ( N_GND_M3_noxref_d N_noxref_6_c_1156_n ) capacitor c=0.00255985f \
 //x=5.8 //y=0.865 //x2=6.255 //y2=1.21
cc_75 ( N_GND_c_75_p N_noxref_6_c_1157_n ) capacitor c=0.00135046f //x=15.895 \
 //y=0 //x2=15.715 //y2=0.865
cc_76 ( N_GND_M9_noxref_d N_noxref_6_c_1157_n ) capacitor c=0.00220047f \
 //x=15.79 //y=0.865 //x2=15.715 //y2=0.865
cc_77 ( N_GND_M9_noxref_d N_noxref_6_c_1159_n ) capacitor c=0.00255985f \
 //x=15.79 //y=0.865 //x2=15.715 //y2=1.21
cc_78 ( N_GND_c_6_p N_noxref_6_c_1160_n ) capacitor c=0.0018059f //x=14.8 \
 //y=0 //x2=15.715 //y2=1.52
cc_79 ( N_GND_c_6_p N_noxref_6_c_1161_n ) capacitor c=0.0114883f //x=14.8 \
 //y=0 //x2=15.715 //y2=1.915
cc_80 ( N_GND_M9_noxref_d N_noxref_6_c_1162_n ) capacitor c=0.0131326f \
 //x=15.79 //y=0.865 //x2=16.09 //y2=0.71
cc_81 ( N_GND_M9_noxref_d N_noxref_6_c_1163_n ) capacitor c=0.00193127f \
 //x=15.79 //y=0.865 //x2=16.09 //y2=1.365
cc_82 ( N_GND_c_82_p N_noxref_6_c_1164_n ) capacitor c=0.00130622f //x=17.96 \
 //y=0 //x2=16.245 //y2=0.865
cc_83 ( N_GND_M9_noxref_d N_noxref_6_c_1164_n ) capacitor c=0.00257848f \
 //x=15.79 //y=0.865 //x2=16.245 //y2=0.865
cc_84 ( N_GND_M9_noxref_d N_noxref_6_c_1166_n ) capacitor c=0.00255985f \
 //x=15.79 //y=0.865 //x2=16.245 //y2=1.21
cc_85 ( N_GND_c_3_p N_noxref_6_M2_noxref_d ) capacitor c=0.00591582f //x=4.81 \
 //y=0 //x2=3.395 //y2=0.915
cc_86 ( N_GND_c_8_p N_noxref_7_c_1395_n ) capacitor c=0.0143714f //x=21.09 \
 //y=0 //x2=19.125 //y2=3.33
cc_87 ( N_GND_c_82_p N_noxref_7_c_1395_n ) capacitor c=0.00157139f //x=17.96 \
 //y=0 //x2=19.125 //y2=3.33
cc_88 ( N_GND_c_88_p N_noxref_7_c_1395_n ) capacitor c=0.00189853f //x=19.225 \
 //y=0 //x2=19.125 //y2=3.33
cc_89 ( N_GND_c_7_p N_noxref_7_c_1395_n ) capacitor c=0.00820844f //x=18.13 \
 //y=0 //x2=19.125 //y2=3.33
cc_90 ( N_GND_c_8_p N_noxref_7_c_1399_n ) capacitor c=0.00174211f //x=21.09 \
 //y=0 //x2=17.505 //y2=3.33
cc_91 ( N_GND_c_7_p N_noxref_7_c_1400_n ) capacitor c=0.0462817f //x=18.13 \
 //y=0 //x2=17.305 //y2=1.655
cc_92 ( N_GND_c_6_p N_noxref_7_c_1401_n ) capacitor c=9.64732e-19 //x=14.8 \
 //y=0 //x2=17.39 //y2=3.33
cc_93 ( N_GND_c_7_p N_noxref_7_c_1402_n ) capacitor c=0.0179404f //x=18.13 \
 //y=0 //x2=19.24 //y2=2.08
cc_94 ( N_GND_c_88_p N_noxref_7_c_1403_n ) capacitor c=0.00135046f //x=19.225 \
 //y=0 //x2=19.045 //y2=0.865
cc_95 ( N_GND_M11_noxref_d N_noxref_7_c_1403_n ) capacitor c=0.00220047f \
 //x=19.12 //y=0.865 //x2=19.045 //y2=0.865
cc_96 ( N_GND_M11_noxref_d N_noxref_7_c_1405_n ) capacitor c=0.00255985f \
 //x=19.12 //y=0.865 //x2=19.045 //y2=1.21
cc_97 ( N_GND_c_7_p N_noxref_7_c_1406_n ) capacitor c=0.0018059f //x=18.13 \
 //y=0 //x2=19.045 //y2=1.52
cc_98 ( N_GND_c_7_p N_noxref_7_c_1407_n ) capacitor c=0.0114883f //x=18.13 \
 //y=0 //x2=19.045 //y2=1.915
cc_99 ( N_GND_M11_noxref_d N_noxref_7_c_1408_n ) capacitor c=0.0131326f \
 //x=19.12 //y=0.865 //x2=19.42 //y2=0.71
cc_100 ( N_GND_M11_noxref_d N_noxref_7_c_1409_n ) capacitor c=0.00193127f \
 //x=19.12 //y=0.865 //x2=19.42 //y2=1.365
cc_101 ( N_GND_c_2_p N_noxref_7_c_1410_n ) capacitor c=0.00130622f //x=21.09 \
 //y=0 //x2=19.575 //y2=0.865
cc_102 ( N_GND_M11_noxref_d N_noxref_7_c_1410_n ) capacitor c=0.00257848f \
 //x=19.12 //y=0.865 //x2=19.575 //y2=0.865
cc_103 ( N_GND_M11_noxref_d N_noxref_7_c_1412_n ) capacitor c=0.00255985f \
 //x=19.12 //y=0.865 //x2=19.575 //y2=1.21
cc_104 ( N_GND_c_6_p N_noxref_7_M10_noxref_d ) capacitor c=8.58106e-19 \
 //x=14.8 //y=0 //x2=16.76 //y2=0.905
cc_105 ( N_GND_c_7_p N_noxref_7_M10_noxref_d ) capacitor c=0.00616547f \
 //x=18.13 //y=0 //x2=16.76 //y2=0.905
cc_106 ( N_GND_M9_noxref_d N_noxref_7_M10_noxref_d ) capacitor c=0.00143464f \
 //x=15.79 //y=0.865 //x2=16.76 //y2=0.905
cc_107 ( N_GND_c_8_p N_noxref_8_c_1542_n ) capacitor c=0.0147496f //x=21.09 \
 //y=0 //x2=9.875 //y2=4.07
cc_108 ( N_GND_c_8_p N_noxref_8_c_1543_n ) capacitor c=0.0015877f //x=21.09 \
 //y=0 //x2=1.225 //y2=4.07
cc_109 ( N_GND_c_8_p N_noxref_8_c_1544_n ) capacitor c=0.0131174f //x=21.09 \
 //y=0 //x2=19.865 //y2=4.07
cc_110 ( N_GND_c_1_p N_noxref_8_c_1545_n ) capacitor c=0.0180363f //x=0.74 \
 //y=0 //x2=1.11 //y2=2.08
cc_111 ( N_GND_c_4_p N_noxref_8_c_1546_n ) capacitor c=9.2064e-19 //x=8.14 \
 //y=0 //x2=9.99 //y2=2.08
cc_112 ( N_GND_c_5_p N_noxref_8_c_1546_n ) capacitor c=9.53263e-19 //x=11.47 \
 //y=0 //x2=9.99 //y2=2.08
cc_113 ( N_GND_c_6_p N_noxref_8_c_1548_n ) capacitor c=0.0462817f //x=14.8 \
 //y=0 //x2=13.975 //y2=1.655
cc_114 ( N_GND_c_5_p N_noxref_8_c_1549_n ) capacitor c=9.64732e-19 //x=11.47 \
 //y=0 //x2=14.06 //y2=4.07
cc_115 ( N_GND_c_2_p N_noxref_8_c_1550_n ) capacitor c=9.53263e-19 //x=21.09 \
 //y=0 //x2=19.98 //y2=2.08
cc_116 ( N_GND_c_7_p N_noxref_8_c_1550_n ) capacitor c=9.2064e-19 //x=18.13 \
 //y=0 //x2=19.98 //y2=2.08
cc_117 ( N_GND_c_117_p N_noxref_8_c_1552_n ) capacitor c=0.00132755f //x=0.99 \
 //y=0 //x2=0.81 //y2=0.875
cc_118 ( N_GND_M0_noxref_d N_noxref_8_c_1552_n ) capacitor c=0.00211996f \
 //x=0.885 //y=0.875 //x2=0.81 //y2=0.875
cc_119 ( N_GND_M0_noxref_d N_noxref_8_c_1554_n ) capacitor c=0.00255985f \
 //x=0.885 //y=0.875 //x2=0.81 //y2=1.22
cc_120 ( N_GND_c_1_p N_noxref_8_c_1555_n ) capacitor c=0.00295461f //x=0.74 \
 //y=0 //x2=0.81 //y2=1.53
cc_121 ( N_GND_c_1_p N_noxref_8_c_1556_n ) capacitor c=0.0134214f //x=0.74 \
 //y=0 //x2=0.81 //y2=1.915
cc_122 ( N_GND_M0_noxref_d N_noxref_8_c_1557_n ) capacitor c=0.0131341f \
 //x=0.885 //y=0.875 //x2=1.185 //y2=0.72
cc_123 ( N_GND_M0_noxref_d N_noxref_8_c_1558_n ) capacitor c=0.00193146f \
 //x=0.885 //y=0.875 //x2=1.185 //y2=1.375
cc_124 ( N_GND_c_9_p N_noxref_8_c_1559_n ) capacitor c=0.00129018f //x=4.64 \
 //y=0 //x2=1.34 //y2=0.875
cc_125 ( N_GND_M0_noxref_d N_noxref_8_c_1559_n ) capacitor c=0.00257848f \
 //x=0.885 //y=0.875 //x2=1.34 //y2=0.875
cc_126 ( N_GND_M0_noxref_d N_noxref_8_c_1561_n ) capacitor c=0.00255985f \
 //x=0.885 //y=0.875 //x2=1.34 //y2=1.22
cc_127 ( N_GND_c_5_p N_noxref_8_M8_noxref_d ) capacitor c=8.58106e-19 \
 //x=11.47 //y=0 //x2=13.43 //y2=0.905
cc_128 ( N_GND_c_6_p N_noxref_8_M8_noxref_d ) capacitor c=0.00616547f //x=14.8 \
 //y=0 //x2=13.43 //y2=0.905
cc_129 ( N_GND_M7_noxref_d N_noxref_8_M8_noxref_d ) capacitor c=0.00143464f \
 //x=12.46 //y=0.865 //x2=13.43 //y2=0.905
cc_130 ( N_GND_c_8_p N_Q_c_1900_n ) capacitor c=0.0187193f //x=21.09 //y=0 \
 //x2=20.605 //y2=3.7
cc_131 ( N_GND_c_8_p N_Q_c_1901_n ) capacitor c=0.00157091f //x=21.09 //y=0 \
 //x2=16.765 //y2=3.7
cc_132 ( N_GND_c_7_p Q ) capacitor c=9.64732e-19 //x=18.13 //y=0 //x2=20.72 \
 //y2=2.22
cc_133 ( N_GND_c_6_p N_Q_c_1903_n ) capacitor c=9.2064e-19 //x=14.8 //y=0 \
 //x2=16.65 //y2=2.08
cc_134 ( N_GND_c_7_p N_Q_c_1903_n ) capacitor c=9.53263e-19 //x=18.13 //y=0 \
 //x2=16.65 //y2=2.08
cc_135 ( N_GND_c_2_p N_Q_c_1905_n ) capacitor c=0.0468439f //x=21.09 //y=0 \
 //x2=20.635 //y2=1.655
cc_136 ( N_GND_c_2_p N_Q_M12_noxref_d ) capacitor c=0.00618259f //x=21.09 \
 //y=0 //x2=20.09 //y2=0.905
cc_137 ( N_GND_c_7_p N_Q_M12_noxref_d ) capacitor c=8.58106e-19 //x=18.13 \
 //y=0 //x2=20.09 //y2=0.905
cc_138 ( N_GND_M11_noxref_d N_Q_M12_noxref_d ) capacitor c=0.00143464f \
 //x=19.12 //y=0.865 //x2=20.09 //y2=0.905
cc_139 ( N_GND_c_8_p N_noxref_10_c_2058_n ) capacitor c=0.00618812f //x=21.09 \
 //y=0 //x2=1.475 //y2=1.59
cc_140 ( N_GND_c_117_p N_noxref_10_c_2058_n ) capacitor c=0.00110021f //x=0.99 \
 //y=0 //x2=1.475 //y2=1.59
cc_141 ( N_GND_c_9_p N_noxref_10_c_2058_n ) capacitor c=0.00179185f //x=4.64 \
 //y=0 //x2=1.475 //y2=1.59
cc_142 ( N_GND_M0_noxref_d N_noxref_10_c_2058_n ) capacitor c=0.00894788f \
 //x=0.885 //y=0.875 //x2=1.475 //y2=1.59
cc_143 ( N_GND_c_8_p N_noxref_10_c_2062_n ) capacitor c=0.00575184f //x=21.09 \
 //y=0 //x2=1.56 //y2=0.625
cc_144 ( N_GND_c_9_p N_noxref_10_c_2062_n ) capacitor c=0.0140218f //x=4.64 \
 //y=0 //x2=1.56 //y2=0.625
cc_145 ( N_GND_M0_noxref_d N_noxref_10_c_2062_n ) capacitor c=0.033954f \
 //x=0.885 //y=0.875 //x2=1.56 //y2=0.625
cc_146 ( N_GND_c_8_p N_noxref_10_c_2065_n ) capacitor c=0.0139021f //x=21.09 \
 //y=0 //x2=2.445 //y2=0.54
cc_147 ( N_GND_c_9_p N_noxref_10_c_2065_n ) capacitor c=0.0356078f //x=4.64 \
 //y=0 //x2=2.445 //y2=0.54
cc_148 ( N_GND_c_2_p N_noxref_10_c_2065_n ) capacitor c=0.00177725f //x=21.09 \
 //y=0 //x2=2.445 //y2=0.54
cc_149 ( N_GND_c_8_p N_noxref_10_M0_noxref_s ) capacitor c=0.0125336f \
 //x=21.09 //y=0 //x2=0.455 //y2=0.375
cc_150 ( N_GND_c_117_p N_noxref_10_M0_noxref_s ) capacitor c=0.0140218f \
 //x=0.99 //y=0 //x2=0.455 //y2=0.375
cc_151 ( N_GND_c_1_p N_noxref_10_M0_noxref_s ) capacitor c=0.0712607f //x=0.74 \
 //y=0 //x2=0.455 //y2=0.375
cc_152 ( N_GND_c_9_p N_noxref_10_M0_noxref_s ) capacitor c=0.0131422f //x=4.64 \
 //y=0 //x2=0.455 //y2=0.375
cc_153 ( N_GND_c_3_p N_noxref_10_M0_noxref_s ) capacitor c=3.31601e-19 \
 //x=4.81 //y=0 //x2=0.455 //y2=0.375
cc_154 ( N_GND_M0_noxref_d N_noxref_10_M0_noxref_s ) capacitor c=0.033718f \
 //x=0.885 //y=0.875 //x2=0.455 //y2=0.375
cc_155 ( N_GND_c_8_p N_noxref_11_c_2105_n ) capacitor c=0.00402784f //x=21.09 \
 //y=0 //x2=3.015 //y2=0.995
cc_156 ( N_GND_c_9_p N_noxref_11_c_2105_n ) capacitor c=0.00829979f //x=4.64 \
 //y=0 //x2=3.015 //y2=0.995
cc_157 ( N_GND_c_8_p N_noxref_11_c_2107_n ) capacitor c=0.00575184f //x=21.09 \
 //y=0 //x2=3.1 //y2=0.625
cc_158 ( N_GND_c_9_p N_noxref_11_c_2107_n ) capacitor c=0.0140218f //x=4.64 \
 //y=0 //x2=3.1 //y2=0.625
cc_159 ( N_GND_M0_noxref_d N_noxref_11_c_2107_n ) capacitor c=6.21394e-19 \
 //x=0.885 //y=0.875 //x2=3.1 //y2=0.625
cc_160 ( N_GND_c_8_p N_noxref_11_c_2110_n ) capacitor c=0.0118365f //x=21.09 \
 //y=0 //x2=3.985 //y2=0.54
cc_161 ( N_GND_c_9_p N_noxref_11_c_2110_n ) capacitor c=0.0365413f //x=4.64 \
 //y=0 //x2=3.985 //y2=0.54
cc_162 ( N_GND_c_2_p N_noxref_11_c_2110_n ) capacitor c=0.00189848f //x=21.09 \
 //y=0 //x2=3.985 //y2=0.54
cc_163 ( N_GND_c_8_p N_noxref_11_c_2113_n ) capacitor c=0.00287549f //x=21.09 \
 //y=0 //x2=4.07 //y2=0.625
cc_164 ( N_GND_c_9_p N_noxref_11_c_2113_n ) capacitor c=0.0142658f //x=4.64 \
 //y=0 //x2=4.07 //y2=0.625
cc_165 ( N_GND_c_3_p N_noxref_11_c_2113_n ) capacitor c=0.0404137f //x=4.81 \
 //y=0 //x2=4.07 //y2=0.625
cc_166 ( N_GND_M0_noxref_d N_noxref_11_M1_noxref_d ) capacitor c=0.00162435f \
 //x=0.885 //y=0.875 //x2=1.86 //y2=0.91
cc_167 ( N_GND_c_1_p N_noxref_11_M2_noxref_s ) capacitor c=8.16352e-19 \
 //x=0.74 //y=0 //x2=2.965 //y2=0.375
cc_168 ( N_GND_c_3_p N_noxref_11_M2_noxref_s ) capacitor c=0.00183576f \
 //x=4.81 //y=0 //x2=2.965 //y2=0.375
cc_169 ( N_GND_c_3_p N_D_c_2158_n ) capacitor c=9.2064e-19 //x=4.81 //y=0 \
 //x2=6.66 //y2=2.08
cc_170 ( N_GND_c_4_p N_D_c_2158_n ) capacitor c=9.53263e-19 //x=8.14 //y=0 \
 //x2=6.66 //y2=2.08
cc_171 ( N_GND_c_8_p N_noxref_13_c_2231_n ) capacitor c=0.00552526f //x=21.09 \
 //y=0 //x2=6.39 //y2=1.58
cc_172 ( N_GND_c_10_p N_noxref_13_c_2231_n ) capacitor c=0.00113001f //x=5.905 \
 //y=0 //x2=6.39 //y2=1.58
cc_173 ( N_GND_c_11_p N_noxref_13_c_2231_n ) capacitor c=0.0018242f //x=7.97 \
 //y=0 //x2=6.39 //y2=1.58
cc_174 ( N_GND_M3_noxref_d N_noxref_13_c_2231_n ) capacitor c=0.00897209f \
 //x=5.8 //y=0.865 //x2=6.39 //y2=1.58
cc_175 ( N_GND_c_8_p N_noxref_13_c_2235_n ) capacitor c=0.00293348f //x=21.09 \
 //y=0 //x2=6.475 //y2=0.615
cc_176 ( N_GND_c_11_p N_noxref_13_c_2235_n ) capacitor c=0.0149357f //x=7.97 \
 //y=0 //x2=6.475 //y2=0.615
cc_177 ( N_GND_M3_noxref_d N_noxref_13_c_2235_n ) capacitor c=0.033812f \
 //x=5.8 //y=0.865 //x2=6.475 //y2=0.615
cc_178 ( N_GND_c_3_p N_noxref_13_c_2238_n ) capacitor c=2.91423e-19 //x=4.81 \
 //y=0 //x2=6.475 //y2=1.495
cc_179 ( N_GND_c_8_p N_noxref_13_c_2239_n ) capacitor c=0.0120397f //x=21.09 \
 //y=0 //x2=7.36 //y2=0.53
cc_180 ( N_GND_c_11_p N_noxref_13_c_2239_n ) capacitor c=0.037553f //x=7.97 \
 //y=0 //x2=7.36 //y2=0.53
cc_181 ( N_GND_c_2_p N_noxref_13_c_2239_n ) capacitor c=0.00198885f //x=21.09 \
 //y=0 //x2=7.36 //y2=0.53
cc_182 ( N_GND_c_8_p N_noxref_13_c_2242_n ) capacitor c=0.00292576f //x=21.09 \
 //y=0 //x2=7.445 //y2=0.615
cc_183 ( N_GND_c_11_p N_noxref_13_c_2242_n ) capacitor c=0.0148673f //x=7.97 \
 //y=0 //x2=7.445 //y2=0.615
cc_184 ( N_GND_c_4_p N_noxref_13_c_2242_n ) capacitor c=0.0431718f //x=8.14 \
 //y=0 //x2=7.445 //y2=0.615
cc_185 ( N_GND_c_8_p N_noxref_13_M3_noxref_s ) capacitor c=0.00293348f \
 //x=21.09 //y=0 //x2=5.37 //y2=0.365
cc_186 ( N_GND_c_10_p N_noxref_13_M3_noxref_s ) capacitor c=0.0149357f \
 //x=5.905 //y=0 //x2=5.37 //y2=0.365
cc_187 ( N_GND_c_3_p N_noxref_13_M3_noxref_s ) capacitor c=0.0583534f //x=4.81 \
 //y=0 //x2=5.37 //y2=0.365
cc_188 ( N_GND_c_4_p N_noxref_13_M3_noxref_s ) capacitor c=0.00198043f \
 //x=8.14 //y=0 //x2=5.37 //y2=0.365
cc_189 ( N_GND_M3_noxref_d N_noxref_13_M3_noxref_s ) capacitor c=0.0334197f \
 //x=5.8 //y=0.865 //x2=5.37 //y2=0.365
cc_190 ( N_GND_c_8_p N_noxref_14_c_2283_n ) capacitor c=0.00556119f //x=21.09 \
 //y=0 //x2=9.72 //y2=1.58
cc_191 ( N_GND_c_16_p N_noxref_14_c_2283_n ) capacitor c=0.00113001f //x=9.235 \
 //y=0 //x2=9.72 //y2=1.58
cc_192 ( N_GND_c_30_p N_noxref_14_c_2283_n ) capacitor c=0.00180846f //x=11.3 \
 //y=0 //x2=9.72 //y2=1.58
cc_193 ( N_GND_M5_noxref_d N_noxref_14_c_2283_n ) capacitor c=0.00897268f \
 //x=9.13 //y=0.865 //x2=9.72 //y2=1.58
cc_194 ( N_GND_c_8_p N_noxref_14_c_2287_n ) capacitor c=0.00302994f //x=21.09 \
 //y=0 //x2=9.805 //y2=0.615
cc_195 ( N_GND_c_30_p N_noxref_14_c_2287_n ) capacitor c=0.0146208f //x=11.3 \
 //y=0 //x2=9.805 //y2=0.615
cc_196 ( N_GND_M5_noxref_d N_noxref_14_c_2287_n ) capacitor c=0.033812f \
 //x=9.13 //y=0.865 //x2=9.805 //y2=0.615
cc_197 ( N_GND_c_4_p N_noxref_14_c_2290_n ) capacitor c=2.91423e-19 //x=8.14 \
 //y=0 //x2=9.805 //y2=1.495
cc_198 ( N_GND_c_8_p N_noxref_14_c_2291_n ) capacitor c=0.0123695f //x=21.09 \
 //y=0 //x2=10.69 //y2=0.53
cc_199 ( N_GND_c_30_p N_noxref_14_c_2291_n ) capacitor c=0.0373121f //x=11.3 \
 //y=0 //x2=10.69 //y2=0.53
cc_200 ( N_GND_c_2_p N_noxref_14_c_2291_n ) capacitor c=0.00198885f //x=21.09 \
 //y=0 //x2=10.69 //y2=0.53
cc_201 ( N_GND_c_8_p N_noxref_14_c_2294_n ) capacitor c=0.00292576f //x=21.09 \
 //y=0 //x2=10.775 //y2=0.615
cc_202 ( N_GND_c_30_p N_noxref_14_c_2294_n ) capacitor c=0.0148673f //x=11.3 \
 //y=0 //x2=10.775 //y2=0.615
cc_203 ( N_GND_c_5_p N_noxref_14_c_2294_n ) capacitor c=0.0431718f //x=11.47 \
 //y=0 //x2=10.775 //y2=0.615
cc_204 ( N_GND_c_8_p N_noxref_14_M5_noxref_s ) capacitor c=0.00293348f \
 //x=21.09 //y=0 //x2=8.7 //y2=0.365
cc_205 ( N_GND_c_16_p N_noxref_14_M5_noxref_s ) capacitor c=0.0149357f \
 //x=9.235 //y=0 //x2=8.7 //y2=0.365
cc_206 ( N_GND_c_4_p N_noxref_14_M5_noxref_s ) capacitor c=0.058339f //x=8.14 \
 //y=0 //x2=8.7 //y2=0.365
cc_207 ( N_GND_c_5_p N_noxref_14_M5_noxref_s ) capacitor c=0.00198043f \
 //x=11.47 //y=0 //x2=8.7 //y2=0.365
cc_208 ( N_GND_M5_noxref_d N_noxref_14_M5_noxref_s ) capacitor c=0.0334197f \
 //x=9.13 //y=0.865 //x2=8.7 //y2=0.365
cc_209 ( N_GND_c_8_p N_noxref_15_c_2336_n ) capacitor c=0.00556119f //x=21.09 \
 //y=0 //x2=13.05 //y2=1.58
cc_210 ( N_GND_c_38_p N_noxref_15_c_2336_n ) capacitor c=0.00113001f \
 //x=12.565 //y=0 //x2=13.05 //y2=1.58
cc_211 ( N_GND_c_51_p N_noxref_15_c_2336_n ) capacitor c=0.00180846f //x=14.63 \
 //y=0 //x2=13.05 //y2=1.58
cc_212 ( N_GND_M7_noxref_d N_noxref_15_c_2336_n ) capacitor c=0.00897268f \
 //x=12.46 //y=0.865 //x2=13.05 //y2=1.58
cc_213 ( N_GND_c_8_p N_noxref_15_c_2340_n ) capacitor c=0.00302994f //x=21.09 \
 //y=0 //x2=13.135 //y2=0.615
cc_214 ( N_GND_c_51_p N_noxref_15_c_2340_n ) capacitor c=0.0146208f //x=14.63 \
 //y=0 //x2=13.135 //y2=0.615
cc_215 ( N_GND_M7_noxref_d N_noxref_15_c_2340_n ) capacitor c=0.033812f \
 //x=12.46 //y=0.865 //x2=13.135 //y2=0.615
cc_216 ( N_GND_c_5_p N_noxref_15_c_2343_n ) capacitor c=2.91423e-19 //x=11.47 \
 //y=0 //x2=13.135 //y2=1.495
cc_217 ( N_GND_c_8_p N_noxref_15_c_2344_n ) capacitor c=0.0124224f //x=21.09 \
 //y=0 //x2=14.02 //y2=0.53
cc_218 ( N_GND_c_51_p N_noxref_15_c_2344_n ) capacitor c=0.0371035f //x=14.63 \
 //y=0 //x2=14.02 //y2=0.53
cc_219 ( N_GND_c_2_p N_noxref_15_c_2344_n ) capacitor c=0.00198885f //x=21.09 \
 //y=0 //x2=14.02 //y2=0.53
cc_220 ( N_GND_c_8_p N_noxref_15_c_2347_n ) capacitor c=0.00303012f //x=21.09 \
 //y=0 //x2=14.105 //y2=0.615
cc_221 ( N_GND_c_51_p N_noxref_15_c_2347_n ) capacitor c=0.0144264f //x=14.63 \
 //y=0 //x2=14.105 //y2=0.615
cc_222 ( N_GND_c_6_p N_noxref_15_c_2347_n ) capacitor c=0.0431718f //x=14.8 \
 //y=0 //x2=14.105 //y2=0.615
cc_223 ( N_GND_c_8_p N_noxref_15_M7_noxref_s ) capacitor c=0.00293348f \
 //x=21.09 //y=0 //x2=12.03 //y2=0.365
cc_224 ( N_GND_c_38_p N_noxref_15_M7_noxref_s ) capacitor c=0.0149357f \
 //x=12.565 //y=0 //x2=12.03 //y2=0.365
cc_225 ( N_GND_c_5_p N_noxref_15_M7_noxref_s ) capacitor c=0.058339f //x=11.47 \
 //y=0 //x2=12.03 //y2=0.365
cc_226 ( N_GND_c_6_p N_noxref_15_M7_noxref_s ) capacitor c=0.00198043f \
 //x=14.8 //y=0 //x2=12.03 //y2=0.365
cc_227 ( N_GND_M7_noxref_d N_noxref_15_M7_noxref_s ) capacitor c=0.0334197f \
 //x=12.46 //y=0.865 //x2=12.03 //y2=0.365
cc_228 ( N_GND_c_8_p N_noxref_16_c_2389_n ) capacitor c=0.00565424f //x=21.09 \
 //y=0 //x2=16.38 //y2=1.58
cc_229 ( N_GND_c_75_p N_noxref_16_c_2389_n ) capacitor c=0.00111428f \
 //x=15.895 //y=0 //x2=16.38 //y2=1.58
cc_230 ( N_GND_c_82_p N_noxref_16_c_2389_n ) capacitor c=0.00180846f //x=17.96 \
 //y=0 //x2=16.38 //y2=1.58
cc_231 ( N_GND_M9_noxref_d N_noxref_16_c_2389_n ) capacitor c=0.00901798f \
 //x=15.79 //y=0.865 //x2=16.38 //y2=1.58
cc_232 ( N_GND_c_8_p N_noxref_16_c_2393_n ) capacitor c=0.0050999f //x=21.09 \
 //y=0 //x2=16.465 //y2=0.615
cc_233 ( N_GND_c_82_p N_noxref_16_c_2393_n ) capacitor c=0.0146208f //x=17.96 \
 //y=0 //x2=16.465 //y2=0.615
cc_234 ( N_GND_M9_noxref_d N_noxref_16_c_2393_n ) capacitor c=0.033812f \
 //x=15.79 //y=0.865 //x2=16.465 //y2=0.615
cc_235 ( N_GND_c_6_p N_noxref_16_c_2396_n ) capacitor c=2.91423e-19 //x=14.8 \
 //y=0 //x2=16.465 //y2=1.495
cc_236 ( N_GND_c_8_p N_noxref_16_c_2397_n ) capacitor c=0.0123615f //x=21.09 \
 //y=0 //x2=17.35 //y2=0.53
cc_237 ( N_GND_c_82_p N_noxref_16_c_2397_n ) capacitor c=0.0373121f //x=17.96 \
 //y=0 //x2=17.35 //y2=0.53
cc_238 ( N_GND_c_2_p N_noxref_16_c_2397_n ) capacitor c=0.00198885f //x=21.09 \
 //y=0 //x2=17.35 //y2=0.53
cc_239 ( N_GND_c_8_p N_noxref_16_c_2400_n ) capacitor c=0.00292576f //x=21.09 \
 //y=0 //x2=17.435 //y2=0.615
cc_240 ( N_GND_c_82_p N_noxref_16_c_2400_n ) capacitor c=0.0148673f //x=17.96 \
 //y=0 //x2=17.435 //y2=0.615
cc_241 ( N_GND_c_7_p N_noxref_16_c_2400_n ) capacitor c=0.0431718f //x=18.13 \
 //y=0 //x2=17.435 //y2=0.615
cc_242 ( N_GND_c_8_p N_noxref_16_M9_noxref_s ) capacitor c=0.00302994f \
 //x=21.09 //y=0 //x2=15.36 //y2=0.365
cc_243 ( N_GND_c_75_p N_noxref_16_M9_noxref_s ) capacitor c=0.0146208f \
 //x=15.895 //y=0 //x2=15.36 //y2=0.365
cc_244 ( N_GND_c_6_p N_noxref_16_M9_noxref_s ) capacitor c=0.058339f //x=14.8 \
 //y=0 //x2=15.36 //y2=0.365
cc_245 ( N_GND_c_7_p N_noxref_16_M9_noxref_s ) capacitor c=0.00198043f \
 //x=18.13 //y=0 //x2=15.36 //y2=0.365
cc_246 ( N_GND_M9_noxref_d N_noxref_16_M9_noxref_s ) capacitor c=0.0334197f \
 //x=15.79 //y=0.865 //x2=15.36 //y2=0.365
cc_247 ( N_GND_c_8_p N_noxref_17_c_2443_n ) capacitor c=0.00556119f //x=21.09 \
 //y=0 //x2=19.71 //y2=1.58
cc_248 ( N_GND_c_88_p N_noxref_17_c_2443_n ) capacitor c=0.00113001f \
 //x=19.225 //y=0 //x2=19.71 //y2=1.58
cc_249 ( N_GND_c_2_p N_noxref_17_c_2443_n ) capacitor c=0.00180846f //x=21.09 \
 //y=0 //x2=19.71 //y2=1.58
cc_250 ( N_GND_M11_noxref_d N_noxref_17_c_2443_n ) capacitor c=0.00897268f \
 //x=19.12 //y=0.865 //x2=19.71 //y2=1.58
cc_251 ( N_GND_c_8_p N_noxref_17_c_2447_n ) capacitor c=0.00302994f //x=21.09 \
 //y=0 //x2=19.795 //y2=0.615
cc_252 ( N_GND_c_2_p N_noxref_17_c_2447_n ) capacitor c=0.0146208f //x=21.09 \
 //y=0 //x2=19.795 //y2=0.615
cc_253 ( N_GND_M11_noxref_d N_noxref_17_c_2447_n ) capacitor c=0.033812f \
 //x=19.12 //y=0.865 //x2=19.795 //y2=0.615
cc_254 ( N_GND_c_7_p N_noxref_17_c_2450_n ) capacitor c=2.91423e-19 //x=18.13 \
 //y=0 //x2=19.795 //y2=1.495
cc_255 ( N_GND_c_8_p N_noxref_17_c_2451_n ) capacitor c=0.0124196f //x=21.09 \
 //y=0 //x2=20.68 //y2=0.53
cc_256 ( N_GND_c_2_p N_noxref_17_c_2451_n ) capacitor c=0.0390924f //x=21.09 \
 //y=0 //x2=20.68 //y2=0.53
cc_257 ( N_GND_c_8_p N_noxref_17_c_2453_n ) capacitor c=0.00302319f //x=21.09 \
 //y=0 //x2=20.765 //y2=0.615
cc_258 ( N_GND_c_2_p N_noxref_17_c_2453_n ) capacitor c=0.0584079f //x=21.09 \
 //y=0 //x2=20.765 //y2=0.615
cc_259 ( N_GND_c_8_p N_noxref_17_M11_noxref_s ) capacitor c=0.00293348f \
 //x=21.09 //y=0 //x2=18.69 //y2=0.365
cc_260 ( N_GND_c_88_p N_noxref_17_M11_noxref_s ) capacitor c=0.0149357f \
 //x=19.225 //y=0 //x2=18.69 //y2=0.365
cc_261 ( N_GND_c_2_p N_noxref_17_M11_noxref_s ) capacitor c=0.00198482f \
 //x=21.09 //y=0 //x2=18.69 //y2=0.365
cc_262 ( N_GND_c_7_p N_noxref_17_M11_noxref_s ) capacitor c=0.058339f \
 //x=18.13 //y=0 //x2=18.69 //y2=0.365
cc_263 ( N_GND_M11_noxref_d N_noxref_17_M11_noxref_s ) capacitor c=0.0334197f \
 //x=19.12 //y=0.865 //x2=18.69 //y2=0.365
cc_264 ( N_VDD_c_266_n N_noxref_3_c_566_n ) capacitor c=6.58823e-19 //x=4.81 \
 //y=7.4 //x2=3.33 //y2=2.08
cc_265 ( N_VDD_c_272_p N_noxref_3_c_584_n ) capacitor c=0.00453663f //x=21.09 \
 //y=7.4 //x2=6.835 //y2=5.2
cc_266 ( N_VDD_c_273_p N_noxref_3_c_584_n ) capacitor c=4.48391e-19 //x=6.395 \
 //y=7.4 //x2=6.835 //y2=5.2
cc_267 ( N_VDD_c_274_p N_noxref_3_c_584_n ) capacitor c=4.48391e-19 //x=7.275 \
 //y=7.4 //x2=6.835 //y2=5.2
cc_268 ( N_VDD_M20_noxref_d N_noxref_3_c_584_n ) capacitor c=0.0124542f \
 //x=6.335 //y=5.02 //x2=6.835 //y2=5.2
cc_269 ( N_VDD_c_266_n N_noxref_3_c_588_n ) capacitor c=0.00985474f //x=4.81 \
 //y=7.4 //x2=6.125 //y2=5.2
cc_270 ( N_VDD_M19_noxref_s N_noxref_3_c_588_n ) capacitor c=0.087833f \
 //x=5.465 //y=5.02 //x2=6.125 //y2=5.2
cc_271 ( N_VDD_c_272_p N_noxref_3_c_590_n ) capacitor c=0.00301575f //x=21.09 \
 //y=7.4 //x2=7.315 //y2=5.2
cc_272 ( N_VDD_c_274_p N_noxref_3_c_590_n ) capacitor c=7.72068e-19 //x=7.275 \
 //y=7.4 //x2=7.315 //y2=5.2
cc_273 ( N_VDD_M22_noxref_d N_noxref_3_c_590_n ) capacitor c=0.0158515f \
 //x=7.215 //y=5.02 //x2=7.315 //y2=5.2
cc_274 ( N_VDD_M23_noxref_s N_noxref_3_c_590_n ) capacitor c=2.44532e-19 \
 //x=8.795 //y=5.02 //x2=7.315 //y2=5.2
cc_275 ( N_VDD_c_266_n N_noxref_3_c_568_n ) capacitor c=0.00151618f //x=4.81 \
 //y=7.4 //x2=7.4 //y2=3.33
cc_276 ( N_VDD_c_267_n N_noxref_3_c_568_n ) capacitor c=0.0429414f //x=8.14 \
 //y=7.4 //x2=7.4 //y2=3.33
cc_277 ( N_VDD_c_272_p N_noxref_3_c_569_n ) capacitor c=0.00125279f //x=21.09 \
 //y=7.4 //x2=9.25 //y2=2.08
cc_278 ( N_VDD_c_285_p N_noxref_3_c_569_n ) capacitor c=2.87256e-19 //x=9.725 \
 //y=7.4 //x2=9.25 //y2=2.08
cc_279 ( N_VDD_c_267_n N_noxref_3_c_569_n ) capacitor c=0.0134208f //x=8.14 \
 //y=7.4 //x2=9.25 //y2=2.08
cc_280 ( N_VDD_c_287_p N_noxref_3_M17_noxref_g ) capacitor c=0.00675175f \
 //x=3.645 //y=7.4 //x2=3.07 //y2=6.02
cc_281 ( N_VDD_M16_noxref_d N_noxref_3_M17_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=3.07 //y2=6.02
cc_282 ( N_VDD_c_287_p N_noxref_3_M18_noxref_g ) capacitor c=0.00675379f \
 //x=3.645 //y=7.4 //x2=3.51 //y2=6.02
cc_283 ( N_VDD_M18_noxref_d N_noxref_3_M18_noxref_g ) capacitor c=0.0394719f \
 //x=3.585 //y=5.02 //x2=3.51 //y2=6.02
cc_284 ( N_VDD_c_285_p N_noxref_3_M23_noxref_g ) capacitor c=0.00726866f \
 //x=9.725 //y=7.4 //x2=9.15 //y2=6.02
cc_285 ( N_VDD_M23_noxref_s N_noxref_3_M23_noxref_g ) capacitor c=0.054195f \
 //x=8.795 //y=5.02 //x2=9.15 //y2=6.02
cc_286 ( N_VDD_c_285_p N_noxref_3_M24_noxref_g ) capacitor c=0.00672952f \
 //x=9.725 //y=7.4 //x2=9.59 //y2=6.02
cc_287 ( N_VDD_M24_noxref_d N_noxref_3_M24_noxref_g ) capacitor c=0.015318f \
 //x=9.665 //y=5.02 //x2=9.59 //y2=6.02
cc_288 ( N_VDD_c_267_n N_noxref_3_c_607_n ) capacitor c=0.0150435f //x=8.14 \
 //y=7.4 //x2=9.25 //y2=4.7
cc_289 ( N_VDD_c_272_p N_noxref_3_M19_noxref_d ) capacitor c=0.00275225f \
 //x=21.09 //y=7.4 //x2=5.895 //y2=5.02
cc_290 ( N_VDD_c_273_p N_noxref_3_M19_noxref_d ) capacitor c=0.0140317f \
 //x=6.395 //y=7.4 //x2=5.895 //y2=5.02
cc_291 ( N_VDD_c_267_n N_noxref_3_M19_noxref_d ) capacitor c=6.94454e-19 \
 //x=8.14 //y=7.4 //x2=5.895 //y2=5.02
cc_292 ( N_VDD_M20_noxref_d N_noxref_3_M19_noxref_d ) capacitor c=0.0664752f \
 //x=6.335 //y=5.02 //x2=5.895 //y2=5.02
cc_293 ( N_VDD_c_272_p N_noxref_3_M21_noxref_d ) capacitor c=0.00275225f \
 //x=21.09 //y=7.4 //x2=6.775 //y2=5.02
cc_294 ( N_VDD_c_274_p N_noxref_3_M21_noxref_d ) capacitor c=0.0140317f \
 //x=7.275 //y=7.4 //x2=6.775 //y2=5.02
cc_295 ( N_VDD_c_267_n N_noxref_3_M21_noxref_d ) capacitor c=0.0120541f \
 //x=8.14 //y=7.4 //x2=6.775 //y2=5.02
cc_296 ( N_VDD_M19_noxref_s N_noxref_3_M21_noxref_d ) capacitor c=0.00111971f \
 //x=5.465 //y=5.02 //x2=6.775 //y2=5.02
cc_297 ( N_VDD_M20_noxref_d N_noxref_3_M21_noxref_d ) capacitor c=0.0664752f \
 //x=6.335 //y=5.02 //x2=6.775 //y2=5.02
cc_298 ( N_VDD_M22_noxref_d N_noxref_3_M21_noxref_d ) capacitor c=0.0664752f \
 //x=7.215 //y=5.02 //x2=6.775 //y2=5.02
cc_299 ( N_VDD_M23_noxref_s N_noxref_3_M21_noxref_d ) capacitor c=4.54516e-19 \
 //x=8.795 //y=5.02 //x2=6.775 //y2=5.02
cc_300 ( N_VDD_c_272_p N_noxref_4_c_808_n ) capacitor c=0.00453663f //x=21.09 \
 //y=7.4 //x2=10.165 //y2=5.2
cc_301 ( N_VDD_c_285_p N_noxref_4_c_808_n ) capacitor c=4.48391e-19 //x=9.725 \
 //y=7.4 //x2=10.165 //y2=5.2
cc_302 ( N_VDD_c_309_p N_noxref_4_c_808_n ) capacitor c=4.48391e-19 //x=10.605 \
 //y=7.4 //x2=10.165 //y2=5.2
cc_303 ( N_VDD_M24_noxref_d N_noxref_4_c_808_n ) capacitor c=0.0124542f \
 //x=9.665 //y=5.02 //x2=10.165 //y2=5.2
cc_304 ( N_VDD_c_267_n N_noxref_4_c_812_n ) capacitor c=0.00985474f //x=8.14 \
 //y=7.4 //x2=9.455 //y2=5.2
cc_305 ( N_VDD_M23_noxref_s N_noxref_4_c_812_n ) capacitor c=0.087833f \
 //x=8.795 //y=5.02 //x2=9.455 //y2=5.2
cc_306 ( N_VDD_c_272_p N_noxref_4_c_814_n ) capacitor c=0.00301575f //x=21.09 \
 //y=7.4 //x2=10.645 //y2=5.2
cc_307 ( N_VDD_c_309_p N_noxref_4_c_814_n ) capacitor c=7.72068e-19 //x=10.605 \
 //y=7.4 //x2=10.645 //y2=5.2
cc_308 ( N_VDD_M26_noxref_d N_noxref_4_c_814_n ) capacitor c=0.0158515f \
 //x=10.545 //y=5.02 //x2=10.645 //y2=5.2
cc_309 ( N_VDD_M27_noxref_s N_noxref_4_c_814_n ) capacitor c=2.44532e-19 \
 //x=12.125 //y=5.02 //x2=10.645 //y2=5.2
cc_310 ( N_VDD_c_267_n N_noxref_4_c_793_n ) capacitor c=0.00151618f //x=8.14 \
 //y=7.4 //x2=10.73 //y2=3.33
cc_311 ( N_VDD_c_268_n N_noxref_4_c_793_n ) capacitor c=0.0427674f //x=11.47 \
 //y=7.4 //x2=10.73 //y2=3.33
cc_312 ( N_VDD_c_272_p N_noxref_4_c_794_n ) capacitor c=0.00125279f //x=21.09 \
 //y=7.4 //x2=12.58 //y2=2.08
cc_313 ( N_VDD_c_320_p N_noxref_4_c_794_n ) capacitor c=2.87256e-19 //x=13.055 \
 //y=7.4 //x2=12.58 //y2=2.08
cc_314 ( N_VDD_c_268_n N_noxref_4_c_794_n ) capacitor c=0.0133228f //x=11.47 \
 //y=7.4 //x2=12.58 //y2=2.08
cc_315 ( N_VDD_c_320_p N_noxref_4_M27_noxref_g ) capacitor c=0.00726866f \
 //x=13.055 //y=7.4 //x2=12.48 //y2=6.02
cc_316 ( N_VDD_M27_noxref_s N_noxref_4_M27_noxref_g ) capacitor c=0.054195f \
 //x=12.125 //y=5.02 //x2=12.48 //y2=6.02
cc_317 ( N_VDD_c_320_p N_noxref_4_M28_noxref_g ) capacitor c=0.00672952f \
 //x=13.055 //y=7.4 //x2=12.92 //y2=6.02
cc_318 ( N_VDD_M28_noxref_d N_noxref_4_M28_noxref_g ) capacitor c=0.015318f \
 //x=12.995 //y=5.02 //x2=12.92 //y2=6.02
cc_319 ( N_VDD_c_268_n N_noxref_4_c_827_n ) capacitor c=0.0149273f //x=11.47 \
 //y=7.4 //x2=12.58 //y2=4.7
cc_320 ( N_VDD_c_272_p N_noxref_4_M23_noxref_d ) capacitor c=0.00275225f \
 //x=21.09 //y=7.4 //x2=9.225 //y2=5.02
cc_321 ( N_VDD_c_285_p N_noxref_4_M23_noxref_d ) capacitor c=0.0140317f \
 //x=9.725 //y=7.4 //x2=9.225 //y2=5.02
cc_322 ( N_VDD_c_268_n N_noxref_4_M23_noxref_d ) capacitor c=6.94454e-19 \
 //x=11.47 //y=7.4 //x2=9.225 //y2=5.02
cc_323 ( N_VDD_M24_noxref_d N_noxref_4_M23_noxref_d ) capacitor c=0.0664752f \
 //x=9.665 //y=5.02 //x2=9.225 //y2=5.02
cc_324 ( N_VDD_c_272_p N_noxref_4_M25_noxref_d ) capacitor c=0.00275225f \
 //x=21.09 //y=7.4 //x2=10.105 //y2=5.02
cc_325 ( N_VDD_c_309_p N_noxref_4_M25_noxref_d ) capacitor c=0.0140317f \
 //x=10.605 //y=7.4 //x2=10.105 //y2=5.02
cc_326 ( N_VDD_c_268_n N_noxref_4_M25_noxref_d ) capacitor c=0.0120541f \
 //x=11.47 //y=7.4 //x2=10.105 //y2=5.02
cc_327 ( N_VDD_M23_noxref_s N_noxref_4_M25_noxref_d ) capacitor c=0.00111971f \
 //x=8.795 //y=5.02 //x2=10.105 //y2=5.02
cc_328 ( N_VDD_M24_noxref_d N_noxref_4_M25_noxref_d ) capacitor c=0.0664752f \
 //x=9.665 //y=5.02 //x2=10.105 //y2=5.02
cc_329 ( N_VDD_M26_noxref_d N_noxref_4_M25_noxref_d ) capacitor c=0.0664752f \
 //x=10.545 //y=5.02 //x2=10.105 //y2=5.02
cc_330 ( N_VDD_M27_noxref_s N_noxref_4_M25_noxref_d ) capacitor c=4.54516e-19 \
 //x=12.125 //y=5.02 //x2=10.105 //y2=5.02
cc_331 ( N_VDD_c_272_p N_CLK_c_940_n ) capacitor c=0.0824294f //x=21.09 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_332 ( N_VDD_c_339_p N_CLK_c_940_n ) capacitor c=0.00258496f //x=4.64 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_333 ( N_VDD_c_340_p N_CLK_c_940_n ) capacitor c=0.00209689f //x=5.515 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_334 ( N_VDD_c_273_p N_CLK_c_940_n ) capacitor c=7.81728e-19 //x=6.395 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_335 ( N_VDD_c_342_p N_CLK_c_940_n ) capacitor c=0.00205475f //x=7.97 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_336 ( N_VDD_c_343_p N_CLK_c_940_n ) capacitor c=0.00209689f //x=8.845 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_337 ( N_VDD_c_285_p N_CLK_c_940_n ) capacitor c=7.81728e-19 //x=9.725 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_338 ( N_VDD_c_345_p N_CLK_c_940_n ) capacitor c=0.00205475f //x=11.3 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_339 ( N_VDD_c_346_p N_CLK_c_940_n ) capacitor c=0.00209689f //x=12.175 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_340 ( N_VDD_c_320_p N_CLK_c_940_n ) capacitor c=7.81728e-19 //x=13.055 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_341 ( N_VDD_c_266_n N_CLK_c_940_n ) capacitor c=0.0389825f //x=4.81 //y=7.4 \
 //x2=13.205 //y2=4.44
cc_342 ( N_VDD_c_267_n N_CLK_c_940_n ) capacitor c=0.0389825f //x=8.14 //y=7.4 \
 //x2=13.205 //y2=4.44
cc_343 ( N_VDD_c_268_n N_CLK_c_940_n ) capacitor c=0.0389825f //x=11.47 \
 //y=7.4 //x2=13.205 //y2=4.44
cc_344 ( N_VDD_M19_noxref_s N_CLK_c_940_n ) capacitor c=0.00541054f //x=5.465 \
 //y=5.02 //x2=13.205 //y2=4.44
cc_345 ( N_VDD_M22_noxref_d N_CLK_c_940_n ) capacitor c=6.7165e-19 //x=7.215 \
 //y=5.02 //x2=13.205 //y2=4.44
cc_346 ( N_VDD_M23_noxref_s N_CLK_c_940_n ) capacitor c=0.00541054f //x=8.795 \
 //y=5.02 //x2=13.205 //y2=4.44
cc_347 ( N_VDD_M26_noxref_d N_CLK_c_940_n ) capacitor c=6.7165e-19 //x=10.545 \
 //y=5.02 //x2=13.205 //y2=4.44
cc_348 ( N_VDD_M27_noxref_s N_CLK_c_940_n ) capacitor c=0.00541054f //x=12.125 \
 //y=5.02 //x2=13.205 //y2=4.44
cc_349 ( N_VDD_c_272_p N_CLK_c_958_n ) capacitor c=0.00146064f //x=21.09 \
 //y=7.4 //x2=2.335 //y2=4.44
cc_350 ( N_VDD_c_272_p N_CLK_c_937_n ) capacitor c=2.03287e-19 //x=21.09 \
 //y=7.4 //x2=2.22 //y2=2.08
cc_351 ( N_VDD_c_264_n N_CLK_c_937_n ) capacitor c=9.53425e-19 //x=0.74 \
 //y=7.4 //x2=2.22 //y2=2.08
cc_352 ( N_VDD_c_268_n N_CLK_c_938_n ) capacitor c=5.27482e-19 //x=11.47 \
 //y=7.4 //x2=13.32 //y2=2.08
cc_353 ( N_VDD_c_269_n N_CLK_c_938_n ) capacitor c=7.54518e-19 //x=14.8 \
 //y=7.4 //x2=13.32 //y2=2.08
cc_354 ( N_VDD_c_361_p N_CLK_M15_noxref_g ) capacitor c=0.00676195f //x=2.765 \
 //y=7.4 //x2=2.19 //y2=6.02
cc_355 ( N_VDD_M14_noxref_d N_CLK_M15_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=2.19 //y2=6.02
cc_356 ( N_VDD_c_361_p N_CLK_M16_noxref_g ) capacitor c=0.00675175f //x=2.765 \
 //y=7.4 //x2=2.63 //y2=6.02
cc_357 ( N_VDD_M16_noxref_d N_CLK_M16_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=2.63 //y2=6.02
cc_358 ( N_VDD_c_365_p N_CLK_M29_noxref_g ) capacitor c=0.00673971f //x=13.935 \
 //y=7.4 //x2=13.36 //y2=6.02
cc_359 ( N_VDD_M28_noxref_d N_CLK_M29_noxref_g ) capacitor c=0.015318f \
 //x=12.995 //y=5.02 //x2=13.36 //y2=6.02
cc_360 ( N_VDD_c_365_p N_CLK_M30_noxref_g ) capacitor c=0.00672952f //x=13.935 \
 //y=7.4 //x2=13.8 //y2=6.02
cc_361 ( N_VDD_c_269_n N_CLK_M30_noxref_g ) capacitor c=0.00864163f //x=14.8 \
 //y=7.4 //x2=13.8 //y2=6.02
cc_362 ( N_VDD_M30_noxref_d N_CLK_M30_noxref_g ) capacitor c=0.0430452f \
 //x=13.875 //y=5.02 //x2=13.8 //y2=6.02
cc_363 ( N_VDD_c_269_n N_noxref_6_c_1142_n ) capacitor c=0.00290959f //x=14.8 \
 //y=7.4 //x2=15.795 //y2=3.7
cc_364 ( N_VDD_c_272_p N_noxref_6_c_1169_n ) capacitor c=0.00449316f //x=21.09 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_365 ( N_VDD_c_372_p N_noxref_6_c_1169_n ) capacitor c=4.32228e-19 //x=1.885 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_366 ( N_VDD_c_361_p N_noxref_6_c_1169_n ) capacitor c=4.31906e-19 //x=2.765 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_367 ( N_VDD_M14_noxref_d N_noxref_6_c_1169_n ) capacitor c=0.0115147f \
 //x=1.825 //y=5.02 //x2=2.325 //y2=5.155
cc_368 ( N_VDD_c_264_n N_noxref_6_c_1173_n ) capacitor c=0.00880189f //x=0.74 \
 //y=7.4 //x2=1.615 //y2=5.155
cc_369 ( N_VDD_M13_noxref_s N_noxref_6_c_1173_n ) capacitor c=0.0831083f \
 //x=0.955 //y=5.02 //x2=1.615 //y2=5.155
cc_370 ( N_VDD_c_272_p N_noxref_6_c_1175_n ) capacitor c=0.0044221f //x=21.09 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_371 ( N_VDD_c_361_p N_noxref_6_c_1175_n ) capacitor c=4.31931e-19 //x=2.765 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_372 ( N_VDD_c_287_p N_noxref_6_c_1175_n ) capacitor c=4.31931e-19 //x=3.645 \
 //y=7.4 //x2=3.205 //y2=5.155
cc_373 ( N_VDD_M16_noxref_d N_noxref_6_c_1175_n ) capacitor c=0.0112985f \
 //x=2.705 //y=5.02 //x2=3.205 //y2=5.155
cc_374 ( N_VDD_c_272_p N_noxref_6_c_1179_n ) capacitor c=0.00434174f //x=21.09 \
 //y=7.4 //x2=3.985 //y2=5.155
cc_375 ( N_VDD_c_287_p N_noxref_6_c_1179_n ) capacitor c=7.46626e-19 //x=3.645 \
 //y=7.4 //x2=3.985 //y2=5.155
cc_376 ( N_VDD_c_339_p N_noxref_6_c_1179_n ) capacitor c=0.00198565f //x=4.64 \
 //y=7.4 //x2=3.985 //y2=5.155
cc_377 ( N_VDD_M18_noxref_d N_noxref_6_c_1179_n ) capacitor c=0.0112985f \
 //x=3.585 //y=5.02 //x2=3.985 //y2=5.155
cc_378 ( N_VDD_c_266_n N_noxref_6_c_1183_n ) capacitor c=0.0426341f //x=4.81 \
 //y=7.4 //x2=4.07 //y2=3.7
cc_379 ( N_VDD_c_272_p N_noxref_6_c_1145_n ) capacitor c=0.00125279f //x=21.09 \
 //y=7.4 //x2=5.92 //y2=2.08
cc_380 ( N_VDD_c_273_p N_noxref_6_c_1145_n ) capacitor c=2.87256e-19 //x=6.395 \
 //y=7.4 //x2=5.92 //y2=2.08
cc_381 ( N_VDD_c_266_n N_noxref_6_c_1145_n ) capacitor c=0.0134665f //x=4.81 \
 //y=7.4 //x2=5.92 //y2=2.08
cc_382 ( N_VDD_c_272_p N_noxref_6_c_1146_n ) capacitor c=0.00126216f //x=21.09 \
 //y=7.4 //x2=15.91 //y2=2.08
cc_383 ( N_VDD_c_390_p N_noxref_6_c_1146_n ) capacitor c=2.87813e-19 \
 //x=16.385 //y=7.4 //x2=15.91 //y2=2.08
cc_384 ( N_VDD_c_269_n N_noxref_6_c_1146_n ) capacitor c=0.0157486f //x=14.8 \
 //y=7.4 //x2=15.91 //y2=2.08
cc_385 ( N_VDD_c_273_p N_noxref_6_M19_noxref_g ) capacitor c=0.00726866f \
 //x=6.395 //y=7.4 //x2=5.82 //y2=6.02
cc_386 ( N_VDD_M19_noxref_s N_noxref_6_M19_noxref_g ) capacitor c=0.054195f \
 //x=5.465 //y=5.02 //x2=5.82 //y2=6.02
cc_387 ( N_VDD_c_273_p N_noxref_6_M20_noxref_g ) capacitor c=0.00672952f \
 //x=6.395 //y=7.4 //x2=6.26 //y2=6.02
cc_388 ( N_VDD_M20_noxref_d N_noxref_6_M20_noxref_g ) capacitor c=0.015318f \
 //x=6.335 //y=5.02 //x2=6.26 //y2=6.02
cc_389 ( N_VDD_c_390_p N_noxref_6_M31_noxref_g ) capacitor c=0.00726866f \
 //x=16.385 //y=7.4 //x2=15.81 //y2=6.02
cc_390 ( N_VDD_M31_noxref_s N_noxref_6_M31_noxref_g ) capacitor c=0.054195f \
 //x=15.455 //y=5.02 //x2=15.81 //y2=6.02
cc_391 ( N_VDD_c_390_p N_noxref_6_M32_noxref_g ) capacitor c=0.00672952f \
 //x=16.385 //y=7.4 //x2=16.25 //y2=6.02
cc_392 ( N_VDD_M32_noxref_d N_noxref_6_M32_noxref_g ) capacitor c=0.015318f \
 //x=16.325 //y=5.02 //x2=16.25 //y2=6.02
cc_393 ( N_VDD_c_266_n N_noxref_6_c_1198_n ) capacitor c=0.015293f //x=4.81 \
 //y=7.4 //x2=5.92 //y2=4.7
cc_394 ( N_VDD_c_269_n N_noxref_6_c_1199_n ) capacitor c=0.0149273f //x=14.8 \
 //y=7.4 //x2=15.91 //y2=4.7
cc_395 ( N_VDD_c_272_p N_noxref_6_M13_noxref_d ) capacitor c=0.00285091f \
 //x=21.09 //y=7.4 //x2=1.385 //y2=5.02
cc_396 ( N_VDD_c_372_p N_noxref_6_M13_noxref_d ) capacitor c=0.0141016f \
 //x=1.885 //y=7.4 //x2=1.385 //y2=5.02
cc_397 ( N_VDD_M14_noxref_d N_noxref_6_M13_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=1.385 //y2=5.02
cc_398 ( N_VDD_c_272_p N_noxref_6_M15_noxref_d ) capacitor c=0.00275186f \
 //x=21.09 //y=7.4 //x2=2.265 //y2=5.02
cc_399 ( N_VDD_c_361_p N_noxref_6_M15_noxref_d ) capacitor c=0.0140346f \
 //x=2.765 //y=7.4 //x2=2.265 //y2=5.02
cc_400 ( N_VDD_c_266_n N_noxref_6_M15_noxref_d ) capacitor c=4.9285e-19 \
 //x=4.81 //y=7.4 //x2=2.265 //y2=5.02
cc_401 ( N_VDD_M13_noxref_s N_noxref_6_M15_noxref_d ) capacitor c=0.00130656f \
 //x=0.955 //y=5.02 //x2=2.265 //y2=5.02
cc_402 ( N_VDD_M14_noxref_d N_noxref_6_M15_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=2.265 //y2=5.02
cc_403 ( N_VDD_M16_noxref_d N_noxref_6_M15_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=2.265 //y2=5.02
cc_404 ( N_VDD_c_272_p N_noxref_6_M17_noxref_d ) capacitor c=0.00275235f \
 //x=21.09 //y=7.4 //x2=3.145 //y2=5.02
cc_405 ( N_VDD_c_287_p N_noxref_6_M17_noxref_d ) capacitor c=0.0137384f \
 //x=3.645 //y=7.4 //x2=3.145 //y2=5.02
cc_406 ( N_VDD_c_266_n N_noxref_6_M17_noxref_d ) capacitor c=0.00939849f \
 //x=4.81 //y=7.4 //x2=3.145 //y2=5.02
cc_407 ( N_VDD_M16_noxref_d N_noxref_6_M17_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=3.145 //y2=5.02
cc_408 ( N_VDD_M18_noxref_d N_noxref_6_M17_noxref_d ) capacitor c=0.0664752f \
 //x=3.585 //y=5.02 //x2=3.145 //y2=5.02
cc_409 ( N_VDD_M19_noxref_s N_noxref_6_M17_noxref_d ) capacitor c=4.52683e-19 \
 //x=5.465 //y=5.02 //x2=3.145 //y2=5.02
cc_410 ( N_VDD_c_272_p N_noxref_7_c_1416_n ) capacitor c=0.00460134f //x=21.09 \
 //y=7.4 //x2=16.825 //y2=5.2
cc_411 ( N_VDD_c_390_p N_noxref_7_c_1416_n ) capacitor c=4.48705e-19 \
 //x=16.385 //y=7.4 //x2=16.825 //y2=5.2
cc_412 ( N_VDD_c_419_p N_noxref_7_c_1416_n ) capacitor c=4.48705e-19 \
 //x=17.265 //y=7.4 //x2=16.825 //y2=5.2
cc_413 ( N_VDD_M32_noxref_d N_noxref_7_c_1416_n ) capacitor c=0.0126924f \
 //x=16.325 //y=5.02 //x2=16.825 //y2=5.2
cc_414 ( N_VDD_c_269_n N_noxref_7_c_1420_n ) capacitor c=0.00985474f //x=14.8 \
 //y=7.4 //x2=16.115 //y2=5.2
cc_415 ( N_VDD_M31_noxref_s N_noxref_7_c_1420_n ) capacitor c=0.087833f \
 //x=15.455 //y=5.02 //x2=16.115 //y2=5.2
cc_416 ( N_VDD_c_272_p N_noxref_7_c_1422_n ) capacitor c=0.00307195f //x=21.09 \
 //y=7.4 //x2=17.305 //y2=5.2
cc_417 ( N_VDD_c_419_p N_noxref_7_c_1422_n ) capacitor c=7.73167e-19 \
 //x=17.265 //y=7.4 //x2=17.305 //y2=5.2
cc_418 ( N_VDD_M34_noxref_d N_noxref_7_c_1422_n ) capacitor c=0.0161518f \
 //x=17.205 //y=5.02 //x2=17.305 //y2=5.2
cc_419 ( N_VDD_M35_noxref_s N_noxref_7_c_1422_n ) capacitor c=2.44532e-19 \
 //x=18.785 //y=5.02 //x2=17.305 //y2=5.2
cc_420 ( N_VDD_c_269_n N_noxref_7_c_1401_n ) capacitor c=0.00151618f //x=14.8 \
 //y=7.4 //x2=17.39 //y2=3.33
cc_421 ( N_VDD_c_270_n N_noxref_7_c_1401_n ) capacitor c=0.0455537f //x=18.13 \
 //y=7.4 //x2=17.39 //y2=3.33
cc_422 ( N_VDD_c_272_p N_noxref_7_c_1402_n ) capacitor c=0.00126216f //x=21.09 \
 //y=7.4 //x2=19.24 //y2=2.08
cc_423 ( N_VDD_c_430_p N_noxref_7_c_1402_n ) capacitor c=2.87813e-19 \
 //x=19.715 //y=7.4 //x2=19.24 //y2=2.08
cc_424 ( N_VDD_c_270_n N_noxref_7_c_1402_n ) capacitor c=0.0160121f //x=18.13 \
 //y=7.4 //x2=19.24 //y2=2.08
cc_425 ( N_VDD_c_430_p N_noxref_7_M35_noxref_g ) capacitor c=0.00726866f \
 //x=19.715 //y=7.4 //x2=19.14 //y2=6.02
cc_426 ( N_VDD_M35_noxref_s N_noxref_7_M35_noxref_g ) capacitor c=0.054195f \
 //x=18.785 //y=5.02 //x2=19.14 //y2=6.02
cc_427 ( N_VDD_c_430_p N_noxref_7_M36_noxref_g ) capacitor c=0.00672952f \
 //x=19.715 //y=7.4 //x2=19.58 //y2=6.02
cc_428 ( N_VDD_M36_noxref_d N_noxref_7_M36_noxref_g ) capacitor c=0.015318f \
 //x=19.655 //y=5.02 //x2=19.58 //y2=6.02
cc_429 ( N_VDD_c_270_n N_noxref_7_c_1435_n ) capacitor c=0.0150435f //x=18.13 \
 //y=7.4 //x2=19.24 //y2=4.7
cc_430 ( N_VDD_c_272_p N_noxref_7_M31_noxref_d ) capacitor c=0.00285083f \
 //x=21.09 //y=7.4 //x2=15.885 //y2=5.02
cc_431 ( N_VDD_c_390_p N_noxref_7_M31_noxref_d ) capacitor c=0.0140984f \
 //x=16.385 //y=7.4 //x2=15.885 //y2=5.02
cc_432 ( N_VDD_c_270_n N_noxref_7_M31_noxref_d ) capacitor c=6.94454e-19 \
 //x=18.13 //y=7.4 //x2=15.885 //y2=5.02
cc_433 ( N_VDD_M32_noxref_d N_noxref_7_M31_noxref_d ) capacitor c=0.0664752f \
 //x=16.325 //y=5.02 //x2=15.885 //y2=5.02
cc_434 ( N_VDD_c_272_p N_noxref_7_M33_noxref_d ) capacitor c=0.00285083f \
 //x=21.09 //y=7.4 //x2=16.765 //y2=5.02
cc_435 ( N_VDD_c_419_p N_noxref_7_M33_noxref_d ) capacitor c=0.0140984f \
 //x=17.265 //y=7.4 //x2=16.765 //y2=5.02
cc_436 ( N_VDD_c_270_n N_noxref_7_M33_noxref_d ) capacitor c=0.0120541f \
 //x=18.13 //y=7.4 //x2=16.765 //y2=5.02
cc_437 ( N_VDD_M31_noxref_s N_noxref_7_M33_noxref_d ) capacitor c=0.00111971f \
 //x=15.455 //y=5.02 //x2=16.765 //y2=5.02
cc_438 ( N_VDD_M32_noxref_d N_noxref_7_M33_noxref_d ) capacitor c=0.0664752f \
 //x=16.325 //y=5.02 //x2=16.765 //y2=5.02
cc_439 ( N_VDD_M34_noxref_d N_noxref_7_M33_noxref_d ) capacitor c=0.0664752f \
 //x=17.205 //y=5.02 //x2=16.765 //y2=5.02
cc_440 ( N_VDD_M35_noxref_s N_noxref_7_M33_noxref_d ) capacitor c=4.54516e-19 \
 //x=18.785 //y=5.02 //x2=16.765 //y2=5.02
cc_441 ( N_VDD_c_272_p N_noxref_8_c_1542_n ) capacitor c=0.035625f //x=21.09 \
 //y=7.4 //x2=9.875 //y2=4.07
cc_442 ( N_VDD_c_372_p N_noxref_8_c_1542_n ) capacitor c=0.00113322f //x=1.885 \
 //y=7.4 //x2=9.875 //y2=4.07
cc_443 ( N_VDD_c_266_n N_noxref_8_c_1542_n ) capacitor c=0.0140578f //x=4.81 \
 //y=7.4 //x2=9.875 //y2=4.07
cc_444 ( N_VDD_c_267_n N_noxref_8_c_1542_n ) capacitor c=0.0140578f //x=8.14 \
 //y=7.4 //x2=9.875 //y2=4.07
cc_445 ( N_VDD_c_272_p N_noxref_8_c_1543_n ) capacitor c=0.00189266f //x=21.09 \
 //y=7.4 //x2=1.225 //y2=4.07
cc_446 ( N_VDD_c_264_n N_noxref_8_c_1543_n ) capacitor c=0.0017219f //x=0.74 \
 //y=7.4 //x2=1.225 //y2=4.07
cc_447 ( N_VDD_M13_noxref_s N_noxref_8_c_1543_n ) capacitor c=0.00128242f \
 //x=0.955 //y=5.02 //x2=1.225 //y2=4.07
cc_448 ( N_VDD_c_272_p N_noxref_8_c_1572_n ) capacitor c=0.0158405f //x=21.09 \
 //y=7.4 //x2=13.945 //y2=4.07
cc_449 ( N_VDD_c_268_n N_noxref_8_c_1572_n ) capacitor c=0.0140578f //x=11.47 \
 //y=7.4 //x2=13.945 //y2=4.07
cc_450 ( N_VDD_c_272_p N_noxref_8_c_1544_n ) capacitor c=0.0403235f //x=21.09 \
 //y=7.4 //x2=19.865 //y2=4.07
cc_451 ( N_VDD_c_458_p N_noxref_8_c_1544_n ) capacitor c=0.00161566f //x=14.63 \
 //y=7.4 //x2=19.865 //y2=4.07
cc_452 ( N_VDD_c_459_p N_noxref_8_c_1544_n ) capacitor c=0.00172186f \
 //x=15.505 //y=7.4 //x2=19.865 //y2=4.07
cc_453 ( N_VDD_c_390_p N_noxref_8_c_1544_n ) capacitor c=6.61469e-19 \
 //x=16.385 //y=7.4 //x2=19.865 //y2=4.07
cc_454 ( N_VDD_c_461_p N_noxref_8_c_1544_n ) capacitor c=0.00168692f //x=17.96 \
 //y=7.4 //x2=19.865 //y2=4.07
cc_455 ( N_VDD_c_462_p N_noxref_8_c_1544_n ) capacitor c=0.00172186f \
 //x=18.835 //y=7.4 //x2=19.865 //y2=4.07
cc_456 ( N_VDD_c_430_p N_noxref_8_c_1544_n ) capacitor c=6.61469e-19 \
 //x=19.715 //y=7.4 //x2=19.865 //y2=4.07
cc_457 ( N_VDD_c_269_n N_noxref_8_c_1544_n ) capacitor c=0.0269494f //x=14.8 \
 //y=7.4 //x2=19.865 //y2=4.07
cc_458 ( N_VDD_c_270_n N_noxref_8_c_1544_n ) capacitor c=0.0269494f //x=18.13 \
 //y=7.4 //x2=19.865 //y2=4.07
cc_459 ( N_VDD_M31_noxref_s N_noxref_8_c_1544_n ) capacitor c=0.00363031f \
 //x=15.455 //y=5.02 //x2=19.865 //y2=4.07
cc_460 ( N_VDD_M34_noxref_d N_noxref_8_c_1544_n ) capacitor c=5.05307e-19 \
 //x=17.205 //y=5.02 //x2=19.865 //y2=4.07
cc_461 ( N_VDD_M35_noxref_s N_noxref_8_c_1544_n ) capacitor c=0.00363031f \
 //x=18.785 //y=5.02 //x2=19.865 //y2=4.07
cc_462 ( N_VDD_c_272_p N_noxref_8_c_1586_n ) capacitor c=0.00172491f //x=21.09 \
 //y=7.4 //x2=14.175 //y2=4.07
cc_463 ( N_VDD_c_269_n N_noxref_8_c_1586_n ) capacitor c=0.00104972f //x=14.8 \
 //y=7.4 //x2=14.175 //y2=4.07
cc_464 ( N_VDD_M30_noxref_d N_noxref_8_c_1586_n ) capacitor c=5.14736e-19 \
 //x=13.875 //y=5.02 //x2=14.175 //y2=4.07
cc_465 ( N_VDD_c_272_p N_noxref_8_c_1545_n ) capacitor c=9.2251e-19 //x=21.09 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_466 ( N_VDD_c_264_n N_noxref_8_c_1545_n ) capacitor c=0.0159723f //x=0.74 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_467 ( N_VDD_M13_noxref_s N_noxref_8_c_1545_n ) capacitor c=0.0122951f \
 //x=0.955 //y=5.02 //x2=1.11 //y2=2.08
cc_468 ( N_VDD_c_267_n N_noxref_8_c_1546_n ) capacitor c=4.57806e-19 //x=8.14 \
 //y=7.4 //x2=9.99 //y2=2.08
cc_469 ( N_VDD_c_268_n N_noxref_8_c_1546_n ) capacitor c=3.69525e-19 //x=11.47 \
 //y=7.4 //x2=9.99 //y2=2.08
cc_470 ( N_VDD_c_272_p N_noxref_8_c_1594_n ) capacitor c=0.00453473f //x=21.09 \
 //y=7.4 //x2=13.495 //y2=5.2
cc_471 ( N_VDD_c_320_p N_noxref_8_c_1594_n ) capacitor c=4.48391e-19 \
 //x=13.055 //y=7.4 //x2=13.495 //y2=5.2
cc_472 ( N_VDD_c_365_p N_noxref_8_c_1594_n ) capacitor c=4.48377e-19 \
 //x=13.935 //y=7.4 //x2=13.495 //y2=5.2
cc_473 ( N_VDD_M28_noxref_d N_noxref_8_c_1594_n ) capacitor c=0.0124506f \
 //x=12.995 //y=5.02 //x2=13.495 //y2=5.2
cc_474 ( N_VDD_c_268_n N_noxref_8_c_1598_n ) capacitor c=0.00985474f //x=11.47 \
 //y=7.4 //x2=12.785 //y2=5.2
cc_475 ( N_VDD_M27_noxref_s N_noxref_8_c_1598_n ) capacitor c=0.087833f \
 //x=12.125 //y=5.02 //x2=12.785 //y2=5.2
cc_476 ( N_VDD_c_272_p N_noxref_8_c_1600_n ) capacitor c=0.00307016f //x=21.09 \
 //y=7.4 //x2=13.975 //y2=5.2
cc_477 ( N_VDD_c_365_p N_noxref_8_c_1600_n ) capacitor c=7.73167e-19 \
 //x=13.935 //y=7.4 //x2=13.975 //y2=5.2
cc_478 ( N_VDD_M30_noxref_d N_noxref_8_c_1600_n ) capacitor c=0.016133f \
 //x=13.875 //y=5.02 //x2=13.975 //y2=5.2
cc_479 ( N_VDD_M31_noxref_s N_noxref_8_c_1600_n ) capacitor c=2.44532e-19 \
 //x=15.455 //y=5.02 //x2=13.975 //y2=5.2
cc_480 ( N_VDD_c_268_n N_noxref_8_c_1549_n ) capacitor c=0.00151618f //x=11.47 \
 //y=7.4 //x2=14.06 //y2=4.07
cc_481 ( N_VDD_c_269_n N_noxref_8_c_1549_n ) capacitor c=0.0451944f //x=14.8 \
 //y=7.4 //x2=14.06 //y2=4.07
cc_482 ( N_VDD_c_265_n N_noxref_8_c_1550_n ) capacitor c=6.61994e-19 //x=21.09 \
 //y=7.4 //x2=19.98 //y2=2.08
cc_483 ( N_VDD_c_270_n N_noxref_8_c_1550_n ) capacitor c=6.2696e-19 //x=18.13 \
 //y=7.4 //x2=19.98 //y2=2.08
cc_484 ( N_VDD_c_372_p N_noxref_8_M13_noxref_g ) capacitor c=0.00749687f \
 //x=1.885 //y=7.4 //x2=1.31 //y2=6.02
cc_485 ( N_VDD_M13_noxref_s N_noxref_8_M13_noxref_g ) capacitor c=0.0477201f \
 //x=0.955 //y=5.02 //x2=1.31 //y2=6.02
cc_486 ( N_VDD_c_372_p N_noxref_8_M14_noxref_g ) capacitor c=0.00675175f \
 //x=1.885 //y=7.4 //x2=1.75 //y2=6.02
cc_487 ( N_VDD_M14_noxref_d N_noxref_8_M14_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=1.75 //y2=6.02
cc_488 ( N_VDD_c_309_p N_noxref_8_M25_noxref_g ) capacitor c=0.00673971f \
 //x=10.605 //y=7.4 //x2=10.03 //y2=6.02
cc_489 ( N_VDD_M24_noxref_d N_noxref_8_M25_noxref_g ) capacitor c=0.015318f \
 //x=9.665 //y=5.02 //x2=10.03 //y2=6.02
cc_490 ( N_VDD_c_309_p N_noxref_8_M26_noxref_g ) capacitor c=0.00672952f \
 //x=10.605 //y=7.4 //x2=10.47 //y2=6.02
cc_491 ( N_VDD_c_268_n N_noxref_8_M26_noxref_g ) capacitor c=0.00864163f \
 //x=11.47 //y=7.4 //x2=10.47 //y2=6.02
cc_492 ( N_VDD_M26_noxref_d N_noxref_8_M26_noxref_g ) capacitor c=0.0430452f \
 //x=10.545 //y=5.02 //x2=10.47 //y2=6.02
cc_493 ( N_VDD_c_500_p N_noxref_8_M37_noxref_g ) capacitor c=0.00673971f \
 //x=20.595 //y=7.4 //x2=20.02 //y2=6.02
cc_494 ( N_VDD_M36_noxref_d N_noxref_8_M37_noxref_g ) capacitor c=0.015318f \
 //x=19.655 //y=5.02 //x2=20.02 //y2=6.02
cc_495 ( N_VDD_c_500_p N_noxref_8_M38_noxref_g ) capacitor c=0.00672952f \
 //x=20.595 //y=7.4 //x2=20.46 //y2=6.02
cc_496 ( N_VDD_c_265_n N_noxref_8_M38_noxref_g ) capacitor c=0.024326f \
 //x=21.09 //y=7.4 //x2=20.46 //y2=6.02
cc_497 ( N_VDD_M38_noxref_d N_noxref_8_M38_noxref_g ) capacitor c=0.0430452f \
 //x=20.535 //y=5.02 //x2=20.46 //y2=6.02
cc_498 ( N_VDD_c_264_n N_noxref_8_c_1622_n ) capacitor c=0.00757682f //x=0.74 \
 //y=7.4 //x2=1.385 //y2=4.79
cc_499 ( N_VDD_M13_noxref_s N_noxref_8_c_1622_n ) capacitor c=0.00445117f \
 //x=0.955 //y=5.02 //x2=1.385 //y2=4.79
cc_500 ( N_VDD_c_272_p N_noxref_8_M27_noxref_d ) capacitor c=0.00275225f \
 //x=21.09 //y=7.4 //x2=12.555 //y2=5.02
cc_501 ( N_VDD_c_320_p N_noxref_8_M27_noxref_d ) capacitor c=0.0140317f \
 //x=13.055 //y=7.4 //x2=12.555 //y2=5.02
cc_502 ( N_VDD_c_269_n N_noxref_8_M27_noxref_d ) capacitor c=6.94454e-19 \
 //x=14.8 //y=7.4 //x2=12.555 //y2=5.02
cc_503 ( N_VDD_M28_noxref_d N_noxref_8_M27_noxref_d ) capacitor c=0.0664752f \
 //x=12.995 //y=5.02 //x2=12.555 //y2=5.02
cc_504 ( N_VDD_c_272_p N_noxref_8_M29_noxref_d ) capacitor c=0.00285083f \
 //x=21.09 //y=7.4 //x2=13.435 //y2=5.02
cc_505 ( N_VDD_c_365_p N_noxref_8_M29_noxref_d ) capacitor c=0.0140984f \
 //x=13.935 //y=7.4 //x2=13.435 //y2=5.02
cc_506 ( N_VDD_c_269_n N_noxref_8_M29_noxref_d ) capacitor c=0.0120541f \
 //x=14.8 //y=7.4 //x2=13.435 //y2=5.02
cc_507 ( N_VDD_M27_noxref_s N_noxref_8_M29_noxref_d ) capacitor c=0.00111971f \
 //x=12.125 //y=5.02 //x2=13.435 //y2=5.02
cc_508 ( N_VDD_M28_noxref_d N_noxref_8_M29_noxref_d ) capacitor c=0.0664752f \
 //x=12.995 //y=5.02 //x2=13.435 //y2=5.02
cc_509 ( N_VDD_M30_noxref_d N_noxref_8_M29_noxref_d ) capacitor c=0.0664752f \
 //x=13.875 //y=5.02 //x2=13.435 //y2=5.02
cc_510 ( N_VDD_M31_noxref_s N_noxref_8_M29_noxref_d ) capacitor c=4.54516e-19 \
 //x=15.455 //y=5.02 //x2=13.435 //y2=5.02
cc_511 ( N_VDD_c_272_p N_Q_c_1900_n ) capacitor c=0.0163573f //x=21.09 //y=7.4 \
 //x2=20.605 //y2=3.7
cc_512 ( N_VDD_M38_noxref_d N_Q_c_1900_n ) capacitor c=4.05358e-19 //x=20.535 \
 //y=5.02 //x2=20.605 //y2=3.7
cc_513 ( N_VDD_c_265_n Q ) capacitor c=0.0466813f //x=21.09 //y=7.4 //x2=20.72 \
 //y2=2.22
cc_514 ( N_VDD_c_270_n Q ) capacitor c=0.00151618f //x=18.13 //y=7.4 \
 //x2=20.72 //y2=2.22
cc_515 ( N_VDD_c_269_n N_Q_c_1903_n ) capacitor c=9.06385e-19 //x=14.8 //y=7.4 \
 //x2=16.65 //y2=2.08
cc_516 ( N_VDD_c_270_n N_Q_c_1903_n ) capacitor c=5.81514e-19 //x=18.13 \
 //y=7.4 //x2=16.65 //y2=2.08
cc_517 ( N_VDD_c_272_p N_Q_c_1915_n ) capacitor c=0.00459955f //x=21.09 \
 //y=7.4 //x2=20.155 //y2=5.2
cc_518 ( N_VDD_c_430_p N_Q_c_1915_n ) capacitor c=4.48705e-19 //x=19.715 \
 //y=7.4 //x2=20.155 //y2=5.2
cc_519 ( N_VDD_c_500_p N_Q_c_1915_n ) capacitor c=4.48693e-19 //x=20.595 \
 //y=7.4 //x2=20.155 //y2=5.2
cc_520 ( N_VDD_M36_noxref_d N_Q_c_1915_n ) capacitor c=0.01269f //x=19.655 \
 //y=5.02 //x2=20.155 //y2=5.2
cc_521 ( N_VDD_c_270_n N_Q_c_1919_n ) capacitor c=0.00985474f //x=18.13 \
 //y=7.4 //x2=19.445 //y2=5.2
cc_522 ( N_VDD_M35_noxref_s N_Q_c_1919_n ) capacitor c=0.087833f //x=18.785 \
 //y=5.02 //x2=19.445 //y2=5.2
cc_523 ( N_VDD_c_272_p N_Q_c_1921_n ) capacitor c=0.00311875f //x=21.09 \
 //y=7.4 //x2=20.635 //y2=5.2
cc_524 ( N_VDD_c_500_p N_Q_c_1921_n ) capacitor c=7.21492e-19 //x=20.595 \
 //y=7.4 //x2=20.635 //y2=5.2
cc_525 ( N_VDD_M38_noxref_d N_Q_c_1921_n ) capacitor c=0.0163364f //x=20.535 \
 //y=5.02 //x2=20.635 //y2=5.2
cc_526 ( N_VDD_c_419_p N_Q_M33_noxref_g ) capacitor c=0.00673971f //x=17.265 \
 //y=7.4 //x2=16.69 //y2=6.02
cc_527 ( N_VDD_M32_noxref_d N_Q_M33_noxref_g ) capacitor c=0.015318f \
 //x=16.325 //y=5.02 //x2=16.69 //y2=6.02
cc_528 ( N_VDD_c_419_p N_Q_M34_noxref_g ) capacitor c=0.00672952f //x=17.265 \
 //y=7.4 //x2=17.13 //y2=6.02
cc_529 ( N_VDD_c_270_n N_Q_M34_noxref_g ) capacitor c=0.00864163f //x=18.13 \
 //y=7.4 //x2=17.13 //y2=6.02
cc_530 ( N_VDD_M34_noxref_d N_Q_M34_noxref_g ) capacitor c=0.0430452f \
 //x=17.205 //y=5.02 //x2=17.13 //y2=6.02
cc_531 ( N_VDD_c_272_p N_Q_M35_noxref_d ) capacitor c=0.00285083f //x=21.09 \
 //y=7.4 //x2=19.215 //y2=5.02
cc_532 ( N_VDD_c_430_p N_Q_M35_noxref_d ) capacitor c=0.0140984f //x=19.715 \
 //y=7.4 //x2=19.215 //y2=5.02
cc_533 ( N_VDD_c_265_n N_Q_M35_noxref_d ) capacitor c=6.94454e-19 //x=21.09 \
 //y=7.4 //x2=19.215 //y2=5.02
cc_534 ( N_VDD_M36_noxref_d N_Q_M35_noxref_d ) capacitor c=0.0664752f \
 //x=19.655 //y=5.02 //x2=19.215 //y2=5.02
cc_535 ( N_VDD_c_272_p N_Q_M37_noxref_d ) capacitor c=0.00294217f //x=21.09 \
 //y=7.4 //x2=20.095 //y2=5.02
cc_536 ( N_VDD_c_500_p N_Q_M37_noxref_d ) capacitor c=0.0138379f //x=20.595 \
 //y=7.4 //x2=20.095 //y2=5.02
cc_537 ( N_VDD_c_265_n N_Q_M37_noxref_d ) capacitor c=0.0123189f //x=21.09 \
 //y=7.4 //x2=20.095 //y2=5.02
cc_538 ( N_VDD_M35_noxref_s N_Q_M37_noxref_d ) capacitor c=0.00111971f \
 //x=18.785 //y=5.02 //x2=20.095 //y2=5.02
cc_539 ( N_VDD_M36_noxref_d N_Q_M37_noxref_d ) capacitor c=0.0664752f \
 //x=19.655 //y=5.02 //x2=20.095 //y2=5.02
cc_540 ( N_VDD_M38_noxref_d N_Q_M37_noxref_d ) capacitor c=0.0664752f \
 //x=20.535 //y=5.02 //x2=20.095 //y2=5.02
cc_541 ( N_VDD_c_266_n N_D_c_2158_n ) capacitor c=4.47073e-19 //x=4.81 //y=7.4 \
 //x2=6.66 //y2=2.08
cc_542 ( N_VDD_c_267_n N_D_c_2158_n ) capacitor c=3.37458e-19 //x=8.14 //y=7.4 \
 //x2=6.66 //y2=2.08
cc_543 ( N_VDD_c_274_p N_D_M21_noxref_g ) capacitor c=0.00673971f //x=7.275 \
 //y=7.4 //x2=6.7 //y2=6.02
cc_544 ( N_VDD_M20_noxref_d N_D_M21_noxref_g ) capacitor c=0.015318f //x=6.335 \
 //y=5.02 //x2=6.7 //y2=6.02
cc_545 ( N_VDD_c_274_p N_D_M22_noxref_g ) capacitor c=0.00672952f //x=7.275 \
 //y=7.4 //x2=7.14 //y2=6.02
cc_546 ( N_VDD_c_267_n N_D_M22_noxref_g ) capacitor c=0.00864163f //x=8.14 \
 //y=7.4 //x2=7.14 //y2=6.02
cc_547 ( N_VDD_M22_noxref_d N_D_M22_noxref_g ) capacitor c=0.0430452f \
 //x=7.215 //y=5.02 //x2=7.14 //y2=6.02
cc_548 ( N_noxref_3_c_561_n N_noxref_4_c_791_n ) capacitor c=0.011463f \
 //x=9.135 //y=3.33 //x2=10.845 //y2=3.33
cc_549 ( N_noxref_3_M24_noxref_g N_noxref_4_c_808_n ) capacitor c=0.0169521f \
 //x=9.59 //y=6.02 //x2=10.165 //y2=5.2
cc_550 ( N_noxref_3_c_569_n N_noxref_4_c_812_n ) capacitor c=0.00539951f \
 //x=9.25 //y=2.08 //x2=9.455 //y2=5.2
cc_551 ( N_noxref_3_M23_noxref_g N_noxref_4_c_812_n ) capacitor c=0.0177326f \
 //x=9.15 //y=6.02 //x2=9.455 //y2=5.2
cc_552 ( N_noxref_3_c_607_n N_noxref_4_c_812_n ) capacitor c=0.00581252f \
 //x=9.25 //y=4.7 //x2=9.455 //y2=5.2
cc_553 ( N_noxref_3_c_568_n N_noxref_4_c_793_n ) capacitor c=3.49822e-19 \
 //x=7.4 //y=3.33 //x2=10.73 //y2=3.33
cc_554 ( N_noxref_3_c_569_n N_noxref_4_c_793_n ) capacitor c=0.00318783f \
 //x=9.25 //y=2.08 //x2=10.73 //y2=3.33
cc_555 ( N_noxref_3_M24_noxref_g N_noxref_4_M23_noxref_d ) capacitor \
 c=0.0173476f //x=9.59 //y=6.02 //x2=9.225 //y2=5.02
cc_556 ( N_noxref_3_c_555_n N_CLK_c_940_n ) capacitor c=0.00360213f //x=7.285 \
 //y=3.33 //x2=13.205 //y2=4.44
cc_557 ( N_noxref_3_c_560_n N_CLK_c_940_n ) capacitor c=4.49102e-19 //x=3.445 \
 //y=3.33 //x2=13.205 //y2=4.44
cc_558 ( N_noxref_3_c_566_n N_CLK_c_940_n ) capacitor c=0.0200057f //x=3.33 \
 //y=2.08 //x2=13.205 //y2=4.44
cc_559 ( N_noxref_3_c_584_n N_CLK_c_940_n ) capacitor c=0.0185297f //x=6.835 \
 //y=5.2 //x2=13.205 //y2=4.44
cc_560 ( N_noxref_3_c_588_n N_CLK_c_940_n ) capacitor c=0.0181237f //x=6.125 \
 //y=5.2 //x2=13.205 //y2=4.44
cc_561 ( N_noxref_3_c_568_n N_CLK_c_940_n ) capacitor c=0.0208321f //x=7.4 \
 //y=3.33 //x2=13.205 //y2=4.44
cc_562 ( N_noxref_3_c_569_n N_CLK_c_940_n ) capacitor c=0.0198304f //x=9.25 \
 //y=2.08 //x2=13.205 //y2=4.44
cc_563 ( N_noxref_3_c_634_p N_CLK_c_940_n ) capacitor c=0.0111881f //x=3.33 \
 //y=4.7 //x2=13.205 //y2=4.44
cc_564 ( N_noxref_3_c_607_n N_CLK_c_940_n ) capacitor c=0.0107057f //x=9.25 \
 //y=4.7 //x2=13.205 //y2=4.44
cc_565 ( N_noxref_3_c_566_n N_CLK_c_958_n ) capacitor c=0.00153281f //x=3.33 \
 //y=2.08 //x2=2.335 //y2=4.44
cc_566 ( N_noxref_3_c_560_n N_CLK_c_937_n ) capacitor c=0.00526349f //x=3.445 \
 //y=3.33 //x2=2.22 //y2=2.08
cc_567 ( N_noxref_3_c_566_n N_CLK_c_937_n ) capacitor c=0.0511464f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_568 ( N_noxref_3_c_639_p N_CLK_c_937_n ) capacitor c=0.00228632f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_569 ( N_noxref_3_c_634_p N_CLK_c_937_n ) capacitor c=0.00218014f //x=3.33 \
 //y=4.7 //x2=2.22 //y2=2.08
cc_570 ( N_noxref_3_M17_noxref_g N_CLK_M15_noxref_g ) capacitor c=0.0101598f \
 //x=3.07 //y=6.02 //x2=2.19 //y2=6.02
cc_571 ( N_noxref_3_M17_noxref_g N_CLK_M16_noxref_g ) capacitor c=0.0602553f \
 //x=3.07 //y=6.02 //x2=2.63 //y2=6.02
cc_572 ( N_noxref_3_M18_noxref_g N_CLK_M16_noxref_g ) capacitor c=0.0101598f \
 //x=3.51 //y=6.02 //x2=2.63 //y2=6.02
cc_573 ( N_noxref_3_c_644_p N_CLK_c_989_n ) capacitor c=0.00456962f //x=3.32 \
 //y=0.915 //x2=2.31 //y2=0.91
cc_574 ( N_noxref_3_c_645_p N_CLK_c_990_n ) capacitor c=0.00438372f //x=3.32 \
 //y=1.26 //x2=2.31 //y2=1.22
cc_575 ( N_noxref_3_c_646_p N_CLK_c_991_n ) capacitor c=0.00438372f //x=3.32 \
 //y=1.57 //x2=2.31 //y2=1.45
cc_576 ( N_noxref_3_c_566_n N_CLK_c_992_n ) capacitor c=0.0023343f //x=3.33 \
 //y=2.08 //x2=2.31 //y2=1.915
cc_577 ( N_noxref_3_c_639_p N_CLK_c_992_n ) capacitor c=0.00933826f //x=3.33 \
 //y=2.08 //x2=2.31 //y2=1.915
cc_578 ( N_noxref_3_c_649_p N_CLK_c_992_n ) capacitor c=0.00438372f //x=3.33 \
 //y=1.915 //x2=2.31 //y2=1.915
cc_579 ( N_noxref_3_c_634_p N_CLK_c_995_n ) capacitor c=0.0611812f //x=3.33 \
 //y=4.7 //x2=2.555 //y2=4.79
cc_580 ( N_noxref_3_c_566_n N_CLK_c_996_n ) capacitor c=0.00142741f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=4.7
cc_581 ( N_noxref_3_c_634_p N_CLK_c_996_n ) capacitor c=0.00487508f //x=3.33 \
 //y=4.7 //x2=2.22 //y2=4.7
cc_582 ( N_noxref_3_c_555_n N_noxref_6_c_1215_n ) capacitor c=0.146341f \
 //x=7.285 //y=3.33 //x2=5.805 //y2=3.7
cc_583 ( N_noxref_3_c_555_n N_noxref_6_c_1216_n ) capacitor c=0.0294746f \
 //x=7.285 //y=3.33 //x2=4.185 //y2=3.7
cc_584 ( N_noxref_3_c_566_n N_noxref_6_c_1216_n ) capacitor c=0.00687545f \
 //x=3.33 //y=2.08 //x2=4.185 //y2=3.7
cc_585 ( N_noxref_3_c_555_n N_noxref_6_c_1142_n ) capacitor c=0.108749f \
 //x=7.285 //y=3.33 //x2=15.795 //y2=3.7
cc_586 ( N_noxref_3_c_561_n N_noxref_6_c_1142_n ) capacitor c=0.175696f \
 //x=9.135 //y=3.33 //x2=15.795 //y2=3.7
cc_587 ( N_noxref_3_c_565_n N_noxref_6_c_1142_n ) capacitor c=0.0267668f \
 //x=7.515 //y=3.33 //x2=15.795 //y2=3.7
cc_588 ( N_noxref_3_c_568_n N_noxref_6_c_1142_n ) capacitor c=0.0206034f \
 //x=7.4 //y=3.33 //x2=15.795 //y2=3.7
cc_589 ( N_noxref_3_c_569_n N_noxref_6_c_1142_n ) capacitor c=0.0205831f \
 //x=9.25 //y=2.08 //x2=15.795 //y2=3.7
cc_590 ( N_noxref_3_c_555_n N_noxref_6_c_1223_n ) capacitor c=0.0266674f \
 //x=7.285 //y=3.33 //x2=6.035 //y2=3.7
cc_591 ( N_noxref_3_M17_noxref_g N_noxref_6_c_1175_n ) capacitor c=0.01736f \
 //x=3.07 //y=6.02 //x2=3.205 //y2=5.155
cc_592 ( N_noxref_3_M18_noxref_g N_noxref_6_c_1179_n ) capacitor c=0.0194981f \
 //x=3.51 //y=6.02 //x2=3.985 //y2=5.155
cc_593 ( N_noxref_3_c_634_p N_noxref_6_c_1179_n ) capacitor c=0.00201851f \
 //x=3.33 //y=4.7 //x2=3.985 //y2=5.155
cc_594 ( N_noxref_3_c_665_p N_noxref_6_c_1144_n ) capacitor c=0.00359704f \
 //x=3.695 //y=1.415 //x2=3.985 //y2=1.665
cc_595 ( N_noxref_3_c_666_p N_noxref_6_c_1144_n ) capacitor c=0.00457401f \
 //x=3.85 //y=1.26 //x2=3.985 //y2=1.665
cc_596 ( N_noxref_3_c_555_n N_noxref_6_c_1229_n ) capacitor c=0.00628992f \
 //x=7.285 //y=3.33 //x2=3.67 //y2=1.665
cc_597 ( N_noxref_3_c_555_n N_noxref_6_c_1183_n ) capacitor c=0.0260398f \
 //x=7.285 //y=3.33 //x2=4.07 //y2=3.7
cc_598 ( N_noxref_3_c_560_n N_noxref_6_c_1183_n ) capacitor c=0.00117715f \
 //x=3.445 //y=3.33 //x2=4.07 //y2=3.7
cc_599 ( N_noxref_3_c_566_n N_noxref_6_c_1183_n ) capacitor c=0.0831612f \
 //x=3.33 //y=2.08 //x2=4.07 //y2=3.7
cc_600 ( N_noxref_3_c_568_n N_noxref_6_c_1183_n ) capacitor c=3.52729e-19 \
 //x=7.4 //y=3.33 //x2=4.07 //y2=3.7
cc_601 ( N_noxref_3_c_639_p N_noxref_6_c_1183_n ) capacitor c=0.00877984f \
 //x=3.33 //y=2.08 //x2=4.07 //y2=3.7
cc_602 ( N_noxref_3_c_649_p N_noxref_6_c_1183_n ) capacitor c=0.00283672f \
 //x=3.33 //y=1.915 //x2=4.07 //y2=3.7
cc_603 ( N_noxref_3_c_634_p N_noxref_6_c_1183_n ) capacitor c=0.013693f \
 //x=3.33 //y=4.7 //x2=4.07 //y2=3.7
cc_604 ( N_noxref_3_c_555_n N_noxref_6_c_1145_n ) capacitor c=0.0257693f \
 //x=7.285 //y=3.33 //x2=5.92 //y2=2.08
cc_605 ( N_noxref_3_c_566_n N_noxref_6_c_1145_n ) capacitor c=9.66956e-19 \
 //x=3.33 //y=2.08 //x2=5.92 //y2=2.08
cc_606 ( N_noxref_3_c_588_n N_noxref_6_c_1145_n ) capacitor c=0.00521572f \
 //x=6.125 //y=5.2 //x2=5.92 //y2=2.08
cc_607 ( N_noxref_3_c_568_n N_noxref_6_c_1145_n ) capacitor c=0.00319084f \
 //x=7.4 //y=3.33 //x2=5.92 //y2=2.08
cc_608 ( N_noxref_3_c_566_n N_noxref_6_c_1241_n ) capacitor c=0.0171303f \
 //x=3.33 //y=2.08 //x2=3.29 //y2=5.155
cc_609 ( N_noxref_3_c_634_p N_noxref_6_c_1241_n ) capacitor c=0.00475601f \
 //x=3.33 //y=4.7 //x2=3.29 //y2=5.155
cc_610 ( N_noxref_3_c_588_n N_noxref_6_M19_noxref_g ) capacitor c=0.0177326f \
 //x=6.125 //y=5.2 //x2=5.82 //y2=6.02
cc_611 ( N_noxref_3_c_584_n N_noxref_6_M20_noxref_g ) capacitor c=0.0169521f \
 //x=6.835 //y=5.2 //x2=6.26 //y2=6.02
cc_612 ( N_noxref_3_M19_noxref_d N_noxref_6_M20_noxref_g ) capacitor \
 c=0.0173476f //x=5.895 //y=5.02 //x2=6.26 //y2=6.02
cc_613 ( N_noxref_3_c_588_n N_noxref_6_c_1198_n ) capacitor c=0.00581252f \
 //x=6.125 //y=5.2 //x2=5.92 //y2=4.7
cc_614 ( N_noxref_3_c_644_p N_noxref_6_M2_noxref_d ) capacitor c=0.00217566f \
 //x=3.32 //y=0.915 //x2=3.395 //y2=0.915
cc_615 ( N_noxref_3_c_645_p N_noxref_6_M2_noxref_d ) capacitor c=0.0034598f \
 //x=3.32 //y=1.26 //x2=3.395 //y2=0.915
cc_616 ( N_noxref_3_c_646_p N_noxref_6_M2_noxref_d ) capacitor c=0.00544291f \
 //x=3.32 //y=1.57 //x2=3.395 //y2=0.915
cc_617 ( N_noxref_3_c_688_p N_noxref_6_M2_noxref_d ) capacitor c=0.00241102f \
 //x=3.695 //y=0.76 //x2=3.395 //y2=0.915
cc_618 ( N_noxref_3_c_665_p N_noxref_6_M2_noxref_d ) capacitor c=0.0140297f \
 //x=3.695 //y=1.415 //x2=3.395 //y2=0.915
cc_619 ( N_noxref_3_c_690_p N_noxref_6_M2_noxref_d ) capacitor c=0.00219619f \
 //x=3.85 //y=0.915 //x2=3.395 //y2=0.915
cc_620 ( N_noxref_3_c_666_p N_noxref_6_M2_noxref_d ) capacitor c=0.00603828f \
 //x=3.85 //y=1.26 //x2=3.395 //y2=0.915
cc_621 ( N_noxref_3_c_649_p N_noxref_6_M2_noxref_d ) capacitor c=0.00661782f \
 //x=3.33 //y=1.915 //x2=3.395 //y2=0.915
cc_622 ( N_noxref_3_M17_noxref_g N_noxref_6_M17_noxref_d ) capacitor \
 c=0.0180032f //x=3.07 //y=6.02 //x2=3.145 //y2=5.02
cc_623 ( N_noxref_3_M18_noxref_g N_noxref_6_M17_noxref_d ) capacitor \
 c=0.0194246f //x=3.51 //y=6.02 //x2=3.145 //y2=5.02
cc_624 ( N_noxref_3_c_555_n N_noxref_8_c_1542_n ) capacitor c=0.0428508f \
 //x=7.285 //y=3.33 //x2=9.875 //y2=4.07
cc_625 ( N_noxref_3_c_560_n N_noxref_8_c_1542_n ) capacitor c=0.0135672f \
 //x=3.445 //y=3.33 //x2=9.875 //y2=4.07
cc_626 ( N_noxref_3_c_561_n N_noxref_8_c_1542_n ) capacitor c=0.0110241f \
 //x=9.135 //y=3.33 //x2=9.875 //y2=4.07
cc_627 ( N_noxref_3_c_565_n N_noxref_8_c_1542_n ) capacitor c=5.70661e-19 \
 //x=7.515 //y=3.33 //x2=9.875 //y2=4.07
cc_628 ( N_noxref_3_c_566_n N_noxref_8_c_1542_n ) capacitor c=0.0206302f \
 //x=3.33 //y=2.08 //x2=9.875 //y2=4.07
cc_629 ( N_noxref_3_c_568_n N_noxref_8_c_1542_n ) capacitor c=0.0181936f \
 //x=7.4 //y=3.33 //x2=9.875 //y2=4.07
cc_630 ( N_noxref_3_c_569_n N_noxref_8_c_1542_n ) capacitor c=0.0184765f \
 //x=9.25 //y=2.08 //x2=9.875 //y2=4.07
cc_631 ( N_noxref_3_c_569_n N_noxref_8_c_1642_n ) capacitor c=0.00179385f \
 //x=9.25 //y=2.08 //x2=10.105 //y2=4.07
cc_632 ( N_noxref_3_c_566_n N_noxref_8_c_1545_n ) capacitor c=0.00175117f \
 //x=3.33 //y=2.08 //x2=1.11 //y2=2.08
cc_633 ( N_noxref_3_c_569_n N_noxref_8_c_1644_n ) capacitor c=0.00400249f \
 //x=9.25 //y=2.08 //x2=9.99 //y2=4.535
cc_634 ( N_noxref_3_c_607_n N_noxref_8_c_1644_n ) capacitor c=0.00417994f \
 //x=9.25 //y=4.7 //x2=9.99 //y2=4.535
cc_635 ( N_noxref_3_c_561_n N_noxref_8_c_1546_n ) capacitor c=0.00318578f \
 //x=9.135 //y=3.33 //x2=9.99 //y2=2.08
cc_636 ( N_noxref_3_c_568_n N_noxref_8_c_1546_n ) capacitor c=9.69022e-19 \
 //x=7.4 //y=3.33 //x2=9.99 //y2=2.08
cc_637 ( N_noxref_3_c_569_n N_noxref_8_c_1546_n ) capacitor c=0.0794726f \
 //x=9.25 //y=2.08 //x2=9.99 //y2=2.08
cc_638 ( N_noxref_3_c_574_n N_noxref_8_c_1546_n ) capacitor c=0.00308814f \
 //x=9.055 //y=1.915 //x2=9.99 //y2=2.08
cc_639 ( N_noxref_3_M23_noxref_g N_noxref_8_M25_noxref_g ) capacitor \
 c=0.0104611f //x=9.15 //y=6.02 //x2=10.03 //y2=6.02
cc_640 ( N_noxref_3_M24_noxref_g N_noxref_8_M25_noxref_g ) capacitor \
 c=0.106811f //x=9.59 //y=6.02 //x2=10.03 //y2=6.02
cc_641 ( N_noxref_3_M24_noxref_g N_noxref_8_M26_noxref_g ) capacitor \
 c=0.0100341f //x=9.59 //y=6.02 //x2=10.47 //y2=6.02
cc_642 ( N_noxref_3_c_570_n N_noxref_8_c_1653_n ) capacitor c=4.86506e-19 \
 //x=9.055 //y=0.865 //x2=10.025 //y2=0.905
cc_643 ( N_noxref_3_c_572_n N_noxref_8_c_1653_n ) capacitor c=0.00152104f \
 //x=9.055 //y=1.21 //x2=10.025 //y2=0.905
cc_644 ( N_noxref_3_c_577_n N_noxref_8_c_1653_n ) capacitor c=0.0151475f \
 //x=9.585 //y=0.865 //x2=10.025 //y2=0.905
cc_645 ( N_noxref_3_c_573_n N_noxref_8_c_1656_n ) capacitor c=0.00109982f \
 //x=9.055 //y=1.52 //x2=10.025 //y2=1.25
cc_646 ( N_noxref_3_c_579_n N_noxref_8_c_1656_n ) capacitor c=0.0111064f \
 //x=9.585 //y=1.21 //x2=10.025 //y2=1.25
cc_647 ( N_noxref_3_c_573_n N_noxref_8_c_1658_n ) capacitor c=9.57794e-19 \
 //x=9.055 //y=1.52 //x2=10.025 //y2=1.56
cc_648 ( N_noxref_3_c_574_n N_noxref_8_c_1658_n ) capacitor c=0.00662747f \
 //x=9.055 //y=1.915 //x2=10.025 //y2=1.56
cc_649 ( N_noxref_3_c_579_n N_noxref_8_c_1658_n ) capacitor c=0.00862358f \
 //x=9.585 //y=1.21 //x2=10.025 //y2=1.56
cc_650 ( N_noxref_3_c_577_n N_noxref_8_c_1661_n ) capacitor c=0.00124821f \
 //x=9.585 //y=0.865 //x2=10.555 //y2=0.905
cc_651 ( N_noxref_3_c_579_n N_noxref_8_c_1662_n ) capacitor c=0.00200715f \
 //x=9.585 //y=1.21 //x2=10.555 //y2=1.25
cc_652 ( N_noxref_3_c_569_n N_noxref_8_c_1663_n ) capacitor c=0.00307062f \
 //x=9.25 //y=2.08 //x2=9.99 //y2=2.08
cc_653 ( N_noxref_3_c_574_n N_noxref_8_c_1663_n ) capacitor c=0.0179092f \
 //x=9.055 //y=1.915 //x2=9.99 //y2=2.08
cc_654 ( N_noxref_3_c_569_n N_noxref_8_c_1665_n ) capacitor c=0.00344981f \
 //x=9.25 //y=2.08 //x2=10.02 //y2=4.7
cc_655 ( N_noxref_3_c_607_n N_noxref_8_c_1665_n ) capacitor c=0.0293367f \
 //x=9.25 //y=4.7 //x2=10.02 //y2=4.7
cc_656 ( N_noxref_3_c_555_n N_noxref_11_c_2110_n ) capacitor c=2.45218e-19 \
 //x=7.285 //y=3.33 //x2=3.985 //y2=0.54
cc_657 ( N_noxref_3_c_566_n N_noxref_11_c_2110_n ) capacitor c=0.00208521f \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_658 ( N_noxref_3_c_644_p N_noxref_11_c_2110_n ) capacitor c=0.0194423f \
 //x=3.32 //y=0.915 //x2=3.985 //y2=0.54
cc_659 ( N_noxref_3_c_690_p N_noxref_11_c_2110_n ) capacitor c=0.00656458f \
 //x=3.85 //y=0.915 //x2=3.985 //y2=0.54
cc_660 ( N_noxref_3_c_639_p N_noxref_11_c_2110_n ) capacitor c=2.20712e-19 \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_661 ( N_noxref_3_c_645_p N_noxref_11_c_2124_n ) capacitor c=0.00538829f \
 //x=3.32 //y=1.26 //x2=3.1 //y2=0.995
cc_662 ( N_noxref_3_c_644_p N_noxref_11_M2_noxref_s ) capacitor c=0.00538829f \
 //x=3.32 //y=0.915 //x2=2.965 //y2=0.375
cc_663 ( N_noxref_3_c_646_p N_noxref_11_M2_noxref_s ) capacitor c=0.00538829f \
 //x=3.32 //y=1.57 //x2=2.965 //y2=0.375
cc_664 ( N_noxref_3_c_690_p N_noxref_11_M2_noxref_s ) capacitor c=0.0143002f \
 //x=3.85 //y=0.915 //x2=2.965 //y2=0.375
cc_665 ( N_noxref_3_c_666_p N_noxref_11_M2_noxref_s ) capacitor c=0.00290153f \
 //x=3.85 //y=1.26 //x2=2.965 //y2=0.375
cc_666 ( N_noxref_3_c_584_n N_D_c_2167_n ) capacitor c=0.0127164f //x=6.835 \
 //y=5.2 //x2=6.66 //y2=4.535
cc_667 ( N_noxref_3_c_568_n N_D_c_2167_n ) capacitor c=0.0101284f //x=7.4 \
 //y=3.33 //x2=6.66 //y2=4.535
cc_668 ( N_noxref_3_c_555_n N_D_c_2158_n ) capacitor c=0.0222863f //x=7.285 \
 //y=3.33 //x2=6.66 //y2=2.08
cc_669 ( N_noxref_3_c_565_n N_D_c_2158_n ) capacitor c=0.00117715f //x=7.515 \
 //y=3.33 //x2=6.66 //y2=2.08
cc_670 ( N_noxref_3_c_568_n N_D_c_2158_n ) capacitor c=0.0730419f //x=7.4 \
 //y=3.33 //x2=6.66 //y2=2.08
cc_671 ( N_noxref_3_c_569_n N_D_c_2158_n ) capacitor c=7.76771e-19 //x=9.25 \
 //y=2.08 //x2=6.66 //y2=2.08
cc_672 ( N_noxref_3_c_584_n N_D_M21_noxref_g ) capacitor c=0.0166421f \
 //x=6.835 //y=5.2 //x2=6.7 //y2=6.02
cc_673 ( N_noxref_3_M21_noxref_d N_D_M21_noxref_g ) capacitor c=0.0173476f \
 //x=6.775 //y=5.02 //x2=6.7 //y2=6.02
cc_674 ( N_noxref_3_c_590_n N_D_M22_noxref_g ) capacitor c=0.018922f //x=7.315 \
 //y=5.2 //x2=7.14 //y2=6.02
cc_675 ( N_noxref_3_M21_noxref_d N_D_M22_noxref_g ) capacitor c=0.0179769f \
 //x=6.775 //y=5.02 //x2=7.14 //y2=6.02
cc_676 ( N_noxref_3_M4_noxref_d N_D_c_2177_n ) capacitor c=0.00217566f \
 //x=6.77 //y=0.905 //x2=6.695 //y2=0.905
cc_677 ( N_noxref_3_M4_noxref_d N_D_c_2178_n ) capacitor c=0.0034598f //x=6.77 \
 //y=0.905 //x2=6.695 //y2=1.25
cc_678 ( N_noxref_3_M4_noxref_d N_D_c_2179_n ) capacitor c=0.0065582f //x=6.77 \
 //y=0.905 //x2=6.695 //y2=1.56
cc_679 ( N_noxref_3_c_568_n N_D_c_2180_n ) capacitor c=0.0142673f //x=7.4 \
 //y=3.33 //x2=7.065 //y2=4.79
cc_680 ( N_noxref_3_c_751_p N_D_c_2180_n ) capacitor c=0.00407665f //x=6.92 \
 //y=5.2 //x2=7.065 //y2=4.79
cc_681 ( N_noxref_3_M4_noxref_d N_D_c_2182_n ) capacitor c=0.00241102f \
 //x=6.77 //y=0.905 //x2=7.07 //y2=0.75
cc_682 ( N_noxref_3_c_567_n N_D_c_2183_n ) capacitor c=0.00359704f //x=7.315 \
 //y=1.655 //x2=7.07 //y2=1.405
cc_683 ( N_noxref_3_M4_noxref_d N_D_c_2183_n ) capacitor c=0.0138845f //x=6.77 \
 //y=0.905 //x2=7.07 //y2=1.405
cc_684 ( N_noxref_3_M4_noxref_d N_D_c_2185_n ) capacitor c=0.00132245f \
 //x=6.77 //y=0.905 //x2=7.225 //y2=0.905
cc_685 ( N_noxref_3_c_567_n N_D_c_2186_n ) capacitor c=0.00457401f //x=7.315 \
 //y=1.655 //x2=7.225 //y2=1.25
cc_686 ( N_noxref_3_M4_noxref_d N_D_c_2186_n ) capacitor c=0.00566463f \
 //x=6.77 //y=0.905 //x2=7.225 //y2=1.25
cc_687 ( N_noxref_3_c_568_n N_D_c_2188_n ) capacitor c=0.00877984f //x=7.4 \
 //y=3.33 //x2=6.66 //y2=2.08
cc_688 ( N_noxref_3_c_568_n N_D_c_2189_n ) capacitor c=0.00306024f //x=7.4 \
 //y=3.33 //x2=6.66 //y2=1.915
cc_689 ( N_noxref_3_M4_noxref_d N_D_c_2189_n ) capacitor c=0.00660593f \
 //x=6.77 //y=0.905 //x2=6.66 //y2=1.915
cc_690 ( N_noxref_3_c_584_n N_D_c_2191_n ) capacitor c=0.00346527f //x=6.835 \
 //y=5.2 //x2=6.69 //y2=4.7
cc_691 ( N_noxref_3_c_568_n N_D_c_2191_n ) capacitor c=0.00533692f //x=7.4 \
 //y=3.33 //x2=6.69 //y2=4.7
cc_692 ( N_noxref_3_c_555_n N_noxref_13_c_2250_n ) capacitor c=0.00241565f \
 //x=7.285 //y=3.33 //x2=5.505 //y2=1.495
cc_693 ( N_noxref_3_c_764_p N_noxref_13_c_2250_n ) capacitor c=3.15806e-19 \
 //x=7.045 //y=1.655 //x2=5.505 //y2=1.495
cc_694 ( N_noxref_3_c_555_n N_noxref_13_c_2231_n ) capacitor c=0.010299f \
 //x=7.285 //y=3.33 //x2=6.39 //y2=1.58
cc_695 ( N_noxref_3_c_555_n N_noxref_13_c_2238_n ) capacitor c=0.00241565f \
 //x=7.285 //y=3.33 //x2=6.475 //y2=1.495
cc_696 ( N_noxref_3_c_764_p N_noxref_13_c_2238_n ) capacitor c=0.020324f \
 //x=7.045 //y=1.655 //x2=6.475 //y2=1.495
cc_697 ( N_noxref_3_c_555_n N_noxref_13_c_2239_n ) capacitor c=7.52304e-19 \
 //x=7.285 //y=3.33 //x2=7.36 //y2=0.53
cc_698 ( N_noxref_3_c_567_n N_noxref_13_c_2239_n ) capacitor c=0.00465965f \
 //x=7.315 //y=1.655 //x2=7.36 //y2=0.53
cc_699 ( N_noxref_3_M4_noxref_d N_noxref_13_c_2239_n ) capacitor c=0.0117692f \
 //x=6.77 //y=0.905 //x2=7.36 //y2=0.53
cc_700 ( N_noxref_3_c_565_n N_noxref_13_M3_noxref_s ) capacitor c=3.47564e-19 \
 //x=7.515 //y=3.33 //x2=5.37 //y2=0.365
cc_701 ( N_noxref_3_c_567_n N_noxref_13_M3_noxref_s ) capacitor c=0.0141735f \
 //x=7.315 //y=1.655 //x2=5.37 //y2=0.365
cc_702 ( N_noxref_3_M4_noxref_d N_noxref_13_M3_noxref_s ) capacitor \
 c=0.0439476f //x=6.77 //y=0.905 //x2=5.37 //y2=0.365
cc_703 ( N_noxref_3_c_561_n N_noxref_14_c_2302_n ) capacitor c=0.00241565f \
 //x=9.135 //y=3.33 //x2=8.835 //y2=1.495
cc_704 ( N_noxref_3_c_567_n N_noxref_14_c_2302_n ) capacitor c=3.22188e-19 \
 //x=7.315 //y=1.655 //x2=8.835 //y2=1.495
cc_705 ( N_noxref_3_c_574_n N_noxref_14_c_2302_n ) capacitor c=0.0034165f \
 //x=9.055 //y=1.915 //x2=8.835 //y2=1.495
cc_706 ( N_noxref_3_c_561_n N_noxref_14_c_2283_n ) capacitor c=0.00649414f \
 //x=9.135 //y=3.33 //x2=9.72 //y2=1.58
cc_707 ( N_noxref_3_c_569_n N_noxref_14_c_2283_n ) capacitor c=0.011692f \
 //x=9.25 //y=2.08 //x2=9.72 //y2=1.58
cc_708 ( N_noxref_3_c_573_n N_noxref_14_c_2283_n ) capacitor c=0.00703567f \
 //x=9.055 //y=1.52 //x2=9.72 //y2=1.58
cc_709 ( N_noxref_3_c_574_n N_noxref_14_c_2283_n ) capacitor c=0.0203514f \
 //x=9.055 //y=1.915 //x2=9.72 //y2=1.58
cc_710 ( N_noxref_3_c_576_n N_noxref_14_c_2283_n ) capacitor c=0.00780629f \
 //x=9.43 //y=1.365 //x2=9.72 //y2=1.58
cc_711 ( N_noxref_3_c_579_n N_noxref_14_c_2283_n ) capacitor c=0.00339872f \
 //x=9.585 //y=1.21 //x2=9.72 //y2=1.58
cc_712 ( N_noxref_3_c_574_n N_noxref_14_c_2290_n ) capacitor c=6.71402e-19 \
 //x=9.055 //y=1.915 //x2=9.805 //y2=1.495
cc_713 ( N_noxref_3_c_570_n N_noxref_14_M5_noxref_s ) capacitor c=0.0326577f \
 //x=9.055 //y=0.865 //x2=8.7 //y2=0.365
cc_714 ( N_noxref_3_c_573_n N_noxref_14_M5_noxref_s ) capacitor c=3.48408e-19 \
 //x=9.055 //y=1.52 //x2=8.7 //y2=0.365
cc_715 ( N_noxref_3_c_577_n N_noxref_14_M5_noxref_s ) capacitor c=0.0120759f \
 //x=9.585 //y=0.865 //x2=8.7 //y2=0.365
cc_716 ( N_noxref_4_c_808_n N_CLK_c_940_n ) capacitor c=0.0185297f //x=10.165 \
 //y=5.2 //x2=13.205 //y2=4.44
cc_717 ( N_noxref_4_c_812_n N_CLK_c_940_n ) capacitor c=0.018142f //x=9.455 \
 //y=5.2 //x2=13.205 //y2=4.44
cc_718 ( N_noxref_4_c_793_n N_CLK_c_940_n ) capacitor c=0.0208321f //x=10.73 \
 //y=3.33 //x2=13.205 //y2=4.44
cc_719 ( N_noxref_4_c_794_n N_CLK_c_940_n ) capacitor c=0.0215137f //x=12.58 \
 //y=2.08 //x2=13.205 //y2=4.44
cc_720 ( N_noxref_4_c_827_n N_CLK_c_940_n ) capacitor c=0.0109968f //x=12.58 \
 //y=4.7 //x2=13.205 //y2=4.44
cc_721 ( N_noxref_4_c_794_n N_CLK_c_1003_n ) capacitor c=0.00400249f //x=12.58 \
 //y=2.08 //x2=13.32 //y2=4.535
cc_722 ( N_noxref_4_c_827_n N_CLK_c_1003_n ) capacitor c=0.00415951f //x=12.58 \
 //y=4.7 //x2=13.32 //y2=4.535
cc_723 ( N_noxref_4_c_787_n N_CLK_c_938_n ) capacitor c=0.00720056f //x=12.465 \
 //y=3.33 //x2=13.32 //y2=2.08
cc_724 ( N_noxref_4_c_793_n N_CLK_c_938_n ) capacitor c=0.00102338f //x=10.73 \
 //y=3.33 //x2=13.32 //y2=2.08
cc_725 ( N_noxref_4_c_794_n N_CLK_c_938_n ) capacitor c=0.0785565f //x=12.58 \
 //y=2.08 //x2=13.32 //y2=2.08
cc_726 ( N_noxref_4_c_799_n N_CLK_c_938_n ) capacitor c=0.00308814f //x=12.385 \
 //y=1.915 //x2=13.32 //y2=2.08
cc_727 ( N_noxref_4_M27_noxref_g N_CLK_M29_noxref_g ) capacitor c=0.0104611f \
 //x=12.48 //y=6.02 //x2=13.36 //y2=6.02
cc_728 ( N_noxref_4_M28_noxref_g N_CLK_M29_noxref_g ) capacitor c=0.106811f \
 //x=12.92 //y=6.02 //x2=13.36 //y2=6.02
cc_729 ( N_noxref_4_M28_noxref_g N_CLK_M30_noxref_g ) capacitor c=0.0100341f \
 //x=12.92 //y=6.02 //x2=13.8 //y2=6.02
cc_730 ( N_noxref_4_c_795_n N_CLK_c_1012_n ) capacitor c=4.86506e-19 \
 //x=12.385 //y=0.865 //x2=13.355 //y2=0.905
cc_731 ( N_noxref_4_c_797_n N_CLK_c_1012_n ) capacitor c=0.00152104f \
 //x=12.385 //y=1.21 //x2=13.355 //y2=0.905
cc_732 ( N_noxref_4_c_802_n N_CLK_c_1012_n ) capacitor c=0.0151475f //x=12.915 \
 //y=0.865 //x2=13.355 //y2=0.905
cc_733 ( N_noxref_4_c_798_n N_CLK_c_1015_n ) capacitor c=0.00109982f \
 //x=12.385 //y=1.52 //x2=13.355 //y2=1.25
cc_734 ( N_noxref_4_c_804_n N_CLK_c_1015_n ) capacitor c=0.0111064f //x=12.915 \
 //y=1.21 //x2=13.355 //y2=1.25
cc_735 ( N_noxref_4_c_798_n N_CLK_c_1017_n ) capacitor c=9.57794e-19 \
 //x=12.385 //y=1.52 //x2=13.355 //y2=1.56
cc_736 ( N_noxref_4_c_799_n N_CLK_c_1017_n ) capacitor c=0.00662747f \
 //x=12.385 //y=1.915 //x2=13.355 //y2=1.56
cc_737 ( N_noxref_4_c_804_n N_CLK_c_1017_n ) capacitor c=0.00862358f \
 //x=12.915 //y=1.21 //x2=13.355 //y2=1.56
cc_738 ( N_noxref_4_c_802_n N_CLK_c_1020_n ) capacitor c=0.00124821f \
 //x=12.915 //y=0.865 //x2=13.885 //y2=0.905
cc_739 ( N_noxref_4_c_804_n N_CLK_c_1021_n ) capacitor c=0.00200715f \
 //x=12.915 //y=1.21 //x2=13.885 //y2=1.25
cc_740 ( N_noxref_4_c_794_n N_CLK_c_1022_n ) capacitor c=0.00307062f //x=12.58 \
 //y=2.08 //x2=13.32 //y2=2.08
cc_741 ( N_noxref_4_c_799_n N_CLK_c_1022_n ) capacitor c=0.0179092f //x=12.385 \
 //y=1.915 //x2=13.32 //y2=2.08
cc_742 ( N_noxref_4_c_794_n N_CLK_c_1024_n ) capacitor c=0.00342116f //x=12.58 \
 //y=2.08 //x2=13.35 //y2=4.7
cc_743 ( N_noxref_4_c_827_n N_CLK_c_1024_n ) capacitor c=0.0292158f //x=12.58 \
 //y=4.7 //x2=13.35 //y2=4.7
cc_744 ( N_noxref_4_c_787_n N_noxref_6_c_1142_n ) capacitor c=0.175696f \
 //x=12.465 //y=3.33 //x2=15.795 //y2=3.7
cc_745 ( N_noxref_4_c_791_n N_noxref_6_c_1142_n ) capacitor c=0.0293967f \
 //x=10.845 //y=3.33 //x2=15.795 //y2=3.7
cc_746 ( N_noxref_4_c_877_p N_noxref_6_c_1142_n ) capacitor c=0.0037701f \
 //x=10.375 //y=1.655 //x2=15.795 //y2=3.7
cc_747 ( N_noxref_4_c_793_n N_noxref_6_c_1142_n ) capacitor c=0.0206034f \
 //x=10.73 //y=3.33 //x2=15.795 //y2=3.7
cc_748 ( N_noxref_4_c_794_n N_noxref_6_c_1142_n ) capacitor c=0.0205831f \
 //x=12.58 //y=2.08 //x2=15.795 //y2=3.7
cc_749 ( N_noxref_4_c_787_n N_noxref_8_c_1572_n ) capacitor c=0.0110241f \
 //x=12.465 //y=3.33 //x2=13.945 //y2=4.07
cc_750 ( N_noxref_4_c_791_n N_noxref_8_c_1572_n ) capacitor c=8.88358e-19 \
 //x=10.845 //y=3.33 //x2=13.945 //y2=4.07
cc_751 ( N_noxref_4_c_793_n N_noxref_8_c_1572_n ) capacitor c=0.0181936f \
 //x=10.73 //y=3.33 //x2=13.945 //y2=4.07
cc_752 ( N_noxref_4_c_794_n N_noxref_8_c_1572_n ) capacitor c=0.0184765f \
 //x=12.58 //y=2.08 //x2=13.945 //y2=4.07
cc_753 ( N_noxref_4_c_793_n N_noxref_8_c_1642_n ) capacitor c=0.00117715f \
 //x=10.73 //y=3.33 //x2=10.105 //y2=4.07
cc_754 ( N_noxref_4_c_808_n N_noxref_8_c_1644_n ) capacitor c=0.0127164f \
 //x=10.165 //y=5.2 //x2=9.99 //y2=4.535
cc_755 ( N_noxref_4_c_793_n N_noxref_8_c_1644_n ) capacitor c=0.0101319f \
 //x=10.73 //y=3.33 //x2=9.99 //y2=4.535
cc_756 ( N_noxref_4_c_791_n N_noxref_8_c_1546_n ) capacitor c=0.00329059f \
 //x=10.845 //y=3.33 //x2=9.99 //y2=2.08
cc_757 ( N_noxref_4_c_793_n N_noxref_8_c_1546_n ) capacitor c=0.0742673f \
 //x=10.73 //y=3.33 //x2=9.99 //y2=2.08
cc_758 ( N_noxref_4_c_794_n N_noxref_8_c_1546_n ) capacitor c=9.69022e-19 \
 //x=12.58 //y=2.08 //x2=9.99 //y2=2.08
cc_759 ( N_noxref_4_M28_noxref_g N_noxref_8_c_1594_n ) capacitor c=0.0169521f \
 //x=12.92 //y=6.02 //x2=13.495 //y2=5.2
cc_760 ( N_noxref_4_c_794_n N_noxref_8_c_1598_n ) capacitor c=0.00539951f \
 //x=12.58 //y=2.08 //x2=12.785 //y2=5.2
cc_761 ( N_noxref_4_M27_noxref_g N_noxref_8_c_1598_n ) capacitor c=0.0177326f \
 //x=12.48 //y=6.02 //x2=12.785 //y2=5.2
cc_762 ( N_noxref_4_c_827_n N_noxref_8_c_1598_n ) capacitor c=0.00581252f \
 //x=12.58 //y=4.7 //x2=12.785 //y2=5.2
cc_763 ( N_noxref_4_c_793_n N_noxref_8_c_1549_n ) capacitor c=3.49822e-19 \
 //x=10.73 //y=3.33 //x2=14.06 //y2=4.07
cc_764 ( N_noxref_4_c_794_n N_noxref_8_c_1549_n ) capacitor c=0.00389543f \
 //x=12.58 //y=2.08 //x2=14.06 //y2=4.07
cc_765 ( N_noxref_4_c_808_n N_noxref_8_M25_noxref_g ) capacitor c=0.0166421f \
 //x=10.165 //y=5.2 //x2=10.03 //y2=6.02
cc_766 ( N_noxref_4_M25_noxref_d N_noxref_8_M25_noxref_g ) capacitor \
 c=0.0173476f //x=10.105 //y=5.02 //x2=10.03 //y2=6.02
cc_767 ( N_noxref_4_c_814_n N_noxref_8_M26_noxref_g ) capacitor c=0.018922f \
 //x=10.645 //y=5.2 //x2=10.47 //y2=6.02
cc_768 ( N_noxref_4_M25_noxref_d N_noxref_8_M26_noxref_g ) capacitor \
 c=0.0179769f //x=10.105 //y=5.02 //x2=10.47 //y2=6.02
cc_769 ( N_noxref_4_M6_noxref_d N_noxref_8_c_1653_n ) capacitor c=0.00217566f \
 //x=10.1 //y=0.905 //x2=10.025 //y2=0.905
cc_770 ( N_noxref_4_M6_noxref_d N_noxref_8_c_1656_n ) capacitor c=0.0034598f \
 //x=10.1 //y=0.905 //x2=10.025 //y2=1.25
cc_771 ( N_noxref_4_M6_noxref_d N_noxref_8_c_1658_n ) capacitor c=0.0065582f \
 //x=10.1 //y=0.905 //x2=10.025 //y2=1.56
cc_772 ( N_noxref_4_c_793_n N_noxref_8_c_1690_n ) capacitor c=0.0142673f \
 //x=10.73 //y=3.33 //x2=10.395 //y2=4.79
cc_773 ( N_noxref_4_c_904_p N_noxref_8_c_1690_n ) capacitor c=0.00407665f \
 //x=10.25 //y=5.2 //x2=10.395 //y2=4.79
cc_774 ( N_noxref_4_M6_noxref_d N_noxref_8_c_1692_n ) capacitor c=0.00241102f \
 //x=10.1 //y=0.905 //x2=10.4 //y2=0.75
cc_775 ( N_noxref_4_c_792_n N_noxref_8_c_1693_n ) capacitor c=0.00359704f \
 //x=10.645 //y=1.655 //x2=10.4 //y2=1.405
cc_776 ( N_noxref_4_M6_noxref_d N_noxref_8_c_1693_n ) capacitor c=0.0138845f \
 //x=10.1 //y=0.905 //x2=10.4 //y2=1.405
cc_777 ( N_noxref_4_M6_noxref_d N_noxref_8_c_1661_n ) capacitor c=0.00132245f \
 //x=10.1 //y=0.905 //x2=10.555 //y2=0.905
cc_778 ( N_noxref_4_c_792_n N_noxref_8_c_1662_n ) capacitor c=0.00457401f \
 //x=10.645 //y=1.655 //x2=10.555 //y2=1.25
cc_779 ( N_noxref_4_M6_noxref_d N_noxref_8_c_1662_n ) capacitor c=0.00566463f \
 //x=10.1 //y=0.905 //x2=10.555 //y2=1.25
cc_780 ( N_noxref_4_c_793_n N_noxref_8_c_1663_n ) capacitor c=0.00877984f \
 //x=10.73 //y=3.33 //x2=9.99 //y2=2.08
cc_781 ( N_noxref_4_c_793_n N_noxref_8_c_1699_n ) capacitor c=0.00306024f \
 //x=10.73 //y=3.33 //x2=9.99 //y2=1.915
cc_782 ( N_noxref_4_M6_noxref_d N_noxref_8_c_1699_n ) capacitor c=0.00660593f \
 //x=10.1 //y=0.905 //x2=9.99 //y2=1.915
cc_783 ( N_noxref_4_c_808_n N_noxref_8_c_1665_n ) capacitor c=0.00346527f \
 //x=10.165 //y=5.2 //x2=10.02 //y2=4.7
cc_784 ( N_noxref_4_c_793_n N_noxref_8_c_1665_n ) capacitor c=0.00517969f \
 //x=10.73 //y=3.33 //x2=10.02 //y2=4.7
cc_785 ( N_noxref_4_M28_noxref_g N_noxref_8_M27_noxref_d ) capacitor \
 c=0.0173476f //x=12.92 //y=6.02 //x2=12.555 //y2=5.02
cc_786 ( N_noxref_4_c_877_p N_noxref_14_c_2302_n ) capacitor c=3.15806e-19 \
 //x=10.375 //y=1.655 //x2=8.835 //y2=1.495
cc_787 ( N_noxref_4_c_877_p N_noxref_14_c_2290_n ) capacitor c=0.0203424f \
 //x=10.375 //y=1.655 //x2=9.805 //y2=1.495
cc_788 ( N_noxref_4_c_792_n N_noxref_14_c_2291_n ) capacitor c=0.0046686f \
 //x=10.645 //y=1.655 //x2=10.69 //y2=0.53
cc_789 ( N_noxref_4_M6_noxref_d N_noxref_14_c_2291_n ) capacitor c=0.0117932f \
 //x=10.1 //y=0.905 //x2=10.69 //y2=0.53
cc_790 ( N_noxref_4_c_791_n N_noxref_14_M5_noxref_s ) capacitor c=3.47564e-19 \
 //x=10.845 //y=3.33 //x2=8.7 //y2=0.365
cc_791 ( N_noxref_4_c_792_n N_noxref_14_M5_noxref_s ) capacitor c=0.0141735f \
 //x=10.645 //y=1.655 //x2=8.7 //y2=0.365
cc_792 ( N_noxref_4_M6_noxref_d N_noxref_14_M5_noxref_s ) capacitor \
 c=0.043966f //x=10.1 //y=0.905 //x2=8.7 //y2=0.365
cc_793 ( N_noxref_4_c_787_n N_noxref_15_c_2355_n ) capacitor c=0.00241565f \
 //x=12.465 //y=3.33 //x2=12.165 //y2=1.495
cc_794 ( N_noxref_4_c_792_n N_noxref_15_c_2355_n ) capacitor c=3.22188e-19 \
 //x=10.645 //y=1.655 //x2=12.165 //y2=1.495
cc_795 ( N_noxref_4_c_799_n N_noxref_15_c_2355_n ) capacitor c=0.0034165f \
 //x=12.385 //y=1.915 //x2=12.165 //y2=1.495
cc_796 ( N_noxref_4_c_787_n N_noxref_15_c_2336_n ) capacitor c=0.00649414f \
 //x=12.465 //y=3.33 //x2=13.05 //y2=1.58
cc_797 ( N_noxref_4_c_794_n N_noxref_15_c_2336_n ) capacitor c=0.011692f \
 //x=12.58 //y=2.08 //x2=13.05 //y2=1.58
cc_798 ( N_noxref_4_c_798_n N_noxref_15_c_2336_n ) capacitor c=0.00703567f \
 //x=12.385 //y=1.52 //x2=13.05 //y2=1.58
cc_799 ( N_noxref_4_c_799_n N_noxref_15_c_2336_n ) capacitor c=0.0203514f \
 //x=12.385 //y=1.915 //x2=13.05 //y2=1.58
cc_800 ( N_noxref_4_c_801_n N_noxref_15_c_2336_n ) capacitor c=0.00780629f \
 //x=12.76 //y=1.365 //x2=13.05 //y2=1.58
cc_801 ( N_noxref_4_c_804_n N_noxref_15_c_2336_n ) capacitor c=0.00339872f \
 //x=12.915 //y=1.21 //x2=13.05 //y2=1.58
cc_802 ( N_noxref_4_c_799_n N_noxref_15_c_2343_n ) capacitor c=6.71402e-19 \
 //x=12.385 //y=1.915 //x2=13.135 //y2=1.495
cc_803 ( N_noxref_4_c_795_n N_noxref_15_M7_noxref_s ) capacitor c=0.0326577f \
 //x=12.385 //y=0.865 //x2=12.03 //y2=0.365
cc_804 ( N_noxref_4_c_798_n N_noxref_15_M7_noxref_s ) capacitor c=3.48408e-19 \
 //x=12.385 //y=1.52 //x2=12.03 //y2=0.365
cc_805 ( N_noxref_4_c_802_n N_noxref_15_M7_noxref_s ) capacitor c=0.0120759f \
 //x=12.915 //y=0.865 //x2=12.03 //y2=0.365
cc_806 ( N_CLK_c_940_n N_noxref_6_c_1215_n ) capacitor c=0.00940379f \
 //x=13.205 //y=4.44 //x2=5.805 //y2=3.7
cc_807 ( N_CLK_c_940_n N_noxref_6_c_1216_n ) capacitor c=7.95009e-19 \
 //x=13.205 //y=4.44 //x2=4.185 //y2=3.7
cc_808 ( N_CLK_c_940_n N_noxref_6_c_1142_n ) capacitor c=0.0492712f //x=13.205 \
 //y=4.44 //x2=15.795 //y2=3.7
cc_809 ( N_CLK_c_938_n N_noxref_6_c_1142_n ) capacitor c=0.0225527f //x=13.32 \
 //y=2.08 //x2=15.795 //y2=3.7
cc_810 ( N_CLK_c_940_n N_noxref_6_c_1223_n ) capacitor c=6.59192e-19 \
 //x=13.205 //y=4.44 //x2=6.035 //y2=3.7
cc_811 ( N_CLK_c_958_n N_noxref_6_c_1169_n ) capacitor c=0.00330099f //x=2.335 \
 //y=4.44 //x2=2.325 //y2=5.155
cc_812 ( N_CLK_c_937_n N_noxref_6_c_1169_n ) capacitor c=0.014564f //x=2.22 \
 //y=2.08 //x2=2.325 //y2=5.155
cc_813 ( N_CLK_M15_noxref_g N_noxref_6_c_1169_n ) capacitor c=0.016514f \
 //x=2.19 //y=6.02 //x2=2.325 //y2=5.155
cc_814 ( N_CLK_c_996_n N_noxref_6_c_1169_n ) capacitor c=0.00322046f //x=2.22 \
 //y=4.7 //x2=2.325 //y2=5.155
cc_815 ( N_CLK_M16_noxref_g N_noxref_6_c_1175_n ) capacitor c=0.01736f \
 //x=2.63 //y=6.02 //x2=3.205 //y2=5.155
cc_816 ( N_CLK_c_940_n N_noxref_6_c_1179_n ) capacitor c=0.0183122f //x=13.205 \
 //y=4.44 //x2=3.985 //y2=5.155
cc_817 ( N_CLK_c_940_n N_noxref_6_c_1183_n ) capacitor c=0.0210274f //x=13.205 \
 //y=4.44 //x2=4.07 //y2=3.7
cc_818 ( N_CLK_c_937_n N_noxref_6_c_1183_n ) capacitor c=0.00319363f //x=2.22 \
 //y=2.08 //x2=4.07 //y2=3.7
cc_819 ( N_CLK_c_940_n N_noxref_6_c_1145_n ) capacitor c=0.0198304f //x=13.205 \
 //y=4.44 //x2=5.92 //y2=2.08
cc_820 ( N_CLK_c_938_n N_noxref_6_c_1146_n ) capacitor c=0.00101176f //x=13.32 \
 //y=2.08 //x2=15.91 //y2=2.08
cc_821 ( N_CLK_c_940_n N_noxref_6_c_1277_n ) capacitor c=0.0311227f //x=13.205 \
 //y=4.44 //x2=2.41 //y2=5.155
cc_822 ( N_CLK_c_995_n N_noxref_6_c_1277_n ) capacitor c=0.00426767f //x=2.555 \
 //y=4.79 //x2=2.41 //y2=5.155
cc_823 ( N_CLK_c_940_n N_noxref_6_c_1198_n ) capacitor c=0.0107057f //x=13.205 \
 //y=4.44 //x2=5.92 //y2=4.7
cc_824 ( N_CLK_M15_noxref_g N_noxref_6_M15_noxref_d ) capacitor c=0.0180032f \
 //x=2.19 //y=6.02 //x2=2.265 //y2=5.02
cc_825 ( N_CLK_M16_noxref_g N_noxref_6_M15_noxref_d ) capacitor c=0.0180032f \
 //x=2.63 //y=6.02 //x2=2.265 //y2=5.02
cc_826 ( N_CLK_c_940_n N_noxref_8_c_1542_n ) capacitor c=0.656956f //x=13.205 \
 //y=4.44 //x2=9.875 //y2=4.07
cc_827 ( N_CLK_c_958_n N_noxref_8_c_1542_n ) capacitor c=0.0291328f //x=2.335 \
 //y=4.44 //x2=9.875 //y2=4.07
cc_828 ( N_CLK_c_937_n N_noxref_8_c_1542_n ) capacitor c=0.0265867f //x=2.22 \
 //y=2.08 //x2=9.875 //y2=4.07
cc_829 ( N_CLK_c_996_n N_noxref_8_c_1542_n ) capacitor c=6.38735e-19 //x=2.22 \
 //y=4.7 //x2=9.875 //y2=4.07
cc_830 ( N_CLK_c_937_n N_noxref_8_c_1543_n ) capacitor c=0.00128547f //x=2.22 \
 //y=2.08 //x2=1.225 //y2=4.07
cc_831 ( N_CLK_c_940_n N_noxref_8_c_1572_n ) capacitor c=0.300301f //x=13.205 \
 //y=4.44 //x2=13.945 //y2=4.07
cc_832 ( N_CLK_c_938_n N_noxref_8_c_1572_n ) capacitor c=0.0187718f //x=13.32 \
 //y=2.08 //x2=13.945 //y2=4.07
cc_833 ( N_CLK_c_1053_p N_noxref_8_c_1572_n ) capacitor c=0.00756255f \
 //x=13.725 //y=4.79 //x2=13.945 //y2=4.07
cc_834 ( N_CLK_c_1024_n N_noxref_8_c_1572_n ) capacitor c=4.6185e-19 //x=13.35 \
 //y=4.7 //x2=13.945 //y2=4.07
cc_835 ( N_CLK_c_940_n N_noxref_8_c_1642_n ) capacitor c=0.0263375f //x=13.205 \
 //y=4.44 //x2=10.105 //y2=4.07
cc_836 ( N_CLK_c_938_n N_noxref_8_c_1586_n ) capacitor c=0.00117715f //x=13.32 \
 //y=2.08 //x2=14.175 //y2=4.07
cc_837 ( N_CLK_c_958_n N_noxref_8_c_1545_n ) capacitor c=0.00551083f //x=2.335 \
 //y=4.44 //x2=1.11 //y2=2.08
cc_838 ( N_CLK_c_937_n N_noxref_8_c_1545_n ) capacitor c=0.0535714f //x=2.22 \
 //y=2.08 //x2=1.11 //y2=2.08
cc_839 ( N_CLK_c_992_n N_noxref_8_c_1545_n ) capacitor c=0.00231304f //x=2.31 \
 //y=1.915 //x2=1.11 //y2=2.08
cc_840 ( N_CLK_c_996_n N_noxref_8_c_1545_n ) capacitor c=0.00183762f //x=2.22 \
 //y=4.7 //x2=1.11 //y2=2.08
cc_841 ( N_CLK_c_940_n N_noxref_8_c_1644_n ) capacitor c=0.0016972f //x=13.205 \
 //y=4.44 //x2=9.99 //y2=4.535
cc_842 ( N_CLK_c_940_n N_noxref_8_c_1546_n ) capacitor c=0.0207534f //x=13.205 \
 //y=4.44 //x2=9.99 //y2=2.08
cc_843 ( N_CLK_c_940_n N_noxref_8_c_1594_n ) capacitor c=0.00325337f \
 //x=13.205 //y=4.44 //x2=13.495 //y2=5.2
cc_844 ( N_CLK_c_1003_n N_noxref_8_c_1594_n ) capacitor c=0.0126974f //x=13.32 \
 //y=4.535 //x2=13.495 //y2=5.2
cc_845 ( N_CLK_c_938_n N_noxref_8_c_1594_n ) capacitor c=3.74769e-19 //x=13.32 \
 //y=2.08 //x2=13.495 //y2=5.2
cc_846 ( N_CLK_M29_noxref_g N_noxref_8_c_1594_n ) capacitor c=0.0166421f \
 //x=13.36 //y=6.02 //x2=13.495 //y2=5.2
cc_847 ( N_CLK_c_1024_n N_noxref_8_c_1594_n ) capacitor c=0.00346519f \
 //x=13.35 //y=4.7 //x2=13.495 //y2=5.2
cc_848 ( N_CLK_c_940_n N_noxref_8_c_1598_n ) capacitor c=0.0172877f //x=13.205 \
 //y=4.44 //x2=12.785 //y2=5.2
cc_849 ( N_CLK_M30_noxref_g N_noxref_8_c_1600_n ) capacitor c=0.0199348f \
 //x=13.8 //y=6.02 //x2=13.975 //y2=5.2
cc_850 ( N_CLK_c_1070_p N_noxref_8_c_1548_n ) capacitor c=0.00359704f \
 //x=13.73 //y=1.405 //x2=13.975 //y2=1.655
cc_851 ( N_CLK_c_1021_n N_noxref_8_c_1548_n ) capacitor c=0.00457401f \
 //x=13.885 //y=1.25 //x2=13.975 //y2=1.655
cc_852 ( N_CLK_c_940_n N_noxref_8_c_1549_n ) capacitor c=0.00707546f \
 //x=13.205 //y=4.44 //x2=14.06 //y2=4.07
cc_853 ( N_CLK_c_1003_n N_noxref_8_c_1549_n ) capacitor c=0.00923416f \
 //x=13.32 //y=4.535 //x2=14.06 //y2=4.07
cc_854 ( N_CLK_c_938_n N_noxref_8_c_1549_n ) capacitor c=0.0757812f //x=13.32 \
 //y=2.08 //x2=14.06 //y2=4.07
cc_855 ( N_CLK_c_1053_p N_noxref_8_c_1549_n ) capacitor c=0.0142673f \
 //x=13.725 //y=4.79 //x2=14.06 //y2=4.07
cc_856 ( N_CLK_c_1022_n N_noxref_8_c_1549_n ) capacitor c=0.00877984f \
 //x=13.32 //y=2.08 //x2=14.06 //y2=4.07
cc_857 ( N_CLK_c_1077_p N_noxref_8_c_1549_n ) capacitor c=0.00306024f \
 //x=13.32 //y=1.915 //x2=14.06 //y2=4.07
cc_858 ( N_CLK_c_1024_n N_noxref_8_c_1549_n ) capacitor c=0.00518077f \
 //x=13.35 //y=4.7 //x2=14.06 //y2=4.07
cc_859 ( N_CLK_c_1053_p N_noxref_8_c_1737_n ) capacitor c=0.00408717f \
 //x=13.725 //y=4.79 //x2=13.58 //y2=5.2
cc_860 ( N_CLK_M15_noxref_g N_noxref_8_M13_noxref_g ) capacitor c=0.0105869f \
 //x=2.19 //y=6.02 //x2=1.31 //y2=6.02
cc_861 ( N_CLK_M15_noxref_g N_noxref_8_M14_noxref_g ) capacitor c=0.10632f \
 //x=2.19 //y=6.02 //x2=1.75 //y2=6.02
cc_862 ( N_CLK_M16_noxref_g N_noxref_8_M14_noxref_g ) capacitor c=0.0101598f \
 //x=2.63 //y=6.02 //x2=1.75 //y2=6.02
cc_863 ( N_CLK_c_1083_p N_noxref_8_c_1552_n ) capacitor c=5.72482e-19 \
 //x=1.785 //y=0.91 //x2=0.81 //y2=0.875
cc_864 ( N_CLK_c_1083_p N_noxref_8_c_1554_n ) capacitor c=0.00149976f \
 //x=1.785 //y=0.91 //x2=0.81 //y2=1.22
cc_865 ( N_CLK_c_1085_p N_noxref_8_c_1555_n ) capacitor c=0.00111227f \
 //x=1.785 //y=1.22 //x2=0.81 //y2=1.53
cc_866 ( N_CLK_c_937_n N_noxref_8_c_1556_n ) capacitor c=0.00238338f //x=2.22 \
 //y=2.08 //x2=0.81 //y2=1.915
cc_867 ( N_CLK_c_992_n N_noxref_8_c_1556_n ) capacitor c=0.00964411f //x=2.31 \
 //y=1.915 //x2=0.81 //y2=1.915
cc_868 ( N_CLK_c_1083_p N_noxref_8_c_1559_n ) capacitor c=0.0160123f //x=1.785 \
 //y=0.91 //x2=1.34 //y2=0.875
cc_869 ( N_CLK_c_989_n N_noxref_8_c_1559_n ) capacitor c=0.00103227f //x=2.31 \
 //y=0.91 //x2=1.34 //y2=0.875
cc_870 ( N_CLK_c_1085_p N_noxref_8_c_1561_n ) capacitor c=0.0124075f //x=1.785 \
 //y=1.22 //x2=1.34 //y2=1.22
cc_871 ( N_CLK_c_990_n N_noxref_8_c_1561_n ) capacitor c=0.0010154f //x=2.31 \
 //y=1.22 //x2=1.34 //y2=1.22
cc_872 ( N_CLK_c_991_n N_noxref_8_c_1561_n ) capacitor c=9.23422e-19 //x=2.31 \
 //y=1.45 //x2=1.34 //y2=1.22
cc_873 ( N_CLK_c_937_n N_noxref_8_c_1751_n ) capacitor c=0.00147352f //x=2.22 \
 //y=2.08 //x2=1.675 //y2=4.79
cc_874 ( N_CLK_c_996_n N_noxref_8_c_1751_n ) capacitor c=0.0168581f //x=2.22 \
 //y=4.7 //x2=1.675 //y2=4.79
cc_875 ( N_CLK_c_937_n N_noxref_8_c_1622_n ) capacitor c=0.00141297f //x=2.22 \
 //y=2.08 //x2=1.385 //y2=4.79
cc_876 ( N_CLK_c_996_n N_noxref_8_c_1622_n ) capacitor c=0.00484466f //x=2.22 \
 //y=4.7 //x2=1.385 //y2=4.79
cc_877 ( N_CLK_c_940_n N_noxref_8_c_1690_n ) capacitor c=0.00960248f \
 //x=13.205 //y=4.44 //x2=10.395 //y2=4.79
cc_878 ( N_CLK_c_940_n N_noxref_8_c_1665_n ) capacitor c=0.00203982f \
 //x=13.205 //y=4.44 //x2=10.02 //y2=4.7
cc_879 ( N_CLK_c_1012_n N_noxref_8_M8_noxref_d ) capacitor c=0.00217566f \
 //x=13.355 //y=0.905 //x2=13.43 //y2=0.905
cc_880 ( N_CLK_c_1015_n N_noxref_8_M8_noxref_d ) capacitor c=0.0034598f \
 //x=13.355 //y=1.25 //x2=13.43 //y2=0.905
cc_881 ( N_CLK_c_1017_n N_noxref_8_M8_noxref_d ) capacitor c=0.0065582f \
 //x=13.355 //y=1.56 //x2=13.43 //y2=0.905
cc_882 ( N_CLK_c_1102_p N_noxref_8_M8_noxref_d ) capacitor c=0.00241102f \
 //x=13.73 //y=0.75 //x2=13.43 //y2=0.905
cc_883 ( N_CLK_c_1070_p N_noxref_8_M8_noxref_d ) capacitor c=0.0138845f \
 //x=13.73 //y=1.405 //x2=13.43 //y2=0.905
cc_884 ( N_CLK_c_1020_n N_noxref_8_M8_noxref_d ) capacitor c=0.00132245f \
 //x=13.885 //y=0.905 //x2=13.43 //y2=0.905
cc_885 ( N_CLK_c_1021_n N_noxref_8_M8_noxref_d ) capacitor c=0.00566463f \
 //x=13.885 //y=1.25 //x2=13.43 //y2=0.905
cc_886 ( N_CLK_c_1077_p N_noxref_8_M8_noxref_d ) capacitor c=0.00660593f \
 //x=13.32 //y=1.915 //x2=13.43 //y2=0.905
cc_887 ( N_CLK_M29_noxref_g N_noxref_8_M29_noxref_d ) capacitor c=0.0173476f \
 //x=13.36 //y=6.02 //x2=13.435 //y2=5.02
cc_888 ( N_CLK_M30_noxref_g N_noxref_8_M29_noxref_d ) capacitor c=0.0179769f \
 //x=13.8 //y=6.02 //x2=13.435 //y2=5.02
cc_889 ( N_CLK_c_1083_p N_noxref_10_c_2065_n ) capacitor c=0.0167228f \
 //x=1.785 //y=0.91 //x2=2.445 //y2=0.54
cc_890 ( N_CLK_c_989_n N_noxref_10_c_2065_n ) capacitor c=0.00534519f //x=2.31 \
 //y=0.91 //x2=2.445 //y2=0.54
cc_891 ( N_CLK_c_937_n N_noxref_10_c_2076_n ) capacitor c=0.012357f //x=2.22 \
 //y=2.08 //x2=2.445 //y2=1.59
cc_892 ( N_CLK_c_1085_p N_noxref_10_c_2076_n ) capacitor c=0.0153476f \
 //x=1.785 //y=1.22 //x2=2.445 //y2=1.59
cc_893 ( N_CLK_c_992_n N_noxref_10_c_2076_n ) capacitor c=0.0230663f //x=2.31 \
 //y=1.915 //x2=2.445 //y2=1.59
cc_894 ( N_CLK_c_1083_p N_noxref_10_M0_noxref_s ) capacitor c=0.00798959f \
 //x=1.785 //y=0.91 //x2=0.455 //y2=0.375
cc_895 ( N_CLK_c_991_n N_noxref_10_M0_noxref_s ) capacitor c=0.00212176f \
 //x=2.31 //y=1.45 //x2=0.455 //y2=0.375
cc_896 ( N_CLK_c_992_n N_noxref_10_M0_noxref_s ) capacitor c=0.00298115f \
 //x=2.31 //y=1.915 //x2=0.455 //y2=0.375
cc_897 ( N_CLK_c_1117_p N_noxref_11_c_2105_n ) capacitor c=2.14837e-19 \
 //x=2.155 //y=0.755 //x2=3.015 //y2=0.995
cc_898 ( N_CLK_c_989_n N_noxref_11_c_2105_n ) capacitor c=0.00123426f //x=2.31 \
 //y=0.91 //x2=3.015 //y2=0.995
cc_899 ( N_CLK_c_990_n N_noxref_11_c_2105_n ) capacitor c=0.0129288f //x=2.31 \
 //y=1.22 //x2=3.015 //y2=0.995
cc_900 ( N_CLK_c_991_n N_noxref_11_c_2105_n ) capacitor c=0.00142359f //x=2.31 \
 //y=1.45 //x2=3.015 //y2=0.995
cc_901 ( N_CLK_c_1083_p N_noxref_11_M1_noxref_d ) capacitor c=0.00223875f \
 //x=1.785 //y=0.91 //x2=1.86 //y2=0.91
cc_902 ( N_CLK_c_1085_p N_noxref_11_M1_noxref_d ) capacitor c=0.00262485f \
 //x=1.785 //y=1.22 //x2=1.86 //y2=0.91
cc_903 ( N_CLK_c_1117_p N_noxref_11_M1_noxref_d ) capacitor c=0.00220746f \
 //x=2.155 //y=0.755 //x2=1.86 //y2=0.91
cc_904 ( N_CLK_c_1124_p N_noxref_11_M1_noxref_d ) capacitor c=0.00194798f \
 //x=2.155 //y=1.375 //x2=1.86 //y2=0.91
cc_905 ( N_CLK_c_989_n N_noxref_11_M1_noxref_d ) capacitor c=0.00198465f \
 //x=2.31 //y=0.91 //x2=1.86 //y2=0.91
cc_906 ( N_CLK_c_990_n N_noxref_11_M1_noxref_d ) capacitor c=0.00128384f \
 //x=2.31 //y=1.22 //x2=1.86 //y2=0.91
cc_907 ( N_CLK_c_989_n N_noxref_11_M2_noxref_s ) capacitor c=7.21316e-19 \
 //x=2.31 //y=0.91 //x2=2.965 //y2=0.375
cc_908 ( N_CLK_c_990_n N_noxref_11_M2_noxref_s ) capacitor c=0.00348171f \
 //x=2.31 //y=1.22 //x2=2.965 //y2=0.375
cc_909 ( N_CLK_c_940_n N_D_c_2167_n ) capacitor c=0.0016972f //x=13.205 \
 //y=4.44 //x2=6.66 //y2=4.535
cc_910 ( N_CLK_c_940_n N_D_c_2158_n ) capacitor c=0.0189188f //x=13.205 \
 //y=4.44 //x2=6.66 //y2=2.08
cc_911 ( N_CLK_c_940_n N_D_c_2180_n ) capacitor c=0.00960248f //x=13.205 \
 //y=4.44 //x2=7.065 //y2=4.79
cc_912 ( N_CLK_c_940_n N_D_c_2191_n ) capacitor c=0.00203982f //x=13.205 \
 //y=4.44 //x2=6.69 //y2=4.7
cc_913 ( N_CLK_c_1017_n N_noxref_15_c_2343_n ) capacitor c=0.00623646f \
 //x=13.355 //y=1.56 //x2=13.135 //y2=1.495
cc_914 ( N_CLK_c_1022_n N_noxref_15_c_2343_n ) capacitor c=0.00176439f \
 //x=13.32 //y=2.08 //x2=13.135 //y2=1.495
cc_915 ( N_CLK_c_938_n N_noxref_15_c_2344_n ) capacitor c=0.0016032f //x=13.32 \
 //y=2.08 //x2=14.02 //y2=0.53
cc_916 ( N_CLK_c_1012_n N_noxref_15_c_2344_n ) capacitor c=0.0188655f \
 //x=13.355 //y=0.905 //x2=14.02 //y2=0.53
cc_917 ( N_CLK_c_1020_n N_noxref_15_c_2344_n ) capacitor c=0.00656458f \
 //x=13.885 //y=0.905 //x2=14.02 //y2=0.53
cc_918 ( N_CLK_c_1022_n N_noxref_15_c_2344_n ) capacitor c=2.1838e-19 \
 //x=13.32 //y=2.08 //x2=14.02 //y2=0.53
cc_919 ( N_CLK_c_1012_n N_noxref_15_M7_noxref_s ) capacitor c=0.00623646f \
 //x=13.355 //y=0.905 //x2=12.03 //y2=0.365
cc_920 ( N_CLK_c_1020_n N_noxref_15_M7_noxref_s ) capacitor c=0.0143002f \
 //x=13.885 //y=0.905 //x2=12.03 //y2=0.365
cc_921 ( N_CLK_c_1021_n N_noxref_15_M7_noxref_s ) capacitor c=0.00290153f \
 //x=13.885 //y=1.25 //x2=12.03 //y2=0.365
cc_922 ( N_noxref_6_M32_noxref_g N_noxref_7_c_1416_n ) capacitor c=0.017965f \
 //x=16.25 //y=6.02 //x2=16.825 //y2=5.2
cc_923 ( N_noxref_6_c_1146_n N_noxref_7_c_1420_n ) capacitor c=0.00530485f \
 //x=15.91 //y=2.08 //x2=16.115 //y2=5.2
cc_924 ( N_noxref_6_M31_noxref_g N_noxref_7_c_1420_n ) capacitor c=0.0177326f \
 //x=15.81 //y=6.02 //x2=16.115 //y2=5.2
cc_925 ( N_noxref_6_c_1199_n N_noxref_7_c_1420_n ) capacitor c=0.00582246f \
 //x=15.91 //y=4.7 //x2=16.115 //y2=5.2
cc_926 ( N_noxref_6_c_1146_n N_noxref_7_c_1401_n ) capacitor c=0.00375655f \
 //x=15.91 //y=2.08 //x2=17.39 //y2=3.33
cc_927 ( N_noxref_6_M32_noxref_g N_noxref_7_M31_noxref_d ) capacitor \
 c=0.0173476f //x=16.25 //y=6.02 //x2=15.885 //y2=5.02
cc_928 ( N_noxref_6_c_1215_n N_noxref_8_c_1542_n ) capacitor c=0.147021f \
 //x=5.805 //y=3.7 //x2=9.875 //y2=4.07
cc_929 ( N_noxref_6_c_1216_n N_noxref_8_c_1542_n ) capacitor c=0.0294294f \
 //x=4.185 //y=3.7 //x2=9.875 //y2=4.07
cc_930 ( N_noxref_6_c_1142_n N_noxref_8_c_1542_n ) capacitor c=0.338937f \
 //x=15.795 //y=3.7 //x2=9.875 //y2=4.07
cc_931 ( N_noxref_6_c_1223_n N_noxref_8_c_1542_n ) capacitor c=0.0264478f \
 //x=6.035 //y=3.7 //x2=9.875 //y2=4.07
cc_932 ( N_noxref_6_c_1173_n N_noxref_8_c_1542_n ) capacitor c=0.0154449f \
 //x=1.615 //y=5.155 //x2=9.875 //y2=4.07
cc_933 ( N_noxref_6_c_1183_n N_noxref_8_c_1542_n ) capacitor c=0.0200328f \
 //x=4.07 //y=3.7 //x2=9.875 //y2=4.07
cc_934 ( N_noxref_6_c_1145_n N_noxref_8_c_1542_n ) capacitor c=0.0203111f \
 //x=5.92 //y=2.08 //x2=9.875 //y2=4.07
cc_935 ( N_noxref_6_c_1142_n N_noxref_8_c_1572_n ) capacitor c=0.339146f \
 //x=15.795 //y=3.7 //x2=13.945 //y2=4.07
cc_936 ( N_noxref_6_c_1142_n N_noxref_8_c_1642_n ) capacitor c=0.0267832f \
 //x=15.795 //y=3.7 //x2=10.105 //y2=4.07
cc_937 ( N_noxref_6_c_1142_n N_noxref_8_c_1544_n ) capacitor c=0.176049f \
 //x=15.795 //y=3.7 //x2=19.865 //y2=4.07
cc_938 ( N_noxref_6_c_1146_n N_noxref_8_c_1544_n ) capacitor c=0.0242341f \
 //x=15.91 //y=2.08 //x2=19.865 //y2=4.07
cc_939 ( N_noxref_6_c_1199_n N_noxref_8_c_1544_n ) capacitor c=0.00703556f \
 //x=15.91 //y=4.7 //x2=19.865 //y2=4.07
cc_940 ( N_noxref_6_c_1142_n N_noxref_8_c_1586_n ) capacitor c=0.0266833f \
 //x=15.795 //y=3.7 //x2=14.175 //y2=4.07
cc_941 ( N_noxref_6_c_1146_n N_noxref_8_c_1586_n ) capacitor c=3.50683e-19 \
 //x=15.91 //y=2.08 //x2=14.175 //y2=4.07
cc_942 ( N_noxref_6_c_1142_n N_noxref_8_c_1546_n ) capacitor c=0.0243898f \
 //x=15.795 //y=3.7 //x2=9.99 //y2=2.08
cc_943 ( N_noxref_6_c_1142_n N_noxref_8_c_1782_n ) capacitor c=0.00433945f \
 //x=15.795 //y=3.7 //x2=13.705 //y2=1.655
cc_944 ( N_noxref_6_c_1142_n N_noxref_8_c_1549_n ) capacitor c=0.0268509f \
 //x=15.795 //y=3.7 //x2=14.06 //y2=4.07
cc_945 ( N_noxref_6_c_1146_n N_noxref_8_c_1549_n ) capacitor c=0.0144279f \
 //x=15.91 //y=2.08 //x2=14.06 //y2=4.07
cc_946 ( N_noxref_6_c_1173_n N_noxref_8_M13_noxref_g ) capacitor c=0.0213876f \
 //x=1.615 //y=5.155 //x2=1.31 //y2=6.02
cc_947 ( N_noxref_6_c_1169_n N_noxref_8_M14_noxref_g ) capacitor c=0.0178794f \
 //x=2.325 //y=5.155 //x2=1.75 //y2=6.02
cc_948 ( N_noxref_6_M13_noxref_d N_noxref_8_M14_noxref_g ) capacitor \
 c=0.0180032f //x=1.385 //y=5.02 //x2=1.75 //y2=6.02
cc_949 ( N_noxref_6_c_1173_n N_noxref_8_c_1751_n ) capacitor c=0.00429591f \
 //x=1.615 //y=5.155 //x2=1.675 //y2=4.79
cc_950 ( N_noxref_6_c_1142_n N_Q_c_1901_n ) capacitor c=0.0244534f //x=15.795 \
 //y=3.7 //x2=16.765 //y2=3.7
cc_951 ( N_noxref_6_c_1146_n N_Q_c_1901_n ) capacitor c=0.00245879f //x=15.91 \
 //y=2.08 //x2=16.765 //y2=3.7
cc_952 ( N_noxref_6_c_1146_n N_Q_c_1941_n ) capacitor c=0.00400249f //x=15.91 \
 //y=2.08 //x2=16.65 //y2=4.535
cc_953 ( N_noxref_6_c_1199_n N_Q_c_1941_n ) capacitor c=0.00417994f //x=15.91 \
 //y=4.7 //x2=16.65 //y2=4.535
cc_954 ( N_noxref_6_c_1142_n N_Q_c_1903_n ) capacitor c=0.00246068f //x=15.795 \
 //y=3.7 //x2=16.65 //y2=2.08
cc_955 ( N_noxref_6_c_1146_n N_Q_c_1903_n ) capacitor c=0.0837791f //x=15.91 \
 //y=2.08 //x2=16.65 //y2=2.08
cc_956 ( N_noxref_6_c_1161_n N_Q_c_1903_n ) capacitor c=0.00308814f //x=15.715 \
 //y=1.915 //x2=16.65 //y2=2.08
cc_957 ( N_noxref_6_M31_noxref_g N_Q_M33_noxref_g ) capacitor c=0.0104611f \
 //x=15.81 //y=6.02 //x2=16.69 //y2=6.02
cc_958 ( N_noxref_6_M32_noxref_g N_Q_M33_noxref_g ) capacitor c=0.106811f \
 //x=16.25 //y=6.02 //x2=16.69 //y2=6.02
cc_959 ( N_noxref_6_M32_noxref_g N_Q_M34_noxref_g ) capacitor c=0.0100341f \
 //x=16.25 //y=6.02 //x2=17.13 //y2=6.02
cc_960 ( N_noxref_6_c_1157_n N_Q_c_1949_n ) capacitor c=4.86506e-19 //x=15.715 \
 //y=0.865 //x2=16.685 //y2=0.905
cc_961 ( N_noxref_6_c_1159_n N_Q_c_1949_n ) capacitor c=0.00152104f //x=15.715 \
 //y=1.21 //x2=16.685 //y2=0.905
cc_962 ( N_noxref_6_c_1164_n N_Q_c_1949_n ) capacitor c=0.0151475f //x=16.245 \
 //y=0.865 //x2=16.685 //y2=0.905
cc_963 ( N_noxref_6_c_1160_n N_Q_c_1952_n ) capacitor c=0.00109982f //x=15.715 \
 //y=1.52 //x2=16.685 //y2=1.25
cc_964 ( N_noxref_6_c_1166_n N_Q_c_1952_n ) capacitor c=0.0111064f //x=16.245 \
 //y=1.21 //x2=16.685 //y2=1.25
cc_965 ( N_noxref_6_c_1160_n N_Q_c_1954_n ) capacitor c=9.57794e-19 //x=15.715 \
 //y=1.52 //x2=16.685 //y2=1.56
cc_966 ( N_noxref_6_c_1161_n N_Q_c_1954_n ) capacitor c=0.00662747f //x=15.715 \
 //y=1.915 //x2=16.685 //y2=1.56
cc_967 ( N_noxref_6_c_1166_n N_Q_c_1954_n ) capacitor c=0.00862358f //x=16.245 \
 //y=1.21 //x2=16.685 //y2=1.56
cc_968 ( N_noxref_6_c_1164_n N_Q_c_1957_n ) capacitor c=0.00124821f //x=16.245 \
 //y=0.865 //x2=17.215 //y2=0.905
cc_969 ( N_noxref_6_c_1166_n N_Q_c_1958_n ) capacitor c=0.00200715f //x=16.245 \
 //y=1.21 //x2=17.215 //y2=1.25
cc_970 ( N_noxref_6_c_1146_n N_Q_c_1959_n ) capacitor c=0.00307062f //x=15.91 \
 //y=2.08 //x2=16.65 //y2=2.08
cc_971 ( N_noxref_6_c_1161_n N_Q_c_1959_n ) capacitor c=0.0179092f //x=15.715 \
 //y=1.915 //x2=16.65 //y2=2.08
cc_972 ( N_noxref_6_c_1146_n N_Q_c_1961_n ) capacitor c=0.00344981f //x=15.91 \
 //y=2.08 //x2=16.68 //y2=4.7
cc_973 ( N_noxref_6_c_1199_n N_Q_c_1961_n ) capacitor c=0.0293367f //x=15.91 \
 //y=4.7 //x2=16.68 //y2=4.7
cc_974 ( N_noxref_6_M2_noxref_d N_noxref_10_M0_noxref_s ) capacitor \
 c=0.00309936f //x=3.395 //y=0.915 //x2=0.455 //y2=0.375
cc_975 ( N_noxref_6_c_1144_n N_noxref_11_c_2110_n ) capacitor c=0.00466084f \
 //x=3.985 //y=1.665 //x2=3.985 //y2=0.54
cc_976 ( N_noxref_6_M2_noxref_d N_noxref_11_c_2110_n ) capacitor c=0.0117786f \
 //x=3.395 //y=0.915 //x2=3.985 //y2=0.54
cc_977 ( N_noxref_6_c_1229_n N_noxref_11_c_2124_n ) capacitor c=0.020048f \
 //x=3.67 //y=1.665 //x2=3.1 //y2=0.995
cc_978 ( N_noxref_6_M2_noxref_d N_noxref_11_M1_noxref_d ) capacitor \
 c=5.27807e-19 //x=3.395 //y=0.915 //x2=1.86 //y2=0.91
cc_979 ( N_noxref_6_c_1144_n N_noxref_11_M2_noxref_s ) capacitor c=0.0207678f \
 //x=3.985 //y=1.665 //x2=2.965 //y2=0.375
cc_980 ( N_noxref_6_M2_noxref_d N_noxref_11_M2_noxref_s ) capacitor \
 c=0.0426444f //x=3.395 //y=0.915 //x2=2.965 //y2=0.375
cc_981 ( N_noxref_6_c_1145_n N_D_c_2167_n ) capacitor c=0.00400249f //x=5.92 \
 //y=2.08 //x2=6.66 //y2=4.535
cc_982 ( N_noxref_6_c_1198_n N_D_c_2167_n ) capacitor c=0.00417994f //x=5.92 \
 //y=4.7 //x2=6.66 //y2=4.535
cc_983 ( N_noxref_6_c_1142_n N_D_c_2158_n ) capacitor c=0.0169594f //x=15.795 \
 //y=3.7 //x2=6.66 //y2=2.08
cc_984 ( N_noxref_6_c_1223_n N_D_c_2158_n ) capacitor c=0.00131333f //x=6.035 \
 //y=3.7 //x2=6.66 //y2=2.08
cc_985 ( N_noxref_6_c_1183_n N_D_c_2158_n ) capacitor c=8.12815e-19 //x=4.07 \
 //y=3.7 //x2=6.66 //y2=2.08
cc_986 ( N_noxref_6_c_1145_n N_D_c_2158_n ) capacitor c=0.0781945f //x=5.92 \
 //y=2.08 //x2=6.66 //y2=2.08
cc_987 ( N_noxref_6_c_1151_n N_D_c_2158_n ) capacitor c=0.00308814f //x=5.725 \
 //y=1.915 //x2=6.66 //y2=2.08
cc_988 ( N_noxref_6_M19_noxref_g N_D_M21_noxref_g ) capacitor c=0.0104611f \
 //x=5.82 //y=6.02 //x2=6.7 //y2=6.02
cc_989 ( N_noxref_6_M20_noxref_g N_D_M21_noxref_g ) capacitor c=0.106811f \
 //x=6.26 //y=6.02 //x2=6.7 //y2=6.02
cc_990 ( N_noxref_6_M20_noxref_g N_D_M22_noxref_g ) capacitor c=0.0100341f \
 //x=6.26 //y=6.02 //x2=7.14 //y2=6.02
cc_991 ( N_noxref_6_c_1147_n N_D_c_2177_n ) capacitor c=4.86506e-19 //x=5.725 \
 //y=0.865 //x2=6.695 //y2=0.905
cc_992 ( N_noxref_6_c_1149_n N_D_c_2177_n ) capacitor c=0.00152104f //x=5.725 \
 //y=1.21 //x2=6.695 //y2=0.905
cc_993 ( N_noxref_6_c_1154_n N_D_c_2177_n ) capacitor c=0.0151475f //x=6.255 \
 //y=0.865 //x2=6.695 //y2=0.905
cc_994 ( N_noxref_6_c_1150_n N_D_c_2178_n ) capacitor c=0.00109982f //x=5.725 \
 //y=1.52 //x2=6.695 //y2=1.25
cc_995 ( N_noxref_6_c_1156_n N_D_c_2178_n ) capacitor c=0.0111064f //x=6.255 \
 //y=1.21 //x2=6.695 //y2=1.25
cc_996 ( N_noxref_6_c_1150_n N_D_c_2179_n ) capacitor c=9.57794e-19 //x=5.725 \
 //y=1.52 //x2=6.695 //y2=1.56
cc_997 ( N_noxref_6_c_1151_n N_D_c_2179_n ) capacitor c=0.00662747f //x=5.725 \
 //y=1.915 //x2=6.695 //y2=1.56
cc_998 ( N_noxref_6_c_1156_n N_D_c_2179_n ) capacitor c=0.00862358f //x=6.255 \
 //y=1.21 //x2=6.695 //y2=1.56
cc_999 ( N_noxref_6_c_1154_n N_D_c_2185_n ) capacitor c=0.00124821f //x=6.255 \
 //y=0.865 //x2=7.225 //y2=0.905
cc_1000 ( N_noxref_6_c_1156_n N_D_c_2186_n ) capacitor c=0.00200715f //x=6.255 \
 //y=1.21 //x2=7.225 //y2=1.25
cc_1001 ( N_noxref_6_c_1145_n N_D_c_2188_n ) capacitor c=0.00307062f //x=5.92 \
 //y=2.08 //x2=6.66 //y2=2.08
cc_1002 ( N_noxref_6_c_1151_n N_D_c_2188_n ) capacitor c=0.0179092f //x=5.725 \
 //y=1.915 //x2=6.66 //y2=2.08
cc_1003 ( N_noxref_6_c_1145_n N_D_c_2191_n ) capacitor c=0.00344981f //x=5.92 \
 //y=2.08 //x2=6.69 //y2=4.7
cc_1004 ( N_noxref_6_c_1198_n N_D_c_2191_n ) capacitor c=0.0293367f //x=5.92 \
 //y=4.7 //x2=6.69 //y2=4.7
cc_1005 ( N_noxref_6_c_1144_n N_noxref_13_c_2250_n ) capacitor c=3.04182e-19 \
 //x=3.985 //y=1.665 //x2=5.505 //y2=1.495
cc_1006 ( N_noxref_6_c_1151_n N_noxref_13_c_2250_n ) capacitor c=0.0034165f \
 //x=5.725 //y=1.915 //x2=5.505 //y2=1.495
cc_1007 ( N_noxref_6_c_1145_n N_noxref_13_c_2231_n ) capacitor c=0.0116993f \
 //x=5.92 //y=2.08 //x2=6.39 //y2=1.58
cc_1008 ( N_noxref_6_c_1150_n N_noxref_13_c_2231_n ) capacitor c=0.00703567f \
 //x=5.725 //y=1.52 //x2=6.39 //y2=1.58
cc_1009 ( N_noxref_6_c_1151_n N_noxref_13_c_2231_n ) capacitor c=0.0203514f \
 //x=5.725 //y=1.915 //x2=6.39 //y2=1.58
cc_1010 ( N_noxref_6_c_1153_n N_noxref_13_c_2231_n ) capacitor c=0.00780629f \
 //x=6.1 //y=1.365 //x2=6.39 //y2=1.58
cc_1011 ( N_noxref_6_c_1156_n N_noxref_13_c_2231_n ) capacitor c=0.00339872f \
 //x=6.255 //y=1.21 //x2=6.39 //y2=1.58
cc_1012 ( N_noxref_6_c_1151_n N_noxref_13_c_2238_n ) capacitor c=6.71402e-19 \
 //x=5.725 //y=1.915 //x2=6.475 //y2=1.495
cc_1013 ( N_noxref_6_c_1147_n N_noxref_13_M3_noxref_s ) capacitor c=0.0327502f \
 //x=5.725 //y=0.865 //x2=5.37 //y2=0.365
cc_1014 ( N_noxref_6_c_1150_n N_noxref_13_M3_noxref_s ) capacitor \
 c=3.48408e-19 //x=5.725 //y=1.52 //x2=5.37 //y2=0.365
cc_1015 ( N_noxref_6_c_1154_n N_noxref_13_M3_noxref_s ) capacitor c=0.0120759f \
 //x=6.255 //y=0.865 //x2=5.37 //y2=0.365
cc_1016 ( N_noxref_6_c_1142_n N_noxref_14_c_2283_n ) capacitor c=0.00299723f \
 //x=15.795 //y=3.7 //x2=9.72 //y2=1.58
cc_1017 ( N_noxref_6_c_1142_n N_noxref_14_c_2290_n ) capacitor c=0.00187232f \
 //x=15.795 //y=3.7 //x2=9.805 //y2=1.495
cc_1018 ( N_noxref_6_c_1142_n N_noxref_14_c_2291_n ) capacitor c=4.7198e-19 \
 //x=15.795 //y=3.7 //x2=10.69 //y2=0.53
cc_1019 ( N_noxref_6_c_1142_n N_noxref_15_c_2336_n ) capacitor c=0.00299723f \
 //x=15.795 //y=3.7 //x2=13.05 //y2=1.58
cc_1020 ( N_noxref_6_c_1142_n N_noxref_15_c_2343_n ) capacitor c=0.00187232f \
 //x=15.795 //y=3.7 //x2=13.135 //y2=1.495
cc_1021 ( N_noxref_6_c_1142_n N_noxref_15_c_2344_n ) capacitor c=4.7198e-19 \
 //x=15.795 //y=3.7 //x2=14.02 //y2=0.53
cc_1022 ( N_noxref_6_c_1142_n N_noxref_15_M7_noxref_s ) capacitor \
 c=3.97107e-19 //x=15.795 //y=3.7 //x2=12.03 //y2=0.365
cc_1023 ( N_noxref_6_c_1142_n N_noxref_16_c_2408_n ) capacitor c=0.00188872f \
 //x=15.795 //y=3.7 //x2=15.495 //y2=1.495
cc_1024 ( N_noxref_6_c_1161_n N_noxref_16_c_2408_n ) capacitor c=0.0034165f \
 //x=15.715 //y=1.915 //x2=15.495 //y2=1.495
cc_1025 ( N_noxref_6_c_1142_n N_noxref_16_c_2389_n ) capacitor c=0.0056636f \
 //x=15.795 //y=3.7 //x2=16.38 //y2=1.58
cc_1026 ( N_noxref_6_c_1146_n N_noxref_16_c_2389_n ) capacitor c=0.011766f \
 //x=15.91 //y=2.08 //x2=16.38 //y2=1.58
cc_1027 ( N_noxref_6_c_1160_n N_noxref_16_c_2389_n ) capacitor c=0.00703567f \
 //x=15.715 //y=1.52 //x2=16.38 //y2=1.58
cc_1028 ( N_noxref_6_c_1161_n N_noxref_16_c_2389_n ) capacitor c=0.0207598f \
 //x=15.715 //y=1.915 //x2=16.38 //y2=1.58
cc_1029 ( N_noxref_6_c_1163_n N_noxref_16_c_2389_n ) capacitor c=0.00780629f \
 //x=16.09 //y=1.365 //x2=16.38 //y2=1.58
cc_1030 ( N_noxref_6_c_1166_n N_noxref_16_c_2389_n ) capacitor c=0.00339872f \
 //x=16.245 //y=1.21 //x2=16.38 //y2=1.58
cc_1031 ( N_noxref_6_c_1161_n N_noxref_16_c_2396_n ) capacitor c=6.71402e-19 \
 //x=15.715 //y=1.915 //x2=16.465 //y2=1.495
cc_1032 ( N_noxref_6_c_1157_n N_noxref_16_M9_noxref_s ) capacitor c=0.0326577f \
 //x=15.715 //y=0.865 //x2=15.36 //y2=0.365
cc_1033 ( N_noxref_6_c_1160_n N_noxref_16_M9_noxref_s ) capacitor \
 c=3.48408e-19 //x=15.715 //y=1.52 //x2=15.36 //y2=0.365
cc_1034 ( N_noxref_6_c_1164_n N_noxref_16_M9_noxref_s ) capacitor c=0.0120759f \
 //x=16.245 //y=0.865 //x2=15.36 //y2=0.365
cc_1035 ( N_noxref_7_c_1395_n N_noxref_8_c_1544_n ) capacitor c=0.0110241f \
 //x=19.125 //y=3.33 //x2=19.865 //y2=4.07
cc_1036 ( N_noxref_7_c_1399_n N_noxref_8_c_1544_n ) capacitor c=8.88358e-19 \
 //x=17.505 //y=3.33 //x2=19.865 //y2=4.07
cc_1037 ( N_noxref_7_c_1416_n N_noxref_8_c_1544_n ) capacitor c=0.0140425f \
 //x=16.825 //y=5.2 //x2=19.865 //y2=4.07
cc_1038 ( N_noxref_7_c_1420_n N_noxref_8_c_1544_n ) capacitor c=0.0135379f \
 //x=16.115 //y=5.2 //x2=19.865 //y2=4.07
cc_1039 ( N_noxref_7_c_1401_n N_noxref_8_c_1544_n ) capacitor c=0.023177f \
 //x=17.39 //y=3.33 //x2=19.865 //y2=4.07
cc_1040 ( N_noxref_7_c_1402_n N_noxref_8_c_1544_n ) capacitor c=0.0242126f \
 //x=19.24 //y=2.08 //x2=19.865 //y2=4.07
cc_1041 ( N_noxref_7_c_1435_n N_noxref_8_c_1544_n ) capacitor c=0.00844647f \
 //x=19.24 //y=4.7 //x2=19.865 //y2=4.07
cc_1042 ( N_noxref_7_c_1401_n N_noxref_8_c_1549_n ) capacitor c=3.49822e-19 \
 //x=17.39 //y=3.33 //x2=14.06 //y2=4.07
cc_1043 ( N_noxref_7_c_1402_n N_noxref_8_c_1797_n ) capacitor c=0.00400249f \
 //x=19.24 //y=2.08 //x2=19.98 //y2=4.535
cc_1044 ( N_noxref_7_c_1435_n N_noxref_8_c_1797_n ) capacitor c=0.00417994f \
 //x=19.24 //y=4.7 //x2=19.98 //y2=4.535
cc_1045 ( N_noxref_7_c_1395_n N_noxref_8_c_1550_n ) capacitor c=0.00720056f \
 //x=19.125 //y=3.33 //x2=19.98 //y2=2.08
cc_1046 ( N_noxref_7_c_1401_n N_noxref_8_c_1550_n ) capacitor c=0.00107361f \
 //x=17.39 //y=3.33 //x2=19.98 //y2=2.08
cc_1047 ( N_noxref_7_c_1402_n N_noxref_8_c_1550_n ) capacitor c=0.0810987f \
 //x=19.24 //y=2.08 //x2=19.98 //y2=2.08
cc_1048 ( N_noxref_7_c_1407_n N_noxref_8_c_1550_n ) capacitor c=0.00308814f \
 //x=19.045 //y=1.915 //x2=19.98 //y2=2.08
cc_1049 ( N_noxref_7_M35_noxref_g N_noxref_8_M37_noxref_g ) capacitor \
 c=0.0104611f //x=19.14 //y=6.02 //x2=20.02 //y2=6.02
cc_1050 ( N_noxref_7_M36_noxref_g N_noxref_8_M37_noxref_g ) capacitor \
 c=0.106811f //x=19.58 //y=6.02 //x2=20.02 //y2=6.02
cc_1051 ( N_noxref_7_M36_noxref_g N_noxref_8_M38_noxref_g ) capacitor \
 c=0.0100341f //x=19.58 //y=6.02 //x2=20.46 //y2=6.02
cc_1052 ( N_noxref_7_c_1403_n N_noxref_8_c_1806_n ) capacitor c=4.86506e-19 \
 //x=19.045 //y=0.865 //x2=20.015 //y2=0.905
cc_1053 ( N_noxref_7_c_1405_n N_noxref_8_c_1806_n ) capacitor c=0.00152104f \
 //x=19.045 //y=1.21 //x2=20.015 //y2=0.905
cc_1054 ( N_noxref_7_c_1410_n N_noxref_8_c_1806_n ) capacitor c=0.0151475f \
 //x=19.575 //y=0.865 //x2=20.015 //y2=0.905
cc_1055 ( N_noxref_7_c_1406_n N_noxref_8_c_1809_n ) capacitor c=0.00109982f \
 //x=19.045 //y=1.52 //x2=20.015 //y2=1.25
cc_1056 ( N_noxref_7_c_1412_n N_noxref_8_c_1809_n ) capacitor c=0.0111064f \
 //x=19.575 //y=1.21 //x2=20.015 //y2=1.25
cc_1057 ( N_noxref_7_c_1406_n N_noxref_8_c_1811_n ) capacitor c=9.57794e-19 \
 //x=19.045 //y=1.52 //x2=20.015 //y2=1.56
cc_1058 ( N_noxref_7_c_1407_n N_noxref_8_c_1811_n ) capacitor c=0.00662747f \
 //x=19.045 //y=1.915 //x2=20.015 //y2=1.56
cc_1059 ( N_noxref_7_c_1412_n N_noxref_8_c_1811_n ) capacitor c=0.00862358f \
 //x=19.575 //y=1.21 //x2=20.015 //y2=1.56
cc_1060 ( N_noxref_7_c_1410_n N_noxref_8_c_1814_n ) capacitor c=0.00124821f \
 //x=19.575 //y=0.865 //x2=20.545 //y2=0.905
cc_1061 ( N_noxref_7_c_1412_n N_noxref_8_c_1815_n ) capacitor c=0.00200715f \
 //x=19.575 //y=1.21 //x2=20.545 //y2=1.25
cc_1062 ( N_noxref_7_c_1402_n N_noxref_8_c_1816_n ) capacitor c=0.00307062f \
 //x=19.24 //y=2.08 //x2=19.98 //y2=2.08
cc_1063 ( N_noxref_7_c_1407_n N_noxref_8_c_1816_n ) capacitor c=0.0179092f \
 //x=19.045 //y=1.915 //x2=19.98 //y2=2.08
cc_1064 ( N_noxref_7_c_1402_n N_noxref_8_c_1818_n ) capacitor c=0.00344981f \
 //x=19.24 //y=2.08 //x2=20.01 //y2=4.7
cc_1065 ( N_noxref_7_c_1435_n N_noxref_8_c_1818_n ) capacitor c=0.0293367f \
 //x=19.24 //y=4.7 //x2=20.01 //y2=4.7
cc_1066 ( N_noxref_7_c_1395_n N_Q_c_1900_n ) capacitor c=0.175696f //x=19.125 \
 //y=3.33 //x2=20.605 //y2=3.7
cc_1067 ( N_noxref_7_c_1399_n N_Q_c_1900_n ) capacitor c=0.0293967f //x=17.505 \
 //y=3.33 //x2=20.605 //y2=3.7
cc_1068 ( N_noxref_7_c_1486_p N_Q_c_1900_n ) capacitor c=0.0037701f //x=17.035 \
 //y=1.655 //x2=20.605 //y2=3.7
cc_1069 ( N_noxref_7_c_1401_n N_Q_c_1900_n ) capacitor c=0.0206034f //x=17.39 \
 //y=3.33 //x2=20.605 //y2=3.7
cc_1070 ( N_noxref_7_c_1402_n N_Q_c_1900_n ) capacitor c=0.0205569f //x=19.24 \
 //y=2.08 //x2=20.605 //y2=3.7
cc_1071 ( N_noxref_7_c_1401_n N_Q_c_1901_n ) capacitor c=0.00117715f //x=17.39 \
 //y=3.33 //x2=16.765 //y2=3.7
cc_1072 ( N_noxref_7_c_1401_n Q ) capacitor c=3.49822e-19 //x=17.39 //y=3.33 \
 //x2=20.72 //y2=2.22
cc_1073 ( N_noxref_7_c_1402_n Q ) capacitor c=0.00407494f //x=19.24 //y=2.08 \
 //x2=20.72 //y2=2.22
cc_1074 ( N_noxref_7_c_1416_n N_Q_c_1941_n ) capacitor c=0.0129336f //x=16.825 \
 //y=5.2 //x2=16.65 //y2=4.535
cc_1075 ( N_noxref_7_c_1401_n N_Q_c_1941_n ) capacitor c=0.0101284f //x=17.39 \
 //y=3.33 //x2=16.65 //y2=4.535
cc_1076 ( N_noxref_7_c_1399_n N_Q_c_1903_n ) capacitor c=0.00720056f \
 //x=17.505 //y=3.33 //x2=16.65 //y2=2.08
cc_1077 ( N_noxref_7_c_1401_n N_Q_c_1903_n ) capacitor c=0.0759968f //x=17.39 \
 //y=3.33 //x2=16.65 //y2=2.08
cc_1078 ( N_noxref_7_c_1402_n N_Q_c_1903_n ) capacitor c=0.001003f //x=19.24 \
 //y=2.08 //x2=16.65 //y2=2.08
cc_1079 ( N_noxref_7_M36_noxref_g N_Q_c_1915_n ) capacitor c=0.017965f \
 //x=19.58 //y=6.02 //x2=20.155 //y2=5.2
cc_1080 ( N_noxref_7_c_1402_n N_Q_c_1919_n ) capacitor c=0.00549854f //x=19.24 \
 //y=2.08 //x2=19.445 //y2=5.2
cc_1081 ( N_noxref_7_M35_noxref_g N_Q_c_1919_n ) capacitor c=0.0177326f \
 //x=19.14 //y=6.02 //x2=19.445 //y2=5.2
cc_1082 ( N_noxref_7_c_1435_n N_Q_c_1919_n ) capacitor c=0.00582246f //x=19.24 \
 //y=4.7 //x2=19.445 //y2=5.2
cc_1083 ( N_noxref_7_c_1416_n N_Q_M33_noxref_g ) capacitor c=0.0166421f \
 //x=16.825 //y=5.2 //x2=16.69 //y2=6.02
cc_1084 ( N_noxref_7_M33_noxref_d N_Q_M33_noxref_g ) capacitor c=0.0173476f \
 //x=16.765 //y=5.02 //x2=16.69 //y2=6.02
cc_1085 ( N_noxref_7_c_1422_n N_Q_M34_noxref_g ) capacitor c=0.0199348f \
 //x=17.305 //y=5.2 //x2=17.13 //y2=6.02
cc_1086 ( N_noxref_7_M33_noxref_d N_Q_M34_noxref_g ) capacitor c=0.0179769f \
 //x=16.765 //y=5.02 //x2=17.13 //y2=6.02
cc_1087 ( N_noxref_7_M10_noxref_d N_Q_c_1949_n ) capacitor c=0.00217566f \
 //x=16.76 //y=0.905 //x2=16.685 //y2=0.905
cc_1088 ( N_noxref_7_M10_noxref_d N_Q_c_1952_n ) capacitor c=0.0034598f \
 //x=16.76 //y=0.905 //x2=16.685 //y2=1.25
cc_1089 ( N_noxref_7_M10_noxref_d N_Q_c_1954_n ) capacitor c=0.0065582f \
 //x=16.76 //y=0.905 //x2=16.685 //y2=1.56
cc_1090 ( N_noxref_7_c_1401_n N_Q_c_1987_n ) capacitor c=0.0142673f //x=17.39 \
 //y=3.33 //x2=17.055 //y2=4.79
cc_1091 ( N_noxref_7_c_1509_p N_Q_c_1987_n ) capacitor c=0.00408717f //x=16.91 \
 //y=5.2 //x2=17.055 //y2=4.79
cc_1092 ( N_noxref_7_M10_noxref_d N_Q_c_1989_n ) capacitor c=0.00241102f \
 //x=16.76 //y=0.905 //x2=17.06 //y2=0.75
cc_1093 ( N_noxref_7_c_1400_n N_Q_c_1990_n ) capacitor c=0.00359704f \
 //x=17.305 //y=1.655 //x2=17.06 //y2=1.405
cc_1094 ( N_noxref_7_M10_noxref_d N_Q_c_1990_n ) capacitor c=0.0138845f \
 //x=16.76 //y=0.905 //x2=17.06 //y2=1.405
cc_1095 ( N_noxref_7_M10_noxref_d N_Q_c_1957_n ) capacitor c=0.00132245f \
 //x=16.76 //y=0.905 //x2=17.215 //y2=0.905
cc_1096 ( N_noxref_7_c_1400_n N_Q_c_1958_n ) capacitor c=0.00457401f \
 //x=17.305 //y=1.655 //x2=17.215 //y2=1.25
cc_1097 ( N_noxref_7_M10_noxref_d N_Q_c_1958_n ) capacitor c=0.00566463f \
 //x=16.76 //y=0.905 //x2=17.215 //y2=1.25
cc_1098 ( N_noxref_7_c_1401_n N_Q_c_1959_n ) capacitor c=0.00877984f //x=17.39 \
 //y=3.33 //x2=16.65 //y2=2.08
cc_1099 ( N_noxref_7_c_1401_n N_Q_c_1996_n ) capacitor c=0.00306024f //x=17.39 \
 //y=3.33 //x2=16.65 //y2=1.915
cc_1100 ( N_noxref_7_M10_noxref_d N_Q_c_1996_n ) capacitor c=0.00660593f \
 //x=16.76 //y=0.905 //x2=16.65 //y2=1.915
cc_1101 ( N_noxref_7_c_1416_n N_Q_c_1961_n ) capacitor c=0.00346635f \
 //x=16.825 //y=5.2 //x2=16.68 //y2=4.7
cc_1102 ( N_noxref_7_c_1401_n N_Q_c_1961_n ) capacitor c=0.00533692f //x=17.39 \
 //y=3.33 //x2=16.68 //y2=4.7
cc_1103 ( N_noxref_7_M36_noxref_g N_Q_M35_noxref_d ) capacitor c=0.0173476f \
 //x=19.58 //y=6.02 //x2=19.215 //y2=5.02
cc_1104 ( N_noxref_7_c_1486_p N_noxref_16_c_2408_n ) capacitor c=3.15806e-19 \
 //x=17.035 //y=1.655 //x2=15.495 //y2=1.495
cc_1105 ( N_noxref_7_c_1486_p N_noxref_16_c_2396_n ) capacitor c=0.0203424f \
 //x=17.035 //y=1.655 //x2=16.465 //y2=1.495
cc_1106 ( N_noxref_7_c_1400_n N_noxref_16_c_2397_n ) capacitor c=0.0046686f \
 //x=17.305 //y=1.655 //x2=17.35 //y2=0.53
cc_1107 ( N_noxref_7_M10_noxref_d N_noxref_16_c_2397_n ) capacitor \
 c=0.0117932f //x=16.76 //y=0.905 //x2=17.35 //y2=0.53
cc_1108 ( N_noxref_7_c_1399_n N_noxref_16_M9_noxref_s ) capacitor \
 c=3.47564e-19 //x=17.505 //y=3.33 //x2=15.36 //y2=0.365
cc_1109 ( N_noxref_7_c_1400_n N_noxref_16_M9_noxref_s ) capacitor c=0.0141735f \
 //x=17.305 //y=1.655 //x2=15.36 //y2=0.365
cc_1110 ( N_noxref_7_M10_noxref_d N_noxref_16_M9_noxref_s ) capacitor \
 c=0.043966f //x=16.76 //y=0.905 //x2=15.36 //y2=0.365
cc_1111 ( N_noxref_7_c_1395_n N_noxref_17_c_2460_n ) capacitor c=0.00241565f \
 //x=19.125 //y=3.33 //x2=18.825 //y2=1.495
cc_1112 ( N_noxref_7_c_1400_n N_noxref_17_c_2460_n ) capacitor c=3.22188e-19 \
 //x=17.305 //y=1.655 //x2=18.825 //y2=1.495
cc_1113 ( N_noxref_7_c_1407_n N_noxref_17_c_2460_n ) capacitor c=0.0034165f \
 //x=19.045 //y=1.915 //x2=18.825 //y2=1.495
cc_1114 ( N_noxref_7_c_1395_n N_noxref_17_c_2443_n ) capacitor c=0.00649414f \
 //x=19.125 //y=3.33 //x2=19.71 //y2=1.58
cc_1115 ( N_noxref_7_c_1402_n N_noxref_17_c_2443_n ) capacitor c=0.011692f \
 //x=19.24 //y=2.08 //x2=19.71 //y2=1.58
cc_1116 ( N_noxref_7_c_1406_n N_noxref_17_c_2443_n ) capacitor c=0.00703567f \
 //x=19.045 //y=1.52 //x2=19.71 //y2=1.58
cc_1117 ( N_noxref_7_c_1407_n N_noxref_17_c_2443_n ) capacitor c=0.0203514f \
 //x=19.045 //y=1.915 //x2=19.71 //y2=1.58
cc_1118 ( N_noxref_7_c_1409_n N_noxref_17_c_2443_n ) capacitor c=0.00780629f \
 //x=19.42 //y=1.365 //x2=19.71 //y2=1.58
cc_1119 ( N_noxref_7_c_1412_n N_noxref_17_c_2443_n ) capacitor c=0.00339872f \
 //x=19.575 //y=1.21 //x2=19.71 //y2=1.58
cc_1120 ( N_noxref_7_c_1407_n N_noxref_17_c_2450_n ) capacitor c=6.71402e-19 \
 //x=19.045 //y=1.915 //x2=19.795 //y2=1.495
cc_1121 ( N_noxref_7_c_1403_n N_noxref_17_M11_noxref_s ) capacitor \
 c=0.0326577f //x=19.045 //y=0.865 //x2=18.69 //y2=0.365
cc_1122 ( N_noxref_7_c_1406_n N_noxref_17_M11_noxref_s ) capacitor \
 c=3.48408e-19 //x=19.045 //y=1.52 //x2=18.69 //y2=0.365
cc_1123 ( N_noxref_7_c_1410_n N_noxref_17_M11_noxref_s ) capacitor \
 c=0.0120759f //x=19.575 //y=0.865 //x2=18.69 //y2=0.365
cc_1124 ( N_noxref_8_c_1544_n N_Q_c_1900_n ) capacitor c=0.304477f //x=19.865 \
 //y=4.07 //x2=20.605 //y2=3.7
cc_1125 ( N_noxref_8_c_1550_n N_Q_c_1900_n ) capacitor c=0.0255669f //x=19.98 \
 //y=2.08 //x2=20.605 //y2=3.7
cc_1126 ( N_noxref_8_c_1822_p N_Q_c_1900_n ) capacitor c=0.00624857f \
 //x=20.385 //y=4.79 //x2=20.605 //y2=3.7
cc_1127 ( N_noxref_8_c_1818_n N_Q_c_1900_n ) capacitor c=3.27069e-19 //x=20.01 \
 //y=4.7 //x2=20.605 //y2=3.7
cc_1128 ( N_noxref_8_c_1544_n N_Q_c_1901_n ) capacitor c=0.0291169f //x=19.865 \
 //y=4.07 //x2=16.765 //y2=3.7
cc_1129 ( N_noxref_8_c_1544_n Q ) capacitor c=0.00642908f //x=19.865 //y=4.07 \
 //x2=20.72 //y2=2.22
cc_1130 ( N_noxref_8_c_1797_n Q ) capacitor c=0.0101115f //x=19.98 //y=4.535 \
 //x2=20.72 //y2=2.22
cc_1131 ( N_noxref_8_c_1550_n Q ) capacitor c=0.0786723f //x=19.98 //y=2.08 \
 //x2=20.72 //y2=2.22
cc_1132 ( N_noxref_8_c_1822_p Q ) capacitor c=0.0142673f //x=20.385 //y=4.79 \
 //x2=20.72 //y2=2.22
cc_1133 ( N_noxref_8_c_1816_n Q ) capacitor c=0.00877984f //x=19.98 //y=2.08 \
 //x2=20.72 //y2=2.22
cc_1134 ( N_noxref_8_c_1830_p Q ) capacitor c=0.00306024f //x=19.98 //y=1.915 \
 //x2=20.72 //y2=2.22
cc_1135 ( N_noxref_8_c_1818_n Q ) capacitor c=0.00533692f //x=20.01 //y=4.7 \
 //x2=20.72 //y2=2.22
cc_1136 ( N_noxref_8_c_1544_n N_Q_c_1941_n ) capacitor c=0.00135863f \
 //x=19.865 //y=4.07 //x2=16.65 //y2=4.535
cc_1137 ( N_noxref_8_c_1544_n N_Q_c_1903_n ) capacitor c=0.022647f //x=19.865 \
 //y=4.07 //x2=16.65 //y2=2.08
cc_1138 ( N_noxref_8_c_1549_n N_Q_c_1903_n ) capacitor c=9.30282e-19 //x=14.06 \
 //y=4.07 //x2=16.65 //y2=2.08
cc_1139 ( N_noxref_8_c_1544_n N_Q_c_1915_n ) capacitor c=0.00208151f \
 //x=19.865 //y=4.07 //x2=20.155 //y2=5.2
cc_1140 ( N_noxref_8_c_1797_n N_Q_c_1915_n ) capacitor c=0.0129205f //x=19.98 \
 //y=4.535 //x2=20.155 //y2=5.2
cc_1141 ( N_noxref_8_M37_noxref_g N_Q_c_1915_n ) capacitor c=0.0166421f \
 //x=20.02 //y=6.02 //x2=20.155 //y2=5.2
cc_1142 ( N_noxref_8_c_1818_n N_Q_c_1915_n ) capacitor c=0.00346627f //x=20.01 \
 //y=4.7 //x2=20.155 //y2=5.2
cc_1143 ( N_noxref_8_c_1544_n N_Q_c_1919_n ) capacitor c=0.01319f //x=19.865 \
 //y=4.07 //x2=19.445 //y2=5.2
cc_1144 ( N_noxref_8_M38_noxref_g N_Q_c_1921_n ) capacitor c=0.0206783f \
 //x=20.46 //y=6.02 //x2=20.635 //y2=5.2
cc_1145 ( N_noxref_8_c_1841_p N_Q_c_1905_n ) capacitor c=0.00359704f //x=20.39 \
 //y=1.405 //x2=20.635 //y2=1.655
cc_1146 ( N_noxref_8_c_1815_n N_Q_c_1905_n ) capacitor c=0.00457401f \
 //x=20.545 //y=1.25 //x2=20.635 //y2=1.655
cc_1147 ( N_noxref_8_c_1822_p N_Q_c_2024_n ) capacitor c=0.00421574f \
 //x=20.385 //y=4.79 //x2=20.24 //y2=5.2
cc_1148 ( N_noxref_8_c_1544_n N_Q_c_1987_n ) capacitor c=0.00756255f \
 //x=19.865 //y=4.07 //x2=17.055 //y2=4.79
cc_1149 ( N_noxref_8_c_1544_n N_Q_c_1961_n ) capacitor c=0.00160199f \
 //x=19.865 //y=4.07 //x2=16.68 //y2=4.7
cc_1150 ( N_noxref_8_c_1806_n N_Q_M12_noxref_d ) capacitor c=0.00217566f \
 //x=20.015 //y=0.905 //x2=20.09 //y2=0.905
cc_1151 ( N_noxref_8_c_1809_n N_Q_M12_noxref_d ) capacitor c=0.0034598f \
 //x=20.015 //y=1.25 //x2=20.09 //y2=0.905
cc_1152 ( N_noxref_8_c_1811_n N_Q_M12_noxref_d ) capacitor c=0.0065582f \
 //x=20.015 //y=1.56 //x2=20.09 //y2=0.905
cc_1153 ( N_noxref_8_c_1849_p N_Q_M12_noxref_d ) capacitor c=0.00241102f \
 //x=20.39 //y=0.75 //x2=20.09 //y2=0.905
cc_1154 ( N_noxref_8_c_1841_p N_Q_M12_noxref_d ) capacitor c=0.0138845f \
 //x=20.39 //y=1.405 //x2=20.09 //y2=0.905
cc_1155 ( N_noxref_8_c_1814_n N_Q_M12_noxref_d ) capacitor c=0.00132245f \
 //x=20.545 //y=0.905 //x2=20.09 //y2=0.905
cc_1156 ( N_noxref_8_c_1815_n N_Q_M12_noxref_d ) capacitor c=0.00566463f \
 //x=20.545 //y=1.25 //x2=20.09 //y2=0.905
cc_1157 ( N_noxref_8_c_1830_p N_Q_M12_noxref_d ) capacitor c=0.00660593f \
 //x=19.98 //y=1.915 //x2=20.09 //y2=0.905
cc_1158 ( N_noxref_8_M37_noxref_g N_Q_M37_noxref_d ) capacitor c=0.0173476f \
 //x=20.02 //y=6.02 //x2=20.095 //y2=5.02
cc_1159 ( N_noxref_8_M38_noxref_g N_Q_M37_noxref_d ) capacitor c=0.0179769f \
 //x=20.46 //y=6.02 //x2=20.095 //y2=5.02
cc_1160 ( N_noxref_8_c_1556_n N_noxref_10_c_2083_n ) capacitor c=0.0034165f \
 //x=0.81 //y=1.915 //x2=0.59 //y2=1.505
cc_1161 ( N_noxref_8_c_1542_n N_noxref_10_c_2058_n ) capacitor c=0.00179505f \
 //x=9.875 //y=4.07 //x2=1.475 //y2=1.59
cc_1162 ( N_noxref_8_c_1543_n N_noxref_10_c_2058_n ) capacitor c=0.00102628f \
 //x=1.225 //y=4.07 //x2=1.475 //y2=1.59
cc_1163 ( N_noxref_8_c_1545_n N_noxref_10_c_2058_n ) capacitor c=0.0122033f \
 //x=1.11 //y=2.08 //x2=1.475 //y2=1.59
cc_1164 ( N_noxref_8_c_1555_n N_noxref_10_c_2058_n ) capacitor c=0.00703864f \
 //x=0.81 //y=1.53 //x2=1.475 //y2=1.59
cc_1165 ( N_noxref_8_c_1556_n N_noxref_10_c_2058_n ) capacitor c=0.0259045f \
 //x=0.81 //y=1.915 //x2=1.475 //y2=1.59
cc_1166 ( N_noxref_8_c_1558_n N_noxref_10_c_2058_n ) capacitor c=0.00708583f \
 //x=1.185 //y=1.375 //x2=1.475 //y2=1.59
cc_1167 ( N_noxref_8_c_1561_n N_noxref_10_c_2058_n ) capacitor c=0.00698822f \
 //x=1.34 //y=1.22 //x2=1.475 //y2=1.59
cc_1168 ( N_noxref_8_c_1542_n N_noxref_10_c_2076_n ) capacitor c=0.0058169f \
 //x=9.875 //y=4.07 //x2=2.445 //y2=1.59
cc_1169 ( N_noxref_8_c_1542_n N_noxref_10_M0_noxref_s ) capacitor \
 c=0.00262629f //x=9.875 //y=4.07 //x2=0.455 //y2=0.375
cc_1170 ( N_noxref_8_c_1552_n N_noxref_10_M0_noxref_s ) capacitor c=0.0327271f \
 //x=0.81 //y=0.875 //x2=0.455 //y2=0.375
cc_1171 ( N_noxref_8_c_1555_n N_noxref_10_M0_noxref_s ) capacitor \
 c=7.99997e-19 //x=0.81 //y=1.53 //x2=0.455 //y2=0.375
cc_1172 ( N_noxref_8_c_1556_n N_noxref_10_M0_noxref_s ) capacitor \
 c=0.00122123f //x=0.81 //y=1.915 //x2=0.455 //y2=0.375
cc_1173 ( N_noxref_8_c_1559_n N_noxref_10_M0_noxref_s ) capacitor c=0.0121427f \
 //x=1.34 //y=0.875 //x2=0.455 //y2=0.375
cc_1174 ( N_noxref_8_c_1542_n N_noxref_11_c_2105_n ) capacitor c=0.0020922f \
 //x=9.875 //y=4.07 //x2=3.015 //y2=0.995
cc_1175 ( N_noxref_8_c_1542_n N_noxref_11_M2_noxref_s ) capacitor \
 c=0.00143334f //x=9.875 //y=4.07 //x2=2.965 //y2=0.375
cc_1176 ( N_noxref_8_c_1542_n N_D_c_2158_n ) capacitor c=0.0169317f //x=9.875 \
 //y=4.07 //x2=6.66 //y2=2.08
cc_1177 ( N_noxref_8_c_1658_n N_noxref_14_c_2290_n ) capacitor c=0.00623646f \
 //x=10.025 //y=1.56 //x2=9.805 //y2=1.495
cc_1178 ( N_noxref_8_c_1663_n N_noxref_14_c_2290_n ) capacitor c=0.00176439f \
 //x=9.99 //y=2.08 //x2=9.805 //y2=1.495
cc_1179 ( N_noxref_8_c_1546_n N_noxref_14_c_2291_n ) capacitor c=0.0016032f \
 //x=9.99 //y=2.08 //x2=10.69 //y2=0.53
cc_1180 ( N_noxref_8_c_1653_n N_noxref_14_c_2291_n ) capacitor c=0.0188655f \
 //x=10.025 //y=0.905 //x2=10.69 //y2=0.53
cc_1181 ( N_noxref_8_c_1661_n N_noxref_14_c_2291_n ) capacitor c=0.00656458f \
 //x=10.555 //y=0.905 //x2=10.69 //y2=0.53
cc_1182 ( N_noxref_8_c_1663_n N_noxref_14_c_2291_n ) capacitor c=2.1838e-19 \
 //x=9.99 //y=2.08 //x2=10.69 //y2=0.53
cc_1183 ( N_noxref_8_c_1653_n N_noxref_14_M5_noxref_s ) capacitor \
 c=0.00623646f //x=10.025 //y=0.905 //x2=8.7 //y2=0.365
cc_1184 ( N_noxref_8_c_1661_n N_noxref_14_M5_noxref_s ) capacitor c=0.0143002f \
 //x=10.555 //y=0.905 //x2=8.7 //y2=0.365
cc_1185 ( N_noxref_8_c_1662_n N_noxref_14_M5_noxref_s ) capacitor \
 c=0.00290153f //x=10.555 //y=1.25 //x2=8.7 //y2=0.365
cc_1186 ( N_noxref_8_c_1782_n N_noxref_15_c_2355_n ) capacitor c=3.15806e-19 \
 //x=13.705 //y=1.655 //x2=12.165 //y2=1.495
cc_1187 ( N_noxref_8_c_1782_n N_noxref_15_c_2343_n ) capacitor c=0.0203424f \
 //x=13.705 //y=1.655 //x2=13.135 //y2=1.495
cc_1188 ( N_noxref_8_c_1548_n N_noxref_15_c_2344_n ) capacitor c=0.00467111f \
 //x=13.975 //y=1.655 //x2=14.02 //y2=0.53
cc_1189 ( N_noxref_8_M8_noxref_d N_noxref_15_c_2344_n ) capacitor c=0.0117932f \
 //x=13.43 //y=0.905 //x2=14.02 //y2=0.53
cc_1190 ( N_noxref_8_c_1548_n N_noxref_15_M7_noxref_s ) capacitor c=0.014284f \
 //x=13.975 //y=1.655 //x2=12.03 //y2=0.365
cc_1191 ( N_noxref_8_M8_noxref_d N_noxref_15_M7_noxref_s ) capacitor \
 c=0.043966f //x=13.43 //y=0.905 //x2=12.03 //y2=0.365
cc_1192 ( N_noxref_8_c_1548_n N_noxref_16_c_2408_n ) capacitor c=3.22188e-19 \
 //x=13.975 //y=1.655 //x2=15.495 //y2=1.495
cc_1193 ( N_noxref_8_c_1544_n N_noxref_16_c_2389_n ) capacitor c=0.00234538f \
 //x=19.865 //y=4.07 //x2=16.38 //y2=1.58
cc_1194 ( N_noxref_8_c_1544_n N_noxref_16_c_2396_n ) capacitor c=9.02759e-19 \
 //x=19.865 //y=4.07 //x2=16.465 //y2=1.495
cc_1195 ( N_noxref_8_c_1811_n N_noxref_17_c_2450_n ) capacitor c=0.00623646f \
 //x=20.015 //y=1.56 //x2=19.795 //y2=1.495
cc_1196 ( N_noxref_8_c_1816_n N_noxref_17_c_2450_n ) capacitor c=0.00176439f \
 //x=19.98 //y=2.08 //x2=19.795 //y2=1.495
cc_1197 ( N_noxref_8_c_1550_n N_noxref_17_c_2451_n ) capacitor c=0.0016032f \
 //x=19.98 //y=2.08 //x2=20.68 //y2=0.53
cc_1198 ( N_noxref_8_c_1806_n N_noxref_17_c_2451_n ) capacitor c=0.0188655f \
 //x=20.015 //y=0.905 //x2=20.68 //y2=0.53
cc_1199 ( N_noxref_8_c_1814_n N_noxref_17_c_2451_n ) capacitor c=0.00656458f \
 //x=20.545 //y=0.905 //x2=20.68 //y2=0.53
cc_1200 ( N_noxref_8_c_1816_n N_noxref_17_c_2451_n ) capacitor c=2.1838e-19 \
 //x=19.98 //y=2.08 //x2=20.68 //y2=0.53
cc_1201 ( N_noxref_8_c_1806_n N_noxref_17_M11_noxref_s ) capacitor \
 c=0.00623646f //x=20.015 //y=0.905 //x2=18.69 //y2=0.365
cc_1202 ( N_noxref_8_c_1814_n N_noxref_17_M11_noxref_s ) capacitor \
 c=0.0143002f //x=20.545 //y=0.905 //x2=18.69 //y2=0.365
cc_1203 ( N_noxref_8_c_1815_n N_noxref_17_M11_noxref_s ) capacitor \
 c=0.00290153f //x=20.545 //y=1.25 //x2=18.69 //y2=0.365
cc_1204 ( N_Q_c_1901_n N_noxref_16_c_2396_n ) capacitor c=5.09612e-19 \
 //x=16.765 //y=3.7 //x2=16.465 //y2=1.495
cc_1205 ( N_Q_c_1954_n N_noxref_16_c_2396_n ) capacitor c=0.00623646f \
 //x=16.685 //y=1.56 //x2=16.465 //y2=1.495
cc_1206 ( N_Q_c_1959_n N_noxref_16_c_2396_n ) capacitor c=0.00176439f \
 //x=16.65 //y=2.08 //x2=16.465 //y2=1.495
cc_1207 ( N_Q_c_1900_n N_noxref_16_c_2397_n ) capacitor c=3.61497e-19 \
 //x=20.605 //y=3.7 //x2=17.35 //y2=0.53
cc_1208 ( N_Q_c_1903_n N_noxref_16_c_2397_n ) capacitor c=0.00160293f \
 //x=16.65 //y=2.08 //x2=17.35 //y2=0.53
cc_1209 ( N_Q_c_1949_n N_noxref_16_c_2397_n ) capacitor c=0.0188655f \
 //x=16.685 //y=0.905 //x2=17.35 //y2=0.53
cc_1210 ( N_Q_c_1957_n N_noxref_16_c_2397_n ) capacitor c=0.00656458f \
 //x=17.215 //y=0.905 //x2=17.35 //y2=0.53
cc_1211 ( N_Q_c_1959_n N_noxref_16_c_2397_n ) capacitor c=2.1838e-19 //x=16.65 \
 //y=2.08 //x2=17.35 //y2=0.53
cc_1212 ( N_Q_c_1949_n N_noxref_16_M9_noxref_s ) capacitor c=0.00623646f \
 //x=16.685 //y=0.905 //x2=15.36 //y2=0.365
cc_1213 ( N_Q_c_1957_n N_noxref_16_M9_noxref_s ) capacitor c=0.0143002f \
 //x=17.215 //y=0.905 //x2=15.36 //y2=0.365
cc_1214 ( N_Q_c_1958_n N_noxref_16_M9_noxref_s ) capacitor c=0.00290153f \
 //x=17.215 //y=1.25 //x2=15.36 //y2=0.365
cc_1215 ( N_Q_c_2048_p N_noxref_17_c_2460_n ) capacitor c=3.15806e-19 \
 //x=20.365 //y=1.655 //x2=18.825 //y2=1.495
cc_1216 ( N_Q_c_1900_n N_noxref_17_c_2443_n ) capacitor c=0.00299723f \
 //x=20.605 //y=3.7 //x2=19.71 //y2=1.58
cc_1217 ( N_Q_c_1900_n N_noxref_17_c_2450_n ) capacitor c=0.00187232f \
 //x=20.605 //y=3.7 //x2=19.795 //y2=1.495
cc_1218 ( N_Q_c_2048_p N_noxref_17_c_2450_n ) capacitor c=0.0203424f \
 //x=20.365 //y=1.655 //x2=19.795 //y2=1.495
cc_1219 ( N_Q_c_1900_n N_noxref_17_c_2451_n ) capacitor c=4.7198e-19 \
 //x=20.605 //y=3.7 //x2=20.68 //y2=0.53
cc_1220 ( N_Q_c_1905_n N_noxref_17_c_2451_n ) capacitor c=0.00467104f \
 //x=20.635 //y=1.655 //x2=20.68 //y2=0.53
cc_1221 ( N_Q_M12_noxref_d N_noxref_17_c_2451_n ) capacitor c=0.0117932f \
 //x=20.09 //y=0.905 //x2=20.68 //y2=0.53
cc_1222 ( N_Q_c_1900_n N_noxref_17_M11_noxref_s ) capacitor c=3.61944e-19 \
 //x=20.605 //y=3.7 //x2=18.69 //y2=0.365
cc_1223 ( N_Q_c_1905_n N_noxref_17_M11_noxref_s ) capacitor c=0.0142774f \
 //x=20.635 //y=1.655 //x2=18.69 //y2=0.365
cc_1224 ( N_Q_M12_noxref_d N_noxref_17_M11_noxref_s ) capacitor c=0.043966f \
 //x=20.09 //y=0.905 //x2=18.69 //y2=0.365
cc_1225 ( N_noxref_10_c_2065_n N_noxref_11_c_2105_n ) capacitor c=0.0136048f \
 //x=2.445 //y=0.54 //x2=3.015 //y2=0.995
cc_1226 ( N_noxref_10_c_2076_n N_noxref_11_c_2105_n ) capacitor c=0.0102225f \
 //x=2.445 //y=1.59 //x2=3.015 //y2=0.995
cc_1227 ( N_noxref_10_M0_noxref_s N_noxref_11_c_2105_n ) capacitor \
 c=0.0228676f //x=0.455 //y=0.375 //x2=3.015 //y2=0.995
cc_1228 ( N_noxref_10_M0_noxref_s N_noxref_11_c_2107_n ) capacitor \
 c=0.0180035f //x=0.455 //y=0.375 //x2=3.1 //y2=0.625
cc_1229 ( N_noxref_10_c_2065_n N_noxref_11_M1_noxref_d ) capacitor \
 c=0.0129526f //x=2.445 //y=0.54 //x2=1.86 //y2=0.91
cc_1230 ( N_noxref_10_c_2076_n N_noxref_11_M1_noxref_d ) capacitor \
 c=0.00908243f //x=2.445 //y=1.59 //x2=1.86 //y2=0.91
cc_1231 ( N_noxref_10_M0_noxref_s N_noxref_11_M1_noxref_d ) capacitor \
 c=0.0159202f //x=0.455 //y=0.375 //x2=1.86 //y2=0.91
cc_1232 ( N_noxref_10_M0_noxref_s N_noxref_11_M2_noxref_s ) capacitor \
 c=0.0213553f //x=0.455 //y=0.375 //x2=2.965 //y2=0.375
cc_1233 ( N_noxref_11_c_2113_n N_noxref_13_M3_noxref_s ) capacitor \
 c=0.00164795f //x=4.07 //y=0.625 //x2=5.37 //y2=0.365
cc_1234 ( N_D_c_2179_n N_noxref_13_c_2238_n ) capacitor c=0.00623646f \
 //x=6.695 //y=1.56 //x2=6.475 //y2=1.495
cc_1235 ( N_D_c_2188_n N_noxref_13_c_2238_n ) capacitor c=0.00176439f //x=6.66 \
 //y=2.08 //x2=6.475 //y2=1.495
cc_1236 ( N_D_c_2158_n N_noxref_13_c_2239_n ) capacitor c=0.00159897f //x=6.66 \
 //y=2.08 //x2=7.36 //y2=0.53
cc_1237 ( N_D_c_2177_n N_noxref_13_c_2239_n ) capacitor c=0.0188655f //x=6.695 \
 //y=0.905 //x2=7.36 //y2=0.53
cc_1238 ( N_D_c_2185_n N_noxref_13_c_2239_n ) capacitor c=0.00656458f \
 //x=7.225 //y=0.905 //x2=7.36 //y2=0.53
cc_1239 ( N_D_c_2188_n N_noxref_13_c_2239_n ) capacitor c=2.1838e-19 //x=6.66 \
 //y=2.08 //x2=7.36 //y2=0.53
cc_1240 ( N_D_c_2177_n N_noxref_13_M3_noxref_s ) capacitor c=0.00623646f \
 //x=6.695 //y=0.905 //x2=5.37 //y2=0.365
cc_1241 ( N_D_c_2185_n N_noxref_13_M3_noxref_s ) capacitor c=0.0143002f \
 //x=7.225 //y=0.905 //x2=5.37 //y2=0.365
cc_1242 ( N_D_c_2186_n N_noxref_13_M3_noxref_s ) capacitor c=0.00290153f \
 //x=7.225 //y=1.25 //x2=5.37 //y2=0.365
cc_1243 ( N_noxref_13_c_2242_n N_noxref_14_M5_noxref_s ) capacitor \
 c=0.00174327f //x=7.445 //y=0.615 //x2=8.7 //y2=0.365
cc_1244 ( N_noxref_14_c_2294_n N_noxref_15_M7_noxref_s ) capacitor \
 c=0.00174327f //x=10.775 //y=0.615 //x2=12.03 //y2=0.365
cc_1245 ( N_noxref_15_c_2347_n N_noxref_16_M9_noxref_s ) capacitor \
 c=0.00174327f //x=14.105 //y=0.615 //x2=15.36 //y2=0.365
cc_1246 ( N_noxref_16_c_2400_n N_noxref_17_M11_noxref_s ) capacitor \
 c=0.00174327f //x=17.435 //y=0.615 //x2=18.69 //y2=0.365
