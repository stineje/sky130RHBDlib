* SPICE3 file created from AND3X1.ext - technology: sky130A

.subckt AND3X1 Y A B C VPB VNB
M1000 VPB.t7 a_147_159# a_277_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_1147_182.t2 a_277_1004.t7 VPB.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPB.t1 a_342_166# a_277_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VNB a_147_159# a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=1.3199p pd=9.67u as=0p ps=0u
M1004 VPB.t3 a_599_943# a_277_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_277_1004.t5 a_147_159# VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_277_1004.t1 a_342_166# VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPB.t4 a_277_1004.t9 a_1147_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_277_1004.t3 a_599_943# VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 a_599_943# a_342_166# 0.18fF
C1 VPB a_342_166# 0.05fF
C2 a_147_159# a_342_166# 0.18fF
C3 a_599_943# VPB 0.06fF
C4 a_599_943# a_147_159# 0.02fF
C5 VPB a_147_159# 0.08fF
R0 a_277_1004.n6 a_277_1004.t9 512.525
R1 a_277_1004.n6 a_277_1004.t7 371.139
R2 a_277_1004.n7 a_277_1004.t8 220.263
R3 a_277_1004.n10 a_277_1004.n8 196.598
R4 a_277_1004.n8 a_277_1004.n5 180.846
R5 a_277_1004.n7 a_277_1004.n6 158.3
R6 a_277_1004.n8 a_277_1004.n7 153.043
R7 a_277_1004.n4 a_277_1004.n3 79.232
R8 a_277_1004.n5 a_277_1004.n4 63.152
R9 a_277_1004.n10 a_277_1004.n9 30
R10 a_277_1004.n11 a_277_1004.n0 24.383
R11 a_277_1004.n11 a_277_1004.n10 23.684
R12 a_277_1004.n5 a_277_1004.n1 16.08
R13 a_277_1004.n4 a_277_1004.n2 16.08
R14 a_277_1004.n1 a_277_1004.t2 14.282
R15 a_277_1004.n1 a_277_1004.t3 14.282
R16 a_277_1004.n2 a_277_1004.t0 14.282
R17 a_277_1004.n2 a_277_1004.t1 14.282
R18 a_277_1004.n3 a_277_1004.t6 14.282
R19 a_277_1004.n3 a_277_1004.t5 14.282
R20 VPB VPB.n145 126.832
R21 VPB.n87 VPB.n85 94.117
R22 VPB.n122 VPB.n121 80.104
R23 VPB.n128 VPB.n127 76
R24 VPB.n138 VPB.n137 76
R25 VPB.n100 VPB.n99 75.654
R26 VPB.n77 VPB.n76 68.979
R27 VPB.n70 VPB.n69 64.528
R28 VPB.n29 VPB.n28 61.764
R29 VPB.n95 VPB.t6 55.106
R30 VPB.n80 VPB.t5 55.106
R31 VPB.n68 VPB.t4 55.106
R32 VPB.n92 VPB.t3 55.106
R33 VPB.n118 VPB.n117 48.952
R34 VPB.n104 VPB.n103 44.502
R35 VPB.n107 VPB.n94 40.824
R36 VPB.n116 VPB.n93 40.824
R37 VPB.n142 VPB.n138 20.452
R38 VPB.n67 VPB.n64 20.452
R39 VPB.n113 VPB.n112 17.801
R40 VPB.n94 VPB.t0 14.282
R41 VPB.n94 VPB.t7 14.282
R42 VPB.n93 VPB.t2 14.282
R43 VPB.n93 VPB.t1 14.282
R44 VPB.n67 VPB.n66 13.653
R45 VPB.n66 VPB.n65 13.653
R46 VPB.n72 VPB.n71 13.653
R47 VPB.n71 VPB.n70 13.653
R48 VPB.n75 VPB.n74 13.653
R49 VPB.n74 VPB.n73 13.653
R50 VPB.n79 VPB.n78 13.653
R51 VPB.n78 VPB.n77 13.653
R52 VPB.n83 VPB.n82 13.653
R53 VPB.n82 VPB.n81 13.653
R54 VPB.n88 VPB.n87 13.653
R55 VPB.n87 VPB.n86 13.653
R56 VPB.n91 VPB.n90 13.653
R57 VPB.n90 VPB.n89 13.653
R58 VPB.n127 VPB.n126 13.653
R59 VPB.n126 VPB.n125 13.653
R60 VPB.n124 VPB.n123 13.653
R61 VPB.n123 VPB.n122 13.653
R62 VPB.n120 VPB.n119 13.653
R63 VPB.n119 VPB.n118 13.653
R64 VPB.n115 VPB.n114 13.653
R65 VPB.n114 VPB.n113 13.653
R66 VPB.n111 VPB.n110 13.653
R67 VPB.n110 VPB.n109 13.653
R68 VPB.n106 VPB.n105 13.653
R69 VPB.n105 VPB.n104 13.653
R70 VPB.n102 VPB.n101 13.653
R71 VPB.n101 VPB.n100 13.653
R72 VPB.n98 VPB.n97 13.653
R73 VPB.n97 VPB.n96 13.653
R74 VPB.n16 VPB.n15 13.653
R75 VPB.n15 VPB.n14 13.653
R76 VPB.n138 VPB.n0 13.653
R77 VPB VPB.n0 13.653
R78 VPB.n109 VPB.n108 13.35
R79 VPB.n142 VPB.n141 13.276
R80 VPB.n141 VPB.n139 13.276
R81 VPB.n43 VPB.n25 13.276
R82 VPB.n25 VPB.n23 13.276
R83 VPB.n75 VPB.n72 13.276
R84 VPB.n79 VPB.n75 13.276
R85 VPB.n84 VPB.n83 13.276
R86 VPB.n88 VPB.n84 13.276
R87 VPB.n91 VPB.n88 13.276
R88 VPB.n127 VPB.n124 13.276
R89 VPB.n124 VPB.n120 13.276
R90 VPB.n115 VPB.n111 13.276
R91 VPB.n106 VPB.n102 13.276
R92 VPB.n102 VPB.n98 13.276
R93 VPB.n138 VPB.n16 13.276
R94 VPB.n64 VPB.n46 13.276
R95 VPB.n46 VPB.n44 13.276
R96 VPB.n51 VPB.n49 12.796
R97 VPB.n51 VPB.n50 12.564
R98 VPB.n95 VPB.n16 12.558
R99 VPB.n92 VPB.n91 12.2
R100 VPB.n59 VPB.n58 12.198
R101 VPB.n57 VPB.n56 12.198
R102 VPB.n54 VPB.n53 12.198
R103 VPB.n83 VPB.n80 10.944
R104 VPB.n68 VPB.n67 10.585
R105 VPB.n116 VPB.n115 9.329
R106 VPB.n111 VPB.n107 8.97
R107 VPB.n64 VPB.n63 7.5
R108 VPB.n49 VPB.n48 7.5
R109 VPB.n53 VPB.n52 7.5
R110 VPB.n56 VPB.n55 7.5
R111 VPB.n46 VPB.n45 7.5
R112 VPB.n61 VPB.n47 7.5
R113 VPB.n25 VPB.n24 7.5
R114 VPB.n38 VPB.n37 7.5
R115 VPB.n32 VPB.n31 7.5
R116 VPB.n34 VPB.n33 7.5
R117 VPB.n27 VPB.n26 7.5
R118 VPB.n43 VPB.n42 7.5
R119 VPB.n141 VPB.n140 7.5
R120 VPB.n12 VPB.n11 7.5
R121 VPB.n6 VPB.n5 7.5
R122 VPB.n8 VPB.n7 7.5
R123 VPB.n2 VPB.n1 7.5
R124 VPB.n143 VPB.n142 7.5
R125 VPB.n84 VPB.n43 7.176
R126 VPB.n39 VPB.n36 6.729
R127 VPB.n35 VPB.n32 6.729
R128 VPB.n30 VPB.n27 6.729
R129 VPB.n13 VPB.n10 6.729
R130 VPB.n9 VPB.n6 6.729
R131 VPB.n4 VPB.n2 6.729
R132 VPB.n30 VPB.n29 6.728
R133 VPB.n35 VPB.n34 6.728
R134 VPB.n39 VPB.n38 6.728
R135 VPB.n42 VPB.n41 6.728
R136 VPB.n4 VPB.n3 6.728
R137 VPB.n9 VPB.n8 6.728
R138 VPB.n13 VPB.n12 6.728
R139 VPB.n144 VPB.n143 6.728
R140 VPB.n63 VPB.n62 6.398
R141 VPB.n107 VPB.n106 4.305
R142 VPB.n120 VPB.n116 3.947
R143 VPB.n72 VPB.n68 2.691
R144 VPB.n80 VPB.n79 2.332
R145 VPB.n61 VPB.n54 1.402
R146 VPB.n61 VPB.n57 1.402
R147 VPB.n61 VPB.n59 1.402
R148 VPB.n61 VPB.n60 1.402
R149 VPB.n127 VPB.n92 1.076
R150 VPB.n62 VPB.n61 0.735
R151 VPB.n61 VPB.n51 0.735
R152 VPB.n98 VPB.n95 0.717
R153 VPB.n40 VPB.n39 0.387
R154 VPB.n40 VPB.n35 0.387
R155 VPB.n40 VPB.n30 0.387
R156 VPB.n41 VPB.n40 0.387
R157 VPB.n145 VPB.n13 0.387
R158 VPB.n145 VPB.n9 0.387
R159 VPB.n145 VPB.n4 0.387
R160 VPB.n145 VPB.n144 0.387
R161 VPB.n21 VPB.n20 0.272
R162 VPB.n137 VPB 0.198
R163 VPB.n18 VPB.n17 0.136
R164 VPB.n19 VPB.n18 0.136
R165 VPB.n20 VPB.n19 0.136
R166 VPB.n22 VPB.n21 0.136
R167 VPB.n128 VPB.n22 0.136
R168 VPB.n130 VPB.n129 0.136
R169 VPB.n131 VPB.n130 0.136
R170 VPB.n132 VPB.n131 0.136
R171 VPB.n133 VPB.n132 0.136
R172 VPB.n134 VPB.n133 0.136
R173 VPB.n135 VPB.n134 0.136
R174 VPB.n136 VPB.n135 0.136
R175 VPB.n137 VPB.n136 0.136
R176 VPB VPB.n128 0.068
R177 VPB.n129 VPB 0.068
R178 a_91_75.t0 a_91_75.n0 117.777
R179 a_91_75.n2 a_91_75.n1 55.228
R180 a_91_75.n4 a_91_75.n3 9.111
R181 a_91_75.n8 a_91_75.n6 7.859
R182 a_91_75.t0 a_91_75.n2 4.04
R183 a_91_75.t0 a_91_75.n8 3.034
R184 a_91_75.n6 a_91_75.n4 1.964
R185 a_91_75.n6 a_91_75.n5 1.964
R186 a_91_75.n8 a_91_75.n7 0.443
R187 a_372_182.n10 a_372_182.n8 82.852
R188 a_372_182.n11 a_372_182.n0 49.6
R189 a_372_182.n7 a_372_182.n6 32.833
R190 a_372_182.n8 a_372_182.t1 32.416
R191 a_372_182.n10 a_372_182.n9 27.2
R192 a_372_182.n3 a_372_182.n2 23.284
R193 a_372_182.n11 a_372_182.n10 22.4
R194 a_372_182.n7 a_372_182.n4 19.017
R195 a_372_182.n6 a_372_182.n5 13.494
R196 a_372_182.t1 a_372_182.n1 7.04
R197 a_372_182.t1 a_372_182.n3 5.727
R198 a_372_182.n8 a_372_182.n7 1.435
R199 a_1147_182.n3 a_1147_182.n1 355.848
R200 a_1147_182.n3 a_1147_182.n2 30
R201 a_1147_182.n4 a_1147_182.n0 24.383
R202 a_1147_182.n4 a_1147_182.n3 23.684
R203 a_1147_182.n1 a_1147_182.t1 14.282
R204 a_1147_182.n1 a_1147_182.t2 14.282
R205 VNB VNB.n130 300.778
R206 VNB.n23 VNB.n22 199.897
R207 VNB.n76 VNB.n74 154.509
R208 VNB.n82 VNB.n81 85.559
R209 VNB.n117 VNB.n116 76
R210 VNB.n107 VNB.n106 76
R211 VNB.n64 VNB.n63 49.896
R212 VNB.n84 VNB.n83 41.971
R213 VNB.n39 VNB.n38 35.01
R214 VNB.t0 VNB.n31 32.601
R215 VNB.n57 VNB.n54 20.452
R216 VNB.n118 VNB.n117 20.452
R217 VNB.n58 VNB.n39 20.094
R218 VNB.n62 VNB.n36 20.094
R219 VNB.n69 VNB.n34 20.094
R220 VNB.n39 VNB.n37 19.017
R221 VNB.n33 VNB.t0 17.353
R222 VNB.n61 VNB.n60 13.653
R223 VNB.n60 VNB.n59 13.653
R224 VNB.n65 VNB.n64 13.653
R225 VNB.n68 VNB.n67 13.653
R226 VNB.n67 VNB.n66 13.653
R227 VNB.n72 VNB.n71 13.653
R228 VNB.n71 VNB.n70 13.653
R229 VNB.n77 VNB.n76 13.653
R230 VNB.n76 VNB.n75 13.653
R231 VNB.n80 VNB.n79 13.653
R232 VNB.n79 VNB.n78 13.653
R233 VNB.n106 VNB.n105 13.653
R234 VNB.n105 VNB.n104 13.653
R235 VNB.n103 VNB.n102 13.653
R236 VNB.n102 VNB.n101 13.653
R237 VNB.n100 VNB.n99 13.653
R238 VNB.n99 VNB.n98 13.653
R239 VNB.n97 VNB.n96 13.653
R240 VNB.n96 VNB.n95 13.653
R241 VNB.n94 VNB.n93 13.653
R242 VNB.n93 VNB.n92 13.653
R243 VNB.n91 VNB.n90 13.653
R244 VNB.n90 VNB.n89 13.653
R245 VNB.n88 VNB.n87 13.653
R246 VNB.n87 VNB.n86 13.653
R247 VNB.n85 VNB.n84 13.653
R248 VNB.n6 VNB.n5 13.653
R249 VNB.n5 VNB.n4 13.653
R250 VNB.n117 VNB.n0 13.653
R251 VNB VNB.n0 13.653
R252 VNB.n57 VNB.n56 13.653
R253 VNB.n56 VNB.n55 13.653
R254 VNB.n125 VNB.n122 13.577
R255 VNB.n42 VNB.n40 13.276
R256 VNB.n54 VNB.n42 13.276
R257 VNB.n15 VNB.n13 13.276
R258 VNB.n28 VNB.n15 13.276
R259 VNB.n68 VNB.n65 13.276
R260 VNB.n73 VNB.n72 13.276
R261 VNB.n77 VNB.n73 13.276
R262 VNB.n80 VNB.n77 13.276
R263 VNB.n106 VNB.n80 13.276
R264 VNB.n106 VNB.n103 13.276
R265 VNB.n103 VNB.n100 13.276
R266 VNB.n100 VNB.n97 13.276
R267 VNB.n97 VNB.n94 13.276
R268 VNB.n94 VNB.n91 13.276
R269 VNB.n91 VNB.n88 13.276
R270 VNB.n88 VNB.n85 13.276
R271 VNB.n117 VNB.n6 13.276
R272 VNB.n3 VNB.n1 13.276
R273 VNB.n118 VNB.n3 13.276
R274 VNB.n62 VNB.n61 13.097
R275 VNB.n34 VNB.n33 12.837
R276 VNB.n82 VNB.n6 12.02
R277 VNB.n72 VNB.n69 9.329
R278 VNB.n58 VNB.n57 8.97
R279 VNB.n33 VNB.n32 7.566
R280 VNB.n127 VNB.n126 7.5
R281 VNB.n21 VNB.n20 7.5
R282 VNB.n17 VNB.n16 7.5
R283 VNB.n15 VNB.n14 7.5
R284 VNB.n28 VNB.n27 7.5
R285 VNB.n119 VNB.n118 7.5
R286 VNB.n3 VNB.n2 7.5
R287 VNB.n124 VNB.n123 7.5
R288 VNB.n48 VNB.n47 7.5
R289 VNB.n44 VNB.n43 7.5
R290 VNB.n42 VNB.n41 7.5
R291 VNB.n54 VNB.n53 7.5
R292 VNB.n73 VNB.n28 7.176
R293 VNB.n129 VNB.n127 7.011
R294 VNB.n24 VNB.n21 7.011
R295 VNB.n19 VNB.n17 7.011
R296 VNB.n50 VNB.n48 7.011
R297 VNB.n46 VNB.n44 7.011
R298 VNB.n27 VNB.n26 7.01
R299 VNB.n19 VNB.n18 7.01
R300 VNB.n24 VNB.n23 7.01
R301 VNB.n53 VNB.n52 7.01
R302 VNB.n46 VNB.n45 7.01
R303 VNB.n50 VNB.n49 7.01
R304 VNB.n129 VNB.n128 7.01
R305 VNB.n125 VNB.n124 6.788
R306 VNB.n120 VNB.n119 6.788
R307 VNB.n30 VNB.n29 4.551
R308 VNB.n61 VNB.n58 4.305
R309 VNB.n69 VNB.n68 3.947
R310 VNB.t0 VNB.n30 2.238
R311 VNB.n85 VNB.n82 1.255
R312 VNB.n130 VNB.n121 0.921
R313 VNB.n130 VNB.n125 0.476
R314 VNB.n130 VNB.n120 0.475
R315 VNB.n36 VNB.n35 0.358
R316 VNB.n11 VNB.n10 0.272
R317 VNB.n25 VNB.n19 0.246
R318 VNB.n26 VNB.n25 0.246
R319 VNB.n25 VNB.n24 0.246
R320 VNB.n51 VNB.n46 0.246
R321 VNB.n52 VNB.n51 0.246
R322 VNB.n51 VNB.n50 0.246
R323 VNB.n130 VNB.n129 0.246
R324 VNB.n116 VNB 0.198
R325 VNB.n65 VNB.n62 0.179
R326 VNB.n8 VNB.n7 0.136
R327 VNB.n9 VNB.n8 0.136
R328 VNB.n10 VNB.n9 0.136
R329 VNB.n12 VNB.n11 0.136
R330 VNB.n107 VNB.n12 0.136
R331 VNB.n109 VNB.n108 0.136
R332 VNB.n110 VNB.n109 0.136
R333 VNB.n111 VNB.n110 0.136
R334 VNB.n112 VNB.n111 0.136
R335 VNB.n113 VNB.n112 0.136
R336 VNB.n114 VNB.n113 0.136
R337 VNB.n115 VNB.n114 0.136
R338 VNB.n116 VNB.n115 0.136
R339 VNB VNB.n107 0.068
R340 VNB.n108 VNB 0.068
C6 VPB VNB 6.39fF
C7 a_1147_182.n0 VNB 0.04fF
C8 a_1147_182.n1 VNB 1.01fF
C9 a_1147_182.n2 VNB 0.04fF
C10 a_1147_182.n3 VNB 0.49fF
C11 a_1147_182.n4 VNB 0.06fF
C12 a_372_182.n0 VNB 0.02fF
C13 a_372_182.n1 VNB 0.09fF
C14 a_372_182.n2 VNB 0.13fF
C15 a_372_182.n3 VNB 0.11fF
C16 a_372_182.t1 VNB 0.30fF
C17 a_372_182.n4 VNB 0.09fF
C18 a_372_182.n5 VNB 0.06fF
C19 a_372_182.n6 VNB 0.01fF
C20 a_372_182.n7 VNB 0.03fF
C21 a_372_182.n8 VNB 0.11fF
C22 a_372_182.n9 VNB 0.02fF
C23 a_372_182.n10 VNB 0.05fF
C24 a_372_182.n11 VNB 0.02fF
C25 a_91_75.n0 VNB 0.03fF
C26 a_91_75.n1 VNB 0.10fF
C27 a_91_75.n2 VNB 0.10fF
C28 a_91_75.n3 VNB 0.04fF
C29 a_91_75.n4 VNB 0.03fF
C30 a_91_75.n5 VNB 0.03fF
C31 a_91_75.n6 VNB 0.11fF
C32 a_91_75.n7 VNB 0.04fF
C33 VPB.n0 VNB 0.03fF
C34 VPB.n1 VNB 0.03fF
C35 VPB.n2 VNB 0.02fF
C36 VPB.n3 VNB 0.17fF
C37 VPB.n5 VNB 0.02fF
C38 VPB.n6 VNB 0.02fF
C39 VPB.n7 VNB 0.02fF
C40 VPB.n8 VNB 0.02fF
C41 VPB.n10 VNB 0.02fF
C42 VPB.n11 VNB 0.02fF
C43 VPB.n12 VNB 0.02fF
C44 VPB.n14 VNB 0.25fF
C45 VPB.n15 VNB 0.02fF
C46 VPB.n16 VNB 0.02fF
C47 VPB.n17 VNB 0.07fF
C48 VPB.n18 VNB 0.02fF
C49 VPB.n19 VNB 0.02fF
C50 VPB.n20 VNB 0.03fF
C51 VPB.n21 VNB 0.03fF
C52 VPB.n22 VNB 0.02fF
C53 VPB.n23 VNB 0.02fF
C54 VPB.n24 VNB 0.02fF
C55 VPB.n25 VNB 0.02fF
C56 VPB.n26 VNB 0.03fF
C57 VPB.n27 VNB 0.02fF
C58 VPB.n28 VNB 0.20fF
C59 VPB.n29 VNB 0.04fF
C60 VPB.n31 VNB 0.02fF
C61 VPB.n32 VNB 0.02fF
C62 VPB.n33 VNB 0.02fF
C63 VPB.n34 VNB 0.02fF
C64 VPB.n36 VNB 0.02fF
C65 VPB.n37 VNB 0.02fF
C66 VPB.n38 VNB 0.02fF
C67 VPB.n40 VNB 0.25fF
C68 VPB.n42 VNB 0.02fF
C69 VPB.n43 VNB 0.02fF
C70 VPB.n44 VNB 0.02fF
C71 VPB.n45 VNB 0.02fF
C72 VPB.n46 VNB 0.02fF
C73 VPB.n47 VNB 0.10fF
C74 VPB.n48 VNB 0.02fF
C75 VPB.n49 VNB 0.02fF
C76 VPB.n50 VNB 0.04fF
C77 VPB.n51 VNB 0.01fF
C78 VPB.n52 VNB 0.02fF
C79 VPB.n53 VNB 0.02fF
C80 VPB.n55 VNB 0.02fF
C81 VPB.n56 VNB 0.02fF
C82 VPB.n58 VNB 0.02fF
C83 VPB.n61 VNB 0.42fF
C84 VPB.n63 VNB 0.03fF
C85 VPB.n64 VNB 0.03fF
C86 VPB.n65 VNB 0.25fF
C87 VPB.n66 VNB 0.03fF
C88 VPB.n67 VNB 0.03fF
C89 VPB.n68 VNB 0.05fF
C90 VPB.n69 VNB 0.12fF
C91 VPB.n70 VNB 0.17fF
C92 VPB.n71 VNB 0.02fF
C93 VPB.n72 VNB 0.01fF
C94 VPB.n73 VNB 0.15fF
C95 VPB.n74 VNB 0.02fF
C96 VPB.n75 VNB 0.02fF
C97 VPB.n76 VNB 0.12fF
C98 VPB.n77 VNB 0.18fF
C99 VPB.n78 VNB 0.02fF
C100 VPB.n79 VNB 0.01fF
C101 VPB.n80 VNB 0.05fF
C102 VPB.n81 VNB 0.25fF
C103 VPB.n82 VNB 0.01fF
C104 VPB.n83 VNB 0.02fF
C105 VPB.n84 VNB 0.03fF
C106 VPB.n85 VNB 0.03fF
C107 VPB.n86 VNB 0.25fF
C108 VPB.n87 VNB 0.01fF
C109 VPB.n88 VNB 0.02fF
C110 VPB.n89 VNB 0.25fF
C111 VPB.n90 VNB 0.02fF
C112 VPB.n91 VNB 0.02fF
C113 VPB.n92 VNB 0.05fF
C114 VPB.n93 VNB 0.09fF
C115 VPB.n94 VNB 0.09fF
C116 VPB.n95 VNB 0.05fF
C117 VPB.n96 VNB 0.19fF
C118 VPB.n97 VNB 0.02fF
C119 VPB.n98 VNB 0.01fF
C120 VPB.n99 VNB 0.12fF
C121 VPB.n100 VNB 0.15fF
C122 VPB.n101 VNB 0.02fF
C123 VPB.n102 VNB 0.02fF
C124 VPB.n103 VNB 0.12fF
C125 VPB.n104 VNB 0.15fF
C126 VPB.n105 VNB 0.02fF
C127 VPB.n106 VNB 0.01fF
C128 VPB.n107 VNB 0.02fF
C129 VPB.n108 VNB 0.12fF
C130 VPB.n109 VNB 0.13fF
C131 VPB.n110 VNB 0.02fF
C132 VPB.n111 VNB 0.02fF
C133 VPB.n112 VNB 0.12fF
C134 VPB.n113 VNB 0.14fF
C135 VPB.n114 VNB 0.02fF
C136 VPB.n115 VNB 0.02fF
C137 VPB.n116 VNB 0.02fF
C138 VPB.n117 VNB 0.12fF
C139 VPB.n118 VNB 0.15fF
C140 VPB.n119 VNB 0.02fF
C141 VPB.n120 VNB 0.01fF
C142 VPB.n121 VNB 0.12fF
C143 VPB.n122 VNB 0.15fF
C144 VPB.n123 VNB 0.02fF
C145 VPB.n124 VNB 0.02fF
C146 VPB.n125 VNB 0.19fF
C147 VPB.n126 VNB 0.02fF
C148 VPB.n127 VNB 0.01fF
C149 VPB.n128 VNB 0.02fF
C150 VPB.n129 VNB 0.02fF
C151 VPB.n130 VNB 0.02fF
C152 VPB.n131 VNB 0.02fF
C153 VPB.n132 VNB 0.02fF
C154 VPB.n133 VNB 0.02fF
C155 VPB.n134 VNB 0.02fF
C156 VPB.n135 VNB 0.02fF
C157 VPB.n136 VNB 0.02fF
C158 VPB.n137 VNB 0.03fF
C159 VPB.n138 VNB 0.03fF
C160 VPB.n139 VNB 0.02fF
C161 VPB.n140 VNB 0.02fF
C162 VPB.n141 VNB 0.02fF
C163 VPB.n142 VNB 0.03fF
C164 VPB.n143 VNB 0.03fF
C165 VPB.n145 VNB 0.39fF
C166 a_277_1004.n0 VNB 0.03fF
C167 a_277_1004.n1 VNB 0.39fF
C168 a_277_1004.n2 VNB 0.39fF
C169 a_277_1004.n3 VNB 0.46fF
C170 a_277_1004.n4 VNB 0.14fF
C171 a_277_1004.n5 VNB 0.23fF
C172 a_277_1004.n6 VNB 0.26fF
C173 a_277_1004.t8 VNB 0.38fF
C174 a_277_1004.n7 VNB 0.42fF
C175 a_277_1004.n8 VNB 0.43fF
C176 a_277_1004.n9 VNB 0.02fF
C177 a_277_1004.n10 VNB 0.20fF
C178 a_277_1004.n11 VNB 0.04fF
.ends
