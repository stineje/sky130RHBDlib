// File: OR3X1.spi.OR3X1.pxi
// Created: Tue Oct 15 15:50:55 2024
// 
simulator lang=spectre
x_PM_OR3X1\%noxref_1 ( N_noxref_1_c_4_p N_noxref_1_c_54_p N_noxref_1_c_14_p \
 N_noxref_1_c_15_p N_noxref_1_c_18_p N_noxref_1_c_19_p N_noxref_1_c_22_p \
 N_noxref_1_c_5_p N_noxref_1_c_6_p N_noxref_1_c_7_p N_noxref_1_c_36_p \
 N_noxref_1_c_1_p N_noxref_1_c_2_p N_noxref_1_c_3_p N_noxref_1_M0_noxref_s \
 N_noxref_1_M3_noxref_s )  PM_OR3X1\%noxref_1
x_PM_OR3X1\%noxref_2 ( N_noxref_2_c_92_p N_noxref_2_c_115_p N_noxref_2_c_89_n \
 N_noxref_2_c_118_p N_noxref_2_c_101_p N_noxref_2_c_90_n N_noxref_2_c_91_n \
 N_noxref_2_M4_noxref_d N_noxref_2_M10_noxref_s N_noxref_2_M11_noxref_d )  \
 PM_OR3X1\%noxref_2
x_PM_OR3X1\%noxref_3 ( N_noxref_3_c_170_n N_noxref_3_c_176_n \
 N_noxref_3_c_179_n N_noxref_3_c_238_p N_noxref_3_c_183_n N_noxref_3_c_187_n \
 N_noxref_3_c_223_n N_noxref_3_c_193_n N_noxref_3_c_291_p N_noxref_3_c_263_p \
 N_noxref_3_M3_noxref_g N_noxref_3_M10_noxref_g N_noxref_3_M11_noxref_g \
 N_noxref_3_c_198_n N_noxref_3_c_312_p N_noxref_3_c_313_p N_noxref_3_c_200_n \
 N_noxref_3_c_233_n N_noxref_3_c_234_n N_noxref_3_c_201_n N_noxref_3_c_304_p \
 N_noxref_3_c_202_n N_noxref_3_c_204_n N_noxref_3_c_205_n \
 N_noxref_3_M0_noxref_d N_noxref_3_M1_noxref_d N_noxref_3_M2_noxref_d \
 N_noxref_3_M8_noxref_d )  PM_OR3X1\%noxref_3
x_PM_OR3X1\%A ( A A A A A A A N_A_c_323_n N_A_c_335_n N_A_M0_noxref_g \
 N_A_M4_noxref_g N_A_M5_noxref_g N_A_c_326_n N_A_c_346_n N_A_c_347_n \
 N_A_c_328_n N_A_c_330_n N_A_c_351_n N_A_c_356_p N_A_c_331_n N_A_c_333_n \
 N_A_c_343_n )  PM_OR3X1\%A
x_PM_OR3X1\%B ( B B B B B B B N_B_c_413_n N_B_c_389_n N_B_M1_noxref_g \
 N_B_M6_noxref_g N_B_M7_noxref_g N_B_c_390_n N_B_c_402_n N_B_c_403_n \
 N_B_c_461_p N_B_c_392_n N_B_c_393_n N_B_c_394_n N_B_c_410_n N_B_c_411_n \
 N_B_c_412_n N_B_c_434_n )  PM_OR3X1\%B
x_PM_OR3X1\%noxref_6 ( N_noxref_6_c_469_n N_noxref_6_c_473_n \
 N_noxref_6_c_474_n N_noxref_6_c_476_n N_noxref_6_M4_noxref_s \
 N_noxref_6_M5_noxref_d N_noxref_6_M7_noxref_d )  PM_OR3X1\%noxref_6
x_PM_OR3X1\%C ( C C C C C C C N_C_c_515_n N_C_M2_noxref_g N_C_M8_noxref_g \
 N_C_M9_noxref_g N_C_c_517_n N_C_c_540_n N_C_c_541_n N_C_c_544_n N_C_c_519_n \
 N_C_c_520_n N_C_c_521_n N_C_c_551_n N_C_c_529_n N_C_c_523_n N_C_c_557_n )  \
 PM_OR3X1\%C
x_PM_OR3X1\%noxref_8 ( N_noxref_8_c_586_n N_noxref_8_c_589_n \
 N_noxref_8_c_590_n N_noxref_8_c_591_n N_noxref_8_M6_noxref_d \
 N_noxref_8_M8_noxref_s N_noxref_8_M9_noxref_d )  PM_OR3X1\%noxref_8
x_PM_OR3X1\%Y ( Y Y Y Y Y Y Y N_Y_c_629_n N_Y_c_653_n N_Y_c_639_n N_Y_c_642_n \
 N_Y_M3_noxref_d N_Y_M10_noxref_d )  PM_OR3X1\%Y
cc_1 ( N_noxref_1_c_1_p N_noxref_2_c_89_n ) capacitor c=0.00989031f //x=0.695 \
 //y=0 //x2=0.74 //y2=7.4
cc_2 ( N_noxref_1_c_2_p N_noxref_2_c_90_n ) capacitor c=0.00855708f //x=4.81 \
 //y=0 //x2=4.81 //y2=7.4
cc_3 ( N_noxref_1_c_3_p N_noxref_2_c_91_n ) capacitor c=0.00989031f //x=6.41 \
 //y=0 //x2=6.29 //y2=7.4
cc_4 ( N_noxref_1_c_4_p N_noxref_3_c_170_n ) capacitor c=0.014587f //x=6.29 \
 //y=0 //x2=5.435 //y2=3.33
cc_5 ( N_noxref_1_c_5_p N_noxref_3_c_170_n ) capacitor c=0.00301933f //x=4.64 \
 //y=0 //x2=5.435 //y2=3.33
cc_6 ( N_noxref_1_c_6_p N_noxref_3_c_170_n ) capacitor c=0.00110325f //x=5.355 \
 //y=0 //x2=5.435 //y2=3.33
cc_7 ( N_noxref_1_c_7_p N_noxref_3_c_170_n ) capacitor c=2.76195e-19 //x=5.84 \
 //y=0.535 //x2=5.435 //y2=3.33
cc_8 ( N_noxref_1_c_2_p N_noxref_3_c_170_n ) capacitor c=0.00820844f //x=4.81 \
 //y=0 //x2=5.435 //y2=3.33
cc_9 ( N_noxref_1_M3_noxref_s N_noxref_3_c_170_n ) capacitor c=0.00164577f \
 //x=5.305 //y=0.37 //x2=5.435 //y2=3.33
cc_10 ( N_noxref_1_c_4_p N_noxref_3_c_176_n ) capacitor c=0.00197108f //x=6.29 \
 //y=0 //x2=3.815 //y2=3.33
cc_11 ( N_noxref_1_c_5_p N_noxref_3_c_176_n ) capacitor c=2.24303e-19 //x=4.64 \
 //y=0 //x2=3.815 //y2=3.33
cc_12 ( N_noxref_1_M0_noxref_s N_noxref_3_c_176_n ) capacitor c=2.00237e-19 \
 //x=0.56 //y=0.365 //x2=3.815 //y2=3.33
cc_13 ( N_noxref_1_c_4_p N_noxref_3_c_179_n ) capacitor c=0.00359057f //x=6.29 \
 //y=0 //x2=2.065 //y2=1.655
cc_14 ( N_noxref_1_c_14_p N_noxref_3_c_179_n ) capacitor c=0.00381844f \
 //x=1.58 //y=0.53 //x2=2.065 //y2=1.655
cc_15 ( N_noxref_1_c_15_p N_noxref_3_c_179_n ) capacitor c=0.00323369f \
 //x=2.065 //y=0.53 //x2=2.065 //y2=1.655
cc_16 ( N_noxref_1_M0_noxref_s N_noxref_3_c_179_n ) capacitor c=0.0173679f \
 //x=0.56 //y=0.365 //x2=2.065 //y2=1.655
cc_17 ( N_noxref_1_c_4_p N_noxref_3_c_183_n ) capacitor c=0.00410159f //x=6.29 \
 //y=0 //x2=3.035 //y2=1.655
cc_18 ( N_noxref_1_c_18_p N_noxref_3_c_183_n ) capacitor c=0.00381844f \
 //x=2.55 //y=0.53 //x2=3.035 //y2=1.655
cc_19 ( N_noxref_1_c_19_p N_noxref_3_c_183_n ) capacitor c=0.00324961f \
 //x=3.035 //y=0.53 //x2=3.035 //y2=1.655
cc_20 ( N_noxref_1_M0_noxref_s N_noxref_3_c_183_n ) capacitor c=0.0175442f \
 //x=0.56 //y=0.365 //x2=3.035 //y2=1.655
cc_21 ( N_noxref_1_c_4_p N_noxref_3_c_187_n ) capacitor c=0.00337239f //x=6.29 \
 //y=0 //x2=3.615 //y2=1.655
cc_22 ( N_noxref_1_c_22_p N_noxref_3_c_187_n ) capacitor c=0.0047981f //x=3.52 \
 //y=0.53 //x2=3.615 //y2=1.655
cc_23 ( N_noxref_1_c_5_p N_noxref_3_c_187_n ) capacitor c=4.94729e-19 //x=4.64 \
 //y=0 //x2=3.615 //y2=1.655
cc_24 ( N_noxref_1_c_2_p N_noxref_3_c_187_n ) capacitor c=0.0293055f //x=4.81 \
 //y=0 //x2=3.615 //y2=1.655
cc_25 ( N_noxref_1_M0_noxref_s N_noxref_3_c_187_n ) capacitor c=0.020002f \
 //x=0.56 //y=0.365 //x2=3.615 //y2=1.655
cc_26 ( N_noxref_1_M3_noxref_s N_noxref_3_c_187_n ) capacitor c=2.64584e-19 \
 //x=5.305 //y=0.37 //x2=3.615 //y2=1.655
cc_27 ( N_noxref_1_c_4_p N_noxref_3_c_193_n ) capacitor c=0.00184963f //x=6.29 \
 //y=0 //x2=5.55 //y2=2.085
cc_28 ( N_noxref_1_c_7_p N_noxref_3_c_193_n ) capacitor c=7.87839e-19 //x=5.84 \
 //y=0.535 //x2=5.55 //y2=2.085
cc_29 ( N_noxref_1_c_2_p N_noxref_3_c_193_n ) capacitor c=0.029021f //x=4.81 \
 //y=0 //x2=5.55 //y2=2.085
cc_30 ( N_noxref_1_c_3_p N_noxref_3_c_193_n ) capacitor c=0.00118981f //x=6.41 \
 //y=0 //x2=5.55 //y2=2.085
cc_31 ( N_noxref_1_M3_noxref_s N_noxref_3_c_193_n ) capacitor c=0.0108503f \
 //x=5.305 //y=0.37 //x2=5.55 //y2=2.085
cc_32 ( N_noxref_1_c_7_p N_noxref_3_c_198_n ) capacitor c=0.0121757f //x=5.84 \
 //y=0.535 //x2=5.66 //y2=0.91
cc_33 ( N_noxref_1_M3_noxref_s N_noxref_3_c_198_n ) capacitor c=0.0317181f \
 //x=5.305 //y=0.37 //x2=5.66 //y2=0.91
cc_34 ( N_noxref_1_c_2_p N_noxref_3_c_200_n ) capacitor c=0.0107331f //x=4.81 \
 //y=0 //x2=5.66 //y2=1.92
cc_35 ( N_noxref_1_M3_noxref_s N_noxref_3_c_201_n ) capacitor c=0.00483274f \
 //x=5.305 //y=0.37 //x2=6.035 //y2=0.755
cc_36 ( N_noxref_1_c_36_p N_noxref_3_c_202_n ) capacitor c=0.0118602f \
 //x=6.325 //y=0.535 //x2=6.19 //y2=0.91
cc_37 ( N_noxref_1_M3_noxref_s N_noxref_3_c_202_n ) capacitor c=0.0143355f \
 //x=5.305 //y=0.37 //x2=6.19 //y2=0.91
cc_38 ( N_noxref_1_M3_noxref_s N_noxref_3_c_204_n ) capacitor c=0.0074042f \
 //x=5.305 //y=0.37 //x2=6.19 //y2=1.255
cc_39 ( N_noxref_1_c_7_p N_noxref_3_c_205_n ) capacitor c=2.1838e-19 //x=5.84 \
 //y=0.535 //x2=5.55 //y2=2.085
cc_40 ( N_noxref_1_c_2_p N_noxref_3_c_205_n ) capacitor c=0.0108179f //x=4.81 \
 //y=0 //x2=5.55 //y2=2.085
cc_41 ( N_noxref_1_M3_noxref_s N_noxref_3_c_205_n ) capacitor c=0.00655738f \
 //x=5.305 //y=0.37 //x2=5.55 //y2=2.085
cc_42 ( N_noxref_1_c_4_p N_noxref_3_M0_noxref_d ) capacitor c=0.00175924f \
 //x=6.29 //y=0 //x2=0.99 //y2=0.905
cc_43 ( N_noxref_1_c_1_p N_noxref_3_M0_noxref_d ) capacitor c=0.00419389f \
 //x=0.695 //y=0 //x2=0.99 //y2=0.905
cc_44 ( N_noxref_1_c_3_p N_noxref_3_M0_noxref_d ) capacitor c=2.31043e-19 \
 //x=6.41 //y=0 //x2=0.99 //y2=0.905
cc_45 ( N_noxref_1_M0_noxref_s N_noxref_3_M0_noxref_d ) capacitor c=0.0775691f \
 //x=0.56 //y=0.365 //x2=0.99 //y2=0.905
cc_46 ( N_noxref_1_c_4_p N_noxref_3_M1_noxref_d ) capacitor c=0.00195394f \
 //x=6.29 //y=0 //x2=1.96 //y2=0.905
cc_47 ( N_noxref_1_c_3_p N_noxref_3_M1_noxref_d ) capacitor c=2.31043e-19 \
 //x=6.41 //y=0 //x2=1.96 //y2=0.905
cc_48 ( N_noxref_1_M0_noxref_s N_noxref_3_M1_noxref_d ) capacitor c=0.0610444f \
 //x=0.56 //y=0.365 //x2=1.96 //y2=0.905
cc_49 ( N_noxref_1_c_4_p N_noxref_3_M2_noxref_d ) capacitor c=0.00193447f \
 //x=6.29 //y=0 //x2=2.93 //y2=0.905
cc_50 ( N_noxref_1_c_2_p N_noxref_3_M2_noxref_d ) capacitor c=0.00374104f \
 //x=4.81 //y=0 //x2=2.93 //y2=0.905
cc_51 ( N_noxref_1_c_3_p N_noxref_3_M2_noxref_d ) capacitor c=2.31043e-19 \
 //x=6.41 //y=0 //x2=2.93 //y2=0.905
cc_52 ( N_noxref_1_M0_noxref_s N_noxref_3_M2_noxref_d ) capacitor c=0.0604189f \
 //x=0.56 //y=0.365 //x2=2.93 //y2=0.905
cc_53 ( N_noxref_1_c_4_p N_A_c_323_n ) capacitor c=6.7762e-19 //x=6.29 //y=0 \
 //x2=1.11 //y2=2.08
cc_54 ( N_noxref_1_c_54_p N_A_c_323_n ) capacitor c=0.00136072f //x=1.095 \
 //y=0.53 //x2=1.11 //y2=2.08
cc_55 ( N_noxref_1_c_1_p N_A_c_323_n ) capacitor c=0.0176887f //x=0.695 //y=0 \
 //x2=1.11 //y2=2.08
cc_56 ( N_noxref_1_c_54_p N_A_c_326_n ) capacitor c=0.0122371f //x=1.095 \
 //y=0.53 //x2=0.915 //y2=0.905
cc_57 ( N_noxref_1_M0_noxref_s N_A_c_326_n ) capacitor c=0.0318083f //x=0.56 \
 //y=0.365 //x2=0.915 //y2=0.905
cc_58 ( N_noxref_1_c_54_p N_A_c_328_n ) capacitor c=2.1838e-19 //x=1.095 \
 //y=0.53 //x2=0.915 //y2=1.915
cc_59 ( N_noxref_1_c_1_p N_A_c_328_n ) capacitor c=0.0198857f //x=0.695 //y=0 \
 //x2=0.915 //y2=1.915
cc_60 ( N_noxref_1_M0_noxref_s N_A_c_330_n ) capacitor c=0.00474433f //x=0.56 \
 //y=0.365 //x2=1.29 //y2=0.75
cc_61 ( N_noxref_1_c_14_p N_A_c_331_n ) capacitor c=0.0113089f //x=1.58 \
 //y=0.53 //x2=1.445 //y2=0.905
cc_62 ( N_noxref_1_M0_noxref_s N_A_c_331_n ) capacitor c=0.00514143f //x=0.56 \
 //y=0.365 //x2=1.445 //y2=0.905
cc_63 ( N_noxref_1_M0_noxref_s N_A_c_333_n ) capacitor c=8.33128e-19 //x=0.56 \
 //y=0.365 //x2=1.445 //y2=1.25
cc_64 ( N_noxref_1_c_1_p N_B_c_389_n ) capacitor c=9.2064e-19 //x=0.695 //y=0 \
 //x2=1.85 //y2=2.08
cc_65 ( N_noxref_1_c_15_p N_B_c_390_n ) capacitor c=0.01113f //x=2.065 \
 //y=0.53 //x2=1.885 //y2=0.905
cc_66 ( N_noxref_1_M0_noxref_s N_B_c_390_n ) capacitor c=0.00590563f //x=0.56 \
 //y=0.365 //x2=1.885 //y2=0.905
cc_67 ( N_noxref_1_M0_noxref_s N_B_c_392_n ) capacitor c=0.00481727f //x=0.56 \
 //y=0.365 //x2=2.26 //y2=0.75
cc_68 ( N_noxref_1_M0_noxref_s N_B_c_393_n ) capacitor c=8.38882e-19 //x=0.56 \
 //y=0.365 //x2=2.26 //y2=1.405
cc_69 ( N_noxref_1_c_18_p N_B_c_394_n ) capacitor c=0.0113819f //x=2.55 \
 //y=0.53 //x2=2.415 //y2=0.905
cc_70 ( N_noxref_1_M0_noxref_s N_B_c_394_n ) capacitor c=0.00513762f //x=0.56 \
 //y=0.365 //x2=2.415 //y2=0.905
cc_71 ( N_noxref_1_c_4_p N_C_c_515_n ) capacitor c=3.7166e-19 //x=6.29 //y=0 \
 //x2=2.96 //y2=2.08
cc_72 ( N_noxref_1_c_2_p N_C_c_515_n ) capacitor c=5.99091e-19 //x=4.81 //y=0 \
 //x2=2.96 //y2=2.08
cc_73 ( N_noxref_1_c_19_p N_C_c_517_n ) capacitor c=0.0108358f //x=3.035 \
 //y=0.53 //x2=2.855 //y2=0.905
cc_74 ( N_noxref_1_M0_noxref_s N_C_c_517_n ) capacitor c=0.00590563f //x=0.56 \
 //y=0.365 //x2=2.855 //y2=0.905
cc_75 ( N_noxref_1_M0_noxref_s N_C_c_519_n ) capacitor c=0.00452306f //x=0.56 \
 //y=0.365 //x2=3.23 //y2=0.75
cc_76 ( N_noxref_1_M0_noxref_s N_C_c_520_n ) capacitor c=0.00316186f //x=0.56 \
 //y=0.365 //x2=3.23 //y2=1.405
cc_77 ( N_noxref_1_c_22_p N_C_c_521_n ) capacitor c=0.0110876f //x=3.52 \
 //y=0.53 //x2=3.385 //y2=0.905
cc_78 ( N_noxref_1_M0_noxref_s N_C_c_521_n ) capacitor c=0.0132184f //x=0.56 \
 //y=0.365 //x2=3.385 //y2=0.905
cc_79 ( N_noxref_1_c_19_p N_C_c_523_n ) capacitor c=2.26024e-19 //x=3.035 \
 //y=0.53 //x2=2.855 //y2=2.08
cc_80 ( N_noxref_1_c_2_p Y ) capacitor c=8.10282e-19 //x=4.81 //y=0 //x2=6.29 \
 //y2=2.22
cc_81 ( N_noxref_1_c_4_p N_Y_c_629_n ) capacitor c=0.00180637f //x=6.29 //y=0 \
 //x2=6.205 //y2=2.08
cc_82 ( N_noxref_1_c_3_p N_Y_c_629_n ) capacitor c=0.0301661f //x=6.41 //y=0 \
 //x2=6.205 //y2=2.08
cc_83 ( N_noxref_1_M3_noxref_s N_Y_c_629_n ) capacitor c=0.00999304f //x=5.305 \
 //y=0.37 //x2=6.205 //y2=2.08
cc_84 ( N_noxref_1_c_4_p N_Y_M3_noxref_d ) capacitor c=0.00194883f //x=6.29 \
 //y=0 //x2=5.735 //y2=0.91
cc_85 ( N_noxref_1_c_7_p N_Y_M3_noxref_d ) capacitor c=0.0146043f //x=5.84 \
 //y=0.535 //x2=5.735 //y2=0.91
cc_86 ( N_noxref_1_c_2_p N_Y_M3_noxref_d ) capacitor c=0.00924905f //x=4.81 \
 //y=0 //x2=5.735 //y2=0.91
cc_87 ( N_noxref_1_c_3_p N_Y_M3_noxref_d ) capacitor c=0.00973758f //x=6.41 \
 //y=0 //x2=5.735 //y2=0.91
cc_88 ( N_noxref_1_M3_noxref_s N_Y_M3_noxref_d ) capacitor c=0.076995f \
 //x=5.305 //y=0.37 //x2=5.735 //y2=0.91
cc_89 ( N_noxref_2_c_92_p N_noxref_3_c_170_n ) capacitor c=0.0112494f //x=6.29 \
 //y=7.4 //x2=5.435 //y2=3.33
cc_90 ( N_noxref_2_c_90_n N_noxref_3_c_170_n ) capacitor c=0.0069465f //x=4.81 \
 //y=7.4 //x2=5.435 //y2=3.33
cc_91 ( N_noxref_2_M10_noxref_s N_noxref_3_c_170_n ) capacitor c=0.00106085f \
 //x=5.35 //y=5.02 //x2=5.435 //y2=3.33
cc_92 ( N_noxref_2_c_92_p N_noxref_3_c_176_n ) capacitor c=0.00139969f \
 //x=6.29 //y=7.4 //x2=3.815 //y2=3.33
cc_93 ( N_noxref_2_c_90_n N_noxref_3_c_223_n ) capacitor c=0.0262421f //x=4.81 \
 //y=7.4 //x2=3.7 //y2=3.33
cc_94 ( N_noxref_2_c_92_p N_noxref_3_c_193_n ) capacitor c=0.00160122f \
 //x=6.29 //y=7.4 //x2=5.55 //y2=2.085
cc_95 ( N_noxref_2_c_90_n N_noxref_3_c_193_n ) capacitor c=0.0272885f //x=4.81 \
 //y=7.4 //x2=5.55 //y2=2.085
cc_96 ( N_noxref_2_c_91_n N_noxref_3_c_193_n ) capacitor c=0.00144809f \
 //x=6.29 //y=7.4 //x2=5.55 //y2=2.085
cc_97 ( N_noxref_2_M10_noxref_s N_noxref_3_c_193_n ) capacitor c=0.00971593f \
 //x=5.35 //y=5.02 //x2=5.55 //y2=2.085
cc_98 ( N_noxref_2_c_101_p N_noxref_3_M10_noxref_g ) capacitor c=0.00748034f \
 //x=6.28 //y=7.4 //x2=5.705 //y2=6.02
cc_99 ( N_noxref_2_c_90_n N_noxref_3_M10_noxref_g ) capacitor c=0.0102569f \
 //x=4.81 //y=7.4 //x2=5.705 //y2=6.02
cc_100 ( N_noxref_2_M10_noxref_s N_noxref_3_M10_noxref_g ) capacitor \
 c=0.0528676f //x=5.35 //y=5.02 //x2=5.705 //y2=6.02
cc_101 ( N_noxref_2_c_101_p N_noxref_3_M11_noxref_g ) capacitor c=0.00697478f \
 //x=6.28 //y=7.4 //x2=6.145 //y2=6.02
cc_102 ( N_noxref_2_M11_noxref_d N_noxref_3_M11_noxref_g ) capacitor \
 c=0.0528676f //x=6.22 //y=5.02 //x2=6.145 //y2=6.02
cc_103 ( N_noxref_2_c_91_n N_noxref_3_c_233_n ) capacitor c=0.0287802f \
 //x=6.29 //y=7.4 //x2=6.07 //y2=4.79
cc_104 ( N_noxref_2_c_90_n N_noxref_3_c_234_n ) capacitor c=0.011132f //x=4.81 \
 //y=7.4 //x2=5.78 //y2=4.79
cc_105 ( N_noxref_2_M10_noxref_s N_noxref_3_c_234_n ) capacitor c=0.00527247f \
 //x=5.35 //y=5.02 //x2=5.78 //y2=4.79
cc_106 ( N_noxref_2_c_90_n N_noxref_3_M8_noxref_d ) capacitor c=0.00966019f \
 //x=4.81 //y=7.4 //x2=3.445 //y2=5.025
cc_107 ( N_noxref_2_M10_noxref_s N_noxref_3_M8_noxref_d ) capacitor \
 c=4.94992e-19 //x=5.35 //y=5.02 //x2=3.445 //y2=5.025
cc_108 ( N_noxref_2_c_89_n N_A_c_323_n ) capacitor c=0.0104719f //x=0.74 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_109 ( N_noxref_2_c_92_p N_A_c_335_n ) capacitor c=3.36335e-19 //x=6.29 \
 //y=7.4 //x2=0.955 //y2=4.705
cc_110 ( N_noxref_2_c_89_n N_A_c_335_n ) capacitor c=0.008636f //x=0.74 \
 //y=7.4 //x2=0.955 //y2=4.705
cc_111 ( N_noxref_2_M4_noxref_d N_A_c_335_n ) capacitor c=2.82936e-19 \
 //x=1.085 //y=5.025 //x2=0.955 //y2=4.705
cc_112 ( N_noxref_2_c_115_p N_A_M4_noxref_g ) capacitor c=0.0067918f //x=1.145 \
 //y=7.4 //x2=1.01 //y2=6.025
cc_113 ( N_noxref_2_c_89_n N_A_M4_noxref_g ) capacitor c=0.0241979f //x=0.74 \
 //y=7.4 //x2=1.01 //y2=6.025
cc_114 ( N_noxref_2_M4_noxref_d N_A_M4_noxref_g ) capacitor c=0.0156786f \
 //x=1.085 //y=5.025 //x2=1.01 //y2=6.025
cc_115 ( N_noxref_2_c_118_p N_A_M5_noxref_g ) capacitor c=0.00678153f //x=4.64 \
 //y=7.4 //x2=1.45 //y2=6.025
cc_116 ( N_noxref_2_M4_noxref_d N_A_M5_noxref_g ) capacitor c=0.019067f \
 //x=1.085 //y=5.025 //x2=1.45 //y2=6.025
cc_117 ( N_noxref_2_c_89_n N_A_c_343_n ) capacitor c=0.00890932f //x=0.74 \
 //y=7.4 //x2=0.955 //y2=4.705
cc_118 ( N_noxref_2_c_89_n N_B_c_389_n ) capacitor c=7.02327e-19 //x=0.74 \
 //y=7.4 //x2=1.85 //y2=2.08
cc_119 ( N_noxref_2_c_118_p N_B_M6_noxref_g ) capacitor c=0.00513565f //x=4.64 \
 //y=7.4 //x2=1.89 //y2=6.025
cc_120 ( N_noxref_2_c_118_p N_B_M7_noxref_g ) capacitor c=0.00512552f //x=4.64 \
 //y=7.4 //x2=2.33 //y2=6.025
cc_121 ( N_noxref_2_c_92_p N_noxref_6_c_469_n ) capacitor c=0.00568164f \
 //x=6.29 //y=7.4 //x2=1.585 //y2=5.21
cc_122 ( N_noxref_2_c_115_p N_noxref_6_c_469_n ) capacitor c=4.37585e-19 \
 //x=1.145 //y=7.4 //x2=1.585 //y2=5.21
cc_123 ( N_noxref_2_c_118_p N_noxref_6_c_469_n ) capacitor c=4.37585e-19 \
 //x=4.64 //y=7.4 //x2=1.585 //y2=5.21
cc_124 ( N_noxref_2_M4_noxref_d N_noxref_6_c_469_n ) capacitor c=0.0130894f \
 //x=1.085 //y=5.025 //x2=1.585 //y2=5.21
cc_125 ( N_noxref_2_c_89_n N_noxref_6_c_473_n ) capacitor c=0.0679103f \
 //x=0.74 //y=7.4 //x2=0.875 //y2=5.21
cc_126 ( N_noxref_2_c_90_n N_noxref_6_c_474_n ) capacitor c=7.99339e-19 \
 //x=4.81 //y=7.4 //x2=2.465 //y2=6.91
cc_127 ( N_noxref_2_c_91_n N_noxref_6_c_474_n ) capacitor c=0.00358655f \
 //x=6.29 //y=7.4 //x2=2.465 //y2=6.91
cc_128 ( N_noxref_2_c_92_p N_noxref_6_c_476_n ) capacitor c=0.0367751f \
 //x=6.29 //y=7.4 //x2=1.755 //y2=6.91
cc_129 ( N_noxref_2_c_118_p N_noxref_6_c_476_n ) capacitor c=0.0586904f \
 //x=4.64 //y=7.4 //x2=1.755 //y2=6.91
cc_130 ( N_noxref_2_c_91_n N_noxref_6_c_476_n ) capacitor c=0.00118659f \
 //x=6.29 //y=7.4 //x2=1.755 //y2=6.91
cc_131 ( N_noxref_2_c_92_p N_noxref_6_M4_noxref_s ) capacitor c=0.00712902f \
 //x=6.29 //y=7.4 //x2=0.655 //y2=5.025
cc_132 ( N_noxref_2_c_115_p N_noxref_6_M4_noxref_s ) capacitor c=0.0141117f \
 //x=1.145 //y=7.4 //x2=0.655 //y2=5.025
cc_133 ( N_noxref_2_c_91_n N_noxref_6_M4_noxref_s ) capacitor c=0.00138926f \
 //x=6.29 //y=7.4 //x2=0.655 //y2=5.025
cc_134 ( N_noxref_2_M4_noxref_d N_noxref_6_M4_noxref_s ) capacitor \
 c=0.0667777f //x=1.085 //y=5.025 //x2=0.655 //y2=5.025
cc_135 ( N_noxref_2_c_89_n N_noxref_6_M5_noxref_d ) capacitor c=8.88629e-19 \
 //x=0.74 //y=7.4 //x2=1.525 //y2=5.025
cc_136 ( N_noxref_2_M4_noxref_d N_noxref_6_M5_noxref_d ) capacitor \
 c=0.0659925f //x=1.085 //y=5.025 //x2=1.525 //y2=5.025
cc_137 ( N_noxref_2_M4_noxref_d N_noxref_6_M7_noxref_d ) capacitor \
 c=0.00107819f //x=1.085 //y=5.025 //x2=2.405 //y2=5.025
cc_138 ( N_noxref_2_c_92_p N_C_c_515_n ) capacitor c=2.78723e-19 //x=6.29 \
 //y=7.4 //x2=2.96 //y2=2.08
cc_139 ( N_noxref_2_c_90_n N_C_c_515_n ) capacitor c=7.00707e-19 //x=4.81 \
 //y=7.4 //x2=2.96 //y2=2.08
cc_140 ( N_noxref_2_c_118_p N_C_M8_noxref_g ) capacitor c=0.00512552f //x=4.64 \
 //y=7.4 //x2=3.37 //y2=6.025
cc_141 ( N_noxref_2_c_118_p N_C_M9_noxref_g ) capacitor c=0.00512552f //x=4.64 \
 //y=7.4 //x2=3.81 //y2=6.025
cc_142 ( N_noxref_2_c_90_n N_C_M9_noxref_g ) capacitor c=0.00342488f //x=4.81 \
 //y=7.4 //x2=3.81 //y2=6.025
cc_143 ( N_noxref_2_c_90_n N_C_c_529_n ) capacitor c=0.0155316f //x=4.81 \
 //y=7.4 //x2=3.735 //y2=4.795
cc_144 ( N_noxref_2_c_92_p N_noxref_8_c_586_n ) capacitor c=0.00436737f \
 //x=6.29 //y=7.4 //x2=3.065 //y2=5.21
cc_145 ( N_noxref_2_c_118_p N_noxref_8_c_586_n ) capacitor c=0.00311573f \
 //x=4.64 //y=7.4 //x2=3.065 //y2=5.21
cc_146 ( N_noxref_2_c_90_n N_noxref_8_c_586_n ) capacitor c=0.00275857f \
 //x=4.81 //y=7.4 //x2=3.065 //y2=5.21
cc_147 ( N_noxref_2_c_89_n N_noxref_8_c_589_n ) capacitor c=9.33216e-19 \
 //x=0.74 //y=7.4 //x2=2.195 //y2=5.21
cc_148 ( N_noxref_2_c_91_n N_noxref_8_c_590_n ) capacitor c=0.00358655f \
 //x=6.29 //y=7.4 //x2=3.945 //y2=6.91
cc_149 ( N_noxref_2_c_92_p N_noxref_8_c_591_n ) capacitor c=0.0327433f \
 //x=6.29 //y=7.4 //x2=3.235 //y2=6.91
cc_150 ( N_noxref_2_c_118_p N_noxref_8_c_591_n ) capacitor c=0.0585561f \
 //x=4.64 //y=7.4 //x2=3.235 //y2=6.91
cc_151 ( N_noxref_2_c_91_n N_noxref_8_c_591_n ) capacitor c=0.00118659f \
 //x=6.29 //y=7.4 //x2=3.235 //y2=6.91
cc_152 ( N_noxref_2_M4_noxref_d N_noxref_8_c_591_n ) capacitor c=9.25055e-19 \
 //x=1.085 //y=5.025 //x2=3.235 //y2=6.91
cc_153 ( N_noxref_2_M4_noxref_d N_noxref_8_M6_noxref_d ) capacitor \
 c=0.00561178f //x=1.085 //y=5.025 //x2=1.965 //y2=5.025
cc_154 ( N_noxref_2_c_90_n N_noxref_8_M9_noxref_d ) capacitor c=0.0520312f \
 //x=4.81 //y=7.4 //x2=3.885 //y2=5.025
cc_155 ( N_noxref_2_M10_noxref_s N_noxref_8_M9_noxref_d ) capacitor \
 c=0.00226909f //x=5.35 //y=5.02 //x2=3.885 //y2=5.025
cc_156 ( N_noxref_2_c_90_n Y ) capacitor c=4.80934e-19 //x=4.81 //y=7.4 \
 //x2=6.29 //y2=2.22
cc_157 ( N_noxref_2_c_91_n Y ) capacitor c=0.0232778f //x=6.29 //y=7.4 \
 //x2=6.29 //y2=2.22
cc_158 ( N_noxref_2_c_92_p N_Y_c_639_n ) capacitor c=0.00190861f //x=6.29 \
 //y=7.4 //x2=6.205 //y2=4.58
cc_159 ( N_noxref_2_c_101_p N_Y_c_639_n ) capacitor c=8.8179e-19 //x=6.28 \
 //y=7.4 //x2=6.205 //y2=4.58
cc_160 ( N_noxref_2_M11_noxref_d N_Y_c_639_n ) capacitor c=0.00641434f \
 //x=6.22 //y=5.02 //x2=6.205 //y2=4.58
cc_161 ( N_noxref_2_c_90_n N_Y_c_642_n ) capacitor c=0.017572f //x=4.81 \
 //y=7.4 //x2=6.01 //y2=4.58
cc_162 ( N_noxref_2_c_92_p N_Y_M10_noxref_d ) capacitor c=0.00708604f //x=6.29 \
 //y=7.4 //x2=5.78 //y2=5.02
cc_163 ( N_noxref_2_c_101_p N_Y_M10_noxref_d ) capacitor c=0.0139004f //x=6.28 \
 //y=7.4 //x2=5.78 //y2=5.02
cc_164 ( N_noxref_2_c_91_n N_Y_M10_noxref_d ) capacitor c=0.0219131f //x=6.29 \
 //y=7.4 //x2=5.78 //y2=5.02
cc_165 ( N_noxref_2_M10_noxref_s N_Y_M10_noxref_d ) capacitor c=0.0843065f \
 //x=5.35 //y=5.02 //x2=5.78 //y2=5.02
cc_166 ( N_noxref_2_M11_noxref_d N_Y_M10_noxref_d ) capacitor c=0.0832641f \
 //x=6.22 //y=5.02 //x2=5.78 //y2=5.02
cc_167 ( N_noxref_3_c_238_p N_A_c_323_n ) capacitor c=0.0112169f //x=1.265 \
 //y=1.655 //x2=1.11 //y2=2.08
cc_168 ( N_noxref_3_M0_noxref_d N_A_c_326_n ) capacitor c=0.0013184f //x=0.99 \
 //y=0.905 //x2=0.915 //y2=0.905
cc_169 ( N_noxref_3_M0_noxref_d N_A_c_346_n ) capacitor c=0.0034598f //x=0.99 \
 //y=0.905 //x2=0.915 //y2=1.25
cc_170 ( N_noxref_3_M0_noxref_d N_A_c_347_n ) capacitor c=0.00300148f //x=0.99 \
 //y=0.905 //x2=0.915 //y2=1.56
cc_171 ( N_noxref_3_c_238_p N_A_c_328_n ) capacitor c=0.00589082f //x=1.265 \
 //y=1.655 //x2=0.915 //y2=1.915
cc_172 ( N_noxref_3_M0_noxref_d N_A_c_328_n ) capacitor c=0.00274546f //x=0.99 \
 //y=0.905 //x2=0.915 //y2=1.915
cc_173 ( N_noxref_3_M0_noxref_d N_A_c_330_n ) capacitor c=0.00241102f //x=0.99 \
 //y=0.905 //x2=1.29 //y2=0.75
cc_174 ( N_noxref_3_M0_noxref_d N_A_c_351_n ) capacitor c=0.0123304f //x=0.99 \
 //y=0.905 //x2=1.29 //y2=1.405
cc_175 ( N_noxref_3_M0_noxref_d N_A_c_331_n ) capacitor c=0.00219619f //x=0.99 \
 //y=0.905 //x2=1.445 //y2=0.905
cc_176 ( N_noxref_3_c_179_n N_A_c_333_n ) capacitor c=0.00431513f //x=2.065 \
 //y=1.655 //x2=1.445 //y2=1.25
cc_177 ( N_noxref_3_M0_noxref_d N_A_c_333_n ) capacitor c=0.00603828f //x=0.99 \
 //y=0.905 //x2=1.445 //y2=1.25
cc_178 ( N_noxref_3_c_179_n N_B_c_389_n ) capacitor c=0.0162392f //x=2.065 \
 //y=1.655 //x2=1.85 //y2=2.08
cc_179 ( N_noxref_3_c_223_n N_B_c_389_n ) capacitor c=0.00270493f //x=3.7 \
 //y=3.33 //x2=1.85 //y2=2.08
cc_180 ( N_noxref_3_M1_noxref_d N_B_c_390_n ) capacitor c=0.00132426f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=0.905
cc_181 ( N_noxref_3_M1_noxref_d N_B_c_402_n ) capacitor c=0.0035101f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=1.255
cc_182 ( N_noxref_3_c_179_n N_B_c_403_n ) capacitor c=0.00158038f //x=2.065 \
 //y=1.655 //x2=1.885 //y2=1.56
cc_183 ( N_noxref_3_M0_noxref_d N_B_c_403_n ) capacitor c=8.74435e-19 //x=0.99 \
 //y=0.905 //x2=1.885 //y2=1.56
cc_184 ( N_noxref_3_M1_noxref_d N_B_c_403_n ) capacitor c=0.00297998f //x=1.96 \
 //y=0.905 //x2=1.885 //y2=1.56
cc_185 ( N_noxref_3_M1_noxref_d N_B_c_392_n ) capacitor c=0.00241102f //x=1.96 \
 //y=0.905 //x2=2.26 //y2=0.75
cc_186 ( N_noxref_3_c_183_n N_B_c_393_n ) capacitor c=0.00430135f //x=3.035 \
 //y=1.655 //x2=2.26 //y2=1.405
cc_187 ( N_noxref_3_M1_noxref_d N_B_c_393_n ) capacitor c=0.0154425f //x=1.96 \
 //y=0.905 //x2=2.26 //y2=1.405
cc_188 ( N_noxref_3_M1_noxref_d N_B_c_394_n ) capacitor c=0.00132831f //x=1.96 \
 //y=0.905 //x2=2.415 //y2=0.905
cc_189 ( N_noxref_3_M1_noxref_d N_B_c_410_n ) capacitor c=0.0035101f //x=1.96 \
 //y=0.905 //x2=2.415 //y2=1.255
cc_190 ( N_noxref_3_c_179_n N_B_c_411_n ) capacitor c=0.00633758f //x=2.065 \
 //y=1.655 //x2=1.85 //y2=2.08
cc_191 ( N_noxref_3_c_179_n N_B_c_412_n ) capacitor c=0.0185539f //x=2.065 \
 //y=1.655 //x2=1.85 //y2=1.915
cc_192 ( N_noxref_3_c_263_p N_noxref_6_c_469_n ) capacitor c=0.00108534f \
 //x=3.7 //y=5.21 //x2=1.585 //y2=5.21
cc_193 ( N_noxref_3_M8_noxref_d N_noxref_6_M7_noxref_d ) capacitor \
 c=0.0049951f //x=3.445 //y=5.025 //x2=2.405 //y2=5.025
cc_194 ( N_noxref_3_c_176_n N_C_c_515_n ) capacitor c=0.00720056f //x=3.815 \
 //y=3.33 //x2=2.96 //y2=2.08
cc_195 ( N_noxref_3_c_183_n N_C_c_515_n ) capacitor c=0.0182656f //x=3.035 \
 //y=1.655 //x2=2.96 //y2=2.08
cc_196 ( N_noxref_3_c_223_n N_C_c_515_n ) capacitor c=0.0909072f //x=3.7 \
 //y=3.33 //x2=2.96 //y2=2.08
cc_197 ( N_noxref_3_c_193_n N_C_c_515_n ) capacitor c=0.00118081f //x=5.55 \
 //y=2.085 //x2=2.96 //y2=2.08
cc_198 ( N_noxref_3_c_223_n N_C_M8_noxref_g ) capacitor c=0.0059988f //x=3.7 \
 //y=3.33 //x2=3.37 //y2=6.025
cc_199 ( N_noxref_3_c_263_p N_C_M8_noxref_g ) capacitor c=0.0132317f //x=3.7 \
 //y=5.21 //x2=3.37 //y2=6.025
cc_200 ( N_noxref_3_c_223_n N_C_M9_noxref_g ) capacitor c=0.0066533f //x=3.7 \
 //y=3.33 //x2=3.81 //y2=6.025
cc_201 ( N_noxref_3_c_263_p N_C_M9_noxref_g ) capacitor c=0.00775053f //x=3.7 \
 //y=5.21 //x2=3.81 //y2=6.025
cc_202 ( N_noxref_3_M8_noxref_d N_C_M9_noxref_g ) capacitor c=0.0136385f \
 //x=3.445 //y=5.025 //x2=3.81 //y2=6.025
cc_203 ( N_noxref_3_M2_noxref_d N_C_c_517_n ) capacitor c=0.00226395f //x=2.93 \
 //y=0.905 //x2=2.855 //y2=0.905
cc_204 ( N_noxref_3_M2_noxref_d N_C_c_540_n ) capacitor c=0.0035101f //x=2.93 \
 //y=0.905 //x2=2.855 //y2=1.255
cc_205 ( N_noxref_3_c_183_n N_C_c_541_n ) capacitor c=0.0013609f //x=3.035 \
 //y=1.655 //x2=2.855 //y2=1.56
cc_206 ( N_noxref_3_M1_noxref_d N_C_c_541_n ) capacitor c=0.00148728f //x=1.96 \
 //y=0.905 //x2=2.855 //y2=1.56
cc_207 ( N_noxref_3_M2_noxref_d N_C_c_541_n ) capacitor c=0.00484362f //x=2.93 \
 //y=0.905 //x2=2.855 //y2=1.56
cc_208 ( N_noxref_3_c_183_n N_C_c_544_n ) capacitor c=0.0216105f //x=3.035 \
 //y=1.655 //x2=2.855 //y2=1.915
cc_209 ( N_noxref_3_c_223_n N_C_c_544_n ) capacitor c=0.00278932f //x=3.7 \
 //y=3.33 //x2=2.855 //y2=1.915
cc_210 ( N_noxref_3_M2_noxref_d N_C_c_544_n ) capacitor c=3.4952e-19 //x=2.93 \
 //y=0.905 //x2=2.855 //y2=1.915
cc_211 ( N_noxref_3_M2_noxref_d N_C_c_519_n ) capacitor c=0.00241102f //x=2.93 \
 //y=0.905 //x2=3.23 //y2=0.75
cc_212 ( N_noxref_3_c_187_n N_C_c_520_n ) capacitor c=0.00777513f //x=3.615 \
 //y=1.655 //x2=3.23 //y2=1.405
cc_213 ( N_noxref_3_M2_noxref_d N_C_c_520_n ) capacitor c=0.0156879f //x=2.93 \
 //y=0.905 //x2=3.23 //y2=1.405
cc_214 ( N_noxref_3_M2_noxref_d N_C_c_521_n ) capacitor c=0.00132831f //x=2.93 \
 //y=0.905 //x2=3.385 //y2=0.905
cc_215 ( N_noxref_3_M2_noxref_d N_C_c_551_n ) capacitor c=0.0035101f //x=2.93 \
 //y=0.905 //x2=3.385 //y2=1.255
cc_216 ( N_noxref_3_c_223_n N_C_c_529_n ) capacitor c=0.0150293f //x=3.7 \
 //y=3.33 //x2=3.735 //y2=4.795
cc_217 ( N_noxref_3_c_263_p N_C_c_529_n ) capacitor c=0.00302595f //x=3.7 \
 //y=5.21 //x2=3.735 //y2=4.795
cc_218 ( N_noxref_3_c_183_n N_C_c_523_n ) capacitor c=0.003666f //x=3.035 \
 //y=1.655 //x2=2.855 //y2=2.08
cc_219 ( N_noxref_3_c_223_n N_C_c_523_n ) capacitor c=0.00882918f //x=3.7 \
 //y=3.33 //x2=2.855 //y2=2.08
cc_220 ( N_noxref_3_c_291_p N_C_c_523_n ) capacitor c=0.00470847f //x=3.12 \
 //y=1.655 //x2=2.855 //y2=2.08
cc_221 ( N_noxref_3_c_223_n N_C_c_557_n ) capacitor c=0.00513934f //x=3.7 \
 //y=3.33 //x2=2.96 //y2=4.705
cc_222 ( N_noxref_3_c_263_p N_noxref_8_c_586_n ) capacitor c=0.0344081f \
 //x=3.7 //y=5.21 //x2=3.065 //y2=5.21
cc_223 ( N_noxref_3_c_263_p N_noxref_8_c_590_n ) capacitor c=0.00113815f \
 //x=3.7 //y=5.21 //x2=3.945 //y2=6.91
cc_224 ( N_noxref_3_M8_noxref_d N_noxref_8_c_590_n ) capacitor c=0.011849f \
 //x=3.445 //y=5.025 //x2=3.945 //y2=6.91
cc_225 ( N_noxref_3_M8_noxref_d N_noxref_8_M6_noxref_d ) capacitor \
 c=0.00101354f //x=3.445 //y=5.025 //x2=1.965 //y2=5.025
cc_226 ( N_noxref_3_M8_noxref_d N_noxref_8_M8_noxref_s ) capacitor \
 c=0.0344081f //x=3.445 //y=5.025 //x2=3.015 //y2=5.025
cc_227 ( N_noxref_3_c_170_n N_noxref_8_M9_noxref_d ) capacitor c=0.00131309f \
 //x=5.435 //y=3.33 //x2=3.885 //y2=5.025
cc_228 ( N_noxref_3_M8_noxref_d N_noxref_8_M9_noxref_d ) capacitor \
 c=0.0458293f //x=3.445 //y=5.025 //x2=3.885 //y2=5.025
cc_229 ( N_noxref_3_c_170_n Y ) capacitor c=0.00584488f //x=5.435 //y=3.33 \
 //x2=6.29 //y2=2.22
cc_230 ( N_noxref_3_c_223_n Y ) capacitor c=0.00118081f //x=3.7 //y=3.33 \
 //x2=6.29 //y2=2.22
cc_231 ( N_noxref_3_c_193_n Y ) capacitor c=0.0711303f //x=5.55 //y=2.085 \
 //x2=6.29 //y2=2.22
cc_232 ( N_noxref_3_c_205_n Y ) capacitor c=8.49451e-19 //x=5.55 //y=2.085 \
 //x2=6.29 //y2=2.22
cc_233 ( N_noxref_3_c_304_p N_Y_c_629_n ) capacitor c=0.0023507f //x=6.035 \
 //y=1.41 //x2=6.205 //y2=2.08
cc_234 ( N_noxref_3_c_205_n N_Y_c_653_n ) capacitor c=0.0167852f //x=5.55 \
 //y=2.085 //x2=6.005 //y2=2.08
cc_235 ( N_noxref_3_c_233_n N_Y_c_639_n ) capacitor c=0.0101013f //x=6.07 \
 //y=4.79 //x2=6.205 //y2=4.58
cc_236 ( N_noxref_3_c_193_n N_Y_c_642_n ) capacitor c=0.0250789f //x=5.55 \
 //y=2.085 //x2=6.01 //y2=4.58
cc_237 ( N_noxref_3_c_234_n N_Y_c_642_n ) capacitor c=0.00962086f //x=5.78 \
 //y=4.79 //x2=6.01 //y2=4.58
cc_238 ( N_noxref_3_c_223_n N_Y_M3_noxref_d ) capacitor c=2.60259e-19 //x=3.7 \
 //y=3.33 //x2=5.735 //y2=0.91
cc_239 ( N_noxref_3_c_193_n N_Y_M3_noxref_d ) capacitor c=0.0175773f //x=5.55 \
 //y=2.085 //x2=5.735 //y2=0.91
cc_240 ( N_noxref_3_c_198_n N_Y_M3_noxref_d ) capacitor c=0.00218556f //x=5.66 \
 //y=0.91 //x2=5.735 //y2=0.91
cc_241 ( N_noxref_3_c_312_p N_Y_M3_noxref_d ) capacitor c=0.00347355f //x=5.66 \
 //y=1.255 //x2=5.735 //y2=0.91
cc_242 ( N_noxref_3_c_313_p N_Y_M3_noxref_d ) capacitor c=0.00742431f //x=5.66 \
 //y=1.565 //x2=5.735 //y2=0.91
cc_243 ( N_noxref_3_c_200_n N_Y_M3_noxref_d ) capacitor c=0.00957707f //x=5.66 \
 //y=1.92 //x2=5.735 //y2=0.91
cc_244 ( N_noxref_3_c_201_n N_Y_M3_noxref_d ) capacitor c=0.00220879f \
 //x=6.035 //y=0.755 //x2=5.735 //y2=0.91
cc_245 ( N_noxref_3_c_304_p N_Y_M3_noxref_d ) capacitor c=0.0138447f //x=6.035 \
 //y=1.41 //x2=5.735 //y2=0.91
cc_246 ( N_noxref_3_c_202_n N_Y_M3_noxref_d ) capacitor c=0.00218624f //x=6.19 \
 //y=0.91 //x2=5.735 //y2=0.91
cc_247 ( N_noxref_3_c_204_n N_Y_M3_noxref_d ) capacitor c=0.00601286f //x=6.19 \
 //y=1.255 //x2=5.735 //y2=0.91
cc_248 ( N_noxref_3_M10_noxref_g N_Y_M10_noxref_d ) capacitor c=0.0219309f \
 //x=5.705 //y=6.02 //x2=5.78 //y2=5.02
cc_249 ( N_noxref_3_M11_noxref_g N_Y_M10_noxref_d ) capacitor c=0.021902f \
 //x=6.145 //y=6.02 //x2=5.78 //y2=5.02
cc_250 ( N_noxref_3_c_233_n N_Y_M10_noxref_d ) capacitor c=0.0148755f //x=6.07 \
 //y=4.79 //x2=5.78 //y2=5.02
cc_251 ( N_noxref_3_c_234_n N_Y_M10_noxref_d ) capacitor c=0.00307344f \
 //x=5.78 //y=4.79 //x2=5.78 //y2=5.02
cc_252 ( N_A_c_335_n N_B_c_413_n ) capacitor c=0.0481157f //x=0.955 //y=4.705 \
 //x2=1.85 //y2=4.54
cc_253 ( N_A_c_356_p N_B_c_413_n ) capacitor c=0.00146509f //x=1.375 //y=4.795 \
 //x2=1.85 //y2=4.54
cc_254 ( N_A_c_343_n N_B_c_413_n ) capacitor c=0.00112871f //x=0.955 //y=4.705 \
 //x2=1.85 //y2=4.54
cc_255 ( N_A_c_323_n N_B_c_389_n ) capacitor c=0.0453706f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=2.08
cc_256 ( N_A_c_328_n N_B_c_389_n ) capacitor c=0.00308814f //x=0.915 //y=1.915 \
 //x2=1.85 //y2=2.08
cc_257 ( N_A_M4_noxref_g N_B_M6_noxref_g ) capacitor c=0.0100243f //x=1.01 \
 //y=6.025 //x2=1.89 //y2=6.025
cc_258 ( N_A_M5_noxref_g N_B_M6_noxref_g ) capacitor c=0.107798f //x=1.45 \
 //y=6.025 //x2=1.89 //y2=6.025
cc_259 ( N_A_M5_noxref_g N_B_M7_noxref_g ) capacitor c=0.0094155f //x=1.45 \
 //y=6.025 //x2=2.33 //y2=6.025
cc_260 ( N_A_c_326_n N_B_c_390_n ) capacitor c=0.00125788f //x=0.915 //y=0.905 \
 //x2=1.885 //y2=0.905
cc_261 ( N_A_c_331_n N_B_c_390_n ) capacitor c=0.0126654f //x=1.445 //y=0.905 \
 //x2=1.885 //y2=0.905
cc_262 ( N_A_c_346_n N_B_c_402_n ) capacitor c=0.00148539f //x=0.915 //y=1.25 \
 //x2=1.885 //y2=1.255
cc_263 ( N_A_c_347_n N_B_c_402_n ) capacitor c=0.00105591f //x=0.915 //y=1.56 \
 //x2=1.885 //y2=1.255
cc_264 ( N_A_c_333_n N_B_c_402_n ) capacitor c=0.0126654f //x=1.445 //y=1.25 \
 //x2=1.885 //y2=1.255
cc_265 ( N_A_c_347_n N_B_c_403_n ) capacitor c=0.00109549f //x=0.915 //y=1.56 \
 //x2=1.885 //y2=1.56
cc_266 ( N_A_c_333_n N_B_c_403_n ) capacitor c=0.00886999f //x=1.445 //y=1.25 \
 //x2=1.885 //y2=1.56
cc_267 ( N_A_c_333_n N_B_c_393_n ) capacitor c=0.00123863f //x=1.445 //y=1.25 \
 //x2=2.26 //y2=1.405
cc_268 ( N_A_c_331_n N_B_c_394_n ) capacitor c=0.00132934f //x=1.445 //y=0.905 \
 //x2=2.415 //y2=0.905
cc_269 ( N_A_c_333_n N_B_c_410_n ) capacitor c=0.00150734f //x=1.445 //y=1.25 \
 //x2=2.415 //y2=1.255
cc_270 ( N_A_c_323_n N_B_c_411_n ) capacitor c=0.00307062f //x=1.11 //y=2.08 \
 //x2=1.85 //y2=2.08
cc_271 ( N_A_c_328_n N_B_c_411_n ) capacitor c=0.0176046f //x=0.915 //y=1.915 \
 //x2=1.85 //y2=2.08
cc_272 ( N_A_c_328_n N_B_c_412_n ) capacitor c=0.00577193f //x=0.915 //y=1.915 \
 //x2=1.85 //y2=1.915
cc_273 ( N_A_c_335_n N_B_c_434_n ) capacitor c=0.00336963f //x=0.955 //y=4.705 \
 //x2=1.885 //y2=4.705
cc_274 ( N_A_c_356_p N_B_c_434_n ) capacitor c=0.0197705f //x=1.375 //y=4.795 \
 //x2=1.885 //y2=4.705
cc_275 ( N_A_c_343_n N_B_c_434_n ) capacitor c=0.00546725f //x=0.955 //y=4.705 \
 //x2=1.885 //y2=4.705
cc_276 ( N_A_c_335_n N_noxref_6_c_469_n ) capacitor c=0.00628365f //x=0.955 \
 //y=4.705 //x2=1.585 //y2=5.21
cc_277 ( N_A_M4_noxref_g N_noxref_6_c_469_n ) capacitor c=0.0182391f //x=1.01 \
 //y=6.025 //x2=1.585 //y2=5.21
cc_278 ( N_A_M5_noxref_g N_noxref_6_c_469_n ) capacitor c=0.0203804f //x=1.45 \
 //y=6.025 //x2=1.585 //y2=5.21
cc_279 ( N_A_c_356_p N_noxref_6_c_469_n ) capacitor c=0.00343485f //x=1.375 \
 //y=4.795 //x2=1.585 //y2=5.21
cc_280 ( N_A_c_343_n N_noxref_6_c_469_n ) capacitor c=0.0017421f //x=0.955 \
 //y=4.705 //x2=1.585 //y2=5.21
cc_281 ( N_A_c_335_n N_noxref_6_c_473_n ) capacitor c=0.0120346f //x=0.955 \
 //y=4.705 //x2=0.875 //y2=5.21
cc_282 ( N_A_c_343_n N_noxref_6_c_473_n ) capacitor c=0.00518332f //x=0.955 \
 //y=4.705 //x2=0.875 //y2=5.21
cc_283 ( N_A_M4_noxref_g N_noxref_6_M4_noxref_s ) capacitor c=0.0473218f \
 //x=1.01 //y=6.025 //x2=0.655 //y2=5.025
cc_284 ( N_A_M5_noxref_g N_noxref_6_M5_noxref_d ) capacitor c=0.0170604f \
 //x=1.45 //y=6.025 //x2=1.525 //y2=5.025
cc_285 ( N_A_c_323_n N_C_c_515_n ) capacitor c=0.00247242f //x=1.11 //y=2.08 \
 //x2=2.96 //y2=2.08
cc_286 ( N_B_M6_noxref_g N_noxref_6_c_469_n ) capacitor c=0.0170604f //x=1.89 \
 //y=6.025 //x2=1.585 //y2=5.21
cc_287 ( N_B_c_434_n N_noxref_6_c_469_n ) capacitor c=2.24869e-19 //x=1.885 \
 //y=4.705 //x2=1.585 //y2=5.21
cc_288 ( N_B_c_413_n N_noxref_6_c_474_n ) capacitor c=8.92402e-19 //x=1.85 \
 //y=4.54 //x2=2.465 //y2=6.91
cc_289 ( N_B_M6_noxref_g N_noxref_6_c_474_n ) capacitor c=0.0148484f //x=1.89 \
 //y=6.025 //x2=2.465 //y2=6.91
cc_290 ( N_B_M7_noxref_g N_noxref_6_c_474_n ) capacitor c=0.0160244f //x=2.33 \
 //y=6.025 //x2=2.465 //y2=6.91
cc_291 ( N_B_M7_noxref_g N_noxref_6_M7_noxref_d ) capacitor c=0.0216879f \
 //x=2.33 //y=6.025 //x2=2.405 //y2=5.025
cc_292 ( N_B_c_413_n N_C_c_515_n ) capacitor c=0.00562297f //x=1.85 //y=4.54 \
 //x2=2.96 //y2=2.08
cc_293 ( N_B_c_389_n N_C_c_515_n ) capacitor c=0.0530421f //x=1.85 //y=2.08 \
 //x2=2.96 //y2=2.08
cc_294 ( N_B_c_411_n N_C_c_515_n ) capacitor c=3.80079e-19 //x=1.85 //y=2.08 \
 //x2=2.96 //y2=2.08
cc_295 ( N_B_c_434_n N_C_c_515_n ) capacitor c=4.01223e-19 //x=1.885 //y=4.705 \
 //x2=2.96 //y2=2.08
cc_296 ( N_B_M7_noxref_g N_C_M8_noxref_g ) capacitor c=0.0343614f //x=2.33 \
 //y=6.025 //x2=3.37 //y2=6.025
cc_297 ( N_B_c_390_n N_C_c_517_n ) capacitor c=0.00131574f //x=1.885 //y=0.905 \
 //x2=2.855 //y2=0.905
cc_298 ( N_B_c_394_n N_C_c_517_n ) capacitor c=0.00886682f //x=2.415 //y=0.905 \
 //x2=2.855 //y2=0.905
cc_299 ( N_B_c_402_n N_C_c_540_n ) capacitor c=0.00150456f //x=1.885 //y=1.255 \
 //x2=2.855 //y2=1.255
cc_300 ( N_B_c_410_n N_C_c_540_n ) capacitor c=0.00886682f //x=2.415 //y=1.255 \
 //x2=2.855 //y2=1.255
cc_301 ( N_B_c_403_n N_C_c_541_n ) capacitor c=0.00276257f //x=1.885 //y=1.56 \
 //x2=2.855 //y2=1.56
cc_302 ( N_B_c_393_n N_C_c_541_n ) capacitor c=0.0177628f //x=2.26 //y=1.405 \
 //x2=2.855 //y2=1.56
cc_303 ( N_B_c_412_n N_C_c_544_n ) capacitor c=0.00494016f //x=1.85 //y=1.915 \
 //x2=2.855 //y2=1.915
cc_304 ( N_B_c_393_n N_C_c_520_n ) capacitor c=0.00123863f //x=2.26 //y=1.405 \
 //x2=3.23 //y2=1.405
cc_305 ( N_B_c_394_n N_C_c_521_n ) capacitor c=0.00132934f //x=2.415 //y=0.905 \
 //x2=3.385 //y2=0.905
cc_306 ( N_B_c_410_n N_C_c_551_n ) capacitor c=0.00150456f //x=2.415 //y=1.255 \
 //x2=3.385 //y2=1.255
cc_307 ( N_B_c_389_n N_C_c_523_n ) capacitor c=0.00235136f //x=1.85 //y=2.08 \
 //x2=2.855 //y2=2.08
cc_308 ( N_B_c_411_n N_C_c_523_n ) capacitor c=0.00922588f //x=1.85 //y=2.08 \
 //x2=2.855 //y2=2.08
cc_309 ( N_B_c_413_n N_C_c_557_n ) capacitor c=0.00227279f //x=1.85 //y=4.54 \
 //x2=2.96 //y2=4.705
cc_310 ( N_B_c_461_p N_C_c_557_n ) capacitor c=0.0106154f //x=2.255 //y=4.795 \
 //x2=2.96 //y2=4.705
cc_311 ( N_B_c_434_n N_C_c_557_n ) capacitor c=0.00510965f //x=1.885 //y=4.705 \
 //x2=2.96 //y2=4.705
cc_312 ( N_B_M7_noxref_g N_noxref_8_c_586_n ) capacitor c=0.0222373f //x=2.33 \
 //y=6.025 //x2=3.065 //y2=5.21
cc_313 ( N_B_M6_noxref_g N_noxref_8_c_589_n ) capacitor c=0.0132989f //x=1.89 \
 //y=6.025 //x2=2.195 //y2=5.21
cc_314 ( N_B_c_461_p N_noxref_8_c_589_n ) capacitor c=0.00410596f //x=2.255 \
 //y=4.795 //x2=2.195 //y2=5.21
cc_315 ( N_B_M7_noxref_g N_noxref_8_c_591_n ) capacitor c=0.00102459f //x=2.33 \
 //y=6.025 //x2=3.235 //y2=6.91
cc_316 ( N_B_M7_noxref_g N_noxref_8_M6_noxref_d ) capacitor c=0.0134276f \
 //x=2.33 //y=6.025 //x2=1.965 //y2=5.025
cc_317 ( N_B_M7_noxref_g N_noxref_8_M8_noxref_s ) capacitor c=0.00207713f \
 //x=2.33 //y=6.025 //x2=3.015 //y2=5.025
cc_318 ( N_noxref_6_c_474_n N_C_M8_noxref_g ) capacitor c=0.00102459f \
 //x=2.465 //y=6.91 //x2=3.37 //y2=6.025
cc_319 ( N_noxref_6_c_474_n N_noxref_8_c_586_n ) capacitor c=0.00112299f \
 //x=2.465 //y=6.91 //x2=3.065 //y2=5.21
cc_320 ( N_noxref_6_M7_noxref_d N_noxref_8_c_586_n ) capacitor c=0.0129087f \
 //x=2.405 //y=5.025 //x2=3.065 //y2=5.21
cc_321 ( N_noxref_6_c_469_n N_noxref_8_c_589_n ) capacitor c=0.0351721f \
 //x=1.585 //y=5.21 //x2=2.195 //y2=5.21
cc_322 ( N_noxref_6_c_474_n N_noxref_8_c_591_n ) capacitor c=0.027433f \
 //x=2.465 //y=6.91 //x2=3.235 //y2=6.91
cc_323 ( N_noxref_6_c_474_n N_noxref_8_M6_noxref_d ) capacitor c=0.0118172f \
 //x=2.465 //y=6.91 //x2=1.965 //y2=5.025
cc_324 ( N_noxref_6_M4_noxref_s N_noxref_8_M6_noxref_d ) capacitor \
 c=0.00107541f //x=0.655 //y=5.025 //x2=1.965 //y2=5.025
cc_325 ( N_noxref_6_M5_noxref_d N_noxref_8_M6_noxref_d ) capacitor \
 c=0.0351721f //x=1.525 //y=5.025 //x2=1.965 //y2=5.025
cc_326 ( N_noxref_6_M7_noxref_d N_noxref_8_M6_noxref_d ) capacitor \
 c=0.0458293f //x=2.405 //y=5.025 //x2=1.965 //y2=5.025
cc_327 ( N_noxref_6_M5_noxref_d N_noxref_8_M8_noxref_s ) capacitor \
 c=0.00194853f //x=1.525 //y=5.025 //x2=3.015 //y2=5.025
cc_328 ( N_noxref_6_M7_noxref_d N_noxref_8_M8_noxref_s ) capacitor c=0.027433f \
 //x=2.405 //y=5.025 //x2=3.015 //y2=5.025
cc_329 ( N_noxref_6_M7_noxref_d N_noxref_8_M9_noxref_d ) capacitor \
 c=9.17547e-19 //x=2.405 //y=5.025 //x2=3.885 //y2=5.025
cc_330 ( N_C_c_515_n N_noxref_8_c_586_n ) capacitor c=0.012085f //x=2.96 \
 //y=2.08 //x2=3.065 //y2=5.21
cc_331 ( N_C_M8_noxref_g N_noxref_8_c_586_n ) capacitor c=0.0286624f //x=3.37 \
 //y=6.025 //x2=3.065 //y2=5.21
cc_332 ( N_C_c_557_n N_noxref_8_c_586_n ) capacitor c=0.0140071f //x=2.96 \
 //y=4.705 //x2=3.065 //y2=5.21
cc_333 ( N_C_M8_noxref_g N_noxref_8_c_590_n ) capacitor c=0.016576f //x=3.37 \
 //y=6.025 //x2=3.945 //y2=6.91
cc_334 ( N_C_M9_noxref_g N_noxref_8_c_590_n ) capacitor c=0.0166873f //x=3.81 \
 //y=6.025 //x2=3.945 //y2=6.91
cc_335 ( N_C_M9_noxref_g N_noxref_8_M9_noxref_d ) capacitor c=0.0351101f \
 //x=3.81 //y=6.025 //x2=3.885 //y2=5.025
