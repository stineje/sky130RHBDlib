// File: nmos_side_left.spi.NMOS_SIDE_LEFT.pxi
// Created: Tue Oct 15 15:58:18 2024
// 
simulator lang=spectre
cc_1 ( noxref_1 noxref_2 ) capacitor c=0.0395419f //x=0.435 //y=0.535 //x2=0 \
 //y2=0
cc_2 ( noxref_1 noxref_3 ) capacitor c=0.0216501f //x=0.435 //y=0.535 \
 //x2=0.622 //y2=0.925
cc_3 ( noxref_2 noxref_3 ) capacitor c=0.0927044f //x=0 //y=0 //x2=0.622 \
 //y2=0.925
