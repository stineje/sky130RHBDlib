magic
tech sky130A
magscale 1 2
timestamp 1652367678
<< metal1 >>
rect 1869 501 2114 535
use aoai4x1_pcell  aoai4x1_pcell_0
timestamp 1652367627
transform 1 0 0 0 1 0
box -87 -34 2085 1550
use invx1_pcell  invx1_pcell_0
timestamp 1652329846
transform 1 0 1998 0 1 0
box -87 -34 531 1550
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform -1 0 1850 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform 1 0 2146 0 1 518
box -53 -33 29 33
<< end >>
