magic
tech sky130A
magscale 1 2
timestamp 1669564332
<< nwell >>
rect -87 786 2307 1550
<< pwell >>
rect -34 -34 2254 544
<< nmos >>
rect 155 297 185 350
tri 185 297 201 313 sw
rect 155 267 261 297
tri 261 267 291 297 sw
rect 155 166 185 267
tri 185 251 201 267 nw
tri 245 251 261 267 ne
tri 185 166 201 182 sw
tri 245 166 261 182 se
rect 261 166 291 267
tri 155 136 185 166 ne
rect 185 136 261 166
tri 261 136 291 166 nw
rect 612 288 642 349
tri 642 288 658 304 sw
rect 806 296 836 349
tri 836 296 852 312 sw
rect 612 258 718 288
tri 718 258 748 288 sw
rect 806 266 912 296
tri 912 266 942 296 sw
rect 612 157 642 258
tri 642 242 658 258 nw
tri 702 242 718 258 ne
tri 642 157 658 173 sw
tri 702 157 718 173 se
rect 718 157 748 258
rect 806 165 836 266
tri 836 250 852 266 nw
tri 896 250 912 266 ne
tri 836 165 852 181 sw
tri 896 165 912 181 se
rect 912 165 942 266
tri 612 127 642 157 ne
rect 642 127 718 157
tri 718 127 748 157 nw
tri 806 135 836 165 ne
rect 836 135 912 165
tri 912 135 942 165 nw
rect 1278 288 1308 349
tri 1308 288 1324 304 sw
rect 1472 296 1502 349
tri 1502 296 1518 312 sw
rect 1278 258 1384 288
tri 1384 258 1414 288 sw
rect 1472 266 1578 296
tri 1578 266 1608 296 sw
rect 1278 157 1308 258
tri 1308 242 1324 258 nw
tri 1368 242 1384 258 ne
tri 1308 157 1324 173 sw
tri 1368 157 1384 173 se
rect 1384 157 1414 258
rect 1472 165 1502 266
tri 1502 250 1518 266 nw
tri 1562 250 1578 266 ne
tri 1502 165 1518 181 sw
tri 1562 165 1578 181 se
rect 1578 165 1608 266
tri 1278 127 1308 157 ne
rect 1308 127 1384 157
tri 1384 127 1414 157 nw
tri 1472 135 1502 165 ne
rect 1502 135 1578 165
tri 1578 135 1608 165 nw
tri 2019 297 2035 313 se
rect 2035 297 2065 350
tri 1929 267 1959 297 se
rect 1959 267 2065 297
rect 1929 166 1959 267
tri 1959 251 1975 267 nw
tri 2019 251 2035 267 ne
tri 1959 166 1975 182 sw
tri 2019 166 2035 182 se
rect 2035 166 2065 267
tri 1929 136 1959 166 ne
rect 1959 136 2035 166
tri 2035 136 2065 166 nw
<< pmos >>
rect 164 1004 194 1404
rect 252 1004 282 1404
rect 631 1004 661 1404
rect 719 1004 749 1404
rect 807 1004 837 1404
rect 895 1004 925 1404
rect 1297 1004 1327 1404
rect 1385 1004 1415 1404
rect 1473 1004 1503 1404
rect 1561 1004 1591 1404
rect 1938 1004 1968 1404
rect 2026 1004 2056 1404
<< ndiff >>
rect 99 334 155 350
rect 99 300 109 334
rect 143 300 155 334
rect 99 262 155 300
rect 185 334 345 350
rect 185 313 303 334
tri 185 297 201 313 ne
rect 201 300 303 313
rect 337 300 345 334
rect 201 297 345 300
tri 261 267 291 297 ne
rect 99 228 109 262
rect 143 228 155 262
rect 99 194 155 228
rect 99 160 109 194
rect 143 160 155 194
tri 185 251 201 267 se
rect 201 251 245 267
tri 245 251 261 267 sw
rect 185 218 261 251
rect 185 184 205 218
rect 239 184 261 218
rect 185 182 261 184
tri 185 166 201 182 ne
rect 201 166 245 182
tri 245 166 261 182 nw
rect 291 262 345 297
rect 291 228 303 262
rect 337 228 345 262
rect 291 194 345 228
rect 99 136 155 160
tri 155 136 185 166 sw
tri 261 136 291 166 se
rect 291 160 303 194
rect 337 160 345 194
rect 291 136 345 160
rect 99 124 345 136
rect 99 90 109 124
rect 143 90 205 124
rect 239 90 303 124
rect 337 90 345 124
rect 99 74 345 90
rect 556 333 612 349
rect 556 299 566 333
rect 600 299 612 333
rect 556 261 612 299
rect 642 333 806 349
rect 642 304 663 333
tri 642 288 658 304 ne
rect 658 299 663 304
rect 697 299 760 333
rect 794 299 806 333
rect 658 288 806 299
rect 836 312 998 349
tri 836 296 852 312 ne
rect 852 296 998 312
rect 556 227 566 261
rect 600 227 612 261
tri 718 258 748 288 ne
rect 748 261 806 288
tri 912 266 942 296 ne
rect 556 193 612 227
rect 556 159 566 193
rect 600 159 612 193
rect 556 127 612 159
tri 642 242 658 258 se
rect 658 242 702 258
tri 702 242 718 258 sw
rect 642 208 718 242
rect 642 174 663 208
rect 697 174 718 208
rect 642 173 718 174
tri 642 157 658 173 ne
rect 658 157 702 173
tri 702 157 718 173 nw
rect 748 227 760 261
rect 794 227 806 261
rect 748 193 806 227
rect 748 159 760 193
rect 794 159 806 193
tri 836 250 852 266 se
rect 852 250 896 266
tri 896 250 912 266 sw
rect 836 217 912 250
rect 836 183 857 217
rect 891 183 912 217
rect 836 181 912 183
tri 836 165 852 181 ne
rect 852 165 896 181
tri 896 165 912 181 nw
rect 942 261 998 296
rect 942 227 954 261
rect 988 227 998 261
rect 942 193 998 227
tri 612 127 642 157 sw
tri 718 127 748 157 se
rect 748 135 806 159
tri 806 135 836 165 sw
tri 912 135 942 165 se
rect 942 159 954 193
rect 988 159 998 193
rect 942 135 998 159
rect 748 127 998 135
rect 556 123 998 127
rect 556 89 566 123
rect 600 89 760 123
rect 794 89 857 123
rect 891 89 954 123
rect 988 89 998 123
rect 556 73 998 89
rect 1222 333 1278 349
rect 1222 299 1232 333
rect 1266 299 1278 333
rect 1222 261 1278 299
rect 1308 333 1472 349
rect 1308 304 1329 333
tri 1308 288 1324 304 ne
rect 1324 299 1329 304
rect 1363 299 1426 333
rect 1460 299 1472 333
rect 1324 288 1472 299
rect 1502 312 1664 349
tri 1502 296 1518 312 ne
rect 1518 296 1664 312
rect 1222 227 1232 261
rect 1266 227 1278 261
tri 1384 258 1414 288 ne
rect 1414 261 1472 288
tri 1578 266 1608 296 ne
rect 1222 193 1278 227
rect 1222 159 1232 193
rect 1266 159 1278 193
rect 1222 127 1278 159
tri 1308 242 1324 258 se
rect 1324 242 1368 258
tri 1368 242 1384 258 sw
rect 1308 208 1384 242
rect 1308 174 1329 208
rect 1363 174 1384 208
rect 1308 173 1384 174
tri 1308 157 1324 173 ne
rect 1324 157 1368 173
tri 1368 157 1384 173 nw
rect 1414 227 1426 261
rect 1460 227 1472 261
rect 1414 193 1472 227
rect 1414 159 1426 193
rect 1460 159 1472 193
tri 1502 250 1518 266 se
rect 1518 250 1562 266
tri 1562 250 1578 266 sw
rect 1502 217 1578 250
rect 1502 183 1523 217
rect 1557 183 1578 217
rect 1502 181 1578 183
tri 1502 165 1518 181 ne
rect 1518 165 1562 181
tri 1562 165 1578 181 nw
rect 1608 261 1664 296
rect 1608 227 1620 261
rect 1654 227 1664 261
rect 1608 193 1664 227
tri 1278 127 1308 157 sw
tri 1384 127 1414 157 se
rect 1414 135 1472 159
tri 1472 135 1502 165 sw
tri 1578 135 1608 165 se
rect 1608 159 1620 193
rect 1654 159 1664 193
rect 1608 135 1664 159
rect 1414 127 1664 135
rect 1222 123 1664 127
rect 1222 89 1232 123
rect 1266 89 1426 123
rect 1460 89 1523 123
rect 1557 89 1620 123
rect 1654 89 1664 123
rect 1222 73 1664 89
rect 1875 334 2035 350
rect 1875 300 1883 334
rect 1917 313 2035 334
rect 1917 300 2019 313
rect 1875 297 2019 300
tri 2019 297 2035 313 nw
rect 2065 334 2121 350
rect 2065 300 2077 334
rect 2111 300 2121 334
rect 1875 262 1929 297
tri 1929 267 1959 297 nw
rect 1875 228 1883 262
rect 1917 228 1929 262
rect 1875 194 1929 228
rect 1875 160 1883 194
rect 1917 160 1929 194
tri 1959 251 1975 267 se
rect 1975 251 2019 267
tri 2019 251 2035 267 sw
rect 1959 218 2035 251
rect 1959 184 1981 218
rect 2015 184 2035 218
rect 1959 182 2035 184
tri 1959 166 1975 182 ne
rect 1975 166 2019 182
tri 2019 166 2035 182 nw
rect 2065 262 2121 300
rect 2065 228 2077 262
rect 2111 228 2121 262
rect 2065 194 2121 228
rect 1875 136 1929 160
tri 1929 136 1959 166 sw
tri 2035 136 2065 166 se
rect 2065 160 2077 194
rect 2111 160 2121 194
rect 2065 136 2121 160
rect 1875 124 2121 136
rect 1875 90 1883 124
rect 1917 90 1981 124
rect 2015 90 2077 124
rect 2111 90 2121 124
rect 1875 74 2121 90
<< pdiff >>
rect 108 1366 164 1404
rect 108 1332 118 1366
rect 152 1332 164 1366
rect 108 1298 164 1332
rect 108 1264 118 1298
rect 152 1264 164 1298
rect 108 1230 164 1264
rect 108 1196 118 1230
rect 152 1196 164 1230
rect 108 1162 164 1196
rect 108 1128 118 1162
rect 152 1128 164 1162
rect 108 1093 164 1128
rect 108 1059 118 1093
rect 152 1059 164 1093
rect 108 1004 164 1059
rect 194 1366 252 1404
rect 194 1332 206 1366
rect 240 1332 252 1366
rect 194 1298 252 1332
rect 194 1264 206 1298
rect 240 1264 252 1298
rect 194 1230 252 1264
rect 194 1196 206 1230
rect 240 1196 252 1230
rect 194 1162 252 1196
rect 194 1128 206 1162
rect 240 1128 252 1162
rect 194 1093 252 1128
rect 194 1059 206 1093
rect 240 1059 252 1093
rect 194 1004 252 1059
rect 282 1366 336 1404
rect 282 1332 294 1366
rect 328 1332 336 1366
rect 282 1298 336 1332
rect 282 1264 294 1298
rect 328 1264 336 1298
rect 282 1230 336 1264
rect 282 1196 294 1230
rect 328 1196 336 1230
rect 282 1162 336 1196
rect 282 1128 294 1162
rect 328 1128 336 1162
rect 282 1093 336 1128
rect 282 1059 294 1093
rect 328 1059 336 1093
rect 282 1004 336 1059
rect 575 1364 631 1404
rect 575 1330 585 1364
rect 619 1330 631 1364
rect 575 1296 631 1330
rect 575 1262 585 1296
rect 619 1262 631 1296
rect 575 1228 631 1262
rect 575 1194 585 1228
rect 619 1194 631 1228
rect 575 1160 631 1194
rect 575 1126 585 1160
rect 619 1126 631 1160
rect 575 1092 631 1126
rect 575 1058 585 1092
rect 619 1058 631 1092
rect 575 1004 631 1058
rect 661 1296 719 1404
rect 661 1262 673 1296
rect 707 1262 719 1296
rect 661 1228 719 1262
rect 661 1194 673 1228
rect 707 1194 719 1228
rect 661 1160 719 1194
rect 661 1126 673 1160
rect 707 1126 719 1160
rect 661 1004 719 1126
rect 749 1364 807 1404
rect 749 1330 761 1364
rect 795 1330 807 1364
rect 749 1296 807 1330
rect 749 1262 761 1296
rect 795 1262 807 1296
rect 749 1228 807 1262
rect 749 1194 761 1228
rect 795 1194 807 1228
rect 749 1160 807 1194
rect 749 1126 761 1160
rect 795 1126 807 1160
rect 749 1092 807 1126
rect 749 1058 761 1092
rect 795 1058 807 1092
rect 749 1004 807 1058
rect 837 1296 895 1404
rect 837 1262 849 1296
rect 883 1262 895 1296
rect 837 1228 895 1262
rect 837 1194 849 1228
rect 883 1194 895 1228
rect 837 1160 895 1194
rect 837 1126 849 1160
rect 883 1126 895 1160
rect 837 1092 895 1126
rect 837 1058 849 1092
rect 883 1058 895 1092
rect 837 1004 895 1058
rect 925 1364 979 1404
rect 925 1330 937 1364
rect 971 1330 979 1364
rect 925 1296 979 1330
rect 925 1262 937 1296
rect 971 1262 979 1296
rect 925 1228 979 1262
rect 925 1194 937 1228
rect 971 1194 979 1228
rect 925 1160 979 1194
rect 925 1126 937 1160
rect 971 1126 979 1160
rect 925 1004 979 1126
rect 1241 1364 1297 1404
rect 1241 1330 1251 1364
rect 1285 1330 1297 1364
rect 1241 1296 1297 1330
rect 1241 1262 1251 1296
rect 1285 1262 1297 1296
rect 1241 1228 1297 1262
rect 1241 1194 1251 1228
rect 1285 1194 1297 1228
rect 1241 1160 1297 1194
rect 1241 1126 1251 1160
rect 1285 1126 1297 1160
rect 1241 1092 1297 1126
rect 1241 1058 1251 1092
rect 1285 1058 1297 1092
rect 1241 1004 1297 1058
rect 1327 1296 1385 1404
rect 1327 1262 1339 1296
rect 1373 1262 1385 1296
rect 1327 1228 1385 1262
rect 1327 1194 1339 1228
rect 1373 1194 1385 1228
rect 1327 1160 1385 1194
rect 1327 1126 1339 1160
rect 1373 1126 1385 1160
rect 1327 1004 1385 1126
rect 1415 1364 1473 1404
rect 1415 1330 1427 1364
rect 1461 1330 1473 1364
rect 1415 1296 1473 1330
rect 1415 1262 1427 1296
rect 1461 1262 1473 1296
rect 1415 1228 1473 1262
rect 1415 1194 1427 1228
rect 1461 1194 1473 1228
rect 1415 1160 1473 1194
rect 1415 1126 1427 1160
rect 1461 1126 1473 1160
rect 1415 1092 1473 1126
rect 1415 1058 1427 1092
rect 1461 1058 1473 1092
rect 1415 1004 1473 1058
rect 1503 1296 1561 1404
rect 1503 1262 1515 1296
rect 1549 1262 1561 1296
rect 1503 1228 1561 1262
rect 1503 1194 1515 1228
rect 1549 1194 1561 1228
rect 1503 1160 1561 1194
rect 1503 1126 1515 1160
rect 1549 1126 1561 1160
rect 1503 1092 1561 1126
rect 1503 1058 1515 1092
rect 1549 1058 1561 1092
rect 1503 1004 1561 1058
rect 1591 1364 1645 1404
rect 1591 1330 1603 1364
rect 1637 1330 1645 1364
rect 1591 1296 1645 1330
rect 1591 1262 1603 1296
rect 1637 1262 1645 1296
rect 1591 1228 1645 1262
rect 1591 1194 1603 1228
rect 1637 1194 1645 1228
rect 1591 1160 1645 1194
rect 1591 1126 1603 1160
rect 1637 1126 1645 1160
rect 1591 1004 1645 1126
rect 1884 1366 1938 1404
rect 1884 1332 1892 1366
rect 1926 1332 1938 1366
rect 1884 1298 1938 1332
rect 1884 1264 1892 1298
rect 1926 1264 1938 1298
rect 1884 1230 1938 1264
rect 1884 1196 1892 1230
rect 1926 1196 1938 1230
rect 1884 1162 1938 1196
rect 1884 1128 1892 1162
rect 1926 1128 1938 1162
rect 1884 1093 1938 1128
rect 1884 1059 1892 1093
rect 1926 1059 1938 1093
rect 1884 1004 1938 1059
rect 1968 1366 2026 1404
rect 1968 1332 1980 1366
rect 2014 1332 2026 1366
rect 1968 1298 2026 1332
rect 1968 1264 1980 1298
rect 2014 1264 2026 1298
rect 1968 1230 2026 1264
rect 1968 1196 1980 1230
rect 2014 1196 2026 1230
rect 1968 1162 2026 1196
rect 1968 1128 1980 1162
rect 2014 1128 2026 1162
rect 1968 1093 2026 1128
rect 1968 1059 1980 1093
rect 2014 1059 2026 1093
rect 1968 1004 2026 1059
rect 2056 1366 2112 1404
rect 2056 1332 2068 1366
rect 2102 1332 2112 1366
rect 2056 1298 2112 1332
rect 2056 1264 2068 1298
rect 2102 1264 2112 1298
rect 2056 1230 2112 1264
rect 2056 1196 2068 1230
rect 2102 1196 2112 1230
rect 2056 1162 2112 1196
rect 2056 1128 2068 1162
rect 2102 1128 2112 1162
rect 2056 1093 2112 1128
rect 2056 1059 2068 1093
rect 2102 1059 2112 1093
rect 2056 1004 2112 1059
<< ndiffc >>
rect 109 300 143 334
rect 303 300 337 334
rect 109 228 143 262
rect 109 160 143 194
rect 205 184 239 218
rect 303 228 337 262
rect 303 160 337 194
rect 109 90 143 124
rect 205 90 239 124
rect 303 90 337 124
rect 566 299 600 333
rect 663 299 697 333
rect 760 299 794 333
rect 566 227 600 261
rect 566 159 600 193
rect 663 174 697 208
rect 760 227 794 261
rect 760 159 794 193
rect 857 183 891 217
rect 954 227 988 261
rect 954 159 988 193
rect 566 89 600 123
rect 760 89 794 123
rect 857 89 891 123
rect 954 89 988 123
rect 1232 299 1266 333
rect 1329 299 1363 333
rect 1426 299 1460 333
rect 1232 227 1266 261
rect 1232 159 1266 193
rect 1329 174 1363 208
rect 1426 227 1460 261
rect 1426 159 1460 193
rect 1523 183 1557 217
rect 1620 227 1654 261
rect 1620 159 1654 193
rect 1232 89 1266 123
rect 1426 89 1460 123
rect 1523 89 1557 123
rect 1620 89 1654 123
rect 1883 300 1917 334
rect 2077 300 2111 334
rect 1883 228 1917 262
rect 1883 160 1917 194
rect 1981 184 2015 218
rect 2077 228 2111 262
rect 2077 160 2111 194
rect 1883 90 1917 124
rect 1981 90 2015 124
rect 2077 90 2111 124
<< pdiffc >>
rect 118 1332 152 1366
rect 118 1264 152 1298
rect 118 1196 152 1230
rect 118 1128 152 1162
rect 118 1059 152 1093
rect 206 1332 240 1366
rect 206 1264 240 1298
rect 206 1196 240 1230
rect 206 1128 240 1162
rect 206 1059 240 1093
rect 294 1332 328 1366
rect 294 1264 328 1298
rect 294 1196 328 1230
rect 294 1128 328 1162
rect 294 1059 328 1093
rect 585 1330 619 1364
rect 585 1262 619 1296
rect 585 1194 619 1228
rect 585 1126 619 1160
rect 585 1058 619 1092
rect 673 1262 707 1296
rect 673 1194 707 1228
rect 673 1126 707 1160
rect 761 1330 795 1364
rect 761 1262 795 1296
rect 761 1194 795 1228
rect 761 1126 795 1160
rect 761 1058 795 1092
rect 849 1262 883 1296
rect 849 1194 883 1228
rect 849 1126 883 1160
rect 849 1058 883 1092
rect 937 1330 971 1364
rect 937 1262 971 1296
rect 937 1194 971 1228
rect 937 1126 971 1160
rect 1251 1330 1285 1364
rect 1251 1262 1285 1296
rect 1251 1194 1285 1228
rect 1251 1126 1285 1160
rect 1251 1058 1285 1092
rect 1339 1262 1373 1296
rect 1339 1194 1373 1228
rect 1339 1126 1373 1160
rect 1427 1330 1461 1364
rect 1427 1262 1461 1296
rect 1427 1194 1461 1228
rect 1427 1126 1461 1160
rect 1427 1058 1461 1092
rect 1515 1262 1549 1296
rect 1515 1194 1549 1228
rect 1515 1126 1549 1160
rect 1515 1058 1549 1092
rect 1603 1330 1637 1364
rect 1603 1262 1637 1296
rect 1603 1194 1637 1228
rect 1603 1126 1637 1160
rect 1892 1332 1926 1366
rect 1892 1264 1926 1298
rect 1892 1196 1926 1230
rect 1892 1128 1926 1162
rect 1892 1059 1926 1093
rect 1980 1332 2014 1366
rect 1980 1264 2014 1298
rect 1980 1196 2014 1230
rect 1980 1128 2014 1162
rect 1980 1059 2014 1093
rect 2068 1332 2102 1366
rect 2068 1264 2102 1298
rect 2068 1196 2102 1230
rect 2068 1128 2102 1162
rect 2068 1059 2102 1093
<< psubdiff >>
rect -34 482 2254 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 410 461 478 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 410 427 427 461
rect 461 427 478 461
rect 1076 461 1144 482
rect -34 313 34 353
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 410 313 478 353
rect 1076 427 1093 461
rect 1127 427 1144 461
rect 1742 461 1810 482
rect 1076 387 1144 427
rect 1076 353 1093 387
rect 1127 353 1144 387
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect -34 17 34 57
rect 410 57 427 91
rect 461 57 478 91
rect 1076 313 1144 353
rect 1742 427 1759 461
rect 1793 427 1810 461
rect 2186 461 2254 482
rect 1742 387 1810 427
rect 1742 353 1759 387
rect 1793 353 1810 387
rect 1076 279 1093 313
rect 1127 279 1144 313
rect 1076 239 1144 279
rect 1076 205 1093 239
rect 1127 205 1144 239
rect 1076 165 1144 205
rect 1076 131 1093 165
rect 1127 131 1144 165
rect 1076 91 1144 131
rect 410 17 478 57
rect 1076 57 1093 91
rect 1127 57 1144 91
rect 1742 313 1810 353
rect 2186 427 2203 461
rect 2237 427 2254 461
rect 2186 387 2254 427
rect 2186 353 2203 387
rect 2237 353 2254 387
rect 1742 279 1759 313
rect 1793 279 1810 313
rect 1742 239 1810 279
rect 1742 205 1759 239
rect 1793 205 1810 239
rect 1742 165 1810 205
rect 1742 131 1759 165
rect 1793 131 1810 165
rect 1742 91 1810 131
rect 1076 17 1144 57
rect 1742 57 1759 91
rect 1793 57 1810 91
rect 2186 313 2254 353
rect 2186 279 2203 313
rect 2237 279 2254 313
rect 2186 239 2254 279
rect 2186 205 2203 239
rect 2237 205 2254 239
rect 2186 165 2254 205
rect 2186 131 2203 165
rect 2237 131 2254 165
rect 2186 91 2254 131
rect 1742 17 1810 57
rect 2186 57 2203 91
rect 2237 57 2254 91
rect 2186 17 2254 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2254 17
rect -34 -34 2254 -17
<< nsubdiff >>
rect -34 1497 2254 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2254 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 410 1423 478 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 1076 1423 1144 1463
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 410 979 478 1019
rect 1076 1389 1093 1423
rect 1127 1389 1144 1423
rect 1742 1423 1810 1463
rect 1076 1349 1144 1389
rect 1076 1315 1093 1349
rect 1127 1315 1144 1349
rect 1076 1275 1144 1315
rect 1076 1241 1093 1275
rect 1127 1241 1144 1275
rect 1076 1201 1144 1241
rect 1076 1167 1093 1201
rect 1127 1167 1144 1201
rect 1076 1127 1144 1167
rect 1076 1093 1093 1127
rect 1127 1093 1144 1127
rect 1076 1053 1144 1093
rect 1076 1019 1093 1053
rect 1127 1019 1144 1053
rect 410 945 427 979
rect 461 945 478 979
rect -34 871 -17 905
rect 17 884 34 905
rect 410 905 478 945
rect 1076 979 1144 1019
rect 1742 1389 1759 1423
rect 1793 1389 1810 1423
rect 2186 1423 2254 1463
rect 1742 1349 1810 1389
rect 1742 1315 1759 1349
rect 1793 1315 1810 1349
rect 1742 1275 1810 1315
rect 1742 1241 1759 1275
rect 1793 1241 1810 1275
rect 1742 1201 1810 1241
rect 1742 1167 1759 1201
rect 1793 1167 1810 1201
rect 1742 1127 1810 1167
rect 1742 1093 1759 1127
rect 1793 1093 1810 1127
rect 1742 1053 1810 1093
rect 1742 1019 1759 1053
rect 1793 1019 1810 1053
rect 1076 945 1093 979
rect 1127 945 1144 979
rect 410 884 427 905
rect 17 871 427 884
rect 461 884 478 905
rect 1076 905 1144 945
rect 1742 979 1810 1019
rect 2186 1389 2203 1423
rect 2237 1389 2254 1423
rect 2186 1349 2254 1389
rect 2186 1315 2203 1349
rect 2237 1315 2254 1349
rect 2186 1275 2254 1315
rect 2186 1241 2203 1275
rect 2237 1241 2254 1275
rect 2186 1201 2254 1241
rect 2186 1167 2203 1201
rect 2237 1167 2254 1201
rect 2186 1127 2254 1167
rect 2186 1093 2203 1127
rect 2237 1093 2254 1127
rect 2186 1053 2254 1093
rect 2186 1019 2203 1053
rect 2237 1019 2254 1053
rect 1742 945 1759 979
rect 1793 945 1810 979
rect 1076 884 1093 905
rect 461 871 1093 884
rect 1127 884 1144 905
rect 1742 905 1810 945
rect 2186 979 2254 1019
rect 2186 945 2203 979
rect 2237 945 2254 979
rect 1742 884 1759 905
rect 1127 871 1759 884
rect 1793 884 1810 905
rect 2186 905 2254 945
rect 2186 884 2203 905
rect 1793 871 2203 884
rect 2237 871 2254 905
rect -34 822 2254 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 427 427 461 461
rect 427 353 461 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1093 427 1127 461
rect 1093 353 1127 387
rect 427 279 461 313
rect 427 205 461 239
rect 427 131 461 165
rect 427 57 461 91
rect 1759 427 1793 461
rect 1759 353 1793 387
rect 1093 279 1127 313
rect 1093 205 1127 239
rect 1093 131 1127 165
rect 1093 57 1127 91
rect 2203 427 2237 461
rect 2203 353 2237 387
rect 1759 279 1793 313
rect 1759 205 1793 239
rect 1759 131 1793 165
rect 1759 57 1793 91
rect 2203 279 2237 313
rect 2203 205 2237 239
rect 2203 131 2237 165
rect 2203 57 2237 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 427 1389 461 1423
rect 427 1315 461 1349
rect 427 1241 461 1275
rect 427 1167 461 1201
rect 427 1093 461 1127
rect 427 1019 461 1053
rect -17 945 17 979
rect 1093 1389 1127 1423
rect 1093 1315 1127 1349
rect 1093 1241 1127 1275
rect 1093 1167 1127 1201
rect 1093 1093 1127 1127
rect 1093 1019 1127 1053
rect 427 945 461 979
rect -17 871 17 905
rect 1759 1389 1793 1423
rect 1759 1315 1793 1349
rect 1759 1241 1793 1275
rect 1759 1167 1793 1201
rect 1759 1093 1793 1127
rect 1759 1019 1793 1053
rect 1093 945 1127 979
rect 427 871 461 905
rect 2203 1389 2237 1423
rect 2203 1315 2237 1349
rect 2203 1241 2237 1275
rect 2203 1167 2237 1201
rect 2203 1093 2237 1127
rect 2203 1019 2237 1053
rect 1759 945 1793 979
rect 1093 871 1127 905
rect 2203 945 2237 979
rect 1759 871 1793 905
rect 2203 871 2237 905
<< poly >>
rect 164 1404 194 1430
rect 252 1404 282 1430
rect 631 1404 661 1430
rect 719 1404 749 1430
rect 807 1404 837 1430
rect 895 1404 925 1430
rect 164 973 194 1004
rect 252 973 282 1004
rect 121 957 282 973
rect 121 923 131 957
rect 165 943 282 957
rect 1297 1404 1327 1430
rect 1385 1404 1415 1430
rect 1473 1404 1503 1430
rect 1561 1404 1591 1430
rect 165 923 175 943
rect 121 907 175 923
rect 631 973 661 1004
rect 719 973 749 1004
rect 631 957 749 973
rect 631 943 649 957
rect 639 923 649 943
rect 683 943 749 957
rect 807 973 837 1004
rect 895 973 925 1004
rect 807 957 925 973
rect 807 943 871 957
rect 683 923 693 943
rect 639 907 693 923
rect 861 923 871 943
rect 905 943 925 957
rect 1938 1404 1968 1430
rect 2026 1404 2056 1430
rect 905 923 915 943
rect 861 907 915 923
rect 1297 973 1327 1004
rect 1385 973 1415 1004
rect 1297 957 1415 973
rect 1297 943 1315 957
rect 1305 923 1315 943
rect 1349 943 1415 957
rect 1473 973 1503 1004
rect 1561 973 1591 1004
rect 1473 957 1591 973
rect 1473 943 1537 957
rect 1349 923 1359 943
rect 1305 907 1359 923
rect 1527 923 1537 943
rect 1571 943 1591 957
rect 1571 923 1581 943
rect 1527 907 1581 923
rect 1938 973 1968 1004
rect 2026 973 2056 1004
rect 1938 957 2099 973
rect 1938 943 2055 957
rect 2045 923 2055 943
rect 2089 923 2099 957
rect 2045 907 2099 923
rect 121 434 175 450
rect 121 400 131 434
rect 165 413 175 434
rect 165 400 185 413
rect 121 384 185 400
rect 155 350 185 384
rect 639 433 693 449
rect 639 413 649 433
rect 612 399 649 413
rect 683 399 693 433
rect 861 433 915 449
rect 861 413 871 433
rect 612 383 693 399
rect 806 399 871 413
rect 905 399 915 433
rect 806 383 915 399
rect 1305 433 1359 449
rect 1305 413 1315 433
rect 612 349 642 383
rect 806 349 836 383
rect 1278 399 1315 413
rect 1349 399 1359 433
rect 1527 433 1581 449
rect 1527 413 1537 433
rect 1278 383 1359 399
rect 1472 399 1537 413
rect 1571 399 1581 433
rect 1472 383 1581 399
rect 2045 434 2099 450
rect 2045 413 2055 434
rect 1278 349 1308 383
rect 1472 349 1502 383
rect 2035 400 2055 413
rect 2089 400 2099 434
rect 2035 384 2099 400
rect 2035 350 2065 384
<< polycont >>
rect 131 923 165 957
rect 649 923 683 957
rect 871 923 905 957
rect 1315 923 1349 957
rect 1537 923 1571 957
rect 2055 923 2089 957
rect 131 400 165 434
rect 649 399 683 433
rect 871 399 905 433
rect 1315 399 1349 433
rect 1537 399 1571 433
rect 2055 400 2089 434
<< locali >>
rect -34 1497 2254 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2254 1497
rect -34 1446 2254 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 118 1366 152 1446
rect 118 1298 152 1332
rect 118 1230 152 1264
rect 118 1162 152 1196
rect 118 1093 152 1128
rect 118 1037 152 1059
rect 206 1366 240 1404
rect 206 1298 240 1332
rect 206 1230 240 1264
rect 206 1162 240 1196
rect 206 1093 240 1128
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 131 957 165 973
rect 131 831 165 923
rect 206 933 240 1059
rect 294 1366 328 1446
rect 294 1298 328 1332
rect 294 1230 328 1264
rect 294 1162 328 1196
rect 294 1093 328 1128
rect 294 1037 328 1059
rect 410 1423 478 1446
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect 585 1364 619 1380
rect 585 1296 619 1330
rect 585 1228 619 1262
rect 585 1160 619 1194
rect 585 1092 619 1126
rect 673 1296 707 1446
rect 1076 1423 1144 1446
rect 673 1228 707 1262
rect 673 1160 707 1194
rect 673 1110 707 1126
rect 761 1364 971 1398
rect 761 1296 795 1330
rect 761 1228 795 1262
rect 761 1160 795 1194
rect 761 1092 795 1126
rect 585 1024 795 1058
rect 849 1296 883 1312
rect 849 1228 883 1262
rect 849 1160 883 1194
rect 849 1092 883 1126
rect 937 1296 971 1330
rect 937 1228 971 1262
rect 937 1160 971 1194
rect 937 1110 971 1126
rect 1076 1389 1093 1423
rect 1127 1389 1144 1423
rect 1076 1349 1144 1389
rect 1076 1315 1093 1349
rect 1127 1315 1144 1349
rect 1076 1275 1144 1315
rect 1076 1241 1093 1275
rect 1127 1241 1144 1275
rect 1076 1201 1144 1241
rect 1076 1167 1093 1201
rect 1127 1167 1144 1201
rect 1076 1127 1144 1167
rect 1076 1093 1093 1127
rect 1127 1093 1144 1127
rect 849 1024 979 1058
rect 410 979 478 1019
rect 410 945 427 979
rect 461 945 478 979
rect 206 899 313 933
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 131 434 165 797
rect 279 535 313 899
rect 410 905 478 945
rect 410 871 427 905
rect 461 871 478 905
rect 410 822 478 871
rect 649 957 683 973
rect 649 831 683 923
rect 279 433 313 501
rect 131 384 165 400
rect 205 399 313 433
rect 410 461 478 544
rect 410 427 427 461
rect 461 427 478 461
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect -34 34 34 57
rect 109 334 143 350
rect 109 262 143 300
rect 109 194 143 228
rect 205 218 239 399
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect 649 433 683 797
rect 871 957 905 973
rect 871 831 905 923
rect 871 781 905 797
rect 945 757 979 1024
rect 1076 1053 1144 1093
rect 1076 1019 1093 1053
rect 1127 1019 1144 1053
rect 1251 1364 1285 1380
rect 1251 1296 1285 1330
rect 1251 1228 1285 1262
rect 1251 1160 1285 1194
rect 1251 1092 1285 1126
rect 1339 1296 1373 1446
rect 1742 1423 1810 1446
rect 1339 1228 1373 1262
rect 1339 1160 1373 1194
rect 1339 1110 1373 1126
rect 1427 1364 1637 1398
rect 1427 1296 1461 1330
rect 1427 1228 1461 1262
rect 1427 1160 1461 1194
rect 1427 1092 1461 1126
rect 1251 1024 1461 1058
rect 1515 1296 1549 1312
rect 1515 1228 1549 1262
rect 1515 1160 1549 1194
rect 1515 1092 1549 1126
rect 1603 1296 1637 1330
rect 1603 1228 1637 1262
rect 1603 1160 1637 1194
rect 1603 1110 1637 1126
rect 1742 1389 1759 1423
rect 1793 1389 1810 1423
rect 1742 1349 1810 1389
rect 1742 1315 1759 1349
rect 1793 1315 1810 1349
rect 1742 1275 1810 1315
rect 1742 1241 1759 1275
rect 1793 1241 1810 1275
rect 1742 1201 1810 1241
rect 1742 1167 1759 1201
rect 1793 1167 1810 1201
rect 1742 1127 1810 1167
rect 1742 1093 1759 1127
rect 1793 1093 1810 1127
rect 1515 1024 1645 1058
rect 1076 979 1144 1019
rect 1076 945 1093 979
rect 1127 945 1144 979
rect 1076 905 1144 945
rect 1076 871 1093 905
rect 1127 871 1144 905
rect 1076 822 1144 871
rect 1315 957 1349 973
rect 1315 905 1349 923
rect 1315 855 1349 871
rect 1537 957 1571 973
rect 649 383 683 399
rect 871 609 905 625
rect 871 433 905 575
rect 871 383 905 399
rect 205 168 239 184
rect 303 334 337 350
rect 303 262 337 300
rect 303 194 337 228
rect 109 124 143 160
rect 303 124 337 160
rect 143 90 205 124
rect 239 90 303 124
rect 109 34 143 90
rect 206 34 240 90
rect 303 34 337 90
rect 410 313 478 353
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect 410 57 427 91
rect 461 57 478 91
rect 566 333 600 349
rect 760 333 794 349
rect 945 347 979 723
rect 1315 683 1349 699
rect 600 299 663 333
rect 697 299 760 333
rect 566 261 600 299
rect 566 193 600 227
rect 760 261 794 299
rect 566 123 600 159
rect 566 73 600 89
rect 663 208 697 224
rect 410 34 478 57
rect 663 34 697 174
rect 760 193 794 227
rect 857 313 979 347
rect 1076 461 1144 544
rect 1076 427 1093 461
rect 1127 427 1144 461
rect 1076 387 1144 427
rect 1076 353 1093 387
rect 1127 353 1144 387
rect 1315 433 1349 649
rect 1315 383 1349 399
rect 1537 535 1571 923
rect 1537 433 1571 501
rect 1537 383 1571 399
rect 1611 757 1645 1024
rect 1742 1053 1810 1093
rect 1742 1019 1759 1053
rect 1793 1019 1810 1053
rect 1892 1366 1926 1446
rect 1892 1298 1926 1332
rect 1892 1230 1926 1264
rect 1892 1162 1926 1196
rect 1892 1093 1926 1128
rect 1892 1037 1926 1059
rect 1980 1366 2014 1404
rect 1980 1298 2014 1332
rect 1980 1230 2014 1264
rect 1980 1162 2014 1196
rect 1980 1093 2014 1128
rect 1742 979 1810 1019
rect 1742 945 1759 979
rect 1793 945 1810 979
rect 1742 905 1810 945
rect 1980 933 2014 1059
rect 2068 1366 2102 1446
rect 2068 1298 2102 1332
rect 2068 1230 2102 1264
rect 2068 1162 2102 1196
rect 2068 1093 2102 1128
rect 2068 1037 2102 1059
rect 2186 1423 2254 1446
rect 2186 1389 2203 1423
rect 2237 1389 2254 1423
rect 2186 1349 2254 1389
rect 2186 1315 2203 1349
rect 2237 1315 2254 1349
rect 2186 1275 2254 1315
rect 2186 1241 2203 1275
rect 2237 1241 2254 1275
rect 2186 1201 2254 1241
rect 2186 1167 2203 1201
rect 2237 1167 2254 1201
rect 2186 1127 2254 1167
rect 2186 1093 2203 1127
rect 2237 1093 2254 1127
rect 2186 1053 2254 1093
rect 2186 1019 2203 1053
rect 2237 1019 2254 1053
rect 2186 979 2254 1019
rect 1742 871 1759 905
rect 1793 871 1810 905
rect 1742 822 1810 871
rect 1907 905 2014 933
rect 1941 899 2014 905
rect 2055 957 2089 973
rect 1076 313 1144 353
rect 857 217 891 313
rect 1076 279 1093 313
rect 1127 279 1144 313
rect 857 167 891 183
rect 954 261 988 277
rect 954 193 988 227
rect 760 123 794 159
rect 954 123 988 159
rect 794 89 857 123
rect 891 89 954 123
rect 760 73 794 89
rect 954 73 988 89
rect 1076 239 1144 279
rect 1076 205 1093 239
rect 1127 205 1144 239
rect 1076 165 1144 205
rect 1076 131 1093 165
rect 1127 131 1144 165
rect 1076 91 1144 131
rect 1076 57 1093 91
rect 1127 57 1144 91
rect 1232 333 1266 349
rect 1426 333 1460 349
rect 1611 347 1645 723
rect 1907 609 1941 871
rect 1266 299 1329 333
rect 1363 299 1426 333
rect 1232 261 1266 299
rect 1232 193 1266 227
rect 1426 261 1460 299
rect 1232 123 1266 159
rect 1232 73 1266 89
rect 1329 208 1363 224
rect 1076 34 1144 57
rect 1329 34 1363 174
rect 1426 193 1460 227
rect 1523 313 1645 347
rect 1742 461 1810 544
rect 1742 427 1759 461
rect 1793 427 1810 461
rect 1742 387 1810 427
rect 1907 433 1941 575
rect 2055 831 2089 923
rect 2186 945 2203 979
rect 2237 945 2254 979
rect 2186 905 2254 945
rect 2186 871 2203 905
rect 2237 871 2254 905
rect 2186 822 2254 871
rect 2055 683 2089 797
rect 2055 434 2089 649
rect 1907 399 2015 433
rect 1742 353 1759 387
rect 1793 353 1810 387
rect 1742 313 1810 353
rect 1523 217 1557 313
rect 1742 279 1759 313
rect 1793 279 1810 313
rect 1523 167 1557 183
rect 1620 261 1654 277
rect 1620 193 1654 227
rect 1426 123 1460 159
rect 1620 123 1654 159
rect 1460 89 1523 123
rect 1557 89 1620 123
rect 1426 73 1460 89
rect 1620 73 1654 89
rect 1742 239 1810 279
rect 1742 205 1759 239
rect 1793 205 1810 239
rect 1742 165 1810 205
rect 1742 131 1759 165
rect 1793 131 1810 165
rect 1742 91 1810 131
rect 1742 57 1759 91
rect 1793 57 1810 91
rect 1742 34 1810 57
rect 1883 334 1917 350
rect 1883 262 1917 300
rect 1883 194 1917 228
rect 1981 218 2015 399
rect 2055 384 2089 400
rect 2186 461 2254 544
rect 2186 427 2203 461
rect 2237 427 2254 461
rect 2186 387 2254 427
rect 2186 353 2203 387
rect 2237 353 2254 387
rect 1981 168 2015 184
rect 2077 334 2111 350
rect 2077 262 2111 300
rect 2077 194 2111 228
rect 1883 124 1917 160
rect 2077 124 2111 160
rect 1917 90 1981 124
rect 2015 90 2077 124
rect 1883 34 1917 90
rect 1980 34 2014 90
rect 2077 34 2111 90
rect 2186 313 2254 353
rect 2186 279 2203 313
rect 2237 279 2254 313
rect 2186 239 2254 279
rect 2186 205 2203 239
rect 2237 205 2254 239
rect 2186 165 2254 205
rect 2186 131 2203 165
rect 2237 131 2254 165
rect 2186 91 2254 131
rect 2186 57 2203 91
rect 2237 57 2254 91
rect 2186 34 2254 57
rect -34 17 2254 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2254 17
rect -34 -34 2254 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 131 797 165 831
rect 649 797 683 831
rect 279 501 313 535
rect 871 797 905 831
rect 1315 871 1349 905
rect 945 723 979 757
rect 871 575 905 609
rect 1315 649 1349 683
rect 1537 501 1571 535
rect 1907 871 1941 905
rect 1611 723 1645 757
rect 1907 575 1941 609
rect 2055 797 2089 831
rect 2055 649 2089 683
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
<< metal1 >>
rect -34 1497 2254 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2254 1497
rect -34 1446 2254 1463
rect 1309 905 1355 911
rect 1901 905 1947 911
rect 1303 871 1315 905
rect 1349 871 1907 905
rect 1941 871 1953 905
rect 1309 865 1355 871
rect 1901 865 1947 871
rect 125 831 171 837
rect 643 831 689 837
rect 865 831 911 837
rect 2049 831 2095 837
rect 119 797 131 831
rect 165 797 649 831
rect 683 797 695 831
rect 859 797 871 831
rect 905 797 2055 831
rect 2089 797 2101 831
rect 125 791 171 797
rect 643 791 689 797
rect 865 791 911 797
rect 2049 791 2095 797
rect 939 757 985 763
rect 1605 757 1651 763
rect 933 723 945 757
rect 979 723 1611 757
rect 1645 723 1657 757
rect 939 717 985 723
rect 1605 717 1651 723
rect 1309 683 1355 689
rect 2049 683 2095 689
rect 1303 649 1315 683
rect 1349 649 2055 683
rect 2089 649 2101 683
rect 1309 643 1355 649
rect 2049 643 2095 649
rect 865 609 911 615
rect 1901 609 1947 615
rect 859 575 871 609
rect 905 575 1907 609
rect 1941 575 1953 609
rect 865 569 911 575
rect 1901 569 1947 575
rect 273 535 319 541
rect 1531 535 1577 541
rect 267 501 279 535
rect 313 501 1537 535
rect 1571 501 1583 535
rect 273 495 319 501
rect 1531 495 1577 501
rect -34 17 2254 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2254 17
rect -34 -34 2254 -17
<< labels >>
rlabel metal1 1611 723 1645 757 1 Y
port 1 n
rlabel metal1 1611 501 1645 535 1 Y
port 2 n
rlabel metal1 1611 427 1645 461 1 Y
port 3 n
rlabel metal1 1611 945 1645 979 1 Y
port 4 n
rlabel metal1 945 723 979 757 1 Y
port 5 n
rlabel metal1 945 649 979 683 1 Y
port 6 n
rlabel metal1 945 427 979 461 1 Y
port 7 n
rlabel metal1 945 871 979 905 1 Y
port 8 n
rlabel metal1 131 871 165 905 1 A
port 9 n
rlabel metal1 131 797 165 831 1 A
port 10 n
rlabel metal1 131 723 165 757 1 A
port 11 n
rlabel metal1 131 649 165 683 1 A
port 12 n
rlabel metal1 131 575 165 609 1 A
port 13 n
rlabel metal1 131 501 165 535 1 A
port 14 n
rlabel metal1 649 501 683 535 1 A
port 15 n
rlabel metal1 649 575 683 609 1 A
port 16 n
rlabel metal1 649 649 683 683 1 A
port 17 n
rlabel metal1 649 723 683 757 1 A
port 18 n
rlabel metal1 649 797 683 831 1 A
port 19 n
rlabel metal1 649 871 683 905 1 A
port 20 n
rlabel metal1 2055 649 2089 683 1 B
port 21 n
rlabel metal1 2055 575 2089 609 1 B
port 22 n
rlabel metal1 2055 723 2089 757 1 B
port 23 n
rlabel metal1 2055 501 2089 535 1 B
port 24 n
rlabel metal1 2055 797 2089 831 1 B
port 25 n
rlabel metal1 2055 871 2089 905 1 B
port 26 n
rlabel metal1 871 797 905 831 1 B
port 27 n
rlabel metal1 1315 649 1349 683 1 B
port 28 n
rlabel metal1 1315 427 1349 461 1 B
port 29 n
rlabel metal1 871 871 905 905 1 B
port 30 n
rlabel metal1 -34 1446 2254 1514 1 VPWR
port 31 n
rlabel metal1 -34 -34 2254 34 1 VGND
port 32 n
rlabel nwell 57 1463 91 1497 1 VPB
port 33 n
rlabel pwell 57 -17 91 17 1 VNB
port 34 n
<< end >>
