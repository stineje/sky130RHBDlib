magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -66 377 3906 897
<< pwell >>
rect 1843 236 3125 291
rect 111 221 3125 236
rect 3399 221 3836 283
rect 111 43 3836 221
rect -26 -43 3866 43
<< locali >>
rect 21 236 223 302
rect 399 401 476 515
rect 582 532 641 652
rect 399 367 635 401
rect 976 367 1127 505
rect 399 289 449 367
rect 601 310 1127 367
rect 3097 391 3228 499
rect 3764 103 3815 751
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3840 831
rect 61 655 127 741
rect 284 735 474 741
rect 284 701 290 735
rect 324 701 362 735
rect 396 701 434 735
rect 468 701 474 735
rect 284 691 474 701
rect 512 707 711 741
rect 512 655 546 707
rect 61 621 546 655
rect 61 372 95 621
rect 146 551 546 585
rect 146 451 212 551
rect 61 338 293 372
rect 133 87 199 199
rect 259 183 293 338
rect 329 253 363 551
rect 512 496 546 551
rect 677 645 711 707
rect 747 735 925 741
rect 781 701 819 735
rect 853 701 891 735
rect 747 681 925 701
rect 961 727 1201 761
rect 961 645 995 727
rect 677 611 995 645
rect 1031 575 1097 691
rect 1151 633 1201 727
rect 677 541 1097 575
rect 677 496 711 541
rect 512 462 711 496
rect 793 498 935 505
rect 793 464 895 498
rect 929 464 935 498
rect 793 458 935 464
rect 793 403 860 458
rect 496 269 562 331
rect 496 253 1107 269
rect 329 235 1107 253
rect 329 219 562 235
rect 259 123 497 183
rect 729 87 795 199
rect 133 53 795 87
rect 831 113 1021 199
rect 831 79 837 113
rect 871 79 909 113
rect 943 79 981 113
rect 1015 79 1021 113
rect 1057 103 1107 235
rect 1167 201 1201 633
rect 1151 103 1201 201
rect 1237 727 1443 761
rect 831 73 1021 79
rect 1237 87 1271 727
rect 1307 577 1373 691
rect 1409 647 1443 727
rect 1481 735 1671 741
rect 1481 701 1487 735
rect 1521 701 1559 735
rect 1593 701 1631 735
rect 1665 701 1671 735
rect 1481 683 1671 701
rect 1707 727 1957 761
rect 1707 647 1741 727
rect 1409 613 1741 647
rect 1777 577 1843 691
rect 1307 543 1843 577
rect 1307 199 1341 543
rect 1390 417 1456 507
rect 1390 383 1521 417
rect 1409 269 1451 347
rect 1487 339 1521 383
rect 1557 409 1623 507
rect 1659 498 1752 507
rect 1659 464 1663 498
rect 1697 464 1752 498
rect 1659 445 1752 464
rect 1809 479 1843 543
rect 1891 661 1957 727
rect 1993 737 2183 747
rect 1993 703 1999 737
rect 2033 703 2071 737
rect 2105 703 2143 737
rect 2177 703 2183 737
rect 1993 697 2183 703
rect 2603 735 2793 741
rect 2603 701 2609 735
rect 2643 701 2681 735
rect 2715 701 2753 735
rect 2787 701 2793 735
rect 3055 735 3233 741
rect 2603 674 2793 701
rect 2829 671 3019 705
rect 1891 627 2562 661
rect 2829 638 2863 671
rect 1891 539 1957 627
rect 2192 535 2288 591
rect 2098 479 2156 511
rect 1809 445 2156 479
rect 2192 409 2226 535
rect 2324 491 2358 627
rect 1557 375 2226 409
rect 1487 305 2156 339
rect 1409 235 1927 269
rect 1307 123 1373 199
rect 1409 87 1451 235
rect 1237 53 1451 87
rect 1623 113 1813 199
rect 1861 177 1927 235
rect 1623 79 1629 113
rect 1663 79 1701 113
rect 1735 79 1773 113
rect 1807 79 1813 113
rect 1623 73 1813 79
rect 1968 113 2086 269
rect 1968 79 1974 113
rect 2008 79 2046 113
rect 2080 79 2086 113
rect 1968 73 2086 79
rect 2122 87 2156 305
rect 2192 257 2226 375
rect 2262 457 2358 491
rect 2262 293 2296 457
rect 2394 421 2460 591
rect 2496 457 2562 627
rect 2606 604 2863 638
rect 2606 421 2640 604
rect 2899 568 2949 635
rect 2332 387 2640 421
rect 2676 534 2949 568
rect 2332 273 2366 387
rect 2676 379 2742 534
rect 2808 464 2815 498
rect 2849 464 2874 498
rect 2808 379 2874 464
rect 2402 343 2604 351
rect 2402 309 2879 343
rect 2192 123 2265 257
rect 2332 123 2421 273
rect 2457 87 2491 309
rect 2122 53 2491 87
rect 2617 113 2807 273
rect 2617 79 2623 113
rect 2657 79 2695 113
rect 2729 79 2767 113
rect 2801 79 2807 113
rect 2845 141 2879 309
rect 2915 269 2949 534
rect 2985 455 3019 671
rect 3089 701 3127 735
rect 3161 701 3199 735
rect 3546 735 3728 751
rect 3546 701 3548 735
rect 3582 701 3620 735
rect 3654 701 3692 735
rect 3726 701 3728 735
rect 3055 535 3233 701
rect 2985 355 3051 455
rect 3269 425 3319 701
rect 3413 461 3510 601
rect 3269 391 3440 425
rect 2985 321 3370 355
rect 3406 285 3440 391
rect 2915 235 3107 269
rect 3041 177 3107 235
rect 3151 251 3440 285
rect 3476 363 3510 461
rect 3546 435 3728 701
rect 3476 297 3723 363
rect 3151 141 3217 251
rect 3476 215 3510 297
rect 2845 107 3217 141
rect 3255 113 3373 199
rect 3421 165 3510 215
rect 2617 73 2807 79
rect 3255 79 3261 113
rect 3295 79 3333 113
rect 3367 79 3373 113
rect 3255 73 3373 79
rect 3546 113 3728 261
rect 3546 79 3548 113
rect 3582 79 3620 113
rect 3654 79 3692 113
rect 3726 79 3728 113
rect 3546 73 3728 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3840 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 290 701 324 735
rect 362 701 396 735
rect 434 701 468 735
rect 747 701 781 735
rect 819 701 853 735
rect 891 701 925 735
rect 895 464 929 498
rect 837 79 871 113
rect 909 79 943 113
rect 981 79 1015 113
rect 1487 701 1521 735
rect 1559 701 1593 735
rect 1631 701 1665 735
rect 1663 464 1697 498
rect 1999 703 2033 737
rect 2071 703 2105 737
rect 2143 703 2177 737
rect 2609 701 2643 735
rect 2681 701 2715 735
rect 2753 701 2787 735
rect 1629 79 1663 113
rect 1701 79 1735 113
rect 1773 79 1807 113
rect 1974 79 2008 113
rect 2046 79 2080 113
rect 2815 464 2849 498
rect 2623 79 2657 113
rect 2695 79 2729 113
rect 2767 79 2801 113
rect 3055 701 3089 735
rect 3127 701 3161 735
rect 3199 701 3233 735
rect 3548 701 3582 735
rect 3620 701 3654 735
rect 3692 701 3726 735
rect 3261 79 3295 113
rect 3333 79 3367 113
rect 3548 79 3582 113
rect 3620 79 3654 113
rect 3692 79 3726 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
<< metal1 >>
rect 0 831 3840 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3840 831
rect 0 791 3840 797
rect 0 737 3840 763
rect 0 735 1999 737
rect 0 701 290 735
rect 324 701 362 735
rect 396 701 434 735
rect 468 701 747 735
rect 781 701 819 735
rect 853 701 891 735
rect 925 701 1487 735
rect 1521 701 1559 735
rect 1593 701 1631 735
rect 1665 703 1999 735
rect 2033 703 2071 737
rect 2105 703 2143 737
rect 2177 735 3840 737
rect 2177 703 2609 735
rect 1665 701 2609 703
rect 2643 701 2681 735
rect 2715 701 2753 735
rect 2787 701 3055 735
rect 3089 701 3127 735
rect 3161 701 3199 735
rect 3233 701 3548 735
rect 3582 701 3620 735
rect 3654 701 3692 735
rect 3726 701 3840 735
rect 0 689 3840 701
rect 883 498 941 504
rect 883 464 895 498
rect 929 495 941 498
rect 1651 498 1709 504
rect 1651 495 1663 498
rect 929 467 1663 495
rect 929 464 941 467
rect 883 458 941 464
rect 1651 464 1663 467
rect 1697 495 1709 498
rect 2803 498 2861 504
rect 2803 495 2815 498
rect 1697 467 2815 495
rect 1697 464 1709 467
rect 1651 458 1709 464
rect 2803 464 2815 467
rect 2849 464 2861 498
rect 2803 458 2861 464
rect 0 113 3840 125
rect 0 79 837 113
rect 871 79 909 113
rect 943 79 981 113
rect 1015 79 1629 113
rect 1663 79 1701 113
rect 1735 79 1773 113
rect 1807 79 1974 113
rect 2008 79 2046 113
rect 2080 79 2623 113
rect 2657 79 2695 113
rect 2729 79 2767 113
rect 2801 79 3261 113
rect 3295 79 3333 113
rect 3367 79 3548 113
rect 3582 79 3620 113
rect 3654 79 3692 113
rect 3726 79 3840 113
rect 0 51 3840 79
rect 0 17 3840 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3840 17
rect 0 -23 3840 -17
<< labels >>
rlabel locali s 3097 391 3228 499 6 CLK
port 1 nsew clock input
rlabel locali s 582 532 641 652 6 D
port 2 nsew signal input
rlabel metal1 s 2803 458 2861 467 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1651 458 1709 467 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 883 458 941 467 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 883 467 2861 495 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 2803 495 2861 504 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 1651 495 1709 504 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 883 495 941 504 6 RESET_B
port 3 nsew signal input
rlabel locali s 21 236 223 302 6 SCD
port 4 nsew signal input
rlabel locali s 601 310 1127 367 6 SCE
port 5 nsew signal input
rlabel locali s 399 289 449 367 6 SCE
port 5 nsew signal input
rlabel locali s 976 367 1127 505 6 SCE
port 5 nsew signal input
rlabel locali s 399 367 635 401 6 SCE
port 5 nsew signal input
rlabel locali s 399 401 476 515 6 SCE
port 5 nsew signal input
rlabel metal1 s 0 51 3840 125 6 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 -23 3840 23 8 VNB
port 7 nsew ground bidirectional
rlabel pwell s -26 -43 3866 43 8 VNB
port 7 nsew ground bidirectional
rlabel pwell s 111 43 3836 221 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 3399 221 3836 283 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 111 221 3125 236 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1843 236 3125 291 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 791 3840 837 6 VPB
port 8 nsew power bidirectional
rlabel nwell s -66 377 3906 897 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 689 3840 763 6 VPWR
port 9 nsew power bidirectional
rlabel locali s 3764 103 3815 751 6 Q
port 10 nsew signal output
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 3840 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 444346
string GDS_START 407998
<< end >>
