VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AOAI4X1
  CLASS CORE ;
  FOREIGN AOAI4X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.990 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN YN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.351900 ;
    PORT
      LAYER li1 ;
        RECT 7.805 5.285 7.975 7.020 ;
        RECT 8.685 5.285 8.855 7.020 ;
        RECT 7.805 5.115 9.335 5.285 ;
        RECT 9.165 1.740 9.335 5.115 ;
        RECT 8.725 1.570 9.335 1.740 ;
        RECT 8.725 0.835 8.895 1.570 ;
    END
  END YN
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.033250 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.915 1.195 4.865 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 1.795 4.710 1.965 4.865 ;
        RECT 1.765 4.535 1.965 4.710 ;
        RECT 1.765 1.915 1.935 4.535 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.026450 ;
    PORT
      LAYER li1 ;
        RECT 5.130 4.710 5.300 4.870 ;
        RECT 5.095 4.540 5.300 4.710 ;
        RECT 5.095 1.915 5.265 4.540 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.027250 ;
    PORT
      LAYER li1 ;
        RECT 8.455 4.710 8.625 4.865 ;
        RECT 8.425 4.535 8.625 4.710 ;
        RECT 8.425 1.915 8.595 4.535 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 10.425 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 10.160 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.135 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.555 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 4.475 5.555 4.645 7.230 ;
        RECT 6.490 4.110 6.830 7.230 ;
        RECT 7.365 5.135 7.535 7.230 ;
        RECT 8.245 5.555 8.415 7.230 ;
        RECT 9.125 5.555 9.295 7.230 ;
        RECT 9.820 4.110 10.160 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 10.160 7.570 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 10.160 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 3.940 0.615 4.110 1.745 ;
        RECT 4.910 0.615 5.080 1.390 ;
        RECT 5.880 0.615 6.050 1.390 ;
        RECT 3.940 0.445 6.050 0.615 ;
        RECT 3.940 0.170 4.110 0.445 ;
        RECT 4.425 0.170 4.595 0.445 ;
        RECT 4.910 0.170 5.080 0.445 ;
        RECT 5.395 0.170 5.565 0.445 ;
        RECT 5.880 0.170 6.050 0.445 ;
        RECT 6.490 0.170 6.830 2.720 ;
        RECT 7.755 0.170 7.925 1.120 ;
        RECT 9.820 0.170 10.160 2.720 ;
        RECT -0.170 -0.170 10.160 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 10.160 0.170 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 1.145 5.285 1.315 7.020 ;
        RECT 2.025 5.285 2.195 7.020 ;
        RECT 4.035 5.295 4.205 7.025 ;
        RECT 4.915 6.825 5.965 6.995 ;
        RECT 4.915 5.295 5.085 6.825 ;
        RECT 1.145 5.115 2.675 5.285 ;
        RECT 4.035 5.125 5.085 5.295 ;
        RECT 5.355 5.295 5.525 6.565 ;
        RECT 5.795 5.555 5.965 6.825 ;
        RECT 5.355 5.125 6.005 5.295 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 2.505 1.740 2.675 5.115 ;
        RECT 4.200 4.710 4.370 4.870 ;
        RECT 4.200 4.540 4.525 4.710 ;
        RECT 4.355 1.915 4.525 4.540 ;
        RECT 5.835 1.740 6.005 5.125 ;
        RECT 7.685 1.915 7.855 4.865 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.065 1.570 2.675 1.740 ;
        RECT 4.425 1.570 6.005 1.740 ;
        RECT 7.270 1.665 7.440 1.745 ;
        RECT 8.240 1.665 8.410 1.745 ;
        RECT 2.065 0.835 2.235 1.570 ;
        RECT 2.550 0.615 2.720 1.385 ;
        RECT 4.425 0.835 4.595 1.570 ;
        RECT 5.395 0.835 5.565 1.570 ;
        RECT 7.270 1.495 8.410 1.665 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
        RECT 7.270 0.365 7.440 1.495 ;
        RECT 8.240 0.615 8.410 1.495 ;
        RECT 9.210 0.615 9.380 1.385 ;
        RECT 8.240 0.445 9.380 0.615 ;
        RECT 8.240 0.365 8.410 0.445 ;
        RECT 9.210 0.365 9.380 0.445 ;
      LAYER mcon ;
        RECT 2.505 2.505 2.675 2.675 ;
        RECT 4.355 2.505 4.525 2.675 ;
        RECT 5.835 2.505 6.005 2.675 ;
        RECT 7.685 2.505 7.855 2.675 ;
      LAYER met1 ;
        RECT 2.475 2.675 2.705 2.705 ;
        RECT 4.325 2.675 4.555 2.705 ;
        RECT 5.805 2.675 6.035 2.705 ;
        RECT 7.655 2.675 7.885 2.705 ;
        RECT 2.445 2.505 4.585 2.675 ;
        RECT 5.775 2.505 7.915 2.675 ;
        RECT 2.475 2.475 2.705 2.505 ;
        RECT 4.325 2.475 4.555 2.505 ;
        RECT 5.805 2.475 6.035 2.505 ;
        RECT 7.655 2.475 7.885 2.505 ;
  END
END AOAI4X1
END LIBRARY

