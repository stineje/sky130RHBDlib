* SPICE3 file created from AND3X1.ext - technology: sky130A

.subckt AND3X1 Y A B C VDD VSS
X0 VDD B a_277_1050 VDD sky130_fd_pr__pfet_01v8 ad=0.00336 pd=2.736 as=0 ps=0 w=2 l=0.15 M=2
X1 VDD C a_277_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X2 Y a_277_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0058 pd=4.58 as=0 ps=0 w=2 l=0.15 M=2
X3 a_277_1050 C a_372_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X4 a_277_1050 A VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X5 VSS A a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0.0013199 pd=9.67 as=0 ps=0 w=3 l=0.15
X6 a_372_210 B a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X7 Y a_277_1050 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0 ps=0 w=3 l=0.15
C0 VDD a_277_1050 2.88f
C1 VDD VSS 2.51f
.ends
