magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 19 21 917 203
rect 29 -17 63 21
<< locali >>
rect 121 51 179 478
rect 392 265 451 471
rect 377 199 451 265
rect 485 199 547 471
rect 581 199 639 348
rect 673 191 755 348
rect 789 199 903 348
rect 701 165 755 191
rect 701 58 799 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 327 87 527
rect 17 17 87 177
rect 213 299 263 527
rect 299 299 357 493
rect 299 265 341 299
rect 213 215 341 265
rect 213 89 265 173
rect 299 157 341 215
rect 614 417 680 493
rect 718 451 784 527
rect 818 417 903 493
rect 614 383 903 417
rect 299 123 667 157
rect 213 17 402 89
rect 436 51 484 123
rect 518 17 584 89
rect 618 51 667 123
rect 833 17 903 161
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 701 58 799 165 6 A1
port 1 nsew signal input
rlabel locali s 701 165 755 191 6 A1
port 1 nsew signal input
rlabel locali s 673 191 755 348 6 A1
port 1 nsew signal input
rlabel locali s 789 199 903 348 6 A2
port 2 nsew signal input
rlabel locali s 581 199 639 348 6 B1
port 3 nsew signal input
rlabel locali s 485 199 547 471 6 C1
port 4 nsew signal input
rlabel locali s 377 199 451 265 6 D1
port 5 nsew signal input
rlabel locali s 392 265 451 471 6 D1
port 5 nsew signal input
rlabel metal1 s 0 -48 920 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 19 21 917 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 121 51 179 478 6 X
port 10 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 3763378
string GDS_START 3754318
<< end >>
