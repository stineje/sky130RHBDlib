* SPICE3 file created from TMRDFFSNQNX1.ext - technology: sky130A

.subckt TMRDFFSNQNX1 QN D CLK SN
X0  m1_13561_871# votern3x1_pcell_0/nmos_top_0/a_0_0#  nshort w=3 l=0.15
X1  m1_13561_871# votern3x1_pcell_0/nmos_bottom_1/a_0_0#  nshort w=3 l=0.15
X2  m1_4152_649# votern3x1_pcell_0/nmos_bottom_2/a_0_0#  nshort w=3 l=0.15
X3 votern3x1_pcell_0/a_805_1331# m1_13561_871#   pshort w=2 l=0.15
X4 QN m1_4152_649# votern3x1_pcell_0/nmos_bottom_1/a_0_0#  nshort w=3 l=0.15
X5 votern3x1_pcell_0/a_805_1331# m1_9056_501#   pshort w=2 l=0.15
X6 votern3x1_pcell_0/a_893_1059# m1_4152_649# votern3x1_pcell_0/a_805_1331#  pshort w=2 l=0.15
X7 votern3x1_pcell_0/a_893_1059# m1_13561_871# votern3x1_pcell_0/a_805_1331#  pshort w=2 l=0.15
X8 QN m1_4152_649# votern3x1_pcell_0/a_893_1059#  pshort w=2 l=0.15
X9 QN m1_9056_501# votern3x1_pcell_0/a_893_1059#  pshort w=2 l=0.15
X10 QN m1_9056_501# votern3x1_pcell_0/nmos_top_0/a_0_0#  nshort w=3 l=0.15
X11 QN m1_9056_501# votern3x1_pcell_0/nmos_bottom_2/a_0_0#  nshort w=3 l=0.15
X12  dffsnx1_pcell_1/m1_406_797# dffsnx1_pcell_1/nand2x1_pcell_2/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X13 m1_9056_501# m1_8522_797# dffsnx1_pcell_1/nand2x1_pcell_2/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X14  dffsnx1_pcell_1/m1_406_797# m1_9056_501#  pshort w=2 l=0.15
X15  m1_8522_797# m1_9056_501#  pshort w=2 l=0.15
X16  D dffsnx1_pcell_1/nand2x1_pcell_5/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X17 dffsnx1_pcell_1/m1_537_501# dffsnx1_pcell_1/m1_406_797# dffsnx1_pcell_1/nand2x1_pcell_5/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X18  D dffsnx1_pcell_1/m1_537_501#  pshort w=2 l=0.15
X19  dffsnx1_pcell_1/m1_406_797# dffsnx1_pcell_1/m1_537_501#  pshort w=2 l=0.15
X20  dffsnx1_pcell_1/m1_537_501# dffsnx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X21 dffsnx1_pcell_1/m1_406_797# dffsnx1_pcell_1/m1_1351_723# dffsnx1_pcell_1/nand3x1_pcell_0/li_393_182#  nshort w=3 l=0.15
X22 dffsnx1_pcell_1/nand3x1_pcell_0/li_393_182# CLK dffsnx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X23  dffsnx1_pcell_1/m1_537_501# dffsnx1_pcell_1/m1_406_797#  pshort w=2 l=0.15
X24  CLK dffsnx1_pcell_1/m1_406_797#  pshort w=2 l=0.15
X25  dffsnx1_pcell_1/m1_1351_723# dffsnx1_pcell_1/m1_406_797#  pshort w=2 l=0.15
X26  m1_9056_501# dffsnx1_pcell_1/nand3x1_pcell_1/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X27 m1_8522_797# dffsnx1_pcell_1/m1_1351_723# dffsnx1_pcell_1/nand3x1_pcell_1/li_393_182#  nshort w=3 l=0.15
X28 dffsnx1_pcell_1/nand3x1_pcell_1/li_393_182# SN dffsnx1_pcell_1/nand3x1_pcell_1/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X29  m1_9056_501# m1_8522_797#  pshort w=2 l=0.15
X30  SN m1_8522_797#  pshort w=2 l=0.15
X31  dffsnx1_pcell_1/m1_1351_723# m1_8522_797#  pshort w=2 l=0.15
X32  dffsnx1_pcell_1/m1_537_501# dffsnx1_pcell_1/nand3x1_pcell_2/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X33 dffsnx1_pcell_1/m1_2461_501# dffsnx1_pcell_1/m1_1351_723# dffsnx1_pcell_1/nand3x1_pcell_2/li_393_182#  nshort w=3 l=0.15
X34 dffsnx1_pcell_1/nand3x1_pcell_2/li_393_182# SN dffsnx1_pcell_1/nand3x1_pcell_2/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X35  dffsnx1_pcell_1/m1_537_501# dffsnx1_pcell_1/m1_2461_501#  pshort w=2 l=0.15
X36  SN dffsnx1_pcell_1/m1_2461_501#  pshort w=2 l=0.15
X37  dffsnx1_pcell_1/m1_1351_723# dffsnx1_pcell_1/m1_2461_501#  pshort w=2 l=0.15
X38  dffsnx1_pcell_1/m1_2461_501# dffsnx1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X39 dffsnx1_pcell_1/m1_1351_723# CLK dffsnx1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X40  dffsnx1_pcell_1/m1_2461_501# dffsnx1_pcell_1/m1_1351_723#  pshort w=2 l=0.15
X41  CLK dffsnx1_pcell_1/m1_1351_723#  pshort w=2 l=0.15
X42  dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X43 m1_4152_649# m1_3606_797# dffsnx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X44  dffsnx1_pcell_0/m1_406_797# m1_4152_649#  pshort w=2 l=0.15
X45  m1_3606_797# m1_4152_649#  pshort w=2 l=0.15
X46  D dffsnx1_pcell_0/nand2x1_pcell_5/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X47 dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/nand2x1_pcell_5/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X48  D dffsnx1_pcell_0/m1_537_501#  pshort w=2 l=0.15
X49  dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/m1_537_501#  pshort w=2 l=0.15
X50  dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X51 dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/nand3x1_pcell_0/li_393_182#  nshort w=3 l=0.15
X52 dffsnx1_pcell_0/nand3x1_pcell_0/li_393_182# CLK dffsnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X53  dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/m1_406_797#  pshort w=2 l=0.15
X54  CLK dffsnx1_pcell_0/m1_406_797#  pshort w=2 l=0.15
X55  dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/m1_406_797#  pshort w=2 l=0.15
X56  m1_4152_649# dffsnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X57 m1_3606_797# dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/nand3x1_pcell_1/li_393_182#  nshort w=3 l=0.15
X58 dffsnx1_pcell_0/nand3x1_pcell_1/li_393_182# SN dffsnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X59  m1_4152_649# m1_3606_797#  pshort w=2 l=0.15
X60  SN m1_3606_797#  pshort w=2 l=0.15
X61  dffsnx1_pcell_0/m1_1351_723# m1_3606_797#  pshort w=2 l=0.15
X62  dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/nand3x1_pcell_2/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X63 dffsnx1_pcell_0/m1_2461_501# dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/nand3x1_pcell_2/li_393_182#  nshort w=3 l=0.15
X64 dffsnx1_pcell_0/nand3x1_pcell_2/li_393_182# SN dffsnx1_pcell_0/nand3x1_pcell_2/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X65  dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/m1_2461_501#  pshort w=2 l=0.15
X66  SN dffsnx1_pcell_0/m1_2461_501#  pshort w=2 l=0.15
X67  dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/m1_2461_501#  pshort w=2 l=0.15
X68  dffsnx1_pcell_0/m1_2461_501# dffsnx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X69 dffsnx1_pcell_0/m1_1351_723# CLK dffsnx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X70  dffsnx1_pcell_0/m1_2461_501# dffsnx1_pcell_0/m1_1351_723#  pshort w=2 l=0.15
X71  CLK dffsnx1_pcell_0/m1_1351_723#  pshort w=2 l=0.15
X72  dffsnx1_pcell_2/m1_406_797# dffsnx1_pcell_2/nand2x1_pcell_2/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X73 m1_13561_871# m1_13413_797# dffsnx1_pcell_2/nand2x1_pcell_2/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X74  dffsnx1_pcell_2/m1_406_797# m1_13561_871#  pshort w=2 l=0.15
X75  m1_13413_797# m1_13561_871#  pshort w=2 l=0.15
X76  D dffsnx1_pcell_2/nand2x1_pcell_5/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X77 dffsnx1_pcell_2/m1_537_501# dffsnx1_pcell_2/m1_406_797# dffsnx1_pcell_2/nand2x1_pcell_5/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X78  D dffsnx1_pcell_2/m1_537_501#  pshort w=2 l=0.15
X79  dffsnx1_pcell_2/m1_406_797# dffsnx1_pcell_2/m1_537_501#  pshort w=2 l=0.15
X80  dffsnx1_pcell_2/m1_537_501# dffsnx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X81 dffsnx1_pcell_2/m1_406_797# dffsnx1_pcell_2/m1_1351_723# dffsnx1_pcell_2/nand3x1_pcell_0/li_393_182#  nshort w=3 l=0.15
X82 dffsnx1_pcell_2/nand3x1_pcell_0/li_393_182# CLK dffsnx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X83  dffsnx1_pcell_2/m1_537_501# dffsnx1_pcell_2/m1_406_797#  pshort w=2 l=0.15
X84  CLK dffsnx1_pcell_2/m1_406_797#  pshort w=2 l=0.15
X85  dffsnx1_pcell_2/m1_1351_723# dffsnx1_pcell_2/m1_406_797#  pshort w=2 l=0.15
X86  m1_13561_871# dffsnx1_pcell_2/nand3x1_pcell_1/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X87 m1_13413_797# dffsnx1_pcell_2/m1_1351_723# dffsnx1_pcell_2/nand3x1_pcell_1/li_393_182#  nshort w=3 l=0.15
X88 dffsnx1_pcell_2/nand3x1_pcell_1/li_393_182# SN dffsnx1_pcell_2/nand3x1_pcell_1/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X89  m1_13561_871# m1_13413_797#  pshort w=2 l=0.15
X90  SN m1_13413_797#  pshort w=2 l=0.15
X91  dffsnx1_pcell_2/m1_1351_723# m1_13413_797#  pshort w=2 l=0.15
X92  dffsnx1_pcell_2/m1_537_501# dffsnx1_pcell_2/nand3x1_pcell_2/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X93 dffsnx1_pcell_2/m1_2461_501# dffsnx1_pcell_2/m1_1351_723# dffsnx1_pcell_2/nand3x1_pcell_2/li_393_182#  nshort w=3 l=0.15
X94 dffsnx1_pcell_2/nand3x1_pcell_2/li_393_182# SN dffsnx1_pcell_2/nand3x1_pcell_2/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X95  dffsnx1_pcell_2/m1_537_501# dffsnx1_pcell_2/m1_2461_501#  pshort w=2 l=0.15
X96  SN dffsnx1_pcell_2/m1_2461_501#  pshort w=2 l=0.15
X97  dffsnx1_pcell_2/m1_1351_723# dffsnx1_pcell_2/m1_2461_501#  pshort w=2 l=0.15
X98  dffsnx1_pcell_2/m1_2461_501# dffsnx1_pcell_2/nand2x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X99 dffsnx1_pcell_2/m1_1351_723# CLK dffsnx1_pcell_2/nand2x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X100  dffsnx1_pcell_2/m1_2461_501# dffsnx1_pcell_2/m1_1351_723#  pshort w=2 l=0.15
X101  CLK dffsnx1_pcell_2/m1_1351_723#  pshort w=2 l=0.15
C0 CLK  4.72fF
.ends
