magic
tech sky130A
magscale 1 2
timestamp 1669200967
<< nwell >>
rect -87 786 1863 1550
<< pwell >>
rect -34 -34 1810 544
<< nmos >>
rect 168 288 198 349
tri 198 288 214 304 sw
rect 362 296 392 349
tri 392 296 408 312 sw
rect 168 258 274 288
tri 274 258 304 288 sw
rect 362 266 468 296
tri 468 266 498 296 sw
rect 168 157 198 258
tri 198 242 214 258 nw
tri 258 242 274 258 ne
tri 198 157 214 173 sw
tri 258 157 274 173 se
rect 274 157 304 258
rect 362 165 392 266
tri 392 250 408 266 nw
tri 452 250 468 266 ne
tri 392 165 408 181 sw
tri 452 165 468 181 se
rect 468 165 498 266
tri 168 127 198 157 ne
rect 198 127 274 157
tri 274 127 304 157 nw
tri 362 135 392 165 ne
rect 392 135 468 165
tri 468 135 498 165 nw
rect 834 296 864 349
tri 864 296 880 312 sw
rect 1028 296 1058 349
tri 1058 296 1074 312 sw
rect 834 266 940 296
tri 940 266 970 296 sw
rect 834 165 864 266
tri 864 250 880 266 nw
tri 924 250 940 266 ne
tri 864 165 880 181 sw
tri 924 165 940 181 se
rect 940 165 970 266
rect 1028 266 1134 296
tri 1134 266 1164 296 sw
rect 1028 251 1059 266
tri 1059 251 1074 266 nw
tri 1118 251 1133 266 ne
rect 1133 251 1164 266
tri 834 135 864 165 ne
rect 864 135 940 165
tri 940 135 970 165 nw
rect 1028 165 1058 251
tri 1058 165 1074 181 sw
tri 1118 165 1134 181 se
rect 1134 165 1164 251
tri 1028 135 1058 165 ne
rect 1058 135 1134 165
tri 1134 135 1164 165 nw
rect 1487 297 1517 350
tri 1517 297 1533 313 sw
rect 1487 267 1593 297
tri 1593 267 1623 297 sw
rect 1487 166 1517 267
tri 1517 251 1533 267 nw
tri 1577 251 1593 267 ne
tri 1517 166 1533 182 sw
tri 1577 166 1593 182 se
rect 1593 166 1623 267
tri 1487 136 1517 166 ne
rect 1517 136 1593 166
tri 1593 136 1623 166 nw
<< pmos >>
rect 187 1004 217 1404
rect 275 1004 305 1404
rect 363 1004 393 1404
rect 451 1004 481 1404
rect 853 1005 883 1405
rect 941 1005 971 1405
rect 1029 1005 1059 1405
rect 1117 1005 1147 1405
rect 1496 1004 1526 1404
rect 1584 1004 1614 1404
<< ndiff >>
rect 112 333 168 349
rect 112 299 122 333
rect 156 299 168 333
rect 112 261 168 299
rect 198 333 362 349
rect 198 304 219 333
tri 198 288 214 304 ne
rect 214 299 219 304
rect 253 299 316 333
rect 350 299 362 333
rect 214 288 362 299
rect 392 312 554 349
tri 392 296 408 312 ne
rect 408 296 554 312
rect 112 227 122 261
rect 156 227 168 261
tri 274 258 304 288 ne
rect 304 261 362 288
tri 468 266 498 296 ne
rect 112 193 168 227
rect 112 159 122 193
rect 156 159 168 193
rect 112 127 168 159
tri 198 242 214 258 se
rect 214 242 258 258
tri 258 242 274 258 sw
rect 198 208 274 242
rect 198 174 219 208
rect 253 174 274 208
rect 198 173 274 174
tri 198 157 214 173 ne
rect 214 157 258 173
tri 258 157 274 173 nw
rect 304 227 316 261
rect 350 227 362 261
rect 304 193 362 227
rect 304 159 316 193
rect 350 159 362 193
tri 392 250 408 266 se
rect 408 250 452 266
tri 452 250 468 266 sw
rect 392 217 468 250
rect 392 183 413 217
rect 447 183 468 217
rect 392 181 468 183
tri 392 165 408 181 ne
rect 408 165 452 181
tri 452 165 468 181 nw
rect 498 261 554 296
rect 498 227 510 261
rect 544 227 554 261
rect 498 193 554 227
tri 168 127 198 157 sw
tri 274 127 304 157 se
rect 304 135 362 159
tri 362 135 392 165 sw
tri 468 135 498 165 se
rect 498 159 510 193
rect 544 159 554 193
rect 498 135 554 159
rect 304 127 554 135
rect 112 123 554 127
rect 112 89 122 123
rect 156 89 316 123
rect 350 89 413 123
rect 447 89 510 123
rect 544 89 554 123
rect 112 73 554 89
rect 778 333 834 349
rect 778 299 788 333
rect 822 299 834 333
rect 778 261 834 299
rect 864 312 1028 349
tri 864 296 880 312 ne
rect 880 296 1028 312
rect 1058 312 1220 349
tri 1058 296 1074 312 ne
rect 1074 296 1220 312
tri 940 266 970 296 ne
rect 778 227 788 261
rect 822 227 834 261
rect 778 193 834 227
rect 778 159 788 193
rect 822 159 834 193
tri 864 250 880 266 se
rect 880 250 924 266
tri 924 250 940 266 sw
rect 864 217 940 250
rect 864 183 885 217
rect 919 183 940 217
rect 864 181 940 183
tri 864 165 880 181 ne
rect 880 165 924 181
tri 924 165 940 181 nw
rect 970 261 1028 296
tri 1134 266 1164 296 ne
rect 970 227 982 261
rect 1016 227 1028 261
tri 1059 251 1074 266 se
rect 1074 251 1118 266
tri 1118 251 1133 266 sw
rect 1164 261 1220 296
rect 970 193 1028 227
rect 778 135 834 159
tri 834 135 864 165 sw
tri 940 135 970 165 se
rect 970 159 982 193
rect 1016 159 1028 193
rect 1058 217 1134 251
rect 1058 183 1079 217
rect 1113 183 1134 217
rect 1058 181 1134 183
tri 1058 165 1074 181 ne
rect 1074 165 1118 181
tri 1118 165 1134 181 nw
rect 1164 227 1176 261
rect 1210 227 1220 261
rect 1164 193 1220 227
rect 970 135 1028 159
tri 1028 135 1058 165 sw
tri 1134 135 1164 165 se
rect 1164 159 1176 193
rect 1210 159 1220 193
rect 1164 135 1220 159
rect 778 123 1220 135
rect 778 89 788 123
rect 822 89 885 123
rect 919 89 982 123
rect 1016 89 1079 123
rect 1113 89 1176 123
rect 1210 89 1220 123
rect 778 73 1220 89
rect 1431 334 1487 350
rect 1431 300 1441 334
rect 1475 300 1487 334
rect 1431 262 1487 300
rect 1517 334 1677 350
rect 1517 313 1635 334
tri 1517 297 1533 313 ne
rect 1533 300 1635 313
rect 1669 300 1677 334
rect 1533 297 1677 300
tri 1593 267 1623 297 ne
rect 1431 228 1441 262
rect 1475 228 1487 262
rect 1431 194 1487 228
rect 1431 160 1441 194
rect 1475 160 1487 194
tri 1517 251 1533 267 se
rect 1533 251 1577 267
tri 1577 251 1593 267 sw
rect 1517 218 1593 251
rect 1517 184 1537 218
rect 1571 184 1593 218
rect 1517 182 1593 184
tri 1517 166 1533 182 ne
rect 1533 166 1577 182
tri 1577 166 1593 182 nw
rect 1623 262 1677 297
rect 1623 228 1635 262
rect 1669 228 1677 262
rect 1623 194 1677 228
rect 1431 136 1487 160
tri 1487 136 1517 166 sw
tri 1593 136 1623 166 se
rect 1623 160 1635 194
rect 1669 160 1677 194
rect 1623 136 1677 160
rect 1431 124 1677 136
rect 1431 90 1441 124
rect 1475 90 1537 124
rect 1571 90 1635 124
rect 1669 90 1677 124
rect 1431 74 1677 90
<< pdiff >>
rect 131 1366 187 1404
rect 131 1332 141 1366
rect 175 1332 187 1366
rect 131 1298 187 1332
rect 131 1264 141 1298
rect 175 1264 187 1298
rect 131 1230 187 1264
rect 131 1196 141 1230
rect 175 1196 187 1230
rect 131 1162 187 1196
rect 131 1128 141 1162
rect 175 1128 187 1162
rect 131 1093 187 1128
rect 131 1059 141 1093
rect 175 1059 187 1093
rect 131 1004 187 1059
rect 217 1366 275 1404
rect 217 1332 229 1366
rect 263 1332 275 1366
rect 217 1298 275 1332
rect 217 1264 229 1298
rect 263 1264 275 1298
rect 217 1230 275 1264
rect 217 1196 229 1230
rect 263 1196 275 1230
rect 217 1162 275 1196
rect 217 1128 229 1162
rect 263 1128 275 1162
rect 217 1093 275 1128
rect 217 1059 229 1093
rect 263 1059 275 1093
rect 217 1004 275 1059
rect 305 1366 363 1404
rect 305 1332 317 1366
rect 351 1332 363 1366
rect 305 1298 363 1332
rect 305 1264 317 1298
rect 351 1264 363 1298
rect 305 1230 363 1264
rect 305 1196 317 1230
rect 351 1196 363 1230
rect 305 1162 363 1196
rect 305 1128 317 1162
rect 351 1128 363 1162
rect 305 1004 363 1128
rect 393 1366 451 1404
rect 393 1332 405 1366
rect 439 1332 451 1366
rect 393 1298 451 1332
rect 393 1264 405 1298
rect 439 1264 451 1298
rect 393 1230 451 1264
rect 393 1196 405 1230
rect 439 1196 451 1230
rect 393 1162 451 1196
rect 393 1128 405 1162
rect 439 1128 451 1162
rect 393 1093 451 1128
rect 393 1059 405 1093
rect 439 1059 451 1093
rect 393 1004 451 1059
rect 481 1366 535 1404
rect 481 1332 493 1366
rect 527 1332 535 1366
rect 481 1298 535 1332
rect 481 1264 493 1298
rect 527 1264 535 1298
rect 481 1230 535 1264
rect 481 1196 493 1230
rect 527 1196 535 1230
rect 481 1162 535 1196
rect 481 1128 493 1162
rect 527 1128 535 1162
rect 481 1004 535 1128
rect 797 1365 853 1405
rect 797 1331 807 1365
rect 841 1331 853 1365
rect 797 1297 853 1331
rect 797 1263 807 1297
rect 841 1263 853 1297
rect 797 1229 853 1263
rect 797 1195 807 1229
rect 841 1195 853 1229
rect 797 1161 853 1195
rect 797 1127 807 1161
rect 841 1127 853 1161
rect 797 1093 853 1127
rect 797 1059 807 1093
rect 841 1059 853 1093
rect 797 1005 853 1059
rect 883 1365 941 1405
rect 883 1331 895 1365
rect 929 1331 941 1365
rect 883 1297 941 1331
rect 883 1263 895 1297
rect 929 1263 941 1297
rect 883 1229 941 1263
rect 883 1195 895 1229
rect 929 1195 941 1229
rect 883 1161 941 1195
rect 883 1127 895 1161
rect 929 1127 941 1161
rect 883 1005 941 1127
rect 971 1365 1029 1405
rect 971 1331 983 1365
rect 1017 1331 1029 1365
rect 971 1297 1029 1331
rect 971 1263 983 1297
rect 1017 1263 1029 1297
rect 971 1229 1029 1263
rect 971 1195 983 1229
rect 1017 1195 1029 1229
rect 971 1161 1029 1195
rect 971 1127 983 1161
rect 1017 1127 1029 1161
rect 971 1093 1029 1127
rect 971 1059 983 1093
rect 1017 1059 1029 1093
rect 971 1005 1029 1059
rect 1059 1297 1117 1405
rect 1059 1263 1071 1297
rect 1105 1263 1117 1297
rect 1059 1229 1117 1263
rect 1059 1195 1071 1229
rect 1105 1195 1117 1229
rect 1059 1161 1117 1195
rect 1059 1127 1071 1161
rect 1105 1127 1117 1161
rect 1059 1093 1117 1127
rect 1059 1059 1071 1093
rect 1105 1059 1117 1093
rect 1059 1005 1117 1059
rect 1147 1365 1201 1405
rect 1147 1331 1159 1365
rect 1193 1331 1201 1365
rect 1147 1297 1201 1331
rect 1147 1263 1159 1297
rect 1193 1263 1201 1297
rect 1147 1229 1201 1263
rect 1147 1195 1159 1229
rect 1193 1195 1201 1229
rect 1147 1161 1201 1195
rect 1147 1127 1159 1161
rect 1193 1127 1201 1161
rect 1147 1005 1201 1127
rect 1440 1366 1496 1404
rect 1440 1332 1450 1366
rect 1484 1332 1496 1366
rect 1440 1298 1496 1332
rect 1440 1264 1450 1298
rect 1484 1264 1496 1298
rect 1440 1230 1496 1264
rect 1440 1196 1450 1230
rect 1484 1196 1496 1230
rect 1440 1162 1496 1196
rect 1440 1128 1450 1162
rect 1484 1128 1496 1162
rect 1440 1093 1496 1128
rect 1440 1059 1450 1093
rect 1484 1059 1496 1093
rect 1440 1004 1496 1059
rect 1526 1366 1584 1404
rect 1526 1332 1538 1366
rect 1572 1332 1584 1366
rect 1526 1298 1584 1332
rect 1526 1264 1538 1298
rect 1572 1264 1584 1298
rect 1526 1230 1584 1264
rect 1526 1196 1538 1230
rect 1572 1196 1584 1230
rect 1526 1162 1584 1196
rect 1526 1128 1538 1162
rect 1572 1128 1584 1162
rect 1526 1093 1584 1128
rect 1526 1059 1538 1093
rect 1572 1059 1584 1093
rect 1526 1004 1584 1059
rect 1614 1366 1668 1404
rect 1614 1332 1626 1366
rect 1660 1332 1668 1366
rect 1614 1298 1668 1332
rect 1614 1264 1626 1298
rect 1660 1264 1668 1298
rect 1614 1230 1668 1264
rect 1614 1196 1626 1230
rect 1660 1196 1668 1230
rect 1614 1162 1668 1196
rect 1614 1128 1626 1162
rect 1660 1128 1668 1162
rect 1614 1093 1668 1128
rect 1614 1059 1626 1093
rect 1660 1059 1668 1093
rect 1614 1004 1668 1059
<< ndiffc >>
rect 122 299 156 333
rect 219 299 253 333
rect 316 299 350 333
rect 122 227 156 261
rect 122 159 156 193
rect 219 174 253 208
rect 316 227 350 261
rect 316 159 350 193
rect 413 183 447 217
rect 510 227 544 261
rect 510 159 544 193
rect 122 89 156 123
rect 316 89 350 123
rect 413 89 447 123
rect 510 89 544 123
rect 788 299 822 333
rect 788 227 822 261
rect 788 159 822 193
rect 885 183 919 217
rect 982 227 1016 261
rect 982 159 1016 193
rect 1079 183 1113 217
rect 1176 227 1210 261
rect 1176 159 1210 193
rect 788 89 822 123
rect 885 89 919 123
rect 982 89 1016 123
rect 1079 89 1113 123
rect 1176 89 1210 123
rect 1441 300 1475 334
rect 1635 300 1669 334
rect 1441 228 1475 262
rect 1441 160 1475 194
rect 1537 184 1571 218
rect 1635 228 1669 262
rect 1635 160 1669 194
rect 1441 90 1475 124
rect 1537 90 1571 124
rect 1635 90 1669 124
<< pdiffc >>
rect 141 1332 175 1366
rect 141 1264 175 1298
rect 141 1196 175 1230
rect 141 1128 175 1162
rect 141 1059 175 1093
rect 229 1332 263 1366
rect 229 1264 263 1298
rect 229 1196 263 1230
rect 229 1128 263 1162
rect 229 1059 263 1093
rect 317 1332 351 1366
rect 317 1264 351 1298
rect 317 1196 351 1230
rect 317 1128 351 1162
rect 405 1332 439 1366
rect 405 1264 439 1298
rect 405 1196 439 1230
rect 405 1128 439 1162
rect 405 1059 439 1093
rect 493 1332 527 1366
rect 493 1264 527 1298
rect 493 1196 527 1230
rect 493 1128 527 1162
rect 807 1331 841 1365
rect 807 1263 841 1297
rect 807 1195 841 1229
rect 807 1127 841 1161
rect 807 1059 841 1093
rect 895 1331 929 1365
rect 895 1263 929 1297
rect 895 1195 929 1229
rect 895 1127 929 1161
rect 983 1331 1017 1365
rect 983 1263 1017 1297
rect 983 1195 1017 1229
rect 983 1127 1017 1161
rect 983 1059 1017 1093
rect 1071 1263 1105 1297
rect 1071 1195 1105 1229
rect 1071 1127 1105 1161
rect 1071 1059 1105 1093
rect 1159 1331 1193 1365
rect 1159 1263 1193 1297
rect 1159 1195 1193 1229
rect 1159 1127 1193 1161
rect 1450 1332 1484 1366
rect 1450 1264 1484 1298
rect 1450 1196 1484 1230
rect 1450 1128 1484 1162
rect 1450 1059 1484 1093
rect 1538 1332 1572 1366
rect 1538 1264 1572 1298
rect 1538 1196 1572 1230
rect 1538 1128 1572 1162
rect 1538 1059 1572 1093
rect 1626 1332 1660 1366
rect 1626 1264 1660 1298
rect 1626 1196 1660 1230
rect 1626 1128 1660 1162
rect 1626 1059 1660 1093
<< psubdiff >>
rect -34 482 1810 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 632 461 700 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 632 427 649 461
rect 683 427 700 461
rect 1298 461 1366 482
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 632 313 700 353
rect 1298 427 1315 461
rect 1349 427 1366 461
rect 1742 461 1810 482
rect 1298 387 1366 427
rect 1298 353 1315 387
rect 1349 353 1366 387
rect 1742 427 1759 461
rect 1793 427 1810 461
rect 632 279 649 313
rect 683 279 700 313
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect -34 17 34 57
rect 632 57 649 91
rect 683 57 700 91
rect 1298 313 1366 353
rect 1742 387 1810 427
rect 1742 353 1759 387
rect 1793 353 1810 387
rect 1298 279 1315 313
rect 1349 279 1366 313
rect 1298 239 1366 279
rect 1298 205 1315 239
rect 1349 205 1366 239
rect 1298 165 1366 205
rect 1298 131 1315 165
rect 1349 131 1366 165
rect 1298 91 1366 131
rect 632 17 700 57
rect 1298 57 1315 91
rect 1349 57 1366 91
rect 1742 313 1810 353
rect 1742 279 1759 313
rect 1793 279 1810 313
rect 1742 239 1810 279
rect 1742 205 1759 239
rect 1793 205 1810 239
rect 1742 165 1810 205
rect 1742 131 1759 165
rect 1793 131 1810 165
rect 1742 91 1810 131
rect 1298 17 1366 57
rect 1742 57 1759 91
rect 1793 57 1810 91
rect 1742 17 1810 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1810 17
rect -34 -34 1810 -17
<< nsubdiff >>
rect -34 1497 1810 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1810 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 632 1423 700 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 1298 1423 1366 1463
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 632 979 700 1019
rect 1298 1389 1315 1423
rect 1349 1389 1366 1423
rect 1742 1423 1810 1463
rect 1298 1349 1366 1389
rect 1298 1315 1315 1349
rect 1349 1315 1366 1349
rect 1298 1275 1366 1315
rect 1298 1241 1315 1275
rect 1349 1241 1366 1275
rect 1298 1201 1366 1241
rect 1298 1167 1315 1201
rect 1349 1167 1366 1201
rect 1298 1127 1366 1167
rect 1298 1093 1315 1127
rect 1349 1093 1366 1127
rect 1298 1053 1366 1093
rect 1298 1019 1315 1053
rect 1349 1019 1366 1053
rect 632 945 649 979
rect 683 945 700 979
rect -34 871 -17 905
rect 17 884 34 905
rect 632 905 700 945
rect 1298 979 1366 1019
rect 1742 1389 1759 1423
rect 1793 1389 1810 1423
rect 1742 1349 1810 1389
rect 1742 1315 1759 1349
rect 1793 1315 1810 1349
rect 1742 1275 1810 1315
rect 1742 1241 1759 1275
rect 1793 1241 1810 1275
rect 1742 1201 1810 1241
rect 1742 1167 1759 1201
rect 1793 1167 1810 1201
rect 1742 1127 1810 1167
rect 1742 1093 1759 1127
rect 1793 1093 1810 1127
rect 1742 1053 1810 1093
rect 1742 1019 1759 1053
rect 1793 1019 1810 1053
rect 1298 945 1315 979
rect 1349 945 1366 979
rect 632 884 649 905
rect 17 871 649 884
rect 683 884 700 905
rect 1298 905 1366 945
rect 1742 979 1810 1019
rect 1742 945 1759 979
rect 1793 945 1810 979
rect 1298 884 1315 905
rect 683 871 1315 884
rect 1349 884 1366 905
rect 1742 905 1810 945
rect 1742 884 1759 905
rect 1349 871 1759 884
rect 1793 871 1810 905
rect -34 822 1810 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 649 427 683 461
rect 649 353 683 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1315 427 1349 461
rect 1315 353 1349 387
rect 1759 427 1793 461
rect 649 279 683 313
rect 649 205 683 239
rect 649 131 683 165
rect 649 57 683 91
rect 1759 353 1793 387
rect 1315 279 1349 313
rect 1315 205 1349 239
rect 1315 131 1349 165
rect 1315 57 1349 91
rect 1759 279 1793 313
rect 1759 205 1793 239
rect 1759 131 1793 165
rect 1759 57 1793 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 649 1389 683 1423
rect 649 1315 683 1349
rect 649 1241 683 1275
rect 649 1167 683 1201
rect 649 1093 683 1127
rect 649 1019 683 1053
rect -17 945 17 979
rect 1315 1389 1349 1423
rect 1315 1315 1349 1349
rect 1315 1241 1349 1275
rect 1315 1167 1349 1201
rect 1315 1093 1349 1127
rect 1315 1019 1349 1053
rect 649 945 683 979
rect -17 871 17 905
rect 1759 1389 1793 1423
rect 1759 1315 1793 1349
rect 1759 1241 1793 1275
rect 1759 1167 1793 1201
rect 1759 1093 1793 1127
rect 1759 1019 1793 1053
rect 1315 945 1349 979
rect 649 871 683 905
rect 1759 945 1793 979
rect 1315 871 1349 905
rect 1759 871 1793 905
<< poly >>
rect 187 1404 217 1430
rect 275 1404 305 1430
rect 363 1404 393 1430
rect 451 1404 481 1430
rect 853 1405 883 1431
rect 941 1405 971 1431
rect 1029 1405 1059 1431
rect 1117 1405 1147 1431
rect 187 973 217 1004
rect 275 973 305 1004
rect 363 973 393 1004
rect 451 973 481 1004
rect 187 957 305 973
rect 187 943 205 957
rect 195 923 205 943
rect 239 943 305 957
rect 349 957 481 973
rect 239 923 249 943
rect 195 907 249 923
rect 349 923 359 957
rect 393 943 481 957
rect 1496 1404 1526 1430
rect 1584 1404 1614 1430
rect 853 974 883 1005
rect 941 974 971 1005
rect 1029 974 1059 1005
rect 1117 974 1147 1005
rect 393 923 403 943
rect 349 907 403 923
rect 830 958 971 974
rect 830 924 840 958
rect 874 944 971 958
rect 1016 958 1147 974
rect 874 924 884 944
rect 830 908 884 924
rect 1016 924 1026 958
rect 1060 944 1147 958
rect 1496 973 1526 1004
rect 1584 973 1614 1004
rect 1060 924 1070 944
rect 1016 908 1070 924
rect 1453 957 1614 973
rect 1453 923 1463 957
rect 1497 943 1614 957
rect 1497 923 1507 943
rect 1453 907 1507 923
rect 195 433 249 449
rect 195 413 205 433
rect 168 399 205 413
rect 239 399 249 433
rect 168 383 249 399
rect 343 433 397 449
rect 343 399 353 433
rect 387 399 397 433
rect 343 383 397 399
rect 861 433 915 449
rect 861 413 871 433
rect 168 349 198 383
rect 362 349 392 383
rect 834 399 871 413
rect 905 399 915 433
rect 834 383 915 399
rect 1009 433 1063 449
rect 1009 399 1019 433
rect 1053 399 1063 433
rect 1009 383 1063 399
rect 834 349 864 383
rect 1028 349 1058 383
rect 1453 434 1507 450
rect 1453 400 1463 434
rect 1497 413 1507 434
rect 1497 400 1517 413
rect 1453 384 1517 400
rect 1487 350 1517 384
<< polycont >>
rect 205 923 239 957
rect 359 923 393 957
rect 840 924 874 958
rect 1026 924 1060 958
rect 1463 923 1497 957
rect 205 399 239 433
rect 353 399 387 433
rect 871 399 905 433
rect 1019 399 1053 433
rect 1463 400 1497 434
<< locali >>
rect -34 1497 1810 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1810 1497
rect -34 1446 1810 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 141 1366 175 1446
rect 141 1298 175 1332
rect 141 1230 175 1264
rect 141 1162 175 1196
rect 141 1093 175 1128
rect 141 1027 175 1059
rect 229 1366 263 1404
rect 229 1298 263 1332
rect 229 1230 263 1264
rect 229 1162 263 1196
rect 229 1093 263 1128
rect 317 1366 351 1446
rect 317 1298 351 1332
rect 317 1230 351 1264
rect 317 1162 351 1196
rect 317 1111 351 1128
rect 405 1366 439 1404
rect 405 1298 439 1332
rect 405 1230 439 1264
rect 405 1162 439 1196
rect 229 1057 263 1059
rect 405 1093 439 1128
rect 493 1366 527 1446
rect 493 1298 527 1332
rect 493 1230 527 1264
rect 493 1162 527 1196
rect 493 1111 527 1128
rect 632 1423 700 1446
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 405 1057 439 1059
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 229 1023 535 1057
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect 359 957 393 973
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 923
rect 205 383 239 399
rect 353 923 359 942
rect 353 907 393 923
rect 353 433 387 907
rect 353 383 387 399
rect 501 535 535 1023
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect 807 1365 841 1405
rect 807 1297 841 1331
rect 807 1229 841 1263
rect 807 1161 841 1195
rect 807 1093 841 1127
rect 895 1365 929 1446
rect 1298 1423 1366 1446
rect 895 1297 929 1331
rect 895 1229 929 1263
rect 895 1161 929 1195
rect 895 1111 929 1127
rect 983 1365 1193 1399
rect 983 1297 1017 1331
rect 983 1229 1017 1263
rect 983 1161 1017 1195
rect 983 1093 1017 1127
rect 807 1025 1017 1059
rect 1071 1297 1105 1313
rect 1071 1229 1105 1263
rect 1071 1161 1105 1195
rect 1071 1093 1105 1127
rect 1159 1297 1193 1331
rect 1159 1229 1193 1263
rect 1159 1161 1193 1195
rect 1159 1111 1193 1127
rect 1298 1389 1315 1423
rect 1349 1389 1366 1423
rect 1298 1349 1366 1389
rect 1298 1315 1315 1349
rect 1349 1315 1366 1349
rect 1298 1275 1366 1315
rect 1298 1241 1315 1275
rect 1349 1241 1366 1275
rect 1298 1201 1366 1241
rect 1298 1167 1315 1201
rect 1349 1167 1366 1201
rect 1298 1127 1366 1167
rect 1298 1093 1315 1127
rect 1349 1093 1366 1127
rect 1071 1025 1201 1059
rect 632 979 700 1019
rect 632 945 649 979
rect 683 945 700 979
rect 632 905 700 945
rect 840 958 874 974
rect 1026 958 1060 974
rect 874 924 905 942
rect 840 908 905 924
rect 632 871 649 905
rect 683 871 700 905
rect 632 822 700 871
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 122 333 156 349
rect 316 333 350 349
rect 501 348 535 501
rect 156 299 219 333
rect 253 299 316 333
rect 122 261 156 299
rect 122 193 156 227
rect 316 261 350 299
rect 122 123 156 159
rect 122 73 156 89
rect 219 208 253 224
rect -34 34 34 57
rect 219 34 253 174
rect 316 193 350 227
rect 413 314 535 348
rect 632 461 700 544
rect 632 427 649 461
rect 683 427 700 461
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect 871 535 905 908
rect 871 433 905 501
rect 871 383 905 399
rect 1019 924 1026 942
rect 1019 908 1060 924
rect 1019 433 1053 908
rect 1019 383 1053 399
rect 1167 535 1201 1025
rect 1298 1053 1366 1093
rect 1298 1019 1315 1053
rect 1349 1019 1366 1053
rect 1450 1366 1484 1446
rect 1450 1298 1484 1332
rect 1450 1230 1484 1264
rect 1450 1162 1484 1196
rect 1450 1093 1484 1128
rect 1450 1037 1484 1059
rect 1538 1366 1572 1404
rect 1538 1298 1572 1332
rect 1538 1230 1572 1264
rect 1538 1162 1572 1196
rect 1538 1093 1572 1128
rect 1298 979 1366 1019
rect 1298 945 1315 979
rect 1349 945 1366 979
rect 1298 905 1366 945
rect 1298 871 1315 905
rect 1349 871 1366 905
rect 1298 822 1366 871
rect 1463 957 1497 973
rect 413 217 447 314
rect 632 313 700 353
rect 632 279 649 313
rect 683 279 700 313
rect 413 167 447 183
rect 510 261 544 277
rect 510 193 544 227
rect 316 123 350 159
rect 510 123 544 159
rect 350 89 413 123
rect 447 89 510 123
rect 316 73 350 89
rect 510 73 544 89
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect 632 57 649 91
rect 683 57 700 91
rect 632 34 700 57
rect 788 333 822 349
rect 1167 348 1201 501
rect 788 261 822 299
rect 788 193 822 227
rect 885 314 1201 348
rect 1298 461 1366 544
rect 1298 427 1315 461
rect 1349 427 1366 461
rect 1298 387 1366 427
rect 1298 353 1315 387
rect 1349 353 1366 387
rect 1463 535 1497 923
rect 1538 933 1572 1059
rect 1626 1366 1660 1446
rect 1626 1298 1660 1332
rect 1626 1230 1660 1264
rect 1626 1162 1660 1196
rect 1626 1093 1660 1128
rect 1626 1037 1660 1059
rect 1742 1423 1810 1446
rect 1742 1389 1759 1423
rect 1793 1389 1810 1423
rect 1742 1349 1810 1389
rect 1742 1315 1759 1349
rect 1793 1315 1810 1349
rect 1742 1275 1810 1315
rect 1742 1241 1759 1275
rect 1793 1241 1810 1275
rect 1742 1201 1810 1241
rect 1742 1167 1759 1201
rect 1793 1167 1810 1201
rect 1742 1127 1810 1167
rect 1742 1093 1759 1127
rect 1793 1093 1810 1127
rect 1742 1053 1810 1093
rect 1742 1019 1759 1053
rect 1793 1019 1810 1053
rect 1742 979 1810 1019
rect 1742 945 1759 979
rect 1793 945 1810 979
rect 1538 899 1645 933
rect 1463 434 1497 501
rect 1611 433 1645 899
rect 1742 905 1810 945
rect 1742 871 1759 905
rect 1793 871 1810 905
rect 1742 822 1810 871
rect 1463 384 1497 400
rect 1537 399 1645 433
rect 1742 461 1810 544
rect 1742 427 1759 461
rect 1793 427 1810 461
rect 885 217 919 314
rect 885 167 919 183
rect 982 261 1016 278
rect 982 193 1016 227
rect 788 123 822 159
rect 1079 217 1113 314
rect 1298 313 1366 353
rect 1298 279 1315 313
rect 1349 279 1366 313
rect 1079 167 1113 183
rect 1176 261 1210 278
rect 1176 193 1210 227
rect 982 123 1016 159
rect 1176 123 1210 159
rect 822 89 885 123
rect 919 89 982 123
rect 1016 89 1079 123
rect 1113 89 1176 123
rect 788 34 822 89
rect 885 34 919 89
rect 982 34 1016 89
rect 1079 34 1113 89
rect 1176 34 1210 89
rect 1298 239 1366 279
rect 1298 205 1315 239
rect 1349 205 1366 239
rect 1298 165 1366 205
rect 1298 131 1315 165
rect 1349 131 1366 165
rect 1298 91 1366 131
rect 1298 57 1315 91
rect 1349 57 1366 91
rect 1298 34 1366 57
rect 1441 334 1475 350
rect 1441 262 1475 300
rect 1441 194 1475 228
rect 1537 218 1571 399
rect 1742 387 1810 427
rect 1742 353 1759 387
rect 1793 353 1810 387
rect 1537 168 1571 184
rect 1635 334 1669 350
rect 1635 262 1669 300
rect 1635 194 1669 228
rect 1441 124 1475 160
rect 1635 124 1669 160
rect 1475 90 1537 124
rect 1571 90 1635 124
rect 1441 34 1475 90
rect 1538 34 1572 90
rect 1635 34 1669 90
rect 1742 313 1810 353
rect 1742 279 1759 313
rect 1793 279 1810 313
rect 1742 239 1810 279
rect 1742 205 1759 239
rect 1793 205 1810 239
rect 1742 165 1810 205
rect 1742 131 1759 165
rect 1793 131 1810 165
rect 1742 91 1810 131
rect 1742 57 1759 91
rect 1793 57 1810 91
rect 1742 34 1810 57
rect -34 17 1810 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1810 17
rect -34 -34 1810 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 501 501 535 535
rect 871 501 905 535
rect 1167 501 1201 535
rect 1463 501 1497 535
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
<< metal1 >>
rect -34 1497 1810 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1810 1497
rect -34 1446 1810 1463
rect 495 535 541 541
rect 865 535 911 541
rect 1161 535 1207 541
rect 1457 535 1503 541
rect 489 501 501 535
rect 535 501 871 535
rect 905 501 917 535
rect 1155 501 1167 535
rect 1201 501 1463 535
rect 1497 501 1509 535
rect 495 495 541 501
rect 865 495 911 501
rect 1161 495 1207 501
rect 1457 495 1503 501
rect -34 17 1810 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1810 17
rect -34 -34 1810 -17
<< labels >>
rlabel metal1 1611 797 1645 831 1 Y
port 1 n
rlabel metal1 1611 723 1645 757 1 Y
port 2 n
rlabel metal1 1611 649 1645 683 1 Y
port 3 n
rlabel metal1 1611 575 1645 609 1 Y
port 4 n
rlabel metal1 1611 501 1645 535 1 Y
port 5 n
rlabel metal1 1611 427 1645 461 1 Y
port 6 n
rlabel metal1 1611 871 1645 905 1 Y
port 7 n
rlabel metal1 205 575 239 609 1 A
port 8 n
rlabel metal1 205 501 239 535 1 A
port 9 n
rlabel metal1 205 427 239 461 1 A
port 10 n
rlabel metal1 205 649 239 683 1 A
port 11 n
rlabel metal1 205 723 239 757 1 A
port 12 n
rlabel metal1 205 797 239 831 1 A
port 13 n
rlabel metal1 205 871 239 905 1 A
port 14 n
rlabel metal1 353 649 387 683 1 B
port 15 n
rlabel metal1 353 575 387 609 1 B
port 16 n
rlabel metal1 353 501 387 535 1 B
port 17 n
rlabel metal1 353 427 387 461 1 B
port 18 n
rlabel metal1 353 723 387 757 1 B
port 19 n
rlabel metal1 353 797 387 831 1 B
port 20 n
rlabel metal1 353 871 387 905 1 B
port 21 n
rlabel metal1 1019 723 1053 757 1 C
port 22 n
rlabel metal1 1019 649 1053 683 1 C
port 23 n
rlabel metal1 1019 575 1053 609 1 C
port 24 n
rlabel metal1 1019 501 1053 535 1 C
port 25 n
rlabel metal1 1019 427 1053 461 1 C
port 26 n
rlabel metal1 1019 797 1053 831 1 C
port 27 n
rlabel metal1 1019 871 1053 905 1 C
port 28 n
rlabel metal1 -34 1446 1810 1514 1 VPWR
port 29 n
rlabel metal1 -34 -34 1810 34 1 VGND
port 30 n
rlabel nwell 57 1463 91 1497 1 VPB
port 31 n
rlabel pwell 57 -17 91 17 1 VNB
port 32 n
<< end >>
