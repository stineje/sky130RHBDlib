// File: TIELO.spi.pex
// Created: Tue Oct 15 15:51:21 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_TIELO\%GND ( 1 7 19 23 35 41 48 )
c21 ( 48 0 ) capacitor c=0.0630778f //x=0.495 //y=0.365
c22 ( 41 0 ) capacitor c=0.237416f //x=1.6 //y=0
c23 ( 35 0 ) capacitor c=0.192997f //x=0.63 //y=0
c24 ( 26 0 ) capacitor c=0.00576908f //x=1.6 //y=0.445
c25 ( 23 0 ) capacitor c=0.00782031f //x=1.515 //y=0.53
c26 ( 22 0 ) capacitor c=0.00468229f //x=1.11 //y=0.445
c27 ( 19 0 ) capacitor c=0.00697428f //x=1.025 //y=0.53
c28 ( 14 0 ) capacitor c=0.00578481f //x=0.63 //y=0.445
c29 ( 7 0 ) capacitor c=0.11015f //x=1.48 //y=0
r30 (  40 41 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=1.48 //y=0 //x2=1.6 //y2=0
r31 (  38 40 ) resistor r=13.2661 //w=0.357 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=0 //x2=1.48 //y2=0
r32 (  37 38 ) resistor r=13.2661 //w=0.357 //l=0.37 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.11 //y2=0
r33 (  35 37 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=0.63 //y=0 //x2=0.74 //y2=0
r34 (  27 48 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.6 //y=0.615 //x2=1.6 //y2=0.53
r35 (  27 48 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.615 //x2=1.6 //y2=1.22
r36 (  26 48 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.6 //y=0.445 //x2=1.6 //y2=0.53
r37 (  25 41 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.6 //y=0.17 //x2=1.6 //y2=0
r38 (  25 26 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0.445
r39 (  24 48 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.195 //y=0.53 //x2=1.11 //y2=0.53
r40 (  23 48 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.53 //x2=1.6 //y2=0.53
r41 (  23 24 ) resistor r=21.9037 //w=0.187 //l=0.32 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.53 //x2=1.195 //y2=0.53
r42 (  22 48 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.11 //y=0.445 //x2=1.11 //y2=0.53
r43 (  21 38 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.11 //y=0.17 //x2=1.11 //y2=0
r44 (  21 22 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=1.11 //y=0.17 //x2=1.11 //y2=0.445
r45 (  20 48 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.715 //y=0.53 //x2=0.63 //y2=0.53
r46 (  19 48 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.025 //y=0.53 //x2=1.11 //y2=0.53
r47 (  19 20 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=1.025 //y=0.53 //x2=0.715 //y2=0.53
r48 (  15 48 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=0.63 //y=0.615 //x2=0.63 //y2=0.53
r49 (  15 48 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.615 //x2=0.63 //y2=1.22
r50 (  14 48 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=0.63 //y=0.445 //x2=0.63 //y2=0.53
r51 (  13 35 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=0.63 //y=0.17 //x2=0.63 //y2=0
r52 (  13 14 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0.445
r53 (  7 40 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=1.48 //y=0 //x2=1.48 //y2=0
r54 (  3 37 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=0.74 \
 //y=0 //x2=0.74 //y2=0
r55 (  1 7 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=1.11 //y=0 //x2=1.48 //y2=0
r56 (  1 3 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=1.11 //y=0 //x2=0.74 //y2=0
ends PM_TIELO\%GND

subckt PM_TIELO\%VDD ( 1 7 19 32 34 35 36 )
c22 ( 36 0 ) capacitor c=0.0502376f //x=1.405 //y=5.02
c23 ( 35 0 ) capacitor c=0.0446708f //x=0.535 //y=5.02
c24 ( 34 0 ) capacitor c=0.239567f //x=1.48 //y=7.4
c25 ( 32 0 ) capacitor c=0.232766f //x=0.74 //y=7.4
c26 ( 19 0 ) capacitor c=0.0288572f //x=1.465 //y=7.4
c27 ( 7 0 ) capacitor c=0.110692f //x=1.48 //y=7.4
r28 (  21 34 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.55 //y=7.23 //x2=1.55 //y2=7.4
r29 (  21 36 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.55 //y=7.23 //x2=1.55 //y2=6.405
r30 (  20 32 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.755 //y=7.4 //x2=0.67 //y2=7.4
r31 (  19 34 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.465 //y=7.4 //x2=1.55 //y2=7.4
r32 (  19 20 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.465 //y=7.4 //x2=0.755 //y2=7.4
r33 (  13 32 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=0.67 //y=7.23 //x2=0.67 //y2=7.4
r34 (  13 35 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.67 //y=7.23 //x2=0.67 //y2=6.405
r35 (  7 34 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=1.48 //y=7.4 //x2=1.48 //y2=7.4
r36 (  3 32 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=0.74 \
 //y=7.4 //x2=0.74 //y2=7.4
r37 (  1 7 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=1.11 //y=7.4 //x2=1.48 //y2=7.4
r38 (  1 3 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=1.11 //y=7.4 //x2=0.74 //y2=7.4
ends PM_TIELO\%VDD

subckt PM_TIELO\%YN ( 1 2 3 11 )
c15 ( 11 0 ) capacitor c=0.0602601f //x=0.925 //y=0.905
r16 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.59 //x2=1.11 //y2=2.96
r17 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.22 //x2=1.11 //y2=2.59
r18 (  1 11 ) resistor r=83.508 //w=0.187 //l=1.22 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.22 //x2=1.11 //y2=1
ends PM_TIELO\%YN

subckt PM_TIELO\%noxref_4 ( 1 3 5 15 16 17 18 19 20 21 25 26 27 29 35 36 38 46 )
c46 ( 46 0 ) capacitor c=0.0267071f //x=0.965 //y=5.02
c47 ( 38 0 ) capacitor c=0.0528519f //x=0.74 //y=2.08
c48 ( 36 0 ) capacitor c=0.0450427f //x=1.38 //y=1.25
c49 ( 35 0 ) capacitor c=0.0200386f //x=1.38 //y=0.905
c50 ( 29 0 ) capacitor c=0.0155406f //x=1.225 //y=1.405
c51 ( 27 0 ) capacitor c=0.0157804f //x=1.225 //y=0.75
c52 ( 26 0 ) capacitor c=0.0524209f //x=0.965 //y=4.79
c53 ( 25 0 ) capacitor c=0.0362815f //x=1.255 //y=4.79
c54 ( 21 0 ) capacitor c=0.0290017f //x=0.85 //y=1.915
c55 ( 20 0 ) capacitor c=0.0250027f //x=0.85 //y=1.56
c56 ( 19 0 ) capacitor c=0.0234316f //x=0.85 //y=1.25
c57 ( 18 0 ) capacitor c=0.0200596f //x=0.85 //y=0.905
c58 ( 17 0 ) capacitor c=0.153902f //x=1.33 //y=6.02
c59 ( 16 0 ) capacitor c=0.153904f //x=0.89 //y=6.02
c60 ( 5 0 ) capacitor c=0.0128331f //x=1.025 //y=4.7
c61 ( 3 0 ) capacitor c=0.131408f //x=0.74 //y=2.08
c62 ( 1 0 ) capacitor c=0.0038963f //x=0.74 //y=4.615
r63 (  38 39 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=0.74 //y=2.08 //x2=0.85 //y2=2.08
r64 (  36 45 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=1.25 //x2=1.34 //y2=1.405
r65 (  35 44 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.905 //x2=1.34 //y2=0.75
r66 (  35 36 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.905 //x2=1.38 //y2=1.25
r67 (  30 43 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=1.405 //x2=0.89 //y2=1.405
r68 (  29 45 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=1.405 //x2=1.34 //y2=1.405
r69 (  28 42 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=0.75 //x2=0.89 //y2=0.75
r70 (  27 44 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.75 //x2=1.34 //y2=0.75
r71 (  27 28 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.75 //x2=1.005 //y2=0.75
r72 (  25 32 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.255 //y=4.79 //x2=1.33 //y2=4.865
r73 (  25 26 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.255 //y=4.79 //x2=0.965 //y2=4.79
r74 (  22 26 ) resistor r=23.4449 //w=0.285 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=0.89 //y=4.865 //x2=0.965 //y2=4.79
r75 (  22 41 ) resistor r=25.3684 //w=0.285 //l=0.22798 //layer=ply \
 //thickness=0.18 //x=0.89 //y=4.865 //x2=0.74 //y2=4.7
r76 (  21 39 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.915 //x2=0.85 //y2=2.08
r77 (  20 43 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.56 //x2=0.89 //y2=1.405
r78 (  20 21 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.56 //x2=0.85 //y2=1.915
r79 (  19 43 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.25 //x2=0.89 //y2=1.405
r80 (  18 42 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.905 //x2=0.89 //y2=0.75
r81 (  18 19 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.905 //x2=0.85 //y2=1.25
r82 (  17 32 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.33 //y=6.02 //x2=1.33 //y2=4.865
r83 (  16 22 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=0.89 //y=6.02 //x2=0.89 //y2=4.865
r84 (  15 29 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.405 //x2=1.225 //y2=1.405
r85 (  15 30 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.405 //x2=1.005 //y2=1.405
r86 (  14 41 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=4.7 //x2=0.74 //y2=4.7
r87 (  7 46 ) resistor r=64.3422 //w=0.187 //l=0.94 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.785 //x2=1.11 //y2=5.725
r88 (  6 14 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.825 //y=4.7 //x2=0.74 //y2=4.74
r89 (  5 7 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.025 //y=4.7 //x2=1.11 //y2=4.785
r90 (  5 6 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=1.025 //y=4.7 //x2=0.825 //y2=4.7
r91 (  3 38 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=2.08 //x2=0.74 //y2=2.08
r92 (  1 14 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.74 //y=4.615 //x2=0.74 //y2=4.74
r93 (  1 3 ) resistor r=173.519 //w=0.187 //l=2.535 //layer=li //thickness=0.1 \
 //x=0.74 //y=4.615 //x2=0.74 //y2=2.08
ends PM_TIELO\%noxref_4

