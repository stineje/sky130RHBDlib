* SPICE3 file created from TIELO.ext - technology: sky130A

.subckt TIELO YN VDD GND
X0 VDD a_121_383 a_121_383 VDD pshort w=2 l=0.15 M=2
X1 YN a_121_383 GND GND nshort w=3 l=0.15
.ends
