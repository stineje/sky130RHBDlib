* SPICE3 file created from TMRDFFSNQX1.ext - technology: sky130A

.subckt TMRDFFSNQX1 Q D CLK SN VDD GND
X0 GND m1_13413_871# voter3x1_pcell_0/votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X1 GND m1_13413_871# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X2 GND m1_3606_649# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X3 voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# m1_13413_871# VDD VDD pshort w=2 l=0.15
X4 voter3x1_pcell_0/m1_1867_797# m1_3606_649# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X5 voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# m1_9639_501# VDD VDD pshort w=2 l=0.15
X6 voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# m1_3606_649# voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X7 voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# m1_13413_871# voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X8 voter3x1_pcell_0/m1_1867_797# m1_3606_649# voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X9 voter3x1_pcell_0/m1_1867_797# m1_9639_501# voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X10 voter3x1_pcell_0/m1_1867_797# m1_9639_501# voter3x1_pcell_0/votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X11 voter3x1_pcell_0/m1_1867_797# m1_9639_501# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X12 Q voter3x1_pcell_0/m1_1867_797# GND GND nshort w=3 l=0.15
X13 VDD voter3x1_pcell_0/m1_1867_797# Q VDD pshort w=2 l=0.15
X14 GND dffsnx1_pcell_1/m1_406_797# dffsnx1_pcell_1/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X15 m1_8629_501# m1_9639_501# dffsnx1_pcell_1/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X16 VDD dffsnx1_pcell_1/m1_406_797# m1_8629_501# VDD pshort w=2 l=0.15
X17 VDD m1_9639_501# m1_8629_501# VDD pshort w=2 l=0.15
X18 GND D dffsnx1_pcell_1/nand2x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X19 dffsnx1_pcell_1/m1_537_501# dffsnx1_pcell_1/m1_406_797# dffsnx1_pcell_1/nand2x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X20 VDD D dffsnx1_pcell_1/m1_537_501# VDD pshort w=2 l=0.15
X21 VDD dffsnx1_pcell_1/m1_406_797# dffsnx1_pcell_1/m1_537_501# VDD pshort w=2 l=0.15
X22 GND dffsnx1_pcell_1/m1_537_501# dffsnx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X23 dffsnx1_pcell_1/m1_406_797# dffsnx1_pcell_1/m1_1351_723# dffsnx1_pcell_1/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X24 dffsnx1_pcell_1/nand3x1_pcell_0/li_393_182# CLK dffsnx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X25 VDD dffsnx1_pcell_1/m1_537_501# dffsnx1_pcell_1/m1_406_797# VDD pshort w=2 l=0.15
X26 VDD CLK dffsnx1_pcell_1/m1_406_797# VDD pshort w=2 l=0.15
X27 VDD dffsnx1_pcell_1/m1_1351_723# dffsnx1_pcell_1/m1_406_797# VDD pshort w=2 l=0.15
X28 GND m1_8629_501# dffsnx1_pcell_1/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X29 m1_9639_501# dffsnx1_pcell_1/m1_1351_723# dffsnx1_pcell_1/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X30 dffsnx1_pcell_1/nand3x1_pcell_1/li_393_182# SN dffsnx1_pcell_1/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X31 VDD m1_8629_501# m1_9639_501# VDD pshort w=2 l=0.15
X32 VDD SN m1_9639_501# VDD pshort w=2 l=0.15
X33 VDD dffsnx1_pcell_1/m1_1351_723# m1_9639_501# VDD pshort w=2 l=0.15
X34 GND dffsnx1_pcell_1/m1_537_501# dffsnx1_pcell_1/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X35 dffsnx1_pcell_1/m1_2461_501# dffsnx1_pcell_1/m1_1351_723# dffsnx1_pcell_1/nand3x1_pcell_2/li_393_182# GND nshort w=3 l=0.15
X36 dffsnx1_pcell_1/nand3x1_pcell_2/li_393_182# SN dffsnx1_pcell_1/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X37 VDD dffsnx1_pcell_1/m1_537_501# dffsnx1_pcell_1/m1_2461_501# VDD pshort w=2 l=0.15
X38 VDD SN dffsnx1_pcell_1/m1_2461_501# VDD pshort w=2 l=0.15
X39 VDD dffsnx1_pcell_1/m1_1351_723# dffsnx1_pcell_1/m1_2461_501# VDD pshort w=2 l=0.15
X40 GND dffsnx1_pcell_1/m1_2461_501# dffsnx1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X41 dffsnx1_pcell_1/m1_1351_723# CLK dffsnx1_pcell_1/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X42 VDD dffsnx1_pcell_1/m1_2461_501# dffsnx1_pcell_1/m1_1351_723# VDD pshort w=2 l=0.15
X43 VDD CLK dffsnx1_pcell_1/m1_1351_723# VDD pshort w=2 l=0.15
X44 GND dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X45 m1_3813_797# m1_3606_649# dffsnx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X46 VDD dffsnx1_pcell_0/m1_406_797# m1_3813_797# VDD pshort w=2 l=0.15
X47 VDD m1_3606_649# m1_3813_797# VDD pshort w=2 l=0.15
X48 GND D dffsnx1_pcell_0/nand2x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X49 dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/nand2x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X50 VDD D dffsnx1_pcell_0/m1_537_501# VDD pshort w=2 l=0.15
X51 VDD dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/m1_537_501# VDD pshort w=2 l=0.15
X52 GND dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X53 dffsnx1_pcell_0/m1_406_797# dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X54 dffsnx1_pcell_0/nand3x1_pcell_0/li_393_182# CLK dffsnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X55 VDD dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/m1_406_797# VDD pshort w=2 l=0.15
X56 VDD CLK dffsnx1_pcell_0/m1_406_797# VDD pshort w=2 l=0.15
X57 VDD dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/m1_406_797# VDD pshort w=2 l=0.15
X58 GND m1_3813_797# dffsnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X59 m1_3606_649# dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X60 dffsnx1_pcell_0/nand3x1_pcell_1/li_393_182# SN dffsnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X61 VDD m1_3813_797# m1_3606_649# VDD pshort w=2 l=0.15
X62 VDD SN m1_3606_649# VDD pshort w=2 l=0.15
X63 VDD dffsnx1_pcell_0/m1_1351_723# m1_3606_649# VDD pshort w=2 l=0.15
X64 GND dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X65 dffsnx1_pcell_0/m1_2461_501# dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/nand3x1_pcell_2/li_393_182# GND nshort w=3 l=0.15
X66 dffsnx1_pcell_0/nand3x1_pcell_2/li_393_182# SN dffsnx1_pcell_0/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X67 VDD dffsnx1_pcell_0/m1_537_501# dffsnx1_pcell_0/m1_2461_501# VDD pshort w=2 l=0.15
X68 VDD SN dffsnx1_pcell_0/m1_2461_501# VDD pshort w=2 l=0.15
X69 VDD dffsnx1_pcell_0/m1_1351_723# dffsnx1_pcell_0/m1_2461_501# VDD pshort w=2 l=0.15
X70 GND dffsnx1_pcell_0/m1_2461_501# dffsnx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X71 dffsnx1_pcell_0/m1_1351_723# CLK dffsnx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X72 VDD dffsnx1_pcell_0/m1_2461_501# dffsnx1_pcell_0/m1_1351_723# VDD pshort w=2 l=0.15
X73 VDD CLK dffsnx1_pcell_0/m1_1351_723# VDD pshort w=2 l=0.15
X74 GND dffsnx1_pcell_2/m1_406_797# dffsnx1_pcell_2/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X75 m1_13561_945# m1_13413_871# dffsnx1_pcell_2/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X76 VDD dffsnx1_pcell_2/m1_406_797# m1_13561_945# VDD pshort w=2 l=0.15
X77 VDD m1_13413_871# m1_13561_945# VDD pshort w=2 l=0.15
X78 GND D dffsnx1_pcell_2/nand2x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X79 dffsnx1_pcell_2/m1_537_501# dffsnx1_pcell_2/m1_406_797# dffsnx1_pcell_2/nand2x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X80 VDD D dffsnx1_pcell_2/m1_537_501# VDD pshort w=2 l=0.15
X81 VDD dffsnx1_pcell_2/m1_406_797# dffsnx1_pcell_2/m1_537_501# VDD pshort w=2 l=0.15
X82 GND dffsnx1_pcell_2/m1_537_501# dffsnx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X83 dffsnx1_pcell_2/m1_406_797# dffsnx1_pcell_2/m1_1351_723# dffsnx1_pcell_2/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X84 dffsnx1_pcell_2/nand3x1_pcell_0/li_393_182# CLK dffsnx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X85 VDD dffsnx1_pcell_2/m1_537_501# dffsnx1_pcell_2/m1_406_797# VDD pshort w=2 l=0.15
X86 VDD CLK dffsnx1_pcell_2/m1_406_797# VDD pshort w=2 l=0.15
X87 VDD dffsnx1_pcell_2/m1_1351_723# dffsnx1_pcell_2/m1_406_797# VDD pshort w=2 l=0.15
X88 GND m1_13561_945# dffsnx1_pcell_2/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X89 m1_13413_871# dffsnx1_pcell_2/m1_1351_723# dffsnx1_pcell_2/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X90 dffsnx1_pcell_2/nand3x1_pcell_1/li_393_182# SN dffsnx1_pcell_2/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X91 VDD m1_13561_945# m1_13413_871# VDD pshort w=2 l=0.15
X92 VDD SN m1_13413_871# VDD pshort w=2 l=0.15
X93 VDD dffsnx1_pcell_2/m1_1351_723# m1_13413_871# VDD pshort w=2 l=0.15
X94 GND dffsnx1_pcell_2/m1_537_501# dffsnx1_pcell_2/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X95 dffsnx1_pcell_2/m1_2461_501# dffsnx1_pcell_2/m1_1351_723# dffsnx1_pcell_2/nand3x1_pcell_2/li_393_182# GND nshort w=3 l=0.15
X96 dffsnx1_pcell_2/nand3x1_pcell_2/li_393_182# SN dffsnx1_pcell_2/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X97 VDD dffsnx1_pcell_2/m1_537_501# dffsnx1_pcell_2/m1_2461_501# VDD pshort w=2 l=0.15
X98 VDD SN dffsnx1_pcell_2/m1_2461_501# VDD pshort w=2 l=0.15
X99 VDD dffsnx1_pcell_2/m1_1351_723# dffsnx1_pcell_2/m1_2461_501# VDD pshort w=2 l=0.15
X100 GND dffsnx1_pcell_2/m1_2461_501# dffsnx1_pcell_2/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X101 dffsnx1_pcell_2/m1_1351_723# CLK dffsnx1_pcell_2/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X102 VDD dffsnx1_pcell_2/m1_2461_501# dffsnx1_pcell_2/m1_1351_723# VDD pshort w=2 l=0.15
X103 VDD CLK dffsnx1_pcell_2/m1_1351_723# VDD pshort w=2 l=0.15
C0 VDD CLK 4.72fF
C1 m1_9639_501# VDD 2.06fF
.ends
