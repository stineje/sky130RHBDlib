magic
tech sky130A
magscale 1 2
timestamp 1648064633
<< nwell >>
rect 84 903 582 1575
rect 83 832 582 903
<< pdiffc >>
rect 141 1105 175 1139
rect 229 1105 263 1139
rect 405 1105 439 1139
<< psubdiff >>
rect 31 510 635 572
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 635 47
<< nsubdiff >>
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 635 1539
rect 31 868 635 930
<< psubdiffcont >>
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
<< poly >>
rect 168 403 198 441
rect 362 410 392 411
<< locali >>
rect 31 1539 635 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 635 1539
rect 31 1492 635 1505
rect 141 1139 175 1157
rect 141 1073 175 1105
rect 229 1139 263 1157
rect 229 1103 263 1105
rect 405 1139 439 1157
rect 405 1103 439 1105
rect 229 1069 535 1103
rect 353 954 361 988
rect 205 461 239 954
rect 353 469 387 954
rect 353 461 357 469
rect 501 376 535 1069
rect 413 342 535 376
rect 413 261 447 342
rect 219 62 253 195
rect 31 47 635 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 635 47
rect 31 0 635 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 361 1505 395 1539
rect 433 1505 467 1539
rect 505 1505 539 1539
rect 577 1505 611 1539
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 361 13 395 47
rect 433 13 467 47
rect 505 13 539 47
rect 577 13 611 47
<< metal1 >>
rect 31 1539 635 1554
rect 31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 361 1539
rect 395 1505 433 1539
rect 467 1505 505 1539
rect 539 1505 577 1539
rect 611 1505 635 1539
rect 31 1492 635 1505
rect 31 47 635 62
rect 31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 361 47
rect 395 13 433 47
rect 467 13 505 47
rect 539 13 577 47
rect 611 13 635 47
rect 31 0 635 13
use diff_ring_side  diff_ring_side_1
timestamp 1648063806
transform 1 0 0 0 1 0
box -84 0 84 1575
use nmos_bottom  nmos_bottom_0
timestamp 1648062456
transform -1 0 360 0 1 101
box 0 0 248 302
use poly_li1_contact  poly_li1_contact_0
timestamp 1648060378
transform 0 1 223 -1 0 987
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_1
timestamp 1648060378
transform 0 1 223 -1 0 445
box -32 -28 34 26
use pmos2  pmos2_0
timestamp 1648061063
transform 1 0 43 0 1 1450
box 52 -461 352 42
use poly_li1_contact  poly_li1_contact_3
timestamp 1648060378
transform 0 1 377 -1 0 987
box -32 -28 34 26
use poly_li1_contact  poly_li1_contact_2
timestamp 1648060378
transform 0 -1 369 1 0 443
box -32 -28 34 26
use pmos2  pmos2_1
timestamp 1648061063
transform 1 0 219 0 1 1450
box 52 -461 352 42
use nmos_top_trim1  nmos_top_trim1_0
timestamp 1648061897
transform -1 0 554 0 1 101
box 0 0 248 309
use diff_ring_side  diff_ring_side_0
timestamp 1648063806
transform 1 0 666 0 1 0
box -84 0 84 1575
<< end >>
