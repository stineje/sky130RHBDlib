magic
tech sky130A
magscale 1 2
timestamp 1652328683
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 131 871 165 905
rect 723 871 757 905
rect 131 797 165 831
rect 723 797 757 831
rect 131 723 165 757
rect 723 723 757 757
rect 131 649 165 683
rect 723 649 757 683
rect 131 575 165 609
rect 723 575 757 609
rect 131 501 165 535
rect 723 501 757 535
rect 131 427 165 461
rect 723 427 757 461
<< metal1 >>
rect -34 1446 922 1514
rect -34 -34 922 34
use bufx1  bufx1_0 pcells
timestamp 1652328347
transform 1 0 0 0 1 0
box -87 -34 975 1550
<< labels >>
rlabel locali 723 427 757 461 1 Y
port 1 nsew signal output
rlabel locali 723 501 757 535 1 Y
port 1 nsew signal output
rlabel locali 723 575 757 609 1 Y
port 1 nsew signal output
rlabel locali 723 649 757 683 1 Y
port 1 nsew signal output
rlabel locali 723 723 757 757 1 Y
port 1 nsew signal output
rlabel locali 723 797 757 831 1 Y
port 1 nsew signal output
rlabel locali 723 871 757 905 1 Y
port 1 nsew signal output
rlabel locali 131 427 165 461 1 A
port 2 nsew signal input
rlabel locali 131 501 165 535 1 A
port 2 nsew signal input
rlabel locali 131 575 165 609 1 A
port 2 nsew signal input
rlabel locali 131 649 165 683 1 A
port 2 nsew signal input
rlabel locali 131 723 165 757 1 A
port 2 nsew signal input
rlabel locali 131 797 165 831 1 A
port 2 nsew signal input
rlabel locali 131 871 165 905 1 A
port 2 nsew signal input
rlabel metal1 -34 1446 922 1514 1 VPWR
port 3 nsew power bidirectional abutment
rlabel metal1 -34 -34 922 34 1 VGND
port 4 nsew ground bidirectional abutment
rlabel nwell 57 1463 91 1497 1 VPB
port 5 nsew power bidirectional
rlabel pwell 57 -17 91 17 1 VNB
port 6 nsew ground bidirectional
<< properties >>
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
