magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 1 21 2203 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 751 47 781 177
rect 835 47 865 177
rect 919 47 949 177
rect 1003 47 1033 177
rect 1087 47 1117 177
rect 1171 47 1201 177
rect 1255 47 1285 177
rect 1339 47 1369 177
rect 1423 47 1453 177
rect 1507 47 1537 177
rect 1591 47 1621 177
rect 1675 47 1705 177
rect 1759 47 1789 177
rect 1843 47 1873 177
rect 1927 47 1957 177
rect 2011 47 2041 177
rect 2095 47 2125 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 751 297 781 497
rect 835 297 865 497
rect 919 297 949 497
rect 1003 297 1033 497
rect 1087 297 1117 497
rect 1171 297 1201 497
rect 1255 297 1285 497
rect 1339 297 1369 497
rect 1423 297 1453 497
rect 1507 297 1537 497
rect 1591 297 1621 497
rect 1675 297 1705 497
rect 1759 297 1789 497
rect 1843 297 1873 497
rect 1927 297 1957 497
rect 2011 297 2041 497
rect 2095 297 2125 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 97 163 177
rect 109 63 119 97
rect 153 63 163 97
rect 109 47 163 63
rect 193 165 247 177
rect 193 131 203 165
rect 237 131 247 165
rect 193 97 247 131
rect 193 63 203 97
rect 237 63 247 97
rect 193 47 247 63
rect 277 97 331 177
rect 277 63 287 97
rect 321 63 331 97
rect 277 47 331 63
rect 361 165 415 177
rect 361 131 371 165
rect 405 131 415 165
rect 361 97 415 131
rect 361 63 371 97
rect 405 63 415 97
rect 361 47 415 63
rect 445 97 499 177
rect 445 63 455 97
rect 489 63 499 97
rect 445 47 499 63
rect 529 165 583 177
rect 529 131 539 165
rect 573 131 583 165
rect 529 97 583 131
rect 529 63 539 97
rect 573 63 583 97
rect 529 47 583 63
rect 613 97 667 177
rect 613 63 623 97
rect 657 63 667 97
rect 613 47 667 63
rect 697 165 751 177
rect 697 131 707 165
rect 741 131 751 165
rect 697 97 751 131
rect 697 63 707 97
rect 741 63 751 97
rect 697 47 751 63
rect 781 97 835 177
rect 781 63 791 97
rect 825 63 835 97
rect 781 47 835 63
rect 865 165 919 177
rect 865 131 875 165
rect 909 131 919 165
rect 865 97 919 131
rect 865 63 875 97
rect 909 63 919 97
rect 865 47 919 63
rect 949 97 1003 177
rect 949 63 959 97
rect 993 63 1003 97
rect 949 47 1003 63
rect 1033 165 1087 177
rect 1033 131 1043 165
rect 1077 131 1087 165
rect 1033 97 1087 131
rect 1033 63 1043 97
rect 1077 63 1087 97
rect 1033 47 1087 63
rect 1117 97 1171 177
rect 1117 63 1127 97
rect 1161 63 1171 97
rect 1117 47 1171 63
rect 1201 165 1255 177
rect 1201 131 1211 165
rect 1245 131 1255 165
rect 1201 97 1255 131
rect 1201 63 1211 97
rect 1245 63 1255 97
rect 1201 47 1255 63
rect 1285 97 1339 177
rect 1285 63 1295 97
rect 1329 63 1339 97
rect 1285 47 1339 63
rect 1369 165 1423 177
rect 1369 131 1379 165
rect 1413 131 1423 165
rect 1369 97 1423 131
rect 1369 63 1379 97
rect 1413 63 1423 97
rect 1369 47 1423 63
rect 1453 97 1507 177
rect 1453 63 1463 97
rect 1497 63 1507 97
rect 1453 47 1507 63
rect 1537 165 1591 177
rect 1537 131 1547 165
rect 1581 131 1591 165
rect 1537 97 1591 131
rect 1537 63 1547 97
rect 1581 63 1591 97
rect 1537 47 1591 63
rect 1621 97 1675 177
rect 1621 63 1631 97
rect 1665 63 1675 97
rect 1621 47 1675 63
rect 1705 165 1759 177
rect 1705 131 1715 165
rect 1749 131 1759 165
rect 1705 97 1759 131
rect 1705 63 1715 97
rect 1749 63 1759 97
rect 1705 47 1759 63
rect 1789 97 1843 177
rect 1789 63 1799 97
rect 1833 63 1843 97
rect 1789 47 1843 63
rect 1873 165 1927 177
rect 1873 131 1883 165
rect 1917 131 1927 165
rect 1873 97 1927 131
rect 1873 63 1883 97
rect 1917 63 1927 97
rect 1873 47 1927 63
rect 1957 97 2011 177
rect 1957 63 1967 97
rect 2001 63 2011 97
rect 1957 47 2011 63
rect 2041 165 2095 177
rect 2041 131 2051 165
rect 2085 131 2095 165
rect 2041 97 2095 131
rect 2041 63 2051 97
rect 2085 63 2095 97
rect 2041 47 2095 63
rect 2125 97 2177 177
rect 2125 63 2135 97
rect 2169 63 2177 97
rect 2125 47 2177 63
<< pdiff >>
rect 27 479 79 497
rect 27 445 35 479
rect 69 445 79 479
rect 27 411 79 445
rect 27 377 35 411
rect 69 377 79 411
rect 27 343 79 377
rect 27 309 35 343
rect 69 309 79 343
rect 27 297 79 309
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 297 163 383
rect 193 479 247 497
rect 193 445 203 479
rect 237 445 247 479
rect 193 411 247 445
rect 193 377 203 411
rect 237 377 247 411
rect 193 343 247 377
rect 193 309 203 343
rect 237 309 247 343
rect 193 297 247 309
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 297 331 383
rect 361 479 415 497
rect 361 445 371 479
rect 405 445 415 479
rect 361 411 415 445
rect 361 377 371 411
rect 405 377 415 411
rect 361 343 415 377
rect 361 309 371 343
rect 405 309 415 343
rect 361 297 415 309
rect 445 485 499 497
rect 445 451 455 485
rect 489 451 499 485
rect 445 417 499 451
rect 445 383 455 417
rect 489 383 499 417
rect 445 297 499 383
rect 529 479 583 497
rect 529 445 539 479
rect 573 445 583 479
rect 529 411 583 445
rect 529 377 539 411
rect 573 377 583 411
rect 529 343 583 377
rect 529 309 539 343
rect 573 309 583 343
rect 529 297 583 309
rect 613 485 667 497
rect 613 451 623 485
rect 657 451 667 485
rect 613 417 667 451
rect 613 383 623 417
rect 657 383 667 417
rect 613 297 667 383
rect 697 479 751 497
rect 697 445 707 479
rect 741 445 751 479
rect 697 411 751 445
rect 697 377 707 411
rect 741 377 751 411
rect 697 343 751 377
rect 697 309 707 343
rect 741 309 751 343
rect 697 297 751 309
rect 781 485 835 497
rect 781 451 791 485
rect 825 451 835 485
rect 781 417 835 451
rect 781 383 791 417
rect 825 383 835 417
rect 781 297 835 383
rect 865 479 919 497
rect 865 445 875 479
rect 909 445 919 479
rect 865 411 919 445
rect 865 377 875 411
rect 909 377 919 411
rect 865 343 919 377
rect 865 309 875 343
rect 909 309 919 343
rect 865 297 919 309
rect 949 485 1003 497
rect 949 451 959 485
rect 993 451 1003 485
rect 949 417 1003 451
rect 949 383 959 417
rect 993 383 1003 417
rect 949 297 1003 383
rect 1033 479 1087 497
rect 1033 445 1043 479
rect 1077 445 1087 479
rect 1033 411 1087 445
rect 1033 377 1043 411
rect 1077 377 1087 411
rect 1033 343 1087 377
rect 1033 309 1043 343
rect 1077 309 1087 343
rect 1033 297 1087 309
rect 1117 485 1171 497
rect 1117 451 1127 485
rect 1161 451 1171 485
rect 1117 417 1171 451
rect 1117 383 1127 417
rect 1161 383 1171 417
rect 1117 297 1171 383
rect 1201 479 1255 497
rect 1201 445 1211 479
rect 1245 445 1255 479
rect 1201 411 1255 445
rect 1201 377 1211 411
rect 1245 377 1255 411
rect 1201 343 1255 377
rect 1201 309 1211 343
rect 1245 309 1255 343
rect 1201 297 1255 309
rect 1285 485 1339 497
rect 1285 451 1295 485
rect 1329 451 1339 485
rect 1285 417 1339 451
rect 1285 383 1295 417
rect 1329 383 1339 417
rect 1285 297 1339 383
rect 1369 479 1423 497
rect 1369 445 1379 479
rect 1413 445 1423 479
rect 1369 411 1423 445
rect 1369 377 1379 411
rect 1413 377 1423 411
rect 1369 343 1423 377
rect 1369 309 1379 343
rect 1413 309 1423 343
rect 1369 297 1423 309
rect 1453 485 1507 497
rect 1453 451 1463 485
rect 1497 451 1507 485
rect 1453 417 1507 451
rect 1453 383 1463 417
rect 1497 383 1507 417
rect 1453 297 1507 383
rect 1537 479 1591 497
rect 1537 445 1547 479
rect 1581 445 1591 479
rect 1537 411 1591 445
rect 1537 377 1547 411
rect 1581 377 1591 411
rect 1537 343 1591 377
rect 1537 309 1547 343
rect 1581 309 1591 343
rect 1537 297 1591 309
rect 1621 485 1675 497
rect 1621 451 1631 485
rect 1665 451 1675 485
rect 1621 417 1675 451
rect 1621 383 1631 417
rect 1665 383 1675 417
rect 1621 297 1675 383
rect 1705 479 1759 497
rect 1705 445 1715 479
rect 1749 445 1759 479
rect 1705 411 1759 445
rect 1705 377 1715 411
rect 1749 377 1759 411
rect 1705 343 1759 377
rect 1705 309 1715 343
rect 1749 309 1759 343
rect 1705 297 1759 309
rect 1789 485 1843 497
rect 1789 451 1799 485
rect 1833 451 1843 485
rect 1789 417 1843 451
rect 1789 383 1799 417
rect 1833 383 1843 417
rect 1789 297 1843 383
rect 1873 479 1927 497
rect 1873 445 1883 479
rect 1917 445 1927 479
rect 1873 411 1927 445
rect 1873 377 1883 411
rect 1917 377 1927 411
rect 1873 343 1927 377
rect 1873 309 1883 343
rect 1917 309 1927 343
rect 1873 297 1927 309
rect 1957 485 2011 497
rect 1957 451 1967 485
rect 2001 451 2011 485
rect 1957 417 2011 451
rect 1957 383 1967 417
rect 2001 383 2011 417
rect 1957 297 2011 383
rect 2041 479 2095 497
rect 2041 445 2051 479
rect 2085 445 2095 479
rect 2041 411 2095 445
rect 2041 377 2051 411
rect 2085 377 2095 411
rect 2041 343 2095 377
rect 2041 309 2051 343
rect 2085 309 2095 343
rect 2041 297 2095 309
rect 2125 485 2177 497
rect 2125 451 2135 485
rect 2169 451 2177 485
rect 2125 417 2177 451
rect 2125 383 2135 417
rect 2169 383 2177 417
rect 2125 297 2177 383
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 119 63 153 97
rect 203 131 237 165
rect 203 63 237 97
rect 287 63 321 97
rect 371 131 405 165
rect 371 63 405 97
rect 455 63 489 97
rect 539 131 573 165
rect 539 63 573 97
rect 623 63 657 97
rect 707 131 741 165
rect 707 63 741 97
rect 791 63 825 97
rect 875 131 909 165
rect 875 63 909 97
rect 959 63 993 97
rect 1043 131 1077 165
rect 1043 63 1077 97
rect 1127 63 1161 97
rect 1211 131 1245 165
rect 1211 63 1245 97
rect 1295 63 1329 97
rect 1379 131 1413 165
rect 1379 63 1413 97
rect 1463 63 1497 97
rect 1547 131 1581 165
rect 1547 63 1581 97
rect 1631 63 1665 97
rect 1715 131 1749 165
rect 1715 63 1749 97
rect 1799 63 1833 97
rect 1883 131 1917 165
rect 1883 63 1917 97
rect 1967 63 2001 97
rect 2051 131 2085 165
rect 2051 63 2085 97
rect 2135 63 2169 97
<< pdiffc >>
rect 35 445 69 479
rect 35 377 69 411
rect 35 309 69 343
rect 119 451 153 485
rect 119 383 153 417
rect 203 445 237 479
rect 203 377 237 411
rect 203 309 237 343
rect 287 451 321 485
rect 287 383 321 417
rect 371 445 405 479
rect 371 377 405 411
rect 371 309 405 343
rect 455 451 489 485
rect 455 383 489 417
rect 539 445 573 479
rect 539 377 573 411
rect 539 309 573 343
rect 623 451 657 485
rect 623 383 657 417
rect 707 445 741 479
rect 707 377 741 411
rect 707 309 741 343
rect 791 451 825 485
rect 791 383 825 417
rect 875 445 909 479
rect 875 377 909 411
rect 875 309 909 343
rect 959 451 993 485
rect 959 383 993 417
rect 1043 445 1077 479
rect 1043 377 1077 411
rect 1043 309 1077 343
rect 1127 451 1161 485
rect 1127 383 1161 417
rect 1211 445 1245 479
rect 1211 377 1245 411
rect 1211 309 1245 343
rect 1295 451 1329 485
rect 1295 383 1329 417
rect 1379 445 1413 479
rect 1379 377 1413 411
rect 1379 309 1413 343
rect 1463 451 1497 485
rect 1463 383 1497 417
rect 1547 445 1581 479
rect 1547 377 1581 411
rect 1547 309 1581 343
rect 1631 451 1665 485
rect 1631 383 1665 417
rect 1715 445 1749 479
rect 1715 377 1749 411
rect 1715 309 1749 343
rect 1799 451 1833 485
rect 1799 383 1833 417
rect 1883 445 1917 479
rect 1883 377 1917 411
rect 1883 309 1917 343
rect 1967 451 2001 485
rect 1967 383 2001 417
rect 2051 445 2085 479
rect 2051 377 2085 411
rect 2051 309 2085 343
rect 2135 451 2169 485
rect 2135 383 2169 417
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 751 497 781 523
rect 835 497 865 523
rect 919 497 949 523
rect 1003 497 1033 523
rect 1087 497 1117 523
rect 1171 497 1201 523
rect 1255 497 1285 523
rect 1339 497 1369 523
rect 1423 497 1453 523
rect 1507 497 1537 523
rect 1591 497 1621 523
rect 1675 497 1705 523
rect 1759 497 1789 523
rect 1843 497 1873 523
rect 1927 497 1957 523
rect 2011 497 2041 523
rect 2095 497 2125 523
rect 79 259 109 297
rect 163 259 193 297
rect 247 259 277 297
rect 79 249 277 259
rect 79 215 119 249
rect 153 215 187 249
rect 221 215 277 249
rect 79 205 277 215
rect 79 177 109 205
rect 163 177 193 205
rect 247 177 277 205
rect 331 259 361 297
rect 415 259 445 297
rect 499 259 529 297
rect 583 259 613 297
rect 667 259 697 297
rect 751 259 781 297
rect 331 249 781 259
rect 331 215 355 249
rect 389 215 423 249
rect 457 215 491 249
rect 525 215 559 249
rect 593 215 627 249
rect 661 215 695 249
rect 729 215 781 249
rect 331 205 781 215
rect 331 177 361 205
rect 415 177 445 205
rect 499 177 529 205
rect 583 177 613 205
rect 667 177 697 205
rect 751 177 781 205
rect 835 259 865 297
rect 919 259 949 297
rect 1003 259 1033 297
rect 1087 259 1117 297
rect 1171 259 1201 297
rect 1255 259 1285 297
rect 1339 259 1369 297
rect 1423 259 1453 297
rect 1507 259 1537 297
rect 1591 259 1621 297
rect 1675 259 1705 297
rect 1759 259 1789 297
rect 1843 259 1873 297
rect 1927 259 1957 297
rect 2011 259 2041 297
rect 2095 259 2125 297
rect 835 249 2125 259
rect 835 215 855 249
rect 889 215 923 249
rect 957 215 991 249
rect 1025 215 1059 249
rect 1093 215 1127 249
rect 1161 215 1195 249
rect 1229 215 1263 249
rect 1297 215 1331 249
rect 1365 215 1399 249
rect 1433 215 1467 249
rect 1501 215 1535 249
rect 1569 215 1603 249
rect 1637 215 1671 249
rect 1705 215 1739 249
rect 1773 215 1807 249
rect 1841 215 1875 249
rect 1909 215 1943 249
rect 1977 215 2011 249
rect 2045 215 2125 249
rect 835 205 2125 215
rect 835 177 865 205
rect 919 177 949 205
rect 1003 177 1033 205
rect 1087 177 1117 205
rect 1171 177 1201 205
rect 1255 177 1285 205
rect 1339 177 1369 205
rect 1423 177 1453 205
rect 1507 177 1537 205
rect 1591 177 1621 205
rect 1675 177 1705 205
rect 1759 177 1789 205
rect 1843 177 1873 205
rect 1927 177 1957 205
rect 2011 177 2041 205
rect 2095 177 2125 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 751 21 781 47
rect 835 21 865 47
rect 919 21 949 47
rect 1003 21 1033 47
rect 1087 21 1117 47
rect 1171 21 1201 47
rect 1255 21 1285 47
rect 1339 21 1369 47
rect 1423 21 1453 47
rect 1507 21 1537 47
rect 1591 21 1621 47
rect 1675 21 1705 47
rect 1759 21 1789 47
rect 1843 21 1873 47
rect 1927 21 1957 47
rect 2011 21 2041 47
rect 2095 21 2125 47
<< polycont >>
rect 119 215 153 249
rect 187 215 221 249
rect 355 215 389 249
rect 423 215 457 249
rect 491 215 525 249
rect 559 215 593 249
rect 627 215 661 249
rect 695 215 729 249
rect 855 215 889 249
rect 923 215 957 249
rect 991 215 1025 249
rect 1059 215 1093 249
rect 1127 215 1161 249
rect 1195 215 1229 249
rect 1263 215 1297 249
rect 1331 215 1365 249
rect 1399 215 1433 249
rect 1467 215 1501 249
rect 1535 215 1569 249
rect 1603 215 1637 249
rect 1671 215 1705 249
rect 1739 215 1773 249
rect 1807 215 1841 249
rect 1875 215 1909 249
rect 1943 215 1977 249
rect 2011 215 2045 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 19 479 85 493
rect 19 445 35 479
rect 69 445 85 479
rect 19 411 85 445
rect 19 377 35 411
rect 69 377 85 411
rect 19 343 85 377
rect 119 485 153 527
rect 119 417 153 451
rect 119 357 153 383
rect 187 479 253 493
rect 187 445 203 479
rect 237 445 253 479
rect 187 411 253 445
rect 187 377 203 411
rect 237 377 253 411
rect 19 309 35 343
rect 69 323 85 343
rect 187 343 253 377
rect 287 485 321 527
rect 287 417 321 451
rect 287 357 321 383
rect 355 479 421 493
rect 355 445 371 479
rect 405 445 421 479
rect 355 411 421 445
rect 355 377 371 411
rect 405 377 421 411
rect 187 323 203 343
rect 69 309 203 323
rect 237 323 253 343
rect 355 343 421 377
rect 455 485 489 527
rect 455 417 489 451
rect 455 367 489 383
rect 523 479 589 493
rect 523 445 539 479
rect 573 445 589 479
rect 523 411 589 445
rect 523 377 539 411
rect 573 377 589 411
rect 237 309 321 323
rect 19 289 321 309
rect 355 309 371 343
rect 405 323 421 343
rect 523 343 589 377
rect 623 485 657 527
rect 623 417 657 451
rect 623 367 657 383
rect 691 479 757 493
rect 691 445 707 479
rect 741 445 757 479
rect 691 411 757 445
rect 691 377 707 411
rect 741 377 757 411
rect 523 323 539 343
rect 405 309 539 323
rect 573 323 589 343
rect 691 343 757 377
rect 791 485 825 527
rect 791 417 825 451
rect 791 367 825 383
rect 859 479 925 493
rect 859 445 875 479
rect 909 445 925 479
rect 859 411 925 445
rect 859 377 875 411
rect 909 377 925 411
rect 691 323 707 343
rect 573 309 707 323
rect 741 323 757 343
rect 859 343 925 377
rect 959 485 993 527
rect 959 417 993 451
rect 959 367 993 383
rect 1027 479 1093 493
rect 1027 445 1043 479
rect 1077 445 1093 479
rect 1027 411 1093 445
rect 1027 377 1043 411
rect 1077 377 1093 411
rect 741 309 825 323
rect 355 289 825 309
rect 859 309 875 343
rect 909 323 925 343
rect 1027 343 1093 377
rect 1127 485 1161 527
rect 1127 417 1161 451
rect 1127 367 1161 383
rect 1195 479 1261 493
rect 1195 445 1211 479
rect 1245 445 1261 479
rect 1195 411 1261 445
rect 1195 377 1211 411
rect 1245 377 1261 411
rect 1027 323 1043 343
rect 909 309 1043 323
rect 1077 323 1093 343
rect 1195 343 1261 377
rect 1295 485 1329 527
rect 1295 417 1329 451
rect 1295 367 1329 383
rect 1363 479 1429 493
rect 1363 445 1379 479
rect 1413 445 1429 479
rect 1363 411 1429 445
rect 1363 377 1379 411
rect 1413 377 1429 411
rect 1195 323 1211 343
rect 1077 309 1211 323
rect 1245 323 1261 343
rect 1363 343 1429 377
rect 1463 485 1497 527
rect 1463 417 1497 451
rect 1463 367 1497 383
rect 1531 479 1597 493
rect 1531 445 1547 479
rect 1581 445 1597 479
rect 1531 411 1597 445
rect 1531 377 1547 411
rect 1581 377 1597 411
rect 1363 323 1379 343
rect 1245 309 1379 323
rect 1413 323 1429 343
rect 1531 343 1597 377
rect 1631 485 1665 527
rect 1631 417 1665 451
rect 1631 367 1665 383
rect 1699 479 1765 493
rect 1699 445 1715 479
rect 1749 445 1765 479
rect 1699 411 1765 445
rect 1699 377 1715 411
rect 1749 377 1765 411
rect 1531 323 1547 343
rect 1413 309 1547 323
rect 1581 323 1597 343
rect 1699 343 1765 377
rect 1799 485 1833 527
rect 1799 417 1833 451
rect 1799 367 1833 383
rect 1867 479 1933 493
rect 1867 445 1883 479
rect 1917 445 1933 479
rect 1867 411 1933 445
rect 1867 377 1883 411
rect 1917 377 1933 411
rect 1699 323 1715 343
rect 1581 309 1715 323
rect 1749 323 1765 343
rect 1867 343 1933 377
rect 1967 485 2001 527
rect 1967 417 2001 451
rect 1967 367 2001 383
rect 2035 479 2101 493
rect 2035 445 2051 479
rect 2085 445 2101 479
rect 2035 411 2101 445
rect 2035 377 2051 411
rect 2085 377 2101 411
rect 1867 323 1883 343
rect 1749 309 1883 323
rect 1917 323 1933 343
rect 2035 343 2101 377
rect 2135 485 2169 527
rect 2135 417 2169 451
rect 2135 367 2169 383
rect 2035 323 2051 343
rect 1917 309 2051 323
rect 2085 323 2101 343
rect 2085 309 2191 323
rect 859 289 2191 309
rect 287 255 321 289
rect 790 255 825 289
rect 18 249 253 255
rect 18 215 119 249
rect 153 215 187 249
rect 221 215 253 249
rect 287 249 749 255
rect 287 215 355 249
rect 389 215 423 249
rect 457 215 491 249
rect 525 215 559 249
rect 593 215 627 249
rect 661 215 695 249
rect 729 215 749 249
rect 790 249 2102 255
rect 790 215 855 249
rect 889 215 923 249
rect 957 215 991 249
rect 1025 215 1059 249
rect 1093 215 1127 249
rect 1161 215 1195 249
rect 1229 215 1263 249
rect 1297 215 1331 249
rect 1365 215 1399 249
rect 1433 215 1467 249
rect 1501 215 1535 249
rect 1569 215 1603 249
rect 1637 215 1671 249
rect 1705 215 1739 249
rect 1773 215 1807 249
rect 1841 215 1875 249
rect 1909 215 1943 249
rect 1977 215 2011 249
rect 2045 215 2102 249
rect 287 181 321 215
rect 790 181 825 215
rect 2136 181 2191 289
rect 19 165 321 181
rect 19 131 35 165
rect 69 147 203 165
rect 69 131 85 147
rect 19 97 85 131
rect 187 131 203 147
rect 237 147 321 165
rect 355 165 825 181
rect 237 131 253 147
rect 19 63 35 97
rect 69 63 85 97
rect 19 52 85 63
rect 119 97 153 113
rect 119 17 153 63
rect 187 97 253 131
rect 355 131 371 165
rect 405 147 539 165
rect 405 131 421 147
rect 187 63 203 97
rect 237 63 253 97
rect 187 52 253 63
rect 287 97 321 113
rect 287 17 321 63
rect 355 97 421 131
rect 523 131 539 147
rect 573 147 707 165
rect 573 131 589 147
rect 355 63 371 97
rect 405 63 421 97
rect 355 52 421 63
rect 455 97 489 113
rect 455 17 489 63
rect 523 97 589 131
rect 691 131 707 147
rect 741 147 825 165
rect 859 165 2191 181
rect 741 131 757 147
rect 523 63 539 97
rect 573 63 589 97
rect 523 52 589 63
rect 623 97 657 113
rect 623 17 657 63
rect 691 97 757 131
rect 859 131 875 165
rect 909 147 1043 165
rect 909 131 925 147
rect 691 63 707 97
rect 741 63 757 97
rect 691 52 757 63
rect 791 97 825 113
rect 791 17 825 63
rect 859 97 925 131
rect 1027 131 1043 147
rect 1077 147 1211 165
rect 1077 131 1093 147
rect 859 63 875 97
rect 909 63 925 97
rect 859 52 925 63
rect 959 97 993 113
rect 859 51 909 52
rect 959 17 993 63
rect 1027 97 1093 131
rect 1195 131 1211 147
rect 1245 147 1379 165
rect 1245 131 1261 147
rect 1027 63 1043 97
rect 1077 63 1093 97
rect 1027 52 1093 63
rect 1127 97 1161 113
rect 1043 51 1077 52
rect 1127 17 1161 63
rect 1195 97 1261 131
rect 1363 131 1379 147
rect 1413 147 1547 165
rect 1413 131 1429 147
rect 1195 63 1211 97
rect 1245 63 1261 97
rect 1195 52 1261 63
rect 1295 97 1329 113
rect 1211 51 1245 52
rect 1295 17 1329 63
rect 1363 97 1429 131
rect 1531 131 1547 147
rect 1581 147 1715 165
rect 1581 131 1597 147
rect 1363 63 1379 97
rect 1413 63 1429 97
rect 1363 52 1429 63
rect 1463 97 1497 113
rect 1463 17 1497 63
rect 1531 97 1597 131
rect 1699 131 1715 147
rect 1749 147 1883 165
rect 1749 131 1765 147
rect 1531 63 1547 97
rect 1581 63 1597 97
rect 1531 52 1597 63
rect 1631 97 1665 113
rect 1631 17 1665 63
rect 1699 97 1765 131
rect 1867 131 1883 147
rect 1917 147 2051 165
rect 1917 131 1933 147
rect 1699 63 1715 97
rect 1749 63 1765 97
rect 1699 52 1765 63
rect 1799 97 1833 113
rect 1799 17 1833 63
rect 1867 97 1933 131
rect 2035 131 2051 147
rect 2085 147 2191 165
rect 2085 131 2101 147
rect 1867 63 1883 97
rect 1917 63 1933 97
rect 1867 52 1933 63
rect 1967 97 2001 113
rect 1967 17 2001 63
rect 2035 97 2101 131
rect 2035 63 2051 97
rect 2085 63 2101 97
rect 2035 52 2101 63
rect 2135 97 2169 113
rect 2135 17 2169 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 2146 221 2180 255 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel locali s 2146 289 2180 323 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 bufinv_16
rlabel metal1 s 0 -48 2208 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2208 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 2208 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 3223662
string GDS_START 3206836
string path 0.000 0.000 55.200 0.000 
<< end >>
