* SPICE3 file created from DFFSNRNQNX1.ext - technology: sky130A

.subckt DFFSNRNQNX1 QN D CLK SN RN VDD GND
X0  D nand3x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X1 m1_867_576# m1_716_723# nand3x1_pcell_0/li_393_182#  nshort w=3 l=0.15
X2 nand3x1_pcell_0/li_393_182# RN nand3x1_pcell_0/nmos_bottom_0/a_0_0#  nshort w=3 l=0.15
X3 VDD D m1_867_576# VDD pshort w=2 l=0.15
X4 VDD RN m1_867_576# VDD pshort w=2 l=0.15
X5 VDD m1_716_723# m1_867_576# VDD pshort w=2 l=0.15
X6 GND m1_867_576# nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X7 m1_716_723# m1_1680_797# nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X8 nand3x1_pcell_1/li_393_182# CLK nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X9 VDD m1_867_576# m1_716_723# VDD pshort w=2 l=0.15
X10 VDD CLK m1_716_723# VDD pshort w=2 l=0.15
X11 VDD m1_1680_797# m1_716_723# VDD pshort w=2 l=0.15
X12 li1_M1_contact_9/VSUBS m1_867_576# nand3x1_pcell_2/nmos_bottom_0/a_0_0# li1_M1_contact_9/VSUBS nshort w=3 l=0.15
X13 m1_2791_575# m1_1680_797# nand3x1_pcell_2/li_393_182# li1_M1_contact_9/VSUBS nshort w=3 l=0.15
X14 nand3x1_pcell_2/li_393_182# SN nand3x1_pcell_2/nmos_bottom_0/a_0_0# li1_M1_contact_9/VSUBS nshort w=3 l=0.15
X15 VDD m1_867_576# m1_2791_575# VDD pshort w=2 l=0.15
X16 VDD SN m1_2791_575# VDD pshort w=2 l=0.15
X17 VDD m1_1680_797# m1_2791_575# VDD pshort w=2 l=0.15
X18 li1_M1_contact_9/VSUBS m1_2791_575# nand3x1_pcell_3/nmos_bottom_0/a_0_0# li1_M1_contact_9/VSUBS nshort w=3 l=0.15
X19 m1_1680_797# RN nand3x1_pcell_3/li_393_182# li1_M1_contact_9/VSUBS nshort w=3 l=0.15
X20 nand3x1_pcell_3/li_393_182# CLK nand3x1_pcell_3/nmos_bottom_0/a_0_0# li1_M1_contact_9/VSUBS nshort w=3 l=0.15
X21 VDD m1_2791_575# m1_1680_797# VDD pshort w=2 l=0.15
X22 VDD CLK m1_1680_797# VDD pshort w=2 l=0.15
X23 VDD RN m1_1680_797# VDD pshort w=2 l=0.15
X24 �7h� m1_716_723# nand3x1_pcell_4/nmos_bottom_0/a_0_0# �7h� nshort w=3 l=0.15
X25 QN m1_4567_723# nand3x1_pcell_4/li_393_182# �7h� nshort w=3 l=0.15
X26 nand3x1_pcell_4/li_393_182# RN nand3x1_pcell_4/nmos_bottom_0/a_0_0# �7h� nshort w=3 l=0.15
X27 VDD m1_716_723# QN VDD pshort w=2 l=0.15
X28 VDD RN QN VDD pshort w=2 l=0.15
X29 VDD m1_4567_723# QN VDD pshort w=2 l=0.15
X30 nand3x1_pcell_5/pmos2_2/VSUBS QN nand3x1_pcell_5/nmos_bottom_0/a_0_0# nand3x1_pcell_5/pmos2_2/VSUBS nshort w=3 l=0.15
X31 m1_4567_723# m1_1680_797# nand3x1_pcell_5/li_393_182# nand3x1_pcell_5/pmos2_2/VSUBS nshort w=3 l=0.15
X32 nand3x1_pcell_5/li_393_182# SN nand3x1_pcell_5/nmos_bottom_0/a_0_0# nand3x1_pcell_5/pmos2_2/VSUBS nshort w=3 l=0.15
X33 VDD QN m1_4567_723# VDD pshort w=2 l=0.15
X34 VDD SN m1_4567_723# VDD pshort w=2 l=0.15
X35 VDD m1_1680_797# m1_4567_723# VDD pshort w=2 l=0.15
C0 m1_1680_797# VDD 2.43fF
C1 VDD nand3x1_pcell_5/pmos2_2/VSUBS 6.34fF
.ends
