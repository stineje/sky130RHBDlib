* SPICE3 file created from AOA4X1.ext - technology: sky130A

.subckt AOA4X1 Y A B C D VDD GND
M1000 a_864_209.t1 C.t0 a_797_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 GND A.t1 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=3.4356p pd=24.18u as=0p ps=0u
M1002 GND a_864_209.t4 a_1444_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD.t2 a_217_1050.t5 a_797_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1549_1050.t1 D.t0 VDD.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VDD.t5 A.t0 a_217_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y.t1 a_1549_1050.t5 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VDD.t11 B.t0 a_217_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VDD.t8 a_864_209.t5 a_1549_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_1549_1050.t7 GND.t4 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1010 VDD.t3 a_1549_1050.t6 Y.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_217_1050.t2 A.t2 VDD.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_797_1051.t1 C.t1 a_864_209.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_797_1051.t3 a_217_1050.t7 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t4 D.t2 a_1549_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_217_1050.t1 B.t2 VDD.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1549_1050.t3 a_864_209.t6 VDD.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 B VDD 0.07fF
C1 D VDD 0.07fF
C2 Y VDD 0.78fF
C3 C VDD 0.07fF
C4 B A 0.27fF
C5 VDD A 0.08fF
R0 C.n0 C.t1 470.752
R1 C.n0 C.t0 384.527
R2 C.n1 C.t2 241.172
R3 C.n1 C.n0 110.173
R4 C.n2 C.n1 76
R5 C.n2 C 0.046
R6 a_797_1051.n0 a_797_1051.t1 101.66
R7 a_797_1051.n0 a_797_1051.t2 101.66
R8 a_797_1051.t0 a_797_1051.n0 14.294
R9 a_797_1051.n0 a_797_1051.t3 14.282
R10 a_864_209.n0 a_864_209.t5 480.392
R11 a_864_209.n0 a_864_209.t6 403.272
R12 a_864_209.n10 a_864_209.n9 244.994
R13 a_864_209.n1 a_864_209.t4 203.821
R14 a_864_209.n1 a_864_209.n0 178.106
R15 a_864_209.n9 a_864_209.n1 153.315
R16 a_864_209.n8 a_864_209.n7 133.539
R17 a_864_209.n9 a_864_209.n8 82.528
R18 a_864_209.n4 a_864_209.n2 80.526
R19 a_864_209.n8 a_864_209.n4 48.405
R20 a_864_209.n4 a_864_209.n3 30
R21 a_864_209.n7 a_864_209.n6 22.578
R22 a_864_209.n10 a_864_209.t0 14.282
R23 a_864_209.t1 a_864_209.n10 14.282
R24 a_864_209.n7 a_864_209.n5 8.58
R25 a_217_1050.n4 a_217_1050.t7 486.819
R26 a_217_1050.n4 a_217_1050.t5 384.527
R27 a_217_1050.n6 a_217_1050.n3 232.158
R28 a_217_1050.n5 a_217_1050.t6 197.395
R29 a_217_1050.n5 a_217_1050.n4 186.206
R30 a_217_1050.n6 a_217_1050.n5 153.315
R31 a_217_1050.n8 a_217_1050.n6 130.933
R32 a_217_1050.n3 a_217_1050.n2 76.002
R33 a_217_1050.n8 a_217_1050.n7 30
R34 a_217_1050.n9 a_217_1050.n0 24.383
R35 a_217_1050.n9 a_217_1050.n8 23.684
R36 a_217_1050.n1 a_217_1050.t4 14.282
R37 a_217_1050.n1 a_217_1050.t1 14.282
R38 a_217_1050.n2 a_217_1050.t0 14.282
R39 a_217_1050.n2 a_217_1050.t2 14.282
R40 a_217_1050.n3 a_217_1050.n1 12.85
R41 VDD.n129 VDD.n127 144.705
R42 VDD.n214 VDD.n212 144.705
R43 VDD.n68 VDD.n66 144.705
R44 VDD.n26 VDD.n25 77.792
R45 VDD.n35 VDD.n34 77.792
R46 VDD.n29 VDD.n23 76.145
R47 VDD.n29 VDD.n28 76
R48 VDD.n33 VDD.n32 76
R49 VDD.n39 VDD.n38 76
R50 VDD.n43 VDD.n42 76
R51 VDD.n70 VDD.n69 76
R52 VDD.n75 VDD.n74 76
R53 VDD.n80 VDD.n79 76
R54 VDD.n86 VDD.n85 76
R55 VDD.n91 VDD.n90 76
R56 VDD.n96 VDD.n95 76
R57 VDD.n101 VDD.n100 76
R58 VDD.n105 VDD.n104 76
R59 VDD.n131 VDD.n130 76
R60 VDD.n244 VDD.n243 76
R61 VDD.n240 VDD.n239 76
R62 VDD.n236 VDD.n235 76
R63 VDD.n232 VDD.n231 76
R64 VDD.n227 VDD.n226 76
R65 VDD.n220 VDD.n219 76
R66 VDD.n216 VDD.n215 76
R67 VDD.n189 VDD.n188 76
R68 VDD.n185 VDD.n184 76
R69 VDD.n180 VDD.n179 76
R70 VDD.n175 VDD.n174 76
R71 VDD.n169 VDD.n168 76
R72 VDD.n164 VDD.n163 76
R73 VDD.n159 VDD.n158 76
R74 VDD.n154 VDD.n153 76
R75 VDD.n155 VDD.t10 55.106
R76 VDD.n97 VDD.t7 55.106
R77 VDD.n37 VDD.t0 55.106
R78 VDD.n24 VDD.t3 55.106
R79 VDD.n181 VDD.t11 55.106
R80 VDD.n71 VDD.t4 55.106
R81 VDD.n222 VDD.n221 41.183
R82 VDD.n171 VDD.n170 40.824
R83 VDD.n82 VDD.n81 40.824
R84 VDD.n110 VDD.n109 36.774
R85 VDD.n48 VDD.n47 36.774
R86 VDD.n205 VDD.n204 36.774
R87 VDD.n77 VDD.n76 36.608
R88 VDD.n177 VDD.n176 36.608
R89 VDD.n93 VDD.n92 32.032
R90 VDD.n224 VDD.n223 32.032
R91 VDD.n161 VDD.n160 32.032
R92 VDD.n153 VDD.n150 21.841
R93 VDD.n23 VDD.n20 21.841
R94 VDD.n170 VDD.t6 14.282
R95 VDD.n170 VDD.t5 14.282
R96 VDD.n221 VDD.t1 14.282
R97 VDD.n221 VDD.t2 14.282
R98 VDD.n81 VDD.t9 14.282
R99 VDD.n81 VDD.t8 14.282
R100 VDD.n150 VDD.n133 14.167
R101 VDD.n133 VDD.n132 14.167
R102 VDD.n125 VDD.n107 14.167
R103 VDD.n107 VDD.n106 14.167
R104 VDD.n64 VDD.n45 14.167
R105 VDD.n45 VDD.n44 14.167
R106 VDD.n210 VDD.n191 14.167
R107 VDD.n191 VDD.n190 14.167
R108 VDD.n20 VDD.n19 14.167
R109 VDD.n19 VDD.n17 14.167
R110 VDD.n69 VDD.n65 14.167
R111 VDD.n130 VDD.n126 14.167
R112 VDD.n215 VDD.n211 14.167
R113 VDD.n23 VDD.n22 13.653
R114 VDD.n22 VDD.n21 13.653
R115 VDD.n28 VDD.n27 13.653
R116 VDD.n27 VDD.n26 13.653
R117 VDD.n32 VDD.n31 13.653
R118 VDD.n31 VDD.n30 13.653
R119 VDD.n38 VDD.n36 13.653
R120 VDD.n36 VDD.n35 13.653
R121 VDD.n42 VDD.n41 13.653
R122 VDD.n41 VDD.n40 13.653
R123 VDD.n69 VDD.n68 13.653
R124 VDD.n68 VDD.n67 13.653
R125 VDD.n74 VDD.n73 13.653
R126 VDD.n73 VDD.n72 13.653
R127 VDD.n79 VDD.n78 13.653
R128 VDD.n78 VDD.n77 13.653
R129 VDD.n85 VDD.n84 13.653
R130 VDD.n84 VDD.n83 13.653
R131 VDD.n90 VDD.n89 13.653
R132 VDD.n89 VDD.n88 13.653
R133 VDD.n95 VDD.n94 13.653
R134 VDD.n94 VDD.n93 13.653
R135 VDD.n100 VDD.n99 13.653
R136 VDD.n99 VDD.n98 13.653
R137 VDD.n104 VDD.n103 13.653
R138 VDD.n103 VDD.n102 13.653
R139 VDD.n130 VDD.n129 13.653
R140 VDD.n129 VDD.n128 13.653
R141 VDD.n243 VDD.n242 13.653
R142 VDD.n242 VDD.n241 13.653
R143 VDD.n239 VDD.n238 13.653
R144 VDD.n238 VDD.n237 13.653
R145 VDD.n235 VDD.n234 13.653
R146 VDD.n234 VDD.n233 13.653
R147 VDD.n231 VDD.n230 13.653
R148 VDD.n230 VDD.n229 13.653
R149 VDD.n226 VDD.n225 13.653
R150 VDD.n225 VDD.n224 13.653
R151 VDD.n219 VDD.n218 13.653
R152 VDD.n218 VDD.n217 13.653
R153 VDD.n215 VDD.n214 13.653
R154 VDD.n214 VDD.n213 13.653
R155 VDD.n188 VDD.n187 13.653
R156 VDD.n187 VDD.n186 13.653
R157 VDD.n184 VDD.n183 13.653
R158 VDD.n183 VDD.n182 13.653
R159 VDD.n179 VDD.n178 13.653
R160 VDD.n178 VDD.n177 13.653
R161 VDD.n174 VDD.n173 13.653
R162 VDD.n173 VDD.n172 13.653
R163 VDD.n168 VDD.n167 13.653
R164 VDD.n167 VDD.n166 13.653
R165 VDD.n163 VDD.n162 13.653
R166 VDD.n162 VDD.n161 13.653
R167 VDD.n158 VDD.n157 13.653
R168 VDD.n157 VDD.n156 13.653
R169 VDD.n153 VDD.n152 13.653
R170 VDD.n152 VDD.n151 13.653
R171 VDD.n4 VDD.n2 12.915
R172 VDD.n4 VDD.n3 12.66
R173 VDD.n13 VDD.n12 12.343
R174 VDD.n10 VDD.n9 12.343
R175 VDD.n7 VDD.n6 12.343
R176 VDD.n85 VDD.n82 8.658
R177 VDD.n174 VDD.n171 8.658
R178 VDD.n126 VDD.n125 7.674
R179 VDD.n65 VDD.n64 7.674
R180 VDD.n211 VDD.n210 7.674
R181 VDD.n59 VDD.n58 7.5
R182 VDD.n53 VDD.n52 7.5
R183 VDD.n55 VDD.n54 7.5
R184 VDD.n50 VDD.n49 7.5
R185 VDD.n64 VDD.n63 7.5
R186 VDD.n120 VDD.n119 7.5
R187 VDD.n114 VDD.n113 7.5
R188 VDD.n116 VDD.n115 7.5
R189 VDD.n122 VDD.n112 7.5
R190 VDD.n122 VDD.n110 7.5
R191 VDD.n125 VDD.n124 7.5
R192 VDD.n195 VDD.n194 7.5
R193 VDD.n198 VDD.n197 7.5
R194 VDD.n200 VDD.n199 7.5
R195 VDD.n203 VDD.n202 7.5
R196 VDD.n210 VDD.n209 7.5
R197 VDD.n145 VDD.n144 7.5
R198 VDD.n139 VDD.n138 7.5
R199 VDD.n141 VDD.n140 7.5
R200 VDD.n147 VDD.n137 7.5
R201 VDD.n147 VDD.n135 7.5
R202 VDD.n150 VDD.n149 7.5
R203 VDD.n20 VDD.n16 7.5
R204 VDD.n2 VDD.n1 7.5
R205 VDD.n6 VDD.n5 7.5
R206 VDD.n9 VDD.n8 7.5
R207 VDD.n19 VDD.n18 7.5
R208 VDD.n14 VDD.n0 7.5
R209 VDD.n51 VDD.n48 6.772
R210 VDD.n62 VDD.n46 6.772
R211 VDD.n60 VDD.n57 6.772
R212 VDD.n56 VDD.n53 6.772
R213 VDD.n123 VDD.n108 6.772
R214 VDD.n121 VDD.n118 6.772
R215 VDD.n117 VDD.n114 6.772
R216 VDD.n148 VDD.n134 6.772
R217 VDD.n146 VDD.n143 6.772
R218 VDD.n142 VDD.n139 6.772
R219 VDD.n51 VDD.n50 6.772
R220 VDD.n56 VDD.n55 6.772
R221 VDD.n60 VDD.n59 6.772
R222 VDD.n63 VDD.n62 6.772
R223 VDD.n117 VDD.n116 6.772
R224 VDD.n121 VDD.n120 6.772
R225 VDD.n124 VDD.n123 6.772
R226 VDD.n142 VDD.n141 6.772
R227 VDD.n146 VDD.n145 6.772
R228 VDD.n149 VDD.n148 6.772
R229 VDD.n209 VDD.n208 6.772
R230 VDD.n196 VDD.n193 6.772
R231 VDD.n201 VDD.n198 6.772
R232 VDD.n206 VDD.n203 6.772
R233 VDD.n206 VDD.n205 6.772
R234 VDD.n201 VDD.n200 6.772
R235 VDD.n196 VDD.n195 6.772
R236 VDD.n208 VDD.n192 6.772
R237 VDD.n16 VDD.n15 6.458
R238 VDD.n112 VDD.n111 6.202
R239 VDD.n137 VDD.n136 6.202
R240 VDD.n226 VDD.n222 5.903
R241 VDD.n88 VDD.n87 4.576
R242 VDD.n229 VDD.n228 4.576
R243 VDD.n166 VDD.n165 4.576
R244 VDD.n100 VDD.n97 2.754
R245 VDD.n158 VDD.n155 2.754
R246 VDD.n74 VDD.n71 2.361
R247 VDD.n184 VDD.n181 2.361
R248 VDD.n28 VDD.n24 1.967
R249 VDD.n38 VDD.n37 1.967
R250 VDD.n14 VDD.n7 1.329
R251 VDD.n14 VDD.n10 1.329
R252 VDD.n14 VDD.n11 1.329
R253 VDD.n14 VDD.n13 1.329
R254 VDD.n15 VDD.n14 0.696
R255 VDD.n14 VDD.n4 0.696
R256 VDD.n61 VDD.n60 0.365
R257 VDD.n61 VDD.n56 0.365
R258 VDD.n61 VDD.n51 0.365
R259 VDD.n62 VDD.n61 0.365
R260 VDD.n122 VDD.n121 0.365
R261 VDD.n122 VDD.n117 0.365
R262 VDD.n123 VDD.n122 0.365
R263 VDD.n147 VDD.n146 0.365
R264 VDD.n147 VDD.n142 0.365
R265 VDD.n148 VDD.n147 0.365
R266 VDD.n207 VDD.n206 0.365
R267 VDD.n207 VDD.n201 0.365
R268 VDD.n207 VDD.n196 0.365
R269 VDD.n208 VDD.n207 0.365
R270 VDD.n70 VDD.n43 0.29
R271 VDD.n131 VDD.n105 0.29
R272 VDD.n216 VDD.n189 0.29
R273 VDD.n154 VDD 0.207
R274 VDD.n91 VDD.n86 0.181
R275 VDD.n236 VDD.n232 0.181
R276 VDD.n175 VDD.n169 0.181
R277 VDD.n33 VDD.n29 0.157
R278 VDD.n39 VDD.n33 0.157
R279 VDD.n43 VDD.n39 0.145
R280 VDD.n75 VDD.n70 0.145
R281 VDD.n80 VDD.n75 0.145
R282 VDD.n86 VDD.n80 0.145
R283 VDD.n96 VDD.n91 0.145
R284 VDD.n101 VDD.n96 0.145
R285 VDD.n105 VDD.n101 0.145
R286 VDD.n244 VDD.n240 0.145
R287 VDD.n240 VDD.n236 0.145
R288 VDD.n232 VDD.n227 0.145
R289 VDD.n227 VDD.n220 0.145
R290 VDD.n220 VDD.n216 0.145
R291 VDD.n189 VDD.n185 0.145
R292 VDD.n185 VDD.n180 0.145
R293 VDD.n180 VDD.n175 0.145
R294 VDD.n169 VDD.n164 0.145
R295 VDD.n164 VDD.n159 0.145
R296 VDD.n159 VDD.n154 0.145
R297 VDD VDD.n131 0.078
R298 VDD VDD.n244 0.066
R299 D.n0 D.t2 472.359
R300 D.n0 D.t0 384.527
R301 D.n1 D.t1 267.725
R302 D.n1 D.n0 83.507
R303 D.n2 D.n1 76
R304 D.n2 D 0.046
R305 a_1549_1050.n0 a_1549_1050.t6 512.525
R306 a_1549_1050.n0 a_1549_1050.t5 371.139
R307 a_1549_1050.n8 a_1549_1050.n6 232.158
R308 a_1549_1050.n1 a_1549_1050.n0 226.306
R309 a_1549_1050.n1 a_1549_1050.t7 157.328
R310 a_1549_1050.n6 a_1549_1050.n1 153.043
R311 a_1549_1050.n6 a_1549_1050.n5 130.933
R312 a_1549_1050.n8 a_1549_1050.n7 76.002
R313 a_1549_1050.n5 a_1549_1050.n4 30
R314 a_1549_1050.n3 a_1549_1050.n2 24.383
R315 a_1549_1050.n5 a_1549_1050.n3 23.684
R316 a_1549_1050.n7 a_1549_1050.t4 14.282
R317 a_1549_1050.n7 a_1549_1050.t3 14.282
R318 a_1549_1050.n9 a_1549_1050.t0 14.282
R319 a_1549_1050.t1 a_1549_1050.n9 14.282
R320 a_1549_1050.n9 a_1549_1050.n8 12.848
R321 A.n0 A.t0 480.392
R322 A.n0 A.t2 403.272
R323 A.n1 A.t1 230.374
R324 A.n1 A.n0 151.553
R325 A.n2 A.n1 76
R326 A.n2 A 0.046
R327 Y.n5 Y.n0 210.56
R328 Y.n5 Y.n4 152.462
R329 Y.n6 Y.n5 76
R330 Y.n4 Y.n3 30
R331 Y.n2 Y.n1 24.383
R332 Y.n4 Y.n2 23.684
R333 Y.n0 Y.t0 14.282
R334 Y.n0 Y.t1 14.282
R335 Y.n6 Y 0.046
R336 GND.n30 GND.n28 219.745
R337 GND.n100 GND.n99 219.745
R338 GND.n63 GND.n62 219.745
R339 GND.n30 GND.n29 85.529
R340 GND.n100 GND.n98 85.529
R341 GND.n63 GND.n61 85.529
R342 GND.n9 GND.n1 76.145
R343 GND.n70 GND.n69 76
R344 GND.n9 GND.n8 76
R345 GND.n17 GND.n16 76
R346 GND.n24 GND.n23 76
R347 GND.n27 GND.n26 76
R348 GND.n34 GND.n33 76
R349 GND.n37 GND.n36 76
R350 GND.n40 GND.n39 76
R351 GND.n43 GND.n42 76
R352 GND.n46 GND.n45 76
R353 GND.n54 GND.n53 76
R354 GND.n57 GND.n56 76
R355 GND.n60 GND.n59 76
R356 GND.n67 GND.n66 76
R357 GND.n137 GND.n136 76
R358 GND.n130 GND.n129 76
R359 GND.n124 GND.n123 76
R360 GND.n118 GND.n117 76
R361 GND.n115 GND.n114 76
R362 GND.n110 GND.n109 76
R363 GND.n103 GND.n102 76
R364 GND.n96 GND.n95 76
R365 GND.n93 GND.n92 76
R366 GND.n90 GND.n89 76
R367 GND.n87 GND.n86 76
R368 GND.n84 GND.n83 76
R369 GND.n81 GND.n80 76
R370 GND.n73 GND.n72 76
R371 GND.n51 GND.n50 63.835
R372 GND.n78 GND.n77 63.835
R373 GND.n5 GND.n4 35.01
R374 GND.n3 GND.n2 29.127
R375 GND.n50 GND.n49 28.421
R376 GND.n77 GND.n76 28.421
R377 GND.n50 GND.n48 25.263
R378 GND.n77 GND.n75 25.263
R379 GND.n48 GND.n47 24.383
R380 GND.n75 GND.n74 24.383
R381 GND.n12 GND.t4 20.794
R382 GND.n6 GND.n5 19.735
R383 GND.n14 GND.n13 19.735
R384 GND.n22 GND.n21 19.735
R385 GND.n112 GND.n111 19.735
R386 GND.n122 GND.n121 19.735
R387 GND.n128 GND.n127 19.735
R388 GND.n134 GND.n133 19.735
R389 GND.n108 GND.n107 19.735
R390 GND.n127 GND.t2 19.724
R391 GND.n111 GND.t1 19.724
R392 GND.n5 GND.n3 19.017
R393 GND.n33 GND.n31 14.167
R394 GND.n66 GND.n64 14.167
R395 GND.n102 GND.n101 14.167
R396 GND.n72 GND.n71 13.653
R397 GND.n80 GND.n79 13.653
R398 GND.n83 GND.n82 13.653
R399 GND.n86 GND.n85 13.653
R400 GND.n89 GND.n88 13.653
R401 GND.n92 GND.n91 13.653
R402 GND.n95 GND.n94 13.653
R403 GND.n102 GND.n97 13.653
R404 GND.n109 GND.n104 13.653
R405 GND.n114 GND.n113 13.653
R406 GND.n117 GND.n116 13.653
R407 GND.n123 GND.n119 13.653
R408 GND.n129 GND.n125 13.653
R409 GND.n136 GND.n135 13.653
R410 GND.n66 GND.n65 13.653
R411 GND.n59 GND.n58 13.653
R412 GND.n56 GND.n55 13.653
R413 GND.n53 GND.n52 13.653
R414 GND.n45 GND.n44 13.653
R415 GND.n42 GND.n41 13.653
R416 GND.n39 GND.n38 13.653
R417 GND.n36 GND.n35 13.653
R418 GND.n33 GND.n32 13.653
R419 GND.n26 GND.n25 13.653
R420 GND.n23 GND.n18 13.653
R421 GND.n16 GND.n15 13.653
R422 GND.n8 GND.n7 13.653
R423 GND.n21 GND.n20 12.837
R424 GND.n107 GND.n106 12.837
R425 GND.n133 GND.n132 11.605
R426 GND.n132 GND.n131 9.809
R427 GND.n123 GND.n122 8.854
R428 GND.n20 GND.n19 7.566
R429 GND.n106 GND.n105 7.566
R430 GND.n31 GND.n30 7.312
R431 GND.n101 GND.n100 7.312
R432 GND.n64 GND.n63 7.312
R433 GND.t2 GND.n126 7.04
R434 GND.n121 GND.n120 5.774
R435 GND.n11 GND.n10 4.551
R436 GND.n8 GND.n6 3.935
R437 GND.n53 GND.n51 3.935
R438 GND.n129 GND.n128 3.935
R439 GND.n114 GND.n112 3.935
R440 GND.n80 GND.n78 3.935
R441 GND.n23 GND.n22 3.541
R442 GND.t4 GND.n11 2.238
R443 GND.n136 GND.n134 0.983
R444 GND.n109 GND.n108 0.983
R445 GND.n1 GND.n0 0.596
R446 GND.n69 GND.n68 0.596
R447 GND.n13 GND.n12 0.358
R448 GND.n34 GND.n27 0.29
R449 GND.n67 GND.n60 0.29
R450 GND.n103 GND.n96 0.29
R451 GND.n70 GND 0.207
R452 GND.n16 GND.n14 0.196
R453 GND.n46 GND.n43 0.181
R454 GND.n124 GND.n118 0.181
R455 GND.n87 GND.n84 0.181
R456 GND.n17 GND.n9 0.157
R457 GND.n24 GND.n17 0.157
R458 GND.n27 GND.n24 0.145
R459 GND.n37 GND.n34 0.145
R460 GND.n40 GND.n37 0.145
R461 GND.n43 GND.n40 0.145
R462 GND.n54 GND.n46 0.145
R463 GND.n57 GND.n54 0.145
R464 GND.n60 GND.n57 0.145
R465 GND.n137 GND.n130 0.145
R466 GND.n130 GND.n124 0.145
R467 GND.n118 GND.n115 0.145
R468 GND.n115 GND.n110 0.145
R469 GND.n110 GND.n103 0.145
R470 GND.n96 GND.n93 0.145
R471 GND.n93 GND.n90 0.145
R472 GND.n90 GND.n87 0.145
R473 GND.n84 GND.n81 0.145
R474 GND.n81 GND.n73 0.145
R475 GND.n73 GND.n70 0.145
R476 GND GND.n67 0.078
R477 GND GND.n137 0.066
R478 a_112_101.n12 a_112_101.n11 26.811
R479 a_112_101.n6 a_112_101.n5 24.977
R480 a_112_101.n2 a_112_101.n1 24.877
R481 a_112_101.t0 a_112_101.n2 12.677
R482 a_112_101.t0 a_112_101.n3 11.595
R483 a_112_101.t1 a_112_101.n8 8.137
R484 a_112_101.t0 a_112_101.n4 7.273
R485 a_112_101.t0 a_112_101.n0 6.109
R486 a_112_101.t1 a_112_101.n7 4.864
R487 a_112_101.t0 a_112_101.n12 2.074
R488 a_112_101.n7 a_112_101.n6 1.13
R489 a_112_101.n12 a_112_101.t1 0.937
R490 a_112_101.t1 a_112_101.n10 0.804
R491 a_112_101.n10 a_112_101.n9 0.136
R492 a_1444_101.t0 a_1444_101.n1 34.62
R493 a_1444_101.t0 a_1444_101.n0 8.137
R494 a_1444_101.t0 a_1444_101.n2 4.69
R495 B.n0 B.t0 472.359
R496 B.n0 B.t2 384.527
R497 B.n1 B.t1 214.619
R498 B.n1 B.n0 136.613
R499 B.n2 B.n1 76
R500 B.n2 B 0.046
C6 VDD GND 9.85fF
C7 a_1444_101.n0 GND 0.05fF
C8 a_1444_101.n1 GND 0.12fF
C9 a_1444_101.n2 GND 0.04fF
C10 a_112_101.n0 GND 0.02fF
C11 a_112_101.n1 GND 0.10fF
C12 a_112_101.n2 GND 0.06fF
C13 a_112_101.n3 GND 0.06fF
C14 a_112_101.n4 GND 0.00fF
C15 a_112_101.n5 GND 0.04fF
C16 a_112_101.n6 GND 0.05fF
C17 a_112_101.n7 GND 0.02fF
C18 a_112_101.n8 GND 0.05fF
C19 a_112_101.n9 GND 0.07fF
C20 a_112_101.n10 GND 0.17fF
C21 a_112_101.t1 GND 0.22fF
C22 a_112_101.n11 GND 0.09fF
C23 a_112_101.n12 GND 0.00fF
C24 Y.n0 GND 0.83fF
C25 Y.n1 GND 0.04fF
C26 Y.n2 GND 0.06fF
C27 Y.n3 GND 0.04fF
C28 Y.n4 GND 0.24fF
C29 Y.n5 GND 0.47fF
C30 Y.n6 GND 0.01fF
C31 a_1549_1050.n0 GND 0.35fF
C32 a_1549_1050.n1 GND 0.45fF
C33 a_1549_1050.n2 GND 0.03fF
C34 a_1549_1050.n3 GND 0.04fF
C35 a_1549_1050.n4 GND 0.03fF
C36 a_1549_1050.n5 GND 0.16fF
C37 a_1549_1050.n6 GND 0.46fF
C38 a_1549_1050.n7 GND 0.50fF
C39 a_1549_1050.n8 GND 0.31fF
C40 a_1549_1050.n9 GND 0.42fF
C41 VDD.n0 GND 0.11fF
C42 VDD.n1 GND 0.02fF
C43 VDD.n2 GND 0.02fF
C44 VDD.n3 GND 0.04fF
C45 VDD.n4 GND 0.01fF
C46 VDD.n5 GND 0.02fF
C47 VDD.n6 GND 0.02fF
C48 VDD.n8 GND 0.02fF
C49 VDD.n9 GND 0.02fF
C50 VDD.n12 GND 0.02fF
C51 VDD.n14 GND 0.42fF
C52 VDD.n16 GND 0.03fF
C53 VDD.n17 GND 0.02fF
C54 VDD.n18 GND 0.02fF
C55 VDD.n19 GND 0.02fF
C56 VDD.n20 GND 0.03fF
C57 VDD.n21 GND 0.25fF
C58 VDD.n22 GND 0.02fF
C59 VDD.n23 GND 0.03fF
C60 VDD.n24 GND 0.05fF
C61 VDD.n25 GND 0.14fF
C62 VDD.n26 GND 0.19fF
C63 VDD.n27 GND 0.01fF
C64 VDD.n28 GND 0.01fF
C65 VDD.n29 GND 0.06fF
C66 VDD.n30 GND 0.16fF
C67 VDD.n31 GND 0.01fF
C68 VDD.n32 GND 0.02fF
C69 VDD.n33 GND 0.02fF
C70 VDD.n34 GND 0.14fF
C71 VDD.n35 GND 0.19fF
C72 VDD.n36 GND 0.01fF
C73 VDD.n37 GND 0.06fF
C74 VDD.n38 GND 0.01fF
C75 VDD.n39 GND 0.02fF
C76 VDD.n40 GND 0.25fF
C77 VDD.n41 GND 0.01fF
C78 VDD.n42 GND 0.02fF
C79 VDD.n43 GND 0.03fF
C80 VDD.n44 GND 0.02fF
C81 VDD.n45 GND 0.02fF
C82 VDD.n46 GND 0.02fF
C83 VDD.n47 GND 0.17fF
C84 VDD.n48 GND 0.04fF
C85 VDD.n49 GND 0.03fF
C86 VDD.n50 GND 0.02fF
C87 VDD.n52 GND 0.02fF
C88 VDD.n53 GND 0.02fF
C89 VDD.n54 GND 0.02fF
C90 VDD.n55 GND 0.02fF
C91 VDD.n57 GND 0.02fF
C92 VDD.n58 GND 0.02fF
C93 VDD.n59 GND 0.02fF
C94 VDD.n61 GND 0.25fF
C95 VDD.n63 GND 0.02fF
C96 VDD.n64 GND 0.02fF
C97 VDD.n65 GND 0.03fF
C98 VDD.n66 GND 0.02fF
C99 VDD.n67 GND 0.25fF
C100 VDD.n68 GND 0.01fF
C101 VDD.n69 GND 0.02fF
C102 VDD.n70 GND 0.03fF
C103 VDD.n71 GND 0.05fF
C104 VDD.n72 GND 0.23fF
C105 VDD.n73 GND 0.01fF
C106 VDD.n74 GND 0.01fF
C107 VDD.n75 GND 0.02fF
C108 VDD.n76 GND 0.13fF
C109 VDD.n77 GND 0.16fF
C110 VDD.n78 GND 0.01fF
C111 VDD.n79 GND 0.02fF
C112 VDD.n80 GND 0.02fF
C113 VDD.n81 GND 0.10fF
C114 VDD.n82 GND 0.02fF
C115 VDD.n83 GND 0.28fF
C116 VDD.n84 GND 0.01fF
C117 VDD.n85 GND 0.02fF
C118 VDD.n86 GND 0.02fF
C119 VDD.n87 GND 0.16fF
C120 VDD.n88 GND 0.13fF
C121 VDD.n89 GND 0.01fF
C122 VDD.n90 GND 0.02fF
C123 VDD.n91 GND 0.02fF
C124 VDD.n92 GND 0.13fF
C125 VDD.n93 GND 0.15fF
C126 VDD.n94 GND 0.01fF
C127 VDD.n95 GND 0.02fF
C128 VDD.n96 GND 0.02fF
C129 VDD.n97 GND 0.06fF
C130 VDD.n98 GND 0.23fF
C131 VDD.n99 GND 0.01fF
C132 VDD.n100 GND 0.01fF
C133 VDD.n101 GND 0.02fF
C134 VDD.n102 GND 0.25fF
C135 VDD.n103 GND 0.01fF
C136 VDD.n104 GND 0.02fF
C137 VDD.n105 GND 0.03fF
C138 VDD.n106 GND 0.02fF
C139 VDD.n107 GND 0.02fF
C140 VDD.n108 GND 0.02fF
C141 VDD.n109 GND 0.20fF
C142 VDD.n110 GND 0.04fF
C143 VDD.n111 GND 0.03fF
C144 VDD.n112 GND 0.02fF
C145 VDD.n113 GND 0.02fF
C146 VDD.n114 GND 0.02fF
C147 VDD.n115 GND 0.02fF
C148 VDD.n116 GND 0.02fF
C149 VDD.n118 GND 0.02fF
C150 VDD.n119 GND 0.02fF
C151 VDD.n120 GND 0.02fF
C152 VDD.n122 GND 0.25fF
C153 VDD.n124 GND 0.02fF
C154 VDD.n125 GND 0.02fF
C155 VDD.n126 GND 0.03fF
C156 VDD.n127 GND 0.02fF
C157 VDD.n128 GND 0.25fF
C158 VDD.n129 GND 0.01fF
C159 VDD.n130 GND 0.02fF
C160 VDD.n131 GND 0.03fF
C161 VDD.n132 GND 0.02fF
C162 VDD.n133 GND 0.02fF
C163 VDD.n134 GND 0.02fF
C164 VDD.n135 GND 0.14fF
C165 VDD.n136 GND 0.03fF
C166 VDD.n137 GND 0.02fF
C167 VDD.n138 GND 0.02fF
C168 VDD.n139 GND 0.02fF
C169 VDD.n140 GND 0.02fF
C170 VDD.n141 GND 0.02fF
C171 VDD.n143 GND 0.02fF
C172 VDD.n144 GND 0.02fF
C173 VDD.n145 GND 0.02fF
C174 VDD.n147 GND 0.42fF
C175 VDD.n149 GND 0.03fF
C176 VDD.n150 GND 0.03fF
C177 VDD.n151 GND 0.25fF
C178 VDD.n152 GND 0.02fF
C179 VDD.n153 GND 0.03fF
C180 VDD.n154 GND 0.03fF
C181 VDD.n155 GND 0.06fF
C182 VDD.n156 GND 0.23fF
C183 VDD.n157 GND 0.01fF
C184 VDD.n158 GND 0.01fF
C185 VDD.n159 GND 0.02fF
C186 VDD.n160 GND 0.13fF
C187 VDD.n161 GND 0.15fF
C188 VDD.n162 GND 0.01fF
C189 VDD.n163 GND 0.02fF
C190 VDD.n164 GND 0.02fF
C191 VDD.n165 GND 0.16fF
C192 VDD.n166 GND 0.13fF
C193 VDD.n167 GND 0.01fF
C194 VDD.n168 GND 0.02fF
C195 VDD.n169 GND 0.02fF
C196 VDD.n170 GND 0.10fF
C197 VDD.n171 GND 0.02fF
C198 VDD.n172 GND 0.28fF
C199 VDD.n173 GND 0.01fF
C200 VDD.n174 GND 0.02fF
C201 VDD.n175 GND 0.02fF
C202 VDD.n176 GND 0.13fF
C203 VDD.n177 GND 0.16fF
C204 VDD.n178 GND 0.01fF
C205 VDD.n179 GND 0.02fF
C206 VDD.n180 GND 0.02fF
C207 VDD.n181 GND 0.05fF
C208 VDD.n182 GND 0.23fF
C209 VDD.n183 GND 0.01fF
C210 VDD.n184 GND 0.01fF
C211 VDD.n185 GND 0.02fF
C212 VDD.n186 GND 0.25fF
C213 VDD.n187 GND 0.01fF
C214 VDD.n188 GND 0.02fF
C215 VDD.n189 GND 0.03fF
C216 VDD.n190 GND 0.02fF
C217 VDD.n191 GND 0.02fF
C218 VDD.n192 GND 0.02fF
C219 VDD.n193 GND 0.02fF
C220 VDD.n194 GND 0.02fF
C221 VDD.n195 GND 0.02fF
C222 VDD.n197 GND 0.02fF
C223 VDD.n198 GND 0.02fF
C224 VDD.n199 GND 0.02fF
C225 VDD.n200 GND 0.02fF
C226 VDD.n202 GND 0.03fF
C227 VDD.n203 GND 0.02fF
C228 VDD.n204 GND 0.20fF
C229 VDD.n205 GND 0.04fF
C230 VDD.n207 GND 0.25fF
C231 VDD.n209 GND 0.02fF
C232 VDD.n210 GND 0.02fF
C233 VDD.n211 GND 0.03fF
C234 VDD.n212 GND 0.02fF
C235 VDD.n213 GND 0.25fF
C236 VDD.n214 GND 0.01fF
C237 VDD.n215 GND 0.02fF
C238 VDD.n216 GND 0.03fF
C239 VDD.n217 GND 0.23fF
C240 VDD.n218 GND 0.01fF
C241 VDD.n219 GND 0.02fF
C242 VDD.n220 GND 0.02fF
C243 VDD.n221 GND 0.10fF
C244 VDD.n222 GND 0.02fF
C245 VDD.n223 GND 0.13fF
C246 VDD.n224 GND 0.15fF
C247 VDD.n225 GND 0.01fF
C248 VDD.n226 GND 0.02fF
C249 VDD.n227 GND 0.02fF
C250 VDD.n228 GND 0.16fF
C251 VDD.n229 GND 0.13fF
C252 VDD.n230 GND 0.01fF
C253 VDD.n231 GND 0.02fF
C254 VDD.n232 GND 0.02fF
C255 VDD.n233 GND 0.28fF
C256 VDD.n234 GND 0.01fF
C257 VDD.n235 GND 0.02fF
C258 VDD.n236 GND 0.02fF
C259 VDD.n237 GND 0.25fF
C260 VDD.n238 GND 0.01fF
C261 VDD.n239 GND 0.02fF
C262 VDD.n240 GND 0.02fF
C263 VDD.n241 GND 0.25fF
C264 VDD.n242 GND 0.01fF
C265 VDD.n243 GND 0.02fF
C266 VDD.n244 GND 0.02fF
C267 a_217_1050.n0 GND 0.03fF
C268 a_217_1050.n1 GND 0.42fF
C269 a_217_1050.n2 GND 0.50fF
C270 a_217_1050.n3 GND 0.32fF
C271 a_217_1050.n4 GND 0.36fF
C272 a_217_1050.t6 GND 0.37fF
C273 a_217_1050.n5 GND 0.45fF
C274 a_217_1050.n6 GND 0.48fF
C275 a_217_1050.n7 GND 0.03fF
C276 a_217_1050.n8 GND 0.16fF
C277 a_217_1050.n9 GND 0.04fF
C278 a_864_209.n0 GND 0.39fF
C279 a_864_209.n1 GND 0.46fF
C280 a_864_209.n2 GND 0.05fF
C281 a_864_209.n3 GND 0.03fF
C282 a_864_209.n4 GND 0.10fF
C283 a_864_209.n5 GND 0.04fF
C284 a_864_209.n6 GND 0.05fF
C285 a_864_209.n7 GND 0.16fF
C286 a_864_209.n8 GND 0.27fF
C287 a_864_209.n9 GND 0.47fF
C288 a_864_209.n10 GND 0.63fF
C289 a_797_1051.n0 GND 0.54fF
.ends
