* SPICE3 file created from TMRDFFSNRNQX1.ext - technology: sky130A

.subckt TMRDFFSNRNQX1 Q D CLK SN RN VDD VSS
X0 a_13105_989 RN a_14802_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X1 VDD RN a_15669_1050 VDD sky130_fd_pr__pfet_01v8 ad=0.004346 pd=3.5146 as=0 ps=0 w=2 l=0.15 M=2
X2 a_599_989 CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X3 VDD RN a_9897_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X4 VSS a_599_989 a_3939_103 VSS sky130_fd_pr__nfet_01v8 ad=0.0049019 pd=4.107 as=0 ps=0 w=3 l=0.15
X5 VDD CLK a_1561_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X6 a_11821_1050 a_12143_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X7 a_7333_989 RN a_9030_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X8 VDD a_13105_989 a_13745_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X9 VDD a_277_1050 a_2201_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X10 a_7333_989 CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X11 a_10219_989 SN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X12 VDD a_7333_989 a_6371_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X13 VDD CLK a_12143_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X14 a_13105_989 RN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X15 a_5182_210 SN a_4901_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X16 a_7106_210 CLK a_6825_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X17 a_1334_210 CLK a_1053_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X18 VDD RN a_277_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X19 a_15669_1050 a_15991_989 a_15764_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X20 a_3258_210 CLK a_2977_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X21 a_6371_989 a_6049_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X22 a_13745_1050 a_13105_989 a_13840_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X23 VSS a_6049_1050 a_6825_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X24 VDD a_7973_1050 a_7333_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X25 VDD a_9897_1050 a_10219_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X26 a_17533_1051 a_15991_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X27 a_599_989 a_1561_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X28 VSS a_4125_1050 a_4901_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X29 a_15991_989 a_15669_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X30 VDD RN a_1561_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X31 a_9897_1050 a_6371_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X32 a_4125_1050 a_599_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X33 VDD SN a_2201_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X34 a_4125_1050 a_4447_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X35 VSS a_4447_989 a_18760_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X36 VSS a_15991_989 a_18094_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X37 VDD a_6371_989 a_6049_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X38 a_18197_1051 a_15991_989 a_17533_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X39 a_6144_210 RN a_5863_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X40 VSS D a_11635_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X41 VDD a_599_989 a_277_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X42 a_15991_989 a_13105_989 a_16726_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X43 a_8068_210 SN a_7787_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X44 a_13745_1050 SN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X45 VSS a_6049_1050 a_7787_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X46 a_17533_1051 a_10219_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X47 a_12143_989 a_11821_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X48 VSS a_6371_989 a_9711_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X49 VDD a_13745_1050 a_13105_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X50 a_17708_209 a_10219_989 a_18760_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X51 a_15991_989 SN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X52 VSS D a_5863_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X53 a_15669_1050 a_12143_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X54 a_4125_1050 RN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X55 VDD a_17708_209 Q VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.0058 ps=4.58 w=2 l=0.15 M=2
X56 VDD a_1561_989 a_2201_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X57 VDD RN a_6049_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X58 a_277_1050 a_599_989 a_372_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X59 a_7973_1050 a_7333_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X60 a_9897_1050 a_10219_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X61 VDD a_13105_989 a_15991_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X62 a_1561_989 a_2201_1050 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X63 a_9030_210 CLK a_8749_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X64 a_18197_1051 a_4447_989 a_17533_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X65 VDD a_4125_1050 a_4447_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X66 a_6371_989 CLK VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X67 a_6049_1050 D VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X68 VSS a_11821_1050 a_12597_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X69 VSS a_13745_1050 a_14521_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X70 a_17708_209 a_10219_989 a_18197_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X71 VSS a_9897_1050 a_10673_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X72 a_277_1050 D VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X73 VSS a_7973_1050 a_8749_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X74 Q a_17708_209 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0 ps=0 w=3 l=0.15
X75 VDD CLK a_13105_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X76 VDD a_11821_1050 a_13745_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X77 a_10219_989 a_7333_989 VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X78 VDD a_13105_989 a_12143_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X79 VSS D a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X80 VDD a_277_1050 a_599_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X81 a_11916_210 RN a_11635_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X82 VDD RN a_11821_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X83 a_9992_210 RN a_9711_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X84 VDD SN a_4447_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X85 a_18197_1051 a_4447_989 a_17708_209 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X86 VDD a_15991_989 a_15669_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X87 VSS a_15991_989 a_17428_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X88 VDD RN a_7333_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X89 VDD SN a_7973_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X90 VSS a_11821_1050 a_13559_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X91 VSS a_12143_989 a_15483_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X92 a_14802_210 CLK a_14521_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X93 a_17708_209 a_4447_989 a_18094_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X94 a_10954_210 SN a_10673_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X95 a_16726_210 SN a_16445_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X96 a_12878_210 CLK a_12597_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X97 VDD a_1561_989 a_4447_989 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X98 VSS a_15669_1050 a_16445_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X99 a_2201_1050 a_1561_989 a_2296_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X100 a_372_210 RN a_91_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X101 VDD a_6049_1050 a_7973_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X102 a_4125_1050 a_4447_989 a_4220_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X103 a_11821_1050 D VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X104 a_13840_210 SN a_13559_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X105 a_15764_210 RN a_15483_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X106 VSS a_277_1050 a_2015_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X107 a_599_989 a_1561_989 a_1334_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X108 a_6371_989 a_7333_989 a_7106_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X109 a_1561_989 RN a_3258_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X110 a_4447_989 a_1561_989 a_5182_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X111 a_11821_1050 a_12143_989 a_11916_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X112 a_17708_209 a_10219_989 a_17428_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X113 a_6049_1050 a_6371_989 a_6144_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X114 a_9897_1050 a_10219_989 a_9992_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X115 a_7973_1050 a_7333_989 a_8068_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X116 VSS a_2201_1050 a_2977_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X117 VSS a_277_1050 a_1053_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X118 a_4220_210 RN a_3939_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X119 a_10219_989 a_7333_989 a_10954_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X120 a_2296_210 SN a_2015_103 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X121 a_12143_989 a_13105_989 a_12878_210 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
C0 CLK D 12.06f
C1 a_4447_989 RN 4.97f
C2 a_7333_989 VDD 3.43f
C3 a_4447_989 a_12143_989 4.03f
C4 a_10219_989 RN 2.33f
C5 VDD a_11821_1050 3.19f
C6 a_4447_989 a_10219_989 3.51f
C7 CLK VDD 8.69f
C8 RN SN 16.07f
C9 a_4447_989 SN 3.36f
C10 a_7973_1050 VDD 2.84f
C11 VDD a_9897_1050 2.84f
C12 a_1561_989 CLK 2.10f
C13 VDD a_13105_989 3.43f
C14 VDD a_6371_989 3.14f
C15 a_4447_989 CLK 2.02f
C16 VDD D 11.48f
C17 a_10219_989 CLK 3.88f
C18 VDD a_13745_1050 2.84f
C19 a_277_1050 VDD 3.19f
C20 a_4447_989 a_6371_989 4.03f
C21 a_2201_1050 VDD 2.84f
C22 a_1561_989 D 4.57f
C23 a_12143_989 a_13105_989 3.35f
C24 a_599_989 VDD 3.14f
C25 a_10219_989 a_13105_989 4.57f
C26 a_6049_1050 VDD 3.19f
C27 a_7333_989 CLK 2.10f
C28 RN D 2.36f
C29 VDD a_17533_1051 3.12f
C30 a_15991_989 VDD 3.96f
C31 a_1561_989 VDD 3.43f
C32 VDD a_15669_1050 2.84f
C33 a_1561_989 a_599_989 3.35f
C34 RN VDD 2.65f
C35 a_7333_989 a_6371_989 3.35f
C36 a_4447_989 VDD 3.52f
C37 a_12143_989 VDD 3.14f
C38 a_4125_1050 VDD 2.84f
C39 a_10219_989 VDD 9.84f
C40 a_7333_989 D 4.57f
C41 SN VSS 7.77f
C42 RN VSS 8.35f
C43 VDD VSS 32.47f
C44 a_4447_989 VSS 5.93f **FLOATING
.ends
