* SPICE3 file created from TMRDFFSNRNQNX1.ext - technology: sky130A

.subckt TMRDFFSNRNQNX1 Q D CLK SN RN VDD GND
X0 GND m1_4715_501# votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X1 GND m1_4715_501# votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X2 GND m1_16259_427# votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X3 votern3x1_pcell_0/a_805_1331# m1_4715_501# VDD VDD pshort w=2 l=0.15
X4 Q m1_16259_427# votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X5 votern3x1_pcell_0/a_805_1331# m1_10453_649# VDD VDD pshort w=2 l=0.15
X6 votern3x1_pcell_0/a_893_1059# m1_16259_427# votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X7 votern3x1_pcell_0/a_893_1059# m1_4715_501# votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X8 Q m1_16259_427# votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X9 Q m1_10453_649# votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X10 Q m1_10453_649# votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X11 Q m1_10453_649# votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X12 GND D dffsnrnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X13 dffsnrnx1_pcell_0/m1_831_501# dffsnrnx1_pcell_0/m1_716_649# dffsnrnx1_pcell_0/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X14 dffsnrnx1_pcell_0/nand3x1_pcell_0/li_393_182# RN dffsnrnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X15 VDD D dffsnrnx1_pcell_0/m1_831_501# VDD pshort w=2 l=0.15
X16 VDD RN dffsnrnx1_pcell_0/m1_831_501# VDD pshort w=2 l=0.15
X17 VDD dffsnrnx1_pcell_0/m1_716_649# dffsnrnx1_pcell_0/m1_831_501# VDD pshort w=2 l=0.15
X18 GND dffsnrnx1_pcell_0/m1_831_501# dffsnrnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X19 dffsnrnx1_pcell_0/m1_716_649# dffsnrnx1_pcell_0/m1_1660_723# dffsnrnx1_pcell_0/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X20 dffsnrnx1_pcell_0/nand3x1_pcell_1/li_393_182# CLK dffsnrnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X21 VDD dffsnrnx1_pcell_0/m1_831_501# dffsnrnx1_pcell_0/m1_716_649# VDD pshort w=2 l=0.15
X22 VDD CLK dffsnrnx1_pcell_0/m1_716_649# VDD pshort w=2 l=0.15
X23 VDD dffsnrnx1_pcell_0/m1_1660_723# dffsnrnx1_pcell_0/m1_716_649# VDD pshort w=2 l=0.15
X24 GND dffsnrnx1_pcell_0/m1_831_501# dffsnrnx1_pcell_0/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X25 dffsnrnx1_pcell_0/m1_2757_501# dffsnrnx1_pcell_0/m1_1660_723# dffsnrnx1_pcell_0/nand3x1_pcell_2/li_393_182# GND nshort w=3 l=0.15
X26 dffsnrnx1_pcell_0/nand3x1_pcell_2/li_393_182# SN dffsnrnx1_pcell_0/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X27 VDD dffsnrnx1_pcell_0/m1_831_501# dffsnrnx1_pcell_0/m1_2757_501# VDD pshort w=2 l=0.15
X28 VDD SN dffsnrnx1_pcell_0/m1_2757_501# VDD pshort w=2 l=0.15
X29 VDD dffsnrnx1_pcell_0/m1_1660_723# dffsnrnx1_pcell_0/m1_2757_501# VDD pshort w=2 l=0.15
X30 GND dffsnrnx1_pcell_0/m1_2757_501# dffsnrnx1_pcell_0/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X31 dffsnrnx1_pcell_0/m1_1660_723# RN dffsnrnx1_pcell_0/nand3x1_pcell_3/li_393_182# GND nshort w=3 l=0.15
X32 dffsnrnx1_pcell_0/nand3x1_pcell_3/li_393_182# CLK dffsnrnx1_pcell_0/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X33 VDD dffsnrnx1_pcell_0/m1_2757_501# dffsnrnx1_pcell_0/m1_1660_723# VDD pshort w=2 l=0.15
X34 VDD CLK dffsnrnx1_pcell_0/m1_1660_723# VDD pshort w=2 l=0.15
X35 VDD RN dffsnrnx1_pcell_0/m1_1660_723# VDD pshort w=2 l=0.15
X36 GND dffsnrnx1_pcell_0/m1_716_649# dffsnrnx1_pcell_0/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X37 m1_4715_501# m1_4567_649# dffsnrnx1_pcell_0/nand3x1_pcell_4/li_393_182# GND nshort w=3 l=0.15
X38 dffsnrnx1_pcell_0/nand3x1_pcell_4/li_393_182# RN dffsnrnx1_pcell_0/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X39 VDD dffsnrnx1_pcell_0/m1_716_649# m1_4715_501# VDD pshort w=2 l=0.15
X40 VDD RN m1_4715_501# VDD pshort w=2 l=0.15
X41 VDD m1_4567_649# m1_4715_501# VDD pshort w=2 l=0.15
X42 GND m1_4715_501# dffsnrnx1_pcell_0/nand3x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X43 m1_4567_649# dffsnrnx1_pcell_0/m1_1660_723# dffsnrnx1_pcell_0/nand3x1_pcell_5/li_393_182# GND nshort w=3 l=0.15
X44 dffsnrnx1_pcell_0/nand3x1_pcell_5/li_393_182# SN dffsnrnx1_pcell_0/nand3x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X45 VDD m1_4715_501# m1_4567_649# VDD pshort w=2 l=0.15
X46 VDD SN m1_4567_649# VDD pshort w=2 l=0.15
X47 VDD dffsnrnx1_pcell_0/m1_1660_723# m1_4567_649# VDD pshort w=2 l=0.15
X48 GND D dffsnrnx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X49 dffsnrnx1_pcell_1/m1_831_501# dffsnrnx1_pcell_1/m1_716_649# dffsnrnx1_pcell_1/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X50 dffsnrnx1_pcell_1/nand3x1_pcell_0/li_393_182# RN dffsnrnx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X51 VDD D dffsnrnx1_pcell_1/m1_831_501# VDD pshort w=2 l=0.15
X52 VDD RN dffsnrnx1_pcell_1/m1_831_501# VDD pshort w=2 l=0.15
X53 VDD dffsnrnx1_pcell_1/m1_716_649# dffsnrnx1_pcell_1/m1_831_501# VDD pshort w=2 l=0.15
X54 GND dffsnrnx1_pcell_1/m1_831_501# dffsnrnx1_pcell_1/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X55 dffsnrnx1_pcell_1/m1_716_649# dffsnrnx1_pcell_1/m1_1660_723# dffsnrnx1_pcell_1/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X56 dffsnrnx1_pcell_1/nand3x1_pcell_1/li_393_182# CLK dffsnrnx1_pcell_1/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X57 VDD dffsnrnx1_pcell_1/m1_831_501# dffsnrnx1_pcell_1/m1_716_649# VDD pshort w=2 l=0.15
X58 VDD CLK dffsnrnx1_pcell_1/m1_716_649# VDD pshort w=2 l=0.15
X59 VDD dffsnrnx1_pcell_1/m1_1660_723# dffsnrnx1_pcell_1/m1_716_649# VDD pshort w=2 l=0.15
X60 GND dffsnrnx1_pcell_1/m1_831_501# dffsnrnx1_pcell_1/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X61 dffsnrnx1_pcell_1/m1_2757_501# dffsnrnx1_pcell_1/m1_1660_723# dffsnrnx1_pcell_1/nand3x1_pcell_2/li_393_182# GND nshort w=3 l=0.15
X62 dffsnrnx1_pcell_1/nand3x1_pcell_2/li_393_182# SN dffsnrnx1_pcell_1/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X63 VDD dffsnrnx1_pcell_1/m1_831_501# dffsnrnx1_pcell_1/m1_2757_501# VDD pshort w=2 l=0.15
X64 VDD SN dffsnrnx1_pcell_1/m1_2757_501# VDD pshort w=2 l=0.15
X65 VDD dffsnrnx1_pcell_1/m1_1660_723# dffsnrnx1_pcell_1/m1_2757_501# VDD pshort w=2 l=0.15
X66 GND dffsnrnx1_pcell_1/m1_2757_501# dffsnrnx1_pcell_1/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X67 dffsnrnx1_pcell_1/m1_1660_723# RN dffsnrnx1_pcell_1/nand3x1_pcell_3/li_393_182# GND nshort w=3 l=0.15
X68 dffsnrnx1_pcell_1/nand3x1_pcell_3/li_393_182# CLK dffsnrnx1_pcell_1/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X69 VDD dffsnrnx1_pcell_1/m1_2757_501# dffsnrnx1_pcell_1/m1_1660_723# VDD pshort w=2 l=0.15
X70 VDD CLK dffsnrnx1_pcell_1/m1_1660_723# VDD pshort w=2 l=0.15
X71 VDD RN dffsnrnx1_pcell_1/m1_1660_723# VDD pshort w=2 l=0.15
X72 GND dffsnrnx1_pcell_1/m1_716_649# dffsnrnx1_pcell_1/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X73 m1_10453_649# m1_10339_501# dffsnrnx1_pcell_1/nand3x1_pcell_4/li_393_182# GND nshort w=3 l=0.15
X74 dffsnrnx1_pcell_1/nand3x1_pcell_4/li_393_182# RN dffsnrnx1_pcell_1/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X75 VDD dffsnrnx1_pcell_1/m1_716_649# m1_10453_649# VDD pshort w=2 l=0.15
X76 VDD RN m1_10453_649# VDD pshort w=2 l=0.15
X77 VDD m1_10339_501# m1_10453_649# VDD pshort w=2 l=0.15
X78 GND m1_10453_649# dffsnrnx1_pcell_1/nand3x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X79 m1_10339_501# dffsnrnx1_pcell_1/m1_1660_723# dffsnrnx1_pcell_1/nand3x1_pcell_5/li_393_182# GND nshort w=3 l=0.15
X80 dffsnrnx1_pcell_1/nand3x1_pcell_5/li_393_182# SN dffsnrnx1_pcell_1/nand3x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X81 VDD m1_10453_649# m1_10339_501# VDD pshort w=2 l=0.15
X82 VDD SN m1_10339_501# VDD pshort w=2 l=0.15
X83 VDD dffsnrnx1_pcell_1/m1_1660_723# m1_10339_501# VDD pshort w=2 l=0.15
X84 GND D dffsnrnx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X85 dffsnrnx1_pcell_2/m1_831_501# dffsnrnx1_pcell_2/m1_716_649# dffsnrnx1_pcell_2/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X86 dffsnrnx1_pcell_2/nand3x1_pcell_0/li_393_182# RN dffsnrnx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X87 VDD D dffsnrnx1_pcell_2/m1_831_501# VDD pshort w=2 l=0.15
X88 VDD RN dffsnrnx1_pcell_2/m1_831_501# VDD pshort w=2 l=0.15
X89 VDD dffsnrnx1_pcell_2/m1_716_649# dffsnrnx1_pcell_2/m1_831_501# VDD pshort w=2 l=0.15
X90 GND dffsnrnx1_pcell_2/m1_831_501# dffsnrnx1_pcell_2/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X91 dffsnrnx1_pcell_2/m1_716_649# dffsnrnx1_pcell_2/m1_1660_723# dffsnrnx1_pcell_2/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X92 dffsnrnx1_pcell_2/nand3x1_pcell_1/li_393_182# CLK dffsnrnx1_pcell_2/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X93 VDD dffsnrnx1_pcell_2/m1_831_501# dffsnrnx1_pcell_2/m1_716_649# VDD pshort w=2 l=0.15
X94 VDD CLK dffsnrnx1_pcell_2/m1_716_649# VDD pshort w=2 l=0.15
X95 VDD dffsnrnx1_pcell_2/m1_1660_723# dffsnrnx1_pcell_2/m1_716_649# VDD pshort w=2 l=0.15
X96 GND dffsnrnx1_pcell_2/m1_831_501# dffsnrnx1_pcell_2/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X97 dffsnrnx1_pcell_2/m1_2757_501# dffsnrnx1_pcell_2/m1_1660_723# dffsnrnx1_pcell_2/nand3x1_pcell_2/li_393_182# GND nshort w=3 l=0.15
X98 dffsnrnx1_pcell_2/nand3x1_pcell_2/li_393_182# SN dffsnrnx1_pcell_2/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X99 VDD dffsnrnx1_pcell_2/m1_831_501# dffsnrnx1_pcell_2/m1_2757_501# VDD pshort w=2 l=0.15
X100 VDD SN dffsnrnx1_pcell_2/m1_2757_501# VDD pshort w=2 l=0.15
X101 VDD dffsnrnx1_pcell_2/m1_1660_723# dffsnrnx1_pcell_2/m1_2757_501# VDD pshort w=2 l=0.15
X102 GND dffsnrnx1_pcell_2/m1_2757_501# dffsnrnx1_pcell_2/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X103 dffsnrnx1_pcell_2/m1_1660_723# RN dffsnrnx1_pcell_2/nand3x1_pcell_3/li_393_182# GND nshort w=3 l=0.15
X104 dffsnrnx1_pcell_2/nand3x1_pcell_3/li_393_182# CLK dffsnrnx1_pcell_2/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X105 VDD dffsnrnx1_pcell_2/m1_2757_501# dffsnrnx1_pcell_2/m1_1660_723# VDD pshort w=2 l=0.15
X106 VDD CLK dffsnrnx1_pcell_2/m1_1660_723# VDD pshort w=2 l=0.15
X107 VDD RN dffsnrnx1_pcell_2/m1_1660_723# VDD pshort w=2 l=0.15
X108 GND dffsnrnx1_pcell_2/m1_716_649# dffsnrnx1_pcell_2/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X109 m1_16259_427# m1_16111_501# dffsnrnx1_pcell_2/nand3x1_pcell_4/li_393_182# GND nshort w=3 l=0.15
X110 dffsnrnx1_pcell_2/nand3x1_pcell_4/li_393_182# RN dffsnrnx1_pcell_2/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X111 VDD dffsnrnx1_pcell_2/m1_716_649# m1_16259_427# VDD pshort w=2 l=0.15
X112 VDD RN m1_16259_427# VDD pshort w=2 l=0.15
X113 VDD m1_16111_501# m1_16259_427# VDD pshort w=2 l=0.15
X114 GND m1_16259_427# dffsnrnx1_pcell_2/nand3x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X115 m1_16111_501# dffsnrnx1_pcell_2/m1_1660_723# dffsnrnx1_pcell_2/nand3x1_pcell_5/li_393_182# GND nshort w=3 l=0.15
X116 dffsnrnx1_pcell_2/nand3x1_pcell_5/li_393_182# SN dffsnrnx1_pcell_2/nand3x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X117 VDD m1_16259_427# m1_16111_501# VDD pshort w=2 l=0.15
X118 VDD SN m1_16111_501# VDD pshort w=2 l=0.15
X119 VDD dffsnrnx1_pcell_2/m1_1660_723# m1_16111_501# VDD pshort w=2 l=0.15
C0 dffsnrnx1_pcell_1/m1_716_649# dffsnrnx1_pcell_1/m1_1660_723# 3.19fF
C1 dffsnrnx1_pcell_2/m1_716_649# m1_10453_649# 2.03fF
C2 D m1_4715_501# 3.05fF
C3 VDD m1_10453_649# 4.09fF
C4 CLK m1_10453_649# 3.04fF
C5 SN RN 5.64fF
C6 SN dffsnrnx1_pcell_0/m1_716_649# 2.04fF
C7 dffsnrnx1_pcell_1/m1_716_649# SN 3.98fF
C8 dffsnrnx1_pcell_2/m1_1660_723# dffsnrnx1_pcell_2/m1_716_649# 3.19fF
C9 SN dffsnrnx1_pcell_2/m1_716_649# 3.98fF
C10 dffsnrnx1_pcell_1/m1_1660_723# D 4.46fF
C11 SN CLK 2.43fF
C12 dffsnrnx1_pcell_0/m1_716_649# dffsnrnx1_pcell_0/m1_1660_723# 3.19fF
C13 m1_4715_501# m1_10453_649# 5.26fF
C14 VDD RN 2.54fF
C15 CLK RN 2.23fF
C16 SN D 2.38fF
C17 VDD CLK 7.04fF
C18 SN m1_4715_501# 4.68fF
C19 D dffsnrnx1_pcell_0/m1_1660_723# 4.47fF
C20 D RN 2.05fF
C21 D VDD 5.91fF
C22 dffsnrnx1_pcell_2/m1_1660_723# m1_10453_649# 4.46fF
C23 D CLK 11.68fF
C24 SN m1_10453_649# 2.65fF
C25 VDD m1_4715_501# 7.21fF
C26 CLK m1_4715_501# 11.67fF
C27 VDD GND 3.87fF
.ends
