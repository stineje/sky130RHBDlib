// File: FA.spi.FA.pxi
// Created: Tue Oct 15 15:48:52 2024
// 
simulator lang=spectre
x_PM_FA\%GND ( GND N_GND_c_16_p N_GND_c_71_p N_GND_c_79_p N_GND_c_435_p \
 N_GND_c_95_p N_GND_c_82_p N_GND_c_22_p N_GND_c_23_p N_GND_c_24_p N_GND_c_25_p \
 N_GND_c_453_p N_GND_c_26_p N_GND_c_27_p N_GND_c_28_p N_GND_c_29_p \
 N_GND_c_30_p N_GND_c_188_p N_GND_c_477_p N_GND_c_31_p N_GND_c_32_p \
 N_GND_c_33_p N_GND_c_34_p N_GND_c_35_p N_GND_c_36_p N_GND_c_495_p \
 N_GND_c_37_p N_GND_c_38_p N_GND_c_520_p N_GND_c_39_p N_GND_c_40_p \
 N_GND_c_41_p N_GND_c_42_p N_GND_c_517_p N_GND_c_43_p N_GND_c_297_p \
 N_GND_c_543_p N_GND_c_44_p N_GND_c_45_p N_GND_c_46_p N_GND_c_331_p \
 N_GND_c_540_p N_GND_c_311_p N_GND_c_319_p N_GND_c_333_p N_GND_c_334_p \
 N_GND_c_335_p N_GND_c_352_p N_GND_c_367_p N_GND_c_371_p N_GND_c_379_p \
 N_GND_c_380_p N_GND_c_381_p N_GND_c_405_p N_GND_c_1_p N_GND_c_2_p N_GND_c_3_p \
 N_GND_c_4_p N_GND_c_5_p N_GND_c_6_p N_GND_c_7_p N_GND_c_8_p N_GND_c_9_p \
 N_GND_c_10_p N_GND_c_11_p N_GND_c_12_p N_GND_c_13_p N_GND_c_14_p N_GND_c_15_p \
 N_GND_M0_noxref_s N_GND_M1_noxref_d N_GND_M3_noxref_d N_GND_M5_noxref_s \
 N_GND_M6_noxref_s N_GND_M7_noxref_d N_GND_M9_noxref_d N_GND_M11_noxref_s \
 N_GND_M12_noxref_d N_GND_M14_noxref_s N_GND_M15_noxref_d N_GND_M17_noxref_s \
 N_GND_M18_noxref_s N_GND_M20_noxref_s )  PM_FA\%GND
x_PM_FA\%VDD ( VDD N_VDD_c_573_p N_VDD_c_574_p N_VDD_c_575_p N_VDD_c_576_p \
 N_VDD_c_599_p N_VDD_c_629_p N_VDD_c_619_p N_VDD_c_651_p N_VDD_c_639_p \
 N_VDD_c_659_p N_VDD_c_660_p N_VDD_c_661_p N_VDD_c_662_p N_VDD_c_663_p \
 N_VDD_c_664_p N_VDD_c_665_p N_VDD_c_666_p N_VDD_c_667_p N_VDD_c_668_p \
 N_VDD_c_669_p N_VDD_c_670_p N_VDD_c_671_p N_VDD_c_759_p N_VDD_c_672_p \
 N_VDD_c_673_p N_VDD_c_674_p N_VDD_c_675_p N_VDD_c_676_p N_VDD_c_677_p \
 N_VDD_c_601_p N_VDD_c_905_p N_VDD_c_935_p N_VDD_c_938_p N_VDD_c_980_p \
 N_VDD_c_558_n N_VDD_c_559_n N_VDD_c_560_n N_VDD_c_561_n N_VDD_c_562_n \
 N_VDD_c_563_n N_VDD_c_564_n N_VDD_c_565_n N_VDD_c_566_n N_VDD_c_567_n \
 N_VDD_c_568_n N_VDD_c_569_n N_VDD_c_570_n N_VDD_c_571_n N_VDD_c_572_n \
 N_VDD_M21_noxref_s N_VDD_M22_noxref_d N_VDD_M23_noxref_d N_VDD_M27_noxref_d \
 N_VDD_M31_noxref_s N_VDD_M32_noxref_d N_VDD_M33_noxref_s N_VDD_M34_noxref_d \
 N_VDD_M35_noxref_d N_VDD_M39_noxref_d N_VDD_M43_noxref_s N_VDD_M44_noxref_d \
 N_VDD_M45_noxref_s N_VDD_M46_noxref_d N_VDD_M48_noxref_d N_VDD_M49_noxref_s \
 N_VDD_M50_noxref_d N_VDD_M51_noxref_s N_VDD_M52_noxref_d N_VDD_M54_noxref_d \
 N_VDD_M55_noxref_s N_VDD_M56_noxref_d N_VDD_M57_noxref_d N_VDD_M61_noxref_s \
 N_VDD_M62_noxref_d )  PM_FA\%VDD
x_PM_FA\%A ( N_A_c_1088_n N_A_c_1090_n N_A_c_1092_n N_A_c_1094_n N_A_c_1132_n \
 N_A_c_1134_n A A A A A A A A A A A A A A A A A A N_A_c_1142_n N_A_c_1260_p \
 N_A_M0_noxref_g N_A_M1_noxref_g N_A_M16_noxref_g N_A_M21_noxref_g \
 N_A_M22_noxref_g N_A_M23_noxref_g N_A_M24_noxref_g N_A_M53_noxref_g \
 N_A_M54_noxref_g N_A_c_1147_n N_A_c_1229_p N_A_c_1230_p N_A_c_1149_n \
 N_A_c_1199_n N_A_c_1200_n N_A_c_1150_n N_A_c_1212_p N_A_c_1151_n N_A_c_1153_n \
 N_A_c_1154_n N_A_c_1156_n N_A_c_1281_p N_A_c_1157_n N_A_c_1158_n N_A_c_1159_n \
 N_A_c_1160_n N_A_c_1162_n N_A_c_1295_p N_A_c_1297_p N_A_c_1298_p N_A_c_1380_p \
 N_A_c_1389_p N_A_c_1373_p N_A_c_1305_p N_A_c_1308_p N_A_c_1163_n N_A_c_1202_n \
 N_A_c_1274_p N_A_c_1382_p N_A_c_1261_p )  PM_FA\%A
x_PM_FA\%noxref_4 ( N_noxref_4_c_1465_n N_noxref_4_c_1471_n \
 N_noxref_4_c_1474_n N_noxref_4_c_1514_n N_noxref_4_c_1488_n \
 N_noxref_4_c_1491_n N_noxref_4_c_1477_n N_noxref_4_c_1480_n \
 N_noxref_4_M4_noxref_g N_noxref_4_M29_noxref_g N_noxref_4_M30_noxref_g \
 N_noxref_4_c_1552_p N_noxref_4_c_1554_p N_noxref_4_c_1555_p \
 N_noxref_4_c_1526_n N_noxref_4_c_1608_p N_noxref_4_c_1527_n \
 N_noxref_4_c_1561_p N_noxref_4_c_1564_p N_noxref_4_c_1569_p \
 N_noxref_4_M0_noxref_d N_noxref_4_M21_noxref_d )  PM_FA\%noxref_4
x_PM_FA\%noxref_5 ( N_noxref_5_c_1646_n N_noxref_5_c_1651_n \
 N_noxref_5_c_1670_n N_noxref_5_c_1689_n N_noxref_5_c_1652_n \
 N_noxref_5_c_1626_n N_noxref_5_c_1627_n N_noxref_5_c_1628_n \
 N_noxref_5_c_1629_n N_noxref_5_c_1656_n N_noxref_5_c_1657_n \
 N_noxref_5_M3_noxref_g N_noxref_5_M25_noxref_g N_noxref_5_M26_noxref_g \
 N_noxref_5_c_1632_n N_noxref_5_c_1634_n N_noxref_5_c_1635_n \
 N_noxref_5_c_1636_n N_noxref_5_c_1637_n N_noxref_5_c_1638_n \
 N_noxref_5_c_1639_n N_noxref_5_c_1641_n N_noxref_5_c_1681_n \
 N_noxref_5_M5_noxref_d N_noxref_5_M31_noxref_d )  PM_FA\%noxref_5
x_PM_FA\%B ( N_B_c_1801_n N_B_c_1910_n N_B_c_1830_n N_B_c_1837_n N_B_c_1839_n \
 N_B_c_1876_n N_B_c_1880_n B B B B B B B B B B B B B B B N_B_c_1803_n \
 N_B_c_1805_n N_B_c_1810_n N_B_M2_noxref_g N_B_M5_noxref_g N_B_M15_noxref_g \
 N_B_M27_noxref_g N_B_M28_noxref_g N_B_M31_noxref_g N_B_M32_noxref_g \
 N_B_M51_noxref_g N_B_M52_noxref_g N_B_c_1931_n N_B_c_1934_n N_B_c_1936_n \
 N_B_c_1939_n N_B_c_2077_p N_B_c_1943_n N_B_c_1944_n N_B_c_1945_n N_B_c_1811_n \
 N_B_c_1813_n N_B_c_2011_n N_B_c_1904_n N_B_c_1814_n N_B_c_2015_n N_B_c_1905_n \
 N_B_c_1815_n N_B_c_2019_n N_B_c_2020_n N_B_c_1817_n N_B_c_1818_n N_B_c_1820_n \
 N_B_c_1950_n N_B_c_1821_n N_B_c_1822_n N_B_c_1823_n N_B_c_1824_n N_B_c_1826_n \
 N_B_c_1907_n N_B_c_1827_n N_B_c_1908_n )  PM_FA\%B
x_PM_FA\%noxref_7 ( N_noxref_7_c_2293_n N_noxref_7_c_2272_n \
 N_noxref_7_c_2182_n N_noxref_7_c_2297_n N_noxref_7_c_2183_n \
 N_noxref_7_c_2187_n N_noxref_7_c_2188_n N_noxref_7_c_2230_n \
 N_noxref_7_c_2231_n N_noxref_7_c_2233_n N_noxref_7_c_2189_n \
 N_noxref_7_c_2277_n N_noxref_7_c_2190_n N_noxref_7_c_2236_n \
 N_noxref_7_c_2238_n N_noxref_7_c_2191_n N_noxref_7_c_2281_n \
 N_noxref_7_c_2239_n N_noxref_7_c_2193_n N_noxref_7_c_2198_n \
 N_noxref_7_c_2392_n N_noxref_7_c_2199_n N_noxref_7_M6_noxref_g \
 N_noxref_7_M7_noxref_g N_noxref_7_M13_noxref_g N_noxref_7_M33_noxref_g \
 N_noxref_7_M34_noxref_g N_noxref_7_M35_noxref_g N_noxref_7_M36_noxref_g \
 N_noxref_7_M47_noxref_g N_noxref_7_M48_noxref_g N_noxref_7_c_2201_n \
 N_noxref_7_c_2441_p N_noxref_7_c_2442_p N_noxref_7_c_2203_n \
 N_noxref_7_c_2263_n N_noxref_7_c_2264_n N_noxref_7_c_2204_n \
 N_noxref_7_c_2287_n N_noxref_7_c_2205_n N_noxref_7_c_2207_n \
 N_noxref_7_c_2208_n N_noxref_7_c_2210_n N_noxref_7_c_2496_p \
 N_noxref_7_c_2211_n N_noxref_7_c_2212_n N_noxref_7_c_2213_n \
 N_noxref_7_c_2214_n N_noxref_7_c_2216_n N_noxref_7_c_2506_p \
 N_noxref_7_c_2508_p N_noxref_7_c_2509_p N_noxref_7_c_2402_n \
 N_noxref_7_c_2541_p N_noxref_7_c_2289_n N_noxref_7_c_2515_p \
 N_noxref_7_c_2518_p N_noxref_7_c_2217_n N_noxref_7_c_2266_n \
 N_noxref_7_c_2291_n N_noxref_7_c_2292_n N_noxref_7_c_2405_n \
 N_noxref_7_M2_noxref_d N_noxref_7_M4_noxref_d N_noxref_7_M25_noxref_d \
 N_noxref_7_M29_noxref_d )  PM_FA\%noxref_7
x_PM_FA\%noxref_8 ( N_noxref_8_c_2602_n N_noxref_8_c_2604_n \
 N_noxref_8_c_2605_n N_noxref_8_c_2658_n N_noxref_8_c_2617_n \
 N_noxref_8_c_2619_n N_noxref_8_c_2607_n N_noxref_8_c_2610_n \
 N_noxref_8_M10_noxref_g N_noxref_8_M41_noxref_g N_noxref_8_M42_noxref_g \
 N_noxref_8_c_2708_p N_noxref_8_c_2709_p N_noxref_8_c_2710_p \
 N_noxref_8_c_2636_n N_noxref_8_c_2712_p N_noxref_8_c_2637_n \
 N_noxref_8_c_2714_p N_noxref_8_c_2705_p N_noxref_8_c_2647_n \
 N_noxref_8_M6_noxref_d N_noxref_8_M33_noxref_d )  PM_FA\%noxref_8
x_PM_FA\%SUM ( N_SUM_c_2794_n N_SUM_c_2795_n SUM SUM SUM SUM SUM \
 N_SUM_c_2779_n N_SUM_c_2781_n N_SUM_c_2765_n N_SUM_c_2792_n N_SUM_c_2782_n \
 N_SUM_c_2784_n N_SUM_c_2766_n N_SUM_c_2793_n N_SUM_M8_noxref_d \
 N_SUM_M10_noxref_d N_SUM_M37_noxref_d N_SUM_M41_noxref_d )  PM_FA\%SUM
x_PM_FA\%noxref_10 ( N_noxref_10_c_2933_n N_noxref_10_c_2955_n \
 N_noxref_10_c_2964_n N_noxref_10_c_2984_n N_noxref_10_c_2935_n \
 N_noxref_10_c_2913_n N_noxref_10_c_2914_n N_noxref_10_c_2915_n \
 N_noxref_10_c_2916_n N_noxref_10_c_2939_n N_noxref_10_c_2940_n \
 N_noxref_10_M9_noxref_g N_noxref_10_M37_noxref_g N_noxref_10_M38_noxref_g \
 N_noxref_10_c_2919_n N_noxref_10_c_2921_n N_noxref_10_c_2922_n \
 N_noxref_10_c_2923_n N_noxref_10_c_2924_n N_noxref_10_c_2925_n \
 N_noxref_10_c_2926_n N_noxref_10_c_2928_n N_noxref_10_c_2960_n \
 N_noxref_10_M11_noxref_d N_noxref_10_M43_noxref_d )  PM_FA\%noxref_10
x_PM_FA\%CIN ( N_CIN_c_3085_n N_CIN_c_3175_n N_CIN_c_3115_n N_CIN_c_3116_n \
 N_CIN_c_3087_n N_CIN_c_3118_n CIN CIN CIN CIN CIN CIN CIN CIN CIN CIN CIN CIN \
 CIN CIN N_CIN_c_3088_n N_CIN_c_3090_n N_CIN_c_3095_n N_CIN_M8_noxref_g \
 N_CIN_M11_noxref_g N_CIN_M12_noxref_g N_CIN_M39_noxref_g N_CIN_M40_noxref_g \
 N_CIN_M43_noxref_g N_CIN_M44_noxref_g N_CIN_M45_noxref_g N_CIN_M46_noxref_g \
 N_CIN_c_3193_n N_CIN_c_3196_n N_CIN_c_3198_n N_CIN_c_3150_n N_CIN_c_3257_n \
 N_CIN_c_3151_n N_CIN_c_3204_n N_CIN_c_3205_n N_CIN_c_3096_n N_CIN_c_3098_n \
 N_CIN_c_3294_n N_CIN_c_3140_n N_CIN_c_3099_n N_CIN_c_3298_n N_CIN_c_3141_n \
 N_CIN_c_3100_n N_CIN_c_3302_n N_CIN_c_3303_n N_CIN_c_3102_n N_CIN_c_3103_n \
 N_CIN_c_3105_n N_CIN_c_3208_n N_CIN_c_3106_n N_CIN_c_3107_n N_CIN_c_3108_n \
 N_CIN_c_3109_n N_CIN_c_3111_n N_CIN_c_3143_n N_CIN_c_3112_n N_CIN_c_3144_n )  \
 PM_FA\%CIN
x_PM_FA\%noxref_12 ( N_noxref_12_c_3336_n N_noxref_12_c_3394_n \
 N_noxref_12_c_3359_n N_noxref_12_c_3363_n N_noxref_12_c_3365_n \
 N_noxref_12_c_3337_n N_noxref_12_c_3395_n N_noxref_12_c_3368_n \
 N_noxref_12_c_3339_n N_noxref_12_c_3426_n N_noxref_12_M14_noxref_g \
 N_noxref_12_M49_noxref_g N_noxref_12_M50_noxref_g N_noxref_12_c_3344_n \
 N_noxref_12_c_3457_p N_noxref_12_c_3458_p N_noxref_12_c_3346_n \
 N_noxref_12_c_3379_n N_noxref_12_c_3380_n N_noxref_12_c_3347_n \
 N_noxref_12_c_3399_n N_noxref_12_c_3348_n N_noxref_12_c_3350_n \
 N_noxref_12_c_3351_n N_noxref_12_M13_noxref_d N_noxref_12_M45_noxref_d \
 N_noxref_12_M47_noxref_d )  PM_FA\%noxref_12
x_PM_FA\%noxref_13 ( N_noxref_13_c_3497_n N_noxref_13_c_3500_n \
 N_noxref_13_c_3502_n N_noxref_13_c_3506_n N_noxref_13_c_3508_n \
 N_noxref_13_c_3475_n N_noxref_13_c_3579_p N_noxref_13_c_3477_n \
 N_noxref_13_c_3478_n N_noxref_13_c_3554_n N_noxref_13_M17_noxref_g \
 N_noxref_13_M55_noxref_g N_noxref_13_M56_noxref_g N_noxref_13_c_3483_n \
 N_noxref_13_c_3598_p N_noxref_13_c_3599_p N_noxref_13_c_3485_n \
 N_noxref_13_c_3522_n N_noxref_13_c_3523_n N_noxref_13_c_3486_n \
 N_noxref_13_c_3586_p N_noxref_13_c_3487_n N_noxref_13_c_3489_n \
 N_noxref_13_c_3490_n N_noxref_13_M16_noxref_d N_noxref_13_M51_noxref_d \
 N_noxref_13_M53_noxref_d )  PM_FA\%noxref_13
x_PM_FA\%noxref_14 ( N_noxref_14_c_3617_n N_noxref_14_c_3675_n \
 N_noxref_14_c_3629_n N_noxref_14_c_3693_n N_noxref_14_c_3650_n \
 N_noxref_14_c_3652_n N_noxref_14_c_3631_n N_noxref_14_c_3632_n \
 N_noxref_14_c_3656_n N_noxref_14_M18_noxref_g N_noxref_14_M57_noxref_g \
 N_noxref_14_M58_noxref_g N_noxref_14_c_3635_n N_noxref_14_c_3744_p \
 N_noxref_14_c_3745_p N_noxref_14_c_3637_n N_noxref_14_c_3639_n \
 N_noxref_14_c_3768_p N_noxref_14_c_3734_p N_noxref_14_c_3640_n \
 N_noxref_14_c_3642_n N_noxref_14_c_3664_n N_noxref_14_M14_noxref_d \
 N_noxref_14_M49_noxref_d )  PM_FA\%noxref_14
x_PM_FA\%noxref_15 ( N_noxref_15_c_3782_n N_noxref_15_c_3803_n \
 N_noxref_15_c_3783_n N_noxref_15_c_3824_n N_noxref_15_c_3805_n \
 N_noxref_15_c_3808_n N_noxref_15_c_3786_n N_noxref_15_c_3856_n \
 N_noxref_15_c_3787_n N_noxref_15_M19_noxref_g N_noxref_15_M59_noxref_g \
 N_noxref_15_M60_noxref_g N_noxref_15_c_3789_n N_noxref_15_c_3867_n \
 N_noxref_15_c_3870_n N_noxref_15_c_3891_p N_noxref_15_c_3791_n \
 N_noxref_15_c_3792_n N_noxref_15_c_3793_n N_noxref_15_c_3874_n \
 N_noxref_15_c_3875_n N_noxref_15_c_3877_n N_noxref_15_c_3878_n \
 N_noxref_15_M17_noxref_d N_noxref_15_M55_noxref_d )  PM_FA\%noxref_15
x_PM_FA\%noxref_16 ( N_noxref_16_c_3919_n N_noxref_16_c_3925_n \
 N_noxref_16_c_3927_n N_noxref_16_c_3986_n N_noxref_16_c_3964_n \
 N_noxref_16_c_3966_n N_noxref_16_c_3931_n N_noxref_16_c_3936_n \
 N_noxref_16_c_3937_n N_noxref_16_M20_noxref_g N_noxref_16_M61_noxref_g \
 N_noxref_16_M62_noxref_g N_noxref_16_c_3942_n N_noxref_16_c_4047_p \
 N_noxref_16_c_4048_p N_noxref_16_c_3944_n N_noxref_16_c_3978_n \
 N_noxref_16_c_3979_n N_noxref_16_c_3945_n N_noxref_16_c_4039_p \
 N_noxref_16_c_3946_n N_noxref_16_c_3948_n N_noxref_16_c_3949_n \
 N_noxref_16_M18_noxref_d N_noxref_16_M19_noxref_d N_noxref_16_M59_noxref_d )  \
 PM_FA\%noxref_16
x_PM_FA\%noxref_17 ( N_noxref_17_c_4059_n N_noxref_17_c_4064_n \
 N_noxref_17_c_4066_n N_noxref_17_c_4067_n N_noxref_17_M23_noxref_s \
 N_noxref_17_M24_noxref_d N_noxref_17_M26_noxref_d )  PM_FA\%noxref_17
x_PM_FA\%noxref_18 ( N_noxref_18_c_4098_n N_noxref_18_c_4099_n \
 N_noxref_18_c_4103_n N_noxref_18_c_4106_n N_noxref_18_c_4107_n \
 N_noxref_18_c_4110_n N_noxref_18_M1_noxref_s )  PM_FA\%noxref_18
x_PM_FA\%noxref_19 ( N_noxref_19_c_4149_n N_noxref_19_c_4154_n \
 N_noxref_19_c_4155_n N_noxref_19_c_4156_n N_noxref_19_M27_noxref_s \
 N_noxref_19_M28_noxref_d N_noxref_19_M30_noxref_d )  PM_FA\%noxref_19
x_PM_FA\%noxref_20 ( N_noxref_20_c_4211_n N_noxref_20_c_4190_n \
 N_noxref_20_c_4194_n N_noxref_20_c_4197_n N_noxref_20_c_4198_n \
 N_noxref_20_c_4201_n N_noxref_20_M3_noxref_s )  PM_FA\%noxref_20
x_PM_FA\%noxref_21 ( N_noxref_21_c_4240_n N_noxref_21_c_4245_n \
 N_noxref_21_c_4247_n N_noxref_21_c_4248_n N_noxref_21_M35_noxref_s \
 N_noxref_21_M36_noxref_d N_noxref_21_M38_noxref_d )  PM_FA\%noxref_21
x_PM_FA\%noxref_22 ( N_noxref_22_c_4277_n N_noxref_22_c_4278_n \
 N_noxref_22_c_4282_n N_noxref_22_c_4285_n N_noxref_22_c_4286_n \
 N_noxref_22_c_4289_n N_noxref_22_M7_noxref_s )  PM_FA\%noxref_22
x_PM_FA\%noxref_23 ( N_noxref_23_c_4326_n N_noxref_23_c_4331_n \
 N_noxref_23_c_4332_n N_noxref_23_c_4333_n N_noxref_23_M39_noxref_s \
 N_noxref_23_M40_noxref_d N_noxref_23_M42_noxref_d )  PM_FA\%noxref_23
x_PM_FA\%noxref_24 ( N_noxref_24_c_4386_n N_noxref_24_c_4365_n \
 N_noxref_24_c_4369_n N_noxref_24_c_4372_n N_noxref_24_c_4373_n \
 N_noxref_24_c_4376_n N_noxref_24_M9_noxref_s )  PM_FA\%noxref_24
x_PM_FA\%noxref_25 ( N_noxref_25_c_4415_n N_noxref_25_c_4416_n \
 N_noxref_25_c_4420_n N_noxref_25_c_4423_n N_noxref_25_c_4424_n \
 N_noxref_25_c_4427_n N_noxref_25_M12_noxref_s )  PM_FA\%noxref_25
x_PM_FA\%noxref_26 ( N_noxref_26_c_4468_n N_noxref_26_c_4469_n \
 N_noxref_26_c_4473_n N_noxref_26_c_4476_n N_noxref_26_c_4477_n \
 N_noxref_26_c_4480_n N_noxref_26_M15_noxref_s )  PM_FA\%noxref_26
x_PM_FA\%noxref_27 ( N_noxref_27_c_4525_n N_noxref_27_c_4530_n \
 N_noxref_27_c_4532_n N_noxref_27_c_4533_n N_noxref_27_M57_noxref_s \
 N_noxref_27_M58_noxref_d N_noxref_27_M60_noxref_d )  PM_FA\%noxref_27
x_PM_FA\%COUT ( COUT COUT COUT COUT COUT COUT COUT N_COUT_c_4568_n \
 N_COUT_c_4592_n N_COUT_c_4578_n N_COUT_c_4581_n N_COUT_M20_noxref_d \
 N_COUT_M61_noxref_d )  PM_FA\%COUT
cc_1 ( N_GND_c_1_p N_VDD_c_558_n ) capacitor c=0.00989031f //x=38.48 //y=0 \
 //x2=38.48 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_559_n ) capacitor c=0.00989031f //x=0.63 //y=0 \
 //x2=0.74 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_560_n ) capacitor c=0.00582097f //x=2.22 //y=0 \
 //x2=2.22 //y2=7.4
cc_4 ( N_GND_c_4_p N_VDD_c_561_n ) capacitor c=0.0057235f //x=5.55 //y=0 \
 //x2=5.55 //y2=7.4
cc_5 ( N_GND_c_5_p N_VDD_c_562_n ) capacitor c=0.00474727f //x=8.88 //y=0 \
 //x2=8.88 //y2=7.4
cc_6 ( N_GND_c_6_p N_VDD_c_563_n ) capacitor c=0.0085201f //x=11.1 //y=0 \
 //x2=11.1 //y2=7.4
cc_7 ( N_GND_c_7_p N_VDD_c_564_n ) capacitor c=0.00582097f //x=13.32 //y=0 \
 //x2=13.32 //y2=7.4
cc_8 ( N_GND_c_8_p N_VDD_c_565_n ) capacitor c=0.0057235f //x=16.65 //y=0 \
 //x2=16.65 //y2=7.4
cc_9 ( N_GND_c_9_p N_VDD_c_566_n ) capacitor c=0.00478842f //x=19.98 //y=0 \
 //x2=19.98 //y2=7.4
cc_10 ( N_GND_c_10_p N_VDD_c_567_n ) capacitor c=0.00969007f //x=22.2 //y=0 \
 //x2=22.2 //y2=7.4
cc_11 ( N_GND_c_11_p N_VDD_c_568_n ) capacitor c=0.00855708f //x=25.53 //y=0 \
 //x2=25.53 //y2=7.4
cc_12 ( N_GND_c_12_p N_VDD_c_569_n ) capacitor c=0.00850989f //x=27.75 //y=0 \
 //x2=27.75 //y2=7.4
cc_13 ( N_GND_c_13_p N_VDD_c_570_n ) capacitor c=0.00829849f //x=31.08 //y=0 \
 //x2=31.08 //y2=7.4
cc_14 ( N_GND_c_14_p N_VDD_c_571_n ) capacitor c=0.00829849f //x=33.3 //y=0 \
 //x2=33.3 //y2=7.4
cc_15 ( N_GND_c_15_p N_VDD_c_572_n ) capacitor c=0.00855708f //x=36.63 //y=0 \
 //x2=36.63 //y2=7.4
cc_16 ( N_GND_c_16_p N_A_c_1088_n ) capacitor c=0.00375365f //x=38.48 //y=0 \
 //x2=3.215 //y2=4.07
cc_17 ( N_GND_c_3_p N_A_c_1088_n ) capacitor c=0.00249386f //x=2.22 //y=0 \
 //x2=3.215 //y2=4.07
cc_18 ( N_GND_c_16_p N_A_c_1090_n ) capacitor c=0.00155455f //x=38.48 //y=0 \
 //x2=0.855 //y2=4.07
cc_19 ( N_GND_M0_noxref_s N_A_c_1090_n ) capacitor c=5.91312e-19 //x=0.495 \
 //y=0.37 //x2=0.855 //y2=4.07
cc_20 ( N_GND_c_16_p N_A_c_1092_n ) capacitor c=2.19685e-19 //x=38.48 //y=0 \
 //x2=3.33 //y2=2.105
cc_21 ( N_GND_c_3_p N_A_c_1092_n ) capacitor c=0.00219549f //x=2.22 //y=0 \
 //x2=3.33 //y2=2.105
cc_22 ( N_GND_c_22_p N_A_c_1094_n ) capacitor c=0.00586301f //x=5.38 //y=0 \
 //x2=29.515 //y2=1.85
cc_23 ( N_GND_c_23_p N_A_c_1094_n ) capacitor c=0.00449081f //x=6.645 //y=0 \
 //x2=29.515 //y2=1.85
cc_24 ( N_GND_c_24_p N_A_c_1094_n ) capacitor c=0.00586301f //x=8.71 //y=0 \
 //x2=29.515 //y2=1.85
cc_25 ( N_GND_c_25_p N_A_c_1094_n ) capacitor c=0.00249862f //x=9.415 //y=0 \
 //x2=29.515 //y2=1.85
cc_26 ( N_GND_c_26_p N_A_c_1094_n ) capacitor c=0.00231363f //x=9.9 //y=0.535 \
 //x2=29.515 //y2=1.85
cc_27 ( N_GND_c_27_p N_A_c_1094_n ) capacitor c=0.00421577f //x=10.385 \
 //y=0.535 //x2=29.515 //y2=1.85
cc_28 ( N_GND_c_28_p N_A_c_1094_n ) capacitor c=0.00259291f //x=10.93 //y=0 \
 //x2=29.515 //y2=1.85
cc_29 ( N_GND_c_29_p N_A_c_1094_n ) capacitor c=0.00259291f //x=11.645 //y=0 \
 //x2=29.515 //y2=1.85
cc_30 ( N_GND_c_30_p N_A_c_1094_n ) capacitor c=0.00486004f //x=12.13 \
 //y=0.535 //x2=29.515 //y2=1.85
cc_31 ( N_GND_c_31_p N_A_c_1094_n ) capacitor c=0.00249862f //x=13.15 //y=0 \
 //x2=29.515 //y2=1.85
cc_32 ( N_GND_c_32_p N_A_c_1094_n ) capacitor c=0.00449081f //x=14.415 //y=0 \
 //x2=29.515 //y2=1.85
cc_33 ( N_GND_c_33_p N_A_c_1094_n ) capacitor c=0.00586301f //x=16.48 //y=0 \
 //x2=29.515 //y2=1.85
cc_34 ( N_GND_c_34_p N_A_c_1094_n ) capacitor c=0.00449081f //x=17.745 //y=0 \
 //x2=29.515 //y2=1.85
cc_35 ( N_GND_c_35_p N_A_c_1094_n ) capacitor c=0.00586301f //x=19.81 //y=0 \
 //x2=29.515 //y2=1.85
cc_36 ( N_GND_c_36_p N_A_c_1094_n ) capacitor c=0.00249862f //x=20.515 //y=0 \
 //x2=29.515 //y2=1.85
cc_37 ( N_GND_c_37_p N_A_c_1094_n ) capacitor c=0.00231363f //x=21 //y=0.535 \
 //x2=29.515 //y2=1.85
cc_38 ( N_GND_c_38_p N_A_c_1094_n ) capacitor c=0.00421577f //x=21.485 \
 //y=0.535 //x2=29.515 //y2=1.85
cc_39 ( N_GND_c_39_p N_A_c_1094_n ) capacitor c=0.00259291f //x=22.03 //y=0 \
 //x2=29.515 //y2=1.85
cc_40 ( N_GND_c_40_p N_A_c_1094_n ) capacitor c=0.00448875f //x=23.295 //y=0 \
 //x2=29.515 //y2=1.85
cc_41 ( N_GND_c_41_p N_A_c_1094_n ) capacitor c=0.00576163f //x=25.36 //y=0 \
 //x2=29.515 //y2=1.85
cc_42 ( N_GND_c_42_p N_A_c_1094_n ) capacitor c=0.00259291f //x=26.075 //y=0 \
 //x2=29.515 //y2=1.85
cc_43 ( N_GND_c_43_p N_A_c_1094_n ) capacitor c=0.00465172f //x=26.56 \
 //y=0.535 //x2=29.515 //y2=1.85
cc_44 ( N_GND_c_44_p N_A_c_1094_n ) capacitor c=0.00249862f //x=27.58 //y=0 \
 //x2=29.515 //y2=1.85
cc_45 ( N_GND_c_45_p N_A_c_1094_n ) capacitor c=0.00448875f //x=28.845 //y=0 \
 //x2=29.515 //y2=1.85
cc_46 ( N_GND_c_46_p N_A_c_1094_n ) capacitor c=0.00117121f //x=30.91 //y=0 \
 //x2=29.515 //y2=1.85
cc_47 ( N_GND_c_4_p N_A_c_1094_n ) capacitor c=0.0427295f //x=5.55 //y=0 \
 //x2=29.515 //y2=1.85
cc_48 ( N_GND_c_5_p N_A_c_1094_n ) capacitor c=0.0428613f //x=8.88 //y=0 \
 //x2=29.515 //y2=1.85
cc_49 ( N_GND_c_6_p N_A_c_1094_n ) capacitor c=0.0459641f //x=11.1 //y=0 \
 //x2=29.515 //y2=1.85
cc_50 ( N_GND_c_7_p N_A_c_1094_n ) capacitor c=0.0392964f //x=13.32 //y=0 \
 //x2=29.515 //y2=1.85
cc_51 ( N_GND_c_8_p N_A_c_1094_n ) capacitor c=0.0380496f //x=16.65 //y=0 \
 //x2=29.515 //y2=1.85
cc_52 ( N_GND_c_9_p N_A_c_1094_n ) capacitor c=0.0370781f //x=19.98 //y=0 \
 //x2=29.515 //y2=1.85
cc_53 ( N_GND_c_10_p N_A_c_1094_n ) capacitor c=0.0391552f //x=22.2 //y=0 \
 //x2=29.515 //y2=1.85
cc_54 ( N_GND_c_11_p N_A_c_1094_n ) capacitor c=0.0439804f //x=25.53 //y=0 \
 //x2=29.515 //y2=1.85
cc_55 ( N_GND_c_12_p N_A_c_1094_n ) capacitor c=0.0447716f //x=27.75 //y=0 \
 //x2=29.515 //y2=1.85
cc_56 ( N_GND_M5_noxref_s N_A_c_1094_n ) capacitor c=0.0183637f //x=9.375 \
 //y=0.37 //x2=29.515 //y2=1.85
cc_57 ( N_GND_M6_noxref_s N_A_c_1094_n ) capacitor c=0.0200331f //x=11.595 \
 //y=0.37 //x2=29.515 //y2=1.85
cc_58 ( N_GND_M11_noxref_s N_A_c_1094_n ) capacitor c=0.0183637f //x=20.475 \
 //y=0.37 //x2=29.515 //y2=1.85
cc_59 ( N_GND_M14_noxref_s N_A_c_1094_n ) capacitor c=0.0200331f //x=26.025 \
 //y=0.37 //x2=29.515 //y2=1.85
cc_60 ( N_GND_c_16_p N_A_c_1132_n ) capacitor c=0.327127f //x=38.48 //y=0 \
 //x2=3.415 //y2=1.85
cc_61 ( N_GND_c_3_p N_A_c_1132_n ) capacitor c=0.00642784f //x=2.22 //y=0 \
 //x2=3.415 //y2=1.85
cc_62 ( N_GND_c_16_p N_A_c_1134_n ) capacitor c=2.30154e-19 //x=38.48 //y=0 \
 //x2=29.6 //y2=2.105
cc_63 ( N_GND_c_3_p A ) capacitor c=0.00676236f //x=2.22 //y=0 //x2=3.33 \
 //y2=2.96
cc_64 ( N_GND_c_12_p A ) capacitor c=4.34469e-19 //x=27.75 //y=0 //x2=29.6 \
 //y2=2.59
cc_65 ( N_GND_c_13_p A ) capacitor c=6.38128e-19 //x=31.08 //y=0 //x2=29.6 \
 //y2=2.59
cc_66 ( N_GND_c_3_p A ) capacitor c=0.00822147f //x=2.22 //y=0 //x2=3.33 \
 //y2=2.22
cc_67 ( N_GND_M1_noxref_d A ) capacitor c=2.10573e-19 //x=3.21 //y=0.87 \
 //x2=3.33 //y2=2.22
cc_68 ( N_GND_c_12_p A ) capacitor c=3.61829e-19 //x=27.75 //y=0 //x2=29.6 \
 //y2=2.22
cc_69 ( N_GND_c_13_p A ) capacitor c=5.01476e-19 //x=31.08 //y=0 //x2=29.6 \
 //y2=2.22
cc_70 ( N_GND_c_16_p N_A_c_1142_n ) capacitor c=0.00187124f //x=38.48 //y=0 \
 //x2=0.74 //y2=2.085
cc_71 ( N_GND_c_71_p N_A_c_1142_n ) capacitor c=8.01092e-19 //x=1.03 //y=0.535 \
 //x2=0.74 //y2=2.085
cc_72 ( N_GND_c_2_p N_A_c_1142_n ) capacitor c=0.0285526f //x=0.63 //y=0 \
 //x2=0.74 //y2=2.085
cc_73 ( N_GND_c_3_p N_A_c_1142_n ) capacitor c=0.00143388f //x=2.22 //y=0 \
 //x2=0.74 //y2=2.085
cc_74 ( N_GND_M0_noxref_s N_A_c_1142_n ) capacitor c=0.0110965f //x=0.495 \
 //y=0.37 //x2=0.74 //y2=2.085
cc_75 ( N_GND_c_71_p N_A_c_1147_n ) capacitor c=0.0120496f //x=1.03 //y=0.535 \
 //x2=0.85 //y2=0.91
cc_76 ( N_GND_M0_noxref_s N_A_c_1147_n ) capacitor c=0.0316686f //x=0.495 \
 //y=0.37 //x2=0.85 //y2=0.91
cc_77 ( N_GND_c_2_p N_A_c_1149_n ) capacitor c=0.0114366f //x=0.63 //y=0 \
 //x2=0.85 //y2=1.92
cc_78 ( N_GND_M0_noxref_s N_A_c_1150_n ) capacitor c=0.00483274f //x=0.495 \
 //y=0.37 //x2=1.225 //y2=0.755
cc_79 ( N_GND_c_79_p N_A_c_1151_n ) capacitor c=0.0118602f //x=1.515 //y=0.535 \
 //x2=1.38 //y2=0.91
cc_80 ( N_GND_M0_noxref_s N_A_c_1151_n ) capacitor c=0.0143355f //x=0.495 \
 //y=0.37 //x2=1.38 //y2=0.91
cc_81 ( N_GND_M0_noxref_s N_A_c_1153_n ) capacitor c=0.0074042f //x=0.495 \
 //y=0.37 //x2=1.38 //y2=1.255
cc_82 ( N_GND_c_82_p N_A_c_1154_n ) capacitor c=0.00134217f //x=3.315 //y=0 \
 //x2=3.135 //y2=0.87
cc_83 ( N_GND_M1_noxref_d N_A_c_1154_n ) capacitor c=0.00220047f //x=3.21 \
 //y=0.87 //x2=3.135 //y2=0.87
cc_84 ( N_GND_M1_noxref_d N_A_c_1156_n ) capacitor c=0.00255985f //x=3.21 \
 //y=0.87 //x2=3.135 //y2=1.215
cc_85 ( N_GND_c_3_p N_A_c_1157_n ) capacitor c=0.00733575f //x=2.22 //y=0 \
 //x2=3.135 //y2=1.92
cc_86 ( N_GND_M1_noxref_d N_A_c_1158_n ) capacitor c=0.013135f //x=3.21 \
 //y=0.87 //x2=3.51 //y2=0.715
cc_87 ( N_GND_M1_noxref_d N_A_c_1159_n ) capacitor c=0.00193136f //x=3.21 \
 //y=0.87 //x2=3.51 //y2=1.37
cc_88 ( N_GND_c_22_p N_A_c_1160_n ) capacitor c=0.00129817f //x=5.38 //y=0 \
 //x2=3.665 //y2=0.87
cc_89 ( N_GND_M1_noxref_d N_A_c_1160_n ) capacitor c=0.00257848f //x=3.21 \
 //y=0.87 //x2=3.665 //y2=0.87
cc_90 ( N_GND_M1_noxref_d N_A_c_1162_n ) capacitor c=0.00255985f //x=3.21 \
 //y=0.87 //x2=3.665 //y2=1.215
cc_91 ( N_GND_c_71_p N_A_c_1163_n ) capacitor c=2.1838e-19 //x=1.03 //y=0.535 \
 //x2=0.74 //y2=2.085
cc_92 ( N_GND_c_2_p N_A_c_1163_n ) capacitor c=0.00769211f //x=0.63 //y=0 \
 //x2=0.74 //y2=2.085
cc_93 ( N_GND_M0_noxref_s N_A_c_1163_n ) capacitor c=0.00655738f //x=0.495 \
 //y=0.37 //x2=0.74 //y2=2.085
cc_94 ( N_GND_c_16_p N_noxref_4_c_1465_n ) capacitor c=0.0225635f //x=38.48 \
 //y=0 //x2=7.655 //y2=2.59
cc_95 ( N_GND_c_95_p N_noxref_4_c_1465_n ) capacitor c=0.0015622f //x=2.05 \
 //y=0 //x2=7.655 //y2=2.59
cc_96 ( N_GND_c_82_p N_noxref_4_c_1465_n ) capacitor c=0.00277229f //x=3.315 \
 //y=0 //x2=7.655 //y2=2.59
cc_97 ( N_GND_c_3_p N_noxref_4_c_1465_n ) capacitor c=0.038878f //x=2.22 //y=0 \
 //x2=7.655 //y2=2.59
cc_98 ( N_GND_c_4_p N_noxref_4_c_1465_n ) capacitor c=0.0262396f //x=5.55 \
 //y=0 //x2=7.655 //y2=2.59
cc_99 ( N_GND_M0_noxref_s N_noxref_4_c_1465_n ) capacitor c=0.00248261f \
 //x=0.495 //y=0.37 //x2=7.655 //y2=2.59
cc_100 ( N_GND_c_16_p N_noxref_4_c_1471_n ) capacitor c=0.00231366f //x=38.48 \
 //y=0 //x2=1.595 //y2=2.59
cc_101 ( N_GND_c_3_p N_noxref_4_c_1471_n ) capacitor c=0.00209945f //x=2.22 \
 //y=0 //x2=1.595 //y2=2.59
cc_102 ( N_GND_M0_noxref_s N_noxref_4_c_1471_n ) capacitor c=0.00120637f \
 //x=0.495 //y=0.37 //x2=1.595 //y2=2.59
cc_103 ( N_GND_c_16_p N_noxref_4_c_1474_n ) capacitor c=0.00129718f //x=38.48 \
 //y=0 //x2=1.395 //y2=2.08
cc_104 ( N_GND_c_3_p N_noxref_4_c_1474_n ) capacitor c=0.0254284f //x=2.22 \
 //y=0 //x2=1.395 //y2=2.08
cc_105 ( N_GND_M0_noxref_s N_noxref_4_c_1474_n ) capacitor c=0.00949589f \
 //x=0.495 //y=0.37 //x2=1.395 //y2=2.08
cc_106 ( N_GND_c_2_p N_noxref_4_c_1477_n ) capacitor c=0.00113816f //x=0.63 \
 //y=0 //x2=1.48 //y2=2.59
cc_107 ( N_GND_c_3_p N_noxref_4_c_1477_n ) capacitor c=5.56859e-19 //x=2.22 \
 //y=0 //x2=1.48 //y2=2.59
cc_108 ( N_GND_M0_noxref_s N_noxref_4_c_1477_n ) capacitor c=2.30929e-19 \
 //x=0.495 //y=0.37 //x2=1.48 //y2=2.59
cc_109 ( N_GND_c_4_p N_noxref_4_c_1480_n ) capacitor c=6.69104e-19 //x=5.55 \
 //y=0 //x2=7.77 //y2=2.085
cc_110 ( N_GND_c_5_p N_noxref_4_c_1480_n ) capacitor c=0.00180575f //x=8.88 \
 //y=0 //x2=7.77 //y2=2.085
cc_111 ( N_GND_c_16_p N_noxref_4_M0_noxref_d ) capacitor c=0.00136354f \
 //x=38.48 //y=0 //x2=0.925 //y2=0.91
cc_112 ( N_GND_c_71_p N_noxref_4_M0_noxref_d ) capacitor c=0.0151737f //x=1.03 \
 //y=0.535 //x2=0.925 //y2=0.91
cc_113 ( N_GND_c_2_p N_noxref_4_M0_noxref_d ) capacitor c=0.00942176f //x=0.63 \
 //y=0 //x2=0.925 //y2=0.91
cc_114 ( N_GND_c_3_p N_noxref_4_M0_noxref_d ) capacitor c=0.00934943f //x=2.22 \
 //y=0 //x2=0.925 //y2=0.91
cc_115 ( N_GND_M0_noxref_s N_noxref_4_M0_noxref_d ) capacitor c=0.076995f \
 //x=0.495 //y=0.37 //x2=0.925 //y2=0.91
cc_116 ( N_GND_c_4_p N_noxref_5_c_1626_n ) capacitor c=0.0146874f //x=5.55 \
 //y=0 //x2=6.66 //y2=2.085
cc_117 ( N_GND_c_6_p N_noxref_5_c_1627_n ) capacitor c=0.00152332f //x=11.1 \
 //y=0 //x2=9.62 //y2=3.33
cc_118 ( N_GND_M5_noxref_s N_noxref_5_c_1628_n ) capacitor c=0.00157668f \
 //x=9.375 //y=0.37 //x2=9.905 //y2=2.08
cc_119 ( N_GND_c_26_p N_noxref_5_c_1629_n ) capacitor c=0.00157668f //x=9.9 \
 //y=0.535 //x2=9.705 //y2=2.08
cc_120 ( N_GND_c_5_p N_noxref_5_c_1629_n ) capacitor c=0.0288208f //x=8.88 \
 //y=0 //x2=9.705 //y2=2.08
cc_121 ( N_GND_M5_noxref_s N_noxref_5_c_1629_n ) capacitor c=0.00514876f \
 //x=9.375 //y=0.37 //x2=9.705 //y2=2.08
cc_122 ( N_GND_c_23_p N_noxref_5_c_1632_n ) capacitor c=0.00134217f //x=6.645 \
 //y=0 //x2=6.465 //y2=0.87
cc_123 ( N_GND_M3_noxref_d N_noxref_5_c_1632_n ) capacitor c=0.00220047f \
 //x=6.54 //y=0.87 //x2=6.465 //y2=0.87
cc_124 ( N_GND_M3_noxref_d N_noxref_5_c_1634_n ) capacitor c=0.00255985f \
 //x=6.54 //y=0.87 //x2=6.465 //y2=1.215
cc_125 ( N_GND_c_4_p N_noxref_5_c_1635_n ) capacitor c=0.00176175f //x=5.55 \
 //y=0 //x2=6.465 //y2=1.525
cc_126 ( N_GND_c_4_p N_noxref_5_c_1636_n ) capacitor c=0.00752966f //x=5.55 \
 //y=0 //x2=6.465 //y2=1.92
cc_127 ( N_GND_M3_noxref_d N_noxref_5_c_1637_n ) capacitor c=0.013135f \
 //x=6.54 //y=0.87 //x2=6.84 //y2=0.715
cc_128 ( N_GND_M3_noxref_d N_noxref_5_c_1638_n ) capacitor c=0.00193136f \
 //x=6.54 //y=0.87 //x2=6.84 //y2=1.37
cc_129 ( N_GND_c_24_p N_noxref_5_c_1639_n ) capacitor c=0.00129817f //x=8.71 \
 //y=0 //x2=6.995 //y2=0.87
cc_130 ( N_GND_M3_noxref_d N_noxref_5_c_1639_n ) capacitor c=0.00257848f \
 //x=6.54 //y=0.87 //x2=6.995 //y2=0.87
cc_131 ( N_GND_M3_noxref_d N_noxref_5_c_1641_n ) capacitor c=0.00255985f \
 //x=6.54 //y=0.87 //x2=6.995 //y2=1.215
cc_132 ( N_GND_c_16_p N_noxref_5_M5_noxref_d ) capacitor c=0.00108086f \
 //x=38.48 //y=0 //x2=9.795 //y2=0.91
cc_133 ( N_GND_c_5_p N_noxref_5_M5_noxref_d ) capacitor c=0.00686786f //x=8.88 \
 //y=0 //x2=9.795 //y2=0.91
cc_134 ( N_GND_c_6_p N_noxref_5_M5_noxref_d ) capacitor c=0.00737105f //x=11.1 \
 //y=0 //x2=9.795 //y2=0.91
cc_135 ( N_GND_M5_noxref_s N_noxref_5_M5_noxref_d ) capacitor c=0.0916952f \
 //x=9.375 //y=0.37 //x2=9.795 //y2=0.91
cc_136 ( N_GND_c_4_p N_B_c_1801_n ) capacitor c=0.00750857f //x=5.55 //y=0 \
 //x2=10.245 //y2=2.96
cc_137 ( N_GND_c_5_p N_B_c_1801_n ) capacitor c=0.0110081f //x=8.88 //y=0 \
 //x2=10.245 //y2=2.96
cc_138 ( N_GND_c_3_p N_B_c_1803_n ) capacitor c=5.75615e-19 //x=2.22 //y=0 \
 //x2=4.44 //y2=2.085
cc_139 ( N_GND_c_4_p N_B_c_1803_n ) capacitor c=0.00175406f //x=5.55 //y=0 \
 //x2=4.44 //y2=2.085
cc_140 ( N_GND_c_16_p N_B_c_1805_n ) capacitor c=0.00115109f //x=38.48 //y=0 \
 //x2=10.36 //y2=2.085
cc_141 ( N_GND_c_27_p N_B_c_1805_n ) capacitor c=4.37745e-19 //x=10.385 \
 //y=0.535 //x2=10.36 //y2=2.085
cc_142 ( N_GND_c_5_p N_B_c_1805_n ) capacitor c=0.00179096f //x=8.88 //y=0 \
 //x2=10.36 //y2=2.085
cc_143 ( N_GND_c_6_p N_B_c_1805_n ) capacitor c=0.0276202f //x=11.1 //y=0 \
 //x2=10.36 //y2=2.085
cc_144 ( N_GND_M5_noxref_s N_B_c_1805_n ) capacitor c=0.00773905f //x=9.375 \
 //y=0.37 //x2=10.36 //y2=2.085
cc_145 ( N_GND_c_12_p N_B_c_1810_n ) capacitor c=0.0170136f //x=27.75 //y=0 \
 //x2=28.86 //y2=2.08
cc_146 ( N_GND_c_26_p N_B_c_1811_n ) capacitor c=0.0119174f //x=9.9 //y=0.535 \
 //x2=9.72 //y2=0.91
cc_147 ( N_GND_M5_noxref_s N_B_c_1811_n ) capacitor c=0.0143355f //x=9.375 \
 //y=0.37 //x2=9.72 //y2=0.91
cc_148 ( N_GND_M5_noxref_s N_B_c_1813_n ) capacitor c=0.0074042f //x=9.375 \
 //y=0.37 //x2=9.72 //y2=1.255
cc_149 ( N_GND_M5_noxref_s N_B_c_1814_n ) capacitor c=0.00489f //x=9.375 \
 //y=0.37 //x2=10.095 //y2=0.755
cc_150 ( N_GND_c_27_p N_B_c_1815_n ) capacitor c=0.0123171f //x=10.385 \
 //y=0.535 //x2=10.25 //y2=0.91
cc_151 ( N_GND_M5_noxref_s N_B_c_1815_n ) capacitor c=0.0317181f //x=9.375 \
 //y=0.37 //x2=10.25 //y2=0.91
cc_152 ( N_GND_c_6_p N_B_c_1817_n ) capacitor c=0.00175661f //x=11.1 //y=0 \
 //x2=10.25 //y2=1.92
cc_153 ( N_GND_c_45_p N_B_c_1818_n ) capacitor c=0.00135046f //x=28.845 //y=0 \
 //x2=28.665 //y2=0.865
cc_154 ( N_GND_M15_noxref_d N_B_c_1818_n ) capacitor c=0.00220047f //x=28.74 \
 //y=0.865 //x2=28.665 //y2=0.865
cc_155 ( N_GND_M15_noxref_d N_B_c_1820_n ) capacitor c=0.00255985f //x=28.74 \
 //y=0.865 //x2=28.665 //y2=1.21
cc_156 ( N_GND_c_12_p N_B_c_1821_n ) capacitor c=0.00754269f //x=27.75 //y=0 \
 //x2=28.665 //y2=1.915
cc_157 ( N_GND_M15_noxref_d N_B_c_1822_n ) capacitor c=0.0131326f //x=28.74 \
 //y=0.865 //x2=29.04 //y2=0.71
cc_158 ( N_GND_M15_noxref_d N_B_c_1823_n ) capacitor c=0.00193127f //x=28.74 \
 //y=0.865 //x2=29.04 //y2=1.365
cc_159 ( N_GND_c_46_p N_B_c_1824_n ) capacitor c=0.00130622f //x=30.91 //y=0 \
 //x2=29.195 //y2=0.865
cc_160 ( N_GND_M15_noxref_d N_B_c_1824_n ) capacitor c=0.00257848f //x=28.74 \
 //y=0.865 //x2=29.195 //y2=0.865
cc_161 ( N_GND_M15_noxref_d N_B_c_1826_n ) capacitor c=0.00255985f //x=28.74 \
 //y=0.865 //x2=29.195 //y2=1.21
cc_162 ( N_GND_c_27_p N_B_c_1827_n ) capacitor c=2.1838e-19 //x=10.385 \
 //y=0.535 //x2=10.25 //y2=2.085
cc_163 ( N_GND_c_6_p N_B_c_1827_n ) capacitor c=0.00758987f //x=11.1 //y=0 \
 //x2=10.25 //y2=2.085
cc_164 ( N_GND_M5_noxref_s N_B_c_1827_n ) capacitor c=0.00628106f //x=9.375 \
 //y=0.37 //x2=10.25 //y2=2.085
cc_165 ( N_GND_c_6_p N_noxref_7_c_2182_n ) capacitor c=0.00424907f //x=11.1 \
 //y=0 //x2=11.725 //y2=3.7
cc_166 ( N_GND_c_7_p N_noxref_7_c_2183_n ) capacitor c=0.0263477f //x=13.32 \
 //y=0 //x2=23.935 //y2=2.22
cc_167 ( N_GND_c_8_p N_noxref_7_c_2183_n ) capacitor c=0.0263477f //x=16.65 \
 //y=0 //x2=23.935 //y2=2.22
cc_168 ( N_GND_c_9_p N_noxref_7_c_2183_n ) capacitor c=0.0272821f //x=19.98 \
 //y=0 //x2=23.935 //y2=2.22
cc_169 ( N_GND_c_10_p N_noxref_7_c_2183_n ) capacitor c=0.0328483f //x=22.2 \
 //y=0 //x2=23.935 //y2=2.22
cc_170 ( N_GND_c_6_p N_noxref_7_c_2187_n ) capacitor c=0.00785146f //x=11.1 \
 //y=0 //x2=11.955 //y2=2.22
cc_171 ( N_GND_c_7_p N_noxref_7_c_2188_n ) capacitor c=0.00249386f //x=13.32 \
 //y=0 //x2=14.315 //y2=4.07
cc_172 ( N_GND_c_4_p N_noxref_7_c_2189_n ) capacitor c=0.0398042f //x=5.55 \
 //y=0 //x2=4.725 //y2=1.655
cc_173 ( N_GND_c_3_p N_noxref_7_c_2190_n ) capacitor c=5.00558e-19 //x=2.22 \
 //y=0 //x2=4.81 //y2=3.7
cc_174 ( N_GND_c_5_p N_noxref_7_c_2191_n ) capacitor c=0.0420788f //x=8.88 \
 //y=0 //x2=8.055 //y2=1.655
cc_175 ( N_GND_M5_noxref_s N_noxref_7_c_2191_n ) capacitor c=3.42693e-19 \
 //x=9.375 //y=0.37 //x2=8.055 //y2=1.655
cc_176 ( N_GND_c_16_p N_noxref_7_c_2193_n ) capacitor c=0.00115146f //x=38.48 \
 //y=0 //x2=11.84 //y2=2.085
cc_177 ( N_GND_c_30_p N_noxref_7_c_2193_n ) capacitor c=4.37744e-19 //x=12.13 \
 //y=0.535 //x2=11.84 //y2=2.085
cc_178 ( N_GND_c_6_p N_noxref_7_c_2193_n ) capacitor c=0.0263296f //x=11.1 \
 //y=0 //x2=11.84 //y2=2.085
cc_179 ( N_GND_c_7_p N_noxref_7_c_2193_n ) capacitor c=9.68873e-19 //x=13.32 \
 //y=0 //x2=11.84 //y2=2.085
cc_180 ( N_GND_M6_noxref_s N_noxref_7_c_2193_n ) capacitor c=0.00818136f \
 //x=11.595 //y=0.37 //x2=11.84 //y2=2.085
cc_181 ( N_GND_c_7_p N_noxref_7_c_2198_n ) capacitor c=0.0125895f //x=13.32 \
 //y=0 //x2=14.43 //y2=2.085
cc_182 ( N_GND_c_10_p N_noxref_7_c_2199_n ) capacitor c=6.92793e-19 //x=22.2 \
 //y=0 //x2=24.05 //y2=2.08
cc_183 ( N_GND_c_11_p N_noxref_7_c_2199_n ) capacitor c=0.00118341f //x=25.53 \
 //y=0 //x2=24.05 //y2=2.08
cc_184 ( N_GND_c_30_p N_noxref_7_c_2201_n ) capacitor c=0.0123171f //x=12.13 \
 //y=0.535 //x2=11.95 //y2=0.91
cc_185 ( N_GND_M6_noxref_s N_noxref_7_c_2201_n ) capacitor c=0.0316686f \
 //x=11.595 //y=0.37 //x2=11.95 //y2=0.91
cc_186 ( N_GND_c_6_p N_noxref_7_c_2203_n ) capacitor c=0.00175661f //x=11.1 \
 //y=0 //x2=11.95 //y2=1.92
cc_187 ( N_GND_M6_noxref_s N_noxref_7_c_2204_n ) capacitor c=0.00489f \
 //x=11.595 //y=0.37 //x2=12.325 //y2=0.755
cc_188 ( N_GND_c_188_p N_noxref_7_c_2205_n ) capacitor c=0.0119174f //x=12.615 \
 //y=0.535 //x2=12.48 //y2=0.91
cc_189 ( N_GND_M6_noxref_s N_noxref_7_c_2205_n ) capacitor c=0.0143355f \
 //x=11.595 //y=0.37 //x2=12.48 //y2=0.91
cc_190 ( N_GND_M6_noxref_s N_noxref_7_c_2207_n ) capacitor c=0.0074042f \
 //x=11.595 //y=0.37 //x2=12.48 //y2=1.255
cc_191 ( N_GND_c_32_p N_noxref_7_c_2208_n ) capacitor c=0.00134217f //x=14.415 \
 //y=0 //x2=14.235 //y2=0.87
cc_192 ( N_GND_M7_noxref_d N_noxref_7_c_2208_n ) capacitor c=0.00220047f \
 //x=14.31 //y=0.87 //x2=14.235 //y2=0.87
cc_193 ( N_GND_M7_noxref_d N_noxref_7_c_2210_n ) capacitor c=0.00255985f \
 //x=14.31 //y=0.87 //x2=14.235 //y2=1.215
cc_194 ( N_GND_c_7_p N_noxref_7_c_2211_n ) capacitor c=0.00786098f //x=13.32 \
 //y=0 //x2=14.235 //y2=1.92
cc_195 ( N_GND_M7_noxref_d N_noxref_7_c_2212_n ) capacitor c=0.013135f \
 //x=14.31 //y=0.87 //x2=14.61 //y2=0.715
cc_196 ( N_GND_M7_noxref_d N_noxref_7_c_2213_n ) capacitor c=0.00193136f \
 //x=14.31 //y=0.87 //x2=14.61 //y2=1.37
cc_197 ( N_GND_c_33_p N_noxref_7_c_2214_n ) capacitor c=0.00129817f //x=16.48 \
 //y=0 //x2=14.765 //y2=0.87
cc_198 ( N_GND_M7_noxref_d N_noxref_7_c_2214_n ) capacitor c=0.00257848f \
 //x=14.31 //y=0.87 //x2=14.765 //y2=0.87
cc_199 ( N_GND_M7_noxref_d N_noxref_7_c_2216_n ) capacitor c=0.00255985f \
 //x=14.31 //y=0.87 //x2=14.765 //y2=1.215
cc_200 ( N_GND_c_30_p N_noxref_7_c_2217_n ) capacitor c=2.1838e-19 //x=12.13 \
 //y=0.535 //x2=11.84 //y2=2.085
cc_201 ( N_GND_c_6_p N_noxref_7_c_2217_n ) capacitor c=0.00703903f //x=11.1 \
 //y=0 //x2=11.84 //y2=2.085
cc_202 ( N_GND_M6_noxref_s N_noxref_7_c_2217_n ) capacitor c=0.00628106f \
 //x=11.595 //y=0.37 //x2=11.84 //y2=2.085
cc_203 ( N_GND_c_3_p N_noxref_7_M2_noxref_d ) capacitor c=8.60262e-19 //x=2.22 \
 //y=0 //x2=4.18 //y2=0.91
cc_204 ( N_GND_c_4_p N_noxref_7_M2_noxref_d ) capacitor c=0.00605305f //x=5.55 \
 //y=0 //x2=4.18 //y2=0.91
cc_205 ( N_GND_M1_noxref_d N_noxref_7_M2_noxref_d ) capacitor c=0.00143464f \
 //x=3.21 //y=0.87 //x2=4.18 //y2=0.91
cc_206 ( N_GND_c_4_p N_noxref_7_M4_noxref_d ) capacitor c=8.60262e-19 //x=5.55 \
 //y=0 //x2=7.51 //y2=0.91
cc_207 ( N_GND_c_5_p N_noxref_7_M4_noxref_d ) capacitor c=0.00605305f //x=8.88 \
 //y=0 //x2=7.51 //y2=0.91
cc_208 ( N_GND_M3_noxref_d N_noxref_7_M4_noxref_d ) capacitor c=0.00143464f \
 //x=6.54 //y=0.87 //x2=7.51 //y2=0.91
cc_209 ( N_GND_M5_noxref_s N_noxref_7_M4_noxref_d ) capacitor c=2.07711e-19 \
 //x=9.375 //y=0.37 //x2=7.51 //y2=0.91
cc_210 ( N_GND_c_7_p N_noxref_8_c_2602_n ) capacitor c=0.0266307f //x=13.32 \
 //y=0 //x2=18.755 //y2=2.59
cc_211 ( N_GND_c_8_p N_noxref_8_c_2602_n ) capacitor c=0.0215583f //x=16.65 \
 //y=0 //x2=18.755 //y2=2.59
cc_212 ( N_GND_c_7_p N_noxref_8_c_2604_n ) capacitor c=0.00209945f //x=13.32 \
 //y=0 //x2=12.695 //y2=2.59
cc_213 ( N_GND_c_7_p N_noxref_8_c_2605_n ) capacitor c=0.0233691f //x=13.32 \
 //y=0 //x2=12.495 //y2=2.08
cc_214 ( N_GND_M6_noxref_s N_noxref_8_c_2605_n ) capacitor c=0.00938913f \
 //x=11.595 //y=0.37 //x2=12.495 //y2=2.08
cc_215 ( N_GND_c_6_p N_noxref_8_c_2607_n ) capacitor c=9.87351e-19 //x=11.1 \
 //y=0 //x2=12.58 //y2=2.59
cc_216 ( N_GND_c_7_p N_noxref_8_c_2607_n ) capacitor c=5.56859e-19 //x=13.32 \
 //y=0 //x2=12.58 //y2=2.59
cc_217 ( N_GND_M6_noxref_s N_noxref_8_c_2607_n ) capacitor c=2.30929e-19 \
 //x=11.595 //y=0.37 //x2=12.58 //y2=2.59
cc_218 ( N_GND_c_8_p N_noxref_8_c_2610_n ) capacitor c=4.76105e-19 //x=16.65 \
 //y=0 //x2=18.87 //y2=2.085
cc_219 ( N_GND_c_9_p N_noxref_8_c_2610_n ) capacitor c=0.00140512f //x=19.98 \
 //y=0 //x2=18.87 //y2=2.085
cc_220 ( N_GND_c_16_p N_noxref_8_M6_noxref_d ) capacitor c=0.00108086f \
 //x=38.48 //y=0 //x2=12.025 //y2=0.91
cc_221 ( N_GND_c_30_p N_noxref_8_M6_noxref_d ) capacitor c=0.0147002f \
 //x=12.13 //y=0.535 //x2=12.025 //y2=0.91
cc_222 ( N_GND_c_6_p N_noxref_8_M6_noxref_d ) capacitor c=0.00721466f //x=11.1 \
 //y=0 //x2=12.025 //y2=0.91
cc_223 ( N_GND_c_7_p N_noxref_8_M6_noxref_d ) capacitor c=0.00687171f \
 //x=13.32 //y=0 //x2=12.025 //y2=0.91
cc_224 ( N_GND_M6_noxref_s N_noxref_8_M6_noxref_d ) capacitor c=0.076995f \
 //x=11.595 //y=0.37 //x2=12.025 //y2=0.91
cc_225 ( N_GND_c_8_p N_SUM_c_2765_n ) capacitor c=0.0377958f //x=16.65 //y=0 \
 //x2=15.825 //y2=1.655
cc_226 ( N_GND_c_9_p N_SUM_c_2766_n ) capacitor c=0.0397037f //x=19.98 //y=0 \
 //x2=19.155 //y2=1.655
cc_227 ( N_GND_M11_noxref_s N_SUM_c_2766_n ) capacitor c=3.42693e-19 \
 //x=20.475 //y=0.37 //x2=19.155 //y2=1.655
cc_228 ( N_GND_c_7_p N_SUM_M8_noxref_d ) capacitor c=8.60262e-19 //x=13.32 \
 //y=0 //x2=15.28 //y2=0.91
cc_229 ( N_GND_c_8_p N_SUM_M8_noxref_d ) capacitor c=0.00605305f //x=16.65 \
 //y=0 //x2=15.28 //y2=0.91
cc_230 ( N_GND_M7_noxref_d N_SUM_M8_noxref_d ) capacitor c=0.00143464f \
 //x=14.31 //y=0.87 //x2=15.28 //y2=0.91
cc_231 ( N_GND_c_8_p N_SUM_M10_noxref_d ) capacitor c=8.60262e-19 //x=16.65 \
 //y=0 //x2=18.61 //y2=0.91
cc_232 ( N_GND_c_9_p N_SUM_M10_noxref_d ) capacitor c=0.00605305f //x=19.98 \
 //y=0 //x2=18.61 //y2=0.91
cc_233 ( N_GND_M9_noxref_d N_SUM_M10_noxref_d ) capacitor c=0.00143464f \
 //x=17.64 //y=0.87 //x2=18.61 //y2=0.91
cc_234 ( N_GND_M11_noxref_s N_SUM_M10_noxref_d ) capacitor c=2.07711e-19 \
 //x=20.475 //y=0.37 //x2=18.61 //y2=0.91
cc_235 ( N_GND_c_8_p N_noxref_10_c_2913_n ) capacitor c=0.012648f //x=16.65 \
 //y=0 //x2=17.76 //y2=2.085
cc_236 ( N_GND_c_10_p N_noxref_10_c_2914_n ) capacitor c=9.6767e-19 //x=22.2 \
 //y=0 //x2=20.72 //y2=3.33
cc_237 ( N_GND_M11_noxref_s N_noxref_10_c_2915_n ) capacitor c=0.00188935f \
 //x=20.475 //y=0.37 //x2=21.005 //y2=2.08
cc_238 ( N_GND_c_37_p N_noxref_10_c_2916_n ) capacitor c=0.00188935f //x=21 \
 //y=0.535 //x2=20.805 //y2=2.08
cc_239 ( N_GND_c_9_p N_noxref_10_c_2916_n ) capacitor c=0.0263707f //x=19.98 \
 //y=0 //x2=20.805 //y2=2.08
cc_240 ( N_GND_M11_noxref_s N_noxref_10_c_2916_n ) capacitor c=0.00561042f \
 //x=20.475 //y=0.37 //x2=20.805 //y2=2.08
cc_241 ( N_GND_c_34_p N_noxref_10_c_2919_n ) capacitor c=0.00134217f \
 //x=17.745 //y=0 //x2=17.565 //y2=0.87
cc_242 ( N_GND_M9_noxref_d N_noxref_10_c_2919_n ) capacitor c=0.00220047f \
 //x=17.64 //y=0.87 //x2=17.565 //y2=0.87
cc_243 ( N_GND_M9_noxref_d N_noxref_10_c_2921_n ) capacitor c=0.00255985f \
 //x=17.64 //y=0.87 //x2=17.565 //y2=1.215
cc_244 ( N_GND_c_8_p N_noxref_10_c_2922_n ) capacitor c=0.00176175f //x=16.65 \
 //y=0 //x2=17.565 //y2=1.525
cc_245 ( N_GND_c_8_p N_noxref_10_c_2923_n ) capacitor c=0.0080354f //x=16.65 \
 //y=0 //x2=17.565 //y2=1.92
cc_246 ( N_GND_M9_noxref_d N_noxref_10_c_2924_n ) capacitor c=0.013135f \
 //x=17.64 //y=0.87 //x2=17.94 //y2=0.715
cc_247 ( N_GND_M9_noxref_d N_noxref_10_c_2925_n ) capacitor c=0.00193136f \
 //x=17.64 //y=0.87 //x2=17.94 //y2=1.37
cc_248 ( N_GND_c_35_p N_noxref_10_c_2926_n ) capacitor c=0.00129817f //x=19.81 \
 //y=0 //x2=18.095 //y2=0.87
cc_249 ( N_GND_M9_noxref_d N_noxref_10_c_2926_n ) capacitor c=0.00257848f \
 //x=17.64 //y=0.87 //x2=18.095 //y2=0.87
cc_250 ( N_GND_M9_noxref_d N_noxref_10_c_2928_n ) capacitor c=0.00255985f \
 //x=17.64 //y=0.87 //x2=18.095 //y2=1.215
cc_251 ( N_GND_c_16_p N_noxref_10_M11_noxref_d ) capacitor c=0.00108086f \
 //x=38.48 //y=0 //x2=20.895 //y2=0.91
cc_252 ( N_GND_c_9_p N_noxref_10_M11_noxref_d ) capacitor c=0.00686786f \
 //x=19.98 //y=0 //x2=20.895 //y2=0.91
cc_253 ( N_GND_c_10_p N_noxref_10_M11_noxref_d ) capacitor c=0.00721119f \
 //x=22.2 //y=0 //x2=20.895 //y2=0.91
cc_254 ( N_GND_M11_noxref_s N_noxref_10_M11_noxref_d ) capacitor c=0.0916952f \
 //x=20.475 //y=0.37 //x2=20.895 //y2=0.91
cc_255 ( N_GND_c_8_p N_CIN_c_3085_n ) capacitor c=0.00750857f //x=16.65 //y=0 \
 //x2=21.345 //y2=2.96
cc_256 ( N_GND_c_9_p N_CIN_c_3085_n ) capacitor c=0.00949826f //x=19.98 //y=0 \
 //x2=21.345 //y2=2.96
cc_257 ( N_GND_c_10_p N_CIN_c_3087_n ) capacitor c=0.00169673f //x=22.2 //y=0 \
 //x2=23.195 //y2=4.44
cc_258 ( N_GND_c_7_p N_CIN_c_3088_n ) capacitor c=4.86635e-19 //x=13.32 //y=0 \
 //x2=15.54 //y2=2.085
cc_259 ( N_GND_c_8_p N_CIN_c_3088_n ) capacitor c=0.00121037f //x=16.65 //y=0 \
 //x2=15.54 //y2=2.085
cc_260 ( N_GND_c_16_p N_CIN_c_3090_n ) capacitor c=0.00115146f //x=38.48 //y=0 \
 //x2=21.46 //y2=2.085
cc_261 ( N_GND_c_38_p N_CIN_c_3090_n ) capacitor c=4.37744e-19 //x=21.485 \
 //y=0.535 //x2=21.46 //y2=2.085
cc_262 ( N_GND_c_9_p N_CIN_c_3090_n ) capacitor c=0.00103703f //x=19.98 //y=0 \
 //x2=21.46 //y2=2.085
cc_263 ( N_GND_c_10_p N_CIN_c_3090_n ) capacitor c=0.0261601f //x=22.2 //y=0 \
 //x2=21.46 //y2=2.085
cc_264 ( N_GND_M11_noxref_s N_CIN_c_3090_n ) capacitor c=0.00772882f \
 //x=20.475 //y=0.37 //x2=21.46 //y2=2.085
cc_265 ( N_GND_c_10_p N_CIN_c_3095_n ) capacitor c=0.0152752f //x=22.2 //y=0 \
 //x2=23.31 //y2=2.08
cc_266 ( N_GND_c_37_p N_CIN_c_3096_n ) capacitor c=0.0119174f //x=21 //y=0.535 \
 //x2=20.82 //y2=0.91
cc_267 ( N_GND_M11_noxref_s N_CIN_c_3096_n ) capacitor c=0.0143355f //x=20.475 \
 //y=0.37 //x2=20.82 //y2=0.91
cc_268 ( N_GND_M11_noxref_s N_CIN_c_3098_n ) capacitor c=0.0074042f //x=20.475 \
 //y=0.37 //x2=20.82 //y2=1.255
cc_269 ( N_GND_M11_noxref_s N_CIN_c_3099_n ) capacitor c=0.00489f //x=20.475 \
 //y=0.37 //x2=21.195 //y2=0.755
cc_270 ( N_GND_c_38_p N_CIN_c_3100_n ) capacitor c=0.0123171f //x=21.485 \
 //y=0.535 //x2=21.35 //y2=0.91
cc_271 ( N_GND_M11_noxref_s N_CIN_c_3100_n ) capacitor c=0.0317792f //x=20.475 \
 //y=0.37 //x2=21.35 //y2=0.91
cc_272 ( N_GND_c_10_p N_CIN_c_3102_n ) capacitor c=0.00189677f //x=22.2 //y=0 \
 //x2=21.35 //y2=1.92
cc_273 ( N_GND_c_40_p N_CIN_c_3103_n ) capacitor c=0.00135046f //x=23.295 \
 //y=0 //x2=23.115 //y2=0.865
cc_274 ( N_GND_M12_noxref_d N_CIN_c_3103_n ) capacitor c=0.00220047f //x=23.19 \
 //y=0.865 //x2=23.115 //y2=0.865
cc_275 ( N_GND_M12_noxref_d N_CIN_c_3105_n ) capacitor c=0.00255985f //x=23.19 \
 //y=0.865 //x2=23.115 //y2=1.21
cc_276 ( N_GND_c_10_p N_CIN_c_3106_n ) capacitor c=0.00676835f //x=22.2 //y=0 \
 //x2=23.115 //y2=1.915
cc_277 ( N_GND_M12_noxref_d N_CIN_c_3107_n ) capacitor c=0.0131326f //x=23.19 \
 //y=0.865 //x2=23.49 //y2=0.71
cc_278 ( N_GND_M12_noxref_d N_CIN_c_3108_n ) capacitor c=0.00193127f //x=23.19 \
 //y=0.865 //x2=23.49 //y2=1.365
cc_279 ( N_GND_c_41_p N_CIN_c_3109_n ) capacitor c=0.00130622f //x=25.36 //y=0 \
 //x2=23.645 //y2=0.865
cc_280 ( N_GND_M12_noxref_d N_CIN_c_3109_n ) capacitor c=0.00257848f //x=23.19 \
 //y=0.865 //x2=23.645 //y2=0.865
cc_281 ( N_GND_M12_noxref_d N_CIN_c_3111_n ) capacitor c=0.00255985f //x=23.19 \
 //y=0.865 //x2=23.645 //y2=1.21
cc_282 ( N_GND_c_38_p N_CIN_c_3112_n ) capacitor c=2.1838e-19 //x=21.485 \
 //y=0.535 //x2=21.35 //y2=2.085
cc_283 ( N_GND_c_10_p N_CIN_c_3112_n ) capacitor c=0.00845889f //x=22.2 //y=0 \
 //x2=21.35 //y2=2.085
cc_284 ( N_GND_M11_noxref_s N_CIN_c_3112_n ) capacitor c=0.00628106f \
 //x=20.475 //y=0.37 //x2=21.35 //y2=2.085
cc_285 ( N_GND_c_11_p N_noxref_12_c_3336_n ) capacitor c=0.00645253f //x=25.53 \
 //y=0 //x2=26.155 //y2=3.33
cc_286 ( N_GND_c_11_p N_noxref_12_c_3337_n ) capacitor c=0.0428814f //x=25.53 \
 //y=0 //x2=24.705 //y2=1.655
cc_287 ( N_GND_M14_noxref_s N_noxref_12_c_3337_n ) capacitor c=3.37896e-19 \
 //x=26.025 //y=0.37 //x2=24.705 //y2=1.655
cc_288 ( N_GND_c_16_p N_noxref_12_c_3339_n ) capacitor c=0.00115146f //x=38.48 \
 //y=0 //x2=26.27 //y2=2.085
cc_289 ( N_GND_c_43_p N_noxref_12_c_3339_n ) capacitor c=4.37744e-19 //x=26.56 \
 //y=0.535 //x2=26.27 //y2=2.085
cc_290 ( N_GND_c_11_p N_noxref_12_c_3339_n ) capacitor c=0.0285768f //x=25.53 \
 //y=0 //x2=26.27 //y2=2.085
cc_291 ( N_GND_c_12_p N_noxref_12_c_3339_n ) capacitor c=0.00130094f //x=27.75 \
 //y=0 //x2=26.27 //y2=2.085
cc_292 ( N_GND_M14_noxref_s N_noxref_12_c_3339_n ) capacitor c=0.00779289f \
 //x=26.025 //y=0.37 //x2=26.27 //y2=2.085
cc_293 ( N_GND_c_43_p N_noxref_12_c_3344_n ) capacitor c=0.0123171f //x=26.56 \
 //y=0.535 //x2=26.38 //y2=0.91
cc_294 ( N_GND_M14_noxref_s N_noxref_12_c_3344_n ) capacitor c=0.0317689f \
 //x=26.025 //y=0.37 //x2=26.38 //y2=0.91
cc_295 ( N_GND_c_11_p N_noxref_12_c_3346_n ) capacitor c=0.00361526f //x=25.53 \
 //y=0 //x2=26.38 //y2=1.92
cc_296 ( N_GND_M14_noxref_s N_noxref_12_c_3347_n ) capacitor c=0.00489f \
 //x=26.025 //y=0.37 //x2=26.755 //y2=0.755
cc_297 ( N_GND_c_297_p N_noxref_12_c_3348_n ) capacitor c=0.0119174f \
 //x=27.045 //y=0.535 //x2=26.91 //y2=0.91
cc_298 ( N_GND_M14_noxref_s N_noxref_12_c_3348_n ) capacitor c=0.0143355f \
 //x=26.025 //y=0.37 //x2=26.91 //y2=0.91
cc_299 ( N_GND_M14_noxref_s N_noxref_12_c_3350_n ) capacitor c=0.0074042f \
 //x=26.025 //y=0.37 //x2=26.91 //y2=1.255
cc_300 ( N_GND_c_43_p N_noxref_12_c_3351_n ) capacitor c=2.1838e-19 //x=26.56 \
 //y=0.535 //x2=26.27 //y2=2.085
cc_301 ( N_GND_c_11_p N_noxref_12_c_3351_n ) capacitor c=0.00920617f //x=25.53 \
 //y=0 //x2=26.27 //y2=2.085
cc_302 ( N_GND_M14_noxref_s N_noxref_12_c_3351_n ) capacitor c=0.00628106f \
 //x=26.025 //y=0.37 //x2=26.27 //y2=2.085
cc_303 ( N_GND_c_10_p N_noxref_12_M13_noxref_d ) capacitor c=8.58106e-19 \
 //x=22.2 //y=0 //x2=24.16 //y2=0.905
cc_304 ( N_GND_c_11_p N_noxref_12_M13_noxref_d ) capacitor c=0.00616547f \
 //x=25.53 //y=0 //x2=24.16 //y2=0.905
cc_305 ( N_GND_M12_noxref_d N_noxref_12_M13_noxref_d ) capacitor c=0.00143464f \
 //x=23.19 //y=0.865 //x2=24.16 //y2=0.905
cc_306 ( N_GND_M14_noxref_s N_noxref_12_M13_noxref_d ) capacitor c=2.09402e-19 \
 //x=26.025 //y=0.37 //x2=24.16 //y2=0.905
cc_307 ( N_GND_c_13_p N_noxref_13_c_3475_n ) capacitor c=0.044612f //x=31.08 \
 //y=0 //x2=30.255 //y2=1.655
cc_308 ( N_GND_M17_noxref_s N_noxref_13_c_3475_n ) capacitor c=3.37896e-19 \
 //x=31.575 //y=0.37 //x2=30.255 //y2=1.655
cc_309 ( N_GND_c_12_p N_noxref_13_c_3477_n ) capacitor c=5.0384e-19 //x=27.75 \
 //y=0 //x2=30.34 //y2=3.33
cc_310 ( N_GND_c_16_p N_noxref_13_c_3478_n ) capacitor c=0.00183858f //x=38.48 \
 //y=0 //x2=31.82 //y2=2.085
cc_311 ( N_GND_c_311_p N_noxref_13_c_3478_n ) capacitor c=7.85046e-19 \
 //x=32.11 //y=0.535 //x2=31.82 //y2=2.085
cc_312 ( N_GND_c_13_p N_noxref_13_c_3478_n ) capacitor c=0.0287905f //x=31.08 \
 //y=0 //x2=31.82 //y2=2.085
cc_313 ( N_GND_c_14_p N_noxref_13_c_3478_n ) capacitor c=0.00118911f //x=33.3 \
 //y=0 //x2=31.82 //y2=2.085
cc_314 ( N_GND_M17_noxref_s N_noxref_13_c_3478_n ) capacitor c=0.010785f \
 //x=31.575 //y=0.37 //x2=31.82 //y2=2.085
cc_315 ( N_GND_c_311_p N_noxref_13_c_3483_n ) capacitor c=0.0123171f //x=32.11 \
 //y=0.535 //x2=31.93 //y2=0.91
cc_316 ( N_GND_M17_noxref_s N_noxref_13_c_3483_n ) capacitor c=0.0317792f \
 //x=31.575 //y=0.37 //x2=31.93 //y2=0.91
cc_317 ( N_GND_c_13_p N_noxref_13_c_3485_n ) capacitor c=0.00465161f //x=31.08 \
 //y=0 //x2=31.93 //y2=1.92
cc_318 ( N_GND_M17_noxref_s N_noxref_13_c_3486_n ) capacitor c=0.00489f \
 //x=31.575 //y=0.37 //x2=32.305 //y2=0.755
cc_319 ( N_GND_c_319_p N_noxref_13_c_3487_n ) capacitor c=0.0119174f \
 //x=32.595 //y=0.535 //x2=32.46 //y2=0.91
cc_320 ( N_GND_M17_noxref_s N_noxref_13_c_3487_n ) capacitor c=0.0143355f \
 //x=31.575 //y=0.37 //x2=32.46 //y2=0.91
cc_321 ( N_GND_M17_noxref_s N_noxref_13_c_3489_n ) capacitor c=0.0074042f \
 //x=31.575 //y=0.37 //x2=32.46 //y2=1.255
cc_322 ( N_GND_c_311_p N_noxref_13_c_3490_n ) capacitor c=2.1838e-19 //x=32.11 \
 //y=0.535 //x2=31.82 //y2=2.085
cc_323 ( N_GND_c_13_p N_noxref_13_c_3490_n ) capacitor c=0.00769211f //x=31.08 \
 //y=0 //x2=31.82 //y2=2.085
cc_324 ( N_GND_M17_noxref_s N_noxref_13_c_3490_n ) capacitor c=0.0065286f \
 //x=31.575 //y=0.37 //x2=31.82 //y2=2.085
cc_325 ( N_GND_c_12_p N_noxref_13_M16_noxref_d ) capacitor c=8.58106e-19 \
 //x=27.75 //y=0 //x2=29.71 //y2=0.905
cc_326 ( N_GND_c_13_p N_noxref_13_M16_noxref_d ) capacitor c=0.00616547f \
 //x=31.08 //y=0 //x2=29.71 //y2=0.905
cc_327 ( N_GND_M15_noxref_d N_noxref_13_M16_noxref_d ) capacitor c=0.00143464f \
 //x=28.74 //y=0.865 //x2=29.71 //y2=0.905
cc_328 ( N_GND_M17_noxref_s N_noxref_13_M16_noxref_d ) capacitor c=2.09402e-19 \
 //x=31.575 //y=0.37 //x2=29.71 //y2=0.905
cc_329 ( N_GND_c_16_p N_noxref_14_c_3617_n ) capacitor c=0.0416947f //x=38.48 \
 //y=0 //x2=34.295 //y2=2.96
cc_330 ( N_GND_c_46_p N_noxref_14_c_3617_n ) capacitor c=0.00208984f //x=30.91 \
 //y=0 //x2=34.295 //y2=2.96
cc_331 ( N_GND_c_331_p N_noxref_14_c_3617_n ) capacitor c=0.00134487f \
 //x=31.625 //y=0 //x2=34.295 //y2=2.96
cc_332 ( N_GND_c_311_p N_noxref_14_c_3617_n ) capacitor c=0.00140351f \
 //x=32.11 //y=0.535 //x2=34.295 //y2=2.96
cc_333 ( N_GND_c_333_p N_noxref_14_c_3617_n ) capacitor c=0.00129597f \
 //x=33.13 //y=0 //x2=34.295 //y2=2.96
cc_334 ( N_GND_c_334_p N_noxref_14_c_3617_n ) capacitor c=0.00166275f \
 //x=33.91 //y=0 //x2=34.295 //y2=2.96
cc_335 ( N_GND_c_335_p N_noxref_14_c_3617_n ) capacitor c=0.00160088f \
 //x=34.395 //y=0.53 //x2=34.295 //y2=2.96
cc_336 ( N_GND_c_12_p N_noxref_14_c_3617_n ) capacitor c=0.0110081f //x=27.75 \
 //y=0 //x2=34.295 //y2=2.96
cc_337 ( N_GND_c_13_p N_noxref_14_c_3617_n ) capacitor c=0.0144849f //x=31.08 \
 //y=0 //x2=34.295 //y2=2.96
cc_338 ( N_GND_c_14_p N_noxref_14_c_3617_n ) capacitor c=0.0144849f //x=33.3 \
 //y=0 //x2=34.295 //y2=2.96
cc_339 ( N_GND_M17_noxref_s N_noxref_14_c_3617_n ) capacitor c=0.00500287f \
 //x=31.575 //y=0.37 //x2=34.295 //y2=2.96
cc_340 ( N_GND_M18_noxref_s N_noxref_14_c_3617_n ) capacitor c=0.00335259f \
 //x=33.86 //y=0.365 //x2=34.295 //y2=2.96
cc_341 ( N_GND_c_12_p N_noxref_14_c_3629_n ) capacitor c=0.0289399f //x=27.75 \
 //y=0 //x2=26.925 //y2=2.08
cc_342 ( N_GND_M14_noxref_s N_noxref_14_c_3629_n ) capacitor c=0.00796381f \
 //x=26.025 //y=0.37 //x2=26.925 //y2=2.08
cc_343 ( N_GND_c_11_p N_noxref_14_c_3631_n ) capacitor c=9.12652e-19 //x=25.53 \
 //y=0 //x2=27.01 //y2=2.96
cc_344 ( N_GND_c_16_p N_noxref_14_c_3632_n ) capacitor c=5.88914e-19 //x=38.48 \
 //y=0 //x2=34.41 //y2=2.08
cc_345 ( N_GND_c_335_p N_noxref_14_c_3632_n ) capacitor c=0.00134181f \
 //x=34.395 //y=0.53 //x2=34.41 //y2=2.08
cc_346 ( N_GND_c_14_p N_noxref_14_c_3632_n ) capacitor c=0.0175793f //x=33.3 \
 //y=0 //x2=34.41 //y2=2.08
cc_347 ( N_GND_c_335_p N_noxref_14_c_3635_n ) capacitor c=0.0126019f \
 //x=34.395 //y=0.53 //x2=34.215 //y2=0.905
cc_348 ( N_GND_M18_noxref_s N_noxref_14_c_3635_n ) capacitor c=0.0318086f \
 //x=33.86 //y=0.365 //x2=34.215 //y2=0.905
cc_349 ( N_GND_c_335_p N_noxref_14_c_3637_n ) capacitor c=2.1838e-19 \
 //x=34.395 //y=0.53 //x2=34.215 //y2=1.915
cc_350 ( N_GND_c_14_p N_noxref_14_c_3637_n ) capacitor c=0.0114883f //x=33.3 \
 //y=0 //x2=34.215 //y2=1.915
cc_351 ( N_GND_M18_noxref_s N_noxref_14_c_3639_n ) capacitor c=0.00479092f \
 //x=33.86 //y=0.365 //x2=34.59 //y2=0.75
cc_352 ( N_GND_c_352_p N_noxref_14_c_3640_n ) capacitor c=0.0113555f //x=34.88 \
 //y=0.53 //x2=34.745 //y2=0.905
cc_353 ( N_GND_M18_noxref_s N_noxref_14_c_3640_n ) capacitor c=0.00514143f \
 //x=33.86 //y=0.365 //x2=34.745 //y2=0.905
cc_354 ( N_GND_M18_noxref_s N_noxref_14_c_3642_n ) capacitor c=8.33128e-19 \
 //x=33.86 //y=0.365 //x2=34.745 //y2=1.25
cc_355 ( N_GND_c_16_p N_noxref_14_M14_noxref_d ) capacitor c=0.00108086f \
 //x=38.48 //y=0 //x2=26.455 //y2=0.91
cc_356 ( N_GND_c_43_p N_noxref_14_M14_noxref_d ) capacitor c=0.0147002f \
 //x=26.56 //y=0.535 //x2=26.455 //y2=0.91
cc_357 ( N_GND_c_11_p N_noxref_14_M14_noxref_d ) capacitor c=0.00737694f \
 //x=25.53 //y=0 //x2=26.455 //y2=0.91
cc_358 ( N_GND_c_12_p N_noxref_14_M14_noxref_d ) capacitor c=0.0068044f \
 //x=27.75 //y=0 //x2=26.455 //y2=0.91
cc_359 ( N_GND_M14_noxref_s N_noxref_14_M14_noxref_d ) capacitor c=0.076995f \
 //x=26.025 //y=0.37 //x2=26.455 //y2=0.91
cc_360 ( N_GND_c_16_p N_noxref_15_c_3782_n ) capacitor c=0.0134551f //x=38.48 \
 //y=0 //x2=35.035 //y2=3.33
cc_361 ( N_GND_c_16_p N_noxref_15_c_3783_n ) capacitor c=0.00130393f //x=38.48 \
 //y=0 //x2=32.475 //y2=2.08
cc_362 ( N_GND_c_14_p N_noxref_15_c_3783_n ) capacitor c=0.0296841f //x=33.3 \
 //y=0 //x2=32.475 //y2=2.08
cc_363 ( N_GND_M17_noxref_s N_noxref_15_c_3783_n ) capacitor c=0.00967469f \
 //x=31.575 //y=0.37 //x2=32.475 //y2=2.08
cc_364 ( N_GND_c_13_p N_noxref_15_c_3786_n ) capacitor c=9.49116e-19 //x=31.08 \
 //y=0 //x2=32.56 //y2=3.33
cc_365 ( N_GND_c_14_p N_noxref_15_c_3787_n ) capacitor c=9.2064e-19 //x=33.3 \
 //y=0 //x2=35.15 //y2=2.08
cc_366 ( N_GND_c_15_p N_noxref_15_c_3787_n ) capacitor c=9.53263e-19 //x=36.63 \
 //y=0 //x2=35.15 //y2=2.08
cc_367 ( N_GND_c_367_p N_noxref_15_c_3789_n ) capacitor c=0.0109802f \
 //x=35.365 //y=0.53 //x2=35.185 //y2=0.905
cc_368 ( N_GND_M18_noxref_s N_noxref_15_c_3789_n ) capacitor c=0.00590563f \
 //x=33.86 //y=0.365 //x2=35.185 //y2=0.905
cc_369 ( N_GND_M18_noxref_s N_noxref_15_c_3791_n ) capacitor c=0.00466751f \
 //x=33.86 //y=0.365 //x2=35.56 //y2=0.75
cc_370 ( N_GND_M18_noxref_s N_noxref_15_c_3792_n ) capacitor c=0.00316186f \
 //x=33.86 //y=0.365 //x2=35.56 //y2=1.405
cc_371 ( N_GND_c_371_p N_noxref_15_c_3793_n ) capacitor c=0.0112321f //x=35.85 \
 //y=0.53 //x2=35.715 //y2=0.905
cc_372 ( N_GND_M18_noxref_s N_noxref_15_c_3793_n ) capacitor c=0.0142835f \
 //x=33.86 //y=0.365 //x2=35.715 //y2=0.905
cc_373 ( N_GND_c_16_p N_noxref_15_M17_noxref_d ) capacitor c=0.00124113f \
 //x=38.48 //y=0 //x2=32.005 //y2=0.91
cc_374 ( N_GND_c_311_p N_noxref_15_M17_noxref_d ) capacitor c=0.0150482f \
 //x=32.11 //y=0.535 //x2=32.005 //y2=0.91
cc_375 ( N_GND_c_13_p N_noxref_15_M17_noxref_d ) capacitor c=0.00920923f \
 //x=31.08 //y=0 //x2=32.005 //y2=0.91
cc_376 ( N_GND_c_14_p N_noxref_15_M17_noxref_d ) capacitor c=0.00949241f \
 //x=33.3 //y=0 //x2=32.005 //y2=0.91
cc_377 ( N_GND_M17_noxref_s N_noxref_15_M17_noxref_d ) capacitor c=0.076995f \
 //x=31.575 //y=0.37 //x2=32.005 //y2=0.91
cc_378 ( N_GND_c_16_p N_noxref_16_c_3919_n ) capacitor c=0.0116078f //x=38.48 \
 //y=0 //x2=37.255 //y2=3.33
cc_379 ( N_GND_c_379_p N_noxref_16_c_3919_n ) capacitor c=0.00136402f \
 //x=36.46 //y=0 //x2=37.255 //y2=3.33
cc_380 ( N_GND_c_380_p N_noxref_16_c_3919_n ) capacitor c=0.00110325f \
 //x=37.175 //y=0 //x2=37.255 //y2=3.33
cc_381 ( N_GND_c_381_p N_noxref_16_c_3919_n ) capacitor c=2.76195e-19 \
 //x=37.66 //y=0.535 //x2=37.255 //y2=3.33
cc_382 ( N_GND_c_15_p N_noxref_16_c_3919_n ) capacitor c=0.00820844f //x=36.63 \
 //y=0 //x2=37.255 //y2=3.33
cc_383 ( N_GND_M20_noxref_s N_noxref_16_c_3919_n ) capacitor c=0.00164577f \
 //x=37.125 //y=0.37 //x2=37.255 //y2=3.33
cc_384 ( N_GND_c_16_p N_noxref_16_c_3925_n ) capacitor c=0.00192312f //x=38.48 \
 //y=0 //x2=36.005 //y2=3.33
cc_385 ( N_GND_M18_noxref_s N_noxref_16_c_3925_n ) capacitor c=6.50479e-19 \
 //x=33.86 //y=0.365 //x2=36.005 //y2=3.33
cc_386 ( N_GND_c_16_p N_noxref_16_c_3927_n ) capacitor c=0.00251084f //x=38.48 \
 //y=0 //x2=35.365 //y2=1.655
cc_387 ( N_GND_c_352_p N_noxref_16_c_3927_n ) capacitor c=0.00379295f \
 //x=34.88 //y=0.53 //x2=35.365 //y2=1.655
cc_388 ( N_GND_c_367_p N_noxref_16_c_3927_n ) capacitor c=0.00320231f \
 //x=35.365 //y=0.53 //x2=35.365 //y2=1.655
cc_389 ( N_GND_M18_noxref_s N_noxref_16_c_3927_n ) capacitor c=0.0170293f \
 //x=33.86 //y=0.365 //x2=35.365 //y2=1.655
cc_390 ( N_GND_c_16_p N_noxref_16_c_3931_n ) capacitor c=0.00197099f //x=38.48 \
 //y=0 //x2=35.805 //y2=1.655
cc_391 ( N_GND_c_371_p N_noxref_16_c_3931_n ) capacitor c=0.00479136f \
 //x=35.85 //y=0.53 //x2=35.805 //y2=1.655
cc_392 ( N_GND_c_15_p N_noxref_16_c_3931_n ) capacitor c=0.0464456f //x=36.63 \
 //y=0 //x2=35.805 //y2=1.655
cc_393 ( N_GND_M18_noxref_s N_noxref_16_c_3931_n ) capacitor c=0.0158743f \
 //x=33.86 //y=0.365 //x2=35.805 //y2=1.655
cc_394 ( N_GND_M20_noxref_s N_noxref_16_c_3931_n ) capacitor c=3.53679e-19 \
 //x=37.125 //y=0.37 //x2=35.805 //y2=1.655
cc_395 ( N_GND_c_14_p N_noxref_16_c_3936_n ) capacitor c=0.00101801f //x=33.3 \
 //y=0 //x2=35.89 //y2=3.33
cc_396 ( N_GND_c_16_p N_noxref_16_c_3937_n ) capacitor c=0.00184963f //x=38.48 \
 //y=0 //x2=37.37 //y2=2.085
cc_397 ( N_GND_c_381_p N_noxref_16_c_3937_n ) capacitor c=7.87839e-19 \
 //x=37.66 //y=0.535 //x2=37.37 //y2=2.085
cc_398 ( N_GND_c_1_p N_noxref_16_c_3937_n ) capacitor c=0.00118981f //x=38.48 \
 //y=0 //x2=37.37 //y2=2.085
cc_399 ( N_GND_c_15_p N_noxref_16_c_3937_n ) capacitor c=0.029021f //x=36.63 \
 //y=0 //x2=37.37 //y2=2.085
cc_400 ( N_GND_M20_noxref_s N_noxref_16_c_3937_n ) capacitor c=0.0108503f \
 //x=37.125 //y=0.37 //x2=37.37 //y2=2.085
cc_401 ( N_GND_c_381_p N_noxref_16_c_3942_n ) capacitor c=0.0121757f //x=37.66 \
 //y=0.535 //x2=37.48 //y2=0.91
cc_402 ( N_GND_M20_noxref_s N_noxref_16_c_3942_n ) capacitor c=0.0317181f \
 //x=37.125 //y=0.37 //x2=37.48 //y2=0.91
cc_403 ( N_GND_c_15_p N_noxref_16_c_3944_n ) capacitor c=0.00552709f //x=36.63 \
 //y=0 //x2=37.48 //y2=1.92
cc_404 ( N_GND_M20_noxref_s N_noxref_16_c_3945_n ) capacitor c=0.00483274f \
 //x=37.125 //y=0.37 //x2=37.855 //y2=0.755
cc_405 ( N_GND_c_405_p N_noxref_16_c_3946_n ) capacitor c=0.0118602f \
 //x=38.145 //y=0.535 //x2=38.01 //y2=0.91
cc_406 ( N_GND_M20_noxref_s N_noxref_16_c_3946_n ) capacitor c=0.0143355f \
 //x=37.125 //y=0.37 //x2=38.01 //y2=0.91
cc_407 ( N_GND_M20_noxref_s N_noxref_16_c_3948_n ) capacitor c=0.0074042f \
 //x=37.125 //y=0.37 //x2=38.01 //y2=1.255
cc_408 ( N_GND_c_381_p N_noxref_16_c_3949_n ) capacitor c=2.1838e-19 //x=37.66 \
 //y=0.535 //x2=37.37 //y2=2.085
cc_409 ( N_GND_c_15_p N_noxref_16_c_3949_n ) capacitor c=0.0108179f //x=36.63 \
 //y=0 //x2=37.37 //y2=2.085
cc_410 ( N_GND_M20_noxref_s N_noxref_16_c_3949_n ) capacitor c=0.00655738f \
 //x=37.125 //y=0.37 //x2=37.37 //y2=2.085
cc_411 ( N_GND_c_16_p N_noxref_16_M18_noxref_d ) capacitor c=0.00104706f \
 //x=38.48 //y=0 //x2=34.29 //y2=0.905
cc_412 ( N_GND_c_14_p N_noxref_16_M18_noxref_d ) capacitor c=0.00416273f \
 //x=33.3 //y=0 //x2=34.29 //y2=0.905
cc_413 ( N_GND_c_15_p N_noxref_16_M18_noxref_d ) capacitor c=2.57516e-19 \
 //x=36.63 //y=0 //x2=34.29 //y2=0.905
cc_414 ( N_GND_M18_noxref_s N_noxref_16_M18_noxref_d ) capacitor c=0.0767111f \
 //x=33.86 //y=0.365 //x2=34.29 //y2=0.905
cc_415 ( N_GND_c_16_p N_noxref_16_M19_noxref_d ) capacitor c=0.00195394f \
 //x=38.48 //y=0 //x2=35.26 //y2=0.905
cc_416 ( N_GND_c_15_p N_noxref_16_M19_noxref_d ) capacitor c=0.00609243f \
 //x=36.63 //y=0 //x2=35.26 //y2=0.905
cc_417 ( N_GND_M18_noxref_s N_noxref_16_M19_noxref_d ) capacitor c=0.0610175f \
 //x=33.86 //y=0.365 //x2=35.26 //y2=0.905
cc_418 ( N_GND_M20_noxref_s N_noxref_16_M19_noxref_d ) capacitor c=2.04477e-19 \
 //x=37.125 //y=0.37 //x2=35.26 //y2=0.905
cc_419 ( N_GND_M0_noxref_s N_noxref_18_c_4098_n ) capacitor c=0.0013253f \
 //x=0.495 //y=0.37 //x2=2.915 //y2=1.5
cc_420 ( N_GND_c_16_p N_noxref_18_c_4099_n ) capacitor c=0.00458512f //x=38.48 \
 //y=0 //x2=3.8 //y2=1.585
cc_421 ( N_GND_c_82_p N_noxref_18_c_4099_n ) capacitor c=0.0011383f //x=3.315 \
 //y=0 //x2=3.8 //y2=1.585
cc_422 ( N_GND_c_22_p N_noxref_18_c_4099_n ) capacitor c=0.00206628f //x=5.38 \
 //y=0 //x2=3.8 //y2=1.585
cc_423 ( N_GND_M1_noxref_d N_noxref_18_c_4099_n ) capacitor c=0.00879973f \
 //x=3.21 //y=0.87 //x2=3.8 //y2=1.585
cc_424 ( N_GND_c_16_p N_noxref_18_c_4103_n ) capacitor c=0.00242791f //x=38.48 \
 //y=0 //x2=3.885 //y2=0.62
cc_425 ( N_GND_c_22_p N_noxref_18_c_4103_n ) capacitor c=0.0142763f //x=5.38 \
 //y=0 //x2=3.885 //y2=0.62
cc_426 ( N_GND_M1_noxref_d N_noxref_18_c_4103_n ) capacitor c=0.033812f \
 //x=3.21 //y=0.87 //x2=3.885 //y2=0.62
cc_427 ( N_GND_c_3_p N_noxref_18_c_4106_n ) capacitor c=2.91423e-19 //x=2.22 \
 //y=0 //x2=3.885 //y2=1.5
cc_428 ( N_GND_c_16_p N_noxref_18_c_4107_n ) capacitor c=0.010074f //x=38.48 \
 //y=0 //x2=4.77 //y2=0.535
cc_429 ( N_GND_c_22_p N_noxref_18_c_4107_n ) capacitor c=0.0368958f //x=5.38 \
 //y=0 //x2=4.77 //y2=0.535
cc_430 ( N_GND_c_1_p N_noxref_18_c_4107_n ) capacitor c=0.00195382f //x=38.48 \
 //y=0 //x2=4.77 //y2=0.535
cc_431 ( N_GND_c_16_p N_noxref_18_c_4110_n ) capacitor c=0.00242513f //x=38.48 \
 //y=0 //x2=4.855 //y2=0.62
cc_432 ( N_GND_c_22_p N_noxref_18_c_4110_n ) capacitor c=0.0142124f //x=5.38 \
 //y=0 //x2=4.855 //y2=0.62
cc_433 ( N_GND_c_4_p N_noxref_18_c_4110_n ) capacitor c=0.0431718f //x=5.55 \
 //y=0 //x2=4.855 //y2=0.62
cc_434 ( N_GND_c_16_p N_noxref_18_M1_noxref_s ) capacitor c=0.0026904f \
 //x=38.48 //y=0 //x2=2.78 //y2=0.37
cc_435 ( N_GND_c_435_p N_noxref_18_M1_noxref_s ) capacitor c=0.0013253f \
 //x=1.6 //y=0.45 //x2=2.78 //y2=0.37
cc_436 ( N_GND_c_82_p N_noxref_18_M1_noxref_s ) capacitor c=0.0144735f \
 //x=3.315 //y=0 //x2=2.78 //y2=0.37
cc_437 ( N_GND_c_3_p N_noxref_18_M1_noxref_s ) capacitor c=0.058339f //x=2.22 \
 //y=0 //x2=2.78 //y2=0.37
cc_438 ( N_GND_c_4_p N_noxref_18_M1_noxref_s ) capacitor c=0.00200438f \
 //x=5.55 //y=0 //x2=2.78 //y2=0.37
cc_439 ( N_GND_M1_noxref_d N_noxref_18_M1_noxref_s ) capacitor c=0.0334197f \
 //x=3.21 //y=0.87 //x2=2.78 //y2=0.37
cc_440 ( N_GND_c_16_p N_noxref_20_c_4190_n ) capacitor c=0.00500722f //x=38.48 \
 //y=0 //x2=7.13 //y2=1.585
cc_441 ( N_GND_c_23_p N_noxref_20_c_4190_n ) capacitor c=0.00115012f //x=6.645 \
 //y=0 //x2=7.13 //y2=1.585
cc_442 ( N_GND_c_24_p N_noxref_20_c_4190_n ) capacitor c=0.00206628f //x=8.71 \
 //y=0 //x2=7.13 //y2=1.585
cc_443 ( N_GND_M3_noxref_d N_noxref_20_c_4190_n ) capacitor c=0.00902563f \
 //x=6.54 //y=0.87 //x2=7.13 //y2=1.585
cc_444 ( N_GND_c_16_p N_noxref_20_c_4194_n ) capacitor c=0.00242791f //x=38.48 \
 //y=0 //x2=7.215 //y2=0.62
cc_445 ( N_GND_c_24_p N_noxref_20_c_4194_n ) capacitor c=0.0142763f //x=8.71 \
 //y=0 //x2=7.215 //y2=0.62
cc_446 ( N_GND_M3_noxref_d N_noxref_20_c_4194_n ) capacitor c=0.033812f \
 //x=6.54 //y=0.87 //x2=7.215 //y2=0.62
cc_447 ( N_GND_c_4_p N_noxref_20_c_4197_n ) capacitor c=2.91423e-19 //x=5.55 \
 //y=0 //x2=7.215 //y2=1.5
cc_448 ( N_GND_c_16_p N_noxref_20_c_4198_n ) capacitor c=0.010074f //x=38.48 \
 //y=0 //x2=8.1 //y2=0.535
cc_449 ( N_GND_c_24_p N_noxref_20_c_4198_n ) capacitor c=0.0368958f //x=8.71 \
 //y=0 //x2=8.1 //y2=0.535
cc_450 ( N_GND_c_1_p N_noxref_20_c_4198_n ) capacitor c=0.00195382f //x=38.48 \
 //y=0 //x2=8.1 //y2=0.535
cc_451 ( N_GND_c_16_p N_noxref_20_c_4201_n ) capacitor c=0.00242513f //x=38.48 \
 //y=0 //x2=8.185 //y2=0.62
cc_452 ( N_GND_c_24_p N_noxref_20_c_4201_n ) capacitor c=0.0142124f //x=8.71 \
 //y=0 //x2=8.185 //y2=0.62
cc_453 ( N_GND_c_453_p N_noxref_20_c_4201_n ) capacitor c=9.92084e-19 //x=9.5 \
 //y=0.45 //x2=8.185 //y2=0.62
cc_454 ( N_GND_c_5_p N_noxref_20_c_4201_n ) capacitor c=0.0431718f //x=8.88 \
 //y=0 //x2=8.185 //y2=0.62
cc_455 ( N_GND_c_16_p N_noxref_20_M3_noxref_s ) capacitor c=0.00242791f \
 //x=38.48 //y=0 //x2=6.11 //y2=0.37
cc_456 ( N_GND_c_23_p N_noxref_20_M3_noxref_s ) capacitor c=0.0142763f \
 //x=6.645 //y=0 //x2=6.11 //y2=0.37
cc_457 ( N_GND_c_4_p N_noxref_20_M3_noxref_s ) capacitor c=0.058339f //x=5.55 \
 //y=0 //x2=6.11 //y2=0.37
cc_458 ( N_GND_c_5_p N_noxref_20_M3_noxref_s ) capacitor c=0.00200548f \
 //x=8.88 //y=0 //x2=6.11 //y2=0.37
cc_459 ( N_GND_M3_noxref_d N_noxref_20_M3_noxref_s ) capacitor c=0.0334197f \
 //x=6.54 //y=0.87 //x2=6.11 //y2=0.37
cc_460 ( N_GND_M5_noxref_s N_noxref_20_M3_noxref_s ) capacitor c=9.92084e-19 \
 //x=9.375 //y=0.37 //x2=6.11 //y2=0.37
cc_461 ( N_GND_M6_noxref_s N_noxref_22_c_4277_n ) capacitor c=0.0013253f \
 //x=11.595 //y=0.37 //x2=14.015 //y2=1.5
cc_462 ( N_GND_c_16_p N_noxref_22_c_4278_n ) capacitor c=0.00500722f //x=38.48 \
 //y=0 //x2=14.9 //y2=1.585
cc_463 ( N_GND_c_32_p N_noxref_22_c_4278_n ) capacitor c=0.00115012f \
 //x=14.415 //y=0 //x2=14.9 //y2=1.585
cc_464 ( N_GND_c_33_p N_noxref_22_c_4278_n ) capacitor c=0.00206628f //x=16.48 \
 //y=0 //x2=14.9 //y2=1.585
cc_465 ( N_GND_M7_noxref_d N_noxref_22_c_4278_n ) capacitor c=0.00902563f \
 //x=14.31 //y=0.87 //x2=14.9 //y2=1.585
cc_466 ( N_GND_c_16_p N_noxref_22_c_4282_n ) capacitor c=0.00242791f //x=38.48 \
 //y=0 //x2=14.985 //y2=0.62
cc_467 ( N_GND_c_33_p N_noxref_22_c_4282_n ) capacitor c=0.0142763f //x=16.48 \
 //y=0 //x2=14.985 //y2=0.62
cc_468 ( N_GND_M7_noxref_d N_noxref_22_c_4282_n ) capacitor c=0.033812f \
 //x=14.31 //y=0.87 //x2=14.985 //y2=0.62
cc_469 ( N_GND_c_7_p N_noxref_22_c_4285_n ) capacitor c=2.91423e-19 //x=13.32 \
 //y=0 //x2=14.985 //y2=1.5
cc_470 ( N_GND_c_16_p N_noxref_22_c_4286_n ) capacitor c=0.010074f //x=38.48 \
 //y=0 //x2=15.87 //y2=0.535
cc_471 ( N_GND_c_33_p N_noxref_22_c_4286_n ) capacitor c=0.0368958f //x=16.48 \
 //y=0 //x2=15.87 //y2=0.535
cc_472 ( N_GND_c_1_p N_noxref_22_c_4286_n ) capacitor c=0.00195382f //x=38.48 \
 //y=0 //x2=15.87 //y2=0.535
cc_473 ( N_GND_c_16_p N_noxref_22_c_4289_n ) capacitor c=0.00242513f //x=38.48 \
 //y=0 //x2=15.955 //y2=0.62
cc_474 ( N_GND_c_33_p N_noxref_22_c_4289_n ) capacitor c=0.0142124f //x=16.48 \
 //y=0 //x2=15.955 //y2=0.62
cc_475 ( N_GND_c_8_p N_noxref_22_c_4289_n ) capacitor c=0.0431718f //x=16.65 \
 //y=0 //x2=15.955 //y2=0.62
cc_476 ( N_GND_c_16_p N_noxref_22_M7_noxref_s ) capacitor c=0.00242791f \
 //x=38.48 //y=0 //x2=13.88 //y2=0.37
cc_477 ( N_GND_c_477_p N_noxref_22_M7_noxref_s ) capacitor c=0.0013253f \
 //x=12.7 //y=0.45 //x2=13.88 //y2=0.37
cc_478 ( N_GND_c_32_p N_noxref_22_M7_noxref_s ) capacitor c=0.0142763f \
 //x=14.415 //y=0 //x2=13.88 //y2=0.37
cc_479 ( N_GND_c_7_p N_noxref_22_M7_noxref_s ) capacitor c=0.058339f //x=13.32 \
 //y=0 //x2=13.88 //y2=0.37
cc_480 ( N_GND_c_8_p N_noxref_22_M7_noxref_s ) capacitor c=0.00200438f \
 //x=16.65 //y=0 //x2=13.88 //y2=0.37
cc_481 ( N_GND_M7_noxref_d N_noxref_22_M7_noxref_s ) capacitor c=0.0334197f \
 //x=14.31 //y=0.87 //x2=13.88 //y2=0.37
cc_482 ( N_GND_c_16_p N_noxref_24_c_4365_n ) capacitor c=0.00500722f //x=38.48 \
 //y=0 //x2=18.23 //y2=1.585
cc_483 ( N_GND_c_34_p N_noxref_24_c_4365_n ) capacitor c=0.00115012f \
 //x=17.745 //y=0 //x2=18.23 //y2=1.585
cc_484 ( N_GND_c_35_p N_noxref_24_c_4365_n ) capacitor c=0.00206628f //x=19.81 \
 //y=0 //x2=18.23 //y2=1.585
cc_485 ( N_GND_M9_noxref_d N_noxref_24_c_4365_n ) capacitor c=0.00902563f \
 //x=17.64 //y=0.87 //x2=18.23 //y2=1.585
cc_486 ( N_GND_c_16_p N_noxref_24_c_4369_n ) capacitor c=0.00242791f //x=38.48 \
 //y=0 //x2=18.315 //y2=0.62
cc_487 ( N_GND_c_35_p N_noxref_24_c_4369_n ) capacitor c=0.0142763f //x=19.81 \
 //y=0 //x2=18.315 //y2=0.62
cc_488 ( N_GND_M9_noxref_d N_noxref_24_c_4369_n ) capacitor c=0.033812f \
 //x=17.64 //y=0.87 //x2=18.315 //y2=0.62
cc_489 ( N_GND_c_8_p N_noxref_24_c_4372_n ) capacitor c=2.91423e-19 //x=16.65 \
 //y=0 //x2=18.315 //y2=1.5
cc_490 ( N_GND_c_16_p N_noxref_24_c_4373_n ) capacitor c=0.010074f //x=38.48 \
 //y=0 //x2=19.2 //y2=0.535
cc_491 ( N_GND_c_35_p N_noxref_24_c_4373_n ) capacitor c=0.0368958f //x=19.81 \
 //y=0 //x2=19.2 //y2=0.535
cc_492 ( N_GND_c_1_p N_noxref_24_c_4373_n ) capacitor c=0.00195382f //x=38.48 \
 //y=0 //x2=19.2 //y2=0.535
cc_493 ( N_GND_c_16_p N_noxref_24_c_4376_n ) capacitor c=0.00242513f //x=38.48 \
 //y=0 //x2=19.285 //y2=0.62
cc_494 ( N_GND_c_35_p N_noxref_24_c_4376_n ) capacitor c=0.0142124f //x=19.81 \
 //y=0 //x2=19.285 //y2=0.62
cc_495 ( N_GND_c_495_p N_noxref_24_c_4376_n ) capacitor c=9.92084e-19 //x=20.6 \
 //y=0.45 //x2=19.285 //y2=0.62
cc_496 ( N_GND_c_9_p N_noxref_24_c_4376_n ) capacitor c=0.0431718f //x=19.98 \
 //y=0 //x2=19.285 //y2=0.62
cc_497 ( N_GND_c_16_p N_noxref_24_M9_noxref_s ) capacitor c=0.00242791f \
 //x=38.48 //y=0 //x2=17.21 //y2=0.37
cc_498 ( N_GND_c_34_p N_noxref_24_M9_noxref_s ) capacitor c=0.0142763f \
 //x=17.745 //y=0 //x2=17.21 //y2=0.37
cc_499 ( N_GND_c_8_p N_noxref_24_M9_noxref_s ) capacitor c=0.058339f //x=16.65 \
 //y=0 //x2=17.21 //y2=0.37
cc_500 ( N_GND_c_9_p N_noxref_24_M9_noxref_s ) capacitor c=0.00200493f \
 //x=19.98 //y=0 //x2=17.21 //y2=0.37
cc_501 ( N_GND_M9_noxref_d N_noxref_24_M9_noxref_s ) capacitor c=0.0334197f \
 //x=17.64 //y=0.87 //x2=17.21 //y2=0.37
cc_502 ( N_GND_M11_noxref_s N_noxref_24_M9_noxref_s ) capacitor c=9.92084e-19 \
 //x=20.475 //y=0.37 //x2=17.21 //y2=0.37
cc_503 ( N_GND_M11_noxref_s N_noxref_25_c_4415_n ) capacitor c=0.00130619f \
 //x=20.475 //y=0.37 //x2=22.895 //y2=1.495
cc_504 ( N_GND_c_16_p N_noxref_25_c_4416_n ) capacitor c=0.00501918f //x=38.48 \
 //y=0 //x2=23.78 //y2=1.58
cc_505 ( N_GND_c_40_p N_noxref_25_c_4416_n ) capacitor c=0.00115748f \
 //x=23.295 //y=0 //x2=23.78 //y2=1.58
cc_506 ( N_GND_c_41_p N_noxref_25_c_4416_n ) capacitor c=0.0020762f //x=25.36 \
 //y=0 //x2=23.78 //y2=1.58
cc_507 ( N_GND_M12_noxref_d N_noxref_25_c_4416_n ) capacitor c=0.00902889f \
 //x=23.19 //y=0.865 //x2=23.78 //y2=1.58
cc_508 ( N_GND_c_16_p N_noxref_25_c_4420_n ) capacitor c=0.00244876f //x=38.48 \
 //y=0 //x2=23.865 //y2=0.615
cc_509 ( N_GND_c_41_p N_noxref_25_c_4420_n ) capacitor c=0.014581f //x=25.36 \
 //y=0 //x2=23.865 //y2=0.615
cc_510 ( N_GND_M12_noxref_d N_noxref_25_c_4420_n ) capacitor c=0.033812f \
 //x=23.19 //y=0.865 //x2=23.865 //y2=0.615
cc_511 ( N_GND_c_10_p N_noxref_25_c_4423_n ) capacitor c=2.91423e-19 //x=22.2 \
 //y=0 //x2=23.865 //y2=1.495
cc_512 ( N_GND_c_16_p N_noxref_25_c_4424_n ) capacitor c=0.0101349f //x=38.48 \
 //y=0 //x2=24.75 //y2=0.53
cc_513 ( N_GND_c_41_p N_noxref_25_c_4424_n ) capacitor c=0.037368f //x=25.36 \
 //y=0 //x2=24.75 //y2=0.53
cc_514 ( N_GND_c_1_p N_noxref_25_c_4424_n ) capacitor c=0.00199999f //x=38.48 \
 //y=0 //x2=24.75 //y2=0.53
cc_515 ( N_GND_c_16_p N_noxref_25_c_4427_n ) capacitor c=0.00244627f //x=38.48 \
 //y=0 //x2=24.835 //y2=0.615
cc_516 ( N_GND_c_41_p N_noxref_25_c_4427_n ) capacitor c=0.014516f //x=25.36 \
 //y=0 //x2=24.835 //y2=0.615
cc_517 ( N_GND_c_517_p N_noxref_25_c_4427_n ) capacitor c=9.77746e-19 \
 //x=26.16 //y=0.45 //x2=24.835 //y2=0.615
cc_518 ( N_GND_c_11_p N_noxref_25_c_4427_n ) capacitor c=0.0431718f //x=25.53 \
 //y=0 //x2=24.835 //y2=0.615
cc_519 ( N_GND_c_16_p N_noxref_25_M12_noxref_s ) capacitor c=0.00244876f \
 //x=38.48 //y=0 //x2=22.76 //y2=0.365
cc_520 ( N_GND_c_520_p N_noxref_25_M12_noxref_s ) capacitor c=0.00130619f \
 //x=21.57 //y=0.45 //x2=22.76 //y2=0.365
cc_521 ( N_GND_c_40_p N_noxref_25_M12_noxref_s ) capacitor c=0.014581f \
 //x=23.295 //y=0 //x2=22.76 //y2=0.365
cc_522 ( N_GND_c_10_p N_noxref_25_M12_noxref_s ) capacitor c=0.058339f \
 //x=22.2 //y=0 //x2=22.76 //y2=0.365
cc_523 ( N_GND_c_11_p N_noxref_25_M12_noxref_s ) capacitor c=0.00198098f \
 //x=25.53 //y=0 //x2=22.76 //y2=0.365
cc_524 ( N_GND_M12_noxref_d N_noxref_25_M12_noxref_s ) capacitor c=0.0334197f \
 //x=23.19 //y=0.865 //x2=22.76 //y2=0.365
cc_525 ( N_GND_M14_noxref_s N_noxref_25_M12_noxref_s ) capacitor c=9.77746e-19 \
 //x=26.025 //y=0.37 //x2=22.76 //y2=0.365
cc_526 ( N_GND_M14_noxref_s N_noxref_26_c_4468_n ) capacitor c=0.0013253f \
 //x=26.025 //y=0.37 //x2=28.445 //y2=1.495
cc_527 ( N_GND_c_16_p N_noxref_26_c_4469_n ) capacitor c=0.00501918f //x=38.48 \
 //y=0 //x2=29.33 //y2=1.58
cc_528 ( N_GND_c_45_p N_noxref_26_c_4469_n ) capacitor c=0.00115748f \
 //x=28.845 //y=0 //x2=29.33 //y2=1.58
cc_529 ( N_GND_c_46_p N_noxref_26_c_4469_n ) capacitor c=0.0020762f //x=30.91 \
 //y=0 //x2=29.33 //y2=1.58
cc_530 ( N_GND_M15_noxref_d N_noxref_26_c_4469_n ) capacitor c=0.00902889f \
 //x=28.74 //y=0.865 //x2=29.33 //y2=1.58
cc_531 ( N_GND_c_16_p N_noxref_26_c_4473_n ) capacitor c=0.00244876f //x=38.48 \
 //y=0 //x2=29.415 //y2=0.615
cc_532 ( N_GND_c_46_p N_noxref_26_c_4473_n ) capacitor c=0.0142704f //x=30.91 \
 //y=0 //x2=29.415 //y2=0.615
cc_533 ( N_GND_M15_noxref_d N_noxref_26_c_4473_n ) capacitor c=0.033812f \
 //x=28.74 //y=0.865 //x2=29.415 //y2=0.615
cc_534 ( N_GND_c_12_p N_noxref_26_c_4476_n ) capacitor c=2.91423e-19 //x=27.75 \
 //y=0 //x2=29.415 //y2=1.495
cc_535 ( N_GND_c_16_p N_noxref_26_c_4477_n ) capacitor c=0.0112457f //x=38.48 \
 //y=0 //x2=30.3 //y2=0.53
cc_536 ( N_GND_c_46_p N_noxref_26_c_4477_n ) capacitor c=0.0374193f //x=30.91 \
 //y=0 //x2=30.3 //y2=0.53
cc_537 ( N_GND_c_1_p N_noxref_26_c_4477_n ) capacitor c=0.00199999f //x=38.48 \
 //y=0 //x2=30.3 //y2=0.53
cc_538 ( N_GND_c_16_p N_noxref_26_c_4480_n ) capacitor c=0.00282863f //x=38.48 \
 //y=0 //x2=30.385 //y2=0.615
cc_539 ( N_GND_c_46_p N_noxref_26_c_4480_n ) capacitor c=0.0148003f //x=30.91 \
 //y=0 //x2=30.385 //y2=0.615
cc_540 ( N_GND_c_540_p N_noxref_26_c_4480_n ) capacitor c=9.77746e-19 \
 //x=31.71 //y=0.45 //x2=30.385 //y2=0.615
cc_541 ( N_GND_c_13_p N_noxref_26_c_4480_n ) capacitor c=0.0431718f //x=31.08 \
 //y=0 //x2=30.385 //y2=0.615
cc_542 ( N_GND_c_16_p N_noxref_26_M15_noxref_s ) capacitor c=0.00244876f \
 //x=38.48 //y=0 //x2=28.31 //y2=0.365
cc_543 ( N_GND_c_543_p N_noxref_26_M15_noxref_s ) capacitor c=0.0013253f \
 //x=27.13 //y=0.45 //x2=28.31 //y2=0.365
cc_544 ( N_GND_c_45_p N_noxref_26_M15_noxref_s ) capacitor c=0.014581f \
 //x=28.845 //y=0 //x2=28.31 //y2=0.365
cc_545 ( N_GND_c_12_p N_noxref_26_M15_noxref_s ) capacitor c=0.058339f \
 //x=27.75 //y=0 //x2=28.31 //y2=0.365
cc_546 ( N_GND_c_13_p N_noxref_26_M15_noxref_s ) capacitor c=0.00198098f \
 //x=31.08 //y=0 //x2=28.31 //y2=0.365
cc_547 ( N_GND_M15_noxref_d N_noxref_26_M15_noxref_s ) capacitor c=0.0334197f \
 //x=28.74 //y=0.865 //x2=28.31 //y2=0.365
cc_548 ( N_GND_M17_noxref_s N_noxref_26_M15_noxref_s ) capacitor c=9.77746e-19 \
 //x=31.575 //y=0.37 //x2=28.31 //y2=0.365
cc_549 ( N_GND_c_15_p COUT ) capacitor c=8.10282e-19 //x=36.63 //y=0 \
 //x2=38.11 //y2=2.22
cc_550 ( N_GND_c_16_p N_COUT_c_4568_n ) capacitor c=0.00180637f //x=38.48 \
 //y=0 //x2=38.025 //y2=2.08
cc_551 ( N_GND_c_1_p N_COUT_c_4568_n ) capacitor c=0.0301661f //x=38.48 //y=0 \
 //x2=38.025 //y2=2.08
cc_552 ( N_GND_M20_noxref_s N_COUT_c_4568_n ) capacitor c=0.00999304f \
 //x=37.125 //y=0.37 //x2=38.025 //y2=2.08
cc_553 ( N_GND_c_16_p N_COUT_M20_noxref_d ) capacitor c=0.00194883f //x=38.48 \
 //y=0 //x2=37.555 //y2=0.91
cc_554 ( N_GND_c_381_p N_COUT_M20_noxref_d ) capacitor c=0.0146043f //x=37.66 \
 //y=0.535 //x2=37.555 //y2=0.91
cc_555 ( N_GND_c_1_p N_COUT_M20_noxref_d ) capacitor c=0.00950831f //x=38.48 \
 //y=0 //x2=37.555 //y2=0.91
cc_556 ( N_GND_c_15_p N_COUT_M20_noxref_d ) capacitor c=0.00924905f //x=36.63 \
 //y=0 //x2=37.555 //y2=0.91
cc_557 ( N_GND_M20_noxref_s N_COUT_M20_noxref_d ) capacitor c=0.076995f \
 //x=37.125 //y=0.37 //x2=37.555 //y2=0.91
cc_558 ( N_VDD_c_573_p N_A_c_1088_n ) capacitor c=0.0179155f //x=38.48 //y=7.4 \
 //x2=3.215 //y2=4.07
cc_559 ( N_VDD_c_574_p N_A_c_1088_n ) capacitor c=9.77842e-19 //x=1.47 //y=7.4 \
 //x2=3.215 //y2=4.07
cc_560 ( N_VDD_c_575_p N_A_c_1088_n ) capacitor c=0.00124367f //x=2.05 //y=7.4 \
 //x2=3.215 //y2=4.07
cc_561 ( N_VDD_c_576_p N_A_c_1088_n ) capacitor c=0.00216965f //x=3.365 \
 //y=7.4 //x2=3.215 //y2=4.07
cc_562 ( N_VDD_c_560_n N_A_c_1088_n ) capacitor c=0.0280406f //x=2.22 //y=7.4 \
 //x2=3.215 //y2=4.07
cc_563 ( N_VDD_M22_noxref_d N_A_c_1088_n ) capacitor c=0.00213856f //x=1.41 \
 //y=5.02 //x2=3.215 //y2=4.07
cc_564 ( N_VDD_c_573_p N_A_c_1090_n ) capacitor c=0.00188164f //x=38.48 \
 //y=7.4 //x2=0.855 //y2=4.07
cc_565 ( N_VDD_c_559_n N_A_c_1090_n ) capacitor c=0.00208272f //x=0.74 //y=7.4 \
 //x2=0.855 //y2=4.07
cc_566 ( N_VDD_M21_noxref_s N_A_c_1090_n ) capacitor c=0.00185024f //x=0.54 \
 //y=5.02 //x2=0.855 //y2=4.07
cc_567 ( N_VDD_c_560_n A ) capacitor c=0.0156437f //x=2.22 //y=7.4 //x2=3.33 \
 //y2=2.96
cc_568 ( N_VDD_c_569_n A ) capacitor c=7.46601e-19 //x=27.75 //y=7.4 //x2=29.6 \
 //y2=2.59
cc_569 ( N_VDD_c_570_n A ) capacitor c=6.80078e-19 //x=31.08 //y=7.4 //x2=29.6 \
 //y2=2.59
cc_570 ( N_VDD_M23_noxref_d A ) capacitor c=3.16761e-19 //x=3.305 //y=5.02 \
 //x2=3.33 //y2=2.22
cc_571 ( N_VDD_M52_noxref_d A ) capacitor c=2.91389e-19 //x=29.275 //y=5.02 \
 //x2=29.6 //y2=2.22
cc_572 ( N_VDD_c_573_p N_A_c_1142_n ) capacitor c=0.00157744f //x=38.48 \
 //y=7.4 //x2=0.74 //y2=2.085
cc_573 ( N_VDD_c_559_n N_A_c_1142_n ) capacitor c=0.0272385f //x=0.74 //y=7.4 \
 //x2=0.74 //y2=2.085
cc_574 ( N_VDD_c_560_n N_A_c_1142_n ) capacitor c=0.00139956f //x=2.22 //y=7.4 \
 //x2=0.74 //y2=2.085
cc_575 ( N_VDD_M21_noxref_s N_A_c_1142_n ) capacitor c=0.00896093f //x=0.54 \
 //y=5.02 //x2=0.74 //y2=2.085
cc_576 ( N_VDD_c_574_p N_A_M21_noxref_g ) capacitor c=0.00748034f //x=1.47 \
 //y=7.4 //x2=0.895 //y2=6.02
cc_577 ( N_VDD_c_559_n N_A_M21_noxref_g ) capacitor c=0.0241676f //x=0.74 \
 //y=7.4 //x2=0.895 //y2=6.02
cc_578 ( N_VDD_M21_noxref_s N_A_M21_noxref_g ) capacitor c=0.0528676f //x=0.54 \
 //y=5.02 //x2=0.895 //y2=6.02
cc_579 ( N_VDD_c_574_p N_A_M22_noxref_g ) capacitor c=0.00697478f //x=1.47 \
 //y=7.4 //x2=1.335 //y2=6.02
cc_580 ( N_VDD_M22_noxref_d N_A_M22_noxref_g ) capacitor c=0.0528676f //x=1.41 \
 //y=5.02 //x2=1.335 //y2=6.02
cc_581 ( N_VDD_c_576_p N_A_M23_noxref_g ) capacitor c=0.00673447f //x=3.365 \
 //y=7.4 //x2=3.23 //y2=6.02
cc_582 ( N_VDD_c_560_n N_A_M23_noxref_g ) capacitor c=0.00449901f //x=2.22 \
 //y=7.4 //x2=3.23 //y2=6.02
cc_583 ( N_VDD_M23_noxref_d N_A_M23_noxref_g ) capacitor c=0.0166176f \
 //x=3.305 //y=5.02 //x2=3.23 //y2=6.02
cc_584 ( N_VDD_c_599_p N_A_M24_noxref_g ) capacitor c=0.006727f //x=5.38 \
 //y=7.4 //x2=3.67 //y2=6.02
cc_585 ( N_VDD_M23_noxref_d N_A_M24_noxref_g ) capacitor c=0.0186652f \
 //x=3.305 //y=5.02 //x2=3.67 //y2=6.02
cc_586 ( N_VDD_c_601_p N_A_M53_noxref_g ) capacitor c=0.00673971f //x=30.215 \
 //y=7.4 //x2=29.64 //y2=6.02
cc_587 ( N_VDD_M52_noxref_d N_A_M53_noxref_g ) capacitor c=0.015318f \
 //x=29.275 //y=5.02 //x2=29.64 //y2=6.02
cc_588 ( N_VDD_c_601_p N_A_M54_noxref_g ) capacitor c=0.00672952f //x=30.215 \
 //y=7.4 //x2=30.08 //y2=6.02
cc_589 ( N_VDD_c_570_n N_A_M54_noxref_g ) capacitor c=0.00886951f //x=31.08 \
 //y=7.4 //x2=30.08 //y2=6.02
cc_590 ( N_VDD_M54_noxref_d N_A_M54_noxref_g ) capacitor c=0.0430452f \
 //x=30.155 //y=5.02 //x2=30.08 //y2=6.02
cc_591 ( N_VDD_c_560_n N_A_c_1199_n ) capacitor c=0.0132667f //x=2.22 //y=7.4 \
 //x2=1.26 //y2=4.79
cc_592 ( N_VDD_c_559_n N_A_c_1200_n ) capacitor c=0.011132f //x=0.74 //y=7.4 \
 //x2=0.97 //y2=4.79
cc_593 ( N_VDD_M21_noxref_s N_A_c_1200_n ) capacitor c=0.00524527f //x=0.54 \
 //y=5.02 //x2=0.97 //y2=4.79
cc_594 ( N_VDD_c_560_n N_A_c_1202_n ) capacitor c=0.0125867f //x=2.22 //y=7.4 \
 //x2=3.33 //y2=4.7
cc_595 ( N_VDD_c_560_n N_noxref_4_c_1465_n ) capacitor c=0.00137387f //x=2.22 \
 //y=7.4 //x2=7.655 //y2=2.59
cc_596 ( N_VDD_c_573_p N_noxref_4_c_1488_n ) capacitor c=0.0012271f //x=38.48 \
 //y=7.4 //x2=1.395 //y2=4.58
cc_597 ( N_VDD_c_574_p N_noxref_4_c_1488_n ) capacitor c=9.08147e-19 //x=1.47 \
 //y=7.4 //x2=1.395 //y2=4.58
cc_598 ( N_VDD_M22_noxref_d N_noxref_4_c_1488_n ) capacitor c=0.00609088f \
 //x=1.41 //y=5.02 //x2=1.395 //y2=4.58
cc_599 ( N_VDD_c_559_n N_noxref_4_c_1491_n ) capacitor c=0.0179238f //x=0.74 \
 //y=7.4 //x2=1.2 //y2=4.58
cc_600 ( N_VDD_c_559_n N_noxref_4_c_1477_n ) capacitor c=5.65246e-19 //x=0.74 \
 //y=7.4 //x2=1.48 //y2=2.59
cc_601 ( N_VDD_c_560_n N_noxref_4_c_1477_n ) capacitor c=0.0220651f //x=2.22 \
 //y=7.4 //x2=1.48 //y2=2.59
cc_602 ( N_VDD_c_561_n N_noxref_4_c_1480_n ) capacitor c=0.00210246f //x=5.55 \
 //y=7.4 //x2=7.77 //y2=2.085
cc_603 ( N_VDD_c_562_n N_noxref_4_c_1480_n ) capacitor c=0.00147528f //x=8.88 \
 //y=7.4 //x2=7.77 //y2=2.085
cc_604 ( N_VDD_c_619_p N_noxref_4_M29_noxref_g ) capacitor c=0.00510247f \
 //x=8.71 //y=7.4 //x2=7.44 //y2=6.02
cc_605 ( N_VDD_c_619_p N_noxref_4_M30_noxref_g ) capacitor c=0.00510919f \
 //x=8.71 //y=7.4 //x2=7.88 //y2=6.02
cc_606 ( N_VDD_c_562_n N_noxref_4_M30_noxref_g ) capacitor c=0.00788519f \
 //x=8.88 //y=7.4 //x2=7.88 //y2=6.02
cc_607 ( N_VDD_c_573_p N_noxref_4_M21_noxref_d ) capacitor c=0.00285171f \
 //x=38.48 //y=7.4 //x2=0.97 //y2=5.02
cc_608 ( N_VDD_c_574_p N_noxref_4_M21_noxref_d ) capacitor c=0.0141332f \
 //x=1.47 //y=7.4 //x2=0.97 //y2=5.02
cc_609 ( N_VDD_c_560_n N_noxref_4_M21_noxref_d ) capacitor c=0.0204646f \
 //x=2.22 //y=7.4 //x2=0.97 //y2=5.02
cc_610 ( N_VDD_M21_noxref_s N_noxref_4_M21_noxref_d ) capacitor c=0.0843065f \
 //x=0.54 //y=5.02 //x2=0.97 //y2=5.02
cc_611 ( N_VDD_M22_noxref_d N_noxref_4_M21_noxref_d ) capacitor c=0.0832641f \
 //x=1.41 //y=5.02 //x2=0.97 //y2=5.02
cc_612 ( N_VDD_c_573_p N_noxref_5_c_1646_n ) capacitor c=0.0245984f //x=38.48 \
 //y=7.4 //x2=9.505 //y2=4.07
cc_613 ( N_VDD_c_599_p N_noxref_5_c_1646_n ) capacitor c=0.00187833f //x=5.38 \
 //y=7.4 //x2=9.505 //y2=4.07
cc_614 ( N_VDD_c_629_p N_noxref_5_c_1646_n ) capacitor c=0.00213804f //x=6.695 \
 //y=7.4 //x2=9.505 //y2=4.07
cc_615 ( N_VDD_c_561_n N_noxref_5_c_1646_n ) capacitor c=0.0272145f //x=5.55 \
 //y=7.4 //x2=9.505 //y2=4.07
cc_616 ( N_VDD_c_562_n N_noxref_5_c_1646_n ) capacitor c=0.0144842f //x=8.88 \
 //y=7.4 //x2=9.505 //y2=4.07
cc_617 ( N_VDD_c_573_p N_noxref_5_c_1651_n ) capacitor c=0.00164816f //x=38.48 \
 //y=7.4 //x2=4.555 //y2=4.07
cc_618 ( N_VDD_c_560_n N_noxref_5_c_1652_n ) capacitor c=7.20931e-19 //x=2.22 \
 //y=7.4 //x2=4.44 //y2=4.07
cc_619 ( N_VDD_c_561_n N_noxref_5_c_1652_n ) capacitor c=0.00211919f //x=5.55 \
 //y=7.4 //x2=4.44 //y2=4.07
cc_620 ( N_VDD_c_562_n N_noxref_5_c_1627_n ) capacitor c=0.0195526f //x=8.88 \
 //y=7.4 //x2=9.62 //y2=3.33
cc_621 ( N_VDD_c_563_n N_noxref_5_c_1627_n ) capacitor c=6.39704e-19 //x=11.1 \
 //y=7.4 //x2=9.62 //y2=3.33
cc_622 ( N_VDD_c_563_n N_noxref_5_c_1656_n ) capacitor c=0.015474f //x=11.1 \
 //y=7.4 //x2=9.9 //y2=4.58
cc_623 ( N_VDD_c_573_p N_noxref_5_c_1657_n ) capacitor c=0.00119381f //x=38.48 \
 //y=7.4 //x2=9.705 //y2=4.58
cc_624 ( N_VDD_c_639_p N_noxref_5_c_1657_n ) capacitor c=0.0010061f //x=10.34 \
 //y=7.4 //x2=9.705 //y2=4.58
cc_625 ( N_VDD_M31_noxref_s N_noxref_5_c_1657_n ) capacitor c=0.00562155f \
 //x=9.42 //y=5.02 //x2=9.705 //y2=4.58
cc_626 ( N_VDD_c_599_p N_noxref_5_M25_noxref_g ) capacitor c=0.00510247f \
 //x=5.38 //y=7.4 //x2=4.11 //y2=6.02
cc_627 ( N_VDD_c_599_p N_noxref_5_M26_noxref_g ) capacitor c=0.00510919f \
 //x=5.38 //y=7.4 //x2=4.55 //y2=6.02
cc_628 ( N_VDD_c_561_n N_noxref_5_M26_noxref_g ) capacitor c=0.0122307f \
 //x=5.55 //y=7.4 //x2=4.55 //y2=6.02
cc_629 ( N_VDD_c_573_p N_noxref_5_M31_noxref_d ) capacitor c=0.00275339f \
 //x=38.48 //y=7.4 //x2=9.84 //y2=5.02
cc_630 ( N_VDD_c_639_p N_noxref_5_M31_noxref_d ) capacitor c=0.0140667f \
 //x=10.34 //y=7.4 //x2=9.84 //y2=5.02
cc_631 ( N_VDD_c_562_n N_noxref_5_M31_noxref_d ) capacitor c=0.019987f \
 //x=8.88 //y=7.4 //x2=9.84 //y2=5.02
cc_632 ( N_VDD_M31_noxref_s N_noxref_5_M31_noxref_d ) capacitor c=0.0832641f \
 //x=9.42 //y=5.02 //x2=9.84 //y2=5.02
cc_633 ( N_VDD_M32_noxref_d N_noxref_5_M31_noxref_d ) capacitor c=0.0843065f \
 //x=10.28 //y=5.02 //x2=9.84 //y2=5.02
cc_634 ( N_VDD_c_573_p N_B_c_1830_n ) capacitor c=0.0233843f //x=38.48 //y=7.4 \
 //x2=10.245 //y2=4.44
cc_635 ( N_VDD_c_619_p N_B_c_1830_n ) capacitor c=0.00304371f //x=8.71 //y=7.4 \
 //x2=10.245 //y2=4.44
cc_636 ( N_VDD_c_651_p N_B_c_1830_n ) capacitor c=0.00151604f //x=9.46 //y=7.4 \
 //x2=10.245 //y2=4.44
cc_637 ( N_VDD_c_639_p N_B_c_1830_n ) capacitor c=0.00156466f //x=10.34 \
 //y=7.4 //x2=10.245 //y2=4.44
cc_638 ( N_VDD_c_562_n N_B_c_1830_n ) capacitor c=0.0377357f //x=8.88 //y=7.4 \
 //x2=10.245 //y2=4.44
cc_639 ( N_VDD_c_563_n N_B_c_1830_n ) capacitor c=0.00909033f //x=11.1 //y=7.4 \
 //x2=10.245 //y2=4.44
cc_640 ( N_VDD_M31_noxref_s N_B_c_1830_n ) capacitor c=0.00317238f //x=9.42 \
 //y=5.02 //x2=10.245 //y2=4.44
cc_641 ( N_VDD_c_573_p N_B_c_1837_n ) capacitor c=0.00150124f //x=38.48 \
 //y=7.4 //x2=6.775 //y2=4.44
cc_642 ( N_VDD_c_561_n N_B_c_1837_n ) capacitor c=0.00665137f //x=5.55 //y=7.4 \
 //x2=6.775 //y2=4.44
cc_643 ( N_VDD_c_573_p N_B_c_1839_n ) capacitor c=0.151266f //x=38.48 //y=7.4 \
 //x2=28.745 //y2=4.81
cc_644 ( N_VDD_c_659_p N_B_c_1839_n ) capacitor c=0.00188643f //x=10.93 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_645 ( N_VDD_c_660_p N_B_c_1839_n ) capacitor c=0.00188643f //x=11.69 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_646 ( N_VDD_c_661_p N_B_c_1839_n ) capacitor c=0.00423504f //x=12.57 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_647 ( N_VDD_c_662_p N_B_c_1839_n ) capacitor c=0.00182748f //x=13.15 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_648 ( N_VDD_c_663_p N_B_c_1839_n ) capacitor c=0.00330958f //x=14.465 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_649 ( N_VDD_c_664_p N_B_c_1839_n ) capacitor c=0.00395021f //x=16.48 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_650 ( N_VDD_c_665_p N_B_c_1839_n ) capacitor c=0.00330958f //x=17.795 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_651 ( N_VDD_c_666_p N_B_c_1839_n ) capacitor c=0.00395021f //x=19.81 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_652 ( N_VDD_c_667_p N_B_c_1839_n ) capacitor c=0.00182748f //x=20.56 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_653 ( N_VDD_c_668_p N_B_c_1839_n ) capacitor c=0.00423504f //x=21.44 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_654 ( N_VDD_c_669_p N_B_c_1839_n ) capacitor c=0.00188643f //x=22.03 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_655 ( N_VDD_c_670_p N_B_c_1839_n ) capacitor c=0.00252442f //x=22.905 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_656 ( N_VDD_c_671_p N_B_c_1839_n ) capacitor c=0.00240512f //x=23.785 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_657 ( N_VDD_c_672_p N_B_c_1839_n ) capacitor c=0.00250541f //x=25.36 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_658 ( N_VDD_c_673_p N_B_c_1839_n ) capacitor c=0.00188643f //x=26.12 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_659 ( N_VDD_c_674_p N_B_c_1839_n ) capacitor c=0.00423504f //x=27 //y=7.4 \
 //x2=28.745 //y2=4.81
cc_660 ( N_VDD_c_675_p N_B_c_1839_n ) capacitor c=0.00182748f //x=27.58 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_661 ( N_VDD_c_676_p N_B_c_1839_n ) capacitor c=0.00252442f //x=28.455 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_662 ( N_VDD_c_677_p N_B_c_1839_n ) capacitor c=9.57335e-19 //x=29.335 \
 //y=7.4 //x2=28.745 //y2=4.81
cc_663 ( N_VDD_c_563_n N_B_c_1839_n ) capacitor c=0.0426633f //x=11.1 //y=7.4 \
 //x2=28.745 //y2=4.81
cc_664 ( N_VDD_c_564_n N_B_c_1839_n ) capacitor c=0.0446978f //x=13.32 //y=7.4 \
 //x2=28.745 //y2=4.81
cc_665 ( N_VDD_c_565_n N_B_c_1839_n ) capacitor c=0.0434624f //x=16.65 //y=7.4 \
 //x2=28.745 //y2=4.81
cc_666 ( N_VDD_c_566_n N_B_c_1839_n ) capacitor c=0.0385849f //x=19.98 //y=7.4 \
 //x2=28.745 //y2=4.81
cc_667 ( N_VDD_c_567_n N_B_c_1839_n ) capacitor c=0.0390057f //x=22.2 //y=7.4 \
 //x2=28.745 //y2=4.81
cc_668 ( N_VDD_c_568_n N_B_c_1839_n ) capacitor c=0.0438666f //x=25.53 //y=7.4 \
 //x2=28.745 //y2=4.81
cc_669 ( N_VDD_c_569_n N_B_c_1839_n ) capacitor c=0.0469639f //x=27.75 //y=7.4 \
 //x2=28.745 //y2=4.81
cc_670 ( N_VDD_M32_noxref_d N_B_c_1839_n ) capacitor c=0.00151586f //x=10.28 \
 //y=5.02 //x2=28.745 //y2=4.81
cc_671 ( N_VDD_M33_noxref_s N_B_c_1839_n ) capacitor c=0.00535916f //x=11.64 \
 //y=5.02 //x2=28.745 //y2=4.81
cc_672 ( N_VDD_M34_noxref_d N_B_c_1839_n ) capacitor c=0.00579106f //x=12.51 \
 //y=5.02 //x2=28.745 //y2=4.81
cc_673 ( N_VDD_M43_noxref_s N_B_c_1839_n ) capacitor c=0.00579106f //x=20.52 \
 //y=5.02 //x2=28.745 //y2=4.81
cc_674 ( N_VDD_M44_noxref_d N_B_c_1839_n ) capacitor c=0.00535916f //x=21.38 \
 //y=5.02 //x2=28.745 //y2=4.81
cc_675 ( N_VDD_M45_noxref_s N_B_c_1839_n ) capacitor c=0.00789822f //x=22.855 \
 //y=5.02 //x2=28.745 //y2=4.81
cc_676 ( N_VDD_M48_noxref_d N_B_c_1839_n ) capacitor c=9.73959e-19 //x=24.605 \
 //y=5.02 //x2=28.745 //y2=4.81
cc_677 ( N_VDD_M49_noxref_s N_B_c_1839_n ) capacitor c=0.00535916f //x=26.07 \
 //y=5.02 //x2=28.745 //y2=4.81
cc_678 ( N_VDD_M50_noxref_d N_B_c_1839_n ) capacitor c=0.00579106f //x=26.94 \
 //y=5.02 //x2=28.745 //y2=4.81
cc_679 ( N_VDD_M51_noxref_s N_B_c_1839_n ) capacitor c=0.00789822f //x=28.405 \
 //y=5.02 //x2=28.745 //y2=4.81
cc_680 ( N_VDD_c_573_p N_B_c_1876_n ) capacitor c=0.00205675f //x=38.48 \
 //y=7.4 //x2=10.475 //y2=4.81
cc_681 ( N_VDD_c_639_p N_B_c_1876_n ) capacitor c=7.65571e-19 //x=10.34 \
 //y=7.4 //x2=10.475 //y2=4.81
cc_682 ( N_VDD_c_563_n N_B_c_1876_n ) capacitor c=0.00172533f //x=11.1 //y=7.4 \
 //x2=10.475 //y2=4.81
cc_683 ( N_VDD_M32_noxref_d N_B_c_1876_n ) capacitor c=0.00291231f //x=10.28 \
 //y=5.02 //x2=10.475 //y2=4.81
cc_684 ( N_VDD_c_677_p N_B_c_1880_n ) capacitor c=4.01696e-19 //x=29.335 \
 //y=7.4 //x2=28.86 //y2=4.63
cc_685 ( N_VDD_c_569_n N_B_c_1880_n ) capacitor c=0.00164027f //x=27.75 \
 //y=7.4 //x2=28.86 //y2=4.63
cc_686 ( N_VDD_c_561_n B ) capacitor c=0.0112651f //x=5.55 //y=7.4 //x2=6.66 \
 //y2=4.44
cc_687 ( N_VDD_c_573_p B ) capacitor c=7.93687e-19 //x=38.48 //y=7.4 \
 //x2=28.86 //y2=4.81
cc_688 ( N_VDD_c_569_n B ) capacitor c=0.00693555f //x=27.75 //y=7.4 \
 //x2=28.86 //y2=4.81
cc_689 ( N_VDD_c_573_p N_B_c_1805_n ) capacitor c=6.77658e-19 //x=38.48 \
 //y=7.4 //x2=10.36 //y2=2.085
cc_690 ( N_VDD_c_562_n N_B_c_1805_n ) capacitor c=0.00101567f //x=8.88 //y=7.4 \
 //x2=10.36 //y2=2.085
cc_691 ( N_VDD_c_563_n N_B_c_1805_n ) capacitor c=0.0269017f //x=11.1 //y=7.4 \
 //x2=10.36 //y2=2.085
cc_692 ( N_VDD_M32_noxref_d N_B_c_1805_n ) capacitor c=0.0143271f //x=10.28 \
 //y=5.02 //x2=10.36 //y2=2.085
cc_693 ( N_VDD_c_569_n N_B_c_1810_n ) capacitor c=0.00989948f //x=27.75 \
 //y=7.4 //x2=28.86 //y2=2.08
cc_694 ( N_VDD_c_629_p N_B_M27_noxref_g ) capacitor c=0.00673447f //x=6.695 \
 //y=7.4 //x2=6.56 //y2=6.02
cc_695 ( N_VDD_c_561_n N_B_M27_noxref_g ) capacitor c=0.00661226f //x=5.55 \
 //y=7.4 //x2=6.56 //y2=6.02
cc_696 ( N_VDD_M27_noxref_d N_B_M27_noxref_g ) capacitor c=0.0166176f \
 //x=6.635 //y=5.02 //x2=6.56 //y2=6.02
cc_697 ( N_VDD_c_619_p N_B_M28_noxref_g ) capacitor c=0.006727f //x=8.71 \
 //y=7.4 //x2=7 //y2=6.02
cc_698 ( N_VDD_M27_noxref_d N_B_M28_noxref_g ) capacitor c=0.0186652f \
 //x=6.635 //y=5.02 //x2=7 //y2=6.02
cc_699 ( N_VDD_c_639_p N_B_M31_noxref_g ) capacitor c=0.00697478f //x=10.34 \
 //y=7.4 //x2=9.765 //y2=6.02
cc_700 ( N_VDD_M31_noxref_s N_B_M31_noxref_g ) capacitor c=0.0528676f //x=9.42 \
 //y=5.02 //x2=9.765 //y2=6.02
cc_701 ( N_VDD_c_639_p N_B_M32_noxref_g ) capacitor c=0.00748009f //x=10.34 \
 //y=7.4 //x2=10.205 //y2=6.02
cc_702 ( N_VDD_c_563_n N_B_M32_noxref_g ) capacitor c=0.00563775f //x=11.1 \
 //y=7.4 //x2=10.205 //y2=6.02
cc_703 ( N_VDD_M32_noxref_d N_B_M32_noxref_g ) capacitor c=0.0528676f \
 //x=10.28 //y=5.02 //x2=10.205 //y2=6.02
cc_704 ( N_VDD_c_677_p N_B_M51_noxref_g ) capacitor c=0.00697794f //x=29.335 \
 //y=7.4 //x2=28.76 //y2=6.02
cc_705 ( N_VDD_M51_noxref_s N_B_M51_noxref_g ) capacitor c=0.054195f \
 //x=28.405 //y=5.02 //x2=28.76 //y2=6.02
cc_706 ( N_VDD_c_677_p N_B_M52_noxref_g ) capacitor c=0.00672952f //x=29.335 \
 //y=7.4 //x2=29.2 //y2=6.02
cc_707 ( N_VDD_M52_noxref_d N_B_M52_noxref_g ) capacitor c=0.015318f \
 //x=29.275 //y=5.02 //x2=29.2 //y2=6.02
cc_708 ( N_VDD_c_562_n N_B_c_1904_n ) capacitor c=0.0133962f //x=8.88 //y=7.4 \
 //x2=9.84 //y2=4.79
cc_709 ( N_VDD_c_563_n N_B_c_1905_n ) capacitor c=0.00683901f //x=11.1 //y=7.4 \
 //x2=10.205 //y2=4.865
cc_710 ( N_VDD_M32_noxref_d N_B_c_1905_n ) capacitor c=0.0034545f //x=10.28 \
 //y=5.02 //x2=10.205 //y2=4.865
cc_711 ( N_VDD_c_561_n N_B_c_1907_n ) capacitor c=0.0124704f //x=5.55 //y=7.4 \
 //x2=6.66 //y2=4.7
cc_712 ( N_VDD_c_569_n N_B_c_1908_n ) capacitor c=0.0067953f //x=27.75 //y=7.4 \
 //x2=28.86 //y2=4.7
cc_713 ( N_VDD_c_563_n N_noxref_7_c_2182_n ) capacitor c=0.00788535f //x=11.1 \
 //y=7.4 //x2=11.725 //y2=3.7
cc_714 ( N_VDD_c_567_n N_noxref_7_c_2183_n ) capacitor c=0.00148115f //x=22.2 \
 //y=7.4 //x2=23.935 //y2=2.22
cc_715 ( N_VDD_c_564_n N_noxref_7_c_2188_n ) capacitor c=0.0198302f //x=13.32 \
 //y=7.4 //x2=14.315 //y2=4.07
cc_716 ( N_VDD_c_563_n N_noxref_7_c_2230_n ) capacitor c=0.00156497f //x=11.1 \
 //y=7.4 //x2=11.955 //y2=4.07
cc_717 ( N_VDD_c_573_p N_noxref_7_c_2231_n ) capacitor c=0.00114115f //x=38.48 \
 //y=7.4 //x2=4.725 //y2=5.205
cc_718 ( N_VDD_c_599_p N_noxref_7_c_2231_n ) capacitor c=0.00139027f //x=5.38 \
 //y=7.4 //x2=4.725 //y2=5.205
cc_719 ( N_VDD_c_560_n N_noxref_7_c_2233_n ) capacitor c=8.9933e-19 //x=2.22 \
 //y=7.4 //x2=4.415 //y2=5.205
cc_720 ( N_VDD_c_560_n N_noxref_7_c_2190_n ) capacitor c=0.00163766f //x=2.22 \
 //y=7.4 //x2=4.81 //y2=3.7
cc_721 ( N_VDD_c_561_n N_noxref_7_c_2190_n ) capacitor c=0.0445615f //x=5.55 \
 //y=7.4 //x2=4.81 //y2=3.7
cc_722 ( N_VDD_c_573_p N_noxref_7_c_2236_n ) capacitor c=0.00113725f //x=38.48 \
 //y=7.4 //x2=8.055 //y2=5.205
cc_723 ( N_VDD_c_619_p N_noxref_7_c_2236_n ) capacitor c=0.00138968f //x=8.71 \
 //y=7.4 //x2=8.055 //y2=5.205
cc_724 ( N_VDD_c_561_n N_noxref_7_c_2238_n ) capacitor c=8.9933e-19 //x=5.55 \
 //y=7.4 //x2=7.745 //y2=5.205
cc_725 ( N_VDD_c_561_n N_noxref_7_c_2239_n ) capacitor c=0.00177938f //x=5.55 \
 //y=7.4 //x2=8.14 //y2=3.7
cc_726 ( N_VDD_c_562_n N_noxref_7_c_2239_n ) capacitor c=0.041662f //x=8.88 \
 //y=7.4 //x2=8.14 //y2=3.7
cc_727 ( N_VDD_c_573_p N_noxref_7_c_2193_n ) capacitor c=0.00100981f //x=38.48 \
 //y=7.4 //x2=11.84 //y2=2.085
cc_728 ( N_VDD_c_563_n N_noxref_7_c_2193_n ) capacitor c=0.0246707f //x=11.1 \
 //y=7.4 //x2=11.84 //y2=2.085
cc_729 ( N_VDD_c_564_n N_noxref_7_c_2193_n ) capacitor c=0.00156253f //x=13.32 \
 //y=7.4 //x2=11.84 //y2=2.085
cc_730 ( N_VDD_M33_noxref_s N_noxref_7_c_2193_n ) capacitor c=0.0063632f \
 //x=11.64 //y=5.02 //x2=11.84 //y2=2.085
cc_731 ( N_VDD_c_564_n N_noxref_7_c_2198_n ) capacitor c=0.0140445f //x=13.32 \
 //y=7.4 //x2=14.43 //y2=2.085
cc_732 ( N_VDD_c_567_n N_noxref_7_c_2199_n ) capacitor c=9.1919e-19 //x=22.2 \
 //y=7.4 //x2=24.05 //y2=2.08
cc_733 ( N_VDD_c_568_n N_noxref_7_c_2199_n ) capacitor c=9.05139e-19 //x=25.53 \
 //y=7.4 //x2=24.05 //y2=2.08
cc_734 ( N_VDD_c_661_p N_noxref_7_M33_noxref_g ) capacitor c=0.00748034f \
 //x=12.57 //y=7.4 //x2=11.995 //y2=6.02
cc_735 ( N_VDD_c_563_n N_noxref_7_M33_noxref_g ) capacitor c=0.00599876f \
 //x=11.1 //y=7.4 //x2=11.995 //y2=6.02
cc_736 ( N_VDD_M33_noxref_s N_noxref_7_M33_noxref_g ) capacitor c=0.0528676f \
 //x=11.64 //y=5.02 //x2=11.995 //y2=6.02
cc_737 ( N_VDD_c_661_p N_noxref_7_M34_noxref_g ) capacitor c=0.00697478f \
 //x=12.57 //y=7.4 //x2=12.435 //y2=6.02
cc_738 ( N_VDD_M34_noxref_d N_noxref_7_M34_noxref_g ) capacitor c=0.0528676f \
 //x=12.51 //y=5.02 //x2=12.435 //y2=6.02
cc_739 ( N_VDD_c_663_p N_noxref_7_M35_noxref_g ) capacitor c=0.00673447f \
 //x=14.465 //y=7.4 //x2=14.33 //y2=6.02
cc_740 ( N_VDD_c_564_n N_noxref_7_M35_noxref_g ) capacitor c=0.00449901f \
 //x=13.32 //y=7.4 //x2=14.33 //y2=6.02
cc_741 ( N_VDD_M35_noxref_d N_noxref_7_M35_noxref_g ) capacitor c=0.0166176f \
 //x=14.405 //y=5.02 //x2=14.33 //y2=6.02
cc_742 ( N_VDD_c_664_p N_noxref_7_M36_noxref_g ) capacitor c=0.006727f \
 //x=16.48 //y=7.4 //x2=14.77 //y2=6.02
cc_743 ( N_VDD_M35_noxref_d N_noxref_7_M36_noxref_g ) capacitor c=0.0186652f \
 //x=14.405 //y=5.02 //x2=14.77 //y2=6.02
cc_744 ( N_VDD_c_759_p N_noxref_7_M47_noxref_g ) capacitor c=0.00673971f \
 //x=24.665 //y=7.4 //x2=24.09 //y2=6.02
cc_745 ( N_VDD_M46_noxref_d N_noxref_7_M47_noxref_g ) capacitor c=0.015318f \
 //x=23.725 //y=5.02 //x2=24.09 //y2=6.02
cc_746 ( N_VDD_c_759_p N_noxref_7_M48_noxref_g ) capacitor c=0.00672952f \
 //x=24.665 //y=7.4 //x2=24.53 //y2=6.02
cc_747 ( N_VDD_c_568_n N_noxref_7_M48_noxref_g ) capacitor c=0.00883456f \
 //x=25.53 //y=7.4 //x2=24.53 //y2=6.02
cc_748 ( N_VDD_M48_noxref_d N_noxref_7_M48_noxref_g ) capacitor c=0.0430452f \
 //x=24.605 //y=5.02 //x2=24.53 //y2=6.02
cc_749 ( N_VDD_c_564_n N_noxref_7_c_2263_n ) capacitor c=0.0100096f //x=13.32 \
 //y=7.4 //x2=12.36 //y2=4.79
cc_750 ( N_VDD_c_563_n N_noxref_7_c_2264_n ) capacitor c=0.00683901f //x=11.1 \
 //y=7.4 //x2=12.07 //y2=4.79
cc_751 ( N_VDD_M33_noxref_s N_noxref_7_c_2264_n ) capacitor c=0.00495203f \
 //x=11.64 //y=5.02 //x2=12.07 //y2=4.79
cc_752 ( N_VDD_c_564_n N_noxref_7_c_2266_n ) capacitor c=0.0097362f //x=13.32 \
 //y=7.4 //x2=14.43 //y2=4.7
cc_753 ( N_VDD_c_561_n N_noxref_7_M25_noxref_d ) capacitor c=0.00966019f \
 //x=5.55 //y=7.4 //x2=4.185 //y2=5.02
cc_754 ( N_VDD_M23_noxref_d N_noxref_7_M25_noxref_d ) capacitor c=0.00561178f \
 //x=3.305 //y=5.02 //x2=4.185 //y2=5.02
cc_755 ( N_VDD_c_562_n N_noxref_7_M29_noxref_d ) capacitor c=0.00966019f \
 //x=8.88 //y=7.4 //x2=7.515 //y2=5.02
cc_756 ( N_VDD_M27_noxref_d N_noxref_7_M29_noxref_d ) capacitor c=0.00561178f \
 //x=6.635 //y=5.02 //x2=7.515 //y2=5.02
cc_757 ( N_VDD_M31_noxref_s N_noxref_7_M29_noxref_d ) capacitor c=5.00921e-19 \
 //x=9.42 //y=5.02 //x2=7.515 //y2=5.02
cc_758 ( N_VDD_c_661_p N_noxref_8_c_2617_n ) capacitor c=7.46634e-19 //x=12.57 \
 //y=7.4 //x2=12.495 //y2=4.58
cc_759 ( N_VDD_M34_noxref_d N_noxref_8_c_2617_n ) capacitor c=0.00520568f \
 //x=12.51 //y=5.02 //x2=12.495 //y2=4.58
cc_760 ( N_VDD_c_563_n N_noxref_8_c_2619_n ) capacitor c=0.0169935f //x=11.1 \
 //y=7.4 //x2=12.3 //y2=4.58
cc_761 ( N_VDD_c_563_n N_noxref_8_c_2607_n ) capacitor c=7.07219e-19 //x=11.1 \
 //y=7.4 //x2=12.58 //y2=2.59
cc_762 ( N_VDD_c_564_n N_noxref_8_c_2607_n ) capacitor c=0.021915f //x=13.32 \
 //y=7.4 //x2=12.58 //y2=2.59
cc_763 ( N_VDD_c_565_n N_noxref_8_c_2610_n ) capacitor c=0.00191336f //x=16.65 \
 //y=7.4 //x2=18.87 //y2=2.085
cc_764 ( N_VDD_c_566_n N_noxref_8_c_2610_n ) capacitor c=0.00116549f //x=19.98 \
 //y=7.4 //x2=18.87 //y2=2.085
cc_765 ( N_VDD_c_666_p N_noxref_8_M41_noxref_g ) capacitor c=0.00510247f \
 //x=19.81 //y=7.4 //x2=18.54 //y2=6.02
cc_766 ( N_VDD_c_666_p N_noxref_8_M42_noxref_g ) capacitor c=0.00510919f \
 //x=19.81 //y=7.4 //x2=18.98 //y2=6.02
cc_767 ( N_VDD_c_566_n N_noxref_8_M42_noxref_g ) capacitor c=0.00788519f \
 //x=19.98 //y=7.4 //x2=18.98 //y2=6.02
cc_768 ( N_VDD_c_573_p N_noxref_8_M33_noxref_d ) capacitor c=0.00264616f \
 //x=38.48 //y=7.4 //x2=12.07 //y2=5.02
cc_769 ( N_VDD_c_661_p N_noxref_8_M33_noxref_d ) capacitor c=0.0139918f \
 //x=12.57 //y=7.4 //x2=12.07 //y2=5.02
cc_770 ( N_VDD_c_564_n N_noxref_8_M33_noxref_d ) capacitor c=0.0183803f \
 //x=13.32 //y=7.4 //x2=12.07 //y2=5.02
cc_771 ( N_VDD_M33_noxref_s N_noxref_8_M33_noxref_d ) capacitor c=0.0843065f \
 //x=11.64 //y=5.02 //x2=12.07 //y2=5.02
cc_772 ( N_VDD_M34_noxref_d N_noxref_8_M33_noxref_d ) capacitor c=0.0832641f \
 //x=12.51 //y=5.02 //x2=12.07 //y2=5.02
cc_773 ( N_VDD_c_564_n SUM ) capacitor c=0.00142003f //x=13.32 //y=7.4 \
 //x2=15.91 //y2=3.33
cc_774 ( N_VDD_c_565_n SUM ) capacitor c=0.0423063f //x=16.65 //y=7.4 \
 //x2=15.91 //y2=3.33
cc_775 ( N_VDD_c_565_n SUM ) capacitor c=0.00157398f //x=16.65 //y=7.4 \
 //x2=19.24 //y2=2.59
cc_776 ( N_VDD_c_566_n SUM ) capacitor c=0.0398339f //x=19.98 //y=7.4 \
 //x2=19.24 //y2=2.59
cc_777 ( N_VDD_c_573_p N_SUM_c_2779_n ) capacitor c=0.00113298f //x=38.48 \
 //y=7.4 //x2=15.825 //y2=5.205
cc_778 ( N_VDD_c_664_p N_SUM_c_2779_n ) capacitor c=0.00138901f //x=16.48 \
 //y=7.4 //x2=15.825 //y2=5.205
cc_779 ( N_VDD_c_564_n N_SUM_c_2781_n ) capacitor c=8.9933e-19 //x=13.32 \
 //y=7.4 //x2=15.515 //y2=5.205
cc_780 ( N_VDD_c_573_p N_SUM_c_2782_n ) capacitor c=0.00113298f //x=38.48 \
 //y=7.4 //x2=19.155 //y2=5.205
cc_781 ( N_VDD_c_666_p N_SUM_c_2782_n ) capacitor c=0.00138901f //x=19.81 \
 //y=7.4 //x2=19.155 //y2=5.205
cc_782 ( N_VDD_c_565_n N_SUM_c_2784_n ) capacitor c=8.9933e-19 //x=16.65 \
 //y=7.4 //x2=18.845 //y2=5.205
cc_783 ( N_VDD_c_565_n N_SUM_M37_noxref_d ) capacitor c=0.00966019f //x=16.65 \
 //y=7.4 //x2=15.285 //y2=5.02
cc_784 ( N_VDD_M35_noxref_d N_SUM_M37_noxref_d ) capacitor c=0.00561178f \
 //x=14.405 //y=5.02 //x2=15.285 //y2=5.02
cc_785 ( N_VDD_c_566_n N_SUM_M41_noxref_d ) capacitor c=0.00966019f //x=19.98 \
 //y=7.4 //x2=18.615 //y2=5.02
cc_786 ( N_VDD_M39_noxref_d N_SUM_M41_noxref_d ) capacitor c=0.00561178f \
 //x=17.735 //y=5.02 //x2=18.615 //y2=5.02
cc_787 ( N_VDD_M43_noxref_s N_SUM_M41_noxref_d ) capacitor c=5.00921e-19 \
 //x=20.52 //y=5.02 //x2=18.615 //y2=5.02
cc_788 ( N_VDD_c_565_n N_noxref_10_c_2933_n ) capacitor c=0.0190041f //x=16.65 \
 //y=7.4 //x2=20.605 //y2=4.07
cc_789 ( N_VDD_c_566_n N_noxref_10_c_2933_n ) capacitor c=0.0150593f //x=19.98 \
 //y=7.4 //x2=20.605 //y2=4.07
cc_790 ( N_VDD_c_564_n N_noxref_10_c_2935_n ) capacitor c=5.31823e-19 \
 //x=13.32 //y=7.4 //x2=15.54 //y2=4.07
cc_791 ( N_VDD_c_565_n N_noxref_10_c_2935_n ) capacitor c=0.00180941f \
 //x=16.65 //y=7.4 //x2=15.54 //y2=4.07
cc_792 ( N_VDD_c_566_n N_noxref_10_c_2914_n ) capacitor c=0.0195394f //x=19.98 \
 //y=7.4 //x2=20.72 //y2=3.33
cc_793 ( N_VDD_c_567_n N_noxref_10_c_2914_n ) capacitor c=4.66518e-19 //x=22.2 \
 //y=7.4 //x2=20.72 //y2=3.33
cc_794 ( N_VDD_c_567_n N_noxref_10_c_2939_n ) capacitor c=0.0170839f //x=22.2 \
 //y=7.4 //x2=21 //y2=4.58
cc_795 ( N_VDD_c_668_p N_noxref_10_c_2940_n ) capacitor c=0.00100547f \
 //x=21.44 //y=7.4 //x2=20.805 //y2=4.58
cc_796 ( N_VDD_M43_noxref_s N_noxref_10_c_2940_n ) capacitor c=0.00542914f \
 //x=20.52 //y=5.02 //x2=20.805 //y2=4.58
cc_797 ( N_VDD_c_664_p N_noxref_10_M37_noxref_g ) capacitor c=0.00510247f \
 //x=16.48 //y=7.4 //x2=15.21 //y2=6.02
cc_798 ( N_VDD_c_664_p N_noxref_10_M38_noxref_g ) capacitor c=0.00510919f \
 //x=16.48 //y=7.4 //x2=15.65 //y2=6.02
cc_799 ( N_VDD_c_565_n N_noxref_10_M38_noxref_g ) capacitor c=0.01202f \
 //x=16.65 //y=7.4 //x2=15.65 //y2=6.02
cc_800 ( N_VDD_c_573_p N_noxref_10_M43_noxref_d ) capacitor c=0.00264616f \
 //x=38.48 //y=7.4 //x2=20.94 //y2=5.02
cc_801 ( N_VDD_c_668_p N_noxref_10_M43_noxref_d ) capacitor c=0.0139918f \
 //x=21.44 //y=7.4 //x2=20.94 //y2=5.02
cc_802 ( N_VDD_c_566_n N_noxref_10_M43_noxref_d ) capacitor c=0.0181582f \
 //x=19.98 //y=7.4 //x2=20.94 //y2=5.02
cc_803 ( N_VDD_M43_noxref_s N_noxref_10_M43_noxref_d ) capacitor c=0.0832641f \
 //x=20.52 //y=5.02 //x2=20.94 //y2=5.02
cc_804 ( N_VDD_M44_noxref_d N_noxref_10_M43_noxref_d ) capacitor c=0.0843065f \
 //x=21.38 //y=5.02 //x2=20.94 //y2=5.02
cc_805 ( N_VDD_c_566_n N_CIN_c_3115_n ) capacitor c=0.0250986f //x=19.98 \
 //y=7.4 //x2=21.345 //y2=4.44
cc_806 ( N_VDD_c_565_n N_CIN_c_3116_n ) capacitor c=0.00666294f //x=16.65 \
 //y=7.4 //x2=17.875 //y2=4.44
cc_807 ( N_VDD_c_567_n N_CIN_c_3087_n ) capacitor c=0.0301333f //x=22.2 \
 //y=7.4 //x2=23.195 //y2=4.44
cc_808 ( N_VDD_c_567_n N_CIN_c_3118_n ) capacitor c=0.00113468f //x=22.2 \
 //y=7.4 //x2=21.575 //y2=4.44
cc_809 ( N_VDD_c_565_n CIN ) capacitor c=0.00930479f //x=16.65 //y=7.4 \
 //x2=17.76 //y2=4.44
cc_810 ( N_VDD_c_573_p N_CIN_c_3090_n ) capacitor c=0.00100981f //x=38.48 \
 //y=7.4 //x2=21.46 //y2=2.085
cc_811 ( N_VDD_c_566_n N_CIN_c_3090_n ) capacitor c=7.316e-19 //x=19.98 \
 //y=7.4 //x2=21.46 //y2=2.085
cc_812 ( N_VDD_c_567_n N_CIN_c_3090_n ) capacitor c=0.0225516f //x=22.2 \
 //y=7.4 //x2=21.46 //y2=2.085
cc_813 ( N_VDD_M44_noxref_d N_CIN_c_3090_n ) capacitor c=0.0063632f //x=21.38 \
 //y=5.02 //x2=21.46 //y2=2.085
cc_814 ( N_VDD_c_573_p N_CIN_c_3095_n ) capacitor c=8.0695e-19 //x=38.48 \
 //y=7.4 //x2=23.31 //y2=2.08
cc_815 ( N_VDD_c_567_n N_CIN_c_3095_n ) capacitor c=0.0118247f //x=22.2 \
 //y=7.4 //x2=23.31 //y2=2.08
cc_816 ( N_VDD_c_665_p N_CIN_M39_noxref_g ) capacitor c=0.00673447f //x=17.795 \
 //y=7.4 //x2=17.66 //y2=6.02
cc_817 ( N_VDD_c_565_n N_CIN_M39_noxref_g ) capacitor c=0.00661226f //x=16.65 \
 //y=7.4 //x2=17.66 //y2=6.02
cc_818 ( N_VDD_M39_noxref_d N_CIN_M39_noxref_g ) capacitor c=0.0166176f \
 //x=17.735 //y=5.02 //x2=17.66 //y2=6.02
cc_819 ( N_VDD_c_666_p N_CIN_M40_noxref_g ) capacitor c=0.006727f //x=19.81 \
 //y=7.4 //x2=18.1 //y2=6.02
cc_820 ( N_VDD_M39_noxref_d N_CIN_M40_noxref_g ) capacitor c=0.0186652f \
 //x=17.735 //y=5.02 //x2=18.1 //y2=6.02
cc_821 ( N_VDD_c_668_p N_CIN_M43_noxref_g ) capacitor c=0.00697478f //x=21.44 \
 //y=7.4 //x2=20.865 //y2=6.02
cc_822 ( N_VDD_M43_noxref_s N_CIN_M43_noxref_g ) capacitor c=0.0528676f \
 //x=20.52 //y=5.02 //x2=20.865 //y2=6.02
cc_823 ( N_VDD_c_668_p N_CIN_M44_noxref_g ) capacitor c=0.00748034f //x=21.44 \
 //y=7.4 //x2=21.305 //y2=6.02
cc_824 ( N_VDD_c_567_n N_CIN_M44_noxref_g ) capacitor c=0.00617701f //x=22.2 \
 //y=7.4 //x2=21.305 //y2=6.02
cc_825 ( N_VDD_M44_noxref_d N_CIN_M44_noxref_g ) capacitor c=0.0528676f \
 //x=21.38 //y=5.02 //x2=21.305 //y2=6.02
cc_826 ( N_VDD_c_671_p N_CIN_M45_noxref_g ) capacitor c=0.00726866f //x=23.785 \
 //y=7.4 //x2=23.21 //y2=6.02
cc_827 ( N_VDD_M45_noxref_s N_CIN_M45_noxref_g ) capacitor c=0.054195f \
 //x=22.855 //y=5.02 //x2=23.21 //y2=6.02
cc_828 ( N_VDD_c_671_p N_CIN_M46_noxref_g ) capacitor c=0.00672952f //x=23.785 \
 //y=7.4 //x2=23.65 //y2=6.02
cc_829 ( N_VDD_M46_noxref_d N_CIN_M46_noxref_g ) capacitor c=0.015318f \
 //x=23.725 //y=5.02 //x2=23.65 //y2=6.02
cc_830 ( N_VDD_c_566_n N_CIN_c_3140_n ) capacitor c=0.0117981f //x=19.98 \
 //y=7.4 //x2=20.94 //y2=4.79
cc_831 ( N_VDD_c_567_n N_CIN_c_3141_n ) capacitor c=0.00843885f //x=22.2 \
 //y=7.4 //x2=21.305 //y2=4.865
cc_832 ( N_VDD_M44_noxref_d N_CIN_c_3141_n ) capacitor c=0.00495203f //x=21.38 \
 //y=5.02 //x2=21.305 //y2=4.865
cc_833 ( N_VDD_c_565_n N_CIN_c_3143_n ) capacitor c=0.00997846f //x=16.65 \
 //y=7.4 //x2=17.76 //y2=4.7
cc_834 ( N_VDD_c_567_n N_CIN_c_3144_n ) capacitor c=0.00965617f //x=22.2 \
 //y=7.4 //x2=23.31 //y2=4.7
cc_835 ( N_VDD_c_568_n N_noxref_12_c_3336_n ) capacitor c=0.0050908f //x=25.53 \
 //y=7.4 //x2=26.155 //y2=3.33
cc_836 ( N_VDD_c_573_p N_noxref_12_c_3359_n ) capacitor c=0.00446322f \
 //x=38.48 //y=7.4 //x2=24.225 //y2=5.2
cc_837 ( N_VDD_c_671_p N_noxref_12_c_3359_n ) capacitor c=4.48037e-19 \
 //x=23.785 //y=7.4 //x2=24.225 //y2=5.2
cc_838 ( N_VDD_c_759_p N_noxref_12_c_3359_n ) capacitor c=4.48037e-19 \
 //x=24.665 //y=7.4 //x2=24.225 //y2=5.2
cc_839 ( N_VDD_M46_noxref_d N_noxref_12_c_3359_n ) capacitor c=0.0121037f \
 //x=23.725 //y=5.02 //x2=24.225 //y2=5.2
cc_840 ( N_VDD_c_567_n N_noxref_12_c_3363_n ) capacitor c=0.00985474f //x=22.2 \
 //y=7.4 //x2=23.515 //y2=5.2
cc_841 ( N_VDD_M45_noxref_s N_noxref_12_c_3363_n ) capacitor c=0.087833f \
 //x=22.855 //y=5.02 //x2=23.515 //y2=5.2
cc_842 ( N_VDD_c_573_p N_noxref_12_c_3365_n ) capacitor c=0.00294854f \
 //x=38.48 //y=7.4 //x2=24.705 //y2=5.2
cc_843 ( N_VDD_c_759_p N_noxref_12_c_3365_n ) capacitor c=7.70829e-19 \
 //x=24.665 //y=7.4 //x2=24.705 //y2=5.2
cc_844 ( N_VDD_M48_noxref_d N_noxref_12_c_3365_n ) capacitor c=0.0154095f \
 //x=24.605 //y=5.02 //x2=24.705 //y2=5.2
cc_845 ( N_VDD_c_567_n N_noxref_12_c_3368_n ) capacitor c=0.00138008f //x=22.2 \
 //y=7.4 //x2=24.79 //y2=3.33
cc_846 ( N_VDD_c_568_n N_noxref_12_c_3368_n ) capacitor c=0.043426f //x=25.53 \
 //y=7.4 //x2=24.79 //y2=3.33
cc_847 ( N_VDD_c_573_p N_noxref_12_c_3339_n ) capacitor c=0.00100981f \
 //x=38.48 //y=7.4 //x2=26.27 //y2=2.085
cc_848 ( N_VDD_c_568_n N_noxref_12_c_3339_n ) capacitor c=0.0249238f //x=25.53 \
 //y=7.4 //x2=26.27 //y2=2.085
cc_849 ( N_VDD_c_569_n N_noxref_12_c_3339_n ) capacitor c=0.00131929f \
 //x=27.75 //y=7.4 //x2=26.27 //y2=2.085
cc_850 ( N_VDD_M49_noxref_s N_noxref_12_c_3339_n ) capacitor c=0.00653582f \
 //x=26.07 //y=5.02 //x2=26.27 //y2=2.085
cc_851 ( N_VDD_c_674_p N_noxref_12_M49_noxref_g ) capacitor c=0.00748034f \
 //x=27 //y=7.4 //x2=26.425 //y2=6.02
cc_852 ( N_VDD_c_568_n N_noxref_12_M49_noxref_g ) capacitor c=0.00860016f \
 //x=25.53 //y=7.4 //x2=26.425 //y2=6.02
cc_853 ( N_VDD_M49_noxref_s N_noxref_12_M49_noxref_g ) capacitor c=0.0528676f \
 //x=26.07 //y=5.02 //x2=26.425 //y2=6.02
cc_854 ( N_VDD_c_674_p N_noxref_12_M50_noxref_g ) capacitor c=0.00697478f \
 //x=27 //y=7.4 //x2=26.865 //y2=6.02
cc_855 ( N_VDD_M50_noxref_d N_noxref_12_M50_noxref_g ) capacitor c=0.0528676f \
 //x=26.94 //y=5.02 //x2=26.865 //y2=6.02
cc_856 ( N_VDD_c_569_n N_noxref_12_c_3379_n ) capacitor c=0.00792909f \
 //x=27.75 //y=7.4 //x2=26.79 //y2=4.79
cc_857 ( N_VDD_c_568_n N_noxref_12_c_3380_n ) capacitor c=0.00684036f \
 //x=25.53 //y=7.4 //x2=26.5 //y2=4.79
cc_858 ( N_VDD_M49_noxref_s N_noxref_12_c_3380_n ) capacitor c=0.00495203f \
 //x=26.07 //y=5.02 //x2=26.5 //y2=4.79
cc_859 ( N_VDD_c_573_p N_noxref_12_M45_noxref_d ) capacitor c=0.00264475f \
 //x=38.48 //y=7.4 //x2=23.285 //y2=5.02
cc_860 ( N_VDD_c_671_p N_noxref_12_M45_noxref_d ) capacitor c=0.0139566f \
 //x=23.785 //y=7.4 //x2=23.285 //y2=5.02
cc_861 ( N_VDD_c_568_n N_noxref_12_M45_noxref_d ) capacitor c=6.94454e-19 \
 //x=25.53 //y=7.4 //x2=23.285 //y2=5.02
cc_862 ( N_VDD_M46_noxref_d N_noxref_12_M45_noxref_d ) capacitor c=0.0664752f \
 //x=23.725 //y=5.02 //x2=23.285 //y2=5.02
cc_863 ( N_VDD_c_573_p N_noxref_12_M47_noxref_d ) capacitor c=0.00264475f \
 //x=38.48 //y=7.4 //x2=24.165 //y2=5.02
cc_864 ( N_VDD_c_759_p N_noxref_12_M47_noxref_d ) capacitor c=0.0139566f \
 //x=24.665 //y=7.4 //x2=24.165 //y2=5.02
cc_865 ( N_VDD_c_568_n N_noxref_12_M47_noxref_d ) capacitor c=0.0120541f \
 //x=25.53 //y=7.4 //x2=24.165 //y2=5.02
cc_866 ( N_VDD_M45_noxref_s N_noxref_12_M47_noxref_d ) capacitor c=0.00111971f \
 //x=22.855 //y=5.02 //x2=24.165 //y2=5.02
cc_867 ( N_VDD_M46_noxref_d N_noxref_12_M47_noxref_d ) capacitor c=0.0664752f \
 //x=23.725 //y=5.02 //x2=24.165 //y2=5.02
cc_868 ( N_VDD_M48_noxref_d N_noxref_12_M47_noxref_d ) capacitor c=0.0664752f \
 //x=24.605 //y=5.02 //x2=24.165 //y2=5.02
cc_869 ( N_VDD_M49_noxref_s N_noxref_12_M47_noxref_d ) capacitor c=5.1407e-19 \
 //x=26.07 //y=5.02 //x2=24.165 //y2=5.02
cc_870 ( N_VDD_c_573_p N_noxref_13_c_3497_n ) capacitor c=0.00920591f \
 //x=38.48 //y=7.4 //x2=31.705 //y2=3.33
cc_871 ( N_VDD_c_570_n N_noxref_13_c_3497_n ) capacitor c=0.0069465f //x=31.08 \
 //y=7.4 //x2=31.705 //y2=3.33
cc_872 ( N_VDD_M55_noxref_s N_noxref_13_c_3497_n ) capacitor c=0.00113028f \
 //x=31.62 //y=5.02 //x2=31.705 //y2=3.33
cc_873 ( N_VDD_c_573_p N_noxref_13_c_3500_n ) capacitor c=0.00161874f \
 //x=38.48 //y=7.4 //x2=30.455 //y2=3.33
cc_874 ( N_VDD_M54_noxref_d N_noxref_13_c_3500_n ) capacitor c=3.3085e-19 \
 //x=30.155 //y=5.02 //x2=30.455 //y2=3.33
cc_875 ( N_VDD_c_573_p N_noxref_13_c_3502_n ) capacitor c=0.0047626f //x=38.48 \
 //y=7.4 //x2=29.775 //y2=5.2
cc_876 ( N_VDD_c_677_p N_noxref_13_c_3502_n ) capacitor c=4.3394e-19 \
 //x=29.335 //y=7.4 //x2=29.775 //y2=5.2
cc_877 ( N_VDD_c_601_p N_noxref_13_c_3502_n ) capacitor c=4.3394e-19 \
 //x=30.215 //y=7.4 //x2=29.775 //y2=5.2
cc_878 ( N_VDD_M52_noxref_d N_noxref_13_c_3502_n ) capacitor c=0.012665f \
 //x=29.275 //y=5.02 //x2=29.775 //y2=5.2
cc_879 ( N_VDD_c_569_n N_noxref_13_c_3506_n ) capacitor c=0.00985474f \
 //x=27.75 //y=7.4 //x2=29.065 //y2=5.2
cc_880 ( N_VDD_M51_noxref_s N_noxref_13_c_3506_n ) capacitor c=0.087833f \
 //x=28.405 //y=5.02 //x2=29.065 //y2=5.2
cc_881 ( N_VDD_c_573_p N_noxref_13_c_3508_n ) capacitor c=0.00318278f \
 //x=38.48 //y=7.4 //x2=30.255 //y2=5.2
cc_882 ( N_VDD_c_601_p N_noxref_13_c_3508_n ) capacitor c=7.21492e-19 \
 //x=30.215 //y=7.4 //x2=30.255 //y2=5.2
cc_883 ( N_VDD_M54_noxref_d N_noxref_13_c_3508_n ) capacitor c=0.016468f \
 //x=30.155 //y=5.02 //x2=30.255 //y2=5.2
cc_884 ( N_VDD_c_569_n N_noxref_13_c_3477_n ) capacitor c=0.00137938f \
 //x=27.75 //y=7.4 //x2=30.34 //y2=3.33
cc_885 ( N_VDD_c_570_n N_noxref_13_c_3477_n ) capacitor c=0.0455991f //x=31.08 \
 //y=7.4 //x2=30.34 //y2=3.33
cc_886 ( N_VDD_c_573_p N_noxref_13_c_3478_n ) capacitor c=0.00160122f \
 //x=38.48 //y=7.4 //x2=31.82 //y2=2.085
cc_887 ( N_VDD_c_570_n N_noxref_13_c_3478_n ) capacitor c=0.0272613f //x=31.08 \
 //y=7.4 //x2=31.82 //y2=2.085
cc_888 ( N_VDD_c_571_n N_noxref_13_c_3478_n ) capacitor c=0.00144308f //x=33.3 \
 //y=7.4 //x2=31.82 //y2=2.085
cc_889 ( N_VDD_M55_noxref_s N_noxref_13_c_3478_n ) capacitor c=0.00951228f \
 //x=31.62 //y=5.02 //x2=31.82 //y2=2.085
cc_890 ( N_VDD_c_905_p N_noxref_13_M55_noxref_g ) capacitor c=0.00748034f \
 //x=32.55 //y=7.4 //x2=31.975 //y2=6.02
cc_891 ( N_VDD_c_570_n N_noxref_13_M55_noxref_g ) capacitor c=0.00877732f \
 //x=31.08 //y=7.4 //x2=31.975 //y2=6.02
cc_892 ( N_VDD_M55_noxref_s N_noxref_13_M55_noxref_g ) capacitor c=0.0528676f \
 //x=31.62 //y=5.02 //x2=31.975 //y2=6.02
cc_893 ( N_VDD_c_905_p N_noxref_13_M56_noxref_g ) capacitor c=0.00697478f \
 //x=32.55 //y=7.4 //x2=32.415 //y2=6.02
cc_894 ( N_VDD_M56_noxref_d N_noxref_13_M56_noxref_g ) capacitor c=0.0528676f \
 //x=32.49 //y=5.02 //x2=32.415 //y2=6.02
cc_895 ( N_VDD_c_571_n N_noxref_13_c_3522_n ) capacitor c=0.012136f //x=33.3 \
 //y=7.4 //x2=32.34 //y2=4.79
cc_896 ( N_VDD_c_570_n N_noxref_13_c_3523_n ) capacitor c=0.00800869f \
 //x=31.08 //y=7.4 //x2=32.05 //y2=4.79
cc_897 ( N_VDD_M55_noxref_s N_noxref_13_c_3523_n ) capacitor c=0.00527247f \
 //x=31.62 //y=5.02 //x2=32.05 //y2=4.79
cc_898 ( N_VDD_c_573_p N_noxref_13_M51_noxref_d ) capacitor c=0.0043371f \
 //x=38.48 //y=7.4 //x2=28.835 //y2=5.02
cc_899 ( N_VDD_c_677_p N_noxref_13_M51_noxref_d ) capacitor c=0.013611f \
 //x=29.335 //y=7.4 //x2=28.835 //y2=5.02
cc_900 ( N_VDD_c_570_n N_noxref_13_M51_noxref_d ) capacitor c=6.94454e-19 \
 //x=31.08 //y=7.4 //x2=28.835 //y2=5.02
cc_901 ( N_VDD_M52_noxref_d N_noxref_13_M51_noxref_d ) capacitor c=0.0664752f \
 //x=29.275 //y=5.02 //x2=28.835 //y2=5.02
cc_902 ( N_VDD_c_573_p N_noxref_13_M53_noxref_d ) capacitor c=0.00582647f \
 //x=38.48 //y=7.4 //x2=29.715 //y2=5.02
cc_903 ( N_VDD_c_601_p N_noxref_13_M53_noxref_d ) capacitor c=0.0138379f \
 //x=30.215 //y=7.4 //x2=29.715 //y2=5.02
cc_904 ( N_VDD_c_570_n N_noxref_13_M53_noxref_d ) capacitor c=0.0120541f \
 //x=31.08 //y=7.4 //x2=29.715 //y2=5.02
cc_905 ( N_VDD_M51_noxref_s N_noxref_13_M53_noxref_d ) capacitor c=0.00111971f \
 //x=28.405 //y=5.02 //x2=29.715 //y2=5.02
cc_906 ( N_VDD_M52_noxref_d N_noxref_13_M53_noxref_d ) capacitor c=0.0664752f \
 //x=29.275 //y=5.02 //x2=29.715 //y2=5.02
cc_907 ( N_VDD_M54_noxref_d N_noxref_13_M53_noxref_d ) capacitor c=0.0664752f \
 //x=30.155 //y=5.02 //x2=29.715 //y2=5.02
cc_908 ( N_VDD_M55_noxref_s N_noxref_13_M53_noxref_d ) capacitor c=5.1407e-19 \
 //x=31.62 //y=5.02 //x2=29.715 //y2=5.02
cc_909 ( N_VDD_c_573_p N_noxref_14_c_3617_n ) capacitor c=0.0198728f //x=38.48 \
 //y=7.4 //x2=34.295 //y2=2.96
cc_910 ( N_VDD_c_569_n N_noxref_14_c_3617_n ) capacitor c=0.00344974f \
 //x=27.75 //y=7.4 //x2=34.295 //y2=2.96
cc_911 ( N_VDD_c_674_p N_noxref_14_c_3650_n ) capacitor c=7.46431e-19 //x=27 \
 //y=7.4 //x2=26.925 //y2=4.58
cc_912 ( N_VDD_M50_noxref_d N_noxref_14_c_3650_n ) capacitor c=0.00520568f \
 //x=26.94 //y=5.02 //x2=26.925 //y2=4.58
cc_913 ( N_VDD_c_568_n N_noxref_14_c_3652_n ) capacitor c=0.0170723f //x=25.53 \
 //y=7.4 //x2=26.73 //y2=4.58
cc_914 ( N_VDD_c_568_n N_noxref_14_c_3631_n ) capacitor c=4.80934e-19 \
 //x=25.53 //y=7.4 //x2=27.01 //y2=2.96
cc_915 ( N_VDD_c_569_n N_noxref_14_c_3631_n ) capacitor c=0.0226238f //x=27.75 \
 //y=7.4 //x2=27.01 //y2=2.96
cc_916 ( N_VDD_c_571_n N_noxref_14_c_3632_n ) capacitor c=0.0103855f //x=33.3 \
 //y=7.4 //x2=34.41 //y2=2.08
cc_917 ( N_VDD_c_573_p N_noxref_14_c_3656_n ) capacitor c=2.84083e-19 \
 //x=38.48 //y=7.4 //x2=34.255 //y2=4.705
cc_918 ( N_VDD_c_571_n N_noxref_14_c_3656_n ) capacitor c=0.00860173f //x=33.3 \
 //y=7.4 //x2=34.255 //y2=4.705
cc_919 ( N_VDD_M57_noxref_d N_noxref_14_c_3656_n ) capacitor c=3.49575e-19 \
 //x=34.385 //y=5.025 //x2=34.255 //y2=4.705
cc_920 ( N_VDD_c_935_p N_noxref_14_M57_noxref_g ) capacitor c=0.0067918f \
 //x=34.445 //y=7.4 //x2=34.31 //y2=6.025
cc_921 ( N_VDD_c_571_n N_noxref_14_M57_noxref_g ) capacitor c=0.00730892f \
 //x=33.3 //y=7.4 //x2=34.31 //y2=6.025
cc_922 ( N_VDD_M57_noxref_d N_noxref_14_M57_noxref_g ) capacitor c=0.0156786f \
 //x=34.385 //y=5.025 //x2=34.31 //y2=6.025
cc_923 ( N_VDD_c_938_p N_noxref_14_M58_noxref_g ) capacitor c=0.00678153f \
 //x=36.46 //y=7.4 //x2=34.75 //y2=6.025
cc_924 ( N_VDD_M57_noxref_d N_noxref_14_M58_noxref_g ) capacitor c=0.0183011f \
 //x=34.385 //y=5.025 //x2=34.75 //y2=6.025
cc_925 ( N_VDD_c_571_n N_noxref_14_c_3664_n ) capacitor c=0.00890932f //x=33.3 \
 //y=7.4 //x2=34.255 //y2=4.705
cc_926 ( N_VDD_c_573_p N_noxref_14_M49_noxref_d ) capacitor c=0.00264616f \
 //x=38.48 //y=7.4 //x2=26.5 //y2=5.02
cc_927 ( N_VDD_c_674_p N_noxref_14_M49_noxref_d ) capacitor c=0.0139918f \
 //x=27 //y=7.4 //x2=26.5 //y2=5.02
cc_928 ( N_VDD_c_569_n N_noxref_14_M49_noxref_d ) capacitor c=0.0183306f \
 //x=27.75 //y=7.4 //x2=26.5 //y2=5.02
cc_929 ( N_VDD_M49_noxref_s N_noxref_14_M49_noxref_d ) capacitor c=0.0843065f \
 //x=26.07 //y=5.02 //x2=26.5 //y2=5.02
cc_930 ( N_VDD_M50_noxref_d N_noxref_14_M49_noxref_d ) capacitor c=0.0832641f \
 //x=26.94 //y=5.02 //x2=26.5 //y2=5.02
cc_931 ( N_VDD_c_573_p N_noxref_15_c_3782_n ) capacitor c=0.0153421f //x=38.48 \
 //y=7.4 //x2=35.035 //y2=3.33
cc_932 ( N_VDD_c_571_n N_noxref_15_c_3782_n ) capacitor c=0.0069465f //x=33.3 \
 //y=7.4 //x2=35.035 //y2=3.33
cc_933 ( N_VDD_M56_noxref_d N_noxref_15_c_3782_n ) capacitor c=5.17699e-19 \
 //x=32.49 //y=5.02 //x2=35.035 //y2=3.33
cc_934 ( N_VDD_c_573_p N_noxref_15_c_3803_n ) capacitor c=0.00163324f \
 //x=38.48 //y=7.4 //x2=32.675 //y2=3.33
cc_935 ( N_VDD_M56_noxref_d N_noxref_15_c_3803_n ) capacitor c=7.33386e-19 \
 //x=32.49 //y=5.02 //x2=32.675 //y2=3.33
cc_936 ( N_VDD_c_573_p N_noxref_15_c_3805_n ) capacitor c=0.00128923f \
 //x=38.48 //y=7.4 //x2=32.475 //y2=4.58
cc_937 ( N_VDD_c_905_p N_noxref_15_c_3805_n ) capacitor c=8.8179e-19 //x=32.55 \
 //y=7.4 //x2=32.475 //y2=4.58
cc_938 ( N_VDD_M56_noxref_d N_noxref_15_c_3805_n ) capacitor c=0.00627485f \
 //x=32.49 //y=5.02 //x2=32.475 //y2=4.58
cc_939 ( N_VDD_c_570_n N_noxref_15_c_3808_n ) capacitor c=0.0176572f //x=31.08 \
 //y=7.4 //x2=32.28 //y2=4.58
cc_940 ( N_VDD_c_570_n N_noxref_15_c_3786_n ) capacitor c=4.80934e-19 \
 //x=31.08 //y=7.4 //x2=32.56 //y2=3.33
cc_941 ( N_VDD_c_571_n N_noxref_15_c_3786_n ) capacitor c=0.02304f //x=33.3 \
 //y=7.4 //x2=32.56 //y2=3.33
cc_942 ( N_VDD_c_571_n N_noxref_15_c_3787_n ) capacitor c=7.02327e-19 //x=33.3 \
 //y=7.4 //x2=35.15 //y2=2.08
cc_943 ( N_VDD_c_572_n N_noxref_15_c_3787_n ) capacitor c=6.16704e-19 \
 //x=36.63 //y=7.4 //x2=35.15 //y2=2.08
cc_944 ( N_VDD_c_938_p N_noxref_15_M59_noxref_g ) capacitor c=0.00513565f \
 //x=36.46 //y=7.4 //x2=35.19 //y2=6.025
cc_945 ( N_VDD_c_938_p N_noxref_15_M60_noxref_g ) capacitor c=0.00512552f \
 //x=36.46 //y=7.4 //x2=35.63 //y2=6.025
cc_946 ( N_VDD_c_572_n N_noxref_15_M60_noxref_g ) capacitor c=0.0120232f \
 //x=36.63 //y=7.4 //x2=35.63 //y2=6.025
cc_947 ( N_VDD_c_573_p N_noxref_15_M55_noxref_d ) capacitor c=0.00585331f \
 //x=38.48 //y=7.4 //x2=32.05 //y2=5.02
cc_948 ( N_VDD_c_905_p N_noxref_15_M55_noxref_d ) capacitor c=0.0139004f \
 //x=32.55 //y=7.4 //x2=32.05 //y2=5.02
cc_949 ( N_VDD_c_571_n N_noxref_15_M55_noxref_d ) capacitor c=0.0204646f \
 //x=33.3 //y=7.4 //x2=32.05 //y2=5.02
cc_950 ( N_VDD_M55_noxref_s N_noxref_15_M55_noxref_d ) capacitor c=0.0843065f \
 //x=31.62 //y=5.02 //x2=32.05 //y2=5.02
cc_951 ( N_VDD_M56_noxref_d N_noxref_15_M55_noxref_d ) capacitor c=0.0832641f \
 //x=32.49 //y=5.02 //x2=32.05 //y2=5.02
cc_952 ( N_VDD_c_573_p N_noxref_16_c_3919_n ) capacitor c=0.00920603f \
 //x=38.48 //y=7.4 //x2=37.255 //y2=3.33
cc_953 ( N_VDD_c_572_n N_noxref_16_c_3919_n ) capacitor c=0.0069465f //x=36.63 \
 //y=7.4 //x2=37.255 //y2=3.33
cc_954 ( N_VDD_M61_noxref_s N_noxref_16_c_3919_n ) capacitor c=0.00106085f \
 //x=37.17 //y=5.02 //x2=37.255 //y2=3.33
cc_955 ( N_VDD_c_573_p N_noxref_16_c_3925_n ) capacitor c=0.0014539f //x=38.48 \
 //y=7.4 //x2=36.005 //y2=3.33
cc_956 ( N_VDD_c_573_p N_noxref_16_c_3964_n ) capacitor c=0.00178185f \
 //x=38.48 //y=7.4 //x2=35.805 //y2=5.21
cc_957 ( N_VDD_c_938_p N_noxref_16_c_3964_n ) capacitor c=0.00136949f \
 //x=36.46 //y=7.4 //x2=35.805 //y2=5.21
cc_958 ( N_VDD_c_571_n N_noxref_16_c_3966_n ) capacitor c=8.9933e-19 //x=33.3 \
 //y=7.4 //x2=35.495 //y2=5.21
cc_959 ( N_VDD_c_571_n N_noxref_16_c_3936_n ) capacitor c=0.00163766f //x=33.3 \
 //y=7.4 //x2=35.89 //y2=3.33
cc_960 ( N_VDD_c_572_n N_noxref_16_c_3936_n ) capacitor c=0.0462234f //x=36.63 \
 //y=7.4 //x2=35.89 //y2=3.33
cc_961 ( N_VDD_c_573_p N_noxref_16_c_3937_n ) capacitor c=0.00160122f \
 //x=38.48 //y=7.4 //x2=37.37 //y2=2.085
cc_962 ( N_VDD_c_558_n N_noxref_16_c_3937_n ) capacitor c=0.00144809f \
 //x=38.48 //y=7.4 //x2=37.37 //y2=2.085
cc_963 ( N_VDD_c_572_n N_noxref_16_c_3937_n ) capacitor c=0.0272885f //x=36.63 \
 //y=7.4 //x2=37.37 //y2=2.085
cc_964 ( N_VDD_M61_noxref_s N_noxref_16_c_3937_n ) capacitor c=0.00971593f \
 //x=37.17 //y=5.02 //x2=37.37 //y2=2.085
cc_965 ( N_VDD_c_980_p N_noxref_16_M61_noxref_g ) capacitor c=0.00748034f \
 //x=38.1 //y=7.4 //x2=37.525 //y2=6.02
cc_966 ( N_VDD_c_572_n N_noxref_16_M61_noxref_g ) capacitor c=0.0102569f \
 //x=36.63 //y=7.4 //x2=37.525 //y2=6.02
cc_967 ( N_VDD_M61_noxref_s N_noxref_16_M61_noxref_g ) capacitor c=0.0528676f \
 //x=37.17 //y=5.02 //x2=37.525 //y2=6.02
cc_968 ( N_VDD_c_980_p N_noxref_16_M62_noxref_g ) capacitor c=0.00697478f \
 //x=38.1 //y=7.4 //x2=37.965 //y2=6.02
cc_969 ( N_VDD_M62_noxref_d N_noxref_16_M62_noxref_g ) capacitor c=0.0528676f \
 //x=38.04 //y=5.02 //x2=37.965 //y2=6.02
cc_970 ( N_VDD_c_558_n N_noxref_16_c_3978_n ) capacitor c=0.0287802f //x=38.48 \
 //y=7.4 //x2=37.89 //y2=4.79
cc_971 ( N_VDD_c_572_n N_noxref_16_c_3979_n ) capacitor c=0.011132f //x=36.63 \
 //y=7.4 //x2=37.6 //y2=4.79
cc_972 ( N_VDD_M61_noxref_s N_noxref_16_c_3979_n ) capacitor c=0.00527247f \
 //x=37.17 //y=5.02 //x2=37.6 //y2=4.79
cc_973 ( N_VDD_c_572_n N_noxref_16_M59_noxref_d ) capacitor c=0.00966019f \
 //x=36.63 //y=7.4 //x2=35.265 //y2=5.025
cc_974 ( N_VDD_M57_noxref_d N_noxref_16_M59_noxref_d ) capacitor c=0.00561178f \
 //x=34.385 //y=5.025 //x2=35.265 //y2=5.025
cc_975 ( N_VDD_M61_noxref_s N_noxref_16_M59_noxref_d ) capacitor c=4.94992e-19 \
 //x=37.17 //y=5.02 //x2=35.265 //y2=5.025
cc_976 ( N_VDD_c_573_p N_noxref_17_c_4059_n ) capacitor c=0.00494742f \
 //x=38.48 //y=7.4 //x2=3.805 //y2=5.205
cc_977 ( N_VDD_c_576_p N_noxref_17_c_4059_n ) capacitor c=4.50595e-19 \
 //x=3.365 //y=7.4 //x2=3.805 //y2=5.205
cc_978 ( N_VDD_c_599_p N_noxref_17_c_4059_n ) capacitor c=4.35755e-19 //x=5.38 \
 //y=7.4 //x2=3.805 //y2=5.205
cc_979 ( N_VDD_c_561_n N_noxref_17_c_4059_n ) capacitor c=0.00289291f //x=5.55 \
 //y=7.4 //x2=3.805 //y2=5.205
cc_980 ( N_VDD_M23_noxref_d N_noxref_17_c_4059_n ) capacitor c=0.0124635f \
 //x=3.305 //y=5.02 //x2=3.805 //y2=5.205
cc_981 ( N_VDD_c_560_n N_noxref_17_c_4064_n ) capacitor c=0.0628444f //x=2.22 \
 //y=7.4 //x2=3.095 //y2=5.205
cc_982 ( N_VDD_M22_noxref_d N_noxref_17_c_4064_n ) capacitor c=0.00269577f \
 //x=1.41 //y=5.02 //x2=3.095 //y2=5.205
cc_983 ( N_VDD_c_558_n N_noxref_17_c_4066_n ) capacitor c=0.0023707f //x=38.48 \
 //y=7.4 //x2=4.685 //y2=6.905
cc_984 ( N_VDD_c_573_p N_noxref_17_c_4067_n ) capacitor c=0.0260915f //x=38.48 \
 //y=7.4 //x2=3.975 //y2=6.905
cc_985 ( N_VDD_c_599_p N_noxref_17_c_4067_n ) capacitor c=0.0593394f //x=5.38 \
 //y=7.4 //x2=3.975 //y2=6.905
cc_986 ( N_VDD_c_573_p N_noxref_17_M23_noxref_s ) capacitor c=0.00242367f \
 //x=38.48 //y=7.4 //x2=2.875 //y2=5.02
cc_987 ( N_VDD_c_576_p N_noxref_17_M23_noxref_s ) capacitor c=0.0100244f \
 //x=3.365 //y=7.4 //x2=2.875 //y2=5.02
cc_988 ( N_VDD_M23_noxref_d N_noxref_17_M23_noxref_s ) capacitor c=0.061257f \
 //x=3.305 //y=5.02 //x2=2.875 //y2=5.02
cc_989 ( N_VDD_c_560_n N_noxref_17_M24_noxref_d ) capacitor c=0.00130916f \
 //x=2.22 //y=7.4 //x2=3.745 //y2=5.02
cc_990 ( N_VDD_M23_noxref_d N_noxref_17_M24_noxref_d ) capacitor c=0.0659925f \
 //x=3.305 //y=5.02 //x2=3.745 //y2=5.02
cc_991 ( N_VDD_c_561_n N_noxref_17_M26_noxref_d ) capacitor c=0.0520312f \
 //x=5.55 //y=7.4 //x2=4.625 //y2=5.02
cc_992 ( N_VDD_M23_noxref_d N_noxref_17_M26_noxref_d ) capacitor c=0.00107819f \
 //x=3.305 //y=5.02 //x2=4.625 //y2=5.02
cc_993 ( N_VDD_c_573_p N_noxref_19_c_4149_n ) capacitor c=0.00445614f \
 //x=38.48 //y=7.4 //x2=7.135 //y2=5.205
cc_994 ( N_VDD_c_629_p N_noxref_19_c_4149_n ) capacitor c=4.50436e-19 \
 //x=6.695 //y=7.4 //x2=7.135 //y2=5.205
cc_995 ( N_VDD_c_619_p N_noxref_19_c_4149_n ) capacitor c=4.50291e-19 //x=8.71 \
 //y=7.4 //x2=7.135 //y2=5.205
cc_996 ( N_VDD_c_562_n N_noxref_19_c_4149_n ) capacitor c=0.00289291f //x=8.88 \
 //y=7.4 //x2=7.135 //y2=5.205
cc_997 ( N_VDD_M27_noxref_d N_noxref_19_c_4149_n ) capacitor c=0.0123249f \
 //x=6.635 //y=5.02 //x2=7.135 //y2=5.205
cc_998 ( N_VDD_c_561_n N_noxref_19_c_4154_n ) capacitor c=0.0628444f //x=5.55 \
 //y=7.4 //x2=6.425 //y2=5.205
cc_999 ( N_VDD_c_558_n N_noxref_19_c_4155_n ) capacitor c=0.0023707f //x=38.48 \
 //y=7.4 //x2=8.015 //y2=6.905
cc_1000 ( N_VDD_c_573_p N_noxref_19_c_4156_n ) capacitor c=0.0164961f \
 //x=38.48 //y=7.4 //x2=7.305 //y2=6.905
cc_1001 ( N_VDD_c_619_p N_noxref_19_c_4156_n ) capacitor c=0.0608014f //x=8.71 \
 //y=7.4 //x2=7.305 //y2=6.905
cc_1002 ( N_VDD_c_573_p N_noxref_19_M27_noxref_s ) capacitor c=0.00242367f \
 //x=38.48 //y=7.4 //x2=6.205 //y2=5.02
cc_1003 ( N_VDD_c_629_p N_noxref_19_M27_noxref_s ) capacitor c=0.0100244f \
 //x=6.695 //y=7.4 //x2=6.205 //y2=5.02
cc_1004 ( N_VDD_M27_noxref_d N_noxref_19_M27_noxref_s ) capacitor c=0.061257f \
 //x=6.635 //y=5.02 //x2=6.205 //y2=5.02
cc_1005 ( N_VDD_c_561_n N_noxref_19_M28_noxref_d ) capacitor c=0.00130916f \
 //x=5.55 //y=7.4 //x2=7.075 //y2=5.02
cc_1006 ( N_VDD_M27_noxref_d N_noxref_19_M28_noxref_d ) capacitor c=0.0659925f \
 //x=6.635 //y=5.02 //x2=7.075 //y2=5.02
cc_1007 ( N_VDD_c_562_n N_noxref_19_M30_noxref_d ) capacitor c=0.0520312f \
 //x=8.88 //y=7.4 //x2=7.955 //y2=5.02
cc_1008 ( N_VDD_M27_noxref_d N_noxref_19_M30_noxref_d ) capacitor \
 c=0.00107819f //x=6.635 //y=5.02 //x2=7.955 //y2=5.02
cc_1009 ( N_VDD_M31_noxref_s N_noxref_19_M30_noxref_d ) capacitor \
 c=0.00230193f //x=9.42 //y=5.02 //x2=7.955 //y2=5.02
cc_1010 ( N_VDD_c_573_p N_noxref_21_c_4240_n ) capacitor c=0.00437344f \
 //x=38.48 //y=7.4 //x2=14.905 //y2=5.205
cc_1011 ( N_VDD_c_663_p N_noxref_21_c_4240_n ) capacitor c=4.49935e-19 \
 //x=14.465 //y=7.4 //x2=14.905 //y2=5.205
cc_1012 ( N_VDD_c_664_p N_noxref_21_c_4240_n ) capacitor c=4.49935e-19 \
 //x=16.48 //y=7.4 //x2=14.905 //y2=5.205
cc_1013 ( N_VDD_c_565_n N_noxref_21_c_4240_n ) capacitor c=0.00289291f \
 //x=16.65 //y=7.4 //x2=14.905 //y2=5.205
cc_1014 ( N_VDD_M35_noxref_d N_noxref_21_c_4240_n ) capacitor c=0.0119951f \
 //x=14.405 //y=5.02 //x2=14.905 //y2=5.205
cc_1015 ( N_VDD_c_564_n N_noxref_21_c_4245_n ) capacitor c=0.0628444f \
 //x=13.32 //y=7.4 //x2=14.195 //y2=5.205
cc_1016 ( N_VDD_M34_noxref_d N_noxref_21_c_4245_n ) capacitor c=0.00269577f \
 //x=12.51 //y=5.02 //x2=14.195 //y2=5.205
cc_1017 ( N_VDD_c_558_n N_noxref_21_c_4247_n ) capacitor c=0.0023707f \
 //x=38.48 //y=7.4 //x2=15.785 //y2=6.905
cc_1018 ( N_VDD_c_573_p N_noxref_21_c_4248_n ) capacitor c=0.0158372f \
 //x=38.48 //y=7.4 //x2=15.075 //y2=6.905
cc_1019 ( N_VDD_c_664_p N_noxref_21_c_4248_n ) capacitor c=0.0604917f \
 //x=16.48 //y=7.4 //x2=15.075 //y2=6.905
cc_1020 ( N_VDD_c_573_p N_noxref_21_M35_noxref_s ) capacitor c=0.00227333f \
 //x=38.48 //y=7.4 //x2=13.975 //y2=5.02
cc_1021 ( N_VDD_c_663_p N_noxref_21_M35_noxref_s ) capacitor c=0.00993188f \
 //x=14.465 //y=7.4 //x2=13.975 //y2=5.02
cc_1022 ( N_VDD_M35_noxref_d N_noxref_21_M35_noxref_s ) capacitor c=0.061257f \
 //x=14.405 //y=5.02 //x2=13.975 //y2=5.02
cc_1023 ( N_VDD_c_564_n N_noxref_21_M36_noxref_d ) capacitor c=0.00130916f \
 //x=13.32 //y=7.4 //x2=14.845 //y2=5.02
cc_1024 ( N_VDD_M35_noxref_d N_noxref_21_M36_noxref_d ) capacitor c=0.0659925f \
 //x=14.405 //y=5.02 //x2=14.845 //y2=5.02
cc_1025 ( N_VDD_c_565_n N_noxref_21_M38_noxref_d ) capacitor c=0.0520312f \
 //x=16.65 //y=7.4 //x2=15.725 //y2=5.02
cc_1026 ( N_VDD_M35_noxref_d N_noxref_21_M38_noxref_d ) capacitor \
 c=0.00107819f //x=14.405 //y=5.02 //x2=15.725 //y2=5.02
cc_1027 ( N_VDD_c_573_p N_noxref_23_c_4326_n ) capacitor c=0.00437344f \
 //x=38.48 //y=7.4 //x2=18.235 //y2=5.205
cc_1028 ( N_VDD_c_665_p N_noxref_23_c_4326_n ) capacitor c=4.49935e-19 \
 //x=17.795 //y=7.4 //x2=18.235 //y2=5.205
cc_1029 ( N_VDD_c_666_p N_noxref_23_c_4326_n ) capacitor c=4.49935e-19 \
 //x=19.81 //y=7.4 //x2=18.235 //y2=5.205
cc_1030 ( N_VDD_c_566_n N_noxref_23_c_4326_n ) capacitor c=0.00289291f \
 //x=19.98 //y=7.4 //x2=18.235 //y2=5.205
cc_1031 ( N_VDD_M39_noxref_d N_noxref_23_c_4326_n ) capacitor c=0.0119951f \
 //x=17.735 //y=5.02 //x2=18.235 //y2=5.205
cc_1032 ( N_VDD_c_565_n N_noxref_23_c_4331_n ) capacitor c=0.0628444f \
 //x=16.65 //y=7.4 //x2=17.525 //y2=5.205
cc_1033 ( N_VDD_c_558_n N_noxref_23_c_4332_n ) capacitor c=0.0023707f \
 //x=38.48 //y=7.4 //x2=19.115 //y2=6.905
cc_1034 ( N_VDD_c_573_p N_noxref_23_c_4333_n ) capacitor c=0.0158566f \
 //x=38.48 //y=7.4 //x2=18.405 //y2=6.905
cc_1035 ( N_VDD_c_666_p N_noxref_23_c_4333_n ) capacitor c=0.0604917f \
 //x=19.81 //y=7.4 //x2=18.405 //y2=6.905
cc_1036 ( N_VDD_c_573_p N_noxref_23_M39_noxref_s ) capacitor c=0.00227333f \
 //x=38.48 //y=7.4 //x2=17.305 //y2=5.02
cc_1037 ( N_VDD_c_665_p N_noxref_23_M39_noxref_s ) capacitor c=0.00993188f \
 //x=17.795 //y=7.4 //x2=17.305 //y2=5.02
cc_1038 ( N_VDD_M39_noxref_d N_noxref_23_M39_noxref_s ) capacitor c=0.061257f \
 //x=17.735 //y=5.02 //x2=17.305 //y2=5.02
cc_1039 ( N_VDD_c_565_n N_noxref_23_M40_noxref_d ) capacitor c=0.00130916f \
 //x=16.65 //y=7.4 //x2=18.175 //y2=5.02
cc_1040 ( N_VDD_M39_noxref_d N_noxref_23_M40_noxref_d ) capacitor c=0.0659925f \
 //x=17.735 //y=5.02 //x2=18.175 //y2=5.02
cc_1041 ( N_VDD_c_566_n N_noxref_23_M42_noxref_d ) capacitor c=0.0520312f \
 //x=19.98 //y=7.4 //x2=19.055 //y2=5.02
cc_1042 ( N_VDD_M39_noxref_d N_noxref_23_M42_noxref_d ) capacitor \
 c=0.00107819f //x=17.735 //y=5.02 //x2=19.055 //y2=5.02
cc_1043 ( N_VDD_M43_noxref_s N_noxref_23_M42_noxref_d ) capacitor \
 c=0.00230193f //x=20.52 //y=5.02 //x2=19.055 //y2=5.02
cc_1044 ( N_VDD_c_573_p N_noxref_27_c_4525_n ) capacitor c=0.00464568f \
 //x=38.48 //y=7.4 //x2=34.885 //y2=5.21
cc_1045 ( N_VDD_c_935_p N_noxref_27_c_4525_n ) capacitor c=4.37585e-19 \
 //x=34.445 //y=7.4 //x2=34.885 //y2=5.21
cc_1046 ( N_VDD_c_938_p N_noxref_27_c_4525_n ) capacitor c=4.37585e-19 \
 //x=36.46 //y=7.4 //x2=34.885 //y2=5.21
cc_1047 ( N_VDD_c_572_n N_noxref_27_c_4525_n ) capacitor c=0.00289291f \
 //x=36.63 //y=7.4 //x2=34.885 //y2=5.21
cc_1048 ( N_VDD_M57_noxref_d N_noxref_27_c_4525_n ) capacitor c=0.0128169f \
 //x=34.385 //y=5.025 //x2=34.885 //y2=5.21
cc_1049 ( N_VDD_c_571_n N_noxref_27_c_4530_n ) capacitor c=0.0669114f //x=33.3 \
 //y=7.4 //x2=34.175 //y2=5.21
cc_1050 ( N_VDD_M56_noxref_d N_noxref_27_c_4530_n ) capacitor c=0.00289186f \
 //x=32.49 //y=5.02 //x2=34.175 //y2=5.21
cc_1051 ( N_VDD_c_558_n N_noxref_27_c_4532_n ) capacitor c=0.00243146f \
 //x=38.48 //y=7.4 //x2=35.765 //y2=6.91
cc_1052 ( N_VDD_c_573_p N_noxref_27_c_4533_n ) capacitor c=0.0321225f \
 //x=38.48 //y=7.4 //x2=35.055 //y2=6.91
cc_1053 ( N_VDD_c_938_p N_noxref_27_c_4533_n ) capacitor c=0.0586694f \
 //x=36.46 //y=7.4 //x2=35.055 //y2=6.91
cc_1054 ( N_VDD_c_573_p N_noxref_27_M57_noxref_s ) capacitor c=0.00579087f \
 //x=38.48 //y=7.4 //x2=33.955 //y2=5.025
cc_1055 ( N_VDD_c_935_p N_noxref_27_M57_noxref_s ) capacitor c=0.0141117f \
 //x=34.445 //y=7.4 //x2=33.955 //y2=5.025
cc_1056 ( N_VDD_M57_noxref_d N_noxref_27_M57_noxref_s ) capacitor c=0.0667021f \
 //x=34.385 //y=5.025 //x2=33.955 //y2=5.025
cc_1057 ( N_VDD_c_571_n N_noxref_27_M58_noxref_d ) capacitor c=8.88629e-19 \
 //x=33.3 //y=7.4 //x2=34.825 //y2=5.025
cc_1058 ( N_VDD_M57_noxref_d N_noxref_27_M58_noxref_d ) capacitor c=0.0659925f \
 //x=34.385 //y=5.025 //x2=34.825 //y2=5.025
cc_1059 ( N_VDD_c_572_n N_noxref_27_M60_noxref_d ) capacitor c=0.0520312f \
 //x=36.63 //y=7.4 //x2=35.705 //y2=5.025
cc_1060 ( N_VDD_M57_noxref_d N_noxref_27_M60_noxref_d ) capacitor \
 c=0.00107819f //x=34.385 //y=5.025 //x2=35.705 //y2=5.025
cc_1061 ( N_VDD_M61_noxref_s N_noxref_27_M60_noxref_d ) capacitor \
 c=0.00226909f //x=37.17 //y=5.02 //x2=35.705 //y2=5.025
cc_1062 ( N_VDD_c_558_n COUT ) capacitor c=0.0232778f //x=38.48 //y=7.4 \
 //x2=38.11 //y2=2.22
cc_1063 ( N_VDD_c_572_n COUT ) capacitor c=4.80934e-19 //x=36.63 //y=7.4 \
 //x2=38.11 //y2=2.22
cc_1064 ( N_VDD_c_573_p N_COUT_c_4578_n ) capacitor c=0.00190861f //x=38.48 \
 //y=7.4 //x2=38.025 //y2=4.58
cc_1065 ( N_VDD_c_980_p N_COUT_c_4578_n ) capacitor c=8.8179e-19 //x=38.1 \
 //y=7.4 //x2=38.025 //y2=4.58
cc_1066 ( N_VDD_M62_noxref_d N_COUT_c_4578_n ) capacitor c=0.00641434f \
 //x=38.04 //y=5.02 //x2=38.025 //y2=4.58
cc_1067 ( N_VDD_c_572_n N_COUT_c_4581_n ) capacitor c=0.017572f //x=36.63 \
 //y=7.4 //x2=37.83 //y2=4.58
cc_1068 ( N_VDD_c_573_p N_COUT_M61_noxref_d ) capacitor c=0.00708604f \
 //x=38.48 //y=7.4 //x2=37.6 //y2=5.02
cc_1069 ( N_VDD_c_980_p N_COUT_M61_noxref_d ) capacitor c=0.0139004f //x=38.1 \
 //y=7.4 //x2=37.6 //y2=5.02
cc_1070 ( N_VDD_c_558_n N_COUT_M61_noxref_d ) capacitor c=0.0205533f //x=38.48 \
 //y=7.4 //x2=37.6 //y2=5.02
cc_1071 ( N_VDD_M61_noxref_s N_COUT_M61_noxref_d ) capacitor c=0.0843065f \
 //x=37.17 //y=5.02 //x2=37.6 //y2=5.02
cc_1072 ( N_VDD_M62_noxref_d N_COUT_M61_noxref_d ) capacitor c=0.0832641f \
 //x=38.04 //y=5.02 //x2=37.6 //y2=5.02
cc_1073 ( N_A_c_1088_n N_noxref_4_c_1465_n ) capacitor c=0.0423564f //x=3.215 \
 //y=4.07 //x2=7.655 //y2=2.59
cc_1074 ( N_A_c_1092_n N_noxref_4_c_1465_n ) capacitor c=0.0288754f //x=3.33 \
 //y=2.105 //x2=7.655 //y2=2.59
cc_1075 ( N_A_c_1094_n N_noxref_4_c_1465_n ) capacitor c=0.190545f //x=29.515 \
 //y=1.85 //x2=7.655 //y2=2.59
cc_1076 ( A N_noxref_4_c_1465_n ) capacitor c=0.0232301f //x=3.33 //y=2.96 \
 //x2=7.655 //y2=2.59
cc_1077 ( A N_noxref_4_c_1465_n ) capacitor c=0.00540955f //x=3.33 //y=2.22 \
 //x2=7.655 //y2=2.59
cc_1078 ( N_A_c_1157_n N_noxref_4_c_1465_n ) capacitor c=0.00162683f //x=3.135 \
 //y=1.92 //x2=7.655 //y2=2.59
cc_1079 ( N_A_c_1088_n N_noxref_4_c_1471_n ) capacitor c=0.00521938f //x=3.215 \
 //y=4.07 //x2=1.595 //y2=2.59
cc_1080 ( N_A_c_1142_n N_noxref_4_c_1471_n ) capacitor c=0.00735597f //x=0.74 \
 //y=2.085 //x2=1.595 //y2=2.59
cc_1081 ( A N_noxref_4_c_1474_n ) capacitor c=4.60786e-19 //x=3.33 //y=2.22 \
 //x2=1.395 //y2=2.08
cc_1082 ( N_A_c_1212_p N_noxref_4_c_1474_n ) capacitor c=0.0023507f //x=1.225 \
 //y=1.41 //x2=1.395 //y2=2.08
cc_1083 ( N_A_c_1088_n N_noxref_4_c_1514_n ) capacitor c=0.0023373f //x=3.215 \
 //y=4.07 //x2=1.195 //y2=2.08
cc_1084 ( N_A_c_1163_n N_noxref_4_c_1514_n ) capacitor c=0.0136603f //x=0.74 \
 //y=2.085 //x2=1.195 //y2=2.08
cc_1085 ( N_A_c_1199_n N_noxref_4_c_1488_n ) capacitor c=0.0099173f //x=1.26 \
 //y=4.79 //x2=1.395 //y2=4.58
cc_1086 ( N_A_c_1088_n N_noxref_4_c_1491_n ) capacitor c=0.0123666f //x=3.215 \
 //y=4.07 //x2=1.2 //y2=4.58
cc_1087 ( N_A_c_1142_n N_noxref_4_c_1491_n ) capacitor c=0.0250789f //x=0.74 \
 //y=2.085 //x2=1.2 //y2=4.58
cc_1088 ( N_A_c_1200_n N_noxref_4_c_1491_n ) capacitor c=0.00962086f //x=0.97 \
 //y=4.79 //x2=1.2 //y2=4.58
cc_1089 ( N_A_c_1088_n N_noxref_4_c_1477_n ) capacitor c=0.0269755f //x=3.215 \
 //y=4.07 //x2=1.48 //y2=2.59
cc_1090 ( N_A_c_1090_n N_noxref_4_c_1477_n ) capacitor c=0.00101501f //x=0.855 \
 //y=4.07 //x2=1.48 //y2=2.59
cc_1091 ( A N_noxref_4_c_1477_n ) capacitor c=0.0158483f //x=3.33 //y=2.96 \
 //x2=1.48 //y2=2.59
cc_1092 ( N_A_c_1142_n N_noxref_4_c_1477_n ) capacitor c=0.0684999f //x=0.74 \
 //y=2.085 //x2=1.48 //y2=2.59
cc_1093 ( N_A_c_1163_n N_noxref_4_c_1477_n ) capacitor c=5.85261e-19 //x=0.74 \
 //y=2.085 //x2=1.48 //y2=2.59
cc_1094 ( N_A_c_1094_n N_noxref_4_c_1480_n ) capacitor c=0.00379578f \
 //x=29.515 //y=1.85 //x2=7.77 //y2=2.085
cc_1095 ( N_A_c_1094_n N_noxref_4_c_1526_n ) capacitor c=0.0120069f //x=29.515 \
 //y=1.85 //x2=7.435 //y2=1.92
cc_1096 ( N_A_c_1094_n N_noxref_4_c_1527_n ) capacitor c=2.55476e-19 \
 //x=29.515 //y=1.85 //x2=7.81 //y2=1.41
cc_1097 ( N_A_c_1142_n N_noxref_4_M0_noxref_d ) capacitor c=0.0178551f \
 //x=0.74 //y=2.085 //x2=0.925 //y2=0.91
cc_1098 ( N_A_c_1147_n N_noxref_4_M0_noxref_d ) capacitor c=0.00218556f \
 //x=0.85 //y=0.91 //x2=0.925 //y2=0.91
cc_1099 ( N_A_c_1229_p N_noxref_4_M0_noxref_d ) capacitor c=0.00347355f \
 //x=0.85 //y=1.255 //x2=0.925 //y2=0.91
cc_1100 ( N_A_c_1230_p N_noxref_4_M0_noxref_d ) capacitor c=0.00742431f \
 //x=0.85 //y=1.565 //x2=0.925 //y2=0.91
cc_1101 ( N_A_c_1149_n N_noxref_4_M0_noxref_d ) capacitor c=0.00784742f \
 //x=0.85 //y=1.92 //x2=0.925 //y2=0.91
cc_1102 ( N_A_c_1150_n N_noxref_4_M0_noxref_d ) capacitor c=0.00220879f \
 //x=1.225 //y=0.755 //x2=0.925 //y2=0.91
cc_1103 ( N_A_c_1212_p N_noxref_4_M0_noxref_d ) capacitor c=0.0138447f \
 //x=1.225 //y=1.41 //x2=0.925 //y2=0.91
cc_1104 ( N_A_c_1151_n N_noxref_4_M0_noxref_d ) capacitor c=0.00218624f \
 //x=1.38 //y=0.91 //x2=0.925 //y2=0.91
cc_1105 ( N_A_c_1153_n N_noxref_4_M0_noxref_d ) capacitor c=0.00601286f \
 //x=1.38 //y=1.255 //x2=0.925 //y2=0.91
cc_1106 ( N_A_M21_noxref_g N_noxref_4_M21_noxref_d ) capacitor c=0.0219309f \
 //x=0.895 //y=6.02 //x2=0.97 //y2=5.02
cc_1107 ( N_A_M22_noxref_g N_noxref_4_M21_noxref_d ) capacitor c=0.021902f \
 //x=1.335 //y=6.02 //x2=0.97 //y2=5.02
cc_1108 ( N_A_c_1199_n N_noxref_4_M21_noxref_d ) capacitor c=0.0146106f \
 //x=1.26 //y=4.79 //x2=0.97 //y2=5.02
cc_1109 ( N_A_c_1200_n N_noxref_4_M21_noxref_d ) capacitor c=0.00307344f \
 //x=0.97 //y=4.79 //x2=0.97 //y2=5.02
cc_1110 ( N_A_c_1088_n N_noxref_5_c_1651_n ) capacitor c=0.0159617f //x=3.215 \
 //y=4.07 //x2=4.555 //y2=4.07
cc_1111 ( A N_noxref_5_c_1651_n ) capacitor c=0.00187343f //x=3.33 //y=2.96 \
 //x2=4.555 //y2=4.07
cc_1112 ( N_A_c_1094_n N_noxref_5_c_1670_n ) capacitor c=0.00856657f \
 //x=29.515 //y=1.85 //x2=9.505 //y2=3.33
cc_1113 ( N_A_c_1088_n N_noxref_5_c_1652_n ) capacitor c=0.00186775f //x=3.215 \
 //y=4.07 //x2=4.44 //y2=4.07
cc_1114 ( A N_noxref_5_c_1652_n ) capacitor c=0.0163266f //x=3.33 //y=2.96 \
 //x2=4.44 //y2=4.07
cc_1115 ( N_A_c_1202_n N_noxref_5_c_1652_n ) capacitor c=0.0022916f //x=3.33 \
 //y=4.7 //x2=4.44 //y2=4.07
cc_1116 ( N_A_c_1094_n N_noxref_5_c_1626_n ) capacitor c=0.00383139f \
 //x=29.515 //y=1.85 //x2=6.66 //y2=2.085
cc_1117 ( A N_noxref_5_c_1626_n ) capacitor c=2.12957e-19 //x=3.33 //y=2.96 \
 //x2=6.66 //y2=2.085
cc_1118 ( N_A_c_1094_n N_noxref_5_c_1629_n ) capacitor c=0.0127014f //x=29.515 \
 //y=1.85 //x2=9.705 //y2=2.08
cc_1119 ( N_A_M23_noxref_g N_noxref_5_M25_noxref_g ) capacitor c=0.0100243f \
 //x=3.23 //y=6.02 //x2=4.11 //y2=6.02
cc_1120 ( N_A_M24_noxref_g N_noxref_5_M25_noxref_g ) capacitor c=0.0610135f \
 //x=3.67 //y=6.02 //x2=4.11 //y2=6.02
cc_1121 ( N_A_M24_noxref_g N_noxref_5_M26_noxref_g ) capacitor c=0.0094155f \
 //x=3.67 //y=6.02 //x2=4.55 //y2=6.02
cc_1122 ( N_A_c_1094_n N_noxref_5_c_1636_n ) capacitor c=0.00970238f \
 //x=29.515 //y=1.85 //x2=6.465 //y2=1.92
cc_1123 ( A N_noxref_5_c_1681_n ) capacitor c=0.00227843f //x=3.33 //y=2.96 \
 //x2=4.44 //y2=4.7
cc_1124 ( N_A_c_1202_n N_noxref_5_c_1681_n ) capacitor c=0.066749f //x=3.33 \
 //y=4.7 //x2=4.44 //y2=4.7
cc_1125 ( N_A_c_1094_n N_noxref_5_M5_noxref_d ) capacitor c=0.0222753f \
 //x=29.515 //y=1.85 //x2=9.795 //y2=0.91
cc_1126 ( N_A_c_1094_n N_B_c_1801_n ) capacitor c=0.0867673f //x=29.515 \
 //y=1.85 //x2=10.245 //y2=2.96
cc_1127 ( A N_B_c_1910_n ) capacitor c=0.00526349f //x=3.33 //y=2.96 \
 //x2=4.555 //y2=2.96
cc_1128 ( N_A_c_1094_n N_B_c_1839_n ) capacitor c=0.0133322f //x=29.515 \
 //y=1.85 //x2=28.745 //y2=4.81
cc_1129 ( A N_B_c_1880_n ) capacitor c=0.00161483f //x=29.6 //y=2.59 \
 //x2=28.86 //y2=4.63
cc_1130 ( N_A_c_1260_p N_B_c_1880_n ) capacitor c=0.003112f //x=29.6 //y=4.535 \
 //x2=28.86 //y2=4.63
cc_1131 ( N_A_c_1261_p N_B_c_1880_n ) capacitor c=3.6528e-19 //x=29.63 //y=4.7 \
 //x2=28.86 //y2=4.63
cc_1132 ( N_A_c_1260_p B ) capacitor c=0.00911664f //x=29.6 //y=4.535 \
 //x2=28.86 //y2=4.81
cc_1133 ( N_A_c_1261_p B ) capacitor c=0.00363571f //x=29.63 //y=4.7 \
 //x2=28.86 //y2=4.81
cc_1134 ( N_A_c_1092_n N_B_c_1803_n ) capacitor c=0.00477139f //x=3.33 \
 //y=2.105 //x2=4.44 //y2=2.085
cc_1135 ( N_A_c_1094_n N_B_c_1803_n ) capacitor c=0.0033965f //x=29.515 \
 //y=1.85 //x2=4.44 //y2=2.085
cc_1136 ( A N_B_c_1803_n ) capacitor c=0.0129698f //x=3.33 //y=2.96 //x2=4.44 \
 //y2=2.085
cc_1137 ( A N_B_c_1803_n ) capacitor c=0.00576402f //x=3.33 //y=2.22 //x2=4.44 \
 //y2=2.085
cc_1138 ( N_A_c_1157_n N_B_c_1803_n ) capacitor c=0.00150155f //x=3.135 \
 //y=1.92 //x2=4.44 //y2=2.085
cc_1139 ( N_A_c_1094_n N_B_c_1805_n ) capacitor c=0.00662949f //x=29.515 \
 //y=1.85 //x2=10.36 //y2=2.085
cc_1140 ( N_A_c_1094_n N_B_c_1810_n ) capacitor c=0.00486413f //x=29.515 \
 //y=1.85 //x2=28.86 //y2=2.08
cc_1141 ( N_A_c_1134_n N_B_c_1810_n ) capacitor c=0.00567525f //x=29.6 \
 //y=2.105 //x2=28.86 //y2=2.08
cc_1142 ( A N_B_c_1810_n ) capacitor c=0.068466f //x=29.6 //y=2.59 //x2=28.86 \
 //y2=2.08
cc_1143 ( A N_B_c_1810_n ) capacitor c=0.010409f //x=29.6 //y=2.22 //x2=28.86 \
 //y2=2.08
cc_1144 ( N_A_c_1274_p N_B_c_1810_n ) capacitor c=0.00302966f //x=29.6 \
 //y=2.08 //x2=28.86 //y2=2.08
cc_1145 ( N_A_M53_noxref_g N_B_M51_noxref_g ) capacitor c=0.0104709f //x=29.64 \
 //y=6.02 //x2=28.76 //y2=6.02
cc_1146 ( N_A_M53_noxref_g N_B_M52_noxref_g ) capacitor c=0.106667f //x=29.64 \
 //y=6.02 //x2=29.2 //y2=6.02
cc_1147 ( N_A_M54_noxref_g N_B_M52_noxref_g ) capacitor c=0.0100341f //x=30.08 \
 //y=6.02 //x2=29.2 //y2=6.02
cc_1148 ( N_A_c_1154_n N_B_c_1931_n ) capacitor c=4.86506e-19 //x=3.135 \
 //y=0.87 //x2=4.105 //y2=0.91
cc_1149 ( N_A_c_1156_n N_B_c_1931_n ) capacitor c=0.00152104f //x=3.135 \
 //y=1.215 //x2=4.105 //y2=0.91
cc_1150 ( N_A_c_1160_n N_B_c_1931_n ) capacitor c=0.0157772f //x=3.665 \
 //y=0.87 //x2=4.105 //y2=0.91
cc_1151 ( N_A_c_1281_p N_B_c_1934_n ) capacitor c=0.00109982f //x=3.135 \
 //y=1.525 //x2=4.105 //y2=1.255
cc_1152 ( N_A_c_1162_n N_B_c_1934_n ) capacitor c=0.0117362f //x=3.665 \
 //y=1.215 //x2=4.105 //y2=1.255
cc_1153 ( N_A_c_1281_p N_B_c_1936_n ) capacitor c=9.57794e-19 //x=3.135 \
 //y=1.525 //x2=4.105 //y2=1.565
cc_1154 ( N_A_c_1157_n N_B_c_1936_n ) capacitor c=0.00581686f //x=3.135 \
 //y=1.92 //x2=4.105 //y2=1.565
cc_1155 ( N_A_c_1162_n N_B_c_1936_n ) capacitor c=0.00862358f //x=3.665 \
 //y=1.215 //x2=4.105 //y2=1.565
cc_1156 ( N_A_c_1092_n N_B_c_1939_n ) capacitor c=2.3323e-19 //x=3.33 \
 //y=2.105 //x2=4.105 //y2=1.92
cc_1157 ( N_A_c_1094_n N_B_c_1939_n ) capacitor c=0.0118904f //x=29.515 \
 //y=1.85 //x2=4.105 //y2=1.92
cc_1158 ( A N_B_c_1939_n ) capacitor c=0.00293774f //x=3.33 //y=2.22 \
 //x2=4.105 //y2=1.92
cc_1159 ( N_A_c_1157_n N_B_c_1939_n ) capacitor c=0.0109942f //x=3.135 \
 //y=1.92 //x2=4.105 //y2=1.92
cc_1160 ( N_A_c_1094_n N_B_c_1943_n ) capacitor c=2.55476e-19 //x=29.515 \
 //y=1.85 //x2=4.48 //y2=1.41
cc_1161 ( N_A_c_1160_n N_B_c_1944_n ) capacitor c=0.00124821f //x=3.665 \
 //y=0.87 //x2=4.635 //y2=0.91
cc_1162 ( N_A_c_1162_n N_B_c_1945_n ) capacitor c=0.00200715f //x=3.665 \
 //y=1.215 //x2=4.635 //y2=1.255
cc_1163 ( N_A_c_1094_n N_B_c_1813_n ) capacitor c=0.00259822f //x=29.515 \
 //y=1.85 //x2=9.72 //y2=1.255
cc_1164 ( N_A_c_1094_n N_B_c_1817_n ) capacitor c=0.00943959f //x=29.515 \
 //y=1.85 //x2=10.25 //y2=1.92
cc_1165 ( N_A_c_1295_p N_B_c_1818_n ) capacitor c=4.86506e-19 //x=29.635 \
 //y=0.905 //x2=28.665 //y2=0.865
cc_1166 ( N_A_c_1295_p N_B_c_1820_n ) capacitor c=0.00152104f //x=29.635 \
 //y=0.905 //x2=28.665 //y2=1.21
cc_1167 ( N_A_c_1297_p N_B_c_1950_n ) capacitor c=0.00109982f //x=29.635 \
 //y=1.25 //x2=28.665 //y2=1.52
cc_1168 ( N_A_c_1298_p N_B_c_1950_n ) capacitor c=9.57794e-19 //x=29.635 \
 //y=1.56 //x2=28.665 //y2=1.52
cc_1169 ( N_A_c_1094_n N_B_c_1821_n ) capacitor c=0.0102404f //x=29.515 \
 //y=1.85 //x2=28.665 //y2=1.915
cc_1170 ( N_A_c_1134_n N_B_c_1821_n ) capacitor c=2.82917e-19 //x=29.6 \
 //y=2.105 //x2=28.665 //y2=1.915
cc_1171 ( A N_B_c_1821_n ) capacitor c=0.00397573f //x=29.6 //y=2.22 \
 //x2=28.665 //y2=1.915
cc_1172 ( N_A_c_1298_p N_B_c_1821_n ) capacitor c=0.00535454f //x=29.635 \
 //y=1.56 //x2=28.665 //y2=1.915
cc_1173 ( N_A_c_1274_p N_B_c_1821_n ) capacitor c=0.0168677f //x=29.6 //y=2.08 \
 //x2=28.665 //y2=1.915
cc_1174 ( N_A_c_1295_p N_B_c_1824_n ) capacitor c=0.0151475f //x=29.635 \
 //y=0.905 //x2=29.195 //y2=0.865
cc_1175 ( N_A_c_1305_p N_B_c_1824_n ) capacitor c=0.00124821f //x=30.165 \
 //y=0.905 //x2=29.195 //y2=0.865
cc_1176 ( N_A_c_1297_p N_B_c_1826_n ) capacitor c=0.0111064f //x=29.635 \
 //y=1.25 //x2=29.195 //y2=1.21
cc_1177 ( N_A_c_1298_p N_B_c_1826_n ) capacitor c=0.00862358f //x=29.635 \
 //y=1.56 //x2=29.195 //y2=1.21
cc_1178 ( N_A_c_1308_p N_B_c_1826_n ) capacitor c=0.00200715f //x=30.165 \
 //y=1.25 //x2=29.195 //y2=1.21
cc_1179 ( N_A_c_1094_n N_B_c_1827_n ) capacitor c=0.00252239f //x=29.515 \
 //y=1.85 //x2=10.25 //y2=2.085
cc_1180 ( N_A_c_1260_p N_B_c_1908_n ) capacitor c=0.00289693f //x=29.6 \
 //y=4.535 //x2=28.86 //y2=4.7
cc_1181 ( N_A_c_1261_p N_B_c_1908_n ) capacitor c=0.0284127f //x=29.63 //y=4.7 \
 //x2=28.86 //y2=4.7
cc_1182 ( A N_noxref_7_c_2272_n ) capacitor c=0.00382596f //x=3.33 //y=2.96 \
 //x2=4.925 //y2=3.7
cc_1183 ( N_A_c_1094_n N_noxref_7_c_2182_n ) capacitor c=0.0228923f //x=29.515 \
 //y=1.85 //x2=11.725 //y2=3.7
cc_1184 ( N_A_c_1094_n N_noxref_7_c_2183_n ) capacitor c=1.06178f //x=29.515 \
 //y=1.85 //x2=23.935 //y2=2.22
cc_1185 ( N_A_c_1094_n N_noxref_7_c_2187_n ) capacitor c=0.0290238f //x=29.515 \
 //y=1.85 //x2=11.955 //y2=2.22
cc_1186 ( N_A_c_1094_n N_noxref_7_c_2188_n ) capacitor c=0.00123405f \
 //x=29.515 //y=1.85 //x2=14.315 //y2=4.07
cc_1187 ( N_A_c_1094_n N_noxref_7_c_2277_n ) capacitor c=0.0177017f //x=29.515 \
 //y=1.85 //x2=4.455 //y2=1.655
cc_1188 ( N_A_c_1094_n N_noxref_7_c_2190_n ) capacitor c=0.0204496f //x=29.515 \
 //y=1.85 //x2=4.81 //y2=3.7
cc_1189 ( A N_noxref_7_c_2190_n ) capacitor c=0.0142305f //x=3.33 //y=2.96 \
 //x2=4.81 //y2=3.7
cc_1190 ( A N_noxref_7_c_2190_n ) capacitor c=6.34057e-19 //x=3.33 //y=2.22 \
 //x2=4.81 //y2=3.7
cc_1191 ( N_A_c_1094_n N_noxref_7_c_2281_n ) capacitor c=0.0177017f //x=29.515 \
 //y=1.85 //x2=7.785 //y2=1.655
cc_1192 ( N_A_c_1094_n N_noxref_7_c_2239_n ) capacitor c=0.0221648f //x=29.515 \
 //y=1.85 //x2=8.14 //y2=3.7
cc_1193 ( N_A_c_1094_n N_noxref_7_c_2193_n ) capacitor c=0.00610431f \
 //x=29.515 //y=1.85 //x2=11.84 //y2=2.085
cc_1194 ( N_A_c_1094_n N_noxref_7_c_2198_n ) capacitor c=0.00258069f \
 //x=29.515 //y=1.85 //x2=14.43 //y2=2.085
cc_1195 ( N_A_c_1094_n N_noxref_7_c_2199_n ) capacitor c=0.00687068f \
 //x=29.515 //y=1.85 //x2=24.05 //y2=2.08
cc_1196 ( N_A_c_1094_n N_noxref_7_c_2203_n ) capacitor c=0.00943959f \
 //x=29.515 //y=1.85 //x2=11.95 //y2=1.92
cc_1197 ( N_A_c_1094_n N_noxref_7_c_2287_n ) capacitor c=0.00265163f \
 //x=29.515 //y=1.85 //x2=12.325 //y2=1.41
cc_1198 ( N_A_c_1094_n N_noxref_7_c_2211_n ) capacitor c=0.00969727f \
 //x=29.515 //y=1.85 //x2=14.235 //y2=1.92
cc_1199 ( N_A_c_1094_n N_noxref_7_c_2289_n ) capacitor c=3.9341e-19 //x=29.515 \
 //y=1.85 //x2=24.46 //y2=1.405
cc_1200 ( N_A_c_1094_n N_noxref_7_c_2217_n ) capacitor c=0.00238027f \
 //x=29.515 //y=1.85 //x2=11.84 //y2=2.085
cc_1201 ( N_A_c_1094_n N_noxref_7_c_2291_n ) capacitor c=0.0023336f //x=29.515 \
 //y=1.85 //x2=24.05 //y2=2.08
cc_1202 ( N_A_c_1094_n N_noxref_7_c_2292_n ) capacitor c=0.00862789f \
 //x=29.515 //y=1.85 //x2=24.05 //y2=1.915
cc_1203 ( N_A_c_1094_n N_noxref_8_c_2602_n ) capacitor c=0.0365096f //x=29.515 \
 //y=1.85 //x2=18.755 //y2=2.59
cc_1204 ( N_A_c_1094_n N_noxref_8_c_2604_n ) capacitor c=0.00172092f \
 //x=29.515 //y=1.85 //x2=12.695 //y2=2.59
cc_1205 ( N_A_c_1094_n N_noxref_8_c_2605_n ) capacitor c=0.0086027f //x=29.515 \
 //y=1.85 //x2=12.495 //y2=2.08
cc_1206 ( N_A_c_1094_n N_noxref_8_c_2610_n ) capacitor c=0.00215939f \
 //x=29.515 //y=1.85 //x2=18.87 //y2=2.085
cc_1207 ( N_A_c_1094_n N_noxref_8_c_2636_n ) capacitor c=0.0115949f //x=29.515 \
 //y=1.85 //x2=18.535 //y2=1.92
cc_1208 ( N_A_c_1094_n N_noxref_8_c_2637_n ) capacitor c=2.55476e-19 \
 //x=29.515 //y=1.85 //x2=18.91 //y2=1.41
cc_1209 ( N_A_c_1094_n N_noxref_8_M6_noxref_d ) capacitor c=0.0221578f \
 //x=29.515 //y=1.85 //x2=12.025 //y2=0.91
cc_1210 ( N_A_c_1094_n SUM ) capacitor c=0.0183046f //x=29.515 //y=1.85 \
 //x2=15.91 //y2=3.33
cc_1211 ( N_A_c_1094_n SUM ) capacitor c=0.0183046f //x=29.515 //y=1.85 \
 //x2=19.24 //y2=2.59
cc_1212 ( N_A_c_1094_n N_SUM_c_2792_n ) capacitor c=0.0177017f //x=29.515 \
 //y=1.85 //x2=15.555 //y2=1.655
cc_1213 ( N_A_c_1094_n N_SUM_c_2793_n ) capacitor c=0.0177017f //x=29.515 \
 //y=1.85 //x2=18.885 //y2=1.655
cc_1214 ( N_A_c_1094_n N_noxref_10_c_2913_n ) capacitor c=0.00257101f \
 //x=29.515 //y=1.85 //x2=17.76 //y2=2.085
cc_1215 ( N_A_c_1094_n N_noxref_10_c_2916_n ) capacitor c=0.0086027f \
 //x=29.515 //y=1.85 //x2=20.805 //y2=2.08
cc_1216 ( N_A_c_1094_n N_noxref_10_c_2923_n ) capacitor c=0.00969727f \
 //x=29.515 //y=1.85 //x2=17.565 //y2=1.92
cc_1217 ( N_A_c_1094_n N_noxref_10_M11_noxref_d ) capacitor c=0.0221578f \
 //x=29.515 //y=1.85 //x2=20.895 //y2=0.91
cc_1218 ( N_A_c_1094_n N_CIN_c_3085_n ) capacitor c=0.00999647f //x=29.515 \
 //y=1.85 //x2=21.345 //y2=2.96
cc_1219 ( N_A_c_1094_n N_CIN_c_3087_n ) capacitor c=0.00350019f //x=29.515 \
 //y=1.85 //x2=23.195 //y2=4.44
cc_1220 ( N_A_c_1094_n N_CIN_c_3088_n ) capacitor c=0.00214372f //x=29.515 \
 //y=1.85 //x2=15.54 //y2=2.085
cc_1221 ( N_A_c_1094_n N_CIN_c_3090_n ) capacitor c=0.00433908f //x=29.515 \
 //y=1.85 //x2=21.46 //y2=2.085
cc_1222 ( N_A_c_1094_n N_CIN_c_3095_n ) capacitor c=0.00269974f //x=29.515 \
 //y=1.85 //x2=23.31 //y2=2.08
cc_1223 ( N_A_c_1094_n N_CIN_c_3150_n ) capacitor c=0.0115949f //x=29.515 \
 //y=1.85 //x2=15.205 //y2=1.92
cc_1224 ( N_A_c_1094_n N_CIN_c_3151_n ) capacitor c=2.55476e-19 //x=29.515 \
 //y=1.85 //x2=15.58 //y2=1.41
cc_1225 ( N_A_c_1094_n N_CIN_c_3098_n ) capacitor c=0.00265163f //x=29.515 \
 //y=1.85 //x2=20.82 //y2=1.255
cc_1226 ( N_A_c_1094_n N_CIN_c_3102_n ) capacitor c=0.00943959f //x=29.515 \
 //y=1.85 //x2=21.35 //y2=1.92
cc_1227 ( N_A_c_1094_n N_CIN_c_3106_n ) capacitor c=0.00968474f //x=29.515 \
 //y=1.85 //x2=23.115 //y2=1.915
cc_1228 ( N_A_c_1094_n N_CIN_c_3112_n ) capacitor c=0.00242142f //x=29.515 \
 //y=1.85 //x2=21.35 //y2=2.085
cc_1229 ( N_A_c_1094_n N_noxref_12_c_3336_n ) capacitor c=0.0312312f \
 //x=29.515 //y=1.85 //x2=26.155 //y2=3.33
cc_1230 ( N_A_c_1094_n N_noxref_12_c_3394_n ) capacitor c=0.00507444f \
 //x=29.515 //y=1.85 //x2=24.905 //y2=3.33
cc_1231 ( N_A_c_1094_n N_noxref_12_c_3395_n ) capacitor c=0.0218297f \
 //x=29.515 //y=1.85 //x2=24.435 //y2=1.655
cc_1232 ( N_A_c_1094_n N_noxref_12_c_3368_n ) capacitor c=0.0233185f \
 //x=29.515 //y=1.85 //x2=24.79 //y2=3.33
cc_1233 ( N_A_c_1094_n N_noxref_12_c_3339_n ) capacitor c=0.00719687f \
 //x=29.515 //y=1.85 //x2=26.27 //y2=2.085
cc_1234 ( N_A_c_1094_n N_noxref_12_c_3346_n ) capacitor c=0.00943959f \
 //x=29.515 //y=1.85 //x2=26.38 //y2=1.92
cc_1235 ( N_A_c_1094_n N_noxref_12_c_3399_n ) capacitor c=0.00259822f \
 //x=29.515 //y=1.85 //x2=26.755 //y2=1.41
cc_1236 ( N_A_c_1094_n N_noxref_12_c_3351_n ) capacitor c=0.0029079f \
 //x=29.515 //y=1.85 //x2=26.27 //y2=2.085
cc_1237 ( A N_noxref_13_c_3500_n ) capacitor c=0.00502038f //x=29.6 //y=2.59 \
 //x2=30.455 //y2=3.33
cc_1238 ( A N_noxref_13_c_3502_n ) capacitor c=8.04589e-19 //x=29.6 //y=2.22 \
 //x2=29.775 //y2=5.2
cc_1239 ( N_A_c_1260_p N_noxref_13_c_3502_n ) capacitor c=0.0131536f //x=29.6 \
 //y=4.535 //x2=29.775 //y2=5.2
cc_1240 ( N_A_M53_noxref_g N_noxref_13_c_3502_n ) capacitor c=0.0166421f \
 //x=29.64 //y=6.02 //x2=29.775 //y2=5.2
cc_1241 ( N_A_c_1261_p N_noxref_13_c_3502_n ) capacitor c=0.00339598f \
 //x=29.63 //y=4.7 //x2=29.775 //y2=5.2
cc_1242 ( N_A_M54_noxref_g N_noxref_13_c_3508_n ) capacitor c=0.0215633f \
 //x=30.08 //y=6.02 //x2=30.255 //y2=5.2
cc_1243 ( N_A_c_1373_p N_noxref_13_c_3475_n ) capacitor c=0.00359704f \
 //x=30.01 //y=1.405 //x2=30.255 //y2=1.655
cc_1244 ( N_A_c_1308_p N_noxref_13_c_3475_n ) capacitor c=0.00457401f \
 //x=30.165 //y=1.25 //x2=30.255 //y2=1.655
cc_1245 ( N_A_c_1094_n N_noxref_13_c_3477_n ) capacitor c=0.0076924f \
 //x=29.515 //y=1.85 //x2=30.34 //y2=3.33
cc_1246 ( N_A_c_1134_n N_noxref_13_c_3477_n ) capacitor c=0.00253269f //x=29.6 \
 //y=2.105 //x2=30.34 //y2=3.33
cc_1247 ( A N_noxref_13_c_3477_n ) capacitor c=0.067502f //x=29.6 //y=2.59 \
 //x2=30.34 //y2=3.33
cc_1248 ( A N_noxref_13_c_3477_n ) capacitor c=0.0118048f //x=29.6 //y=2.22 \
 //x2=30.34 //y2=3.33
cc_1249 ( N_A_c_1260_p N_noxref_13_c_3477_n ) capacitor c=0.00982279f //x=29.6 \
 //y=4.535 //x2=30.34 //y2=3.33
cc_1250 ( N_A_c_1380_p N_noxref_13_c_3477_n ) capacitor c=0.0122366f \
 //x=30.005 //y=4.79 //x2=30.34 //y2=3.33
cc_1251 ( N_A_c_1274_p N_noxref_13_c_3477_n ) capacitor c=0.00522025f //x=29.6 \
 //y=2.08 //x2=30.34 //y2=3.33
cc_1252 ( N_A_c_1382_p N_noxref_13_c_3477_n ) capacitor c=0.00264698f //x=29.6 \
 //y=1.915 //x2=30.34 //y2=3.33
cc_1253 ( N_A_c_1261_p N_noxref_13_c_3477_n ) capacitor c=0.00392192f \
 //x=29.63 //y=4.7 //x2=30.34 //y2=3.33
cc_1254 ( A N_noxref_13_c_3478_n ) capacitor c=0.00113455f //x=29.6 //y=2.59 \
 //x2=31.82 //y2=2.085
cc_1255 ( N_A_c_1380_p N_noxref_13_c_3554_n ) capacitor c=0.00421574f \
 //x=30.005 //y=4.79 //x2=29.86 //y2=5.2
cc_1256 ( N_A_c_1295_p N_noxref_13_M16_noxref_d ) capacitor c=0.00217566f \
 //x=29.635 //y=0.905 //x2=29.71 //y2=0.905
cc_1257 ( N_A_c_1297_p N_noxref_13_M16_noxref_d ) capacitor c=0.0034598f \
 //x=29.635 //y=1.25 //x2=29.71 //y2=0.905
cc_1258 ( N_A_c_1298_p N_noxref_13_M16_noxref_d ) capacitor c=0.00663299f \
 //x=29.635 //y=1.56 //x2=29.71 //y2=0.905
cc_1259 ( N_A_c_1389_p N_noxref_13_M16_noxref_d ) capacitor c=0.00241102f \
 //x=30.01 //y=0.75 //x2=29.71 //y2=0.905
cc_1260 ( N_A_c_1373_p N_noxref_13_M16_noxref_d ) capacitor c=0.0138845f \
 //x=30.01 //y=1.405 //x2=29.71 //y2=0.905
cc_1261 ( N_A_c_1305_p N_noxref_13_M16_noxref_d ) capacitor c=0.00132245f \
 //x=30.165 //y=0.905 //x2=29.71 //y2=0.905
cc_1262 ( N_A_c_1308_p N_noxref_13_M16_noxref_d ) capacitor c=0.00566463f \
 //x=30.165 //y=1.25 //x2=29.71 //y2=0.905
cc_1263 ( N_A_c_1382_p N_noxref_13_M16_noxref_d ) capacitor c=0.00660593f \
 //x=29.6 //y=1.915 //x2=29.71 //y2=0.905
cc_1264 ( N_A_M53_noxref_g N_noxref_13_M53_noxref_d ) capacitor c=0.0173476f \
 //x=29.64 //y=6.02 //x2=29.715 //y2=5.02
cc_1265 ( N_A_M54_noxref_g N_noxref_13_M53_noxref_d ) capacitor c=0.0179769f \
 //x=30.08 //y=6.02 //x2=29.715 //y2=5.02
cc_1266 ( N_A_c_1094_n N_noxref_14_c_3617_n ) capacitor c=0.0652984f \
 //x=29.515 //y=1.85 //x2=34.295 //y2=2.96
cc_1267 ( N_A_c_1134_n N_noxref_14_c_3617_n ) capacitor c=0.0129385f //x=29.6 \
 //y=2.105 //x2=34.295 //y2=2.96
cc_1268 ( A N_noxref_14_c_3617_n ) capacitor c=0.0245919f //x=29.6 //y=2.59 \
 //x2=34.295 //y2=2.96
cc_1269 ( A N_noxref_14_c_3617_n ) capacitor c=0.00326621f //x=29.6 //y=2.22 \
 //x2=34.295 //y2=2.96
cc_1270 ( N_A_c_1260_p N_noxref_14_c_3617_n ) capacitor c=5.29067e-19 //x=29.6 \
 //y=4.535 //x2=34.295 //y2=2.96
cc_1271 ( N_A_c_1094_n N_noxref_14_c_3675_n ) capacitor c=0.00784532f \
 //x=29.515 //y=1.85 //x2=27.125 //y2=2.96
cc_1272 ( N_A_c_1094_n N_noxref_14_c_3629_n ) capacitor c=0.0139768f \
 //x=29.515 //y=1.85 //x2=26.925 //y2=2.08
cc_1273 ( N_A_c_1094_n N_noxref_14_c_3652_n ) capacitor c=5.58471e-19 \
 //x=29.515 //y=1.85 //x2=26.73 //y2=4.58
cc_1274 ( A N_noxref_14_c_3631_n ) capacitor c=0.00133278f //x=29.6 //y=2.59 \
 //x2=27.01 //y2=2.96
cc_1275 ( N_A_c_1094_n N_noxref_14_M14_noxref_d ) capacitor c=0.0240156f \
 //x=29.515 //y=1.85 //x2=26.455 //y2=0.91
cc_1276 ( N_A_c_1088_n N_noxref_17_c_4059_n ) capacitor c=0.00258051f \
 //x=3.215 //y=4.07 //x2=3.805 //y2=5.205
cc_1277 ( A N_noxref_17_c_4059_n ) capacitor c=0.0120071f //x=3.33 //y=2.96 \
 //x2=3.805 //y2=5.205
cc_1278 ( A N_noxref_17_c_4059_n ) capacitor c=6.10729e-19 //x=3.33 //y=2.22 \
 //x2=3.805 //y2=5.205
cc_1279 ( N_A_M23_noxref_g N_noxref_17_c_4059_n ) capacitor c=0.0190059f \
 //x=3.23 //y=6.02 //x2=3.805 //y2=5.205
cc_1280 ( N_A_M24_noxref_g N_noxref_17_c_4059_n ) capacitor c=0.0198429f \
 //x=3.67 //y=6.02 //x2=3.805 //y2=5.205
cc_1281 ( N_A_c_1202_n N_noxref_17_c_4059_n ) capacitor c=0.00503467f //x=3.33 \
 //y=4.7 //x2=3.805 //y2=5.205
cc_1282 ( N_A_c_1088_n N_noxref_17_c_4064_n ) capacitor c=0.00663113f \
 //x=3.215 //y=4.07 //x2=3.095 //y2=5.205
cc_1283 ( N_A_M23_noxref_g N_noxref_17_M23_noxref_s ) capacitor c=0.0441361f \
 //x=3.23 //y=6.02 //x2=2.875 //y2=5.02
cc_1284 ( N_A_M24_noxref_g N_noxref_17_M24_noxref_d ) capacitor c=0.0170604f \
 //x=3.67 //y=6.02 //x2=3.745 //y2=5.02
cc_1285 ( N_A_c_1157_n N_noxref_18_c_4098_n ) capacitor c=0.0034165f //x=3.135 \
 //y=1.92 //x2=2.915 //y2=1.5
cc_1286 ( N_A_c_1092_n N_noxref_18_c_4099_n ) capacitor c=6.57795e-19 //x=3.33 \
 //y=2.105 //x2=3.8 //y2=1.585
cc_1287 ( N_A_c_1132_n N_noxref_18_c_4099_n ) capacitor c=0.0201754f //x=3.415 \
 //y=1.85 //x2=3.8 //y2=1.585
cc_1288 ( A N_noxref_18_c_4099_n ) capacitor c=0.0133658f //x=3.33 //y=2.22 \
 //x2=3.8 //y2=1.585
cc_1289 ( N_A_c_1281_p N_noxref_18_c_4099_n ) capacitor c=0.00695056f \
 //x=3.135 //y=1.525 //x2=3.8 //y2=1.585
cc_1290 ( N_A_c_1157_n N_noxref_18_c_4099_n ) capacitor c=0.0172357f //x=3.135 \
 //y=1.92 //x2=3.8 //y2=1.585
cc_1291 ( N_A_c_1159_n N_noxref_18_c_4099_n ) capacitor c=0.00771868f //x=3.51 \
 //y=1.37 //x2=3.8 //y2=1.585
cc_1292 ( N_A_c_1162_n N_noxref_18_c_4099_n ) capacitor c=0.0034036f //x=3.665 \
 //y=1.215 //x2=3.8 //y2=1.585
cc_1293 ( N_A_c_1094_n N_noxref_18_c_4106_n ) capacitor c=0.00952696f \
 //x=29.515 //y=1.85 //x2=3.885 //y2=1.5
cc_1294 ( N_A_c_1157_n N_noxref_18_c_4106_n ) capacitor c=6.71402e-19 \
 //x=3.135 //y=1.92 //x2=3.885 //y2=1.5
cc_1295 ( N_A_c_1094_n N_noxref_18_c_4107_n ) capacitor c=0.00479599f \
 //x=29.515 //y=1.85 //x2=4.77 //y2=0.535
cc_1296 ( N_A_c_1094_n N_noxref_18_M1_noxref_s ) capacitor c=0.00162009f \
 //x=29.515 //y=1.85 //x2=2.78 //y2=0.37
cc_1297 ( N_A_c_1154_n N_noxref_18_M1_noxref_s ) capacitor c=0.0326577f \
 //x=3.135 //y=0.87 //x2=2.78 //y2=0.37
cc_1298 ( N_A_c_1281_p N_noxref_18_M1_noxref_s ) capacitor c=3.48408e-19 \
 //x=3.135 //y=1.525 //x2=2.78 //y2=0.37
cc_1299 ( N_A_c_1160_n N_noxref_18_M1_noxref_s ) capacitor c=0.0120759f \
 //x=3.665 //y=0.87 //x2=2.78 //y2=0.37
cc_1300 ( N_A_c_1094_n N_noxref_20_c_4211_n ) capacitor c=0.00952696f \
 //x=29.515 //y=1.85 //x2=6.245 //y2=1.5
cc_1301 ( N_A_c_1094_n N_noxref_20_c_4190_n ) capacitor c=0.0330561f \
 //x=29.515 //y=1.85 //x2=7.13 //y2=1.585
cc_1302 ( N_A_c_1094_n N_noxref_20_c_4197_n ) capacitor c=0.00952696f \
 //x=29.515 //y=1.85 //x2=7.215 //y2=1.5
cc_1303 ( N_A_c_1094_n N_noxref_20_c_4198_n ) capacitor c=0.00479599f \
 //x=29.515 //y=1.85 //x2=8.1 //y2=0.535
cc_1304 ( N_A_c_1094_n N_noxref_20_M3_noxref_s ) capacitor c=0.00162009f \
 //x=29.515 //y=1.85 //x2=6.11 //y2=0.37
cc_1305 ( N_A_c_1094_n N_noxref_22_c_4277_n ) capacitor c=0.00952696f \
 //x=29.515 //y=1.85 //x2=14.015 //y2=1.5
cc_1306 ( N_A_c_1094_n N_noxref_22_c_4278_n ) capacitor c=0.0330561f \
 //x=29.515 //y=1.85 //x2=14.9 //y2=1.585
cc_1307 ( N_A_c_1094_n N_noxref_22_c_4285_n ) capacitor c=0.00952696f \
 //x=29.515 //y=1.85 //x2=14.985 //y2=1.5
cc_1308 ( N_A_c_1094_n N_noxref_22_c_4286_n ) capacitor c=0.00479599f \
 //x=29.515 //y=1.85 //x2=15.87 //y2=0.535
cc_1309 ( N_A_c_1094_n N_noxref_22_M7_noxref_s ) capacitor c=0.00162009f \
 //x=29.515 //y=1.85 //x2=13.88 //y2=0.37
cc_1310 ( N_A_c_1094_n N_noxref_24_c_4386_n ) capacitor c=0.00952696f \
 //x=29.515 //y=1.85 //x2=17.345 //y2=1.5
cc_1311 ( N_A_c_1094_n N_noxref_24_c_4365_n ) capacitor c=0.0330561f \
 //x=29.515 //y=1.85 //x2=18.23 //y2=1.585
cc_1312 ( N_A_c_1094_n N_noxref_24_c_4372_n ) capacitor c=0.00952696f \
 //x=29.515 //y=1.85 //x2=18.315 //y2=1.5
cc_1313 ( N_A_c_1094_n N_noxref_24_c_4373_n ) capacitor c=0.00479599f \
 //x=29.515 //y=1.85 //x2=19.2 //y2=0.535
cc_1314 ( N_A_c_1094_n N_noxref_24_M9_noxref_s ) capacitor c=0.00162009f \
 //x=29.515 //y=1.85 //x2=17.21 //y2=0.37
cc_1315 ( N_A_c_1094_n N_noxref_25_c_4415_n ) capacitor c=0.00946709f \
 //x=29.515 //y=1.85 //x2=22.895 //y2=1.495
cc_1316 ( N_A_c_1094_n N_noxref_25_c_4416_n ) capacitor c=0.0328762f \
 //x=29.515 //y=1.85 //x2=23.78 //y2=1.58
cc_1317 ( N_A_c_1094_n N_noxref_25_c_4423_n ) capacitor c=0.00946709f \
 //x=29.515 //y=1.85 //x2=23.865 //y2=1.495
cc_1318 ( N_A_c_1094_n N_noxref_25_c_4424_n ) capacitor c=0.00329512f \
 //x=29.515 //y=1.85 //x2=24.75 //y2=0.53
cc_1319 ( N_A_c_1094_n N_noxref_25_M12_noxref_s ) capacitor c=0.00161084f \
 //x=29.515 //y=1.85 //x2=22.76 //y2=0.365
cc_1320 ( N_A_c_1094_n N_noxref_26_c_4468_n ) capacitor c=0.00946709f \
 //x=29.515 //y=1.85 //x2=28.445 //y2=1.495
cc_1321 ( N_A_c_1094_n N_noxref_26_c_4469_n ) capacitor c=0.0324418f \
 //x=29.515 //y=1.85 //x2=29.33 //y2=1.58
cc_1322 ( N_A_c_1094_n N_noxref_26_c_4476_n ) capacitor c=0.00799446f \
 //x=29.515 //y=1.85 //x2=29.415 //y2=1.495
cc_1323 ( A N_noxref_26_c_4476_n ) capacitor c=0.00292347f //x=29.6 //y=2.22 \
 //x2=29.415 //y2=1.495
cc_1324 ( N_A_c_1298_p N_noxref_26_c_4476_n ) capacitor c=0.00623646f \
 //x=29.635 //y=1.56 //x2=29.415 //y2=1.495
cc_1325 ( N_A_c_1274_p N_noxref_26_c_4476_n ) capacitor c=8.6727e-19 //x=29.6 \
 //y=2.08 //x2=29.415 //y2=1.495
cc_1326 ( N_A_c_1094_n N_noxref_26_c_4477_n ) capacitor c=0.00150612f \
 //x=29.515 //y=1.85 //x2=30.3 //y2=0.53
cc_1327 ( N_A_c_1134_n N_noxref_26_c_4477_n ) capacitor c=2.37839e-19 //x=29.6 \
 //y=2.105 //x2=30.3 //y2=0.53
cc_1328 ( A N_noxref_26_c_4477_n ) capacitor c=0.00164051f //x=29.6 //y=2.22 \
 //x2=30.3 //y2=0.53
cc_1329 ( N_A_c_1295_p N_noxref_26_c_4477_n ) capacitor c=0.0183476f \
 //x=29.635 //y=0.905 //x2=30.3 //y2=0.53
cc_1330 ( N_A_c_1305_p N_noxref_26_c_4477_n ) capacitor c=0.00656458f \
 //x=30.165 //y=0.905 //x2=30.3 //y2=0.53
cc_1331 ( N_A_c_1274_p N_noxref_26_c_4477_n ) capacitor c=2.1838e-19 //x=29.6 \
 //y=2.08 //x2=30.3 //y2=0.53
cc_1332 ( N_A_c_1295_p N_noxref_26_M15_noxref_s ) capacitor c=0.00623646f \
 //x=29.635 //y=0.905 //x2=28.31 //y2=0.365
cc_1333 ( N_A_c_1305_p N_noxref_26_M15_noxref_s ) capacitor c=0.0143002f \
 //x=30.165 //y=0.905 //x2=28.31 //y2=0.365
cc_1334 ( N_A_c_1308_p N_noxref_26_M15_noxref_s ) capacitor c=0.00290153f \
 //x=30.165 //y=1.25 //x2=28.31 //y2=0.365
cc_1335 ( N_noxref_4_c_1465_n N_noxref_5_c_1646_n ) capacitor c=7.67045e-19 \
 //x=7.655 //y=2.59 //x2=9.505 //y2=4.07
cc_1336 ( N_noxref_4_c_1480_n N_noxref_5_c_1646_n ) capacitor c=0.0166527f \
 //x=7.77 //y=2.085 //x2=9.505 //y2=4.07
cc_1337 ( N_noxref_4_c_1465_n N_noxref_5_c_1651_n ) capacitor c=6.56372e-19 \
 //x=7.655 //y=2.59 //x2=4.555 //y2=4.07
cc_1338 ( N_noxref_4_c_1465_n N_noxref_5_c_1670_n ) capacitor c=0.00949286f \
 //x=7.655 //y=2.59 //x2=9.505 //y2=3.33
cc_1339 ( N_noxref_4_c_1480_n N_noxref_5_c_1670_n ) capacitor c=0.0158195f \
 //x=7.77 //y=2.085 //x2=9.505 //y2=3.33
cc_1340 ( N_noxref_4_c_1465_n N_noxref_5_c_1689_n ) capacitor c=9.78991e-19 \
 //x=7.655 //y=2.59 //x2=6.775 //y2=3.33
cc_1341 ( N_noxref_4_c_1480_n N_noxref_5_c_1689_n ) capacitor c=7.52994e-19 \
 //x=7.77 //y=2.085 //x2=6.775 //y2=3.33
cc_1342 ( N_noxref_4_c_1465_n N_noxref_5_c_1626_n ) capacitor c=0.0224325f \
 //x=7.655 //y=2.59 //x2=6.66 //y2=2.085
cc_1343 ( N_noxref_4_c_1480_n N_noxref_5_c_1626_n ) capacitor c=0.0237286f \
 //x=7.77 //y=2.085 //x2=6.66 //y2=2.085
cc_1344 ( N_noxref_4_c_1526_n N_noxref_5_c_1626_n ) capacitor c=0.00247765f \
 //x=7.435 //y=1.92 //x2=6.66 //y2=2.085
cc_1345 ( N_noxref_4_c_1480_n N_noxref_5_c_1627_n ) capacitor c=0.00187546f \
 //x=7.77 //y=2.085 //x2=9.62 //y2=3.33
cc_1346 ( N_noxref_4_c_1552_p N_noxref_5_c_1632_n ) capacitor c=4.86506e-19 \
 //x=7.435 //y=0.91 //x2=6.465 //y2=0.87
cc_1347 ( N_noxref_4_c_1552_p N_noxref_5_c_1634_n ) capacitor c=0.00152104f \
 //x=7.435 //y=0.91 //x2=6.465 //y2=1.215
cc_1348 ( N_noxref_4_c_1554_p N_noxref_5_c_1635_n ) capacitor c=0.00109982f \
 //x=7.435 //y=1.255 //x2=6.465 //y2=1.525
cc_1349 ( N_noxref_4_c_1555_p N_noxref_5_c_1635_n ) capacitor c=9.57794e-19 \
 //x=7.435 //y=1.565 //x2=6.465 //y2=1.525
cc_1350 ( N_noxref_4_c_1465_n N_noxref_5_c_1636_n ) capacitor c=0.00394879f \
 //x=7.655 //y=2.59 //x2=6.465 //y2=1.92
cc_1351 ( N_noxref_4_c_1480_n N_noxref_5_c_1636_n ) capacitor c=0.00217068f \
 //x=7.77 //y=2.085 //x2=6.465 //y2=1.92
cc_1352 ( N_noxref_4_c_1555_p N_noxref_5_c_1636_n ) capacitor c=0.00531182f \
 //x=7.435 //y=1.565 //x2=6.465 //y2=1.92
cc_1353 ( N_noxref_4_c_1526_n N_noxref_5_c_1636_n ) capacitor c=0.0118933f \
 //x=7.435 //y=1.92 //x2=6.465 //y2=1.92
cc_1354 ( N_noxref_4_c_1552_p N_noxref_5_c_1639_n ) capacitor c=0.0157772f \
 //x=7.435 //y=0.91 //x2=6.995 //y2=0.87
cc_1355 ( N_noxref_4_c_1561_p N_noxref_5_c_1639_n ) capacitor c=0.00124821f \
 //x=7.965 //y=0.91 //x2=6.995 //y2=0.87
cc_1356 ( N_noxref_4_c_1554_p N_noxref_5_c_1641_n ) capacitor c=0.0117362f \
 //x=7.435 //y=1.255 //x2=6.995 //y2=1.215
cc_1357 ( N_noxref_4_c_1555_p N_noxref_5_c_1641_n ) capacitor c=0.00862358f \
 //x=7.435 //y=1.565 //x2=6.995 //y2=1.215
cc_1358 ( N_noxref_4_c_1564_p N_noxref_5_c_1641_n ) capacitor c=0.00200715f \
 //x=7.965 //y=1.255 //x2=6.995 //y2=1.215
cc_1359 ( N_noxref_4_c_1465_n N_B_c_1801_n ) capacitor c=0.300234f //x=7.655 \
 //y=2.59 //x2=10.245 //y2=2.96
cc_1360 ( N_noxref_4_c_1480_n N_B_c_1801_n ) capacitor c=0.0176337f //x=7.77 \
 //y=2.085 //x2=10.245 //y2=2.96
cc_1361 ( N_noxref_4_c_1465_n N_B_c_1910_n ) capacitor c=0.0290321f //x=7.655 \
 //y=2.59 //x2=4.555 //y2=2.96
cc_1362 ( N_noxref_4_c_1480_n N_B_c_1830_n ) capacitor c=0.01781f //x=7.77 \
 //y=2.085 //x2=10.245 //y2=4.44
cc_1363 ( N_noxref_4_c_1569_p N_B_c_1830_n ) capacitor c=0.0105048f //x=7.77 \
 //y=4.7 //x2=10.245 //y2=4.44
cc_1364 ( N_noxref_4_c_1480_n N_B_c_1837_n ) capacitor c=9.41499e-19 //x=7.77 \
 //y=2.085 //x2=6.775 //y2=4.44
cc_1365 ( N_noxref_4_c_1480_n B ) capacitor c=0.0082518f //x=7.77 //y=2.085 \
 //x2=6.66 //y2=4.44
cc_1366 ( N_noxref_4_c_1569_p B ) capacitor c=0.00226398f //x=7.77 //y=4.7 \
 //x2=6.66 //y2=4.44
cc_1367 ( N_noxref_4_c_1465_n N_B_c_1803_n ) capacitor c=0.0198692f //x=7.655 \
 //y=2.59 //x2=4.44 //y2=2.085
cc_1368 ( N_noxref_4_c_1477_n N_B_c_1803_n ) capacitor c=2.14844e-19 //x=1.48 \
 //y=2.59 //x2=4.44 //y2=2.085
cc_1369 ( N_noxref_4_M29_noxref_g N_B_M27_noxref_g ) capacitor c=0.0100243f \
 //x=7.44 //y=6.02 //x2=6.56 //y2=6.02
cc_1370 ( N_noxref_4_M29_noxref_g N_B_M28_noxref_g ) capacitor c=0.0610135f \
 //x=7.44 //y=6.02 //x2=7 //y2=6.02
cc_1371 ( N_noxref_4_M30_noxref_g N_B_M28_noxref_g ) capacitor c=0.0094155f \
 //x=7.88 //y=6.02 //x2=7 //y2=6.02
cc_1372 ( N_noxref_4_c_1465_n N_B_c_1939_n ) capacitor c=0.0049293f //x=7.655 \
 //y=2.59 //x2=4.105 //y2=1.92
cc_1373 ( N_noxref_4_c_1480_n N_B_c_1907_n ) capacitor c=0.0022916f //x=7.77 \
 //y=2.085 //x2=6.66 //y2=4.7
cc_1374 ( N_noxref_4_c_1569_p N_B_c_1907_n ) capacitor c=0.066749f //x=7.77 \
 //y=4.7 //x2=6.66 //y2=4.7
cc_1375 ( N_noxref_4_c_1465_n N_noxref_7_c_2293_n ) capacitor c=0.00619185f \
 //x=7.655 //y=2.59 //x2=8.025 //y2=3.7
cc_1376 ( N_noxref_4_c_1480_n N_noxref_7_c_2293_n ) capacitor c=0.0167028f \
 //x=7.77 //y=2.085 //x2=8.025 //y2=3.7
cc_1377 ( N_noxref_4_c_1465_n N_noxref_7_c_2272_n ) capacitor c=6.30506e-19 \
 //x=7.655 //y=2.59 //x2=4.925 //y2=3.7
cc_1378 ( N_noxref_4_c_1480_n N_noxref_7_c_2272_n ) capacitor c=2.02744e-19 \
 //x=7.77 //y=2.085 //x2=4.925 //y2=3.7
cc_1379 ( N_noxref_4_c_1480_n N_noxref_7_c_2297_n ) capacitor c=0.00153295f \
 //x=7.77 //y=2.085 //x2=8.255 //y2=3.7
cc_1380 ( N_noxref_4_c_1465_n N_noxref_7_c_2233_n ) capacitor c=4.65436e-19 \
 //x=7.655 //y=2.59 //x2=4.415 //y2=5.205
cc_1381 ( N_noxref_4_c_1465_n N_noxref_7_c_2190_n ) capacitor c=0.0167161f \
 //x=7.655 //y=2.59 //x2=4.81 //y2=3.7
cc_1382 ( N_noxref_4_c_1477_n N_noxref_7_c_2190_n ) capacitor c=2.79968e-19 \
 //x=1.48 //y=2.59 //x2=4.81 //y2=3.7
cc_1383 ( N_noxref_4_c_1480_n N_noxref_7_c_2190_n ) capacitor c=0.00277451f \
 //x=7.77 //y=2.085 //x2=4.81 //y2=3.7
cc_1384 ( N_noxref_4_M30_noxref_g N_noxref_7_c_2236_n ) capacitor c=0.0180846f \
 //x=7.88 //y=6.02 //x2=8.055 //y2=5.205
cc_1385 ( N_noxref_4_c_1569_p N_noxref_7_c_2236_n ) capacitor c=0.00161455f \
 //x=7.77 //y=4.7 //x2=8.055 //y2=5.205
cc_1386 ( N_noxref_4_c_1480_n N_noxref_7_c_2238_n ) capacitor c=0.0129715f \
 //x=7.77 //y=2.085 //x2=7.745 //y2=5.205
cc_1387 ( N_noxref_4_M29_noxref_g N_noxref_7_c_2238_n ) capacitor c=0.0132788f \
 //x=7.44 //y=6.02 //x2=7.745 //y2=5.205
cc_1388 ( N_noxref_4_c_1569_p N_noxref_7_c_2238_n ) capacitor c=0.00554627f \
 //x=7.77 //y=4.7 //x2=7.745 //y2=5.205
cc_1389 ( N_noxref_4_c_1526_n N_noxref_7_c_2191_n ) capacitor c=0.00355555f \
 //x=7.435 //y=1.92 //x2=8.055 //y2=1.655
cc_1390 ( N_noxref_4_c_1527_n N_noxref_7_c_2191_n ) capacitor c=0.00196666f \
 //x=7.81 //y=1.41 //x2=8.055 //y2=1.655
cc_1391 ( N_noxref_4_c_1564_p N_noxref_7_c_2191_n ) capacitor c=0.00423452f \
 //x=7.965 //y=1.255 //x2=8.055 //y2=1.655
cc_1392 ( N_noxref_4_c_1480_n N_noxref_7_c_2281_n ) capacitor c=0.0136356f \
 //x=7.77 //y=2.085 //x2=7.785 //y2=1.655
cc_1393 ( N_noxref_4_c_1526_n N_noxref_7_c_2281_n ) capacitor c=0.0062602f \
 //x=7.435 //y=1.92 //x2=7.785 //y2=1.655
cc_1394 ( N_noxref_4_c_1465_n N_noxref_7_c_2239_n ) capacitor c=0.0100753f \
 //x=7.655 //y=2.59 //x2=8.14 //y2=3.7
cc_1395 ( N_noxref_4_c_1480_n N_noxref_7_c_2239_n ) capacitor c=0.187361f \
 //x=7.77 //y=2.085 //x2=8.14 //y2=3.7
cc_1396 ( N_noxref_4_c_1526_n N_noxref_7_c_2239_n ) capacitor c=0.0168114f \
 //x=7.435 //y=1.92 //x2=8.14 //y2=3.7
cc_1397 ( N_noxref_4_c_1569_p N_noxref_7_c_2239_n ) capacitor c=0.0209809f \
 //x=7.77 //y=4.7 //x2=8.14 //y2=3.7
cc_1398 ( N_noxref_4_c_1552_p N_noxref_7_M4_noxref_d ) capacitor c=0.00217566f \
 //x=7.435 //y=0.91 //x2=7.51 //y2=0.91
cc_1399 ( N_noxref_4_c_1554_p N_noxref_7_M4_noxref_d ) capacitor c=0.0034598f \
 //x=7.435 //y=1.255 //x2=7.51 //y2=0.91
cc_1400 ( N_noxref_4_c_1555_p N_noxref_7_M4_noxref_d ) capacitor c=0.00522042f \
 //x=7.435 //y=1.565 //x2=7.51 //y2=0.91
cc_1401 ( N_noxref_4_c_1526_n N_noxref_7_M4_noxref_d ) capacitor c=0.00643086f \
 //x=7.435 //y=1.92 //x2=7.51 //y2=0.91
cc_1402 ( N_noxref_4_c_1608_p N_noxref_7_M4_noxref_d ) capacitor c=0.00241053f \
 //x=7.81 //y=0.755 //x2=7.51 //y2=0.91
cc_1403 ( N_noxref_4_c_1527_n N_noxref_7_M4_noxref_d ) capacitor c=0.0124466f \
 //x=7.81 //y=1.41 //x2=7.51 //y2=0.91
cc_1404 ( N_noxref_4_c_1561_p N_noxref_7_M4_noxref_d ) capacitor c=0.00132245f \
 //x=7.965 //y=0.91 //x2=7.51 //y2=0.91
cc_1405 ( N_noxref_4_c_1564_p N_noxref_7_M4_noxref_d ) capacitor c=0.00566463f \
 //x=7.965 //y=1.255 //x2=7.51 //y2=0.91
cc_1406 ( N_noxref_4_M30_noxref_g N_noxref_7_M29_noxref_d ) capacitor \
 c=0.0136385f //x=7.88 //y=6.02 //x2=7.515 //y2=5.02
cc_1407 ( N_noxref_4_c_1465_n N_noxref_17_c_4059_n ) capacitor c=0.00680306f \
 //x=7.655 //y=2.59 //x2=3.805 //y2=5.205
cc_1408 ( N_noxref_4_c_1465_n N_noxref_18_c_4098_n ) capacitor c=0.00446497f \
 //x=7.655 //y=2.59 //x2=2.915 //y2=1.5
cc_1409 ( N_noxref_4_c_1465_n N_noxref_18_c_4099_n ) capacitor c=0.00494246f \
 //x=7.655 //y=2.59 //x2=3.8 //y2=1.585
cc_1410 ( N_noxref_4_M29_noxref_g N_noxref_19_c_4149_n ) capacitor \
 c=0.0170604f //x=7.44 //y=6.02 //x2=7.135 //y2=5.205
cc_1411 ( N_noxref_4_M29_noxref_g N_noxref_19_c_4155_n ) capacitor \
 c=0.0144401f //x=7.44 //y=6.02 //x2=8.015 //y2=6.905
cc_1412 ( N_noxref_4_M30_noxref_g N_noxref_19_c_4155_n ) capacitor \
 c=0.0163317f //x=7.88 //y=6.02 //x2=8.015 //y2=6.905
cc_1413 ( N_noxref_4_M30_noxref_g N_noxref_19_M30_noxref_d ) capacitor \
 c=0.0351101f //x=7.88 //y=6.02 //x2=7.955 //y2=5.02
cc_1414 ( N_noxref_4_c_1555_p N_noxref_20_c_4197_n ) capacitor c=0.00628626f \
 //x=7.435 //y=1.565 //x2=7.215 //y2=1.5
cc_1415 ( N_noxref_4_c_1552_p N_noxref_20_c_4198_n ) capacitor c=0.0197911f \
 //x=7.435 //y=0.91 //x2=8.1 //y2=0.535
cc_1416 ( N_noxref_4_c_1561_p N_noxref_20_c_4198_n ) capacitor c=0.00655813f \
 //x=7.965 //y=0.91 //x2=8.1 //y2=0.535
cc_1417 ( N_noxref_4_c_1552_p N_noxref_20_M3_noxref_s ) capacitor \
 c=0.00628626f //x=7.435 //y=0.91 //x2=6.11 //y2=0.37
cc_1418 ( N_noxref_4_c_1561_p N_noxref_20_M3_noxref_s ) capacitor c=0.0143002f \
 //x=7.965 //y=0.91 //x2=6.11 //y2=0.37
cc_1419 ( N_noxref_4_c_1564_p N_noxref_20_M3_noxref_s ) capacitor \
 c=0.00290153f //x=7.965 //y=1.255 //x2=6.11 //y2=0.37
cc_1420 ( N_noxref_5_c_1646_n N_B_c_1801_n ) capacitor c=0.01084f //x=9.505 \
 //y=4.07 //x2=10.245 //y2=2.96
cc_1421 ( N_noxref_5_c_1670_n N_B_c_1801_n ) capacitor c=0.269397f //x=9.505 \
 //y=3.33 //x2=10.245 //y2=2.96
cc_1422 ( N_noxref_5_c_1689_n N_B_c_1801_n ) capacitor c=0.0291219f //x=6.775 \
 //y=3.33 //x2=10.245 //y2=2.96
cc_1423 ( N_noxref_5_c_1626_n N_B_c_1801_n ) capacitor c=0.0215791f //x=6.66 \
 //y=2.085 //x2=10.245 //y2=2.96
cc_1424 ( N_noxref_5_c_1627_n N_B_c_1801_n ) capacitor c=0.0251512f //x=9.62 \
 //y=3.33 //x2=10.245 //y2=2.96
cc_1425 ( N_noxref_5_c_1628_n N_B_c_1801_n ) capacitor c=0.00570105f //x=9.905 \
 //y=2.08 //x2=10.245 //y2=2.96
cc_1426 ( N_noxref_5_c_1651_n N_B_c_1910_n ) capacitor c=0.00956028f //x=4.555 \
 //y=4.07 //x2=4.555 //y2=2.96
cc_1427 ( N_noxref_5_c_1652_n N_B_c_1910_n ) capacitor c=2.06418e-19 //x=4.44 \
 //y=4.07 //x2=4.555 //y2=2.96
cc_1428 ( N_noxref_5_c_1646_n N_B_c_1830_n ) capacitor c=0.267726f //x=9.505 \
 //y=4.07 //x2=10.245 //y2=4.44
cc_1429 ( N_noxref_5_c_1627_n N_B_c_1830_n ) capacitor c=0.0131307f //x=9.62 \
 //y=3.33 //x2=10.245 //y2=4.44
cc_1430 ( N_noxref_5_c_1656_n N_B_c_1830_n ) capacitor c=0.0201293f //x=9.9 \
 //y=4.58 //x2=10.245 //y2=4.44
cc_1431 ( N_noxref_5_c_1657_n N_B_c_1830_n ) capacitor c=0.00582322f //x=9.705 \
 //y=4.58 //x2=10.245 //y2=4.44
cc_1432 ( N_noxref_5_c_1646_n N_B_c_1837_n ) capacitor c=0.0286083f //x=9.505 \
 //y=4.07 //x2=6.775 //y2=4.44
cc_1433 ( N_noxref_5_M31_noxref_d N_B_c_1876_n ) capacitor c=0.00766276f \
 //x=9.84 //y=5.02 //x2=10.475 //y2=4.81
cc_1434 ( N_noxref_5_c_1646_n B ) capacitor c=0.00480464f //x=9.505 //y=4.07 \
 //x2=6.66 //y2=4.44
cc_1435 ( N_noxref_5_c_1626_n B ) capacitor c=0.00883142f //x=6.66 //y=2.085 \
 //x2=6.66 //y2=4.44
cc_1436 ( N_noxref_5_c_1651_n N_B_c_1803_n ) capacitor c=2.06418e-19 //x=4.555 \
 //y=4.07 //x2=4.44 //y2=2.085
cc_1437 ( N_noxref_5_c_1652_n N_B_c_1803_n ) capacitor c=0.00912271f //x=4.44 \
 //y=4.07 //x2=4.44 //y2=2.085
cc_1438 ( N_noxref_5_c_1626_n N_B_c_1803_n ) capacitor c=3.72011e-19 //x=6.66 \
 //y=2.085 //x2=4.44 //y2=2.085
cc_1439 ( N_noxref_5_c_1646_n N_B_c_1805_n ) capacitor c=0.00395405f //x=9.505 \
 //y=4.07 //x2=10.36 //y2=2.085
cc_1440 ( N_noxref_5_c_1670_n N_B_c_1805_n ) capacitor c=0.00734193f //x=9.505 \
 //y=3.33 //x2=10.36 //y2=2.085
cc_1441 ( N_noxref_5_c_1627_n N_B_c_1805_n ) capacitor c=0.0618066f //x=9.62 \
 //y=3.33 //x2=10.36 //y2=2.085
cc_1442 ( N_noxref_5_c_1656_n N_B_c_1805_n ) capacitor c=0.0248246f //x=9.9 \
 //y=4.58 //x2=10.36 //y2=2.085
cc_1443 ( N_noxref_5_M5_noxref_d N_B_c_1805_n ) capacitor c=0.0173675f \
 //x=9.795 //y=0.91 //x2=10.36 //y2=2.085
cc_1444 ( N_noxref_5_M31_noxref_d N_B_c_1805_n ) capacitor c=0.00915986f \
 //x=9.84 //y=5.02 //x2=10.36 //y2=2.085
cc_1445 ( N_noxref_5_M31_noxref_d N_B_M31_noxref_g ) capacitor c=0.021902f \
 //x=9.84 //y=5.02 //x2=9.765 //y2=6.02
cc_1446 ( N_noxref_5_M31_noxref_d N_B_M32_noxref_g ) capacitor c=0.0212035f \
 //x=9.84 //y=5.02 //x2=10.205 //y2=6.02
cc_1447 ( N_noxref_5_M5_noxref_d N_B_c_1811_n ) capacitor c=0.00216577f \
 //x=9.795 //y=0.91 //x2=9.72 //y2=0.91
cc_1448 ( N_noxref_5_c_1628_n N_B_c_1813_n ) capacitor c=0.00242714f //x=9.905 \
 //y=2.08 //x2=9.72 //y2=1.255
cc_1449 ( N_noxref_5_M5_noxref_d N_B_c_1813_n ) capacitor c=0.00599232f \
 //x=9.795 //y=0.91 //x2=9.72 //y2=1.255
cc_1450 ( N_noxref_5_c_1656_n N_B_c_2011_n ) capacitor c=0.00491319f //x=9.9 \
 //y=4.58 //x2=10.13 //y2=4.79
cc_1451 ( N_noxref_5_M31_noxref_d N_B_c_2011_n ) capacitor c=0.0146105f \
 //x=9.84 //y=5.02 //x2=10.13 //y2=4.79
cc_1452 ( N_noxref_5_c_1657_n N_B_c_1904_n ) capacitor c=0.00491319f //x=9.705 \
 //y=4.58 //x2=9.84 //y2=4.79
cc_1453 ( N_noxref_5_M5_noxref_d N_B_c_1814_n ) capacitor c=0.00220879f \
 //x=9.795 //y=0.91 //x2=10.095 //y2=0.755
cc_1454 ( N_noxref_5_M5_noxref_d N_B_c_2015_n ) capacitor c=0.0138055f \
 //x=9.795 //y=0.91 //x2=10.095 //y2=1.41
cc_1455 ( N_noxref_5_c_1656_n N_B_c_1905_n ) capacitor c=0.00917766f //x=9.9 \
 //y=4.58 //x2=10.205 //y2=4.865
cc_1456 ( N_noxref_5_M31_noxref_d N_B_c_1905_n ) capacitor c=0.00307344f \
 //x=9.84 //y=5.02 //x2=10.205 //y2=4.865
cc_1457 ( N_noxref_5_M5_noxref_d N_B_c_1815_n ) capacitor c=0.00220616f \
 //x=9.795 //y=0.91 //x2=10.25 //y2=0.91
cc_1458 ( N_noxref_5_M5_noxref_d N_B_c_2019_n ) capacitor c=0.00347355f \
 //x=9.795 //y=0.91 //x2=10.25 //y2=1.255
cc_1459 ( N_noxref_5_M5_noxref_d N_B_c_2020_n ) capacitor c=0.007449f \
 //x=9.795 //y=0.91 //x2=10.25 //y2=1.565
cc_1460 ( N_noxref_5_M5_noxref_d N_B_c_1817_n ) capacitor c=0.00829952f \
 //x=9.795 //y=0.91 //x2=10.25 //y2=1.92
cc_1461 ( N_noxref_5_c_1646_n N_B_c_1907_n ) capacitor c=6.08197e-19 //x=9.505 \
 //y=4.07 //x2=6.66 //y2=4.7
cc_1462 ( N_noxref_5_c_1627_n N_B_c_1827_n ) capacitor c=5.85261e-19 //x=9.62 \
 //y=3.33 //x2=10.25 //y2=2.085
cc_1463 ( N_noxref_5_c_1628_n N_B_c_1827_n ) capacitor c=0.0146705f //x=9.905 \
 //y=2.08 //x2=10.25 //y2=2.085
cc_1464 ( N_noxref_5_c_1646_n N_noxref_7_c_2293_n ) capacitor c=0.275255f \
 //x=9.505 //y=4.07 //x2=8.025 //y2=3.7
cc_1465 ( N_noxref_5_c_1670_n N_noxref_7_c_2293_n ) capacitor c=0.109685f \
 //x=9.505 //y=3.33 //x2=8.025 //y2=3.7
cc_1466 ( N_noxref_5_c_1689_n N_noxref_7_c_2293_n ) capacitor c=0.0286715f \
 //x=6.775 //y=3.33 //x2=8.025 //y2=3.7
cc_1467 ( N_noxref_5_c_1626_n N_noxref_7_c_2293_n ) capacitor c=0.00490264f \
 //x=6.66 //y=2.085 //x2=8.025 //y2=3.7
cc_1468 ( N_noxref_5_c_1646_n N_noxref_7_c_2272_n ) capacitor c=0.0293663f \
 //x=9.505 //y=4.07 //x2=4.925 //y2=3.7
cc_1469 ( N_noxref_5_c_1646_n N_noxref_7_c_2182_n ) capacitor c=0.142936f \
 //x=9.505 //y=4.07 //x2=11.725 //y2=3.7
cc_1470 ( N_noxref_5_c_1670_n N_noxref_7_c_2182_n ) capacitor c=0.142037f \
 //x=9.505 //y=3.33 //x2=11.725 //y2=3.7
cc_1471 ( N_noxref_5_c_1627_n N_noxref_7_c_2182_n ) capacitor c=0.0221777f \
 //x=9.62 //y=3.33 //x2=11.725 //y2=3.7
cc_1472 ( N_noxref_5_c_1646_n N_noxref_7_c_2297_n ) capacitor c=0.0267435f \
 //x=9.505 //y=4.07 //x2=8.255 //y2=3.7
cc_1473 ( N_noxref_5_c_1670_n N_noxref_7_c_2297_n ) capacitor c=0.0266741f \
 //x=9.505 //y=3.33 //x2=8.255 //y2=3.7
cc_1474 ( N_noxref_5_c_1627_n N_noxref_7_c_2297_n ) capacitor c=5.90394e-19 \
 //x=9.62 //y=3.33 //x2=8.255 //y2=3.7
cc_1475 ( N_noxref_5_c_1646_n N_noxref_7_c_2230_n ) capacitor c=0.00740361f \
 //x=9.505 //y=4.07 //x2=11.955 //y2=4.07
cc_1476 ( N_noxref_5_c_1646_n N_noxref_7_c_2231_n ) capacitor c=0.00431193f \
 //x=9.505 //y=4.07 //x2=4.725 //y2=5.205
cc_1477 ( N_noxref_5_c_1651_n N_noxref_7_c_2231_n ) capacitor c=0.00102585f \
 //x=4.555 //y=4.07 //x2=4.725 //y2=5.205
cc_1478 ( N_noxref_5_M26_noxref_g N_noxref_7_c_2231_n ) capacitor c=0.0187432f \
 //x=4.55 //y=6.02 //x2=4.725 //y2=5.205
cc_1479 ( N_noxref_5_c_1681_n N_noxref_7_c_2231_n ) capacitor c=0.00161455f \
 //x=4.44 //y=4.7 //x2=4.725 //y2=5.205
cc_1480 ( N_noxref_5_c_1651_n N_noxref_7_c_2233_n ) capacitor c=0.00142608f \
 //x=4.555 //y=4.07 //x2=4.415 //y2=5.205
cc_1481 ( N_noxref_5_c_1652_n N_noxref_7_c_2233_n ) capacitor c=0.0123412f \
 //x=4.44 //y=4.07 //x2=4.415 //y2=5.205
cc_1482 ( N_noxref_5_M25_noxref_g N_noxref_7_c_2233_n ) capacitor c=0.0132788f \
 //x=4.11 //y=6.02 //x2=4.415 //y2=5.205
cc_1483 ( N_noxref_5_c_1681_n N_noxref_7_c_2233_n ) capacitor c=0.00557817f \
 //x=4.44 //y=4.7 //x2=4.415 //y2=5.205
cc_1484 ( N_noxref_5_c_1646_n N_noxref_7_c_2190_n ) capacitor c=0.0229481f \
 //x=9.505 //y=4.07 //x2=4.81 //y2=3.7
cc_1485 ( N_noxref_5_c_1651_n N_noxref_7_c_2190_n ) capacitor c=0.00168517f \
 //x=4.555 //y=4.07 //x2=4.81 //y2=3.7
cc_1486 ( N_noxref_5_c_1689_n N_noxref_7_c_2190_n ) capacitor c=0.00286172f \
 //x=6.775 //y=3.33 //x2=4.81 //y2=3.7
cc_1487 ( N_noxref_5_c_1652_n N_noxref_7_c_2190_n ) capacitor c=0.0637046f \
 //x=4.44 //y=4.07 //x2=4.81 //y2=3.7
cc_1488 ( N_noxref_5_c_1626_n N_noxref_7_c_2190_n ) capacitor c=0.00714689f \
 //x=6.66 //y=2.085 //x2=4.81 //y2=3.7
cc_1489 ( N_noxref_5_c_1681_n N_noxref_7_c_2190_n ) capacitor c=0.0232466f \
 //x=4.44 //y=4.7 //x2=4.81 //y2=3.7
cc_1490 ( N_noxref_5_c_1646_n N_noxref_7_c_2239_n ) capacitor c=0.0181107f \
 //x=9.505 //y=4.07 //x2=8.14 //y2=3.7
cc_1491 ( N_noxref_5_c_1670_n N_noxref_7_c_2239_n ) capacitor c=0.0186917f \
 //x=9.505 //y=3.33 //x2=8.14 //y2=3.7
cc_1492 ( N_noxref_5_c_1626_n N_noxref_7_c_2239_n ) capacitor c=0.00336585f \
 //x=6.66 //y=2.085 //x2=8.14 //y2=3.7
cc_1493 ( N_noxref_5_c_1629_n N_noxref_7_c_2239_n ) capacitor c=0.0147021f \
 //x=9.705 //y=2.08 //x2=8.14 //y2=3.7
cc_1494 ( N_noxref_5_M31_noxref_d N_noxref_7_c_2239_n ) capacitor \
 c=0.00109417f //x=9.84 //y=5.02 //x2=8.14 //y2=3.7
cc_1495 ( N_noxref_5_c_1627_n N_noxref_7_c_2193_n ) capacitor c=9.98852e-19 \
 //x=9.62 //y=3.33 //x2=11.84 //y2=2.085
cc_1496 ( N_noxref_5_M26_noxref_g N_noxref_7_M25_noxref_d ) capacitor \
 c=0.0136385f //x=4.55 //y=6.02 //x2=4.185 //y2=5.02
cc_1497 ( N_noxref_5_M31_noxref_d N_noxref_8_M33_noxref_d ) capacitor \
 c=5.05958e-19 //x=9.84 //y=5.02 //x2=12.07 //y2=5.02
cc_1498 ( N_noxref_5_M25_noxref_g N_noxref_17_c_4059_n ) capacitor \
 c=0.0170604f //x=4.11 //y=6.02 //x2=3.805 //y2=5.205
cc_1499 ( N_noxref_5_M25_noxref_g N_noxref_17_c_4066_n ) capacitor \
 c=0.0150677f //x=4.11 //y=6.02 //x2=4.685 //y2=6.905
cc_1500 ( N_noxref_5_M26_noxref_g N_noxref_17_c_4066_n ) capacitor c=0.016333f \
 //x=4.55 //y=6.02 //x2=4.685 //y2=6.905
cc_1501 ( N_noxref_5_M26_noxref_g N_noxref_17_M26_noxref_d ) capacitor \
 c=0.0351101f //x=4.55 //y=6.02 //x2=4.625 //y2=5.02
cc_1502 ( N_noxref_5_c_1646_n N_noxref_19_c_4154_n ) capacitor c=0.0060417f \
 //x=9.505 //y=4.07 //x2=6.425 //y2=5.205
cc_1503 ( N_noxref_5_c_1636_n N_noxref_20_c_4211_n ) capacitor c=0.0034165f \
 //x=6.465 //y=1.92 //x2=6.245 //y2=1.5
cc_1504 ( N_noxref_5_c_1626_n N_noxref_20_c_4190_n ) capacitor c=0.00911914f \
 //x=6.66 //y=2.085 //x2=7.13 //y2=1.585
cc_1505 ( N_noxref_5_c_1635_n N_noxref_20_c_4190_n ) capacitor c=0.00696002f \
 //x=6.465 //y=1.525 //x2=7.13 //y2=1.585
cc_1506 ( N_noxref_5_c_1636_n N_noxref_20_c_4190_n ) capacitor c=0.0163188f \
 //x=6.465 //y=1.92 //x2=7.13 //y2=1.585
cc_1507 ( N_noxref_5_c_1638_n N_noxref_20_c_4190_n ) capacitor c=0.00772214f \
 //x=6.84 //y=1.37 //x2=7.13 //y2=1.585
cc_1508 ( N_noxref_5_c_1641_n N_noxref_20_c_4190_n ) capacitor c=0.0034036f \
 //x=6.995 //y=1.215 //x2=7.13 //y2=1.585
cc_1509 ( N_noxref_5_c_1636_n N_noxref_20_c_4197_n ) capacitor c=6.71402e-19 \
 //x=6.465 //y=1.92 //x2=7.215 //y2=1.5
cc_1510 ( N_noxref_5_c_1632_n N_noxref_20_M3_noxref_s ) capacitor c=0.0326577f \
 //x=6.465 //y=0.87 //x2=6.11 //y2=0.37
cc_1511 ( N_noxref_5_c_1635_n N_noxref_20_M3_noxref_s ) capacitor \
 c=3.48408e-19 //x=6.465 //y=1.525 //x2=6.11 //y2=0.37
cc_1512 ( N_noxref_5_c_1639_n N_noxref_20_M3_noxref_s ) capacitor c=0.0120759f \
 //x=6.995 //y=0.87 //x2=6.11 //y2=0.37
cc_1513 ( N_B_c_1801_n N_noxref_7_c_2293_n ) capacitor c=0.084255f //x=10.245 \
 //y=2.96 //x2=8.025 //y2=3.7
cc_1514 ( N_B_c_1830_n N_noxref_7_c_2293_n ) capacitor c=0.0102755f //x=10.245 \
 //y=4.44 //x2=8.025 //y2=3.7
cc_1515 ( N_B_c_1837_n N_noxref_7_c_2293_n ) capacitor c=0.00181512f //x=6.775 \
 //y=4.44 //x2=8.025 //y2=3.7
cc_1516 ( N_B_c_1801_n N_noxref_7_c_2272_n ) capacitor c=0.0133597f //x=10.245 \
 //y=2.96 //x2=4.925 //y2=3.7
cc_1517 ( N_B_c_1801_n N_noxref_7_c_2182_n ) capacitor c=0.0432502f //x=10.245 \
 //y=2.96 //x2=11.725 //y2=3.7
cc_1518 ( N_B_c_1830_n N_noxref_7_c_2182_n ) capacitor c=0.0417889f //x=10.245 \
 //y=4.44 //x2=11.725 //y2=3.7
cc_1519 ( N_B_c_1839_n N_noxref_7_c_2182_n ) capacitor c=0.0358408f //x=28.745 \
 //y=4.81 //x2=11.725 //y2=3.7
cc_1520 ( N_B_c_1805_n N_noxref_7_c_2182_n ) capacitor c=0.0243649f //x=10.36 \
 //y=2.085 //x2=11.725 //y2=3.7
cc_1521 ( N_B_c_1801_n N_noxref_7_c_2297_n ) capacitor c=5.76919e-19 \
 //x=10.245 //y=2.96 //x2=8.255 //y2=3.7
cc_1522 ( N_B_c_1830_n N_noxref_7_c_2297_n ) capacitor c=5.69512e-19 \
 //x=10.245 //y=4.44 //x2=8.255 //y2=3.7
cc_1523 ( N_B_c_1839_n N_noxref_7_c_2183_n ) capacitor c=0.0162513f //x=28.745 \
 //y=4.81 //x2=23.935 //y2=2.22
cc_1524 ( N_B_c_1839_n N_noxref_7_c_2188_n ) capacitor c=0.112171f //x=28.745 \
 //y=4.81 //x2=14.315 //y2=4.07
cc_1525 ( N_B_c_1839_n N_noxref_7_c_2230_n ) capacitor c=0.0133159f //x=28.745 \
 //y=4.81 //x2=11.955 //y2=4.07
cc_1526 ( N_B_c_1805_n N_noxref_7_c_2230_n ) capacitor c=0.00131283f //x=10.36 \
 //y=2.085 //x2=11.955 //y2=4.07
cc_1527 ( N_B_c_1939_n N_noxref_7_c_2189_n ) capacitor c=0.00355555f //x=4.105 \
 //y=1.92 //x2=4.725 //y2=1.655
cc_1528 ( N_B_c_1943_n N_noxref_7_c_2189_n ) capacitor c=0.00196666f //x=4.48 \
 //y=1.41 //x2=4.725 //y2=1.655
cc_1529 ( N_B_c_1945_n N_noxref_7_c_2189_n ) capacitor c=0.00423452f //x=4.635 \
 //y=1.255 //x2=4.725 //y2=1.655
cc_1530 ( N_B_c_1803_n N_noxref_7_c_2277_n ) capacitor c=0.0132209f //x=4.44 \
 //y=2.085 //x2=4.455 //y2=1.655
cc_1531 ( N_B_c_1939_n N_noxref_7_c_2277_n ) capacitor c=0.0062602f //x=4.105 \
 //y=1.92 //x2=4.455 //y2=1.655
cc_1532 ( N_B_c_1801_n N_noxref_7_c_2190_n ) capacitor c=0.0192028f //x=10.245 \
 //y=2.96 //x2=4.81 //y2=3.7
cc_1533 ( N_B_c_1910_n N_noxref_7_c_2190_n ) capacitor c=0.00244604f //x=4.555 \
 //y=2.96 //x2=4.81 //y2=3.7
cc_1534 ( B N_noxref_7_c_2190_n ) capacitor c=7.44407e-19 //x=6.66 //y=4.44 \
 //x2=4.81 //y2=3.7
cc_1535 ( N_B_c_1803_n N_noxref_7_c_2190_n ) capacitor c=0.078005f //x=4.44 \
 //y=2.085 //x2=4.81 //y2=3.7
cc_1536 ( N_B_c_1939_n N_noxref_7_c_2190_n ) capacitor c=0.0130045f //x=4.105 \
 //y=1.92 //x2=4.81 //y2=3.7
cc_1537 ( N_B_c_1830_n N_noxref_7_c_2236_n ) capacitor c=0.00665427f \
 //x=10.245 //y=4.44 //x2=8.055 //y2=5.205
cc_1538 ( N_B_c_1830_n N_noxref_7_c_2238_n ) capacitor c=0.00351988f \
 //x=10.245 //y=4.44 //x2=7.745 //y2=5.205
cc_1539 ( N_B_c_1801_n N_noxref_7_c_2239_n ) capacitor c=0.020158f //x=10.245 \
 //y=2.96 //x2=8.14 //y2=3.7
cc_1540 ( N_B_c_1830_n N_noxref_7_c_2239_n ) capacitor c=0.0186407f //x=10.245 \
 //y=4.44 //x2=8.14 //y2=3.7
cc_1541 ( B N_noxref_7_c_2239_n ) capacitor c=0.00138227f //x=6.66 //y=4.44 \
 //x2=8.14 //y2=3.7
cc_1542 ( N_B_c_1805_n N_noxref_7_c_2239_n ) capacitor c=0.00125526f //x=10.36 \
 //y=2.085 //x2=8.14 //y2=3.7
cc_1543 ( N_B_c_1801_n N_noxref_7_c_2193_n ) capacitor c=0.00382596f \
 //x=10.245 //y=2.96 //x2=11.84 //y2=2.085
cc_1544 ( N_B_c_1839_n N_noxref_7_c_2193_n ) capacitor c=0.0142866f //x=28.745 \
 //y=4.81 //x2=11.84 //y2=2.085
cc_1545 ( N_B_c_1805_n N_noxref_7_c_2193_n ) capacitor c=0.0180426f //x=10.36 \
 //y=2.085 //x2=11.84 //y2=2.085
cc_1546 ( N_B_c_1839_n N_noxref_7_c_2198_n ) capacitor c=0.0160683f //x=28.745 \
 //y=4.81 //x2=14.43 //y2=2.085
cc_1547 ( N_B_c_1839_n N_noxref_7_c_2392_n ) capacitor c=0.0189082f //x=28.745 \
 //y=4.81 //x2=24.05 //y2=4.535
cc_1548 ( N_B_c_1839_n N_noxref_7_M33_noxref_g ) capacitor c=0.00545663f \
 //x=28.745 //y=4.81 //x2=11.995 //y2=6.02
cc_1549 ( N_B_c_1839_n N_noxref_7_M34_noxref_g ) capacitor c=0.00561282f \
 //x=28.745 //y=4.81 //x2=12.435 //y2=6.02
cc_1550 ( N_B_c_1839_n N_noxref_7_M35_noxref_g ) capacitor c=0.00288572f \
 //x=28.745 //y=4.81 //x2=14.33 //y2=6.02
cc_1551 ( N_B_c_1839_n N_noxref_7_M36_noxref_g ) capacitor c=0.00278062f \
 //x=28.745 //y=4.81 //x2=14.77 //y2=6.02
cc_1552 ( N_B_c_1839_n N_noxref_7_M47_noxref_g ) capacitor c=0.00255691f \
 //x=28.745 //y=4.81 //x2=24.09 //y2=6.02
cc_1553 ( N_B_c_1839_n N_noxref_7_M48_noxref_g ) capacitor c=0.00308796f \
 //x=28.745 //y=4.81 //x2=24.53 //y2=6.02
cc_1554 ( N_B_c_1839_n N_noxref_7_c_2263_n ) capacitor c=0.00173868f \
 //x=28.745 //y=4.81 //x2=12.36 //y2=4.79
cc_1555 ( N_B_c_1839_n N_noxref_7_c_2264_n ) capacitor c=0.00142457f \
 //x=28.745 //y=4.81 //x2=12.07 //y2=4.79
cc_1556 ( N_B_c_1905_n N_noxref_7_c_2264_n ) capacitor c=2.80896e-19 \
 //x=10.205 //y=4.865 //x2=12.07 //y2=4.79
cc_1557 ( N_B_c_1839_n N_noxref_7_c_2402_n ) capacitor c=0.00706443f \
 //x=28.745 //y=4.81 //x2=24.455 //y2=4.79
cc_1558 ( N_B_c_1827_n N_noxref_7_c_2217_n ) capacitor c=2.82709e-19 //x=10.25 \
 //y=2.085 //x2=11.84 //y2=2.085
cc_1559 ( N_B_c_1839_n N_noxref_7_c_2266_n ) capacitor c=0.00566296f \
 //x=28.745 //y=4.81 //x2=14.43 //y2=4.7
cc_1560 ( N_B_c_1839_n N_noxref_7_c_2405_n ) capacitor c=0.00174211f \
 //x=28.745 //y=4.81 //x2=24.08 //y2=4.7
cc_1561 ( N_B_c_1931_n N_noxref_7_M2_noxref_d ) capacitor c=0.00217566f \
 //x=4.105 //y=0.91 //x2=4.18 //y2=0.91
cc_1562 ( N_B_c_1934_n N_noxref_7_M2_noxref_d ) capacitor c=0.0034598f \
 //x=4.105 //y=1.255 //x2=4.18 //y2=0.91
cc_1563 ( N_B_c_1936_n N_noxref_7_M2_noxref_d ) capacitor c=0.00522042f \
 //x=4.105 //y=1.565 //x2=4.18 //y2=0.91
cc_1564 ( N_B_c_1939_n N_noxref_7_M2_noxref_d ) capacitor c=0.00643086f \
 //x=4.105 //y=1.92 //x2=4.18 //y2=0.91
cc_1565 ( N_B_c_2077_p N_noxref_7_M2_noxref_d ) capacitor c=0.00241053f \
 //x=4.48 //y=0.755 //x2=4.18 //y2=0.91
cc_1566 ( N_B_c_1943_n N_noxref_7_M2_noxref_d ) capacitor c=0.0124466f \
 //x=4.48 //y=1.41 //x2=4.18 //y2=0.91
cc_1567 ( N_B_c_1944_n N_noxref_7_M2_noxref_d ) capacitor c=0.00132245f \
 //x=4.635 //y=0.91 //x2=4.18 //y2=0.91
cc_1568 ( N_B_c_1945_n N_noxref_7_M2_noxref_d ) capacitor c=0.00566463f \
 //x=4.635 //y=1.255 //x2=4.18 //y2=0.91
cc_1569 ( N_B_c_1839_n N_noxref_8_c_2602_n ) capacitor c=0.0137923f //x=28.745 \
 //y=4.81 //x2=18.755 //y2=2.59
cc_1570 ( N_B_c_1839_n N_noxref_8_c_2604_n ) capacitor c=5.08263e-19 \
 //x=28.745 //y=4.81 //x2=12.695 //y2=2.59
cc_1571 ( N_B_c_1839_n N_noxref_8_c_2617_n ) capacitor c=0.0126369f //x=28.745 \
 //y=4.81 //x2=12.495 //y2=4.58
cc_1572 ( N_B_c_1805_n N_noxref_8_c_2607_n ) capacitor c=0.00186982f //x=10.36 \
 //y=2.085 //x2=12.58 //y2=2.59
cc_1573 ( N_B_c_1839_n N_noxref_8_c_2610_n ) capacitor c=0.0114176f //x=28.745 \
 //y=4.81 //x2=18.87 //y2=2.085
cc_1574 ( N_B_c_1839_n N_noxref_8_M41_noxref_g ) capacitor c=0.00521961f \
 //x=28.745 //y=4.81 //x2=18.54 //y2=6.02
cc_1575 ( N_B_c_1839_n N_noxref_8_M42_noxref_g ) capacitor c=0.00288572f \
 //x=28.745 //y=4.81 //x2=18.98 //y2=6.02
cc_1576 ( N_B_c_1839_n N_noxref_8_c_2647_n ) capacitor c=0.00280928f \
 //x=28.745 //y=4.81 //x2=18.87 //y2=4.7
cc_1577 ( N_B_c_1839_n N_noxref_8_M33_noxref_d ) capacitor c=0.0200696f \
 //x=28.745 //y=4.81 //x2=12.07 //y2=5.02
cc_1578 ( N_B_c_1839_n N_SUM_c_2794_n ) capacitor c=0.00688342f //x=28.745 \
 //y=4.81 //x2=19.125 //y2=3.7
cc_1579 ( N_B_c_1839_n N_SUM_c_2795_n ) capacitor c=5.85081e-19 //x=28.745 \
 //y=4.81 //x2=16.025 //y2=3.7
cc_1580 ( N_B_c_1839_n SUM ) capacitor c=0.0202834f //x=28.745 //y=4.81 \
 //x2=15.91 //y2=3.33
cc_1581 ( N_B_c_1839_n SUM ) capacitor c=0.0179428f //x=28.745 //y=4.81 \
 //x2=19.24 //y2=2.59
cc_1582 ( N_B_c_1839_n N_SUM_c_2781_n ) capacitor c=0.018342f //x=28.745 \
 //y=4.81 //x2=15.515 //y2=5.205
cc_1583 ( N_B_c_1839_n N_SUM_c_2784_n ) capacitor c=0.018342f //x=28.745 \
 //y=4.81 //x2=18.845 //y2=5.205
cc_1584 ( N_B_c_1839_n N_noxref_10_c_2933_n ) capacitor c=0.100197f //x=28.745 \
 //y=4.81 //x2=20.605 //y2=4.07
cc_1585 ( N_B_c_1839_n N_noxref_10_c_2955_n ) capacitor c=0.0133733f \
 //x=28.745 //y=4.81 //x2=15.655 //y2=4.07
cc_1586 ( N_B_c_1839_n N_noxref_10_c_2935_n ) capacitor c=0.0140678f \
 //x=28.745 //y=4.81 //x2=15.54 //y2=4.07
cc_1587 ( N_B_c_1839_n N_noxref_10_c_2940_n ) capacitor c=0.0102765f \
 //x=28.745 //y=4.81 //x2=20.805 //y2=4.58
cc_1588 ( N_B_c_1839_n N_noxref_10_M37_noxref_g ) capacitor c=0.00521961f \
 //x=28.745 //y=4.81 //x2=15.21 //y2=6.02
cc_1589 ( N_B_c_1839_n N_noxref_10_M38_noxref_g ) capacitor c=0.00288572f \
 //x=28.745 //y=4.81 //x2=15.65 //y2=6.02
cc_1590 ( N_B_c_1839_n N_noxref_10_c_2960_n ) capacitor c=0.00547599f \
 //x=28.745 //y=4.81 //x2=15.54 //y2=4.7
cc_1591 ( N_B_c_1839_n N_noxref_10_M43_noxref_d ) capacitor c=0.0207947f \
 //x=28.745 //y=4.81 //x2=20.94 //y2=5.02
cc_1592 ( N_B_c_1839_n N_CIN_c_3085_n ) capacitor c=8.03833e-19 //x=28.745 \
 //y=4.81 //x2=21.345 //y2=2.96
cc_1593 ( N_B_c_1839_n N_CIN_c_3115_n ) capacitor c=0.300319f //x=28.745 \
 //y=4.81 //x2=21.345 //y2=4.44
cc_1594 ( N_B_c_1839_n N_CIN_c_3116_n ) capacitor c=0.0300123f //x=28.745 \
 //y=4.81 //x2=17.875 //y2=4.44
cc_1595 ( N_B_c_1839_n N_CIN_c_3087_n ) capacitor c=0.172897f //x=28.745 \
 //y=4.81 //x2=23.195 //y2=4.44
cc_1596 ( N_B_c_1839_n N_CIN_c_3118_n ) capacitor c=0.0272073f //x=28.745 \
 //y=4.81 //x2=21.575 //y2=4.44
cc_1597 ( N_B_c_1839_n CIN ) capacitor c=0.0152342f //x=28.745 //y=4.81 \
 //x2=17.76 //y2=4.44
cc_1598 ( N_B_c_1839_n N_CIN_c_3090_n ) capacitor c=0.0134632f //x=28.745 \
 //y=4.81 //x2=21.46 //y2=2.085
cc_1599 ( N_B_c_1839_n N_CIN_c_3095_n ) capacitor c=0.0162486f //x=28.745 \
 //y=4.81 //x2=23.31 //y2=2.08
cc_1600 ( N_B_c_1839_n N_CIN_M39_noxref_g ) capacitor c=0.00288572f //x=28.745 \
 //y=4.81 //x2=17.66 //y2=6.02
cc_1601 ( N_B_c_1839_n N_CIN_M40_noxref_g ) capacitor c=0.00278062f //x=28.745 \
 //y=4.81 //x2=18.1 //y2=6.02
cc_1602 ( N_B_c_1839_n N_CIN_M43_noxref_g ) capacitor c=0.00561282f //x=28.745 \
 //y=4.81 //x2=20.865 //y2=6.02
cc_1603 ( N_B_c_1839_n N_CIN_M44_noxref_g ) capacitor c=0.00545663f //x=28.745 \
 //y=4.81 //x2=21.305 //y2=6.02
cc_1604 ( N_B_c_1839_n N_CIN_M45_noxref_g ) capacitor c=0.00545663f //x=28.745 \
 //y=4.81 //x2=23.21 //y2=6.02
cc_1605 ( N_B_c_1839_n N_CIN_M46_noxref_g ) capacitor c=0.00276989f //x=28.745 \
 //y=4.81 //x2=23.65 //y2=6.02
cc_1606 ( N_B_c_1839_n N_CIN_c_3140_n ) capacitor c=8.54019e-19 //x=28.745 \
 //y=4.81 //x2=20.94 //y2=4.79
cc_1607 ( N_B_c_1839_n N_CIN_c_3141_n ) capacitor c=0.00124888f //x=28.745 \
 //y=4.81 //x2=21.305 //y2=4.865
cc_1608 ( N_B_c_1839_n N_CIN_c_3143_n ) capacitor c=0.00349942f //x=28.745 \
 //y=4.81 //x2=17.76 //y2=4.7
cc_1609 ( N_B_c_1839_n N_CIN_c_3144_n ) capacitor c=0.00578154f //x=28.745 \
 //y=4.81 //x2=23.31 //y2=4.7
cc_1610 ( N_B_c_1839_n N_noxref_12_c_3336_n ) capacitor c=0.0329704f \
 //x=28.745 //y=4.81 //x2=26.155 //y2=3.33
cc_1611 ( N_B_c_1839_n N_noxref_12_c_3394_n ) capacitor c=0.00523f //x=28.745 \
 //y=4.81 //x2=24.905 //y2=3.33
cc_1612 ( N_B_c_1839_n N_noxref_12_c_3363_n ) capacitor c=0.0569486f \
 //x=28.745 //y=4.81 //x2=23.515 //y2=5.2
cc_1613 ( N_B_c_1839_n N_noxref_12_c_3368_n ) capacitor c=0.0245172f \
 //x=28.745 //y=4.81 //x2=24.79 //y2=3.33
cc_1614 ( N_B_c_1839_n N_noxref_12_c_3339_n ) capacitor c=0.0165049f \
 //x=28.745 //y=4.81 //x2=26.27 //y2=2.085
cc_1615 ( N_B_c_1810_n N_noxref_12_c_3339_n ) capacitor c=0.00121909f \
 //x=28.86 //y=2.08 //x2=26.27 //y2=2.085
cc_1616 ( N_B_c_1839_n N_noxref_12_M49_noxref_g ) capacitor c=0.00545663f \
 //x=28.745 //y=4.81 //x2=26.425 //y2=6.02
cc_1617 ( N_B_c_1839_n N_noxref_12_M50_noxref_g ) capacitor c=0.00561282f \
 //x=28.745 //y=4.81 //x2=26.865 //y2=6.02
cc_1618 ( N_B_c_1839_n N_noxref_12_c_3379_n ) capacitor c=0.00343031f \
 //x=28.745 //y=4.81 //x2=26.79 //y2=4.79
cc_1619 ( N_B_c_1839_n N_noxref_12_c_3380_n ) capacitor c=0.00245815f \
 //x=28.745 //y=4.81 //x2=26.5 //y2=4.79
cc_1620 ( N_B_M52_noxref_g N_noxref_13_c_3502_n ) capacitor c=0.0195934f \
 //x=29.2 //y=6.02 //x2=29.775 //y2=5.2
cc_1621 ( N_B_c_1880_n N_noxref_13_c_3506_n ) capacitor c=0.00158553f \
 //x=28.86 //y=4.63 //x2=29.065 //y2=5.2
cc_1622 ( B N_noxref_13_c_3506_n ) capacitor c=0.0071986f //x=28.86 //y=4.81 \
 //x2=29.065 //y2=5.2
cc_1623 ( N_B_M51_noxref_g N_noxref_13_c_3506_n ) capacitor c=0.0177326f \
 //x=28.76 //y=6.02 //x2=29.065 //y2=5.2
cc_1624 ( N_B_c_1908_n N_noxref_13_c_3506_n ) capacitor c=0.00439828f \
 //x=28.86 //y=4.7 //x2=29.065 //y2=5.2
cc_1625 ( N_B_c_1880_n N_noxref_13_c_3477_n ) capacitor c=2.54914e-19 \
 //x=28.86 //y=4.63 //x2=30.34 //y2=3.33
cc_1626 ( B N_noxref_13_c_3477_n ) capacitor c=8.9408e-19 //x=28.86 //y=4.81 \
 //x2=30.34 //y2=3.33
cc_1627 ( N_B_c_1810_n N_noxref_13_c_3477_n ) capacitor c=0.00359535f \
 //x=28.86 //y=2.08 //x2=30.34 //y2=3.33
cc_1628 ( N_B_M52_noxref_g N_noxref_13_M51_noxref_d ) capacitor c=0.0173476f \
 //x=29.2 //y=6.02 //x2=28.835 //y2=5.02
cc_1629 ( N_B_c_1839_n N_noxref_14_c_3617_n ) capacitor c=0.0285469f \
 //x=28.745 //y=4.81 //x2=34.295 //y2=2.96
cc_1630 ( N_B_c_1880_n N_noxref_14_c_3617_n ) capacitor c=0.00357573f \
 //x=28.86 //y=4.63 //x2=34.295 //y2=2.96
cc_1631 ( B N_noxref_14_c_3617_n ) capacitor c=0.00125414f //x=28.86 //y=4.81 \
 //x2=34.295 //y2=2.96
cc_1632 ( N_B_c_1810_n N_noxref_14_c_3617_n ) capacitor c=0.0276355f //x=28.86 \
 //y=2.08 //x2=34.295 //y2=2.96
cc_1633 ( N_B_c_1821_n N_noxref_14_c_3617_n ) capacitor c=0.00345132f \
 //x=28.665 //y=1.915 //x2=34.295 //y2=2.96
cc_1634 ( N_B_c_1839_n N_noxref_14_c_3675_n ) capacitor c=0.00408345f \
 //x=28.745 //y=4.81 //x2=27.125 //y2=2.96
cc_1635 ( N_B_c_1810_n N_noxref_14_c_3675_n ) capacitor c=7.01366e-19 \
 //x=28.86 //y=2.08 //x2=27.125 //y2=2.96
cc_1636 ( N_B_c_1810_n N_noxref_14_c_3629_n ) capacitor c=0.0161038f //x=28.86 \
 //y=2.08 //x2=26.925 //y2=2.08
cc_1637 ( N_B_c_1839_n N_noxref_14_c_3650_n ) capacitor c=0.0166551f \
 //x=28.745 //y=4.81 //x2=26.925 //y2=4.58
cc_1638 ( B N_noxref_14_c_3650_n ) capacitor c=3.31905e-19 //x=28.86 //y=4.81 \
 //x2=26.925 //y2=4.58
cc_1639 ( N_B_c_1839_n N_noxref_14_M49_noxref_d ) capacitor c=0.0226525f \
 //x=28.745 //y=4.81 //x2=26.5 //y2=5.02
cc_1640 ( N_B_c_1936_n N_noxref_18_c_4106_n ) capacitor c=0.00628626f \
 //x=4.105 //y=1.565 //x2=3.885 //y2=1.5
cc_1641 ( N_B_c_1931_n N_noxref_18_c_4107_n ) capacitor c=0.0197911f //x=4.105 \
 //y=0.91 //x2=4.77 //y2=0.535
cc_1642 ( N_B_c_1944_n N_noxref_18_c_4107_n ) capacitor c=0.00655813f \
 //x=4.635 //y=0.91 //x2=4.77 //y2=0.535
cc_1643 ( N_B_c_1931_n N_noxref_18_M1_noxref_s ) capacitor c=0.00628626f \
 //x=4.105 //y=0.91 //x2=2.78 //y2=0.37
cc_1644 ( N_B_c_1944_n N_noxref_18_M1_noxref_s ) capacitor c=0.0143002f \
 //x=4.635 //y=0.91 //x2=2.78 //y2=0.37
cc_1645 ( N_B_c_1945_n N_noxref_18_M1_noxref_s ) capacitor c=0.00290153f \
 //x=4.635 //y=1.255 //x2=2.78 //y2=0.37
cc_1646 ( N_B_c_1830_n N_noxref_19_c_4149_n ) capacitor c=0.0172642f \
 //x=10.245 //y=4.44 //x2=7.135 //y2=5.205
cc_1647 ( N_B_c_1837_n N_noxref_19_c_4149_n ) capacitor c=0.00485884f \
 //x=6.775 //y=4.44 //x2=7.135 //y2=5.205
cc_1648 ( B N_noxref_19_c_4149_n ) capacitor c=0.0111238f //x=6.66 //y=4.44 \
 //x2=7.135 //y2=5.205
cc_1649 ( N_B_M27_noxref_g N_noxref_19_c_4149_n ) capacitor c=0.018644f \
 //x=6.56 //y=6.02 //x2=7.135 //y2=5.205
cc_1650 ( N_B_M28_noxref_g N_noxref_19_c_4149_n ) capacitor c=0.0169648f //x=7 \
 //y=6.02 //x2=7.135 //y2=5.205
cc_1651 ( N_B_c_1907_n N_noxref_19_c_4149_n ) capacitor c=0.00531676f //x=6.66 \
 //y=4.7 //x2=7.135 //y2=5.205
cc_1652 ( N_B_c_1830_n N_noxref_19_c_4155_n ) capacitor c=0.00389598f \
 //x=10.245 //y=4.44 //x2=8.015 //y2=6.905
cc_1653 ( N_B_M27_noxref_g N_noxref_19_M27_noxref_s ) capacitor c=0.0441361f \
 //x=6.56 //y=6.02 //x2=6.205 //y2=5.02
cc_1654 ( N_B_M28_noxref_g N_noxref_19_M28_noxref_d ) capacitor c=0.0170604f \
 //x=7 //y=6.02 //x2=7.075 //y2=5.02
cc_1655 ( N_B_c_1839_n N_noxref_21_c_4245_n ) capacitor c=0.0445529f \
 //x=28.745 //y=4.81 //x2=14.195 //y2=5.205
cc_1656 ( N_B_c_1839_n N_noxref_21_c_4247_n ) capacitor c=0.00525338f \
 //x=28.745 //y=4.81 //x2=15.785 //y2=6.905
cc_1657 ( N_B_c_1839_n N_noxref_23_c_4331_n ) capacitor c=0.0445529f \
 //x=28.745 //y=4.81 //x2=17.525 //y2=5.205
cc_1658 ( N_B_c_1839_n N_noxref_23_c_4332_n ) capacitor c=0.00535477f \
 //x=28.745 //y=4.81 //x2=19.115 //y2=6.905
cc_1659 ( N_B_c_1821_n N_noxref_26_c_4468_n ) capacitor c=0.0034165f \
 //x=28.665 //y=1.915 //x2=28.445 //y2=1.495
cc_1660 ( B N_noxref_26_c_4469_n ) capacitor c=5.58247e-19 //x=28.86 //y=4.81 \
 //x2=29.33 //y2=1.58
cc_1661 ( N_B_c_1810_n N_noxref_26_c_4469_n ) capacitor c=0.00915291f \
 //x=28.86 //y=2.08 //x2=29.33 //y2=1.58
cc_1662 ( N_B_c_1950_n N_noxref_26_c_4469_n ) capacitor c=0.00695513f \
 //x=28.665 //y=1.52 //x2=29.33 //y2=1.58
cc_1663 ( N_B_c_1821_n N_noxref_26_c_4469_n ) capacitor c=0.01618f //x=28.665 \
 //y=1.915 //x2=29.33 //y2=1.58
cc_1664 ( N_B_c_1823_n N_noxref_26_c_4469_n ) capacitor c=0.00772095f \
 //x=29.04 //y=1.365 //x2=29.33 //y2=1.58
cc_1665 ( N_B_c_1826_n N_noxref_26_c_4469_n ) capacitor c=0.00339872f \
 //x=29.195 //y=1.21 //x2=29.33 //y2=1.58
cc_1666 ( N_B_c_1821_n N_noxref_26_c_4476_n ) capacitor c=6.71402e-19 \
 //x=28.665 //y=1.915 //x2=29.415 //y2=1.495
cc_1667 ( N_B_c_1818_n N_noxref_26_M15_noxref_s ) capacitor c=0.0326577f \
 //x=28.665 //y=0.865 //x2=28.31 //y2=0.365
cc_1668 ( N_B_c_1950_n N_noxref_26_M15_noxref_s ) capacitor c=3.48408e-19 \
 //x=28.665 //y=1.52 //x2=28.31 //y2=0.365
cc_1669 ( N_B_c_1824_n N_noxref_26_M15_noxref_s ) capacitor c=0.0120759f \
 //x=29.195 //y=0.865 //x2=28.31 //y2=0.365
cc_1670 ( N_noxref_7_c_2183_n N_noxref_8_c_2602_n ) capacitor c=0.557732f \
 //x=23.935 //y=2.22 //x2=18.755 //y2=2.59
cc_1671 ( N_noxref_7_c_2188_n N_noxref_8_c_2602_n ) capacitor c=0.0417312f \
 //x=14.315 //y=4.07 //x2=18.755 //y2=2.59
cc_1672 ( N_noxref_7_c_2198_n N_noxref_8_c_2602_n ) capacitor c=0.0237012f \
 //x=14.43 //y=2.085 //x2=18.755 //y2=2.59
cc_1673 ( N_noxref_7_c_2183_n N_noxref_8_c_2604_n ) capacitor c=0.0288578f \
 //x=23.935 //y=2.22 //x2=12.695 //y2=2.59
cc_1674 ( N_noxref_7_c_2188_n N_noxref_8_c_2604_n ) capacitor c=0.00501595f \
 //x=14.315 //y=4.07 //x2=12.695 //y2=2.59
cc_1675 ( N_noxref_7_c_2193_n N_noxref_8_c_2604_n ) capacitor c=0.00735597f \
 //x=11.84 //y=2.085 //x2=12.695 //y2=2.59
cc_1676 ( N_noxref_7_c_2183_n N_noxref_8_c_2605_n ) capacitor c=0.00671665f \
 //x=23.935 //y=2.22 //x2=12.495 //y2=2.08
cc_1677 ( N_noxref_7_c_2198_n N_noxref_8_c_2605_n ) capacitor c=0.01579f \
 //x=14.43 //y=2.085 //x2=12.495 //y2=2.08
cc_1678 ( N_noxref_7_c_2287_n N_noxref_8_c_2605_n ) capacitor c=0.00242714f \
 //x=12.325 //y=1.41 //x2=12.495 //y2=2.08
cc_1679 ( N_noxref_7_c_2183_n N_noxref_8_c_2658_n ) capacitor c=0.00627324f \
 //x=23.935 //y=2.22 //x2=12.295 //y2=2.08
cc_1680 ( N_noxref_7_c_2187_n N_noxref_8_c_2658_n ) capacitor c=9.73374e-19 \
 //x=11.955 //y=2.22 //x2=12.295 //y2=2.08
cc_1681 ( N_noxref_7_c_2217_n N_noxref_8_c_2658_n ) capacitor c=0.014524f \
 //x=11.84 //y=2.085 //x2=12.295 //y2=2.08
cc_1682 ( N_noxref_7_c_2263_n N_noxref_8_c_2617_n ) capacitor c=0.0101013f \
 //x=12.36 //y=4.79 //x2=12.495 //y2=4.58
cc_1683 ( N_noxref_7_c_2188_n N_noxref_8_c_2619_n ) capacitor c=0.00826867f \
 //x=14.315 //y=4.07 //x2=12.3 //y2=4.58
cc_1684 ( N_noxref_7_c_2193_n N_noxref_8_c_2619_n ) capacitor c=0.0237053f \
 //x=11.84 //y=2.085 //x2=12.3 //y2=4.58
cc_1685 ( N_noxref_7_c_2264_n N_noxref_8_c_2619_n ) capacitor c=0.00910651f \
 //x=12.07 //y=4.79 //x2=12.3 //y2=4.58
cc_1686 ( N_noxref_7_c_2182_n N_noxref_8_c_2607_n ) capacitor c=0.00494289f \
 //x=11.725 //y=3.7 //x2=12.58 //y2=2.59
cc_1687 ( N_noxref_7_c_2183_n N_noxref_8_c_2607_n ) capacitor c=0.0125569f \
 //x=23.935 //y=2.22 //x2=12.58 //y2=2.59
cc_1688 ( N_noxref_7_c_2187_n N_noxref_8_c_2607_n ) capacitor c=8.96923e-19 \
 //x=11.955 //y=2.22 //x2=12.58 //y2=2.59
cc_1689 ( N_noxref_7_c_2188_n N_noxref_8_c_2607_n ) capacitor c=0.0246041f \
 //x=14.315 //y=4.07 //x2=12.58 //y2=2.59
cc_1690 ( N_noxref_7_c_2230_n N_noxref_8_c_2607_n ) capacitor c=0.00101501f \
 //x=11.955 //y=4.07 //x2=12.58 //y2=2.59
cc_1691 ( N_noxref_7_c_2193_n N_noxref_8_c_2607_n ) capacitor c=0.063977f \
 //x=11.84 //y=2.085 //x2=12.58 //y2=2.59
cc_1692 ( N_noxref_7_c_2217_n N_noxref_8_c_2607_n ) capacitor c=3.84914e-19 \
 //x=11.84 //y=2.085 //x2=12.58 //y2=2.59
cc_1693 ( N_noxref_7_c_2183_n N_noxref_8_c_2610_n ) capacitor c=0.0151933f \
 //x=23.935 //y=2.22 //x2=18.87 //y2=2.085
cc_1694 ( N_noxref_7_c_2183_n N_noxref_8_c_2636_n ) capacitor c=0.0100622f \
 //x=23.935 //y=2.22 //x2=18.535 //y2=1.92
cc_1695 ( N_noxref_7_c_2193_n N_noxref_8_M6_noxref_d ) capacitor c=0.016954f \
 //x=11.84 //y=2.085 //x2=12.025 //y2=0.91
cc_1696 ( N_noxref_7_c_2201_n N_noxref_8_M6_noxref_d ) capacitor c=0.00218556f \
 //x=11.95 //y=0.91 //x2=12.025 //y2=0.91
cc_1697 ( N_noxref_7_c_2441_p N_noxref_8_M6_noxref_d ) capacitor c=0.00347355f \
 //x=11.95 //y=1.255 //x2=12.025 //y2=0.91
cc_1698 ( N_noxref_7_c_2442_p N_noxref_8_M6_noxref_d ) capacitor c=0.00742431f \
 //x=11.95 //y=1.565 //x2=12.025 //y2=0.91
cc_1699 ( N_noxref_7_c_2203_n N_noxref_8_M6_noxref_d ) capacitor c=0.00829952f \
 //x=11.95 //y=1.92 //x2=12.025 //y2=0.91
cc_1700 ( N_noxref_7_c_2204_n N_noxref_8_M6_noxref_d ) capacitor c=0.00220879f \
 //x=12.325 //y=0.755 //x2=12.025 //y2=0.91
cc_1701 ( N_noxref_7_c_2287_n N_noxref_8_M6_noxref_d ) capacitor c=0.0138055f \
 //x=12.325 //y=1.41 //x2=12.025 //y2=0.91
cc_1702 ( N_noxref_7_c_2205_n N_noxref_8_M6_noxref_d ) capacitor c=0.00218624f \
 //x=12.48 //y=0.91 //x2=12.025 //y2=0.91
cc_1703 ( N_noxref_7_c_2207_n N_noxref_8_M6_noxref_d ) capacitor c=0.00601286f \
 //x=12.48 //y=1.255 //x2=12.025 //y2=0.91
cc_1704 ( N_noxref_7_M33_noxref_g N_noxref_8_M33_noxref_d ) capacitor \
 c=0.0221134f //x=11.995 //y=6.02 //x2=12.07 //y2=5.02
cc_1705 ( N_noxref_7_M34_noxref_g N_noxref_8_M33_noxref_d ) capacitor \
 c=0.0220851f //x=12.435 //y=6.02 //x2=12.07 //y2=5.02
cc_1706 ( N_noxref_7_c_2263_n N_noxref_8_M33_noxref_d ) capacitor c=0.0137349f \
 //x=12.36 //y=4.79 //x2=12.07 //y2=5.02
cc_1707 ( N_noxref_7_c_2264_n N_noxref_8_M33_noxref_d ) capacitor \
 c=0.00307344f //x=12.07 //y=4.79 //x2=12.07 //y2=5.02
cc_1708 ( N_noxref_7_c_2182_n N_SUM_c_2795_n ) capacitor c=0.00359266f \
 //x=11.725 //y=3.7 //x2=16.025 //y2=3.7
cc_1709 ( N_noxref_7_c_2198_n N_SUM_c_2795_n ) capacitor c=0.00251749f \
 //x=14.43 //y=2.085 //x2=16.025 //y2=3.7
cc_1710 ( N_noxref_7_c_2183_n SUM ) capacitor c=0.0143521f //x=23.935 //y=2.22 \
 //x2=15.91 //y2=3.33
cc_1711 ( N_noxref_7_c_2198_n SUM ) capacitor c=0.0143506f //x=14.43 //y=2.085 \
 //x2=15.91 //y2=3.33
cc_1712 ( N_noxref_7_c_2183_n SUM ) capacitor c=0.0166927f //x=23.935 //y=2.22 \
 //x2=19.24 //y2=2.59
cc_1713 ( N_noxref_7_c_2188_n N_noxref_10_c_2955_n ) capacitor c=0.0159617f \
 //x=14.315 //y=4.07 //x2=15.655 //y2=4.07
cc_1714 ( N_noxref_7_c_2198_n N_noxref_10_c_2955_n ) capacitor c=0.00187343f \
 //x=14.43 //y=2.085 //x2=15.655 //y2=4.07
cc_1715 ( N_noxref_7_c_2183_n N_noxref_10_c_2964_n ) capacitor c=0.0088156f \
 //x=23.935 //y=2.22 //x2=20.605 //y2=3.33
cc_1716 ( N_noxref_7_c_2188_n N_noxref_10_c_2935_n ) capacitor c=0.00186775f \
 //x=14.315 //y=4.07 //x2=15.54 //y2=4.07
cc_1717 ( N_noxref_7_c_2198_n N_noxref_10_c_2935_n ) capacitor c=0.0146936f \
 //x=14.43 //y=2.085 //x2=15.54 //y2=4.07
cc_1718 ( N_noxref_7_c_2266_n N_noxref_10_c_2935_n ) capacitor c=0.00206818f \
 //x=14.43 //y=4.7 //x2=15.54 //y2=4.07
cc_1719 ( N_noxref_7_c_2183_n N_noxref_10_c_2913_n ) capacitor c=0.0159854f \
 //x=23.935 //y=2.22 //x2=17.76 //y2=2.085
cc_1720 ( N_noxref_7_c_2198_n N_noxref_10_c_2913_n ) capacitor c=2.12957e-19 \
 //x=14.43 //y=2.085 //x2=17.76 //y2=2.085
cc_1721 ( N_noxref_7_c_2183_n N_noxref_10_c_2914_n ) capacitor c=0.0130629f \
 //x=23.935 //y=2.22 //x2=20.72 //y2=3.33
cc_1722 ( N_noxref_7_c_2183_n N_noxref_10_c_2915_n ) capacitor c=0.0104444f \
 //x=23.935 //y=2.22 //x2=21.005 //y2=2.08
cc_1723 ( N_noxref_7_c_2183_n N_noxref_10_c_2916_n ) capacitor c=0.00212379f \
 //x=23.935 //y=2.22 //x2=20.805 //y2=2.08
cc_1724 ( N_noxref_7_M35_noxref_g N_noxref_10_M37_noxref_g ) capacitor \
 c=0.00995478f //x=14.33 //y=6.02 //x2=15.21 //y2=6.02
cc_1725 ( N_noxref_7_M36_noxref_g N_noxref_10_M37_noxref_g ) capacitor \
 c=0.0607725f //x=14.77 //y=6.02 //x2=15.21 //y2=6.02
cc_1726 ( N_noxref_7_M36_noxref_g N_noxref_10_M38_noxref_g ) capacitor \
 c=0.00934598f //x=14.77 //y=6.02 //x2=15.65 //y2=6.02
cc_1727 ( N_noxref_7_c_2183_n N_noxref_10_c_2923_n ) capacitor c=0.00778021f \
 //x=23.935 //y=2.22 //x2=17.565 //y2=1.92
cc_1728 ( N_noxref_7_c_2198_n N_noxref_10_c_2960_n ) capacitor c=0.00205597f \
 //x=14.43 //y=2.085 //x2=15.54 //y2=4.7
cc_1729 ( N_noxref_7_c_2266_n N_noxref_10_c_2960_n ) capacitor c=0.066508f \
 //x=14.43 //y=4.7 //x2=15.54 //y2=4.7
cc_1730 ( N_noxref_7_c_2183_n N_CIN_c_3085_n ) capacitor c=0.136334f \
 //x=23.935 //y=2.22 //x2=21.345 //y2=2.96
cc_1731 ( N_noxref_7_c_2183_n N_CIN_c_3175_n ) capacitor c=9.72687e-19 \
 //x=23.935 //y=2.22 //x2=15.655 //y2=2.96
cc_1732 ( N_noxref_7_c_2198_n N_CIN_c_3175_n ) capacitor c=0.00526349f \
 //x=14.43 //y=2.085 //x2=15.655 //y2=2.96
cc_1733 ( N_noxref_7_c_2183_n N_CIN_c_3115_n ) capacitor c=5.40549e-19 \
 //x=23.935 //y=2.22 //x2=21.345 //y2=4.44
cc_1734 ( N_noxref_7_c_2183_n N_CIN_c_3087_n ) capacitor c=0.0247047f \
 //x=23.935 //y=2.22 //x2=23.195 //y2=4.44
cc_1735 ( N_noxref_7_c_2199_n N_CIN_c_3087_n ) capacitor c=0.0071153f \
 //x=24.05 //y=2.08 //x2=23.195 //y2=4.44
cc_1736 ( N_noxref_7_c_2183_n N_CIN_c_3088_n ) capacitor c=0.0133561f \
 //x=23.935 //y=2.22 //x2=15.54 //y2=2.085
cc_1737 ( N_noxref_7_c_2198_n N_CIN_c_3088_n ) capacitor c=0.0173966f \
 //x=14.43 //y=2.085 //x2=15.54 //y2=2.085
cc_1738 ( N_noxref_7_c_2211_n N_CIN_c_3088_n ) capacitor c=0.00188281f \
 //x=14.235 //y=1.92 //x2=15.54 //y2=2.085
cc_1739 ( N_noxref_7_c_2183_n N_CIN_c_3090_n ) capacitor c=0.0169229f \
 //x=23.935 //y=2.22 //x2=21.46 //y2=2.085
cc_1740 ( N_noxref_7_c_2199_n N_CIN_c_3090_n ) capacitor c=0.0018227f \
 //x=24.05 //y=2.08 //x2=21.46 //y2=2.085
cc_1741 ( N_noxref_7_c_2183_n N_CIN_c_3095_n ) capacitor c=0.0230807f \
 //x=23.935 //y=2.22 //x2=23.31 //y2=2.08
cc_1742 ( N_noxref_7_c_2392_n N_CIN_c_3095_n ) capacitor c=0.00197351f \
 //x=24.05 //y=4.535 //x2=23.31 //y2=2.08
cc_1743 ( N_noxref_7_c_2199_n N_CIN_c_3095_n ) capacitor c=0.0820691f \
 //x=24.05 //y=2.08 //x2=23.31 //y2=2.08
cc_1744 ( N_noxref_7_c_2291_n N_CIN_c_3095_n ) capacitor c=0.00277771f \
 //x=24.05 //y=2.08 //x2=23.31 //y2=2.08
cc_1745 ( N_noxref_7_c_2405_n N_CIN_c_3095_n ) capacitor c=0.00321326f \
 //x=24.08 //y=4.7 //x2=23.31 //y2=2.08
cc_1746 ( N_noxref_7_M47_noxref_g N_CIN_M45_noxref_g ) capacitor c=0.0103916f \
 //x=24.09 //y=6.02 //x2=23.21 //y2=6.02
cc_1747 ( N_noxref_7_M47_noxref_g N_CIN_M46_noxref_g ) capacitor c=0.106731f \
 //x=24.09 //y=6.02 //x2=23.65 //y2=6.02
cc_1748 ( N_noxref_7_M48_noxref_g N_CIN_M46_noxref_g ) capacitor c=0.00996457f \
 //x=24.53 //y=6.02 //x2=23.65 //y2=6.02
cc_1749 ( N_noxref_7_c_2208_n N_CIN_c_3193_n ) capacitor c=4.86506e-19 \
 //x=14.235 //y=0.87 //x2=15.205 //y2=0.91
cc_1750 ( N_noxref_7_c_2210_n N_CIN_c_3193_n ) capacitor c=0.00152104f \
 //x=14.235 //y=1.215 //x2=15.205 //y2=0.91
cc_1751 ( N_noxref_7_c_2214_n N_CIN_c_3193_n ) capacitor c=0.0157772f \
 //x=14.765 //y=0.87 //x2=15.205 //y2=0.91
cc_1752 ( N_noxref_7_c_2496_p N_CIN_c_3196_n ) capacitor c=0.00109982f \
 //x=14.235 //y=1.525 //x2=15.205 //y2=1.255
cc_1753 ( N_noxref_7_c_2216_n N_CIN_c_3196_n ) capacitor c=0.0117362f \
 //x=14.765 //y=1.215 //x2=15.205 //y2=1.255
cc_1754 ( N_noxref_7_c_2496_p N_CIN_c_3198_n ) capacitor c=9.57794e-19 \
 //x=14.235 //y=1.525 //x2=15.205 //y2=1.565
cc_1755 ( N_noxref_7_c_2211_n N_CIN_c_3198_n ) capacitor c=0.00531182f \
 //x=14.235 //y=1.92 //x2=15.205 //y2=1.565
cc_1756 ( N_noxref_7_c_2216_n N_CIN_c_3198_n ) capacitor c=0.00862358f \
 //x=14.765 //y=1.215 //x2=15.205 //y2=1.565
cc_1757 ( N_noxref_7_c_2183_n N_CIN_c_3150_n ) capacitor c=0.0100622f \
 //x=23.935 //y=2.22 //x2=15.205 //y2=1.92
cc_1758 ( N_noxref_7_c_2198_n N_CIN_c_3150_n ) capacitor c=0.00218978f \
 //x=14.43 //y=2.085 //x2=15.205 //y2=1.92
cc_1759 ( N_noxref_7_c_2211_n N_CIN_c_3150_n ) capacitor c=0.0108001f \
 //x=14.235 //y=1.92 //x2=15.205 //y2=1.92
cc_1760 ( N_noxref_7_c_2214_n N_CIN_c_3204_n ) capacitor c=0.00124821f \
 //x=14.765 //y=0.87 //x2=15.735 //y2=0.91
cc_1761 ( N_noxref_7_c_2216_n N_CIN_c_3205_n ) capacitor c=0.00200715f \
 //x=14.765 //y=1.215 //x2=15.735 //y2=1.255
cc_1762 ( N_noxref_7_c_2506_p N_CIN_c_3103_n ) capacitor c=4.86506e-19 \
 //x=24.085 //y=0.905 //x2=23.115 //y2=0.865
cc_1763 ( N_noxref_7_c_2506_p N_CIN_c_3105_n ) capacitor c=0.00152104f \
 //x=24.085 //y=0.905 //x2=23.115 //y2=1.21
cc_1764 ( N_noxref_7_c_2508_p N_CIN_c_3208_n ) capacitor c=0.00109982f \
 //x=24.085 //y=1.25 //x2=23.115 //y2=1.52
cc_1765 ( N_noxref_7_c_2509_p N_CIN_c_3208_n ) capacitor c=9.57794e-19 \
 //x=24.085 //y=1.56 //x2=23.115 //y2=1.52
cc_1766 ( N_noxref_7_c_2183_n N_CIN_c_3106_n ) capacitor c=0.00667419f \
 //x=23.935 //y=2.22 //x2=23.115 //y2=1.915
cc_1767 ( N_noxref_7_c_2199_n N_CIN_c_3106_n ) capacitor c=0.00276811f \
 //x=24.05 //y=2.08 //x2=23.115 //y2=1.915
cc_1768 ( N_noxref_7_c_2509_p N_CIN_c_3106_n ) capacitor c=0.00535454f \
 //x=24.085 //y=1.56 //x2=23.115 //y2=1.915
cc_1769 ( N_noxref_7_c_2291_n N_CIN_c_3106_n ) capacitor c=0.017087f //x=24.05 \
 //y=2.08 //x2=23.115 //y2=1.915
cc_1770 ( N_noxref_7_c_2506_p N_CIN_c_3109_n ) capacitor c=0.0151475f \
 //x=24.085 //y=0.905 //x2=23.645 //y2=0.865
cc_1771 ( N_noxref_7_c_2515_p N_CIN_c_3109_n ) capacitor c=0.00124821f \
 //x=24.615 //y=0.905 //x2=23.645 //y2=0.865
cc_1772 ( N_noxref_7_c_2508_p N_CIN_c_3111_n ) capacitor c=0.0111064f \
 //x=24.085 //y=1.25 //x2=23.645 //y2=1.21
cc_1773 ( N_noxref_7_c_2509_p N_CIN_c_3111_n ) capacitor c=0.00862358f \
 //x=24.085 //y=1.56 //x2=23.645 //y2=1.21
cc_1774 ( N_noxref_7_c_2518_p N_CIN_c_3111_n ) capacitor c=0.00200715f \
 //x=24.615 //y=1.25 //x2=23.645 //y2=1.21
cc_1775 ( N_noxref_7_c_2183_n N_CIN_c_3112_n ) capacitor c=0.00696407f \
 //x=23.935 //y=2.22 //x2=21.35 //y2=2.085
cc_1776 ( N_noxref_7_c_2392_n N_CIN_c_3144_n ) capacitor c=0.00387682f \
 //x=24.05 //y=4.535 //x2=23.31 //y2=4.7
cc_1777 ( N_noxref_7_c_2405_n N_CIN_c_3144_n ) capacitor c=0.0300377f \
 //x=24.08 //y=4.7 //x2=23.31 //y2=4.7
cc_1778 ( N_noxref_7_c_2199_n N_noxref_12_c_3394_n ) capacitor c=0.00502038f \
 //x=24.05 //y=2.08 //x2=24.905 //y2=3.33
cc_1779 ( N_noxref_7_c_2392_n N_noxref_12_c_3359_n ) capacitor c=0.0101261f \
 //x=24.05 //y=4.535 //x2=24.225 //y2=5.2
cc_1780 ( N_noxref_7_M47_noxref_g N_noxref_12_c_3359_n ) capacitor \
 c=0.0166416f //x=24.09 //y=6.02 //x2=24.225 //y2=5.2
cc_1781 ( N_noxref_7_c_2405_n N_noxref_12_c_3359_n ) capacitor c=0.00326711f \
 //x=24.08 //y=4.7 //x2=24.225 //y2=5.2
cc_1782 ( N_noxref_7_M48_noxref_g N_noxref_12_c_3365_n ) capacitor \
 c=0.0177856f //x=24.53 //y=6.02 //x2=24.705 //y2=5.2
cc_1783 ( N_noxref_7_c_2289_n N_noxref_12_c_3337_n ) capacitor c=0.00371277f \
 //x=24.46 //y=1.405 //x2=24.705 //y2=1.655
cc_1784 ( N_noxref_7_c_2518_p N_noxref_12_c_3337_n ) capacitor c=0.00457401f \
 //x=24.615 //y=1.25 //x2=24.705 //y2=1.655
cc_1785 ( N_noxref_7_c_2183_n N_noxref_12_c_3368_n ) capacitor c=0.00652978f \
 //x=23.935 //y=2.22 //x2=24.79 //y2=3.33
cc_1786 ( N_noxref_7_c_2392_n N_noxref_12_c_3368_n ) capacitor c=0.00831972f \
 //x=24.05 //y=4.535 //x2=24.79 //y2=3.33
cc_1787 ( N_noxref_7_c_2199_n N_noxref_12_c_3368_n ) capacitor c=0.0783284f \
 //x=24.05 //y=2.08 //x2=24.79 //y2=3.33
cc_1788 ( N_noxref_7_c_2402_n N_noxref_12_c_3368_n ) capacitor c=0.0112669f \
 //x=24.455 //y=4.79 //x2=24.79 //y2=3.33
cc_1789 ( N_noxref_7_c_2291_n N_noxref_12_c_3368_n ) capacitor c=0.00700867f \
 //x=24.05 //y=2.08 //x2=24.79 //y2=3.33
cc_1790 ( N_noxref_7_c_2292_n N_noxref_12_c_3368_n ) capacitor c=0.001643f \
 //x=24.05 //y=1.915 //x2=24.79 //y2=3.33
cc_1791 ( N_noxref_7_c_2405_n N_noxref_12_c_3368_n ) capacitor c=0.00517969f \
 //x=24.08 //y=4.7 //x2=24.79 //y2=3.33
cc_1792 ( N_noxref_7_c_2199_n N_noxref_12_c_3339_n ) capacitor c=0.00154446f \
 //x=24.05 //y=2.08 //x2=26.27 //y2=2.085
cc_1793 ( N_noxref_7_c_2402_n N_noxref_12_c_3426_n ) capacitor c=0.00371777f \
 //x=24.455 //y=4.79 //x2=24.31 //y2=5.2
cc_1794 ( N_noxref_7_c_2506_p N_noxref_12_M13_noxref_d ) capacitor \
 c=0.00217566f //x=24.085 //y=0.905 //x2=24.16 //y2=0.905
cc_1795 ( N_noxref_7_c_2508_p N_noxref_12_M13_noxref_d ) capacitor \
 c=0.0034598f //x=24.085 //y=1.25 //x2=24.16 //y2=0.905
cc_1796 ( N_noxref_7_c_2509_p N_noxref_12_M13_noxref_d ) capacitor \
 c=0.00669531f //x=24.085 //y=1.56 //x2=24.16 //y2=0.905
cc_1797 ( N_noxref_7_c_2541_p N_noxref_12_M13_noxref_d ) capacitor \
 c=0.00241102f //x=24.46 //y=0.75 //x2=24.16 //y2=0.905
cc_1798 ( N_noxref_7_c_2289_n N_noxref_12_M13_noxref_d ) capacitor \
 c=0.0137169f //x=24.46 //y=1.405 //x2=24.16 //y2=0.905
cc_1799 ( N_noxref_7_c_2515_p N_noxref_12_M13_noxref_d ) capacitor \
 c=0.00132245f //x=24.615 //y=0.905 //x2=24.16 //y2=0.905
cc_1800 ( N_noxref_7_c_2518_p N_noxref_12_M13_noxref_d ) capacitor \
 c=0.00566463f //x=24.615 //y=1.25 //x2=24.16 //y2=0.905
cc_1801 ( N_noxref_7_c_2292_n N_noxref_12_M13_noxref_d ) capacitor \
 c=0.00660593f //x=24.05 //y=1.915 //x2=24.16 //y2=0.905
cc_1802 ( N_noxref_7_M47_noxref_g N_noxref_12_M47_noxref_d ) capacitor \
 c=0.0173476f //x=24.09 //y=6.02 //x2=24.165 //y2=5.02
cc_1803 ( N_noxref_7_M48_noxref_g N_noxref_12_M47_noxref_d ) capacitor \
 c=0.0179769f //x=24.53 //y=6.02 //x2=24.165 //y2=5.02
cc_1804 ( N_noxref_7_c_2233_n N_noxref_17_c_4059_n ) capacitor c=0.0348754f \
 //x=4.415 //y=5.205 //x2=3.805 //y2=5.205
cc_1805 ( N_noxref_7_c_2231_n N_noxref_17_c_4066_n ) capacitor c=0.0015978f \
 //x=4.725 //y=5.205 //x2=4.685 //y2=6.905
cc_1806 ( N_noxref_7_M25_noxref_d N_noxref_17_c_4066_n ) capacitor c=0.01159f \
 //x=4.185 //y=5.02 //x2=4.685 //y2=6.905
cc_1807 ( N_noxref_7_M25_noxref_d N_noxref_17_M23_noxref_s ) capacitor \
 c=0.00107541f //x=4.185 //y=5.02 //x2=2.875 //y2=5.02
cc_1808 ( N_noxref_7_M25_noxref_d N_noxref_17_M24_noxref_d ) capacitor \
 c=0.0348754f //x=4.185 //y=5.02 //x2=3.745 //y2=5.02
cc_1809 ( N_noxref_7_c_2231_n N_noxref_17_M26_noxref_d ) capacitor \
 c=0.0154556f //x=4.725 //y=5.205 //x2=4.625 //y2=5.02
cc_1810 ( N_noxref_7_M25_noxref_d N_noxref_17_M26_noxref_d ) capacitor \
 c=0.0458293f //x=4.185 //y=5.02 //x2=4.625 //y2=5.02
cc_1811 ( N_noxref_7_c_2277_n N_noxref_18_c_4098_n ) capacitor c=2.94752e-19 \
 //x=4.455 //y=1.655 //x2=2.915 //y2=1.5
cc_1812 ( N_noxref_7_c_2277_n N_noxref_18_c_4106_n ) capacitor c=0.0200666f \
 //x=4.455 //y=1.655 //x2=3.885 //y2=1.5
cc_1813 ( N_noxref_7_c_2189_n N_noxref_18_c_4107_n ) capacitor c=0.00506925f \
 //x=4.725 //y=1.655 //x2=4.77 //y2=0.535
cc_1814 ( N_noxref_7_M2_noxref_d N_noxref_18_c_4107_n ) capacitor c=0.0111538f \
 //x=4.18 //y=0.91 //x2=4.77 //y2=0.535
cc_1815 ( N_noxref_7_c_2189_n N_noxref_18_M1_noxref_s ) capacitor c=0.0138559f \
 //x=4.725 //y=1.655 //x2=2.78 //y2=0.37
cc_1816 ( N_noxref_7_M2_noxref_d N_noxref_18_M1_noxref_s ) capacitor \
 c=0.0436902f //x=4.18 //y=0.91 //x2=2.78 //y2=0.37
cc_1817 ( N_noxref_7_c_2238_n N_noxref_19_c_4149_n ) capacitor c=0.0348754f \
 //x=7.745 //y=5.205 //x2=7.135 //y2=5.205
cc_1818 ( N_noxref_7_c_2231_n N_noxref_19_c_4154_n ) capacitor c=2.91997e-19 \
 //x=4.725 //y=5.205 //x2=6.425 //y2=5.205
cc_1819 ( N_noxref_7_c_2236_n N_noxref_19_c_4155_n ) capacitor c=0.00157156f \
 //x=8.055 //y=5.205 //x2=8.015 //y2=6.905
cc_1820 ( N_noxref_7_M29_noxref_d N_noxref_19_c_4155_n ) capacitor c=0.011538f \
 //x=7.515 //y=5.02 //x2=8.015 //y2=6.905
cc_1821 ( N_noxref_7_M25_noxref_d N_noxref_19_M27_noxref_s ) capacitor \
 c=4.36987e-19 //x=4.185 //y=5.02 //x2=6.205 //y2=5.02
cc_1822 ( N_noxref_7_M29_noxref_d N_noxref_19_M27_noxref_s ) capacitor \
 c=0.00107541f //x=7.515 //y=5.02 //x2=6.205 //y2=5.02
cc_1823 ( N_noxref_7_M29_noxref_d N_noxref_19_M28_noxref_d ) capacitor \
 c=0.0348754f //x=7.515 //y=5.02 //x2=7.075 //y2=5.02
cc_1824 ( N_noxref_7_c_2236_n N_noxref_19_M30_noxref_d ) capacitor \
 c=0.0151538f //x=8.055 //y=5.205 //x2=7.955 //y2=5.02
cc_1825 ( N_noxref_7_M29_noxref_d N_noxref_19_M30_noxref_d ) capacitor \
 c=0.0458293f //x=7.515 //y=5.02 //x2=7.955 //y2=5.02
cc_1826 ( N_noxref_7_c_2189_n N_noxref_20_c_4211_n ) capacitor c=3.32751e-19 \
 //x=4.725 //y=1.655 //x2=6.245 //y2=1.5
cc_1827 ( N_noxref_7_c_2281_n N_noxref_20_c_4211_n ) capacitor c=2.94752e-19 \
 //x=7.785 //y=1.655 //x2=6.245 //y2=1.5
cc_1828 ( N_noxref_7_c_2281_n N_noxref_20_c_4197_n ) capacitor c=0.0202508f \
 //x=7.785 //y=1.655 //x2=7.215 //y2=1.5
cc_1829 ( N_noxref_7_c_2191_n N_noxref_20_c_4198_n ) capacitor c=0.00506925f \
 //x=8.055 //y=1.655 //x2=8.1 //y2=0.535
cc_1830 ( N_noxref_7_M4_noxref_d N_noxref_20_c_4198_n ) capacitor c=0.0111538f \
 //x=7.51 //y=0.91 //x2=8.1 //y2=0.535
cc_1831 ( N_noxref_7_c_2191_n N_noxref_20_M3_noxref_s ) capacitor c=0.0138559f \
 //x=8.055 //y=1.655 //x2=6.11 //y2=0.37
cc_1832 ( N_noxref_7_M4_noxref_d N_noxref_20_M3_noxref_s ) capacitor \
 c=0.0438744f //x=7.51 //y=0.91 //x2=6.11 //y2=0.37
cc_1833 ( N_noxref_7_c_2198_n N_noxref_21_c_4240_n ) capacitor c=0.0092378f \
 //x=14.43 //y=2.085 //x2=14.905 //y2=5.205
cc_1834 ( N_noxref_7_M35_noxref_g N_noxref_21_c_4240_n ) capacitor \
 c=0.0177772f //x=14.33 //y=6.02 //x2=14.905 //y2=5.205
cc_1835 ( N_noxref_7_M36_noxref_g N_noxref_21_c_4240_n ) capacitor c=0.015826f \
 //x=14.77 //y=6.02 //x2=14.905 //y2=5.205
cc_1836 ( N_noxref_7_c_2266_n N_noxref_21_c_4240_n ) capacitor c=0.00486914f \
 //x=14.43 //y=4.7 //x2=14.905 //y2=5.205
cc_1837 ( N_noxref_7_M35_noxref_g N_noxref_21_M35_noxref_s ) capacitor \
 c=0.0441361f //x=14.33 //y=6.02 //x2=13.975 //y2=5.02
cc_1838 ( N_noxref_7_M36_noxref_g N_noxref_21_M36_noxref_d ) capacitor \
 c=0.0170604f //x=14.77 //y=6.02 //x2=14.845 //y2=5.02
cc_1839 ( N_noxref_7_c_2211_n N_noxref_22_c_4277_n ) capacitor c=0.0034165f \
 //x=14.235 //y=1.92 //x2=14.015 //y2=1.5
cc_1840 ( N_noxref_7_c_2198_n N_noxref_22_c_4278_n ) capacitor c=0.00955218f \
 //x=14.43 //y=2.085 //x2=14.9 //y2=1.585
cc_1841 ( N_noxref_7_c_2496_p N_noxref_22_c_4278_n ) capacitor c=0.00696002f \
 //x=14.235 //y=1.525 //x2=14.9 //y2=1.585
cc_1842 ( N_noxref_7_c_2211_n N_noxref_22_c_4278_n ) capacitor c=0.0163188f \
 //x=14.235 //y=1.92 //x2=14.9 //y2=1.585
cc_1843 ( N_noxref_7_c_2213_n N_noxref_22_c_4278_n ) capacitor c=0.00772214f \
 //x=14.61 //y=1.37 //x2=14.9 //y2=1.585
cc_1844 ( N_noxref_7_c_2216_n N_noxref_22_c_4278_n ) capacitor c=0.0034036f \
 //x=14.765 //y=1.215 //x2=14.9 //y2=1.585
cc_1845 ( N_noxref_7_c_2211_n N_noxref_22_c_4285_n ) capacitor c=6.71402e-19 \
 //x=14.235 //y=1.92 //x2=14.985 //y2=1.5
cc_1846 ( N_noxref_7_c_2208_n N_noxref_22_M7_noxref_s ) capacitor c=0.0326577f \
 //x=14.235 //y=0.87 //x2=13.88 //y2=0.37
cc_1847 ( N_noxref_7_c_2496_p N_noxref_22_M7_noxref_s ) capacitor \
 c=3.48408e-19 //x=14.235 //y=1.525 //x2=13.88 //y2=0.37
cc_1848 ( N_noxref_7_c_2214_n N_noxref_22_M7_noxref_s ) capacitor c=0.0120759f \
 //x=14.765 //y=0.87 //x2=13.88 //y2=0.37
cc_1849 ( N_noxref_7_c_2509_p N_noxref_25_c_4423_n ) capacitor c=0.00623646f \
 //x=24.085 //y=1.56 //x2=23.865 //y2=1.495
cc_1850 ( N_noxref_7_c_2291_n N_noxref_25_c_4423_n ) capacitor c=0.00157097f \
 //x=24.05 //y=2.08 //x2=23.865 //y2=1.495
cc_1851 ( N_noxref_7_c_2199_n N_noxref_25_c_4424_n ) capacitor c=9.57163e-19 \
 //x=24.05 //y=2.08 //x2=24.75 //y2=0.53
cc_1852 ( N_noxref_7_c_2506_p N_noxref_25_c_4424_n ) capacitor c=0.0188655f \
 //x=24.085 //y=0.905 //x2=24.75 //y2=0.53
cc_1853 ( N_noxref_7_c_2515_p N_noxref_25_c_4424_n ) capacitor c=0.00656458f \
 //x=24.615 //y=0.905 //x2=24.75 //y2=0.53
cc_1854 ( N_noxref_7_c_2291_n N_noxref_25_c_4424_n ) capacitor c=2.1838e-19 \
 //x=24.05 //y=2.08 //x2=24.75 //y2=0.53
cc_1855 ( N_noxref_7_c_2506_p N_noxref_25_M12_noxref_s ) capacitor \
 c=0.00623646f //x=24.085 //y=0.905 //x2=22.76 //y2=0.365
cc_1856 ( N_noxref_7_c_2515_p N_noxref_25_M12_noxref_s ) capacitor \
 c=0.0143002f //x=24.615 //y=0.905 //x2=22.76 //y2=0.365
cc_1857 ( N_noxref_7_c_2518_p N_noxref_25_M12_noxref_s ) capacitor \
 c=0.00290153f //x=24.615 //y=1.25 //x2=22.76 //y2=0.365
cc_1858 ( N_noxref_8_c_2602_n N_SUM_c_2794_n ) capacitor c=0.00619185f \
 //x=18.755 //y=2.59 //x2=19.125 //y2=3.7
cc_1859 ( N_noxref_8_c_2610_n N_SUM_c_2794_n ) capacitor c=0.0182357f \
 //x=18.87 //y=2.085 //x2=19.125 //y2=3.7
cc_1860 ( N_noxref_8_c_2602_n N_SUM_c_2795_n ) capacitor c=6.30506e-19 \
 //x=18.755 //y=2.59 //x2=16.025 //y2=3.7
cc_1861 ( N_noxref_8_c_2610_n N_SUM_c_2795_n ) capacitor c=2.02744e-19 \
 //x=18.87 //y=2.085 //x2=16.025 //y2=3.7
cc_1862 ( N_noxref_8_c_2602_n SUM ) capacitor c=0.0144f //x=18.755 //y=2.59 \
 //x2=15.91 //y2=3.33
cc_1863 ( N_noxref_8_c_2607_n SUM ) capacitor c=2.79968e-19 //x=12.58 //y=2.59 \
 //x2=15.91 //y2=3.33
cc_1864 ( N_noxref_8_c_2610_n SUM ) capacitor c=0.00277451f //x=18.87 \
 //y=2.085 //x2=15.91 //y2=3.33
cc_1865 ( N_noxref_8_c_2602_n SUM ) capacitor c=0.0100753f //x=18.755 //y=2.59 \
 //x2=19.24 //y2=2.59
cc_1866 ( N_noxref_8_c_2610_n SUM ) capacitor c=0.186203f //x=18.87 //y=2.085 \
 //x2=19.24 //y2=2.59
cc_1867 ( N_noxref_8_c_2636_n SUM ) capacitor c=0.0147734f //x=18.535 //y=1.92 \
 //x2=19.24 //y2=2.59
cc_1868 ( N_noxref_8_c_2647_n SUM ) capacitor c=0.0203f //x=18.87 //y=4.7 \
 //x2=19.24 //y2=2.59
cc_1869 ( N_noxref_8_M42_noxref_g N_SUM_c_2782_n ) capacitor c=0.0173253f \
 //x=18.98 //y=6.02 //x2=19.155 //y2=5.205
cc_1870 ( N_noxref_8_c_2647_n N_SUM_c_2782_n ) capacitor c=0.00161455f \
 //x=18.87 //y=4.7 //x2=19.155 //y2=5.205
cc_1871 ( N_noxref_8_c_2610_n N_SUM_c_2784_n ) capacitor c=0.0100636f \
 //x=18.87 //y=2.085 //x2=18.845 //y2=5.205
cc_1872 ( N_noxref_8_M41_noxref_g N_SUM_c_2784_n ) capacitor c=0.0132788f \
 //x=18.54 //y=6.02 //x2=18.845 //y2=5.205
cc_1873 ( N_noxref_8_c_2647_n N_SUM_c_2784_n ) capacitor c=0.00518581f \
 //x=18.87 //y=4.7 //x2=18.845 //y2=5.205
cc_1874 ( N_noxref_8_c_2636_n N_SUM_c_2766_n ) capacitor c=0.00355555f \
 //x=18.535 //y=1.92 //x2=19.155 //y2=1.655
cc_1875 ( N_noxref_8_c_2637_n N_SUM_c_2766_n ) capacitor c=0.00196666f \
 //x=18.91 //y=1.41 //x2=19.155 //y2=1.655
cc_1876 ( N_noxref_8_c_2705_p N_SUM_c_2766_n ) capacitor c=0.00423452f \
 //x=19.065 //y=1.255 //x2=19.155 //y2=1.655
cc_1877 ( N_noxref_8_c_2610_n N_SUM_c_2793_n ) capacitor c=0.0136356f \
 //x=18.87 //y=2.085 //x2=18.885 //y2=1.655
cc_1878 ( N_noxref_8_c_2636_n N_SUM_c_2793_n ) capacitor c=0.00640467f \
 //x=18.535 //y=1.92 //x2=18.885 //y2=1.655
cc_1879 ( N_noxref_8_c_2708_p N_SUM_M10_noxref_d ) capacitor c=0.00217566f \
 //x=18.535 //y=0.91 //x2=18.61 //y2=0.91
cc_1880 ( N_noxref_8_c_2709_p N_SUM_M10_noxref_d ) capacitor c=0.0034598f \
 //x=18.535 //y=1.255 //x2=18.61 //y2=0.91
cc_1881 ( N_noxref_8_c_2710_p N_SUM_M10_noxref_d ) capacitor c=0.00522042f \
 //x=18.535 //y=1.565 //x2=18.61 //y2=0.91
cc_1882 ( N_noxref_8_c_2636_n N_SUM_M10_noxref_d ) capacitor c=0.00643086f \
 //x=18.535 //y=1.92 //x2=18.61 //y2=0.91
cc_1883 ( N_noxref_8_c_2712_p N_SUM_M10_noxref_d ) capacitor c=0.00241053f \
 //x=18.91 //y=0.755 //x2=18.61 //y2=0.91
cc_1884 ( N_noxref_8_c_2637_n N_SUM_M10_noxref_d ) capacitor c=0.0124466f \
 //x=18.91 //y=1.41 //x2=18.61 //y2=0.91
cc_1885 ( N_noxref_8_c_2714_p N_SUM_M10_noxref_d ) capacitor c=0.00132245f \
 //x=19.065 //y=0.91 //x2=18.61 //y2=0.91
cc_1886 ( N_noxref_8_c_2705_p N_SUM_M10_noxref_d ) capacitor c=0.00566463f \
 //x=19.065 //y=1.255 //x2=18.61 //y2=0.91
cc_1887 ( N_noxref_8_M42_noxref_g N_SUM_M41_noxref_d ) capacitor c=0.0136385f \
 //x=18.98 //y=6.02 //x2=18.615 //y2=5.02
cc_1888 ( N_noxref_8_c_2602_n N_noxref_10_c_2933_n ) capacitor c=7.67045e-19 \
 //x=18.755 //y=2.59 //x2=20.605 //y2=4.07
cc_1889 ( N_noxref_8_c_2610_n N_noxref_10_c_2933_n ) capacitor c=0.0166527f \
 //x=18.87 //y=2.085 //x2=20.605 //y2=4.07
cc_1890 ( N_noxref_8_c_2602_n N_noxref_10_c_2955_n ) capacitor c=6.56372e-19 \
 //x=18.755 //y=2.59 //x2=15.655 //y2=4.07
cc_1891 ( N_noxref_8_c_2602_n N_noxref_10_c_2964_n ) capacitor c=0.00949286f \
 //x=18.755 //y=2.59 //x2=20.605 //y2=3.33
cc_1892 ( N_noxref_8_c_2610_n N_noxref_10_c_2964_n ) capacitor c=0.0158195f \
 //x=18.87 //y=2.085 //x2=20.605 //y2=3.33
cc_1893 ( N_noxref_8_c_2602_n N_noxref_10_c_2984_n ) capacitor c=9.78991e-19 \
 //x=18.755 //y=2.59 //x2=17.875 //y2=3.33
cc_1894 ( N_noxref_8_c_2610_n N_noxref_10_c_2984_n ) capacitor c=7.52994e-19 \
 //x=18.87 //y=2.085 //x2=17.875 //y2=3.33
cc_1895 ( N_noxref_8_c_2602_n N_noxref_10_c_2913_n ) capacitor c=0.0201094f \
 //x=18.755 //y=2.59 //x2=17.76 //y2=2.085
cc_1896 ( N_noxref_8_c_2610_n N_noxref_10_c_2913_n ) capacitor c=0.0217425f \
 //x=18.87 //y=2.085 //x2=17.76 //y2=2.085
cc_1897 ( N_noxref_8_c_2636_n N_noxref_10_c_2913_n ) capacitor c=0.00218978f \
 //x=18.535 //y=1.92 //x2=17.76 //y2=2.085
cc_1898 ( N_noxref_8_c_2610_n N_noxref_10_c_2914_n ) capacitor c=0.00201026f \
 //x=18.87 //y=2.085 //x2=20.72 //y2=3.33
cc_1899 ( N_noxref_8_c_2708_p N_noxref_10_c_2919_n ) capacitor c=4.86506e-19 \
 //x=18.535 //y=0.91 //x2=17.565 //y2=0.87
cc_1900 ( N_noxref_8_c_2708_p N_noxref_10_c_2921_n ) capacitor c=0.00152104f \
 //x=18.535 //y=0.91 //x2=17.565 //y2=1.215
cc_1901 ( N_noxref_8_c_2709_p N_noxref_10_c_2922_n ) capacitor c=0.00109982f \
 //x=18.535 //y=1.255 //x2=17.565 //y2=1.525
cc_1902 ( N_noxref_8_c_2710_p N_noxref_10_c_2922_n ) capacitor c=9.57794e-19 \
 //x=18.535 //y=1.565 //x2=17.565 //y2=1.525
cc_1903 ( N_noxref_8_c_2610_n N_noxref_10_c_2923_n ) capacitor c=0.00188281f \
 //x=18.87 //y=2.085 //x2=17.565 //y2=1.92
cc_1904 ( N_noxref_8_c_2710_p N_noxref_10_c_2923_n ) capacitor c=0.00531182f \
 //x=18.535 //y=1.565 //x2=17.565 //y2=1.92
cc_1905 ( N_noxref_8_c_2636_n N_noxref_10_c_2923_n ) capacitor c=0.0108001f \
 //x=18.535 //y=1.92 //x2=17.565 //y2=1.92
cc_1906 ( N_noxref_8_c_2708_p N_noxref_10_c_2926_n ) capacitor c=0.0157772f \
 //x=18.535 //y=0.91 //x2=18.095 //y2=0.87
cc_1907 ( N_noxref_8_c_2714_p N_noxref_10_c_2926_n ) capacitor c=0.00124821f \
 //x=19.065 //y=0.91 //x2=18.095 //y2=0.87
cc_1908 ( N_noxref_8_c_2709_p N_noxref_10_c_2928_n ) capacitor c=0.0117362f \
 //x=18.535 //y=1.255 //x2=18.095 //y2=1.215
cc_1909 ( N_noxref_8_c_2710_p N_noxref_10_c_2928_n ) capacitor c=0.00862358f \
 //x=18.535 //y=1.565 //x2=18.095 //y2=1.215
cc_1910 ( N_noxref_8_c_2705_p N_noxref_10_c_2928_n ) capacitor c=0.00200715f \
 //x=19.065 //y=1.255 //x2=18.095 //y2=1.215
cc_1911 ( N_noxref_8_c_2602_n N_CIN_c_3085_n ) capacitor c=0.300234f \
 //x=18.755 //y=2.59 //x2=21.345 //y2=2.96
cc_1912 ( N_noxref_8_c_2610_n N_CIN_c_3085_n ) capacitor c=0.0176337f \
 //x=18.87 //y=2.085 //x2=21.345 //y2=2.96
cc_1913 ( N_noxref_8_c_2602_n N_CIN_c_3175_n ) capacitor c=0.0290321f \
 //x=18.755 //y=2.59 //x2=15.655 //y2=2.96
cc_1914 ( N_noxref_8_c_2610_n N_CIN_c_3115_n ) capacitor c=0.0156763f \
 //x=18.87 //y=2.085 //x2=21.345 //y2=4.44
cc_1915 ( N_noxref_8_c_2647_n N_CIN_c_3115_n ) capacitor c=0.00715101f \
 //x=18.87 //y=4.7 //x2=21.345 //y2=4.44
cc_1916 ( N_noxref_8_c_2610_n N_CIN_c_3116_n ) capacitor c=9.41499e-19 \
 //x=18.87 //y=2.085 //x2=17.875 //y2=4.44
cc_1917 ( N_noxref_8_c_2610_n CIN ) capacitor c=0.00631381f //x=18.87 \
 //y=2.085 //x2=17.76 //y2=4.44
cc_1918 ( N_noxref_8_c_2647_n CIN ) capacitor c=0.00204153f //x=18.87 //y=4.7 \
 //x2=17.76 //y2=4.44
cc_1919 ( N_noxref_8_c_2602_n N_CIN_c_3088_n ) capacitor c=0.0175708f \
 //x=18.755 //y=2.59 //x2=15.54 //y2=2.085
cc_1920 ( N_noxref_8_c_2607_n N_CIN_c_3088_n ) capacitor c=2.14844e-19 \
 //x=12.58 //y=2.59 //x2=15.54 //y2=2.085
cc_1921 ( N_noxref_8_M41_noxref_g N_CIN_M39_noxref_g ) capacitor c=0.00995478f \
 //x=18.54 //y=6.02 //x2=17.66 //y2=6.02
cc_1922 ( N_noxref_8_M41_noxref_g N_CIN_M40_noxref_g ) capacitor c=0.0607725f \
 //x=18.54 //y=6.02 //x2=18.1 //y2=6.02
cc_1923 ( N_noxref_8_M42_noxref_g N_CIN_M40_noxref_g ) capacitor c=0.00934598f \
 //x=18.98 //y=6.02 //x2=18.1 //y2=6.02
cc_1924 ( N_noxref_8_c_2610_n N_CIN_c_3143_n ) capacitor c=0.00206818f \
 //x=18.87 //y=2.085 //x2=17.76 //y2=4.7
cc_1925 ( N_noxref_8_c_2647_n N_CIN_c_3143_n ) capacitor c=0.066508f //x=18.87 \
 //y=4.7 //x2=17.76 //y2=4.7
cc_1926 ( N_noxref_8_M41_noxref_g N_noxref_23_c_4326_n ) capacitor \
 c=0.0170604f //x=18.54 //y=6.02 //x2=18.235 //y2=5.205
cc_1927 ( N_noxref_8_M41_noxref_g N_noxref_23_c_4332_n ) capacitor \
 c=0.0141512f //x=18.54 //y=6.02 //x2=19.115 //y2=6.905
cc_1928 ( N_noxref_8_M42_noxref_g N_noxref_23_c_4332_n ) capacitor \
 c=0.0163268f //x=18.98 //y=6.02 //x2=19.115 //y2=6.905
cc_1929 ( N_noxref_8_M42_noxref_g N_noxref_23_M42_noxref_d ) capacitor \
 c=0.0351101f //x=18.98 //y=6.02 //x2=19.055 //y2=5.02
cc_1930 ( N_noxref_8_c_2710_p N_noxref_24_c_4372_n ) capacitor c=0.00628626f \
 //x=18.535 //y=1.565 //x2=18.315 //y2=1.5
cc_1931 ( N_noxref_8_c_2708_p N_noxref_24_c_4373_n ) capacitor c=0.0197911f \
 //x=18.535 //y=0.91 //x2=19.2 //y2=0.535
cc_1932 ( N_noxref_8_c_2714_p N_noxref_24_c_4373_n ) capacitor c=0.00655813f \
 //x=19.065 //y=0.91 //x2=19.2 //y2=0.535
cc_1933 ( N_noxref_8_c_2708_p N_noxref_24_M9_noxref_s ) capacitor \
 c=0.00628626f //x=18.535 //y=0.91 //x2=17.21 //y2=0.37
cc_1934 ( N_noxref_8_c_2714_p N_noxref_24_M9_noxref_s ) capacitor c=0.0143002f \
 //x=19.065 //y=0.91 //x2=17.21 //y2=0.37
cc_1935 ( N_noxref_8_c_2705_p N_noxref_24_M9_noxref_s ) capacitor \
 c=0.00290153f //x=19.065 //y=1.255 //x2=17.21 //y2=0.37
cc_1936 ( N_SUM_c_2794_n N_noxref_10_c_2933_n ) capacitor c=0.304758f \
 //x=19.125 //y=3.7 //x2=20.605 //y2=4.07
cc_1937 ( N_SUM_c_2795_n N_noxref_10_c_2933_n ) capacitor c=0.0293663f \
 //x=16.025 //y=3.7 //x2=20.605 //y2=4.07
cc_1938 ( SUM N_noxref_10_c_2933_n ) capacitor c=0.0202742f //x=15.91 //y=3.33 \
 //x2=20.605 //y2=4.07
cc_1939 ( SUM N_noxref_10_c_2933_n ) capacitor c=0.0181107f //x=19.24 //y=2.59 \
 //x2=20.605 //y2=4.07
cc_1940 ( SUM N_noxref_10_c_2955_n ) capacitor c=0.00168517f //x=15.91 \
 //y=3.33 //x2=15.655 //y2=4.07
cc_1941 ( N_SUM_c_2794_n N_noxref_10_c_2964_n ) capacitor c=0.139118f \
 //x=19.125 //y=3.7 //x2=20.605 //y2=3.33
cc_1942 ( SUM N_noxref_10_c_2964_n ) capacitor c=0.0186917f //x=19.24 //y=2.59 \
 //x2=20.605 //y2=3.33
cc_1943 ( N_SUM_c_2794_n N_noxref_10_c_2984_n ) capacitor c=0.0286715f \
 //x=19.125 //y=3.7 //x2=17.875 //y2=3.33
cc_1944 ( SUM N_noxref_10_c_2984_n ) capacitor c=0.00286172f //x=15.91 \
 //y=3.33 //x2=17.875 //y2=3.33
cc_1945 ( SUM N_noxref_10_c_2935_n ) capacitor c=0.0633004f //x=15.91 //y=3.33 \
 //x2=15.54 //y2=4.07
cc_1946 ( N_SUM_c_2781_n N_noxref_10_c_2935_n ) capacitor c=0.00950688f \
 //x=15.515 //y=5.205 //x2=15.54 //y2=4.07
cc_1947 ( N_SUM_c_2794_n N_noxref_10_c_2913_n ) capacitor c=0.00490264f \
 //x=19.125 //y=3.7 //x2=17.76 //y2=2.085
cc_1948 ( SUM N_noxref_10_c_2913_n ) capacitor c=0.00689401f //x=15.91 \
 //y=3.33 //x2=17.76 //y2=2.085
cc_1949 ( SUM N_noxref_10_c_2913_n ) capacitor c=0.00285275f //x=19.24 \
 //y=2.59 //x2=17.76 //y2=2.085
cc_1950 ( N_SUM_c_2794_n N_noxref_10_c_2914_n ) capacitor c=0.00382062f \
 //x=19.125 //y=3.7 //x2=20.72 //y2=3.33
cc_1951 ( SUM N_noxref_10_c_2916_n ) capacitor c=0.0152631f //x=19.24 //y=2.59 \
 //x2=20.805 //y2=2.08
cc_1952 ( N_SUM_c_2781_n N_noxref_10_M37_noxref_g ) capacitor c=0.0132788f \
 //x=15.515 //y=5.205 //x2=15.21 //y2=6.02
cc_1953 ( N_SUM_c_2779_n N_noxref_10_M38_noxref_g ) capacitor c=0.0173253f \
 //x=15.825 //y=5.205 //x2=15.65 //y2=6.02
cc_1954 ( N_SUM_M37_noxref_d N_noxref_10_M38_noxref_g ) capacitor c=0.0136385f \
 //x=15.285 //y=5.02 //x2=15.65 //y2=6.02
cc_1955 ( SUM N_noxref_10_c_2960_n ) capacitor c=0.0203f //x=15.91 //y=3.33 \
 //x2=15.54 //y2=4.7
cc_1956 ( N_SUM_c_2779_n N_noxref_10_c_2960_n ) capacitor c=0.00161455f \
 //x=15.825 //y=5.205 //x2=15.54 //y2=4.7
cc_1957 ( N_SUM_c_2781_n N_noxref_10_c_2960_n ) capacitor c=0.00518581f \
 //x=15.515 //y=5.205 //x2=15.54 //y2=4.7
cc_1958 ( SUM N_noxref_10_M43_noxref_d ) capacitor c=6.37915e-19 //x=19.24 \
 //y=2.59 //x2=20.94 //y2=5.02
cc_1959 ( N_SUM_c_2794_n N_CIN_c_3085_n ) capacitor c=0.085016f //x=19.125 \
 //y=3.7 //x2=21.345 //y2=2.96
cc_1960 ( N_SUM_c_2795_n N_CIN_c_3085_n ) capacitor c=0.0133597f //x=16.025 \
 //y=3.7 //x2=21.345 //y2=2.96
cc_1961 ( SUM N_CIN_c_3085_n ) capacitor c=0.0192028f //x=15.91 //y=3.33 \
 //x2=21.345 //y2=2.96
cc_1962 ( SUM N_CIN_c_3085_n ) capacitor c=0.0186479f //x=19.24 //y=2.59 \
 //x2=21.345 //y2=2.96
cc_1963 ( SUM N_CIN_c_3175_n ) capacitor c=0.00244604f //x=15.91 //y=3.33 \
 //x2=15.655 //y2=2.96
cc_1964 ( N_SUM_c_2794_n N_CIN_c_3115_n ) capacitor c=0.0110294f //x=19.125 \
 //y=3.7 //x2=21.345 //y2=4.44
cc_1965 ( SUM N_CIN_c_3115_n ) capacitor c=0.014393f //x=19.24 //y=2.59 \
 //x2=21.345 //y2=4.44
cc_1966 ( N_SUM_c_2794_n N_CIN_c_3116_n ) capacitor c=0.00181512f //x=19.125 \
 //y=3.7 //x2=17.875 //y2=4.44
cc_1967 ( SUM CIN ) capacitor c=6.40138e-19 //x=15.91 //y=3.33 //x2=17.76 \
 //y2=4.44
cc_1968 ( SUM CIN ) capacitor c=9.00369e-19 //x=19.24 //y=2.59 //x2=17.76 \
 //y2=4.44
cc_1969 ( SUM N_CIN_c_3088_n ) capacitor c=0.0784004f //x=15.91 //y=3.33 \
 //x2=15.54 //y2=2.085
cc_1970 ( N_SUM_c_2792_n N_CIN_c_3088_n ) capacitor c=0.0132209f //x=15.555 \
 //y=1.655 //x2=15.54 //y2=2.085
cc_1971 ( SUM N_CIN_c_3090_n ) capacitor c=0.0015583f //x=19.24 //y=2.59 \
 //x2=21.46 //y2=2.085
cc_1972 ( N_SUM_M8_noxref_d N_CIN_c_3193_n ) capacitor c=0.00217566f //x=15.28 \
 //y=0.91 //x2=15.205 //y2=0.91
cc_1973 ( N_SUM_M8_noxref_d N_CIN_c_3196_n ) capacitor c=0.0034598f //x=15.28 \
 //y=0.91 //x2=15.205 //y2=1.255
cc_1974 ( N_SUM_M8_noxref_d N_CIN_c_3198_n ) capacitor c=0.00522042f //x=15.28 \
 //y=0.91 //x2=15.205 //y2=1.565
cc_1975 ( SUM N_CIN_c_3150_n ) capacitor c=0.0147734f //x=15.91 //y=3.33 \
 //x2=15.205 //y2=1.92
cc_1976 ( N_SUM_c_2765_n N_CIN_c_3150_n ) capacitor c=0.00355555f //x=15.825 \
 //y=1.655 //x2=15.205 //y2=1.92
cc_1977 ( N_SUM_c_2792_n N_CIN_c_3150_n ) capacitor c=0.00640467f //x=15.555 \
 //y=1.655 //x2=15.205 //y2=1.92
cc_1978 ( N_SUM_M8_noxref_d N_CIN_c_3150_n ) capacitor c=0.00643086f //x=15.28 \
 //y=0.91 //x2=15.205 //y2=1.92
cc_1979 ( N_SUM_M8_noxref_d N_CIN_c_3257_n ) capacitor c=0.00241053f //x=15.28 \
 //y=0.91 //x2=15.58 //y2=0.755
cc_1980 ( N_SUM_c_2765_n N_CIN_c_3151_n ) capacitor c=0.00196666f //x=15.825 \
 //y=1.655 //x2=15.58 //y2=1.41
cc_1981 ( N_SUM_M8_noxref_d N_CIN_c_3151_n ) capacitor c=0.0124466f //x=15.28 \
 //y=0.91 //x2=15.58 //y2=1.41
cc_1982 ( N_SUM_M8_noxref_d N_CIN_c_3204_n ) capacitor c=0.00132245f //x=15.28 \
 //y=0.91 //x2=15.735 //y2=0.91
cc_1983 ( N_SUM_c_2765_n N_CIN_c_3205_n ) capacitor c=0.00423452f //x=15.825 \
 //y=1.655 //x2=15.735 //y2=1.255
cc_1984 ( N_SUM_M8_noxref_d N_CIN_c_3205_n ) capacitor c=0.00566463f //x=15.28 \
 //y=0.91 //x2=15.735 //y2=1.255
cc_1985 ( N_SUM_c_2781_n N_noxref_21_c_4240_n ) capacitor c=0.0348754f \
 //x=15.515 //y=5.205 //x2=14.905 //y2=5.205
cc_1986 ( N_SUM_c_2779_n N_noxref_21_c_4247_n ) capacitor c=0.0015364f \
 //x=15.825 //y=5.205 //x2=15.785 //y2=6.905
cc_1987 ( N_SUM_M37_noxref_d N_noxref_21_c_4247_n ) capacitor c=0.0114841f \
 //x=15.285 //y=5.02 //x2=15.785 //y2=6.905
cc_1988 ( N_SUM_M37_noxref_d N_noxref_21_M35_noxref_s ) capacitor \
 c=0.00107541f //x=15.285 //y=5.02 //x2=13.975 //y2=5.02
cc_1989 ( N_SUM_M37_noxref_d N_noxref_21_M36_noxref_d ) capacitor c=0.0348754f \
 //x=15.285 //y=5.02 //x2=14.845 //y2=5.02
cc_1990 ( N_SUM_c_2779_n N_noxref_21_M38_noxref_d ) capacitor c=0.0147101f \
 //x=15.825 //y=5.205 //x2=15.725 //y2=5.02
cc_1991 ( N_SUM_M37_noxref_d N_noxref_21_M38_noxref_d ) capacitor c=0.0458293f \
 //x=15.285 //y=5.02 //x2=15.725 //y2=5.02
cc_1992 ( N_SUM_c_2792_n N_noxref_22_c_4277_n ) capacitor c=2.94752e-19 \
 //x=15.555 //y=1.655 //x2=14.015 //y2=1.5
cc_1993 ( N_SUM_c_2792_n N_noxref_22_c_4285_n ) capacitor c=0.0200666f \
 //x=15.555 //y=1.655 //x2=14.985 //y2=1.5
cc_1994 ( N_SUM_c_2765_n N_noxref_22_c_4286_n ) capacitor c=0.00506925f \
 //x=15.825 //y=1.655 //x2=15.87 //y2=0.535
cc_1995 ( N_SUM_M8_noxref_d N_noxref_22_c_4286_n ) capacitor c=0.0111538f \
 //x=15.28 //y=0.91 //x2=15.87 //y2=0.535
cc_1996 ( N_SUM_c_2765_n N_noxref_22_M7_noxref_s ) capacitor c=0.0138559f \
 //x=15.825 //y=1.655 //x2=13.88 //y2=0.37
cc_1997 ( N_SUM_M8_noxref_d N_noxref_22_M7_noxref_s ) capacitor c=0.0436902f \
 //x=15.28 //y=0.91 //x2=13.88 //y2=0.37
cc_1998 ( N_SUM_c_2784_n N_noxref_23_c_4326_n ) capacitor c=0.0348754f \
 //x=18.845 //y=5.205 //x2=18.235 //y2=5.205
cc_1999 ( N_SUM_c_2779_n N_noxref_23_c_4331_n ) capacitor c=2.91997e-19 \
 //x=15.825 //y=5.205 //x2=17.525 //y2=5.205
cc_2000 ( N_SUM_c_2782_n N_noxref_23_c_4332_n ) capacitor c=0.0015364f \
 //x=19.155 //y=5.205 //x2=19.115 //y2=6.905
cc_2001 ( N_SUM_M41_noxref_d N_noxref_23_c_4332_n ) capacitor c=0.0114841f \
 //x=18.615 //y=5.02 //x2=19.115 //y2=6.905
cc_2002 ( N_SUM_M37_noxref_d N_noxref_23_M39_noxref_s ) capacitor \
 c=4.36987e-19 //x=15.285 //y=5.02 //x2=17.305 //y2=5.02
cc_2003 ( N_SUM_M41_noxref_d N_noxref_23_M39_noxref_s ) capacitor \
 c=0.00107541f //x=18.615 //y=5.02 //x2=17.305 //y2=5.02
cc_2004 ( N_SUM_M41_noxref_d N_noxref_23_M40_noxref_d ) capacitor c=0.0348754f \
 //x=18.615 //y=5.02 //x2=18.175 //y2=5.02
cc_2005 ( N_SUM_c_2782_n N_noxref_23_M42_noxref_d ) capacitor c=0.0147101f \
 //x=19.155 //y=5.205 //x2=19.055 //y2=5.02
cc_2006 ( N_SUM_M41_noxref_d N_noxref_23_M42_noxref_d ) capacitor c=0.0458293f \
 //x=18.615 //y=5.02 //x2=19.055 //y2=5.02
cc_2007 ( N_SUM_c_2765_n N_noxref_24_c_4386_n ) capacitor c=3.32751e-19 \
 //x=15.825 //y=1.655 //x2=17.345 //y2=1.5
cc_2008 ( N_SUM_c_2793_n N_noxref_24_c_4386_n ) capacitor c=2.94752e-19 \
 //x=18.885 //y=1.655 //x2=17.345 //y2=1.5
cc_2009 ( N_SUM_c_2793_n N_noxref_24_c_4372_n ) capacitor c=0.0202508f \
 //x=18.885 //y=1.655 //x2=18.315 //y2=1.5
cc_2010 ( N_SUM_c_2766_n N_noxref_24_c_4373_n ) capacitor c=0.00506925f \
 //x=19.155 //y=1.655 //x2=19.2 //y2=0.535
cc_2011 ( N_SUM_M10_noxref_d N_noxref_24_c_4373_n ) capacitor c=0.0111538f \
 //x=18.61 //y=0.91 //x2=19.2 //y2=0.535
cc_2012 ( N_SUM_c_2766_n N_noxref_24_M9_noxref_s ) capacitor c=0.0138559f \
 //x=19.155 //y=1.655 //x2=17.21 //y2=0.37
cc_2013 ( N_SUM_M10_noxref_d N_noxref_24_M9_noxref_s ) capacitor c=0.0438744f \
 //x=18.61 //y=0.91 //x2=17.21 //y2=0.37
cc_2014 ( N_noxref_10_c_2933_n N_CIN_c_3085_n ) capacitor c=0.0166896f \
 //x=20.605 //y=4.07 //x2=21.345 //y2=2.96
cc_2015 ( N_noxref_10_c_2964_n N_CIN_c_3085_n ) capacitor c=0.269397f \
 //x=20.605 //y=3.33 //x2=21.345 //y2=2.96
cc_2016 ( N_noxref_10_c_2984_n N_CIN_c_3085_n ) capacitor c=0.0291219f \
 //x=17.875 //y=3.33 //x2=21.345 //y2=2.96
cc_2017 ( N_noxref_10_c_2913_n N_CIN_c_3085_n ) capacitor c=0.0215791f \
 //x=17.76 //y=2.085 //x2=21.345 //y2=2.96
cc_2018 ( N_noxref_10_c_2914_n N_CIN_c_3085_n ) capacitor c=0.0244663f \
 //x=20.72 //y=3.33 //x2=21.345 //y2=2.96
cc_2019 ( N_noxref_10_c_2955_n N_CIN_c_3175_n ) capacitor c=0.00956028f \
 //x=15.655 //y=4.07 //x2=15.655 //y2=2.96
cc_2020 ( N_noxref_10_c_2935_n N_CIN_c_3175_n ) capacitor c=2.06418e-19 \
 //x=15.54 //y=4.07 //x2=15.655 //y2=2.96
cc_2021 ( N_noxref_10_c_2933_n N_CIN_c_3115_n ) capacitor c=0.267726f \
 //x=20.605 //y=4.07 //x2=21.345 //y2=4.44
cc_2022 ( N_noxref_10_c_2964_n N_CIN_c_3115_n ) capacitor c=0.00450734f \
 //x=20.605 //y=3.33 //x2=21.345 //y2=4.44
cc_2023 ( N_noxref_10_c_2914_n N_CIN_c_3115_n ) capacitor c=0.0125568f \
 //x=20.72 //y=3.33 //x2=21.345 //y2=4.44
cc_2024 ( N_noxref_10_c_2939_n N_CIN_c_3115_n ) capacitor c=0.0107052f //x=21 \
 //y=4.58 //x2=21.345 //y2=4.44
cc_2025 ( N_noxref_10_c_2940_n N_CIN_c_3115_n ) capacitor c=0.00279065f \
 //x=20.805 //y=4.58 //x2=21.345 //y2=4.44
cc_2026 ( N_noxref_10_c_2933_n N_CIN_c_3116_n ) capacitor c=0.0286083f \
 //x=20.605 //y=4.07 //x2=17.875 //y2=4.44
cc_2027 ( N_noxref_10_c_2914_n N_CIN_c_3118_n ) capacitor c=5.73829e-19 \
 //x=20.72 //y=3.33 //x2=21.575 //y2=4.44
cc_2028 ( N_noxref_10_c_2939_n N_CIN_c_3118_n ) capacitor c=8.69443e-19 //x=21 \
 //y=4.58 //x2=21.575 //y2=4.44
cc_2029 ( N_noxref_10_c_2933_n CIN ) capacitor c=0.00480464f //x=20.605 \
 //y=4.07 //x2=17.76 //y2=4.44
cc_2030 ( N_noxref_10_c_2913_n CIN ) capacitor c=0.00883142f //x=17.76 \
 //y=2.085 //x2=17.76 //y2=4.44
cc_2031 ( N_noxref_10_c_2955_n N_CIN_c_3088_n ) capacitor c=2.06418e-19 \
 //x=15.655 //y=4.07 //x2=15.54 //y2=2.085
cc_2032 ( N_noxref_10_c_2935_n N_CIN_c_3088_n ) capacitor c=0.00912271f \
 //x=15.54 //y=4.07 //x2=15.54 //y2=2.085
cc_2033 ( N_noxref_10_c_2913_n N_CIN_c_3088_n ) capacitor c=3.72011e-19 \
 //x=17.76 //y=2.085 //x2=15.54 //y2=2.085
cc_2034 ( N_noxref_10_c_2933_n N_CIN_c_3090_n ) capacitor c=0.00735597f \
 //x=20.605 //y=4.07 //x2=21.46 //y2=2.085
cc_2035 ( N_noxref_10_c_2964_n N_CIN_c_3090_n ) capacitor c=0.00493066f \
 //x=20.605 //y=3.33 //x2=21.46 //y2=2.085
cc_2036 ( N_noxref_10_c_2914_n N_CIN_c_3090_n ) capacitor c=0.0625765f \
 //x=20.72 //y=3.33 //x2=21.46 //y2=2.085
cc_2037 ( N_noxref_10_c_2939_n N_CIN_c_3090_n ) capacitor c=0.025409f //x=21 \
 //y=4.58 //x2=21.46 //y2=2.085
cc_2038 ( N_noxref_10_M11_noxref_d N_CIN_c_3090_n ) capacitor c=0.0173592f \
 //x=20.895 //y=0.91 //x2=21.46 //y2=2.085
cc_2039 ( N_noxref_10_c_2914_n N_CIN_c_3095_n ) capacitor c=0.00103525f \
 //x=20.72 //y=3.33 //x2=23.31 //y2=2.08
cc_2040 ( N_noxref_10_M43_noxref_d N_CIN_M43_noxref_g ) capacitor c=0.0220851f \
 //x=20.94 //y=5.02 //x2=20.865 //y2=6.02
cc_2041 ( N_noxref_10_M43_noxref_d N_CIN_M44_noxref_g ) capacitor c=0.0221134f \
 //x=20.94 //y=5.02 //x2=21.305 //y2=6.02
cc_2042 ( N_noxref_10_M11_noxref_d N_CIN_c_3096_n ) capacitor c=0.00216577f \
 //x=20.895 //y=0.91 //x2=20.82 //y2=0.91
cc_2043 ( N_noxref_10_c_2915_n N_CIN_c_3098_n ) capacitor c=0.00242714f \
 //x=21.005 //y=2.08 //x2=20.82 //y2=1.255
cc_2044 ( N_noxref_10_M11_noxref_d N_CIN_c_3098_n ) capacitor c=0.00599232f \
 //x=20.895 //y=0.91 //x2=20.82 //y2=1.255
cc_2045 ( N_noxref_10_c_2939_n N_CIN_c_3294_n ) capacitor c=0.00505067f //x=21 \
 //y=4.58 //x2=21.23 //y2=4.79
cc_2046 ( N_noxref_10_M43_noxref_d N_CIN_c_3294_n ) capacitor c=0.0137349f \
 //x=20.94 //y=5.02 //x2=21.23 //y2=4.79
cc_2047 ( N_noxref_10_c_2940_n N_CIN_c_3140_n ) capacitor c=0.00505067f \
 //x=20.805 //y=4.58 //x2=20.94 //y2=4.79
cc_2048 ( N_noxref_10_M11_noxref_d N_CIN_c_3099_n ) capacitor c=0.00220879f \
 //x=20.895 //y=0.91 //x2=21.195 //y2=0.755
cc_2049 ( N_noxref_10_M11_noxref_d N_CIN_c_3298_n ) capacitor c=0.0138055f \
 //x=20.895 //y=0.91 //x2=21.195 //y2=1.41
cc_2050 ( N_noxref_10_c_2939_n N_CIN_c_3141_n ) capacitor c=0.00941483f //x=21 \
 //y=4.58 //x2=21.305 //y2=4.865
cc_2051 ( N_noxref_10_M43_noxref_d N_CIN_c_3141_n ) capacitor c=0.00307344f \
 //x=20.94 //y=5.02 //x2=21.305 //y2=4.865
cc_2052 ( N_noxref_10_M11_noxref_d N_CIN_c_3100_n ) capacitor c=0.00220616f \
 //x=20.895 //y=0.91 //x2=21.35 //y2=0.91
cc_2053 ( N_noxref_10_M11_noxref_d N_CIN_c_3302_n ) capacitor c=0.00347355f \
 //x=20.895 //y=0.91 //x2=21.35 //y2=1.255
cc_2054 ( N_noxref_10_M11_noxref_d N_CIN_c_3303_n ) capacitor c=0.007449f \
 //x=20.895 //y=0.91 //x2=21.35 //y2=1.565
cc_2055 ( N_noxref_10_M11_noxref_d N_CIN_c_3102_n ) capacitor c=0.00829952f \
 //x=20.895 //y=0.91 //x2=21.35 //y2=1.92
cc_2056 ( N_noxref_10_c_2933_n N_CIN_c_3143_n ) capacitor c=4.45507e-19 \
 //x=20.605 //y=4.07 //x2=17.76 //y2=4.7
cc_2057 ( N_noxref_10_c_2914_n N_CIN_c_3112_n ) capacitor c=3.84914e-19 \
 //x=20.72 //y=3.33 //x2=21.35 //y2=2.085
cc_2058 ( N_noxref_10_c_2915_n N_CIN_c_3112_n ) capacitor c=0.014524f \
 //x=21.005 //y=2.08 //x2=21.35 //y2=2.085
cc_2059 ( N_noxref_10_c_2964_n N_noxref_12_c_3394_n ) capacitor c=0.00359266f \
 //x=20.605 //y=3.33 //x2=24.905 //y2=3.33
cc_2060 ( N_noxref_10_M37_noxref_g N_noxref_21_c_4240_n ) capacitor \
 c=0.0170604f //x=15.21 //y=6.02 //x2=14.905 //y2=5.205
cc_2061 ( N_noxref_10_M37_noxref_g N_noxref_21_c_4247_n ) capacitor \
 c=0.0141512f //x=15.21 //y=6.02 //x2=15.785 //y2=6.905
cc_2062 ( N_noxref_10_M38_noxref_g N_noxref_21_c_4247_n ) capacitor \
 c=0.0163268f //x=15.65 //y=6.02 //x2=15.785 //y2=6.905
cc_2063 ( N_noxref_10_M38_noxref_g N_noxref_21_M38_noxref_d ) capacitor \
 c=0.0351101f //x=15.65 //y=6.02 //x2=15.725 //y2=5.02
cc_2064 ( N_noxref_10_c_2923_n N_noxref_24_c_4386_n ) capacitor c=0.0034165f \
 //x=17.565 //y=1.92 //x2=17.345 //y2=1.5
cc_2065 ( N_noxref_10_c_2913_n N_noxref_24_c_4365_n ) capacitor c=0.00911914f \
 //x=17.76 //y=2.085 //x2=18.23 //y2=1.585
cc_2066 ( N_noxref_10_c_2922_n N_noxref_24_c_4365_n ) capacitor c=0.00696002f \
 //x=17.565 //y=1.525 //x2=18.23 //y2=1.585
cc_2067 ( N_noxref_10_c_2923_n N_noxref_24_c_4365_n ) capacitor c=0.0163188f \
 //x=17.565 //y=1.92 //x2=18.23 //y2=1.585
cc_2068 ( N_noxref_10_c_2925_n N_noxref_24_c_4365_n ) capacitor c=0.00772214f \
 //x=17.94 //y=1.37 //x2=18.23 //y2=1.585
cc_2069 ( N_noxref_10_c_2928_n N_noxref_24_c_4365_n ) capacitor c=0.0034036f \
 //x=18.095 //y=1.215 //x2=18.23 //y2=1.585
cc_2070 ( N_noxref_10_c_2923_n N_noxref_24_c_4372_n ) capacitor c=6.71402e-19 \
 //x=17.565 //y=1.92 //x2=18.315 //y2=1.5
cc_2071 ( N_noxref_10_c_2919_n N_noxref_24_M9_noxref_s ) capacitor \
 c=0.0326577f //x=17.565 //y=0.87 //x2=17.21 //y2=0.37
cc_2072 ( N_noxref_10_c_2922_n N_noxref_24_M9_noxref_s ) capacitor \
 c=3.48408e-19 //x=17.565 //y=1.525 //x2=17.21 //y2=0.37
cc_2073 ( N_noxref_10_c_2926_n N_noxref_24_M9_noxref_s ) capacitor \
 c=0.0120759f //x=18.095 //y=0.87 //x2=17.21 //y2=0.37
cc_2074 ( N_CIN_M46_noxref_g N_noxref_12_c_3359_n ) capacitor c=0.0158157f \
 //x=23.65 //y=6.02 //x2=24.225 //y2=5.2
cc_2075 ( N_CIN_c_3095_n N_noxref_12_c_3363_n ) capacitor c=0.00367046f \
 //x=23.31 //y=2.08 //x2=23.515 //y2=5.2
cc_2076 ( N_CIN_M45_noxref_g N_noxref_12_c_3363_n ) capacitor c=0.0177326f \
 //x=23.21 //y=6.02 //x2=23.515 //y2=5.2
cc_2077 ( N_CIN_c_3144_n N_noxref_12_c_3363_n ) capacitor c=0.00542152f \
 //x=23.31 //y=4.7 //x2=23.515 //y2=5.2
cc_2078 ( N_CIN_c_3095_n N_noxref_12_c_3368_n ) capacitor c=0.00422717f \
 //x=23.31 //y=2.08 //x2=24.79 //y2=3.33
cc_2079 ( N_CIN_M46_noxref_g N_noxref_12_M45_noxref_d ) capacitor c=0.0173476f \
 //x=23.65 //y=6.02 //x2=23.285 //y2=5.02
cc_2080 ( N_CIN_c_3198_n N_noxref_22_c_4285_n ) capacitor c=0.00628626f \
 //x=15.205 //y=1.565 //x2=14.985 //y2=1.5
cc_2081 ( N_CIN_c_3193_n N_noxref_22_c_4286_n ) capacitor c=0.0197911f \
 //x=15.205 //y=0.91 //x2=15.87 //y2=0.535
cc_2082 ( N_CIN_c_3204_n N_noxref_22_c_4286_n ) capacitor c=0.00655813f \
 //x=15.735 //y=0.91 //x2=15.87 //y2=0.535
cc_2083 ( N_CIN_c_3193_n N_noxref_22_M7_noxref_s ) capacitor c=0.00628626f \
 //x=15.205 //y=0.91 //x2=13.88 //y2=0.37
cc_2084 ( N_CIN_c_3204_n N_noxref_22_M7_noxref_s ) capacitor c=0.0143002f \
 //x=15.735 //y=0.91 //x2=13.88 //y2=0.37
cc_2085 ( N_CIN_c_3205_n N_noxref_22_M7_noxref_s ) capacitor c=0.00290153f \
 //x=15.735 //y=1.255 //x2=13.88 //y2=0.37
cc_2086 ( CIN N_noxref_23_c_4326_n ) capacitor c=0.00910154f //x=17.76 \
 //y=4.44 //x2=18.235 //y2=5.205
cc_2087 ( N_CIN_M39_noxref_g N_noxref_23_c_4326_n ) capacitor c=0.0177772f \
 //x=17.66 //y=6.02 //x2=18.235 //y2=5.205
cc_2088 ( N_CIN_M40_noxref_g N_noxref_23_c_4326_n ) capacitor c=0.015826f \
 //x=18.1 //y=6.02 //x2=18.235 //y2=5.205
cc_2089 ( N_CIN_c_3143_n N_noxref_23_c_4326_n ) capacitor c=0.00486914f \
 //x=17.76 //y=4.7 //x2=18.235 //y2=5.205
cc_2090 ( N_CIN_M39_noxref_g N_noxref_23_M39_noxref_s ) capacitor c=0.0441361f \
 //x=17.66 //y=6.02 //x2=17.305 //y2=5.02
cc_2091 ( N_CIN_M40_noxref_g N_noxref_23_M40_noxref_d ) capacitor c=0.0170604f \
 //x=18.1 //y=6.02 //x2=18.175 //y2=5.02
cc_2092 ( N_CIN_c_3106_n N_noxref_25_c_4415_n ) capacitor c=0.0034165f \
 //x=23.115 //y=1.915 //x2=22.895 //y2=1.495
cc_2093 ( N_CIN_c_3095_n N_noxref_25_c_4416_n ) capacitor c=0.00915253f \
 //x=23.31 //y=2.08 //x2=23.78 //y2=1.58
cc_2094 ( N_CIN_c_3208_n N_noxref_25_c_4416_n ) capacitor c=0.00695513f \
 //x=23.115 //y=1.52 //x2=23.78 //y2=1.58
cc_2095 ( N_CIN_c_3106_n N_noxref_25_c_4416_n ) capacitor c=0.0163257f \
 //x=23.115 //y=1.915 //x2=23.78 //y2=1.58
cc_2096 ( N_CIN_c_3108_n N_noxref_25_c_4416_n ) capacitor c=0.00772095f \
 //x=23.49 //y=1.365 //x2=23.78 //y2=1.58
cc_2097 ( N_CIN_c_3111_n N_noxref_25_c_4416_n ) capacitor c=0.00339872f \
 //x=23.645 //y=1.21 //x2=23.78 //y2=1.58
cc_2098 ( N_CIN_c_3106_n N_noxref_25_c_4423_n ) capacitor c=6.71402e-19 \
 //x=23.115 //y=1.915 //x2=23.865 //y2=1.495
cc_2099 ( N_CIN_c_3103_n N_noxref_25_M12_noxref_s ) capacitor c=0.0326577f \
 //x=23.115 //y=0.865 //x2=22.76 //y2=0.365
cc_2100 ( N_CIN_c_3208_n N_noxref_25_M12_noxref_s ) capacitor c=3.48408e-19 \
 //x=23.115 //y=1.52 //x2=22.76 //y2=0.365
cc_2101 ( N_CIN_c_3109_n N_noxref_25_M12_noxref_s ) capacitor c=0.0120759f \
 //x=23.645 //y=0.865 //x2=22.76 //y2=0.365
cc_2102 ( N_noxref_12_c_3336_n N_noxref_13_c_3500_n ) capacitor c=0.00359266f \
 //x=26.155 //y=3.33 //x2=30.455 //y2=3.33
cc_2103 ( N_noxref_12_c_3339_n N_noxref_14_c_3675_n ) capacitor c=0.00735597f \
 //x=26.27 //y=2.085 //x2=27.125 //y2=2.96
cc_2104 ( N_noxref_12_c_3399_n N_noxref_14_c_3629_n ) capacitor c=0.00242714f \
 //x=26.755 //y=1.41 //x2=26.925 //y2=2.08
cc_2105 ( N_noxref_12_c_3351_n N_noxref_14_c_3693_n ) capacitor c=0.0131993f \
 //x=26.27 //y=2.085 //x2=26.725 //y2=2.08
cc_2106 ( N_noxref_12_c_3379_n N_noxref_14_c_3650_n ) capacitor c=0.00988771f \
 //x=26.79 //y=4.79 //x2=26.925 //y2=4.58
cc_2107 ( N_noxref_12_c_3339_n N_noxref_14_c_3652_n ) capacitor c=0.023923f \
 //x=26.27 //y=2.085 //x2=26.73 //y2=4.58
cc_2108 ( N_noxref_12_c_3380_n N_noxref_14_c_3652_n ) capacitor c=0.00723812f \
 //x=26.5 //y=4.79 //x2=26.73 //y2=4.58
cc_2109 ( N_noxref_12_c_3336_n N_noxref_14_c_3631_n ) capacitor c=0.00502038f \
 //x=26.155 //y=3.33 //x2=27.01 //y2=2.96
cc_2110 ( N_noxref_12_c_3368_n N_noxref_14_c_3631_n ) capacitor c=0.0012766f \
 //x=24.79 //y=3.33 //x2=27.01 //y2=2.96
cc_2111 ( N_noxref_12_c_3339_n N_noxref_14_c_3631_n ) capacitor c=0.0682571f \
 //x=26.27 //y=2.085 //x2=27.01 //y2=2.96
cc_2112 ( N_noxref_12_c_3351_n N_noxref_14_c_3631_n ) capacitor c=5.85261e-19 \
 //x=26.27 //y=2.085 //x2=27.01 //y2=2.96
cc_2113 ( N_noxref_12_c_3339_n N_noxref_14_M14_noxref_d ) capacitor \
 c=0.0176945f //x=26.27 //y=2.085 //x2=26.455 //y2=0.91
cc_2114 ( N_noxref_12_c_3344_n N_noxref_14_M14_noxref_d ) capacitor \
 c=0.00218556f //x=26.38 //y=0.91 //x2=26.455 //y2=0.91
cc_2115 ( N_noxref_12_c_3457_p N_noxref_14_M14_noxref_d ) capacitor \
 c=0.00347355f //x=26.38 //y=1.255 //x2=26.455 //y2=0.91
cc_2116 ( N_noxref_12_c_3458_p N_noxref_14_M14_noxref_d ) capacitor \
 c=0.00742431f //x=26.38 //y=1.565 //x2=26.455 //y2=0.91
cc_2117 ( N_noxref_12_c_3346_n N_noxref_14_M14_noxref_d ) capacitor \
 c=0.00738639f //x=26.38 //y=1.92 //x2=26.455 //y2=0.91
cc_2118 ( N_noxref_12_c_3347_n N_noxref_14_M14_noxref_d ) capacitor \
 c=0.00220879f //x=26.755 //y=0.755 //x2=26.455 //y2=0.91
cc_2119 ( N_noxref_12_c_3399_n N_noxref_14_M14_noxref_d ) capacitor \
 c=0.0138055f //x=26.755 //y=1.41 //x2=26.455 //y2=0.91
cc_2120 ( N_noxref_12_c_3348_n N_noxref_14_M14_noxref_d ) capacitor \
 c=0.00218624f //x=26.91 //y=0.91 //x2=26.455 //y2=0.91
cc_2121 ( N_noxref_12_c_3350_n N_noxref_14_M14_noxref_d ) capacitor \
 c=0.00601286f //x=26.91 //y=1.255 //x2=26.455 //y2=0.91
cc_2122 ( N_noxref_12_c_3368_n N_noxref_14_M49_noxref_d ) capacitor \
 c=5.78106e-19 //x=24.79 //y=3.33 //x2=26.5 //y2=5.02
cc_2123 ( N_noxref_12_M49_noxref_g N_noxref_14_M49_noxref_d ) capacitor \
 c=0.0221134f //x=26.425 //y=6.02 //x2=26.5 //y2=5.02
cc_2124 ( N_noxref_12_M50_noxref_g N_noxref_14_M49_noxref_d ) capacitor \
 c=0.0220851f //x=26.865 //y=6.02 //x2=26.5 //y2=5.02
cc_2125 ( N_noxref_12_c_3379_n N_noxref_14_M49_noxref_d ) capacitor \
 c=0.0139997f //x=26.79 //y=4.79 //x2=26.5 //y2=5.02
cc_2126 ( N_noxref_12_c_3380_n N_noxref_14_M49_noxref_d ) capacitor \
 c=0.00307344f //x=26.5 //y=4.79 //x2=26.5 //y2=5.02
cc_2127 ( N_noxref_12_c_3395_n N_noxref_25_c_4415_n ) capacitor c=3.15806e-19 \
 //x=24.435 //y=1.655 //x2=22.895 //y2=1.495
cc_2128 ( N_noxref_12_c_3395_n N_noxref_25_c_4423_n ) capacitor c=0.0201674f \
 //x=24.435 //y=1.655 //x2=23.865 //y2=1.495
cc_2129 ( N_noxref_12_c_3337_n N_noxref_25_c_4424_n ) capacitor c=0.00510677f \
 //x=24.705 //y=1.655 //x2=24.75 //y2=0.53
cc_2130 ( N_noxref_12_M13_noxref_d N_noxref_25_c_4424_n ) capacitor \
 c=0.0114445f //x=24.16 //y=0.905 //x2=24.75 //y2=0.53
cc_2131 ( N_noxref_12_c_3337_n N_noxref_25_M12_noxref_s ) capacitor \
 c=0.0135507f //x=24.705 //y=1.655 //x2=22.76 //y2=0.365
cc_2132 ( N_noxref_12_M13_noxref_d N_noxref_25_M12_noxref_s ) capacitor \
 c=0.0437911f //x=24.16 //y=0.905 //x2=22.76 //y2=0.365
cc_2133 ( N_noxref_13_c_3497_n N_noxref_14_c_3617_n ) capacitor c=0.140643f \
 //x=31.705 //y=3.33 //x2=34.295 //y2=2.96
cc_2134 ( N_noxref_13_c_3500_n N_noxref_14_c_3617_n ) capacitor c=0.0292689f \
 //x=30.455 //y=3.33 //x2=34.295 //y2=2.96
cc_2135 ( N_noxref_13_c_3502_n N_noxref_14_c_3617_n ) capacitor c=0.00672451f \
 //x=29.775 //y=5.2 //x2=34.295 //y2=2.96
cc_2136 ( N_noxref_13_c_3506_n N_noxref_14_c_3617_n ) capacitor c=0.00655208f \
 //x=29.065 //y=5.2 //x2=34.295 //y2=2.96
cc_2137 ( N_noxref_13_c_3579_p N_noxref_14_c_3617_n ) capacitor c=0.00745069f \
 //x=29.985 //y=1.655 //x2=34.295 //y2=2.96
cc_2138 ( N_noxref_13_c_3477_n N_noxref_14_c_3617_n ) capacitor c=0.0254565f \
 //x=30.34 //y=3.33 //x2=34.295 //y2=2.96
cc_2139 ( N_noxref_13_c_3478_n N_noxref_14_c_3617_n ) capacitor c=0.0247839f \
 //x=31.82 //y=2.085 //x2=34.295 //y2=2.96
cc_2140 ( N_noxref_13_c_3490_n N_noxref_14_c_3617_n ) capacitor c=0.00335064f \
 //x=31.82 //y=2.085 //x2=34.295 //y2=2.96
cc_2141 ( N_noxref_13_c_3478_n N_noxref_14_c_3632_n ) capacitor c=8.15748e-19 \
 //x=31.82 //y=2.085 //x2=34.41 //y2=2.08
cc_2142 ( N_noxref_13_c_3497_n N_noxref_15_c_3803_n ) capacitor c=0.023945f \
 //x=31.705 //y=3.33 //x2=32.675 //y2=3.33
cc_2143 ( N_noxref_13_c_3478_n N_noxref_15_c_3803_n ) capacitor c=0.00245229f \
 //x=31.82 //y=2.085 //x2=32.675 //y2=3.33
cc_2144 ( N_noxref_13_c_3586_p N_noxref_15_c_3783_n ) capacitor c=0.0023507f \
 //x=32.305 //y=1.41 //x2=32.475 //y2=2.08
cc_2145 ( N_noxref_13_c_3490_n N_noxref_15_c_3824_n ) capacitor c=0.0136603f \
 //x=31.82 //y=2.085 //x2=32.275 //y2=2.08
cc_2146 ( N_noxref_13_c_3522_n N_noxref_15_c_3805_n ) capacitor c=0.0101013f \
 //x=32.34 //y=4.79 //x2=32.475 //y2=4.58
cc_2147 ( N_noxref_13_c_3478_n N_noxref_15_c_3808_n ) capacitor c=0.0250497f \
 //x=31.82 //y=2.085 //x2=32.28 //y2=4.58
cc_2148 ( N_noxref_13_c_3523_n N_noxref_15_c_3808_n ) capacitor c=0.00723812f \
 //x=32.05 //y=4.79 //x2=32.28 //y2=4.58
cc_2149 ( N_noxref_13_c_3497_n N_noxref_15_c_3786_n ) capacitor c=0.00197285f \
 //x=31.705 //y=3.33 //x2=32.56 //y2=3.33
cc_2150 ( N_noxref_13_c_3477_n N_noxref_15_c_3786_n ) capacitor c=7.75719e-19 \
 //x=30.34 //y=3.33 //x2=32.56 //y2=3.33
cc_2151 ( N_noxref_13_c_3478_n N_noxref_15_c_3786_n ) capacitor c=0.0684818f \
 //x=31.82 //y=2.085 //x2=32.56 //y2=3.33
cc_2152 ( N_noxref_13_c_3490_n N_noxref_15_c_3786_n ) capacitor c=5.85261e-19 \
 //x=31.82 //y=2.085 //x2=32.56 //y2=3.33
cc_2153 ( N_noxref_13_c_3477_n N_noxref_15_M17_noxref_d ) capacitor \
 c=3.32322e-19 //x=30.34 //y=3.33 //x2=32.005 //y2=0.91
cc_2154 ( N_noxref_13_c_3478_n N_noxref_15_M17_noxref_d ) capacitor \
 c=0.0174384f //x=31.82 //y=2.085 //x2=32.005 //y2=0.91
cc_2155 ( N_noxref_13_c_3483_n N_noxref_15_M17_noxref_d ) capacitor \
 c=0.00218556f //x=31.93 //y=0.91 //x2=32.005 //y2=0.91
cc_2156 ( N_noxref_13_c_3598_p N_noxref_15_M17_noxref_d ) capacitor \
 c=0.00347355f //x=31.93 //y=1.255 //x2=32.005 //y2=0.91
cc_2157 ( N_noxref_13_c_3599_p N_noxref_15_M17_noxref_d ) capacitor \
 c=0.00742431f //x=31.93 //y=1.565 //x2=32.005 //y2=0.91
cc_2158 ( N_noxref_13_c_3485_n N_noxref_15_M17_noxref_d ) capacitor \
 c=0.00784742f //x=31.93 //y=1.92 //x2=32.005 //y2=0.91
cc_2159 ( N_noxref_13_c_3486_n N_noxref_15_M17_noxref_d ) capacitor \
 c=0.00220879f //x=32.305 //y=0.755 //x2=32.005 //y2=0.91
cc_2160 ( N_noxref_13_c_3586_p N_noxref_15_M17_noxref_d ) capacitor \
 c=0.0138447f //x=32.305 //y=1.41 //x2=32.005 //y2=0.91
cc_2161 ( N_noxref_13_c_3487_n N_noxref_15_M17_noxref_d ) capacitor \
 c=0.00218624f //x=32.46 //y=0.91 //x2=32.005 //y2=0.91
cc_2162 ( N_noxref_13_c_3489_n N_noxref_15_M17_noxref_d ) capacitor \
 c=0.00601286f //x=32.46 //y=1.255 //x2=32.005 //y2=0.91
cc_2163 ( N_noxref_13_c_3477_n N_noxref_15_M55_noxref_d ) capacitor \
 c=6.34797e-19 //x=30.34 //y=3.33 //x2=32.05 //y2=5.02
cc_2164 ( N_noxref_13_M55_noxref_g N_noxref_15_M55_noxref_d ) capacitor \
 c=0.0219309f //x=31.975 //y=6.02 //x2=32.05 //y2=5.02
cc_2165 ( N_noxref_13_M56_noxref_g N_noxref_15_M55_noxref_d ) capacitor \
 c=0.021902f //x=32.415 //y=6.02 //x2=32.05 //y2=5.02
cc_2166 ( N_noxref_13_c_3522_n N_noxref_15_M55_noxref_d ) capacitor \
 c=0.0148755f //x=32.34 //y=4.79 //x2=32.05 //y2=5.02
cc_2167 ( N_noxref_13_c_3523_n N_noxref_15_M55_noxref_d ) capacitor \
 c=0.00307344f //x=32.05 //y=4.79 //x2=32.05 //y2=5.02
cc_2168 ( N_noxref_13_c_3497_n N_noxref_16_c_3925_n ) capacitor c=4.2915e-19 \
 //x=31.705 //y=3.33 //x2=36.005 //y2=3.33
cc_2169 ( N_noxref_13_c_3579_p N_noxref_26_c_4468_n ) capacitor c=3.15806e-19 \
 //x=29.985 //y=1.655 //x2=28.445 //y2=1.495
cc_2170 ( N_noxref_13_c_3579_p N_noxref_26_c_4476_n ) capacitor c=0.0201674f \
 //x=29.985 //y=1.655 //x2=29.415 //y2=1.495
cc_2171 ( N_noxref_13_c_3475_n N_noxref_26_c_4477_n ) capacitor c=0.00464204f \
 //x=30.255 //y=1.655 //x2=30.3 //y2=0.53
cc_2172 ( N_noxref_13_M16_noxref_d N_noxref_26_c_4477_n ) capacitor \
 c=0.0117318f //x=29.71 //y=0.905 //x2=30.3 //y2=0.53
cc_2173 ( N_noxref_13_c_3475_n N_noxref_26_M15_noxref_s ) capacitor \
 c=0.0140283f //x=30.255 //y=1.655 //x2=28.31 //y2=0.365
cc_2174 ( N_noxref_13_M16_noxref_d N_noxref_26_M15_noxref_s ) capacitor \
 c=0.0437911f //x=29.71 //y=0.905 //x2=28.31 //y2=0.365
cc_2175 ( N_noxref_14_c_3617_n N_noxref_15_c_3782_n ) capacitor c=0.173431f \
 //x=34.295 //y=2.96 //x2=35.035 //y2=3.33
cc_2176 ( N_noxref_14_c_3632_n N_noxref_15_c_3782_n ) capacitor c=0.0268861f \
 //x=34.41 //y=2.08 //x2=35.035 //y2=3.33
cc_2177 ( N_noxref_14_c_3656_n N_noxref_15_c_3782_n ) capacitor c=0.00510216f \
 //x=34.255 //y=4.705 //x2=35.035 //y2=3.33
cc_2178 ( N_noxref_14_c_3617_n N_noxref_15_c_3803_n ) capacitor c=0.029061f \
 //x=34.295 //y=2.96 //x2=32.675 //y2=3.33
cc_2179 ( N_noxref_14_c_3632_n N_noxref_15_c_3803_n ) capacitor c=3.78304e-19 \
 //x=34.41 //y=2.08 //x2=32.675 //y2=3.33
cc_2180 ( N_noxref_14_c_3632_n N_noxref_15_c_3783_n ) capacitor c=0.0137292f \
 //x=34.41 //y=2.08 //x2=32.475 //y2=2.08
cc_2181 ( N_noxref_14_c_3617_n N_noxref_15_c_3824_n ) capacitor c=0.00763858f \
 //x=34.295 //y=2.96 //x2=32.275 //y2=2.08
cc_2182 ( N_noxref_14_c_3617_n N_noxref_15_c_3808_n ) capacitor c=0.00318102f \
 //x=34.295 //y=2.96 //x2=32.28 //y2=4.58
cc_2183 ( N_noxref_14_c_3617_n N_noxref_15_c_3786_n ) capacitor c=0.0259021f \
 //x=34.295 //y=2.96 //x2=32.56 //y2=3.33
cc_2184 ( N_noxref_14_c_3656_n N_noxref_15_c_3856_n ) capacitor c=0.0452802f \
 //x=34.255 //y=4.705 //x2=35.15 //y2=4.54
cc_2185 ( N_noxref_14_c_3734_p N_noxref_15_c_3856_n ) capacitor c=0.00146509f \
 //x=34.675 //y=4.795 //x2=35.15 //y2=4.54
cc_2186 ( N_noxref_14_c_3664_n N_noxref_15_c_3856_n ) capacitor c=0.00112871f \
 //x=34.255 //y=4.705 //x2=35.15 //y2=4.54
cc_2187 ( N_noxref_14_c_3617_n N_noxref_15_c_3787_n ) capacitor c=0.00735597f \
 //x=34.295 //y=2.96 //x2=35.15 //y2=2.08
cc_2188 ( N_noxref_14_c_3632_n N_noxref_15_c_3787_n ) capacitor c=0.0433387f \
 //x=34.41 //y=2.08 //x2=35.15 //y2=2.08
cc_2189 ( N_noxref_14_c_3637_n N_noxref_15_c_3787_n ) capacitor c=0.00308814f \
 //x=34.215 //y=1.915 //x2=35.15 //y2=2.08
cc_2190 ( N_noxref_14_M57_noxref_g N_noxref_15_M59_noxref_g ) capacitor \
 c=0.0100243f //x=34.31 //y=6.025 //x2=35.19 //y2=6.025
cc_2191 ( N_noxref_14_M58_noxref_g N_noxref_15_M59_noxref_g ) capacitor \
 c=0.107798f //x=34.75 //y=6.025 //x2=35.19 //y2=6.025
cc_2192 ( N_noxref_14_M58_noxref_g N_noxref_15_M60_noxref_g ) capacitor \
 c=0.0094155f //x=34.75 //y=6.025 //x2=35.63 //y2=6.025
cc_2193 ( N_noxref_14_c_3635_n N_noxref_15_c_3789_n ) capacitor c=0.00125788f \
 //x=34.215 //y=0.905 //x2=35.185 //y2=0.905
cc_2194 ( N_noxref_14_c_3640_n N_noxref_15_c_3789_n ) capacitor c=0.0126654f \
 //x=34.745 //y=0.905 //x2=35.185 //y2=0.905
cc_2195 ( N_noxref_14_c_3744_p N_noxref_15_c_3867_n ) capacitor c=0.00148539f \
 //x=34.215 //y=1.25 //x2=35.185 //y2=1.255
cc_2196 ( N_noxref_14_c_3745_p N_noxref_15_c_3867_n ) capacitor c=0.00105591f \
 //x=34.215 //y=1.56 //x2=35.185 //y2=1.255
cc_2197 ( N_noxref_14_c_3642_n N_noxref_15_c_3867_n ) capacitor c=0.0126654f \
 //x=34.745 //y=1.25 //x2=35.185 //y2=1.255
cc_2198 ( N_noxref_14_c_3745_p N_noxref_15_c_3870_n ) capacitor c=0.00109549f \
 //x=34.215 //y=1.56 //x2=35.185 //y2=1.56
cc_2199 ( N_noxref_14_c_3642_n N_noxref_15_c_3870_n ) capacitor c=0.00886999f \
 //x=34.745 //y=1.25 //x2=35.185 //y2=1.56
cc_2200 ( N_noxref_14_c_3642_n N_noxref_15_c_3792_n ) capacitor c=0.00123863f \
 //x=34.745 //y=1.25 //x2=35.56 //y2=1.405
cc_2201 ( N_noxref_14_c_3640_n N_noxref_15_c_3793_n ) capacitor c=0.00132934f \
 //x=34.745 //y=0.905 //x2=35.715 //y2=0.905
cc_2202 ( N_noxref_14_c_3642_n N_noxref_15_c_3874_n ) capacitor c=0.00150734f \
 //x=34.745 //y=1.25 //x2=35.715 //y2=1.255
cc_2203 ( N_noxref_14_c_3632_n N_noxref_15_c_3875_n ) capacitor c=0.00307062f \
 //x=34.41 //y=2.08 //x2=35.15 //y2=2.08
cc_2204 ( N_noxref_14_c_3637_n N_noxref_15_c_3875_n ) capacitor c=0.0179092f \
 //x=34.215 //y=1.915 //x2=35.15 //y2=2.08
cc_2205 ( N_noxref_14_c_3637_n N_noxref_15_c_3877_n ) capacitor c=0.00577193f \
 //x=34.215 //y=1.915 //x2=35.15 //y2=1.915
cc_2206 ( N_noxref_14_c_3656_n N_noxref_15_c_3878_n ) capacitor c=0.00336963f \
 //x=34.255 //y=4.705 //x2=35.185 //y2=4.705
cc_2207 ( N_noxref_14_c_3734_p N_noxref_15_c_3878_n ) capacitor c=0.020271f \
 //x=34.675 //y=4.795 //x2=35.185 //y2=4.705
cc_2208 ( N_noxref_14_c_3664_n N_noxref_15_c_3878_n ) capacitor c=0.00546725f \
 //x=34.255 //y=4.705 //x2=35.185 //y2=4.705
cc_2209 ( N_noxref_14_c_3642_n N_noxref_16_c_3927_n ) capacitor c=0.00431513f \
 //x=34.745 //y=1.25 //x2=35.365 //y2=1.655
cc_2210 ( N_noxref_14_c_3617_n N_noxref_16_c_3986_n ) capacitor c=0.00116459f \
 //x=34.295 //y=2.96 //x2=34.565 //y2=1.655
cc_2211 ( N_noxref_14_c_3632_n N_noxref_16_c_3986_n ) capacitor c=0.0108811f \
 //x=34.41 //y=2.08 //x2=34.565 //y2=1.655
cc_2212 ( N_noxref_14_c_3637_n N_noxref_16_c_3986_n ) capacitor c=0.00524371f \
 //x=34.215 //y=1.915 //x2=34.565 //y2=1.655
cc_2213 ( N_noxref_14_c_3632_n N_noxref_16_c_3936_n ) capacitor c=0.00373525f \
 //x=34.41 //y=2.08 //x2=35.89 //y2=3.33
cc_2214 ( N_noxref_14_c_3635_n N_noxref_16_M18_noxref_d ) capacitor \
 c=0.0013184f //x=34.215 //y=0.905 //x2=34.29 //y2=0.905
cc_2215 ( N_noxref_14_c_3744_p N_noxref_16_M18_noxref_d ) capacitor \
 c=0.0034598f //x=34.215 //y=1.25 //x2=34.29 //y2=0.905
cc_2216 ( N_noxref_14_c_3745_p N_noxref_16_M18_noxref_d ) capacitor \
 c=0.00300148f //x=34.215 //y=1.56 //x2=34.29 //y2=0.905
cc_2217 ( N_noxref_14_c_3637_n N_noxref_16_M18_noxref_d ) capacitor \
 c=0.00273686f //x=34.215 //y=1.915 //x2=34.29 //y2=0.905
cc_2218 ( N_noxref_14_c_3639_n N_noxref_16_M18_noxref_d ) capacitor \
 c=0.00241102f //x=34.59 //y=0.75 //x2=34.29 //y2=0.905
cc_2219 ( N_noxref_14_c_3768_p N_noxref_16_M18_noxref_d ) capacitor \
 c=0.0123304f //x=34.59 //y=1.405 //x2=34.29 //y2=0.905
cc_2220 ( N_noxref_14_c_3640_n N_noxref_16_M18_noxref_d ) capacitor \
 c=0.00219619f //x=34.745 //y=0.905 //x2=34.29 //y2=0.905
cc_2221 ( N_noxref_14_c_3642_n N_noxref_16_M18_noxref_d ) capacitor \
 c=0.00603828f //x=34.745 //y=1.25 //x2=34.29 //y2=0.905
cc_2222 ( N_noxref_14_c_3617_n N_noxref_26_c_4477_n ) capacitor c=2.8058e-19 \
 //x=34.295 //y=2.96 //x2=30.3 //y2=0.53
cc_2223 ( N_noxref_14_c_3617_n N_noxref_26_M15_noxref_s ) capacitor \
 c=6.20367e-19 //x=34.295 //y=2.96 //x2=28.31 //y2=0.365
cc_2224 ( N_noxref_14_c_3656_n N_noxref_27_c_4525_n ) capacitor c=0.00617454f \
 //x=34.255 //y=4.705 //x2=34.885 //y2=5.21
cc_2225 ( N_noxref_14_M57_noxref_g N_noxref_27_c_4525_n ) capacitor \
 c=0.0182391f //x=34.31 //y=6.025 //x2=34.885 //y2=5.21
cc_2226 ( N_noxref_14_M58_noxref_g N_noxref_27_c_4525_n ) capacitor \
 c=0.0192395f //x=34.75 //y=6.025 //x2=34.885 //y2=5.21
cc_2227 ( N_noxref_14_c_3734_p N_noxref_27_c_4525_n ) capacitor c=0.00346501f \
 //x=34.675 //y=4.795 //x2=34.885 //y2=5.21
cc_2228 ( N_noxref_14_c_3664_n N_noxref_27_c_4525_n ) capacitor c=0.0017421f \
 //x=34.255 //y=4.705 //x2=34.885 //y2=5.21
cc_2229 ( N_noxref_14_c_3656_n N_noxref_27_c_4530_n ) capacitor c=0.0119751f \
 //x=34.255 //y=4.705 //x2=34.175 //y2=5.21
cc_2230 ( N_noxref_14_c_3664_n N_noxref_27_c_4530_n ) capacitor c=0.00524594f \
 //x=34.255 //y=4.705 //x2=34.175 //y2=5.21
cc_2231 ( N_noxref_14_M57_noxref_g N_noxref_27_M57_noxref_s ) capacitor \
 c=0.0473218f //x=34.31 //y=6.025 //x2=33.955 //y2=5.025
cc_2232 ( N_noxref_14_M58_noxref_g N_noxref_27_M58_noxref_d ) capacitor \
 c=0.0170604f //x=34.75 //y=6.025 //x2=34.825 //y2=5.025
cc_2233 ( N_noxref_15_c_3782_n N_noxref_16_c_3925_n ) capacitor c=0.023945f \
 //x=35.035 //y=3.33 //x2=36.005 //y2=3.33
cc_2234 ( N_noxref_15_c_3787_n N_noxref_16_c_3925_n ) capacitor c=0.00197285f \
 //x=35.15 //y=2.08 //x2=36.005 //y2=3.33
cc_2235 ( N_noxref_15_c_3782_n N_noxref_16_c_3927_n ) capacitor c=0.00172904f \
 //x=35.035 //y=3.33 //x2=35.365 //y2=1.655
cc_2236 ( N_noxref_15_c_3787_n N_noxref_16_c_3927_n ) capacitor c=0.0164694f \
 //x=35.15 //y=2.08 //x2=35.365 //y2=1.655
cc_2237 ( N_noxref_15_c_3870_n N_noxref_16_c_3927_n ) capacitor c=0.0021898f \
 //x=35.185 //y=1.56 //x2=35.365 //y2=1.655
cc_2238 ( N_noxref_15_c_3875_n N_noxref_16_c_3927_n ) capacitor c=0.00635719f \
 //x=35.15 //y=2.08 //x2=35.365 //y2=1.655
cc_2239 ( N_noxref_15_c_3877_n N_noxref_16_c_3927_n ) capacitor c=0.0189485f \
 //x=35.15 //y=1.915 //x2=35.365 //y2=1.655
cc_2240 ( N_noxref_15_c_3782_n N_noxref_16_c_3986_n ) capacitor c=0.00581867f \
 //x=35.035 //y=3.33 //x2=34.565 //y2=1.655
cc_2241 ( N_noxref_15_M60_noxref_g N_noxref_16_c_3964_n ) capacitor \
 c=0.0217686f //x=35.63 //y=6.025 //x2=35.805 //y2=5.21
cc_2242 ( N_noxref_15_M59_noxref_g N_noxref_16_c_3966_n ) capacitor \
 c=0.0132788f //x=35.19 //y=6.025 //x2=35.495 //y2=5.21
cc_2243 ( N_noxref_15_c_3891_p N_noxref_16_c_3966_n ) capacitor c=0.00410596f \
 //x=35.555 //y=4.795 //x2=35.495 //y2=5.21
cc_2244 ( N_noxref_15_c_3792_n N_noxref_16_c_3931_n ) capacitor c=0.00801563f \
 //x=35.56 //y=1.405 //x2=35.805 //y2=1.655
cc_2245 ( N_noxref_15_c_3782_n N_noxref_16_c_3936_n ) capacitor c=0.00245229f \
 //x=35.035 //y=3.33 //x2=35.89 //y2=3.33
cc_2246 ( N_noxref_15_c_3856_n N_noxref_16_c_3936_n ) capacitor c=0.0102183f \
 //x=35.15 //y=4.54 //x2=35.89 //y2=3.33
cc_2247 ( N_noxref_15_c_3787_n N_noxref_16_c_3936_n ) capacitor c=0.0816612f \
 //x=35.15 //y=2.08 //x2=35.89 //y2=3.33
cc_2248 ( N_noxref_15_c_3891_p N_noxref_16_c_3936_n ) capacitor c=0.0144455f \
 //x=35.555 //y=4.795 //x2=35.89 //y2=3.33
cc_2249 ( N_noxref_15_c_3875_n N_noxref_16_c_3936_n ) capacitor c=0.00877984f \
 //x=35.15 //y=2.08 //x2=35.89 //y2=3.33
cc_2250 ( N_noxref_15_c_3877_n N_noxref_16_c_3936_n ) capacitor c=0.00306024f \
 //x=35.15 //y=1.915 //x2=35.89 //y2=3.33
cc_2251 ( N_noxref_15_c_3878_n N_noxref_16_c_3936_n ) capacitor c=0.00537091f \
 //x=35.185 //y=4.705 //x2=35.89 //y2=3.33
cc_2252 ( N_noxref_15_c_3787_n N_noxref_16_c_3937_n ) capacitor c=0.00106083f \
 //x=35.15 //y=2.08 //x2=37.37 //y2=2.085
cc_2253 ( N_noxref_15_c_3870_n N_noxref_16_M18_noxref_d ) capacitor \
 c=0.00148728f //x=35.185 //y=1.56 //x2=34.29 //y2=0.905
cc_2254 ( N_noxref_15_c_3789_n N_noxref_16_M19_noxref_d ) capacitor \
 c=0.00226395f //x=35.185 //y=0.905 //x2=35.26 //y2=0.905
cc_2255 ( N_noxref_15_c_3867_n N_noxref_16_M19_noxref_d ) capacitor \
 c=0.0035101f //x=35.185 //y=1.255 //x2=35.26 //y2=0.905
cc_2256 ( N_noxref_15_c_3870_n N_noxref_16_M19_noxref_d ) capacitor \
 c=0.00546704f //x=35.185 //y=1.56 //x2=35.26 //y2=0.905
cc_2257 ( N_noxref_15_c_3791_n N_noxref_16_M19_noxref_d ) capacitor \
 c=0.00241102f //x=35.56 //y=0.75 //x2=35.26 //y2=0.905
cc_2258 ( N_noxref_15_c_3792_n N_noxref_16_M19_noxref_d ) capacitor \
 c=0.0158021f //x=35.56 //y=1.405 //x2=35.26 //y2=0.905
cc_2259 ( N_noxref_15_c_3793_n N_noxref_16_M19_noxref_d ) capacitor \
 c=0.00132831f //x=35.715 //y=0.905 //x2=35.26 //y2=0.905
cc_2260 ( N_noxref_15_c_3874_n N_noxref_16_M19_noxref_d ) capacitor \
 c=0.0035101f //x=35.715 //y=1.255 //x2=35.26 //y2=0.905
cc_2261 ( N_noxref_15_c_3877_n N_noxref_16_M19_noxref_d ) capacitor \
 c=3.4952e-19 //x=35.15 //y=1.915 //x2=35.26 //y2=0.905
cc_2262 ( N_noxref_15_M60_noxref_g N_noxref_16_M59_noxref_d ) capacitor \
 c=0.0136385f //x=35.63 //y=6.025 //x2=35.265 //y2=5.025
cc_2263 ( N_noxref_15_c_3782_n N_noxref_27_c_4525_n ) capacitor c=0.00894443f \
 //x=35.035 //y=3.33 //x2=34.885 //y2=5.21
cc_2264 ( N_noxref_15_M59_noxref_g N_noxref_27_c_4525_n ) capacitor \
 c=0.0170604f //x=35.19 //y=6.025 //x2=34.885 //y2=5.21
cc_2265 ( N_noxref_15_c_3878_n N_noxref_27_c_4525_n ) capacitor c=2.3112e-19 \
 //x=35.185 //y=4.705 //x2=34.885 //y2=5.21
cc_2266 ( N_noxref_15_c_3782_n N_noxref_27_c_4530_n ) capacitor c=0.00198612f \
 //x=35.035 //y=3.33 //x2=34.175 //y2=5.21
cc_2267 ( N_noxref_15_c_3856_n N_noxref_27_c_4532_n ) capacitor c=8.92402e-19 \
 //x=35.15 //y=4.54 //x2=35.765 //y2=6.91
cc_2268 ( N_noxref_15_M59_noxref_g N_noxref_27_c_4532_n ) capacitor \
 c=0.0148484f //x=35.19 //y=6.025 //x2=35.765 //y2=6.91
cc_2269 ( N_noxref_15_M60_noxref_g N_noxref_27_c_4532_n ) capacitor \
 c=0.0163196f //x=35.63 //y=6.025 //x2=35.765 //y2=6.91
cc_2270 ( N_noxref_15_M60_noxref_g N_noxref_27_M60_noxref_d ) capacitor \
 c=0.0351101f //x=35.63 //y=6.025 //x2=35.705 //y2=5.025
cc_2271 ( N_noxref_16_c_3966_n N_noxref_27_c_4525_n ) capacitor c=0.0348754f \
 //x=35.495 //y=5.21 //x2=34.885 //y2=5.21
cc_2272 ( N_noxref_16_c_3964_n N_noxref_27_c_4532_n ) capacitor c=0.00173777f \
 //x=35.805 //y=5.21 //x2=35.765 //y2=6.91
cc_2273 ( N_noxref_16_M59_noxref_d N_noxref_27_c_4532_n ) capacitor \
 c=0.0118172f //x=35.265 //y=5.025 //x2=35.765 //y2=6.91
cc_2274 ( N_noxref_16_M59_noxref_d N_noxref_27_M57_noxref_s ) capacitor \
 c=0.00107541f //x=35.265 //y=5.025 //x2=33.955 //y2=5.025
cc_2275 ( N_noxref_16_M59_noxref_d N_noxref_27_M58_noxref_d ) capacitor \
 c=0.0348754f //x=35.265 //y=5.025 //x2=34.825 //y2=5.025
cc_2276 ( N_noxref_16_c_3964_n N_noxref_27_M60_noxref_d ) capacitor \
 c=0.015774f //x=35.805 //y=5.21 //x2=35.705 //y2=5.025
cc_2277 ( N_noxref_16_M59_noxref_d N_noxref_27_M60_noxref_d ) capacitor \
 c=0.0458293f //x=35.265 //y=5.025 //x2=35.705 //y2=5.025
cc_2278 ( N_noxref_16_c_3919_n COUT ) capacitor c=0.00423952f //x=37.255 \
 //y=3.33 //x2=38.11 //y2=2.22
cc_2279 ( N_noxref_16_c_3936_n COUT ) capacitor c=0.00126776f //x=35.89 \
 //y=3.33 //x2=38.11 //y2=2.22
cc_2280 ( N_noxref_16_c_3937_n COUT ) capacitor c=0.0711303f //x=37.37 \
 //y=2.085 //x2=38.11 //y2=2.22
cc_2281 ( N_noxref_16_c_3949_n COUT ) capacitor c=8.49451e-19 //x=37.37 \
 //y=2.085 //x2=38.11 //y2=2.22
cc_2282 ( N_noxref_16_c_4039_p N_COUT_c_4568_n ) capacitor c=0.0023507f \
 //x=37.855 //y=1.41 //x2=38.025 //y2=2.08
cc_2283 ( N_noxref_16_c_3949_n N_COUT_c_4592_n ) capacitor c=0.0167852f \
 //x=37.37 //y=2.085 //x2=37.825 //y2=2.08
cc_2284 ( N_noxref_16_c_3978_n N_COUT_c_4578_n ) capacitor c=0.0101013f \
 //x=37.89 //y=4.79 //x2=38.025 //y2=4.58
cc_2285 ( N_noxref_16_c_3937_n N_COUT_c_4581_n ) capacitor c=0.0250878f \
 //x=37.37 //y=2.085 //x2=37.83 //y2=4.58
cc_2286 ( N_noxref_16_c_3979_n N_COUT_c_4581_n ) capacitor c=0.00962086f \
 //x=37.6 //y=4.79 //x2=37.83 //y2=4.58
cc_2287 ( N_noxref_16_c_3936_n N_COUT_M20_noxref_d ) capacitor c=3.35192e-19 \
 //x=35.89 //y=3.33 //x2=37.555 //y2=0.91
cc_2288 ( N_noxref_16_c_3937_n N_COUT_M20_noxref_d ) capacitor c=0.0175773f \
 //x=37.37 //y=2.085 //x2=37.555 //y2=0.91
cc_2289 ( N_noxref_16_c_3942_n N_COUT_M20_noxref_d ) capacitor c=0.00218556f \
 //x=37.48 //y=0.91 //x2=37.555 //y2=0.91
cc_2290 ( N_noxref_16_c_4047_p N_COUT_M20_noxref_d ) capacitor c=0.00347355f \
 //x=37.48 //y=1.255 //x2=37.555 //y2=0.91
cc_2291 ( N_noxref_16_c_4048_p N_COUT_M20_noxref_d ) capacitor c=0.00742431f \
 //x=37.48 //y=1.565 //x2=37.555 //y2=0.91
cc_2292 ( N_noxref_16_c_3944_n N_COUT_M20_noxref_d ) capacitor c=0.00957707f \
 //x=37.48 //y=1.92 //x2=37.555 //y2=0.91
cc_2293 ( N_noxref_16_c_3945_n N_COUT_M20_noxref_d ) capacitor c=0.00220879f \
 //x=37.855 //y=0.755 //x2=37.555 //y2=0.91
cc_2294 ( N_noxref_16_c_4039_p N_COUT_M20_noxref_d ) capacitor c=0.0138447f \
 //x=37.855 //y=1.41 //x2=37.555 //y2=0.91
cc_2295 ( N_noxref_16_c_3946_n N_COUT_M20_noxref_d ) capacitor c=0.00218624f \
 //x=38.01 //y=0.91 //x2=37.555 //y2=0.91
cc_2296 ( N_noxref_16_c_3948_n N_COUT_M20_noxref_d ) capacitor c=0.00601286f \
 //x=38.01 //y=1.255 //x2=37.555 //y2=0.91
cc_2297 ( N_noxref_16_c_3936_n N_COUT_M61_noxref_d ) capacitor c=6.2839e-19 \
 //x=35.89 //y=3.33 //x2=37.6 //y2=5.02
cc_2298 ( N_noxref_16_M61_noxref_g N_COUT_M61_noxref_d ) capacitor \
 c=0.0219309f //x=37.525 //y=6.02 //x2=37.6 //y2=5.02
cc_2299 ( N_noxref_16_M62_noxref_g N_COUT_M61_noxref_d ) capacitor c=0.021902f \
 //x=37.965 //y=6.02 //x2=37.6 //y2=5.02
cc_2300 ( N_noxref_16_c_3978_n N_COUT_M61_noxref_d ) capacitor c=0.0148755f \
 //x=37.89 //y=4.79 //x2=37.6 //y2=5.02
cc_2301 ( N_noxref_16_c_3979_n N_COUT_M61_noxref_d ) capacitor c=0.00307344f \
 //x=37.6 //y=4.79 //x2=37.6 //y2=5.02
cc_2302 ( N_noxref_17_M26_noxref_d N_noxref_19_M27_noxref_s ) capacitor \
 c=0.00181587f //x=4.625 //y=5.02 //x2=6.205 //y2=5.02
cc_2303 ( N_noxref_18_c_4110_n N_noxref_20_M3_noxref_s ) capacitor \
 c=0.00174327f //x=4.855 //y=0.62 //x2=6.11 //y2=0.37
cc_2304 ( N_noxref_21_M38_noxref_d N_noxref_23_M39_noxref_s ) capacitor \
 c=0.00181587f //x=15.725 //y=5.02 //x2=17.305 //y2=5.02
cc_2305 ( N_noxref_22_c_4289_n N_noxref_24_M9_noxref_s ) capacitor \
 c=0.00174327f //x=15.955 //y=0.62 //x2=17.21 //y2=0.37
