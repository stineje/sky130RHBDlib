* SPICE3 file created from TMRDFFRNQX1.ext - technology: sky130A

.subckt TMRDFFRNQX1 Q D CLK RN VDD GND
M1000 a_5779_989.t2 RN.t0 VDD.t35 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_9009_1050.t2 a_9331_989.t5 VDD.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 Q.t2 a_15932_209.t7 VDD.t101 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_5457_1050.t6 CLK.t0 VDD.t95 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 GND a_9331_989.t7 a_16318_101.t0 nshort w=-1.605u l=1.765u
+  ad=4.9019p pd=41.07u as=0p ps=0u
M1005 a_15757_1051.t3 a_9331_989.t6 a_16421_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VDD.t64 a_14511_989.t5 a_14189_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VDD.t39 RN.t1 a_147_187.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 GND a_5457_1050.t7 a_8823_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1009 VDD.t23 a_147_187.t8 a_4151_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VDD.t76 a_5327_187.t7 a_7321_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_16421_1051.t6 a_4151_989.t5 a_15932_209.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_14511_989.t0 a_14189_1050.t7 VDD.t10 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_12501_1050.t1 a_10959_989.t8 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 GND a_5457_1050.t8 a_6233_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1015 VDD.t31 RN.t3 a_10959_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_5457_1050.t1 a_5779_989.t7 VDD.t79 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_5327_187.t1 RN.t5 VDD.t43 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 GND a_9009_1050.t8 a_9806_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1019 VDD.t8 a_147_187.t9 a_277_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_15757_1051.t6 a_4151_989.t6 a_16421_1051.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VDD.t60 a_10507_187.t9 a_10637_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VDD.t14 a_12501_1050.t5 a_10507_187.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 GND a_5779_989.t9 a_7216_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1024 VDD.t32 RN.t6 a_10507_187.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 GND a_147_187.t10 a_91_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_14189_1050.t6 a_10637_1050.t7 VDD.t70 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 GND a_7321_1050.t5 a_7861_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_10959_989.t4 a_10637_1050.t8 VDD.t80 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_599_989.t4 D.t1 VDD.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_16421_1051.t7 a_14511_989.t7 a_15932_209.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 Q a_15932_209.t8 GND.t13 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1032 GND a_5327_187.t9 a_5271_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_5327_187.t5 CLK.t3 VDD.t85 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 VDD.t82 a_599_989.t8 a_2141_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_9331_989.t1 a_9009_1050.t7 VDD.t62 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 VDD.t54 CLK.t4 a_277_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VDD.t100 a_5457_1050.t9 a_5779_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 VDD.t57 a_5457_1050.t10 a_9009_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 VDD.t68 a_277_1050.t7 a_3829_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 VDD.t87 CLK.t5 a_10507_187.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 VDD.t36 RN.t8 a_5779_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 VDD.t21 a_9331_989.t8 a_9009_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1043 VDD.t4 CLK.t6 a_10637_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_9331_989.t4 a_5327_187.t8 VDD.t96 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_14189_1050.t2 RN.t9 VDD.t33 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_10959_989.t1 D.t2 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_599_989.t1 RN.t10 VDD.t34 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_3829_1050.t3 a_4151_989.t7 VDD.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_10637_1050.t3 a_10507_187.t10 VDD.t88 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 VDD.t9 a_14511_989.t9 a_15757_1051.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_147_187.t6 CLK.t7 VDD.t90 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 GND a_12501_1050.t6 a_13041_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1053 GND a_277_1050.t8 a_3643_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_4151_989.t0 a_3829_1050.t7 VDD.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 a_9009_1050.t3 a_5457_1050.t11 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 a_15757_1051.t1 a_9331_989.t9 VDD.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 VDD.t65 a_14189_1050.t8 a_14511_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 VDD.t2 a_10959_989.t9 a_12501_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1059 VDD.t7 a_147_187.t11 a_2141_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1060 VDD.t52 a_599_989.t9 a_277_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 VDD.t44 RN.t12 a_9009_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 VDD.t49 D.t4 a_5779_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 VDD.t86 a_2141_1050.t5 a_147_187.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1064 VDD.t67 a_5327_187.t11 a_5457_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 VDD.t77 a_7321_1050.t6 a_5327_187.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 GND a_3829_1050.t8 a_4626_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_14189_1050.t4 a_14511_989.t11 VDD.t74 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_10959_989.t6 RN.t13 VDD.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 GND a_599_989.t10 a_2036_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1070 a_147_187.t2 RN.t14 VDD.t37 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 GND a_10637_1050.t9 a_14003_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1072 GND a_2141_1050.t6 a_2681_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1073 a_4151_989.t2 a_147_187.t12 VDD.t93 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1074 a_7321_1050.t0 a_5327_187.t12 VDD.t75 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 a_15932_209.t2 a_4151_989.t9 a_16421_1051.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1076 VDD.t0 a_10959_989.t10 a_10637_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 a_15757_1051.t7 a_14511_989.t12 VDD.t83 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1078 VDD.t6 a_10507_187.t12 a_14511_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 VDD.t59 a_10507_187.t13 a_12501_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 VDD.t91 a_15932_209.t9 Q.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 GND a_9331_989.t10 a_15652_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1082 GND a_14189_1050.t9 a_14986_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_277_1050.t1 a_147_187.t13 VDD.t94 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 a_16421_1051.t2 a_4151_989.t11 a_15757_1051.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 VDD.t50 a_9009_1050.t9 a_9331_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_10507_187.t4 a_12501_1050.t7 VDD.t78 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 a_10637_1050.t1 a_10959_989.t11 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 a_10507_187.t2 RN.t15 VDD.t47 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 a_7321_1050.t4 a_5779_989.t10 VDD.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 VDD.t20 a_277_1050.t9 a_599_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 a_15932_209.t1 a_14511_989.t13 a_16421_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1092 VDD.t66 a_4151_989.t12 a_3829_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1093 VDD.t40 RN.t17 a_599_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 GND a_277_1050.t11 a_1053_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1095 a_2141_1050.t3 a_599_989.t11 VDD.t81 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1096 VDD.t25 a_5779_989.t11 a_5457_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 VDD.t41 RN.t19 a_5327_187.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 a_16421_1051.t1 a_9331_989.t11 a_15757_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1099 a_277_1050.t5 CLK.t11 VDD.t55 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 a_3829_1050.t5 a_277_1050.t10 VDD.t98 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1101 a_5779_989.t5 a_5457_1050.t12 VDD.t92 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 GND a_4151_989.t13 a_16984_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_10637_1050.t5 CLK.t12 VDD.t58 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 a_10507_187.t5 CLK.t13 VDD.t56 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 VDD.t15 a_10637_1050.t10 a_14189_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 VDD.t69 a_10637_1050.t11 a_10959_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 GND a_10637_1050.t12 a_11413_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1108 VDD.t53 D.t5 a_599_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 VDD.t38 RN.t21 a_3829_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 a_599_989.t5 a_277_1050.t12 VDD.t72 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 VDD.t27 CLK.t15 a_5327_187.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1112 VDD.t29 CLK.t16 a_5457_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1113 a_2141_1050.t1 a_147_187.t14 VDD.t73 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1114 GND a_10959_989.t7 a_12396_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1115 a_277_1050.t3 a_599_989.t12 VDD.t51 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1116 a_3829_1050.t0 RN.t23 VDD.t45 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1117 a_5779_989.t3 D.t6 VDD.t48 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1118 a_9009_1050.t4 RN.t24 VDD.t42 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1119 a_5457_1050.t3 a_5327_187.t14 VDD.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1120 a_5327_187.t6 a_7321_1050.t7 VDD.t97 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1121 VDD.t71 a_5327_187.t15 a_9331_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1122 a_147_187.t4 a_2141_1050.t7 VDD.t63 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1123 GND a_10507_187.t7 a_10451_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1124 VDD.t46 RN.t25 a_14189_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1125 VDD.t19 D.t7 a_10959_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1126 VDD.t28 CLK.t17 a_147_187.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1127 VDD.t84 a_3829_1050.t9 a_4151_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1128 VDD.t99 a_5779_989.t12 a_7321_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1129 VDD.t26 a_9331_989.t13 a_15757_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1130 a_14511_989.t1 a_10507_187.t14 VDD.t61 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1131 a_12501_1050.t3 a_10507_187.t15 VDD.t89 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 CLK VDD 1.71fF
C1 D VDD 0.15fF
C2 RN VDD 0.50fF
C3 Q VDD 0.76fF
C4 CLK D 0.45fF
C5 CLK RN 1.13fF
C6 D RN 12.60fF
R0 a_10959_989.n5 a_10959_989.t9 480.392
R1 a_10959_989.n7 a_10959_989.t11 454.685
R2 a_10959_989.n7 a_10959_989.t10 428.979
R3 a_10959_989.n5 a_10959_989.t8 403.272
R4 a_10959_989.n6 a_10959_989.t7 283.48
R5 a_10959_989.n8 a_10959_989.t12 237.959
R6 a_10959_989.n12 a_10959_989.n10 219.626
R7 a_10959_989.n10 a_10959_989.n4 170.799
R8 a_10959_989.n8 a_10959_989.n7 98.447
R9 a_10959_989.n6 a_10959_989.n5 98.447
R10 a_10959_989.n9 a_10959_989.n8 80.035
R11 a_10959_989.n3 a_10959_989.n2 79.232
R12 a_10959_989.n9 a_10959_989.n6 77.315
R13 a_10959_989.n10 a_10959_989.n9 76
R14 a_10959_989.n4 a_10959_989.n3 63.152
R15 a_10959_989.n4 a_10959_989.n0 16.08
R16 a_10959_989.n3 a_10959_989.n1 16.08
R17 a_10959_989.n12 a_10959_989.n11 15.218
R18 a_10959_989.n0 a_10959_989.t0 14.282
R19 a_10959_989.n0 a_10959_989.t6 14.282
R20 a_10959_989.n1 a_10959_989.t2 14.282
R21 a_10959_989.n1 a_10959_989.t1 14.282
R22 a_10959_989.n2 a_10959_989.t3 14.282
R23 a_10959_989.n2 a_10959_989.t4 14.282
R24 a_10959_989.n13 a_10959_989.n12 12.014
R25 a_12396_101.n10 a_12396_101.n9 93.333
R26 a_12396_101.n2 a_12396_101.n1 41.622
R27 a_12396_101.n13 a_12396_101.n12 26.667
R28 a_12396_101.n6 a_12396_101.n5 24.977
R29 a_12396_101.t0 a_12396_101.n2 21.209
R30 a_12396_101.t0 a_12396_101.n3 11.595
R31 a_12396_101.t1 a_12396_101.n8 8.137
R32 a_12396_101.t0 a_12396_101.n0 6.109
R33 a_12396_101.t1 a_12396_101.n7 4.864
R34 a_12396_101.t0 a_12396_101.n4 3.871
R35 a_12396_101.t0 a_12396_101.n13 2.535
R36 a_12396_101.n13 a_12396_101.t1 1.145
R37 a_12396_101.n7 a_12396_101.n6 1.13
R38 a_12396_101.t1 a_12396_101.n11 0.804
R39 a_12396_101.n11 a_12396_101.n10 0.136
R40 GND.n30 GND.n29 219.745
R41 GND.n60 GND.n58 219.745
R42 GND.n90 GND.n88 219.745
R43 GND.n451 GND.n450 219.745
R44 GND.n493 GND.n491 219.745
R45 GND.n526 GND.n524 219.745
R46 GND.n568 GND.n566 219.745
R47 GND.n610 GND.n608 219.745
R48 GND.n640 GND.n638 219.745
R49 GND.n682 GND.n680 219.745
R50 GND.n724 GND.n722 219.745
R51 GND.n754 GND.n752 219.745
R52 GND.n796 GND.n794 219.745
R53 GND.n381 GND.n379 219.745
R54 GND.n351 GND.n349 219.745
R55 GND.n309 GND.n307 219.745
R56 GND.n264 GND.n262 219.745
R57 GND.n234 GND.n232 219.745
R58 GND.n192 GND.n190 219.745
R59 GND.n150 GND.n148 219.745
R60 GND.n120 GND.n119 219.745
R61 GND.n181 GND.n180 85.559
R62 GND.n223 GND.n222 85.559
R63 GND.n340 GND.n339 85.559
R64 GND.n805 GND.n804 85.559
R65 GND.n763 GND.n762 85.559
R66 GND.n691 GND.n690 85.559
R67 GND.n649 GND.n648 85.559
R68 GND.n577 GND.n576 85.559
R69 GND.n535 GND.n534 85.559
R70 GND.n460 GND.n459 85.559
R71 GND.n418 GND.n417 85.559
R72 GND.n30 GND.n28 85.529
R73 GND.n60 GND.n59 85.529
R74 GND.n90 GND.n89 85.529
R75 GND.n451 GND.n449 85.529
R76 GND.n493 GND.n492 85.529
R77 GND.n526 GND.n525 85.529
R78 GND.n568 GND.n567 85.529
R79 GND.n610 GND.n609 85.529
R80 GND.n640 GND.n639 85.529
R81 GND.n682 GND.n681 85.529
R82 GND.n724 GND.n723 85.529
R83 GND.n754 GND.n753 85.529
R84 GND.n796 GND.n795 85.529
R85 GND.n381 GND.n380 85.529
R86 GND.n351 GND.n350 85.529
R87 GND.n309 GND.n308 85.529
R88 GND.n264 GND.n263 85.529
R89 GND.n234 GND.n233 85.529
R90 GND.n192 GND.n191 85.529
R91 GND.n150 GND.n149 85.529
R92 GND.n120 GND.n118 85.529
R93 GND.n78 GND.n77 84.842
R94 GND.n108 GND.n107 84.842
R95 GND.n138 GND.n137 84.842
R96 GND.n252 GND.n251 84.842
R97 GND.n369 GND.n368 84.842
R98 GND.n732 GND.n731 84.842
R99 GND.n618 GND.n617 84.842
R100 GND.n48 GND.n47 84.842
R101 GND.n9 GND.n1 76.145
R102 GND.n412 GND.n411 76
R103 GND.n73 GND.n72 76
R104 GND.n76 GND.n75 76
R105 GND.n81 GND.n80 76
R106 GND.n84 GND.n83 76
R107 GND.n87 GND.n86 76
R108 GND.n94 GND.n93 76
R109 GND.n97 GND.n96 76
R110 GND.n100 GND.n99 76
R111 GND.n103 GND.n102 76
R112 GND.n106 GND.n105 76
R113 GND.n111 GND.n110 76
R114 GND.n114 GND.n113 76
R115 GND.n117 GND.n116 76
R116 GND.n124 GND.n123 76
R117 GND.n127 GND.n126 76
R118 GND.n130 GND.n129 76
R119 GND.n133 GND.n132 76
R120 GND.n136 GND.n135 76
R121 GND.n141 GND.n140 76
R122 GND.n144 GND.n143 76
R123 GND.n147 GND.n146 76
R124 GND.n154 GND.n153 76
R125 GND.n157 GND.n156 76
R126 GND.n160 GND.n159 76
R127 GND.n163 GND.n162 76
R128 GND.n166 GND.n165 76
R129 GND.n169 GND.n168 76
R130 GND.n172 GND.n171 76
R131 GND.n175 GND.n174 76
R132 GND.n178 GND.n177 76
R133 GND.n183 GND.n182 76
R134 GND.n186 GND.n185 76
R135 GND.n189 GND.n188 76
R136 GND.n196 GND.n195 76
R137 GND.n199 GND.n198 76
R138 GND.n202 GND.n201 76
R139 GND.n205 GND.n204 76
R140 GND.n208 GND.n207 76
R141 GND.n211 GND.n210 76
R142 GND.n214 GND.n213 76
R143 GND.n217 GND.n216 76
R144 GND.n220 GND.n219 76
R145 GND.n225 GND.n224 76
R146 GND.n228 GND.n227 76
R147 GND.n231 GND.n230 76
R148 GND.n238 GND.n237 76
R149 GND.n241 GND.n240 76
R150 GND.n244 GND.n243 76
R151 GND.n247 GND.n246 76
R152 GND.n250 GND.n249 76
R153 GND.n255 GND.n254 76
R154 GND.n258 GND.n257 76
R155 GND.n261 GND.n260 76
R156 GND.n268 GND.n267 76
R157 GND.n271 GND.n270 76
R158 GND.n274 GND.n273 76
R159 GND.n277 GND.n276 76
R160 GND.n280 GND.n279 76
R161 GND.n283 GND.n282 76
R162 GND.n286 GND.n285 76
R163 GND.n289 GND.n288 76
R164 GND.n292 GND.n291 76
R165 GND.n300 GND.n299 76
R166 GND.n303 GND.n302 76
R167 GND.n306 GND.n305 76
R168 GND.n313 GND.n312 76
R169 GND.n316 GND.n315 76
R170 GND.n319 GND.n318 76
R171 GND.n322 GND.n321 76
R172 GND.n325 GND.n324 76
R173 GND.n328 GND.n327 76
R174 GND.n331 GND.n330 76
R175 GND.n334 GND.n333 76
R176 GND.n337 GND.n336 76
R177 GND.n342 GND.n341 76
R178 GND.n345 GND.n344 76
R179 GND.n348 GND.n347 76
R180 GND.n355 GND.n354 76
R181 GND.n358 GND.n357 76
R182 GND.n361 GND.n360 76
R183 GND.n364 GND.n363 76
R184 GND.n367 GND.n366 76
R185 GND.n372 GND.n371 76
R186 GND.n375 GND.n374 76
R187 GND.n378 GND.n377 76
R188 GND.n385 GND.n384 76
R189 GND.n388 GND.n387 76
R190 GND.n391 GND.n390 76
R191 GND.n394 GND.n393 76
R192 GND.n397 GND.n396 76
R193 GND.n400 GND.n399 76
R194 GND.n403 GND.n402 76
R195 GND.n406 GND.n405 76
R196 GND.n409 GND.n408 76
R197 GND.n807 GND.n806 76
R198 GND.n802 GND.n801 76
R199 GND.n799 GND.n798 76
R200 GND.n792 GND.n791 76
R201 GND.n789 GND.n788 76
R202 GND.n786 GND.n785 76
R203 GND.n783 GND.n782 76
R204 GND.n780 GND.n779 76
R205 GND.n777 GND.n776 76
R206 GND.n774 GND.n773 76
R207 GND.n771 GND.n770 76
R208 GND.n768 GND.n767 76
R209 GND.n765 GND.n764 76
R210 GND.n760 GND.n759 76
R211 GND.n757 GND.n756 76
R212 GND.n750 GND.n749 76
R213 GND.n747 GND.n746 76
R214 GND.n744 GND.n743 76
R215 GND.n741 GND.n740 76
R216 GND.n738 GND.n737 76
R217 GND.n735 GND.n734 76
R218 GND.n730 GND.n729 76
R219 GND.n727 GND.n726 76
R220 GND.n720 GND.n719 76
R221 GND.n717 GND.n716 76
R222 GND.n714 GND.n713 76
R223 GND.n711 GND.n710 76
R224 GND.n708 GND.n707 76
R225 GND.n705 GND.n704 76
R226 GND.n702 GND.n701 76
R227 GND.n699 GND.n698 76
R228 GND.n696 GND.n695 76
R229 GND.n693 GND.n692 76
R230 GND.n688 GND.n687 76
R231 GND.n685 GND.n684 76
R232 GND.n678 GND.n677 76
R233 GND.n675 GND.n674 76
R234 GND.n672 GND.n671 76
R235 GND.n669 GND.n668 76
R236 GND.n666 GND.n665 76
R237 GND.n663 GND.n662 76
R238 GND.n660 GND.n659 76
R239 GND.n657 GND.n656 76
R240 GND.n654 GND.n653 76
R241 GND.n651 GND.n650 76
R242 GND.n646 GND.n645 76
R243 GND.n643 GND.n642 76
R244 GND.n636 GND.n635 76
R245 GND.n633 GND.n632 76
R246 GND.n630 GND.n629 76
R247 GND.n627 GND.n626 76
R248 GND.n624 GND.n623 76
R249 GND.n621 GND.n620 76
R250 GND.n616 GND.n615 76
R251 GND.n613 GND.n612 76
R252 GND.n606 GND.n605 76
R253 GND.n603 GND.n602 76
R254 GND.n600 GND.n599 76
R255 GND.n597 GND.n596 76
R256 GND.n594 GND.n593 76
R257 GND.n591 GND.n590 76
R258 GND.n588 GND.n587 76
R259 GND.n585 GND.n584 76
R260 GND.n582 GND.n581 76
R261 GND.n579 GND.n578 76
R262 GND.n574 GND.n573 76
R263 GND.n571 GND.n570 76
R264 GND.n564 GND.n563 76
R265 GND.n561 GND.n560 76
R266 GND.n558 GND.n557 76
R267 GND.n555 GND.n554 76
R268 GND.n552 GND.n551 76
R269 GND.n549 GND.n548 76
R270 GND.n546 GND.n545 76
R271 GND.n543 GND.n542 76
R272 GND.n540 GND.n539 76
R273 GND.n537 GND.n536 76
R274 GND.n532 GND.n531 76
R275 GND.n529 GND.n528 76
R276 GND.n522 GND.n521 76
R277 GND.n519 GND.n518 76
R278 GND.n516 GND.n515 76
R279 GND.n513 GND.n512 76
R280 GND.n510 GND.n509 76
R281 GND.n507 GND.n506 76
R282 GND.n499 GND.n498 76
R283 GND.n496 GND.n495 76
R284 GND.n489 GND.n488 76
R285 GND.n486 GND.n485 76
R286 GND.n483 GND.n482 76
R287 GND.n480 GND.n479 76
R288 GND.n477 GND.n476 76
R289 GND.n474 GND.n473 76
R290 GND.n471 GND.n470 76
R291 GND.n468 GND.n467 76
R292 GND.n465 GND.n464 76
R293 GND.n462 GND.n461 76
R294 GND.n457 GND.n456 76
R295 GND.n454 GND.n453 76
R296 GND.n447 GND.n446 76
R297 GND.n444 GND.n443 76
R298 GND.n441 GND.n440 76
R299 GND.n438 GND.n437 76
R300 GND.n435 GND.n434 76
R301 GND.n432 GND.n431 76
R302 GND.n429 GND.n428 76
R303 GND.n426 GND.n425 76
R304 GND.n423 GND.n422 76
R305 GND.n420 GND.n419 76
R306 GND.n415 GND.n414 76
R307 GND.n9 GND.n8 76
R308 GND.n17 GND.n16 76
R309 GND.n24 GND.n23 76
R310 GND.n27 GND.n26 76
R311 GND.n34 GND.n33 76
R312 GND.n37 GND.n36 76
R313 GND.n40 GND.n39 76
R314 GND.n43 GND.n42 76
R315 GND.n46 GND.n45 76
R316 GND.n51 GND.n50 76
R317 GND.n54 GND.n53 76
R318 GND.n57 GND.n56 76
R319 GND.n64 GND.n63 76
R320 GND.n67 GND.n66 76
R321 GND.n70 GND.n69 76
R322 GND.n298 GND.n297 64.552
R323 GND.n504 GND.n503 63.835
R324 GND.n5 GND.n4 35.01
R325 GND.n3 GND.n2 29.127
R326 GND.n297 GND.n296 28.421
R327 GND.n503 GND.n502 28.421
R328 GND.n297 GND.n295 25.263
R329 GND.n503 GND.n501 25.263
R330 GND.n295 GND.n294 24.383
R331 GND.n501 GND.n500 24.383
R332 GND.n12 GND.t13 20.794
R333 GND.n6 GND.n5 19.735
R334 GND.n14 GND.n13 19.735
R335 GND.n21 GND.n20 19.735
R336 GND.n5 GND.n3 19.017
R337 GND.n33 GND.n31 14.167
R338 GND.n63 GND.n61 14.167
R339 GND.n93 GND.n91 14.167
R340 GND.n123 GND.n121 14.167
R341 GND.n153 GND.n151 14.167
R342 GND.n195 GND.n193 14.167
R343 GND.n237 GND.n235 14.167
R344 GND.n267 GND.n265 14.167
R345 GND.n312 GND.n310 14.167
R346 GND.n354 GND.n352 14.167
R347 GND.n384 GND.n382 14.167
R348 GND.n798 GND.n797 14.167
R349 GND.n756 GND.n755 14.167
R350 GND.n726 GND.n725 14.167
R351 GND.n684 GND.n683 14.167
R352 GND.n642 GND.n641 14.167
R353 GND.n612 GND.n611 14.167
R354 GND.n570 GND.n569 14.167
R355 GND.n528 GND.n527 14.167
R356 GND.n495 GND.n494 14.167
R357 GND.n453 GND.n452 14.167
R358 GND.n414 GND.n413 13.653
R359 GND.n419 GND.n416 13.653
R360 GND.n422 GND.n421 13.653
R361 GND.n425 GND.n424 13.653
R362 GND.n428 GND.n427 13.653
R363 GND.n431 GND.n430 13.653
R364 GND.n434 GND.n433 13.653
R365 GND.n437 GND.n436 13.653
R366 GND.n440 GND.n439 13.653
R367 GND.n443 GND.n442 13.653
R368 GND.n446 GND.n445 13.653
R369 GND.n453 GND.n448 13.653
R370 GND.n456 GND.n455 13.653
R371 GND.n461 GND.n458 13.653
R372 GND.n464 GND.n463 13.653
R373 GND.n467 GND.n466 13.653
R374 GND.n470 GND.n469 13.653
R375 GND.n473 GND.n472 13.653
R376 GND.n476 GND.n475 13.653
R377 GND.n479 GND.n478 13.653
R378 GND.n482 GND.n481 13.653
R379 GND.n485 GND.n484 13.653
R380 GND.n488 GND.n487 13.653
R381 GND.n495 GND.n490 13.653
R382 GND.n498 GND.n497 13.653
R383 GND.n506 GND.n505 13.653
R384 GND.n509 GND.n508 13.653
R385 GND.n512 GND.n511 13.653
R386 GND.n515 GND.n514 13.653
R387 GND.n518 GND.n517 13.653
R388 GND.n521 GND.n520 13.653
R389 GND.n528 GND.n523 13.653
R390 GND.n531 GND.n530 13.653
R391 GND.n536 GND.n533 13.653
R392 GND.n539 GND.n538 13.653
R393 GND.n542 GND.n541 13.653
R394 GND.n545 GND.n544 13.653
R395 GND.n548 GND.n547 13.653
R396 GND.n551 GND.n550 13.653
R397 GND.n554 GND.n553 13.653
R398 GND.n557 GND.n556 13.653
R399 GND.n560 GND.n559 13.653
R400 GND.n563 GND.n562 13.653
R401 GND.n570 GND.n565 13.653
R402 GND.n573 GND.n572 13.653
R403 GND.n578 GND.n575 13.653
R404 GND.n581 GND.n580 13.653
R405 GND.n584 GND.n583 13.653
R406 GND.n587 GND.n586 13.653
R407 GND.n590 GND.n589 13.653
R408 GND.n593 GND.n592 13.653
R409 GND.n596 GND.n595 13.653
R410 GND.n599 GND.n598 13.653
R411 GND.n602 GND.n601 13.653
R412 GND.n605 GND.n604 13.653
R413 GND.n612 GND.n607 13.653
R414 GND.n615 GND.n614 13.653
R415 GND.n620 GND.n619 13.653
R416 GND.n623 GND.n622 13.653
R417 GND.n626 GND.n625 13.653
R418 GND.n629 GND.n628 13.653
R419 GND.n632 GND.n631 13.653
R420 GND.n635 GND.n634 13.653
R421 GND.n642 GND.n637 13.653
R422 GND.n645 GND.n644 13.653
R423 GND.n650 GND.n647 13.653
R424 GND.n653 GND.n652 13.653
R425 GND.n656 GND.n655 13.653
R426 GND.n659 GND.n658 13.653
R427 GND.n662 GND.n661 13.653
R428 GND.n665 GND.n664 13.653
R429 GND.n668 GND.n667 13.653
R430 GND.n671 GND.n670 13.653
R431 GND.n674 GND.n673 13.653
R432 GND.n677 GND.n676 13.653
R433 GND.n684 GND.n679 13.653
R434 GND.n687 GND.n686 13.653
R435 GND.n692 GND.n689 13.653
R436 GND.n695 GND.n694 13.653
R437 GND.n698 GND.n697 13.653
R438 GND.n701 GND.n700 13.653
R439 GND.n704 GND.n703 13.653
R440 GND.n707 GND.n706 13.653
R441 GND.n710 GND.n709 13.653
R442 GND.n713 GND.n712 13.653
R443 GND.n716 GND.n715 13.653
R444 GND.n719 GND.n718 13.653
R445 GND.n726 GND.n721 13.653
R446 GND.n729 GND.n728 13.653
R447 GND.n734 GND.n733 13.653
R448 GND.n737 GND.n736 13.653
R449 GND.n740 GND.n739 13.653
R450 GND.n743 GND.n742 13.653
R451 GND.n746 GND.n745 13.653
R452 GND.n749 GND.n748 13.653
R453 GND.n756 GND.n751 13.653
R454 GND.n759 GND.n758 13.653
R455 GND.n764 GND.n761 13.653
R456 GND.n767 GND.n766 13.653
R457 GND.n770 GND.n769 13.653
R458 GND.n773 GND.n772 13.653
R459 GND.n776 GND.n775 13.653
R460 GND.n779 GND.n778 13.653
R461 GND.n782 GND.n781 13.653
R462 GND.n785 GND.n784 13.653
R463 GND.n788 GND.n787 13.653
R464 GND.n791 GND.n790 13.653
R465 GND.n798 GND.n793 13.653
R466 GND.n801 GND.n800 13.653
R467 GND.n806 GND.n803 13.653
R468 GND.n408 GND.n407 13.653
R469 GND.n405 GND.n404 13.653
R470 GND.n402 GND.n401 13.653
R471 GND.n399 GND.n398 13.653
R472 GND.n396 GND.n395 13.653
R473 GND.n393 GND.n392 13.653
R474 GND.n390 GND.n389 13.653
R475 GND.n387 GND.n386 13.653
R476 GND.n384 GND.n383 13.653
R477 GND.n377 GND.n376 13.653
R478 GND.n374 GND.n373 13.653
R479 GND.n371 GND.n370 13.653
R480 GND.n366 GND.n365 13.653
R481 GND.n363 GND.n362 13.653
R482 GND.n360 GND.n359 13.653
R483 GND.n357 GND.n356 13.653
R484 GND.n354 GND.n353 13.653
R485 GND.n347 GND.n346 13.653
R486 GND.n344 GND.n343 13.653
R487 GND.n341 GND.n338 13.653
R488 GND.n336 GND.n335 13.653
R489 GND.n333 GND.n332 13.653
R490 GND.n330 GND.n329 13.653
R491 GND.n327 GND.n326 13.653
R492 GND.n324 GND.n323 13.653
R493 GND.n321 GND.n320 13.653
R494 GND.n318 GND.n317 13.653
R495 GND.n315 GND.n314 13.653
R496 GND.n312 GND.n311 13.653
R497 GND.n305 GND.n304 13.653
R498 GND.n302 GND.n301 13.653
R499 GND.n299 GND.n293 13.653
R500 GND.n291 GND.n290 13.653
R501 GND.n288 GND.n287 13.653
R502 GND.n285 GND.n284 13.653
R503 GND.n282 GND.n281 13.653
R504 GND.n279 GND.n278 13.653
R505 GND.n276 GND.n275 13.653
R506 GND.n273 GND.n272 13.653
R507 GND.n270 GND.n269 13.653
R508 GND.n267 GND.n266 13.653
R509 GND.n260 GND.n259 13.653
R510 GND.n257 GND.n256 13.653
R511 GND.n254 GND.n253 13.653
R512 GND.n249 GND.n248 13.653
R513 GND.n246 GND.n245 13.653
R514 GND.n243 GND.n242 13.653
R515 GND.n240 GND.n239 13.653
R516 GND.n237 GND.n236 13.653
R517 GND.n230 GND.n229 13.653
R518 GND.n227 GND.n226 13.653
R519 GND.n224 GND.n221 13.653
R520 GND.n219 GND.n218 13.653
R521 GND.n216 GND.n215 13.653
R522 GND.n213 GND.n212 13.653
R523 GND.n210 GND.n209 13.653
R524 GND.n207 GND.n206 13.653
R525 GND.n204 GND.n203 13.653
R526 GND.n201 GND.n200 13.653
R527 GND.n198 GND.n197 13.653
R528 GND.n195 GND.n194 13.653
R529 GND.n188 GND.n187 13.653
R530 GND.n185 GND.n184 13.653
R531 GND.n182 GND.n179 13.653
R532 GND.n177 GND.n176 13.653
R533 GND.n174 GND.n173 13.653
R534 GND.n171 GND.n170 13.653
R535 GND.n168 GND.n167 13.653
R536 GND.n165 GND.n164 13.653
R537 GND.n162 GND.n161 13.653
R538 GND.n159 GND.n158 13.653
R539 GND.n156 GND.n155 13.653
R540 GND.n153 GND.n152 13.653
R541 GND.n146 GND.n145 13.653
R542 GND.n143 GND.n142 13.653
R543 GND.n140 GND.n139 13.653
R544 GND.n135 GND.n134 13.653
R545 GND.n132 GND.n131 13.653
R546 GND.n129 GND.n128 13.653
R547 GND.n126 GND.n125 13.653
R548 GND.n123 GND.n122 13.653
R549 GND.n116 GND.n115 13.653
R550 GND.n113 GND.n112 13.653
R551 GND.n110 GND.n109 13.653
R552 GND.n105 GND.n104 13.653
R553 GND.n102 GND.n101 13.653
R554 GND.n99 GND.n98 13.653
R555 GND.n96 GND.n95 13.653
R556 GND.n93 GND.n92 13.653
R557 GND.n86 GND.n85 13.653
R558 GND.n83 GND.n82 13.653
R559 GND.n80 GND.n79 13.653
R560 GND.n75 GND.n74 13.653
R561 GND.n72 GND.n71 13.653
R562 GND.n8 GND.n7 13.653
R563 GND.n16 GND.n15 13.653
R564 GND.n23 GND.n22 13.653
R565 GND.n26 GND.n25 13.653
R566 GND.n33 GND.n32 13.653
R567 GND.n36 GND.n35 13.653
R568 GND.n39 GND.n38 13.653
R569 GND.n42 GND.n41 13.653
R570 GND.n45 GND.n44 13.653
R571 GND.n50 GND.n49 13.653
R572 GND.n53 GND.n52 13.653
R573 GND.n56 GND.n55 13.653
R574 GND.n63 GND.n62 13.653
R575 GND.n66 GND.n65 13.653
R576 GND.n69 GND.n68 13.653
R577 GND.n20 GND.n19 12.837
R578 GND.n19 GND.n18 7.566
R579 GND.n31 GND.n30 7.312
R580 GND.n61 GND.n60 7.312
R581 GND.n91 GND.n90 7.312
R582 GND.n452 GND.n451 7.312
R583 GND.n494 GND.n493 7.312
R584 GND.n527 GND.n526 7.312
R585 GND.n569 GND.n568 7.312
R586 GND.n611 GND.n610 7.312
R587 GND.n641 GND.n640 7.312
R588 GND.n683 GND.n682 7.312
R589 GND.n725 GND.n724 7.312
R590 GND.n755 GND.n754 7.312
R591 GND.n797 GND.n796 7.312
R592 GND.n382 GND.n381 7.312
R593 GND.n352 GND.n351 7.312
R594 GND.n310 GND.n309 7.312
R595 GND.n265 GND.n264 7.312
R596 GND.n235 GND.n234 7.312
R597 GND.n193 GND.n192 7.312
R598 GND.n151 GND.n150 7.312
R599 GND.n121 GND.n120 7.312
R600 GND.n11 GND.n10 4.551
R601 GND.n8 GND.n6 3.935
R602 GND.n50 GND.n48 3.935
R603 GND.n80 GND.n78 3.935
R604 GND.n110 GND.n108 3.935
R605 GND.n140 GND.n138 3.935
R606 GND.n254 GND.n252 3.935
R607 GND.n371 GND.n369 3.935
R608 GND.n734 GND.n732 3.935
R609 GND.n620 GND.n618 3.935
R610 GND.n506 GND.n504 3.935
R611 GND.n23 GND.n21 3.541
R612 GND.t13 GND.n11 2.238
R613 GND.n411 GND.n410 0.596
R614 GND.n1 GND.n0 0.596
R615 GND.n13 GND.n12 0.358
R616 GND.n34 GND.n27 0.29
R617 GND.n64 GND.n57 0.29
R618 GND.n94 GND.n87 0.29
R619 GND.n124 GND.n117 0.29
R620 GND.n154 GND.n147 0.29
R621 GND.n196 GND.n189 0.29
R622 GND.n238 GND.n231 0.29
R623 GND.n268 GND.n261 0.29
R624 GND.n313 GND.n306 0.29
R625 GND.n355 GND.n348 0.29
R626 GND.n385 GND.n378 0.29
R627 GND.n799 GND.n792 0.29
R628 GND.n757 GND.n750 0.29
R629 GND.n727 GND.n720 0.29
R630 GND.n685 GND.n678 0.29
R631 GND.n643 GND.n636 0.29
R632 GND.n613 GND.n606 0.29
R633 GND.n571 GND.n564 0.29
R634 GND.n529 GND.n522 0.29
R635 GND.n496 GND.n489 0.29
R636 GND.n454 GND.n447 0.29
R637 GND.n412 GND 0.207
R638 GND.n172 GND.n169 0.197
R639 GND.n214 GND.n211 0.197
R640 GND.n286 GND.n283 0.197
R641 GND.n331 GND.n328 0.197
R642 GND.n403 GND.n400 0.197
R643 GND.n777 GND.n774 0.197
R644 GND.n705 GND.n702 0.197
R645 GND.n663 GND.n660 0.197
R646 GND.n591 GND.n588 0.197
R647 GND.n549 GND.n546 0.197
R648 GND.n474 GND.n471 0.197
R649 GND.n432 GND.n429 0.197
R650 GND.n16 GND.n14 0.196
R651 GND.n182 GND.n181 0.196
R652 GND.n224 GND.n223 0.196
R653 GND.n299 GND.n298 0.196
R654 GND.n341 GND.n340 0.196
R655 GND.n806 GND.n805 0.196
R656 GND.n764 GND.n763 0.196
R657 GND.n692 GND.n691 0.196
R658 GND.n650 GND.n649 0.196
R659 GND.n578 GND.n577 0.196
R660 GND.n536 GND.n535 0.196
R661 GND.n461 GND.n460 0.196
R662 GND.n419 GND.n418 0.196
R663 GND.n46 GND.n43 0.181
R664 GND.n76 GND.n73 0.181
R665 GND.n106 GND.n103 0.181
R666 GND.n136 GND.n133 0.181
R667 GND.n250 GND.n247 0.181
R668 GND.n367 GND.n364 0.181
R669 GND.n741 GND.n738 0.181
R670 GND.n627 GND.n624 0.181
R671 GND.n513 GND.n510 0.181
R672 GND.n17 GND.n9 0.157
R673 GND.n24 GND.n17 0.157
R674 GND.n27 GND.n24 0.145
R675 GND.n37 GND.n34 0.145
R676 GND.n40 GND.n37 0.145
R677 GND.n43 GND.n40 0.145
R678 GND.n51 GND.n46 0.145
R679 GND.n54 GND.n51 0.145
R680 GND.n57 GND.n54 0.145
R681 GND.n67 GND.n64 0.145
R682 GND.n70 GND.n67 0.145
R683 GND.n73 GND.n70 0.145
R684 GND.n81 GND.n76 0.145
R685 GND.n84 GND.n81 0.145
R686 GND.n87 GND.n84 0.145
R687 GND.n97 GND.n94 0.145
R688 GND.n100 GND.n97 0.145
R689 GND.n103 GND.n100 0.145
R690 GND.n111 GND.n106 0.145
R691 GND.n114 GND.n111 0.145
R692 GND.n117 GND.n114 0.145
R693 GND.n127 GND.n124 0.145
R694 GND.n130 GND.n127 0.145
R695 GND.n133 GND.n130 0.145
R696 GND.n141 GND.n136 0.145
R697 GND.n144 GND.n141 0.145
R698 GND.n147 GND.n144 0.145
R699 GND.n157 GND.n154 0.145
R700 GND.n160 GND.n157 0.145
R701 GND.n163 GND.n160 0.145
R702 GND.n166 GND.n163 0.145
R703 GND.n169 GND.n166 0.145
R704 GND.n175 GND.n172 0.145
R705 GND.n178 GND.n175 0.145
R706 GND.n183 GND.n178 0.145
R707 GND.n186 GND.n183 0.145
R708 GND.n189 GND.n186 0.145
R709 GND.n199 GND.n196 0.145
R710 GND.n202 GND.n199 0.145
R711 GND.n205 GND.n202 0.145
R712 GND.n208 GND.n205 0.145
R713 GND.n211 GND.n208 0.145
R714 GND.n217 GND.n214 0.145
R715 GND.n220 GND.n217 0.145
R716 GND.n225 GND.n220 0.145
R717 GND.n228 GND.n225 0.145
R718 GND.n231 GND.n228 0.145
R719 GND.n241 GND.n238 0.145
R720 GND.n244 GND.n241 0.145
R721 GND.n247 GND.n244 0.145
R722 GND.n255 GND.n250 0.145
R723 GND.n258 GND.n255 0.145
R724 GND.n261 GND.n258 0.145
R725 GND.n271 GND.n268 0.145
R726 GND.n274 GND.n271 0.145
R727 GND.n277 GND.n274 0.145
R728 GND.n280 GND.n277 0.145
R729 GND.n283 GND.n280 0.145
R730 GND.n289 GND.n286 0.145
R731 GND.n292 GND.n289 0.145
R732 GND.n300 GND.n292 0.145
R733 GND.n303 GND.n300 0.145
R734 GND.n306 GND.n303 0.145
R735 GND.n316 GND.n313 0.145
R736 GND.n319 GND.n316 0.145
R737 GND.n322 GND.n319 0.145
R738 GND.n325 GND.n322 0.145
R739 GND.n328 GND.n325 0.145
R740 GND.n334 GND.n331 0.145
R741 GND.n337 GND.n334 0.145
R742 GND.n342 GND.n337 0.145
R743 GND.n345 GND.n342 0.145
R744 GND.n348 GND.n345 0.145
R745 GND.n358 GND.n355 0.145
R746 GND.n361 GND.n358 0.145
R747 GND.n364 GND.n361 0.145
R748 GND.n372 GND.n367 0.145
R749 GND.n375 GND.n372 0.145
R750 GND.n378 GND.n375 0.145
R751 GND.n388 GND.n385 0.145
R752 GND.n391 GND.n388 0.145
R753 GND.n394 GND.n391 0.145
R754 GND.n397 GND.n394 0.145
R755 GND.n400 GND.n397 0.145
R756 GND.n406 GND.n403 0.145
R757 GND.n409 GND.n406 0.145
R758 GND.n807 GND.n802 0.145
R759 GND.n802 GND.n799 0.145
R760 GND.n792 GND.n789 0.145
R761 GND.n789 GND.n786 0.145
R762 GND.n786 GND.n783 0.145
R763 GND.n783 GND.n780 0.145
R764 GND.n780 GND.n777 0.145
R765 GND.n774 GND.n771 0.145
R766 GND.n771 GND.n768 0.145
R767 GND.n768 GND.n765 0.145
R768 GND.n765 GND.n760 0.145
R769 GND.n760 GND.n757 0.145
R770 GND.n750 GND.n747 0.145
R771 GND.n747 GND.n744 0.145
R772 GND.n744 GND.n741 0.145
R773 GND.n738 GND.n735 0.145
R774 GND.n735 GND.n730 0.145
R775 GND.n730 GND.n727 0.145
R776 GND.n720 GND.n717 0.145
R777 GND.n717 GND.n714 0.145
R778 GND.n714 GND.n711 0.145
R779 GND.n711 GND.n708 0.145
R780 GND.n708 GND.n705 0.145
R781 GND.n702 GND.n699 0.145
R782 GND.n699 GND.n696 0.145
R783 GND.n696 GND.n693 0.145
R784 GND.n693 GND.n688 0.145
R785 GND.n688 GND.n685 0.145
R786 GND.n678 GND.n675 0.145
R787 GND.n675 GND.n672 0.145
R788 GND.n672 GND.n669 0.145
R789 GND.n669 GND.n666 0.145
R790 GND.n666 GND.n663 0.145
R791 GND.n660 GND.n657 0.145
R792 GND.n657 GND.n654 0.145
R793 GND.n654 GND.n651 0.145
R794 GND.n651 GND.n646 0.145
R795 GND.n646 GND.n643 0.145
R796 GND.n636 GND.n633 0.145
R797 GND.n633 GND.n630 0.145
R798 GND.n630 GND.n627 0.145
R799 GND.n624 GND.n621 0.145
R800 GND.n621 GND.n616 0.145
R801 GND.n616 GND.n613 0.145
R802 GND.n606 GND.n603 0.145
R803 GND.n603 GND.n600 0.145
R804 GND.n600 GND.n597 0.145
R805 GND.n597 GND.n594 0.145
R806 GND.n594 GND.n591 0.145
R807 GND.n588 GND.n585 0.145
R808 GND.n585 GND.n582 0.145
R809 GND.n582 GND.n579 0.145
R810 GND.n579 GND.n574 0.145
R811 GND.n574 GND.n571 0.145
R812 GND.n564 GND.n561 0.145
R813 GND.n561 GND.n558 0.145
R814 GND.n558 GND.n555 0.145
R815 GND.n555 GND.n552 0.145
R816 GND.n552 GND.n549 0.145
R817 GND.n546 GND.n543 0.145
R818 GND.n543 GND.n540 0.145
R819 GND.n540 GND.n537 0.145
R820 GND.n537 GND.n532 0.145
R821 GND.n532 GND.n529 0.145
R822 GND.n522 GND.n519 0.145
R823 GND.n519 GND.n516 0.145
R824 GND.n516 GND.n513 0.145
R825 GND.n510 GND.n507 0.145
R826 GND.n507 GND.n499 0.145
R827 GND.n499 GND.n496 0.145
R828 GND.n489 GND.n486 0.145
R829 GND.n486 GND.n483 0.145
R830 GND.n483 GND.n480 0.145
R831 GND.n480 GND.n477 0.145
R832 GND.n477 GND.n474 0.145
R833 GND.n471 GND.n468 0.145
R834 GND.n468 GND.n465 0.145
R835 GND.n465 GND.n462 0.145
R836 GND.n462 GND.n457 0.145
R837 GND.n457 GND.n454 0.145
R838 GND.n447 GND.n444 0.145
R839 GND.n444 GND.n441 0.145
R840 GND.n441 GND.n438 0.145
R841 GND.n438 GND.n435 0.145
R842 GND.n435 GND.n432 0.145
R843 GND.n429 GND.n426 0.145
R844 GND.n426 GND.n423 0.145
R845 GND.n423 GND.n420 0.145
R846 GND.n420 GND.n415 0.145
R847 GND.n415 GND.n412 0.145
R848 GND GND.n807 0.086
R849 GND GND.n409 0.058
R850 RN.n17 RN.t21 479.223
R851 RN.n8 RN.t12 479.223
R852 RN.n0 RN.t25 479.223
R853 RN.n23 RN.t10 454.685
R854 RN.n20 RN.t14 454.685
R855 RN.n14 RN.t0 454.685
R856 RN.n11 RN.t5 454.685
R857 RN.n5 RN.t13 454.685
R858 RN.n2 RN.t15 454.685
R859 RN.n23 RN.t17 428.979
R860 RN.n20 RN.t1 428.979
R861 RN.n14 RN.t8 428.979
R862 RN.n11 RN.t19 428.979
R863 RN.n5 RN.t3 428.979
R864 RN.n2 RN.t6 428.979
R865 RN.n17 RN.t23 375.52
R866 RN.n8 RN.t24 375.52
R867 RN.n0 RN.t9 375.52
R868 RN.n24 RN.n23 178.106
R869 RN.n21 RN.n20 178.106
R870 RN.n15 RN.n14 178.106
R871 RN.n12 RN.n11 178.106
R872 RN.n6 RN.n5 178.106
R873 RN.n3 RN.n2 178.106
R874 RN.n18 RN.n17 175.429
R875 RN.n9 RN.n8 175.429
R876 RN.n1 RN.n0 175.429
R877 RN.n18 RN.t18 162.048
R878 RN.n9 RN.t4 162.048
R879 RN.n1 RN.t22 162.048
R880 RN.n24 RN.t16 158.3
R881 RN.n21 RN.t7 158.3
R882 RN.n15 RN.t2 158.3
R883 RN.n12 RN.t26 158.3
R884 RN.n6 RN.t20 158.3
R885 RN.n3 RN.t11 158.3
R886 RN.n4 RN.n1 78.675
R887 RN.n4 RN.n3 76
R888 RN.n7 RN.n6 76
R889 RN.n10 RN.n9 76
R890 RN.n13 RN.n12 76
R891 RN.n16 RN.n15 76
R892 RN.n19 RN.n18 76
R893 RN.n22 RN.n21 76
R894 RN.n25 RN.n24 76
R895 RN.n10 RN.n7 10.293
R896 RN.n19 RN.n16 10.293
R897 RN.n7 RN.n4 5.94
R898 RN.n16 RN.n13 5.94
R899 RN.n25 RN.n22 5.94
R900 RN.n13 RN.n10 2.675
R901 RN.n22 RN.n19 2.675
R902 RN.n25 RN 0.046
R903 VDD.n891 VDD.n889 144.705
R904 VDD.n972 VDD.n970 144.705
R905 VDD.n1033 VDD.n1031 144.705
R906 VDD.n1114 VDD.n1112 144.705
R907 VDD.n1195 VDD.n1193 144.705
R908 VDD.n1256 VDD.n1254 144.705
R909 VDD.n1337 VDD.n1335 144.705
R910 VDD.n1418 VDD.n1416 144.705
R911 VDD.n1479 VDD.n1477 144.705
R912 VDD.n744 VDD.n742 144.705
R913 VDD.n1560 VDD.n1558 144.705
R914 VDD.n683 VDD.n681 144.705
R915 VDD.n602 VDD.n600 144.705
R916 VDD.n521 VDD.n519 144.705
R917 VDD.n460 VDD.n458 144.705
R918 VDD.n379 VDD.n377 144.705
R919 VDD.n298 VDD.n296 144.705
R920 VDD.n237 VDD.n235 144.705
R921 VDD.n176 VDD.n174 144.705
R922 VDD.n122 VDD.n120 144.705
R923 VDD.n68 VDD.n66 144.705
R924 VDD.n26 VDD.n25 77.792
R925 VDD.n35 VDD.n34 77.792
R926 VDD.n29 VDD.n23 76.145
R927 VDD.n29 VDD.n28 76
R928 VDD.n33 VDD.n32 76
R929 VDD.n39 VDD.n38 76
R930 VDD.n43 VDD.n42 76
R931 VDD.n70 VDD.n69 76
R932 VDD.n74 VDD.n73 76
R933 VDD.n78 VDD.n77 76
R934 VDD.n82 VDD.n81 76
R935 VDD.n86 VDD.n85 76
R936 VDD.n90 VDD.n89 76
R937 VDD.n94 VDD.n93 76
R938 VDD.n98 VDD.n97 76
R939 VDD.n124 VDD.n123 76
R940 VDD.n128 VDD.n127 76
R941 VDD.n132 VDD.n131 76
R942 VDD.n136 VDD.n135 76
R943 VDD.n140 VDD.n139 76
R944 VDD.n144 VDD.n143 76
R945 VDD.n148 VDD.n147 76
R946 VDD.n152 VDD.n151 76
R947 VDD.n178 VDD.n177 76
R948 VDD.n183 VDD.n182 76
R949 VDD.n188 VDD.n187 76
R950 VDD.n194 VDD.n193 76
R951 VDD.n199 VDD.n198 76
R952 VDD.n204 VDD.n203 76
R953 VDD.n209 VDD.n208 76
R954 VDD.n213 VDD.n212 76
R955 VDD.n239 VDD.n238 76
R956 VDD.n244 VDD.n243 76
R957 VDD.n249 VDD.n248 76
R958 VDD.n255 VDD.n254 76
R959 VDD.n260 VDD.n259 76
R960 VDD.n265 VDD.n264 76
R961 VDD.n270 VDD.n269 76
R962 VDD.n274 VDD.n273 76
R963 VDD.n300 VDD.n299 76
R964 VDD.n304 VDD.n303 76
R965 VDD.n308 VDD.n307 76
R966 VDD.n313 VDD.n312 76
R967 VDD.n320 VDD.n319 76
R968 VDD.n325 VDD.n324 76
R969 VDD.n330 VDD.n329 76
R970 VDD.n337 VDD.n336 76
R971 VDD.n342 VDD.n341 76
R972 VDD.n347 VDD.n346 76
R973 VDD.n351 VDD.n350 76
R974 VDD.n355 VDD.n354 76
R975 VDD.n381 VDD.n380 76
R976 VDD.n385 VDD.n384 76
R977 VDD.n389 VDD.n388 76
R978 VDD.n394 VDD.n393 76
R979 VDD.n401 VDD.n400 76
R980 VDD.n406 VDD.n405 76
R981 VDD.n411 VDD.n410 76
R982 VDD.n418 VDD.n417 76
R983 VDD.n423 VDD.n422 76
R984 VDD.n428 VDD.n427 76
R985 VDD.n432 VDD.n431 76
R986 VDD.n436 VDD.n435 76
R987 VDD.n462 VDD.n461 76
R988 VDD.n467 VDD.n466 76
R989 VDD.n472 VDD.n471 76
R990 VDD.n478 VDD.n477 76
R991 VDD.n483 VDD.n482 76
R992 VDD.n488 VDD.n487 76
R993 VDD.n493 VDD.n492 76
R994 VDD.n497 VDD.n496 76
R995 VDD.n523 VDD.n522 76
R996 VDD.n527 VDD.n526 76
R997 VDD.n531 VDD.n530 76
R998 VDD.n536 VDD.n535 76
R999 VDD.n543 VDD.n542 76
R1000 VDD.n548 VDD.n547 76
R1001 VDD.n553 VDD.n552 76
R1002 VDD.n560 VDD.n559 76
R1003 VDD.n565 VDD.n564 76
R1004 VDD.n570 VDD.n569 76
R1005 VDD.n574 VDD.n573 76
R1006 VDD.n578 VDD.n577 76
R1007 VDD.n604 VDD.n603 76
R1008 VDD.n608 VDD.n607 76
R1009 VDD.n612 VDD.n611 76
R1010 VDD.n617 VDD.n616 76
R1011 VDD.n624 VDD.n623 76
R1012 VDD.n629 VDD.n628 76
R1013 VDD.n634 VDD.n633 76
R1014 VDD.n641 VDD.n640 76
R1015 VDD.n646 VDD.n645 76
R1016 VDD.n651 VDD.n650 76
R1017 VDD.n655 VDD.n654 76
R1018 VDD.n659 VDD.n658 76
R1019 VDD.n685 VDD.n684 76
R1020 VDD.n690 VDD.n689 76
R1021 VDD.n695 VDD.n694 76
R1022 VDD.n701 VDD.n700 76
R1023 VDD.n706 VDD.n705 76
R1024 VDD.n711 VDD.n710 76
R1025 VDD.n716 VDD.n715 76
R1026 VDD.n720 VDD.n719 76
R1027 VDD.n746 VDD.n745 76
R1028 VDD.n750 VDD.n749 76
R1029 VDD.n754 VDD.n753 76
R1030 VDD.n759 VDD.n758 76
R1031 VDD.n766 VDD.n765 76
R1032 VDD.n771 VDD.n770 76
R1033 VDD.n776 VDD.n775 76
R1034 VDD.n783 VDD.n782 76
R1035 VDD.n788 VDD.n787 76
R1036 VDD.n1571 VDD.n1570 76
R1037 VDD.n1566 VDD.n1565 76
R1038 VDD.n1562 VDD.n1561 76
R1039 VDD.n1536 VDD.n1535 76
R1040 VDD.n1532 VDD.n1531 76
R1041 VDD.n1528 VDD.n1527 76
R1042 VDD.n1524 VDD.n1523 76
R1043 VDD.n1519 VDD.n1518 76
R1044 VDD.n1512 VDD.n1511 76
R1045 VDD.n1507 VDD.n1506 76
R1046 VDD.n1502 VDD.n1501 76
R1047 VDD.n1495 VDD.n1494 76
R1048 VDD.n1490 VDD.n1489 76
R1049 VDD.n1485 VDD.n1484 76
R1050 VDD.n1481 VDD.n1480 76
R1051 VDD.n1455 VDD.n1454 76
R1052 VDD.n1451 VDD.n1450 76
R1053 VDD.n1446 VDD.n1445 76
R1054 VDD.n1441 VDD.n1440 76
R1055 VDD.n1435 VDD.n1434 76
R1056 VDD.n1430 VDD.n1429 76
R1057 VDD.n1425 VDD.n1424 76
R1058 VDD.n1420 VDD.n1419 76
R1059 VDD.n1394 VDD.n1393 76
R1060 VDD.n1390 VDD.n1389 76
R1061 VDD.n1386 VDD.n1385 76
R1062 VDD.n1382 VDD.n1381 76
R1063 VDD.n1377 VDD.n1376 76
R1064 VDD.n1370 VDD.n1369 76
R1065 VDD.n1365 VDD.n1364 76
R1066 VDD.n1360 VDD.n1359 76
R1067 VDD.n1353 VDD.n1352 76
R1068 VDD.n1348 VDD.n1347 76
R1069 VDD.n1343 VDD.n1342 76
R1070 VDD.n1339 VDD.n1338 76
R1071 VDD.n1313 VDD.n1312 76
R1072 VDD.n1309 VDD.n1308 76
R1073 VDD.n1305 VDD.n1304 76
R1074 VDD.n1301 VDD.n1300 76
R1075 VDD.n1296 VDD.n1295 76
R1076 VDD.n1289 VDD.n1288 76
R1077 VDD.n1284 VDD.n1283 76
R1078 VDD.n1279 VDD.n1278 76
R1079 VDD.n1272 VDD.n1271 76
R1080 VDD.n1267 VDD.n1266 76
R1081 VDD.n1262 VDD.n1261 76
R1082 VDD.n1258 VDD.n1257 76
R1083 VDD.n1232 VDD.n1231 76
R1084 VDD.n1228 VDD.n1227 76
R1085 VDD.n1223 VDD.n1222 76
R1086 VDD.n1218 VDD.n1217 76
R1087 VDD.n1212 VDD.n1211 76
R1088 VDD.n1207 VDD.n1206 76
R1089 VDD.n1202 VDD.n1201 76
R1090 VDD.n1197 VDD.n1196 76
R1091 VDD.n1171 VDD.n1170 76
R1092 VDD.n1167 VDD.n1166 76
R1093 VDD.n1163 VDD.n1162 76
R1094 VDD.n1159 VDD.n1158 76
R1095 VDD.n1154 VDD.n1153 76
R1096 VDD.n1147 VDD.n1146 76
R1097 VDD.n1142 VDD.n1141 76
R1098 VDD.n1137 VDD.n1136 76
R1099 VDD.n1130 VDD.n1129 76
R1100 VDD.n1125 VDD.n1124 76
R1101 VDD.n1120 VDD.n1119 76
R1102 VDD.n1116 VDD.n1115 76
R1103 VDD.n1090 VDD.n1089 76
R1104 VDD.n1086 VDD.n1085 76
R1105 VDD.n1082 VDD.n1081 76
R1106 VDD.n1078 VDD.n1077 76
R1107 VDD.n1073 VDD.n1072 76
R1108 VDD.n1066 VDD.n1065 76
R1109 VDD.n1061 VDD.n1060 76
R1110 VDD.n1056 VDD.n1055 76
R1111 VDD.n1049 VDD.n1048 76
R1112 VDD.n1044 VDD.n1043 76
R1113 VDD.n1039 VDD.n1038 76
R1114 VDD.n1035 VDD.n1034 76
R1115 VDD.n1009 VDD.n1008 76
R1116 VDD.n1005 VDD.n1004 76
R1117 VDD.n1000 VDD.n999 76
R1118 VDD.n995 VDD.n994 76
R1119 VDD.n989 VDD.n988 76
R1120 VDD.n984 VDD.n983 76
R1121 VDD.n979 VDD.n978 76
R1122 VDD.n974 VDD.n973 76
R1123 VDD.n948 VDD.n947 76
R1124 VDD.n944 VDD.n943 76
R1125 VDD.n940 VDD.n939 76
R1126 VDD.n936 VDD.n935 76
R1127 VDD.n931 VDD.n930 76
R1128 VDD.n924 VDD.n923 76
R1129 VDD.n919 VDD.n918 76
R1130 VDD.n914 VDD.n913 76
R1131 VDD.n907 VDD.n906 76
R1132 VDD.n902 VDD.n901 76
R1133 VDD.n897 VDD.n896 76
R1134 VDD.n893 VDD.n892 76
R1135 VDD.n866 VDD.n865 76
R1136 VDD.n862 VDD.n861 76
R1137 VDD.n858 VDD.n857 76
R1138 VDD.n854 VDD.n853 76
R1139 VDD.n849 VDD.n848 76
R1140 VDD.n842 VDD.n841 76
R1141 VDD.n837 VDD.n836 76
R1142 VDD.n832 VDD.n831 76
R1143 VDD.n825 VDD.n824 76
R1144 VDD.n820 VDD.n819 76
R1145 VDD.n815 VDD.n814 76
R1146 VDD.n811 VDD.n810 76
R1147 VDD.n310 VDD.n309 64.064
R1148 VDD.n391 VDD.n390 64.064
R1149 VDD.n533 VDD.n532 64.064
R1150 VDD.n614 VDD.n613 64.064
R1151 VDD.n756 VDD.n755 64.064
R1152 VDD.n1521 VDD.n1520 64.064
R1153 VDD.n1379 VDD.n1378 64.064
R1154 VDD.n1298 VDD.n1297 64.064
R1155 VDD.n1156 VDD.n1155 64.064
R1156 VDD.n1075 VDD.n1074 64.064
R1157 VDD.n933 VDD.n932 64.064
R1158 VDD.n851 VDD.n850 64.064
R1159 VDD.n339 VDD.n338 59.488
R1160 VDD.n420 VDD.n419 59.488
R1161 VDD.n562 VDD.n561 59.488
R1162 VDD.n643 VDD.n642 59.488
R1163 VDD.n785 VDD.n784 59.488
R1164 VDD.n1492 VDD.n1491 59.488
R1165 VDD.n1350 VDD.n1349 59.488
R1166 VDD.n1269 VDD.n1268 59.488
R1167 VDD.n1127 VDD.n1126 59.488
R1168 VDD.n1046 VDD.n1045 59.488
R1169 VDD.n904 VDD.n903 59.488
R1170 VDD.n822 VDD.n821 59.488
R1171 VDD.n205 VDD.t16 55.465
R1172 VDD.n179 VDD.t9 55.465
R1173 VDD.n816 VDD.t94 55.106
R1174 VDD.n898 VDD.t72 55.106
R1175 VDD.n975 VDD.t81 55.106
R1176 VDD.n1040 VDD.t63 55.106
R1177 VDD.n1121 VDD.t98 55.106
R1178 VDD.n1198 VDD.t13 55.106
R1179 VDD.n1263 VDD.t11 55.106
R1180 VDD.n1344 VDD.t92 55.106
R1181 VDD.n1421 VDD.t24 55.106
R1182 VDD.n1486 VDD.t97 55.106
R1183 VDD.n1567 VDD.t5 55.106
R1184 VDD.n712 VDD.t62 55.106
R1185 VDD.n647 VDD.t88 55.106
R1186 VDD.n566 VDD.t80 55.106
R1187 VDD.n489 VDD.t3 55.106
R1188 VDD.n424 VDD.t78 55.106
R1189 VDD.n343 VDD.t70 55.106
R1190 VDD.n266 VDD.t10 55.106
R1191 VDD.n37 VDD.t101 55.106
R1192 VDD.n24 VDD.t91 55.106
R1193 VDD.n857 VDD.t52 55.106
R1194 VDD.n939 VDD.t40 55.106
R1195 VDD.n1081 VDD.t39 55.106
R1196 VDD.n1162 VDD.t66 55.106
R1197 VDD.n1304 VDD.t25 55.106
R1198 VDD.n1385 VDD.t36 55.106
R1199 VDD.n1527 VDD.t41 55.106
R1200 VDD.n753 VDD.t21 55.106
R1201 VDD.n611 VDD.t0 55.106
R1202 VDD.n530 VDD.t31 55.106
R1203 VDD.n388 VDD.t32 55.106
R1204 VDD.n307 VDD.t64 55.106
R1205 VDD.n1001 VDD.t7 55.106
R1206 VDD.n1224 VDD.t23 55.106
R1207 VDD.n1447 VDD.t76 55.106
R1208 VDD.n686 VDD.t71 55.106
R1209 VDD.n463 VDD.t59 55.106
R1210 VDD.n240 VDD.t6 55.106
R1211 VDD.n190 VDD.n189 41.183
R1212 VDD.n827 VDD.n826 40.824
R1213 VDD.n847 VDD.n846 40.824
R1214 VDD.n909 VDD.n908 40.824
R1215 VDD.n929 VDD.n928 40.824
R1216 VDD.n991 VDD.n990 40.824
R1217 VDD.n1051 VDD.n1050 40.824
R1218 VDD.n1071 VDD.n1070 40.824
R1219 VDD.n1132 VDD.n1131 40.824
R1220 VDD.n1152 VDD.n1151 40.824
R1221 VDD.n1214 VDD.n1213 40.824
R1222 VDD.n1274 VDD.n1273 40.824
R1223 VDD.n1294 VDD.n1293 40.824
R1224 VDD.n1355 VDD.n1354 40.824
R1225 VDD.n1375 VDD.n1374 40.824
R1226 VDD.n1437 VDD.n1436 40.824
R1227 VDD.n1497 VDD.n1496 40.824
R1228 VDD.n1517 VDD.n1516 40.824
R1229 VDD.n778 VDD.n777 40.824
R1230 VDD.n764 VDD.n763 40.824
R1231 VDD.n697 VDD.n696 40.824
R1232 VDD.n636 VDD.n635 40.824
R1233 VDD.n622 VDD.n621 40.824
R1234 VDD.n555 VDD.n554 40.824
R1235 VDD.n541 VDD.n540 40.824
R1236 VDD.n474 VDD.n473 40.824
R1237 VDD.n413 VDD.n412 40.824
R1238 VDD.n399 VDD.n398 40.824
R1239 VDD.n332 VDD.n331 40.824
R1240 VDD.n318 VDD.n317 40.824
R1241 VDD.n251 VDD.n250 40.824
R1242 VDD.n953 VDD.n952 36.774
R1243 VDD.n1014 VDD.n1013 36.774
R1244 VDD.n1095 VDD.n1094 36.774
R1245 VDD.n1176 VDD.n1175 36.774
R1246 VDD.n1237 VDD.n1236 36.774
R1247 VDD.n1318 VDD.n1317 36.774
R1248 VDD.n1399 VDD.n1398 36.774
R1249 VDD.n1460 VDD.n1459 36.774
R1250 VDD.n1541 VDD.n1540 36.774
R1251 VDD.n725 VDD.n724 36.774
R1252 VDD.n664 VDD.n663 36.774
R1253 VDD.n583 VDD.n582 36.774
R1254 VDD.n502 VDD.n501 36.774
R1255 VDD.n441 VDD.n440 36.774
R1256 VDD.n360 VDD.n359 36.774
R1257 VDD.n279 VDD.n278 36.774
R1258 VDD.n218 VDD.n217 36.774
R1259 VDD.n157 VDD.n156 36.774
R1260 VDD.n103 VDD.n102 36.774
R1261 VDD.n48 VDD.n47 36.774
R1262 VDD.n882 VDD.n881 36.774
R1263 VDD.n185 VDD.n184 36.608
R1264 VDD.n246 VDD.n245 36.608
R1265 VDD.n469 VDD.n468 36.608
R1266 VDD.n692 VDD.n691 36.608
R1267 VDD.n1443 VDD.n1442 36.608
R1268 VDD.n1220 VDD.n1219 36.608
R1269 VDD.n997 VDD.n996 36.608
R1270 VDD.n201 VDD.n200 32.032
R1271 VDD.n262 VDD.n261 32.032
R1272 VDD.n485 VDD.n484 32.032
R1273 VDD.n708 VDD.n707 32.032
R1274 VDD.n1427 VDD.n1426 32.032
R1275 VDD.n1204 VDD.n1203 32.032
R1276 VDD.n981 VDD.n980 32.032
R1277 VDD.n315 VDD.n314 27.456
R1278 VDD.n396 VDD.n395 27.456
R1279 VDD.n538 VDD.n537 27.456
R1280 VDD.n619 VDD.n618 27.456
R1281 VDD.n761 VDD.n760 27.456
R1282 VDD.n1514 VDD.n1513 27.456
R1283 VDD.n1372 VDD.n1371 27.456
R1284 VDD.n1291 VDD.n1290 27.456
R1285 VDD.n1149 VDD.n1148 27.456
R1286 VDD.n1068 VDD.n1067 27.456
R1287 VDD.n926 VDD.n925 27.456
R1288 VDD.n844 VDD.n843 27.456
R1289 VDD.n334 VDD.n333 22.88
R1290 VDD.n415 VDD.n414 22.88
R1291 VDD.n557 VDD.n556 22.88
R1292 VDD.n638 VDD.n637 22.88
R1293 VDD.n780 VDD.n779 22.88
R1294 VDD.n1499 VDD.n1498 22.88
R1295 VDD.n1357 VDD.n1356 22.88
R1296 VDD.n1276 VDD.n1275 22.88
R1297 VDD.n1134 VDD.n1133 22.88
R1298 VDD.n1053 VDD.n1052 22.88
R1299 VDD.n911 VDD.n910 22.88
R1300 VDD.n829 VDD.n828 22.88
R1301 VDD.n810 VDD.n807 21.841
R1302 VDD.n23 VDD.n20 21.841
R1303 VDD.n826 VDD.t55 14.282
R1304 VDD.n826 VDD.t8 14.282
R1305 VDD.n846 VDD.t51 14.282
R1306 VDD.n846 VDD.t54 14.282
R1307 VDD.n908 VDD.t17 14.282
R1308 VDD.n908 VDD.t20 14.282
R1309 VDD.n928 VDD.t34 14.282
R1310 VDD.n928 VDD.t53 14.282
R1311 VDD.n990 VDD.t73 14.282
R1312 VDD.n990 VDD.t82 14.282
R1313 VDD.n1050 VDD.t90 14.282
R1314 VDD.n1050 VDD.t86 14.282
R1315 VDD.n1070 VDD.t37 14.282
R1316 VDD.n1070 VDD.t28 14.282
R1317 VDD.n1131 VDD.t45 14.282
R1318 VDD.n1131 VDD.t68 14.282
R1319 VDD.n1151 VDD.t12 14.282
R1320 VDD.n1151 VDD.t38 14.282
R1321 VDD.n1213 VDD.t93 14.282
R1322 VDD.n1213 VDD.t84 14.282
R1323 VDD.n1273 VDD.t95 14.282
R1324 VDD.n1273 VDD.t67 14.282
R1325 VDD.n1293 VDD.t79 14.282
R1326 VDD.n1293 VDD.t29 14.282
R1327 VDD.n1354 VDD.t48 14.282
R1328 VDD.n1354 VDD.t100 14.282
R1329 VDD.n1374 VDD.t35 14.282
R1330 VDD.n1374 VDD.t49 14.282
R1331 VDD.n1436 VDD.t75 14.282
R1332 VDD.n1436 VDD.t99 14.282
R1333 VDD.n1496 VDD.t85 14.282
R1334 VDD.n1496 VDD.t77 14.282
R1335 VDD.n1516 VDD.t43 14.282
R1336 VDD.n1516 VDD.t27 14.282
R1337 VDD.n777 VDD.t42 14.282
R1338 VDD.n777 VDD.t57 14.282
R1339 VDD.n763 VDD.t22 14.282
R1340 VDD.n763 VDD.t44 14.282
R1341 VDD.n696 VDD.t96 14.282
R1342 VDD.n696 VDD.t50 14.282
R1343 VDD.n635 VDD.t58 14.282
R1344 VDD.n635 VDD.t60 14.282
R1345 VDD.n621 VDD.t1 14.282
R1346 VDD.n621 VDD.t4 14.282
R1347 VDD.n554 VDD.t18 14.282
R1348 VDD.n554 VDD.t69 14.282
R1349 VDD.n540 VDD.t30 14.282
R1350 VDD.n540 VDD.t19 14.282
R1351 VDD.n473 VDD.t89 14.282
R1352 VDD.n473 VDD.t2 14.282
R1353 VDD.n412 VDD.t56 14.282
R1354 VDD.n412 VDD.t14 14.282
R1355 VDD.n398 VDD.t47 14.282
R1356 VDD.n398 VDD.t87 14.282
R1357 VDD.n331 VDD.t33 14.282
R1358 VDD.n331 VDD.t15 14.282
R1359 VDD.n317 VDD.t74 14.282
R1360 VDD.n317 VDD.t46 14.282
R1361 VDD.n250 VDD.t61 14.282
R1362 VDD.n250 VDD.t65 14.282
R1363 VDD.n189 VDD.t83 14.282
R1364 VDD.n189 VDD.t26 14.282
R1365 VDD.n807 VDD.n790 14.167
R1366 VDD.n790 VDD.n789 14.167
R1367 VDD.n968 VDD.n950 14.167
R1368 VDD.n950 VDD.n949 14.167
R1369 VDD.n1029 VDD.n1011 14.167
R1370 VDD.n1011 VDD.n1010 14.167
R1371 VDD.n1110 VDD.n1092 14.167
R1372 VDD.n1092 VDD.n1091 14.167
R1373 VDD.n1191 VDD.n1173 14.167
R1374 VDD.n1173 VDD.n1172 14.167
R1375 VDD.n1252 VDD.n1234 14.167
R1376 VDD.n1234 VDD.n1233 14.167
R1377 VDD.n1333 VDD.n1315 14.167
R1378 VDD.n1315 VDD.n1314 14.167
R1379 VDD.n1414 VDD.n1396 14.167
R1380 VDD.n1396 VDD.n1395 14.167
R1381 VDD.n1475 VDD.n1457 14.167
R1382 VDD.n1457 VDD.n1456 14.167
R1383 VDD.n1556 VDD.n1538 14.167
R1384 VDD.n1538 VDD.n1537 14.167
R1385 VDD.n740 VDD.n722 14.167
R1386 VDD.n722 VDD.n721 14.167
R1387 VDD.n679 VDD.n661 14.167
R1388 VDD.n661 VDD.n660 14.167
R1389 VDD.n598 VDD.n580 14.167
R1390 VDD.n580 VDD.n579 14.167
R1391 VDD.n517 VDD.n499 14.167
R1392 VDD.n499 VDD.n498 14.167
R1393 VDD.n456 VDD.n438 14.167
R1394 VDD.n438 VDD.n437 14.167
R1395 VDD.n375 VDD.n357 14.167
R1396 VDD.n357 VDD.n356 14.167
R1397 VDD.n294 VDD.n276 14.167
R1398 VDD.n276 VDD.n275 14.167
R1399 VDD.n233 VDD.n215 14.167
R1400 VDD.n215 VDD.n214 14.167
R1401 VDD.n172 VDD.n154 14.167
R1402 VDD.n154 VDD.n153 14.167
R1403 VDD.n118 VDD.n100 14.167
R1404 VDD.n100 VDD.n99 14.167
R1405 VDD.n64 VDD.n45 14.167
R1406 VDD.n45 VDD.n44 14.167
R1407 VDD.n887 VDD.n868 14.167
R1408 VDD.n868 VDD.n867 14.167
R1409 VDD.n20 VDD.n19 14.167
R1410 VDD.n19 VDD.n17 14.167
R1411 VDD.n69 VDD.n65 14.167
R1412 VDD.n123 VDD.n119 14.167
R1413 VDD.n177 VDD.n173 14.167
R1414 VDD.n238 VDD.n234 14.167
R1415 VDD.n299 VDD.n295 14.167
R1416 VDD.n380 VDD.n376 14.167
R1417 VDD.n461 VDD.n457 14.167
R1418 VDD.n522 VDD.n518 14.167
R1419 VDD.n603 VDD.n599 14.167
R1420 VDD.n684 VDD.n680 14.167
R1421 VDD.n745 VDD.n741 14.167
R1422 VDD.n1561 VDD.n1557 14.167
R1423 VDD.n1480 VDD.n1476 14.167
R1424 VDD.n1419 VDD.n1415 14.167
R1425 VDD.n1338 VDD.n1334 14.167
R1426 VDD.n1257 VDD.n1253 14.167
R1427 VDD.n1196 VDD.n1192 14.167
R1428 VDD.n1115 VDD.n1111 14.167
R1429 VDD.n1034 VDD.n1030 14.167
R1430 VDD.n973 VDD.n969 14.167
R1431 VDD.n892 VDD.n888 14.167
R1432 VDD.n327 VDD.n326 13.728
R1433 VDD.n408 VDD.n407 13.728
R1434 VDD.n550 VDD.n549 13.728
R1435 VDD.n631 VDD.n630 13.728
R1436 VDD.n773 VDD.n772 13.728
R1437 VDD.n1504 VDD.n1503 13.728
R1438 VDD.n1362 VDD.n1361 13.728
R1439 VDD.n1281 VDD.n1280 13.728
R1440 VDD.n1139 VDD.n1138 13.728
R1441 VDD.n1058 VDD.n1057 13.728
R1442 VDD.n916 VDD.n915 13.728
R1443 VDD.n834 VDD.n833 13.728
R1444 VDD.n23 VDD.n22 13.653
R1445 VDD.n22 VDD.n21 13.653
R1446 VDD.n28 VDD.n27 13.653
R1447 VDD.n27 VDD.n26 13.653
R1448 VDD.n32 VDD.n31 13.653
R1449 VDD.n31 VDD.n30 13.653
R1450 VDD.n38 VDD.n36 13.653
R1451 VDD.n36 VDD.n35 13.653
R1452 VDD.n42 VDD.n41 13.653
R1453 VDD.n41 VDD.n40 13.653
R1454 VDD.n69 VDD.n68 13.653
R1455 VDD.n68 VDD.n67 13.653
R1456 VDD.n73 VDD.n72 13.653
R1457 VDD.n72 VDD.n71 13.653
R1458 VDD.n77 VDD.n76 13.653
R1459 VDD.n76 VDD.n75 13.653
R1460 VDD.n81 VDD.n80 13.653
R1461 VDD.n80 VDD.n79 13.653
R1462 VDD.n85 VDD.n84 13.653
R1463 VDD.n84 VDD.n83 13.653
R1464 VDD.n89 VDD.n88 13.653
R1465 VDD.n88 VDD.n87 13.653
R1466 VDD.n93 VDD.n92 13.653
R1467 VDD.n92 VDD.n91 13.653
R1468 VDD.n97 VDD.n96 13.653
R1469 VDD.n96 VDD.n95 13.653
R1470 VDD.n123 VDD.n122 13.653
R1471 VDD.n122 VDD.n121 13.653
R1472 VDD.n127 VDD.n126 13.653
R1473 VDD.n126 VDD.n125 13.653
R1474 VDD.n131 VDD.n130 13.653
R1475 VDD.n130 VDD.n129 13.653
R1476 VDD.n135 VDD.n134 13.653
R1477 VDD.n134 VDD.n133 13.653
R1478 VDD.n139 VDD.n138 13.653
R1479 VDD.n138 VDD.n137 13.653
R1480 VDD.n143 VDD.n142 13.653
R1481 VDD.n142 VDD.n141 13.653
R1482 VDD.n147 VDD.n146 13.653
R1483 VDD.n146 VDD.n145 13.653
R1484 VDD.n151 VDD.n150 13.653
R1485 VDD.n150 VDD.n149 13.653
R1486 VDD.n177 VDD.n176 13.653
R1487 VDD.n176 VDD.n175 13.653
R1488 VDD.n182 VDD.n181 13.653
R1489 VDD.n181 VDD.n180 13.653
R1490 VDD.n187 VDD.n186 13.653
R1491 VDD.n186 VDD.n185 13.653
R1492 VDD.n193 VDD.n192 13.653
R1493 VDD.n192 VDD.n191 13.653
R1494 VDD.n198 VDD.n197 13.653
R1495 VDD.n197 VDD.n196 13.653
R1496 VDD.n203 VDD.n202 13.653
R1497 VDD.n202 VDD.n201 13.653
R1498 VDD.n208 VDD.n207 13.653
R1499 VDD.n207 VDD.n206 13.653
R1500 VDD.n212 VDD.n211 13.653
R1501 VDD.n211 VDD.n210 13.653
R1502 VDD.n238 VDD.n237 13.653
R1503 VDD.n237 VDD.n236 13.653
R1504 VDD.n243 VDD.n242 13.653
R1505 VDD.n242 VDD.n241 13.653
R1506 VDD.n248 VDD.n247 13.653
R1507 VDD.n247 VDD.n246 13.653
R1508 VDD.n254 VDD.n253 13.653
R1509 VDD.n253 VDD.n252 13.653
R1510 VDD.n259 VDD.n258 13.653
R1511 VDD.n258 VDD.n257 13.653
R1512 VDD.n264 VDD.n263 13.653
R1513 VDD.n263 VDD.n262 13.653
R1514 VDD.n269 VDD.n268 13.653
R1515 VDD.n268 VDD.n267 13.653
R1516 VDD.n273 VDD.n272 13.653
R1517 VDD.n272 VDD.n271 13.653
R1518 VDD.n299 VDD.n298 13.653
R1519 VDD.n298 VDD.n297 13.653
R1520 VDD.n303 VDD.n302 13.653
R1521 VDD.n302 VDD.n301 13.653
R1522 VDD.n307 VDD.n306 13.653
R1523 VDD.n306 VDD.n305 13.653
R1524 VDD.n312 VDD.n311 13.653
R1525 VDD.n311 VDD.n310 13.653
R1526 VDD.n319 VDD.n316 13.653
R1527 VDD.n316 VDD.n315 13.653
R1528 VDD.n324 VDD.n323 13.653
R1529 VDD.n323 VDD.n322 13.653
R1530 VDD.n329 VDD.n328 13.653
R1531 VDD.n328 VDD.n327 13.653
R1532 VDD.n336 VDD.n335 13.653
R1533 VDD.n335 VDD.n334 13.653
R1534 VDD.n341 VDD.n340 13.653
R1535 VDD.n340 VDD.n339 13.653
R1536 VDD.n346 VDD.n345 13.653
R1537 VDD.n345 VDD.n344 13.653
R1538 VDD.n350 VDD.n349 13.653
R1539 VDD.n349 VDD.n348 13.653
R1540 VDD.n354 VDD.n353 13.653
R1541 VDD.n353 VDD.n352 13.653
R1542 VDD.n380 VDD.n379 13.653
R1543 VDD.n379 VDD.n378 13.653
R1544 VDD.n384 VDD.n383 13.653
R1545 VDD.n383 VDD.n382 13.653
R1546 VDD.n388 VDD.n387 13.653
R1547 VDD.n387 VDD.n386 13.653
R1548 VDD.n393 VDD.n392 13.653
R1549 VDD.n392 VDD.n391 13.653
R1550 VDD.n400 VDD.n397 13.653
R1551 VDD.n397 VDD.n396 13.653
R1552 VDD.n405 VDD.n404 13.653
R1553 VDD.n404 VDD.n403 13.653
R1554 VDD.n410 VDD.n409 13.653
R1555 VDD.n409 VDD.n408 13.653
R1556 VDD.n417 VDD.n416 13.653
R1557 VDD.n416 VDD.n415 13.653
R1558 VDD.n422 VDD.n421 13.653
R1559 VDD.n421 VDD.n420 13.653
R1560 VDD.n427 VDD.n426 13.653
R1561 VDD.n426 VDD.n425 13.653
R1562 VDD.n431 VDD.n430 13.653
R1563 VDD.n430 VDD.n429 13.653
R1564 VDD.n435 VDD.n434 13.653
R1565 VDD.n434 VDD.n433 13.653
R1566 VDD.n461 VDD.n460 13.653
R1567 VDD.n460 VDD.n459 13.653
R1568 VDD.n466 VDD.n465 13.653
R1569 VDD.n465 VDD.n464 13.653
R1570 VDD.n471 VDD.n470 13.653
R1571 VDD.n470 VDD.n469 13.653
R1572 VDD.n477 VDD.n476 13.653
R1573 VDD.n476 VDD.n475 13.653
R1574 VDD.n482 VDD.n481 13.653
R1575 VDD.n481 VDD.n480 13.653
R1576 VDD.n487 VDD.n486 13.653
R1577 VDD.n486 VDD.n485 13.653
R1578 VDD.n492 VDD.n491 13.653
R1579 VDD.n491 VDD.n490 13.653
R1580 VDD.n496 VDD.n495 13.653
R1581 VDD.n495 VDD.n494 13.653
R1582 VDD.n522 VDD.n521 13.653
R1583 VDD.n521 VDD.n520 13.653
R1584 VDD.n526 VDD.n525 13.653
R1585 VDD.n525 VDD.n524 13.653
R1586 VDD.n530 VDD.n529 13.653
R1587 VDD.n529 VDD.n528 13.653
R1588 VDD.n535 VDD.n534 13.653
R1589 VDD.n534 VDD.n533 13.653
R1590 VDD.n542 VDD.n539 13.653
R1591 VDD.n539 VDD.n538 13.653
R1592 VDD.n547 VDD.n546 13.653
R1593 VDD.n546 VDD.n545 13.653
R1594 VDD.n552 VDD.n551 13.653
R1595 VDD.n551 VDD.n550 13.653
R1596 VDD.n559 VDD.n558 13.653
R1597 VDD.n558 VDD.n557 13.653
R1598 VDD.n564 VDD.n563 13.653
R1599 VDD.n563 VDD.n562 13.653
R1600 VDD.n569 VDD.n568 13.653
R1601 VDD.n568 VDD.n567 13.653
R1602 VDD.n573 VDD.n572 13.653
R1603 VDD.n572 VDD.n571 13.653
R1604 VDD.n577 VDD.n576 13.653
R1605 VDD.n576 VDD.n575 13.653
R1606 VDD.n603 VDD.n602 13.653
R1607 VDD.n602 VDD.n601 13.653
R1608 VDD.n607 VDD.n606 13.653
R1609 VDD.n606 VDD.n605 13.653
R1610 VDD.n611 VDD.n610 13.653
R1611 VDD.n610 VDD.n609 13.653
R1612 VDD.n616 VDD.n615 13.653
R1613 VDD.n615 VDD.n614 13.653
R1614 VDD.n623 VDD.n620 13.653
R1615 VDD.n620 VDD.n619 13.653
R1616 VDD.n628 VDD.n627 13.653
R1617 VDD.n627 VDD.n626 13.653
R1618 VDD.n633 VDD.n632 13.653
R1619 VDD.n632 VDD.n631 13.653
R1620 VDD.n640 VDD.n639 13.653
R1621 VDD.n639 VDD.n638 13.653
R1622 VDD.n645 VDD.n644 13.653
R1623 VDD.n644 VDD.n643 13.653
R1624 VDD.n650 VDD.n649 13.653
R1625 VDD.n649 VDD.n648 13.653
R1626 VDD.n654 VDD.n653 13.653
R1627 VDD.n653 VDD.n652 13.653
R1628 VDD.n658 VDD.n657 13.653
R1629 VDD.n657 VDD.n656 13.653
R1630 VDD.n684 VDD.n683 13.653
R1631 VDD.n683 VDD.n682 13.653
R1632 VDD.n689 VDD.n688 13.653
R1633 VDD.n688 VDD.n687 13.653
R1634 VDD.n694 VDD.n693 13.653
R1635 VDD.n693 VDD.n692 13.653
R1636 VDD.n700 VDD.n699 13.653
R1637 VDD.n699 VDD.n698 13.653
R1638 VDD.n705 VDD.n704 13.653
R1639 VDD.n704 VDD.n703 13.653
R1640 VDD.n710 VDD.n709 13.653
R1641 VDD.n709 VDD.n708 13.653
R1642 VDD.n715 VDD.n714 13.653
R1643 VDD.n714 VDD.n713 13.653
R1644 VDD.n719 VDD.n718 13.653
R1645 VDD.n718 VDD.n717 13.653
R1646 VDD.n745 VDD.n744 13.653
R1647 VDD.n744 VDD.n743 13.653
R1648 VDD.n749 VDD.n748 13.653
R1649 VDD.n748 VDD.n747 13.653
R1650 VDD.n753 VDD.n752 13.653
R1651 VDD.n752 VDD.n751 13.653
R1652 VDD.n758 VDD.n757 13.653
R1653 VDD.n757 VDD.n756 13.653
R1654 VDD.n765 VDD.n762 13.653
R1655 VDD.n762 VDD.n761 13.653
R1656 VDD.n770 VDD.n769 13.653
R1657 VDD.n769 VDD.n768 13.653
R1658 VDD.n775 VDD.n774 13.653
R1659 VDD.n774 VDD.n773 13.653
R1660 VDD.n782 VDD.n781 13.653
R1661 VDD.n781 VDD.n780 13.653
R1662 VDD.n787 VDD.n786 13.653
R1663 VDD.n786 VDD.n785 13.653
R1664 VDD.n1570 VDD.n1569 13.653
R1665 VDD.n1569 VDD.n1568 13.653
R1666 VDD.n1565 VDD.n1564 13.653
R1667 VDD.n1564 VDD.n1563 13.653
R1668 VDD.n1561 VDD.n1560 13.653
R1669 VDD.n1560 VDD.n1559 13.653
R1670 VDD.n1535 VDD.n1534 13.653
R1671 VDD.n1534 VDD.n1533 13.653
R1672 VDD.n1531 VDD.n1530 13.653
R1673 VDD.n1530 VDD.n1529 13.653
R1674 VDD.n1527 VDD.n1526 13.653
R1675 VDD.n1526 VDD.n1525 13.653
R1676 VDD.n1523 VDD.n1522 13.653
R1677 VDD.n1522 VDD.n1521 13.653
R1678 VDD.n1518 VDD.n1515 13.653
R1679 VDD.n1515 VDD.n1514 13.653
R1680 VDD.n1511 VDD.n1510 13.653
R1681 VDD.n1510 VDD.n1509 13.653
R1682 VDD.n1506 VDD.n1505 13.653
R1683 VDD.n1505 VDD.n1504 13.653
R1684 VDD.n1501 VDD.n1500 13.653
R1685 VDD.n1500 VDD.n1499 13.653
R1686 VDD.n1494 VDD.n1493 13.653
R1687 VDD.n1493 VDD.n1492 13.653
R1688 VDD.n1489 VDD.n1488 13.653
R1689 VDD.n1488 VDD.n1487 13.653
R1690 VDD.n1484 VDD.n1483 13.653
R1691 VDD.n1483 VDD.n1482 13.653
R1692 VDD.n1480 VDD.n1479 13.653
R1693 VDD.n1479 VDD.n1478 13.653
R1694 VDD.n1454 VDD.n1453 13.653
R1695 VDD.n1453 VDD.n1452 13.653
R1696 VDD.n1450 VDD.n1449 13.653
R1697 VDD.n1449 VDD.n1448 13.653
R1698 VDD.n1445 VDD.n1444 13.653
R1699 VDD.n1444 VDD.n1443 13.653
R1700 VDD.n1440 VDD.n1439 13.653
R1701 VDD.n1439 VDD.n1438 13.653
R1702 VDD.n1434 VDD.n1433 13.653
R1703 VDD.n1433 VDD.n1432 13.653
R1704 VDD.n1429 VDD.n1428 13.653
R1705 VDD.n1428 VDD.n1427 13.653
R1706 VDD.n1424 VDD.n1423 13.653
R1707 VDD.n1423 VDD.n1422 13.653
R1708 VDD.n1419 VDD.n1418 13.653
R1709 VDD.n1418 VDD.n1417 13.653
R1710 VDD.n1393 VDD.n1392 13.653
R1711 VDD.n1392 VDD.n1391 13.653
R1712 VDD.n1389 VDD.n1388 13.653
R1713 VDD.n1388 VDD.n1387 13.653
R1714 VDD.n1385 VDD.n1384 13.653
R1715 VDD.n1384 VDD.n1383 13.653
R1716 VDD.n1381 VDD.n1380 13.653
R1717 VDD.n1380 VDD.n1379 13.653
R1718 VDD.n1376 VDD.n1373 13.653
R1719 VDD.n1373 VDD.n1372 13.653
R1720 VDD.n1369 VDD.n1368 13.653
R1721 VDD.n1368 VDD.n1367 13.653
R1722 VDD.n1364 VDD.n1363 13.653
R1723 VDD.n1363 VDD.n1362 13.653
R1724 VDD.n1359 VDD.n1358 13.653
R1725 VDD.n1358 VDD.n1357 13.653
R1726 VDD.n1352 VDD.n1351 13.653
R1727 VDD.n1351 VDD.n1350 13.653
R1728 VDD.n1347 VDD.n1346 13.653
R1729 VDD.n1346 VDD.n1345 13.653
R1730 VDD.n1342 VDD.n1341 13.653
R1731 VDD.n1341 VDD.n1340 13.653
R1732 VDD.n1338 VDD.n1337 13.653
R1733 VDD.n1337 VDD.n1336 13.653
R1734 VDD.n1312 VDD.n1311 13.653
R1735 VDD.n1311 VDD.n1310 13.653
R1736 VDD.n1308 VDD.n1307 13.653
R1737 VDD.n1307 VDD.n1306 13.653
R1738 VDD.n1304 VDD.n1303 13.653
R1739 VDD.n1303 VDD.n1302 13.653
R1740 VDD.n1300 VDD.n1299 13.653
R1741 VDD.n1299 VDD.n1298 13.653
R1742 VDD.n1295 VDD.n1292 13.653
R1743 VDD.n1292 VDD.n1291 13.653
R1744 VDD.n1288 VDD.n1287 13.653
R1745 VDD.n1287 VDD.n1286 13.653
R1746 VDD.n1283 VDD.n1282 13.653
R1747 VDD.n1282 VDD.n1281 13.653
R1748 VDD.n1278 VDD.n1277 13.653
R1749 VDD.n1277 VDD.n1276 13.653
R1750 VDD.n1271 VDD.n1270 13.653
R1751 VDD.n1270 VDD.n1269 13.653
R1752 VDD.n1266 VDD.n1265 13.653
R1753 VDD.n1265 VDD.n1264 13.653
R1754 VDD.n1261 VDD.n1260 13.653
R1755 VDD.n1260 VDD.n1259 13.653
R1756 VDD.n1257 VDD.n1256 13.653
R1757 VDD.n1256 VDD.n1255 13.653
R1758 VDD.n1231 VDD.n1230 13.653
R1759 VDD.n1230 VDD.n1229 13.653
R1760 VDD.n1227 VDD.n1226 13.653
R1761 VDD.n1226 VDD.n1225 13.653
R1762 VDD.n1222 VDD.n1221 13.653
R1763 VDD.n1221 VDD.n1220 13.653
R1764 VDD.n1217 VDD.n1216 13.653
R1765 VDD.n1216 VDD.n1215 13.653
R1766 VDD.n1211 VDD.n1210 13.653
R1767 VDD.n1210 VDD.n1209 13.653
R1768 VDD.n1206 VDD.n1205 13.653
R1769 VDD.n1205 VDD.n1204 13.653
R1770 VDD.n1201 VDD.n1200 13.653
R1771 VDD.n1200 VDD.n1199 13.653
R1772 VDD.n1196 VDD.n1195 13.653
R1773 VDD.n1195 VDD.n1194 13.653
R1774 VDD.n1170 VDD.n1169 13.653
R1775 VDD.n1169 VDD.n1168 13.653
R1776 VDD.n1166 VDD.n1165 13.653
R1777 VDD.n1165 VDD.n1164 13.653
R1778 VDD.n1162 VDD.n1161 13.653
R1779 VDD.n1161 VDD.n1160 13.653
R1780 VDD.n1158 VDD.n1157 13.653
R1781 VDD.n1157 VDD.n1156 13.653
R1782 VDD.n1153 VDD.n1150 13.653
R1783 VDD.n1150 VDD.n1149 13.653
R1784 VDD.n1146 VDD.n1145 13.653
R1785 VDD.n1145 VDD.n1144 13.653
R1786 VDD.n1141 VDD.n1140 13.653
R1787 VDD.n1140 VDD.n1139 13.653
R1788 VDD.n1136 VDD.n1135 13.653
R1789 VDD.n1135 VDD.n1134 13.653
R1790 VDD.n1129 VDD.n1128 13.653
R1791 VDD.n1128 VDD.n1127 13.653
R1792 VDD.n1124 VDD.n1123 13.653
R1793 VDD.n1123 VDD.n1122 13.653
R1794 VDD.n1119 VDD.n1118 13.653
R1795 VDD.n1118 VDD.n1117 13.653
R1796 VDD.n1115 VDD.n1114 13.653
R1797 VDD.n1114 VDD.n1113 13.653
R1798 VDD.n1089 VDD.n1088 13.653
R1799 VDD.n1088 VDD.n1087 13.653
R1800 VDD.n1085 VDD.n1084 13.653
R1801 VDD.n1084 VDD.n1083 13.653
R1802 VDD.n1081 VDD.n1080 13.653
R1803 VDD.n1080 VDD.n1079 13.653
R1804 VDD.n1077 VDD.n1076 13.653
R1805 VDD.n1076 VDD.n1075 13.653
R1806 VDD.n1072 VDD.n1069 13.653
R1807 VDD.n1069 VDD.n1068 13.653
R1808 VDD.n1065 VDD.n1064 13.653
R1809 VDD.n1064 VDD.n1063 13.653
R1810 VDD.n1060 VDD.n1059 13.653
R1811 VDD.n1059 VDD.n1058 13.653
R1812 VDD.n1055 VDD.n1054 13.653
R1813 VDD.n1054 VDD.n1053 13.653
R1814 VDD.n1048 VDD.n1047 13.653
R1815 VDD.n1047 VDD.n1046 13.653
R1816 VDD.n1043 VDD.n1042 13.653
R1817 VDD.n1042 VDD.n1041 13.653
R1818 VDD.n1038 VDD.n1037 13.653
R1819 VDD.n1037 VDD.n1036 13.653
R1820 VDD.n1034 VDD.n1033 13.653
R1821 VDD.n1033 VDD.n1032 13.653
R1822 VDD.n1008 VDD.n1007 13.653
R1823 VDD.n1007 VDD.n1006 13.653
R1824 VDD.n1004 VDD.n1003 13.653
R1825 VDD.n1003 VDD.n1002 13.653
R1826 VDD.n999 VDD.n998 13.653
R1827 VDD.n998 VDD.n997 13.653
R1828 VDD.n994 VDD.n993 13.653
R1829 VDD.n993 VDD.n992 13.653
R1830 VDD.n988 VDD.n987 13.653
R1831 VDD.n987 VDD.n986 13.653
R1832 VDD.n983 VDD.n982 13.653
R1833 VDD.n982 VDD.n981 13.653
R1834 VDD.n978 VDD.n977 13.653
R1835 VDD.n977 VDD.n976 13.653
R1836 VDD.n973 VDD.n972 13.653
R1837 VDD.n972 VDD.n971 13.653
R1838 VDD.n947 VDD.n946 13.653
R1839 VDD.n946 VDD.n945 13.653
R1840 VDD.n943 VDD.n942 13.653
R1841 VDD.n942 VDD.n941 13.653
R1842 VDD.n939 VDD.n938 13.653
R1843 VDD.n938 VDD.n937 13.653
R1844 VDD.n935 VDD.n934 13.653
R1845 VDD.n934 VDD.n933 13.653
R1846 VDD.n930 VDD.n927 13.653
R1847 VDD.n927 VDD.n926 13.653
R1848 VDD.n923 VDD.n922 13.653
R1849 VDD.n922 VDD.n921 13.653
R1850 VDD.n918 VDD.n917 13.653
R1851 VDD.n917 VDD.n916 13.653
R1852 VDD.n913 VDD.n912 13.653
R1853 VDD.n912 VDD.n911 13.653
R1854 VDD.n906 VDD.n905 13.653
R1855 VDD.n905 VDD.n904 13.653
R1856 VDD.n901 VDD.n900 13.653
R1857 VDD.n900 VDD.n899 13.653
R1858 VDD.n896 VDD.n895 13.653
R1859 VDD.n895 VDD.n894 13.653
R1860 VDD.n892 VDD.n891 13.653
R1861 VDD.n891 VDD.n890 13.653
R1862 VDD.n865 VDD.n864 13.653
R1863 VDD.n864 VDD.n863 13.653
R1864 VDD.n861 VDD.n860 13.653
R1865 VDD.n860 VDD.n859 13.653
R1866 VDD.n857 VDD.n856 13.653
R1867 VDD.n856 VDD.n855 13.653
R1868 VDD.n853 VDD.n852 13.653
R1869 VDD.n852 VDD.n851 13.653
R1870 VDD.n848 VDD.n845 13.653
R1871 VDD.n845 VDD.n844 13.653
R1872 VDD.n841 VDD.n840 13.653
R1873 VDD.n840 VDD.n839 13.653
R1874 VDD.n836 VDD.n835 13.653
R1875 VDD.n835 VDD.n834 13.653
R1876 VDD.n831 VDD.n830 13.653
R1877 VDD.n830 VDD.n829 13.653
R1878 VDD.n824 VDD.n823 13.653
R1879 VDD.n823 VDD.n822 13.653
R1880 VDD.n819 VDD.n818 13.653
R1881 VDD.n818 VDD.n817 13.653
R1882 VDD.n814 VDD.n813 13.653
R1883 VDD.n813 VDD.n812 13.653
R1884 VDD.n810 VDD.n809 13.653
R1885 VDD.n809 VDD.n808 13.653
R1886 VDD.n4 VDD.n2 12.915
R1887 VDD.n4 VDD.n3 12.66
R1888 VDD.n13 VDD.n12 12.343
R1889 VDD.n11 VDD.n10 12.343
R1890 VDD.n7 VDD.n6 12.343
R1891 VDD.n322 VDD.n321 9.152
R1892 VDD.n403 VDD.n402 9.152
R1893 VDD.n545 VDD.n544 9.152
R1894 VDD.n626 VDD.n625 9.152
R1895 VDD.n768 VDD.n767 9.152
R1896 VDD.n1509 VDD.n1508 9.152
R1897 VDD.n1367 VDD.n1366 9.152
R1898 VDD.n1286 VDD.n1285 9.152
R1899 VDD.n1144 VDD.n1143 9.152
R1900 VDD.n1063 VDD.n1062 9.152
R1901 VDD.n921 VDD.n920 9.152
R1902 VDD.n839 VDD.n838 9.152
R1903 VDD.n193 VDD.n190 8.658
R1904 VDD.n254 VDD.n251 8.658
R1905 VDD.n477 VDD.n474 8.658
R1906 VDD.n700 VDD.n697 8.658
R1907 VDD.n1440 VDD.n1437 8.658
R1908 VDD.n1217 VDD.n1214 8.658
R1909 VDD.n994 VDD.n991 8.658
R1910 VDD.n969 VDD.n968 7.674
R1911 VDD.n1030 VDD.n1029 7.674
R1912 VDD.n1111 VDD.n1110 7.674
R1913 VDD.n1192 VDD.n1191 7.674
R1914 VDD.n1253 VDD.n1252 7.674
R1915 VDD.n1334 VDD.n1333 7.674
R1916 VDD.n1415 VDD.n1414 7.674
R1917 VDD.n1476 VDD.n1475 7.674
R1918 VDD.n1557 VDD.n1556 7.674
R1919 VDD.n741 VDD.n740 7.674
R1920 VDD.n680 VDD.n679 7.674
R1921 VDD.n599 VDD.n598 7.674
R1922 VDD.n518 VDD.n517 7.674
R1923 VDD.n457 VDD.n456 7.674
R1924 VDD.n376 VDD.n375 7.674
R1925 VDD.n295 VDD.n294 7.674
R1926 VDD.n234 VDD.n233 7.674
R1927 VDD.n173 VDD.n172 7.674
R1928 VDD.n119 VDD.n118 7.674
R1929 VDD.n65 VDD.n64 7.674
R1930 VDD.n888 VDD.n887 7.674
R1931 VDD.n59 VDD.n58 7.5
R1932 VDD.n53 VDD.n52 7.5
R1933 VDD.n55 VDD.n54 7.5
R1934 VDD.n50 VDD.n49 7.5
R1935 VDD.n64 VDD.n63 7.5
R1936 VDD.n113 VDD.n112 7.5
R1937 VDD.n107 VDD.n106 7.5
R1938 VDD.n109 VDD.n108 7.5
R1939 VDD.n115 VDD.n105 7.5
R1940 VDD.n115 VDD.n103 7.5
R1941 VDD.n118 VDD.n117 7.5
R1942 VDD.n167 VDD.n166 7.5
R1943 VDD.n161 VDD.n160 7.5
R1944 VDD.n163 VDD.n162 7.5
R1945 VDD.n169 VDD.n159 7.5
R1946 VDD.n169 VDD.n157 7.5
R1947 VDD.n172 VDD.n171 7.5
R1948 VDD.n228 VDD.n227 7.5
R1949 VDD.n222 VDD.n221 7.5
R1950 VDD.n224 VDD.n223 7.5
R1951 VDD.n230 VDD.n220 7.5
R1952 VDD.n230 VDD.n218 7.5
R1953 VDD.n233 VDD.n232 7.5
R1954 VDD.n289 VDD.n288 7.5
R1955 VDD.n283 VDD.n282 7.5
R1956 VDD.n285 VDD.n284 7.5
R1957 VDD.n291 VDD.n281 7.5
R1958 VDD.n291 VDD.n279 7.5
R1959 VDD.n294 VDD.n293 7.5
R1960 VDD.n370 VDD.n369 7.5
R1961 VDD.n364 VDD.n363 7.5
R1962 VDD.n366 VDD.n365 7.5
R1963 VDD.n372 VDD.n362 7.5
R1964 VDD.n372 VDD.n360 7.5
R1965 VDD.n375 VDD.n374 7.5
R1966 VDD.n451 VDD.n450 7.5
R1967 VDD.n445 VDD.n444 7.5
R1968 VDD.n447 VDD.n446 7.5
R1969 VDD.n453 VDD.n443 7.5
R1970 VDD.n453 VDD.n441 7.5
R1971 VDD.n456 VDD.n455 7.5
R1972 VDD.n512 VDD.n511 7.5
R1973 VDD.n506 VDD.n505 7.5
R1974 VDD.n508 VDD.n507 7.5
R1975 VDD.n514 VDD.n504 7.5
R1976 VDD.n514 VDD.n502 7.5
R1977 VDD.n517 VDD.n516 7.5
R1978 VDD.n593 VDD.n592 7.5
R1979 VDD.n587 VDD.n586 7.5
R1980 VDD.n589 VDD.n588 7.5
R1981 VDD.n595 VDD.n585 7.5
R1982 VDD.n595 VDD.n583 7.5
R1983 VDD.n598 VDD.n597 7.5
R1984 VDD.n674 VDD.n673 7.5
R1985 VDD.n668 VDD.n667 7.5
R1986 VDD.n670 VDD.n669 7.5
R1987 VDD.n676 VDD.n666 7.5
R1988 VDD.n676 VDD.n664 7.5
R1989 VDD.n679 VDD.n678 7.5
R1990 VDD.n735 VDD.n734 7.5
R1991 VDD.n729 VDD.n728 7.5
R1992 VDD.n731 VDD.n730 7.5
R1993 VDD.n737 VDD.n727 7.5
R1994 VDD.n737 VDD.n725 7.5
R1995 VDD.n740 VDD.n739 7.5
R1996 VDD.n1551 VDD.n1550 7.5
R1997 VDD.n1545 VDD.n1544 7.5
R1998 VDD.n1547 VDD.n1546 7.5
R1999 VDD.n1553 VDD.n1543 7.5
R2000 VDD.n1553 VDD.n1541 7.5
R2001 VDD.n1556 VDD.n1555 7.5
R2002 VDD.n1470 VDD.n1469 7.5
R2003 VDD.n1464 VDD.n1463 7.5
R2004 VDD.n1466 VDD.n1465 7.5
R2005 VDD.n1472 VDD.n1462 7.5
R2006 VDD.n1472 VDD.n1460 7.5
R2007 VDD.n1475 VDD.n1474 7.5
R2008 VDD.n1409 VDD.n1408 7.5
R2009 VDD.n1403 VDD.n1402 7.5
R2010 VDD.n1405 VDD.n1404 7.5
R2011 VDD.n1411 VDD.n1401 7.5
R2012 VDD.n1411 VDD.n1399 7.5
R2013 VDD.n1414 VDD.n1413 7.5
R2014 VDD.n1328 VDD.n1327 7.5
R2015 VDD.n1322 VDD.n1321 7.5
R2016 VDD.n1324 VDD.n1323 7.5
R2017 VDD.n1330 VDD.n1320 7.5
R2018 VDD.n1330 VDD.n1318 7.5
R2019 VDD.n1333 VDD.n1332 7.5
R2020 VDD.n1247 VDD.n1246 7.5
R2021 VDD.n1241 VDD.n1240 7.5
R2022 VDD.n1243 VDD.n1242 7.5
R2023 VDD.n1249 VDD.n1239 7.5
R2024 VDD.n1249 VDD.n1237 7.5
R2025 VDD.n1252 VDD.n1251 7.5
R2026 VDD.n1186 VDD.n1185 7.5
R2027 VDD.n1180 VDD.n1179 7.5
R2028 VDD.n1182 VDD.n1181 7.5
R2029 VDD.n1188 VDD.n1178 7.5
R2030 VDD.n1188 VDD.n1176 7.5
R2031 VDD.n1191 VDD.n1190 7.5
R2032 VDD.n1105 VDD.n1104 7.5
R2033 VDD.n1099 VDD.n1098 7.5
R2034 VDD.n1101 VDD.n1100 7.5
R2035 VDD.n1107 VDD.n1097 7.5
R2036 VDD.n1107 VDD.n1095 7.5
R2037 VDD.n1110 VDD.n1109 7.5
R2038 VDD.n1024 VDD.n1023 7.5
R2039 VDD.n1018 VDD.n1017 7.5
R2040 VDD.n1020 VDD.n1019 7.5
R2041 VDD.n1026 VDD.n1016 7.5
R2042 VDD.n1026 VDD.n1014 7.5
R2043 VDD.n1029 VDD.n1028 7.5
R2044 VDD.n963 VDD.n962 7.5
R2045 VDD.n957 VDD.n956 7.5
R2046 VDD.n959 VDD.n958 7.5
R2047 VDD.n965 VDD.n955 7.5
R2048 VDD.n965 VDD.n953 7.5
R2049 VDD.n968 VDD.n967 7.5
R2050 VDD.n872 VDD.n871 7.5
R2051 VDD.n875 VDD.n874 7.5
R2052 VDD.n877 VDD.n876 7.5
R2053 VDD.n880 VDD.n879 7.5
R2054 VDD.n887 VDD.n886 7.5
R2055 VDD.n802 VDD.n801 7.5
R2056 VDD.n796 VDD.n795 7.5
R2057 VDD.n798 VDD.n797 7.5
R2058 VDD.n804 VDD.n794 7.5
R2059 VDD.n804 VDD.n792 7.5
R2060 VDD.n807 VDD.n806 7.5
R2061 VDD.n20 VDD.n16 7.5
R2062 VDD.n2 VDD.n1 7.5
R2063 VDD.n6 VDD.n5 7.5
R2064 VDD.n10 VDD.n9 7.5
R2065 VDD.n19 VDD.n18 7.5
R2066 VDD.n14 VDD.n0 7.5
R2067 VDD.n51 VDD.n48 6.772
R2068 VDD.n62 VDD.n46 6.772
R2069 VDD.n60 VDD.n57 6.772
R2070 VDD.n56 VDD.n53 6.772
R2071 VDD.n116 VDD.n101 6.772
R2072 VDD.n114 VDD.n111 6.772
R2073 VDD.n110 VDD.n107 6.772
R2074 VDD.n170 VDD.n155 6.772
R2075 VDD.n168 VDD.n165 6.772
R2076 VDD.n164 VDD.n161 6.772
R2077 VDD.n231 VDD.n216 6.772
R2078 VDD.n229 VDD.n226 6.772
R2079 VDD.n225 VDD.n222 6.772
R2080 VDD.n292 VDD.n277 6.772
R2081 VDD.n290 VDD.n287 6.772
R2082 VDD.n286 VDD.n283 6.772
R2083 VDD.n373 VDD.n358 6.772
R2084 VDD.n371 VDD.n368 6.772
R2085 VDD.n367 VDD.n364 6.772
R2086 VDD.n454 VDD.n439 6.772
R2087 VDD.n452 VDD.n449 6.772
R2088 VDD.n448 VDD.n445 6.772
R2089 VDD.n515 VDD.n500 6.772
R2090 VDD.n513 VDD.n510 6.772
R2091 VDD.n509 VDD.n506 6.772
R2092 VDD.n596 VDD.n581 6.772
R2093 VDD.n594 VDD.n591 6.772
R2094 VDD.n590 VDD.n587 6.772
R2095 VDD.n677 VDD.n662 6.772
R2096 VDD.n675 VDD.n672 6.772
R2097 VDD.n671 VDD.n668 6.772
R2098 VDD.n738 VDD.n723 6.772
R2099 VDD.n736 VDD.n733 6.772
R2100 VDD.n732 VDD.n729 6.772
R2101 VDD.n1554 VDD.n1539 6.772
R2102 VDD.n1552 VDD.n1549 6.772
R2103 VDD.n1548 VDD.n1545 6.772
R2104 VDD.n1473 VDD.n1458 6.772
R2105 VDD.n1471 VDD.n1468 6.772
R2106 VDD.n1467 VDD.n1464 6.772
R2107 VDD.n1412 VDD.n1397 6.772
R2108 VDD.n1410 VDD.n1407 6.772
R2109 VDD.n1406 VDD.n1403 6.772
R2110 VDD.n1331 VDD.n1316 6.772
R2111 VDD.n1329 VDD.n1326 6.772
R2112 VDD.n1325 VDD.n1322 6.772
R2113 VDD.n1250 VDD.n1235 6.772
R2114 VDD.n1248 VDD.n1245 6.772
R2115 VDD.n1244 VDD.n1241 6.772
R2116 VDD.n1189 VDD.n1174 6.772
R2117 VDD.n1187 VDD.n1184 6.772
R2118 VDD.n1183 VDD.n1180 6.772
R2119 VDD.n1108 VDD.n1093 6.772
R2120 VDD.n1106 VDD.n1103 6.772
R2121 VDD.n1102 VDD.n1099 6.772
R2122 VDD.n1027 VDD.n1012 6.772
R2123 VDD.n1025 VDD.n1022 6.772
R2124 VDD.n1021 VDD.n1018 6.772
R2125 VDD.n966 VDD.n951 6.772
R2126 VDD.n964 VDD.n961 6.772
R2127 VDD.n960 VDD.n957 6.772
R2128 VDD.n805 VDD.n791 6.772
R2129 VDD.n803 VDD.n800 6.772
R2130 VDD.n799 VDD.n796 6.772
R2131 VDD.n51 VDD.n50 6.772
R2132 VDD.n56 VDD.n55 6.772
R2133 VDD.n60 VDD.n59 6.772
R2134 VDD.n63 VDD.n62 6.772
R2135 VDD.n110 VDD.n109 6.772
R2136 VDD.n114 VDD.n113 6.772
R2137 VDD.n117 VDD.n116 6.772
R2138 VDD.n164 VDD.n163 6.772
R2139 VDD.n168 VDD.n167 6.772
R2140 VDD.n171 VDD.n170 6.772
R2141 VDD.n225 VDD.n224 6.772
R2142 VDD.n229 VDD.n228 6.772
R2143 VDD.n232 VDD.n231 6.772
R2144 VDD.n286 VDD.n285 6.772
R2145 VDD.n290 VDD.n289 6.772
R2146 VDD.n293 VDD.n292 6.772
R2147 VDD.n367 VDD.n366 6.772
R2148 VDD.n371 VDD.n370 6.772
R2149 VDD.n374 VDD.n373 6.772
R2150 VDD.n448 VDD.n447 6.772
R2151 VDD.n452 VDD.n451 6.772
R2152 VDD.n455 VDD.n454 6.772
R2153 VDD.n509 VDD.n508 6.772
R2154 VDD.n513 VDD.n512 6.772
R2155 VDD.n516 VDD.n515 6.772
R2156 VDD.n590 VDD.n589 6.772
R2157 VDD.n594 VDD.n593 6.772
R2158 VDD.n597 VDD.n596 6.772
R2159 VDD.n671 VDD.n670 6.772
R2160 VDD.n675 VDD.n674 6.772
R2161 VDD.n678 VDD.n677 6.772
R2162 VDD.n732 VDD.n731 6.772
R2163 VDD.n736 VDD.n735 6.772
R2164 VDD.n739 VDD.n738 6.772
R2165 VDD.n1548 VDD.n1547 6.772
R2166 VDD.n1552 VDD.n1551 6.772
R2167 VDD.n1555 VDD.n1554 6.772
R2168 VDD.n1467 VDD.n1466 6.772
R2169 VDD.n1471 VDD.n1470 6.772
R2170 VDD.n1474 VDD.n1473 6.772
R2171 VDD.n1406 VDD.n1405 6.772
R2172 VDD.n1410 VDD.n1409 6.772
R2173 VDD.n1413 VDD.n1412 6.772
R2174 VDD.n1325 VDD.n1324 6.772
R2175 VDD.n1329 VDD.n1328 6.772
R2176 VDD.n1332 VDD.n1331 6.772
R2177 VDD.n1244 VDD.n1243 6.772
R2178 VDD.n1248 VDD.n1247 6.772
R2179 VDD.n1251 VDD.n1250 6.772
R2180 VDD.n1183 VDD.n1182 6.772
R2181 VDD.n1187 VDD.n1186 6.772
R2182 VDD.n1190 VDD.n1189 6.772
R2183 VDD.n1102 VDD.n1101 6.772
R2184 VDD.n1106 VDD.n1105 6.772
R2185 VDD.n1109 VDD.n1108 6.772
R2186 VDD.n1021 VDD.n1020 6.772
R2187 VDD.n1025 VDD.n1024 6.772
R2188 VDD.n1028 VDD.n1027 6.772
R2189 VDD.n960 VDD.n959 6.772
R2190 VDD.n964 VDD.n963 6.772
R2191 VDD.n967 VDD.n966 6.772
R2192 VDD.n799 VDD.n798 6.772
R2193 VDD.n803 VDD.n802 6.772
R2194 VDD.n806 VDD.n805 6.772
R2195 VDD.n886 VDD.n885 6.772
R2196 VDD.n873 VDD.n870 6.772
R2197 VDD.n878 VDD.n875 6.772
R2198 VDD.n883 VDD.n880 6.772
R2199 VDD.n883 VDD.n882 6.772
R2200 VDD.n878 VDD.n877 6.772
R2201 VDD.n873 VDD.n872 6.772
R2202 VDD.n885 VDD.n869 6.772
R2203 VDD.n336 VDD.n332 6.69
R2204 VDD.n417 VDD.n413 6.69
R2205 VDD.n559 VDD.n555 6.69
R2206 VDD.n640 VDD.n636 6.69
R2207 VDD.n782 VDD.n778 6.69
R2208 VDD.n1501 VDD.n1497 6.69
R2209 VDD.n1359 VDD.n1355 6.69
R2210 VDD.n1278 VDD.n1274 6.69
R2211 VDD.n1136 VDD.n1132 6.69
R2212 VDD.n1055 VDD.n1051 6.69
R2213 VDD.n913 VDD.n909 6.69
R2214 VDD.n831 VDD.n827 6.69
R2215 VDD.n16 VDD.n15 6.458
R2216 VDD.n319 VDD.n318 6.296
R2217 VDD.n400 VDD.n399 6.296
R2218 VDD.n542 VDD.n541 6.296
R2219 VDD.n623 VDD.n622 6.296
R2220 VDD.n765 VDD.n764 6.296
R2221 VDD.n1518 VDD.n1517 6.296
R2222 VDD.n1376 VDD.n1375 6.296
R2223 VDD.n1295 VDD.n1294 6.296
R2224 VDD.n1153 VDD.n1152 6.296
R2225 VDD.n1072 VDD.n1071 6.296
R2226 VDD.n930 VDD.n929 6.296
R2227 VDD.n848 VDD.n847 6.296
R2228 VDD.n105 VDD.n104 6.202
R2229 VDD.n159 VDD.n158 6.202
R2230 VDD.n220 VDD.n219 6.202
R2231 VDD.n281 VDD.n280 6.202
R2232 VDD.n362 VDD.n361 6.202
R2233 VDD.n443 VDD.n442 6.202
R2234 VDD.n504 VDD.n503 6.202
R2235 VDD.n585 VDD.n584 6.202
R2236 VDD.n666 VDD.n665 6.202
R2237 VDD.n727 VDD.n726 6.202
R2238 VDD.n1543 VDD.n1542 6.202
R2239 VDD.n1462 VDD.n1461 6.202
R2240 VDD.n1401 VDD.n1400 6.202
R2241 VDD.n1320 VDD.n1319 6.202
R2242 VDD.n1239 VDD.n1238 6.202
R2243 VDD.n1178 VDD.n1177 6.202
R2244 VDD.n1097 VDD.n1096 6.202
R2245 VDD.n1016 VDD.n1015 6.202
R2246 VDD.n955 VDD.n954 6.202
R2247 VDD.n794 VDD.n793 6.202
R2248 VDD.n196 VDD.n195 4.576
R2249 VDD.n257 VDD.n256 4.576
R2250 VDD.n480 VDD.n479 4.576
R2251 VDD.n703 VDD.n702 4.576
R2252 VDD.n1432 VDD.n1431 4.576
R2253 VDD.n1209 VDD.n1208 4.576
R2254 VDD.n986 VDD.n985 4.576
R2255 VDD.n208 VDD.n205 2.754
R2256 VDD.n269 VDD.n266 2.754
R2257 VDD.n492 VDD.n489 2.754
R2258 VDD.n715 VDD.n712 2.754
R2259 VDD.n1424 VDD.n1421 2.754
R2260 VDD.n1201 VDD.n1198 2.754
R2261 VDD.n978 VDD.n975 2.754
R2262 VDD.n182 VDD.n179 2.361
R2263 VDD.n243 VDD.n240 2.361
R2264 VDD.n466 VDD.n463 2.361
R2265 VDD.n689 VDD.n686 2.361
R2266 VDD.n1450 VDD.n1447 2.361
R2267 VDD.n1227 VDD.n1224 2.361
R2268 VDD.n1004 VDD.n1001 2.361
R2269 VDD.n28 VDD.n24 1.967
R2270 VDD.n38 VDD.n37 1.967
R2271 VDD.n14 VDD.n7 1.329
R2272 VDD.n14 VDD.n8 1.329
R2273 VDD.n14 VDD.n11 1.329
R2274 VDD.n14 VDD.n13 1.329
R2275 VDD.n15 VDD.n14 0.696
R2276 VDD.n14 VDD.n4 0.696
R2277 VDD.n346 VDD.n343 0.393
R2278 VDD.n427 VDD.n424 0.393
R2279 VDD.n569 VDD.n566 0.393
R2280 VDD.n650 VDD.n647 0.393
R2281 VDD.n1570 VDD.n1567 0.393
R2282 VDD.n1489 VDD.n1486 0.393
R2283 VDD.n1347 VDD.n1344 0.393
R2284 VDD.n1266 VDD.n1263 0.393
R2285 VDD.n1124 VDD.n1121 0.393
R2286 VDD.n1043 VDD.n1040 0.393
R2287 VDD.n901 VDD.n898 0.393
R2288 VDD.n819 VDD.n816 0.393
R2289 VDD.n61 VDD.n60 0.365
R2290 VDD.n61 VDD.n56 0.365
R2291 VDD.n61 VDD.n51 0.365
R2292 VDD.n62 VDD.n61 0.365
R2293 VDD.n115 VDD.n114 0.365
R2294 VDD.n115 VDD.n110 0.365
R2295 VDD.n116 VDD.n115 0.365
R2296 VDD.n169 VDD.n168 0.365
R2297 VDD.n169 VDD.n164 0.365
R2298 VDD.n170 VDD.n169 0.365
R2299 VDD.n230 VDD.n229 0.365
R2300 VDD.n230 VDD.n225 0.365
R2301 VDD.n231 VDD.n230 0.365
R2302 VDD.n291 VDD.n290 0.365
R2303 VDD.n291 VDD.n286 0.365
R2304 VDD.n292 VDD.n291 0.365
R2305 VDD.n372 VDD.n371 0.365
R2306 VDD.n372 VDD.n367 0.365
R2307 VDD.n373 VDD.n372 0.365
R2308 VDD.n453 VDD.n452 0.365
R2309 VDD.n453 VDD.n448 0.365
R2310 VDD.n454 VDD.n453 0.365
R2311 VDD.n514 VDD.n513 0.365
R2312 VDD.n514 VDD.n509 0.365
R2313 VDD.n515 VDD.n514 0.365
R2314 VDD.n595 VDD.n594 0.365
R2315 VDD.n595 VDD.n590 0.365
R2316 VDD.n596 VDD.n595 0.365
R2317 VDD.n676 VDD.n675 0.365
R2318 VDD.n676 VDD.n671 0.365
R2319 VDD.n677 VDD.n676 0.365
R2320 VDD.n737 VDD.n736 0.365
R2321 VDD.n737 VDD.n732 0.365
R2322 VDD.n738 VDD.n737 0.365
R2323 VDD.n1553 VDD.n1552 0.365
R2324 VDD.n1553 VDD.n1548 0.365
R2325 VDD.n1554 VDD.n1553 0.365
R2326 VDD.n1472 VDD.n1471 0.365
R2327 VDD.n1472 VDD.n1467 0.365
R2328 VDD.n1473 VDD.n1472 0.365
R2329 VDD.n1411 VDD.n1410 0.365
R2330 VDD.n1411 VDD.n1406 0.365
R2331 VDD.n1412 VDD.n1411 0.365
R2332 VDD.n1330 VDD.n1329 0.365
R2333 VDD.n1330 VDD.n1325 0.365
R2334 VDD.n1331 VDD.n1330 0.365
R2335 VDD.n1249 VDD.n1248 0.365
R2336 VDD.n1249 VDD.n1244 0.365
R2337 VDD.n1250 VDD.n1249 0.365
R2338 VDD.n1188 VDD.n1187 0.365
R2339 VDD.n1188 VDD.n1183 0.365
R2340 VDD.n1189 VDD.n1188 0.365
R2341 VDD.n1107 VDD.n1106 0.365
R2342 VDD.n1107 VDD.n1102 0.365
R2343 VDD.n1108 VDD.n1107 0.365
R2344 VDD.n1026 VDD.n1025 0.365
R2345 VDD.n1026 VDD.n1021 0.365
R2346 VDD.n1027 VDD.n1026 0.365
R2347 VDD.n965 VDD.n964 0.365
R2348 VDD.n965 VDD.n960 0.365
R2349 VDD.n966 VDD.n965 0.365
R2350 VDD.n804 VDD.n803 0.365
R2351 VDD.n804 VDD.n799 0.365
R2352 VDD.n805 VDD.n804 0.365
R2353 VDD.n884 VDD.n883 0.365
R2354 VDD.n884 VDD.n878 0.365
R2355 VDD.n884 VDD.n873 0.365
R2356 VDD.n885 VDD.n884 0.365
R2357 VDD.n70 VDD.n43 0.29
R2358 VDD.n124 VDD.n98 0.29
R2359 VDD.n178 VDD.n152 0.29
R2360 VDD.n239 VDD.n213 0.29
R2361 VDD.n300 VDD.n274 0.29
R2362 VDD.n381 VDD.n355 0.29
R2363 VDD.n462 VDD.n436 0.29
R2364 VDD.n523 VDD.n497 0.29
R2365 VDD.n604 VDD.n578 0.29
R2366 VDD.n685 VDD.n659 0.29
R2367 VDD.n746 VDD.n720 0.29
R2368 VDD.n1562 VDD.n1536 0.29
R2369 VDD.n1481 VDD.n1455 0.29
R2370 VDD.n1420 VDD.n1394 0.29
R2371 VDD.n1339 VDD.n1313 0.29
R2372 VDD.n1258 VDD.n1232 0.29
R2373 VDD.n1197 VDD.n1171 0.29
R2374 VDD.n1116 VDD.n1090 0.29
R2375 VDD.n1035 VDD.n1009 0.29
R2376 VDD.n974 VDD.n948 0.29
R2377 VDD.n893 VDD.n866 0.29
R2378 VDD.n811 VDD 0.207
R2379 VDD.n330 VDD.n325 0.197
R2380 VDD.n411 VDD.n406 0.197
R2381 VDD.n553 VDD.n548 0.197
R2382 VDD.n634 VDD.n629 0.197
R2383 VDD.n776 VDD.n771 0.197
R2384 VDD.n1512 VDD.n1507 0.197
R2385 VDD.n1370 VDD.n1365 0.197
R2386 VDD.n1289 VDD.n1284 0.197
R2387 VDD.n1147 VDD.n1142 0.197
R2388 VDD.n1066 VDD.n1061 0.197
R2389 VDD.n924 VDD.n919 0.197
R2390 VDD.n842 VDD.n837 0.197
R2391 VDD.n86 VDD.n82 0.181
R2392 VDD.n140 VDD.n136 0.181
R2393 VDD.n199 VDD.n194 0.181
R2394 VDD.n260 VDD.n255 0.181
R2395 VDD.n483 VDD.n478 0.181
R2396 VDD.n706 VDD.n701 0.181
R2397 VDD.n1441 VDD.n1435 0.181
R2398 VDD.n1218 VDD.n1212 0.181
R2399 VDD.n995 VDD.n989 0.181
R2400 VDD.n33 VDD.n29 0.157
R2401 VDD.n39 VDD.n33 0.157
R2402 VDD.n43 VDD.n39 0.145
R2403 VDD.n74 VDD.n70 0.145
R2404 VDD.n78 VDD.n74 0.145
R2405 VDD.n82 VDD.n78 0.145
R2406 VDD.n90 VDD.n86 0.145
R2407 VDD.n94 VDD.n90 0.145
R2408 VDD.n98 VDD.n94 0.145
R2409 VDD.n128 VDD.n124 0.145
R2410 VDD.n132 VDD.n128 0.145
R2411 VDD.n136 VDD.n132 0.145
R2412 VDD.n144 VDD.n140 0.145
R2413 VDD.n148 VDD.n144 0.145
R2414 VDD.n152 VDD.n148 0.145
R2415 VDD.n183 VDD.n178 0.145
R2416 VDD.n188 VDD.n183 0.145
R2417 VDD.n194 VDD.n188 0.145
R2418 VDD.n204 VDD.n199 0.145
R2419 VDD.n209 VDD.n204 0.145
R2420 VDD.n213 VDD.n209 0.145
R2421 VDD.n244 VDD.n239 0.145
R2422 VDD.n249 VDD.n244 0.145
R2423 VDD.n255 VDD.n249 0.145
R2424 VDD.n265 VDD.n260 0.145
R2425 VDD.n270 VDD.n265 0.145
R2426 VDD.n274 VDD.n270 0.145
R2427 VDD.n304 VDD.n300 0.145
R2428 VDD.n308 VDD.n304 0.145
R2429 VDD.n313 VDD.n308 0.145
R2430 VDD.n320 VDD.n313 0.145
R2431 VDD.n325 VDD.n320 0.145
R2432 VDD.n337 VDD.n330 0.145
R2433 VDD.n342 VDD.n337 0.145
R2434 VDD.n347 VDD.n342 0.145
R2435 VDD.n351 VDD.n347 0.145
R2436 VDD.n355 VDD.n351 0.145
R2437 VDD.n385 VDD.n381 0.145
R2438 VDD.n389 VDD.n385 0.145
R2439 VDD.n394 VDD.n389 0.145
R2440 VDD.n401 VDD.n394 0.145
R2441 VDD.n406 VDD.n401 0.145
R2442 VDD.n418 VDD.n411 0.145
R2443 VDD.n423 VDD.n418 0.145
R2444 VDD.n428 VDD.n423 0.145
R2445 VDD.n432 VDD.n428 0.145
R2446 VDD.n436 VDD.n432 0.145
R2447 VDD.n467 VDD.n462 0.145
R2448 VDD.n472 VDD.n467 0.145
R2449 VDD.n478 VDD.n472 0.145
R2450 VDD.n488 VDD.n483 0.145
R2451 VDD.n493 VDD.n488 0.145
R2452 VDD.n497 VDD.n493 0.145
R2453 VDD.n527 VDD.n523 0.145
R2454 VDD.n531 VDD.n527 0.145
R2455 VDD.n536 VDD.n531 0.145
R2456 VDD.n543 VDD.n536 0.145
R2457 VDD.n548 VDD.n543 0.145
R2458 VDD.n560 VDD.n553 0.145
R2459 VDD.n565 VDD.n560 0.145
R2460 VDD.n570 VDD.n565 0.145
R2461 VDD.n574 VDD.n570 0.145
R2462 VDD.n578 VDD.n574 0.145
R2463 VDD.n608 VDD.n604 0.145
R2464 VDD.n612 VDD.n608 0.145
R2465 VDD.n617 VDD.n612 0.145
R2466 VDD.n624 VDD.n617 0.145
R2467 VDD.n629 VDD.n624 0.145
R2468 VDD.n641 VDD.n634 0.145
R2469 VDD.n646 VDD.n641 0.145
R2470 VDD.n651 VDD.n646 0.145
R2471 VDD.n655 VDD.n651 0.145
R2472 VDD.n659 VDD.n655 0.145
R2473 VDD.n690 VDD.n685 0.145
R2474 VDD.n695 VDD.n690 0.145
R2475 VDD.n701 VDD.n695 0.145
R2476 VDD.n711 VDD.n706 0.145
R2477 VDD.n716 VDD.n711 0.145
R2478 VDD.n720 VDD.n716 0.145
R2479 VDD.n750 VDD.n746 0.145
R2480 VDD.n754 VDD.n750 0.145
R2481 VDD.n759 VDD.n754 0.145
R2482 VDD.n766 VDD.n759 0.145
R2483 VDD.n771 VDD.n766 0.145
R2484 VDD.n783 VDD.n776 0.145
R2485 VDD.n788 VDD.n783 0.145
R2486 VDD.n1571 VDD.n1566 0.145
R2487 VDD.n1566 VDD.n1562 0.145
R2488 VDD.n1536 VDD.n1532 0.145
R2489 VDD.n1532 VDD.n1528 0.145
R2490 VDD.n1528 VDD.n1524 0.145
R2491 VDD.n1524 VDD.n1519 0.145
R2492 VDD.n1519 VDD.n1512 0.145
R2493 VDD.n1507 VDD.n1502 0.145
R2494 VDD.n1502 VDD.n1495 0.145
R2495 VDD.n1495 VDD.n1490 0.145
R2496 VDD.n1490 VDD.n1485 0.145
R2497 VDD.n1485 VDD.n1481 0.145
R2498 VDD.n1455 VDD.n1451 0.145
R2499 VDD.n1451 VDD.n1446 0.145
R2500 VDD.n1446 VDD.n1441 0.145
R2501 VDD.n1435 VDD.n1430 0.145
R2502 VDD.n1430 VDD.n1425 0.145
R2503 VDD.n1425 VDD.n1420 0.145
R2504 VDD.n1394 VDD.n1390 0.145
R2505 VDD.n1390 VDD.n1386 0.145
R2506 VDD.n1386 VDD.n1382 0.145
R2507 VDD.n1382 VDD.n1377 0.145
R2508 VDD.n1377 VDD.n1370 0.145
R2509 VDD.n1365 VDD.n1360 0.145
R2510 VDD.n1360 VDD.n1353 0.145
R2511 VDD.n1353 VDD.n1348 0.145
R2512 VDD.n1348 VDD.n1343 0.145
R2513 VDD.n1343 VDD.n1339 0.145
R2514 VDD.n1313 VDD.n1309 0.145
R2515 VDD.n1309 VDD.n1305 0.145
R2516 VDD.n1305 VDD.n1301 0.145
R2517 VDD.n1301 VDD.n1296 0.145
R2518 VDD.n1296 VDD.n1289 0.145
R2519 VDD.n1284 VDD.n1279 0.145
R2520 VDD.n1279 VDD.n1272 0.145
R2521 VDD.n1272 VDD.n1267 0.145
R2522 VDD.n1267 VDD.n1262 0.145
R2523 VDD.n1262 VDD.n1258 0.145
R2524 VDD.n1232 VDD.n1228 0.145
R2525 VDD.n1228 VDD.n1223 0.145
R2526 VDD.n1223 VDD.n1218 0.145
R2527 VDD.n1212 VDD.n1207 0.145
R2528 VDD.n1207 VDD.n1202 0.145
R2529 VDD.n1202 VDD.n1197 0.145
R2530 VDD.n1171 VDD.n1167 0.145
R2531 VDD.n1167 VDD.n1163 0.145
R2532 VDD.n1163 VDD.n1159 0.145
R2533 VDD.n1159 VDD.n1154 0.145
R2534 VDD.n1154 VDD.n1147 0.145
R2535 VDD.n1142 VDD.n1137 0.145
R2536 VDD.n1137 VDD.n1130 0.145
R2537 VDD.n1130 VDD.n1125 0.145
R2538 VDD.n1125 VDD.n1120 0.145
R2539 VDD.n1120 VDD.n1116 0.145
R2540 VDD.n1090 VDD.n1086 0.145
R2541 VDD.n1086 VDD.n1082 0.145
R2542 VDD.n1082 VDD.n1078 0.145
R2543 VDD.n1078 VDD.n1073 0.145
R2544 VDD.n1073 VDD.n1066 0.145
R2545 VDD.n1061 VDD.n1056 0.145
R2546 VDD.n1056 VDD.n1049 0.145
R2547 VDD.n1049 VDD.n1044 0.145
R2548 VDD.n1044 VDD.n1039 0.145
R2549 VDD.n1039 VDD.n1035 0.145
R2550 VDD.n1009 VDD.n1005 0.145
R2551 VDD.n1005 VDD.n1000 0.145
R2552 VDD.n1000 VDD.n995 0.145
R2553 VDD.n989 VDD.n984 0.145
R2554 VDD.n984 VDD.n979 0.145
R2555 VDD.n979 VDD.n974 0.145
R2556 VDD.n948 VDD.n944 0.145
R2557 VDD.n944 VDD.n940 0.145
R2558 VDD.n940 VDD.n936 0.145
R2559 VDD.n936 VDD.n931 0.145
R2560 VDD.n931 VDD.n924 0.145
R2561 VDD.n919 VDD.n914 0.145
R2562 VDD.n914 VDD.n907 0.145
R2563 VDD.n907 VDD.n902 0.145
R2564 VDD.n902 VDD.n897 0.145
R2565 VDD.n897 VDD.n893 0.145
R2566 VDD.n866 VDD.n862 0.145
R2567 VDD.n862 VDD.n858 0.145
R2568 VDD.n858 VDD.n854 0.145
R2569 VDD.n854 VDD.n849 0.145
R2570 VDD.n849 VDD.n842 0.145
R2571 VDD.n837 VDD.n832 0.145
R2572 VDD.n832 VDD.n825 0.145
R2573 VDD.n825 VDD.n820 0.145
R2574 VDD.n820 VDD.n815 0.145
R2575 VDD.n815 VDD.n811 0.145
R2576 VDD VDD.n1571 0.086
R2577 VDD VDD.n788 0.058
R2578 a_5779_989.n0 a_5779_989.t12 480.392
R2579 a_5779_989.n2 a_5779_989.t7 454.685
R2580 a_5779_989.n2 a_5779_989.t11 428.979
R2581 a_5779_989.n0 a_5779_989.t10 403.272
R2582 a_5779_989.n1 a_5779_989.t9 283.48
R2583 a_5779_989.n3 a_5779_989.t8 237.959
R2584 a_5779_989.n9 a_5779_989.n8 213.104
R2585 a_5779_989.n13 a_5779_989.n9 170.799
R2586 a_5779_989.n3 a_5779_989.n2 98.447
R2587 a_5779_989.n1 a_5779_989.n0 98.447
R2588 a_5779_989.n4 a_5779_989.n3 80.035
R2589 a_5779_989.n12 a_5779_989.n11 79.232
R2590 a_5779_989.n4 a_5779_989.n1 77.315
R2591 a_5779_989.n9 a_5779_989.n4 76
R2592 a_5779_989.n13 a_5779_989.n12 63.152
R2593 a_5779_989.n8 a_5779_989.n7 30
R2594 a_5779_989.n6 a_5779_989.n5 24.383
R2595 a_5779_989.n8 a_5779_989.n6 23.684
R2596 a_5779_989.n12 a_5779_989.n10 16.08
R2597 a_5779_989.n14 a_5779_989.n13 16.078
R2598 a_5779_989.n10 a_5779_989.t4 14.282
R2599 a_5779_989.n10 a_5779_989.t3 14.282
R2600 a_5779_989.n11 a_5779_989.t6 14.282
R2601 a_5779_989.n11 a_5779_989.t5 14.282
R2602 a_5779_989.n14 a_5779_989.t1 14.282
R2603 a_5779_989.t2 a_5779_989.n14 14.282
R2604 a_9331_989.n5 a_9331_989.t13 512.525
R2605 a_9331_989.n3 a_9331_989.t6 477.179
R2606 a_9331_989.n8 a_9331_989.t5 454.685
R2607 a_9331_989.n8 a_9331_989.t8 428.979
R2608 a_9331_989.n3 a_9331_989.t11 406.485
R2609 a_9331_989.n5 a_9331_989.t9 371.139
R2610 a_9331_989.n4 a_9331_989.t7 363.924
R2611 a_9331_989.n7 a_9331_989.t10 250.5
R2612 a_9331_989.n9 a_9331_989.t12 211.406
R2613 a_9331_989.n13 a_9331_989.n11 190.561
R2614 a_9331_989.n11 a_9331_989.n2 179.052
R2615 a_9331_989.n9 a_9331_989.n8 125
R2616 a_9331_989.n7 a_9331_989.n6 106.997
R2617 a_9331_989.n6 a_9331_989.n4 101.359
R2618 a_9331_989.n10 a_9331_989.n7 96.087
R2619 a_9331_989.n10 a_9331_989.n9 78.947
R2620 a_9331_989.n2 a_9331_989.n1 76.002
R2621 a_9331_989.n11 a_9331_989.n10 76
R2622 a_9331_989.n6 a_9331_989.n5 71.88
R2623 a_9331_989.n4 a_9331_989.n3 15.776
R2624 a_9331_989.n13 a_9331_989.n12 15.218
R2625 a_9331_989.n0 a_9331_989.t2 14.282
R2626 a_9331_989.n0 a_9331_989.t4 14.282
R2627 a_9331_989.n1 a_9331_989.t0 14.282
R2628 a_9331_989.n1 a_9331_989.t1 14.282
R2629 a_9331_989.n2 a_9331_989.n0 12.85
R2630 a_9331_989.n14 a_9331_989.n13 12.014
R2631 a_9009_1050.n0 a_9009_1050.t9 480.392
R2632 a_9009_1050.n0 a_9009_1050.t7 403.272
R2633 a_9009_1050.n1 a_9009_1050.t8 310.033
R2634 a_9009_1050.n6 a_9009_1050.n5 239.657
R2635 a_9009_1050.n6 a_9009_1050.n1 153.315
R2636 a_9009_1050.n10 a_9009_1050.n6 144.246
R2637 a_9009_1050.n9 a_9009_1050.n8 79.232
R2638 a_9009_1050.n1 a_9009_1050.n0 71.894
R2639 a_9009_1050.n10 a_9009_1050.n9 63.152
R2640 a_9009_1050.n5 a_9009_1050.n4 30
R2641 a_9009_1050.n3 a_9009_1050.n2 24.383
R2642 a_9009_1050.n5 a_9009_1050.n3 23.684
R2643 a_9009_1050.n9 a_9009_1050.n7 16.08
R2644 a_9009_1050.n11 a_9009_1050.n10 16.078
R2645 a_9009_1050.n7 a_9009_1050.t5 14.282
R2646 a_9009_1050.n7 a_9009_1050.t4 14.282
R2647 a_9009_1050.n8 a_9009_1050.t6 14.282
R2648 a_9009_1050.n8 a_9009_1050.t3 14.282
R2649 a_9009_1050.n11 a_9009_1050.t1 14.282
R2650 a_9009_1050.t2 a_9009_1050.n11 14.282
R2651 a_147_187.n4 a_147_187.t9 512.525
R2652 a_147_187.n2 a_147_187.t11 472.359
R2653 a_147_187.n0 a_147_187.t8 472.359
R2654 a_147_187.n2 a_147_187.t14 384.527
R2655 a_147_187.n0 a_147_187.t12 384.527
R2656 a_147_187.n4 a_147_187.t13 371.139
R2657 a_147_187.n5 a_147_187.t10 340.774
R2658 a_147_187.n3 a_147_187.t7 294.278
R2659 a_147_187.n1 a_147_187.t15 294.278
R2660 a_147_187.n12 a_147_187.n11 266.21
R2661 a_147_187.n16 a_147_187.n12 117.693
R2662 a_147_187.n5 a_147_187.n4 109.607
R2663 a_147_187.n6 a_147_187.n5 83.572
R2664 a_147_187.n7 a_147_187.n1 81.396
R2665 a_147_187.n15 a_147_187.n14 79.232
R2666 a_147_187.n6 a_147_187.n3 76
R2667 a_147_187.n12 a_147_187.n7 76
R2668 a_147_187.n16 a_147_187.n15 63.152
R2669 a_147_187.n3 a_147_187.n2 56.954
R2670 a_147_187.n1 a_147_187.n0 56.954
R2671 a_147_187.n11 a_147_187.n10 30
R2672 a_147_187.n9 a_147_187.n8 24.383
R2673 a_147_187.n11 a_147_187.n9 23.684
R2674 a_147_187.n15 a_147_187.n13 16.08
R2675 a_147_187.n17 a_147_187.n16 16.078
R2676 a_147_187.n13 a_147_187.t0 14.282
R2677 a_147_187.n13 a_147_187.t6 14.282
R2678 a_147_187.n14 a_147_187.t5 14.282
R2679 a_147_187.n14 a_147_187.t4 14.282
R2680 a_147_187.t3 a_147_187.n17 14.282
R2681 a_147_187.n17 a_147_187.t2 14.282
R2682 a_147_187.n7 a_147_187.n6 4.035
R2683 a_2036_101.t0 a_2036_101.n1 34.62
R2684 a_2036_101.t0 a_2036_101.n0 8.137
R2685 a_2036_101.t0 a_2036_101.n2 4.69
R2686 a_2141_1050.n0 a_2141_1050.t5 512.525
R2687 a_2141_1050.n0 a_2141_1050.t7 371.139
R2688 a_2141_1050.n1 a_2141_1050.t6 287.668
R2689 a_2141_1050.n3 a_2141_1050.n2 232.331
R2690 a_2141_1050.n1 a_2141_1050.n0 162.713
R2691 a_2141_1050.n3 a_2141_1050.n1 153.315
R2692 a_2141_1050.n5 a_2141_1050.n3 152.499
R2693 a_2141_1050.n5 a_2141_1050.n4 76.002
R2694 a_2141_1050.n4 a_2141_1050.t4 14.282
R2695 a_2141_1050.n4 a_2141_1050.t3 14.282
R2696 a_2141_1050.t2 a_2141_1050.n6 14.282
R2697 a_2141_1050.n6 a_2141_1050.t1 14.282
R2698 a_2141_1050.n6 a_2141_1050.n5 12.848
R2699 a_15932_209.n3 a_15932_209.t9 512.525
R2700 a_15932_209.n3 a_15932_209.t7 371.139
R2701 a_15932_209.n4 a_15932_209.t8 263.54
R2702 a_15932_209.n13 a_15932_209.n5 216.728
R2703 a_15932_209.n5 a_15932_209.n4 153.043
R2704 a_15932_209.n5 a_15932_209.n2 126.664
R2705 a_15932_209.n4 a_15932_209.n3 120.094
R2706 a_15932_209.n12 a_15932_209.n11 114.024
R2707 a_15932_209.n12 a_15932_209.n8 111.94
R2708 a_15932_209.n13 a_15932_209.n12 78.403
R2709 a_15932_209.n2 a_15932_209.n1 75.271
R2710 a_15932_209.n15 a_15932_209.n13 27.275
R2711 a_15932_209.n8 a_15932_209.n7 22.578
R2712 a_15932_209.n11 a_15932_209.n10 22.578
R2713 a_15932_209.n15 a_15932_209.n14 15.001
R2714 a_15932_209.n0 a_15932_209.t6 14.282
R2715 a_15932_209.n0 a_15932_209.t1 14.282
R2716 a_15932_209.n1 a_15932_209.t5 14.282
R2717 a_15932_209.n1 a_15932_209.t2 14.282
R2718 a_15932_209.n16 a_15932_209.n15 12.632
R2719 a_15932_209.n2 a_15932_209.n0 12.119
R2720 a_15932_209.n8 a_15932_209.n6 8.58
R2721 a_15932_209.n11 a_15932_209.n9 8.58
R2722 Q.n2 Q.n1 253.86
R2723 Q.n2 Q.n0 130.901
R2724 Q.n3 Q.n2 76
R2725 Q.n0 Q.t1 14.282
R2726 Q.n0 Q.t2 14.282
R2727 Q.n3 Q 0.046
R2728 CLK.n14 CLK.t4 459.505
R2729 CLK.n11 CLK.t17 459.505
R2730 CLK.n8 CLK.t16 459.505
R2731 CLK.n5 CLK.t15 459.505
R2732 CLK.n2 CLK.t6 459.505
R2733 CLK.n0 CLK.t5 459.505
R2734 CLK.n14 CLK.t11 384.527
R2735 CLK.n11 CLK.t7 384.527
R2736 CLK.n8 CLK.t0 384.527
R2737 CLK.n5 CLK.t3 384.527
R2738 CLK.n2 CLK.t12 384.527
R2739 CLK.n0 CLK.t13 384.527
R2740 CLK.n15 CLK.t8 322.152
R2741 CLK.n12 CLK.t14 322.151
R2742 CLK.n9 CLK.t9 322.151
R2743 CLK.n6 CLK.t2 322.151
R2744 CLK.n3 CLK.t1 322.151
R2745 CLK.n1 CLK.t10 322.151
R2746 CLK.n4 CLK.n1 58.818
R2747 CLK.n16 CLK.n15 49.342
R2748 CLK.n4 CLK.n3 49.342
R2749 CLK.n7 CLK.n6 49.342
R2750 CLK.n10 CLK.n9 49.342
R2751 CLK.n13 CLK.n12 49.342
R2752 CLK.n15 CLK.n14 27.599
R2753 CLK.n1 CLK.n0 27.599
R2754 CLK.n3 CLK.n2 27.599
R2755 CLK.n6 CLK.n5 27.599
R2756 CLK.n9 CLK.n8 27.599
R2757 CLK.n12 CLK.n11 27.599
R2758 CLK.n7 CLK.n4 9.476
R2759 CLK.n10 CLK.n7 9.476
R2760 CLK.n13 CLK.n10 9.476
R2761 CLK.n16 CLK.n13 9.476
R2762 CLK.n16 CLK 0.046
R2763 a_5457_1050.n2 a_5457_1050.t9 512.525
R2764 a_5457_1050.n0 a_5457_1050.t10 512.525
R2765 a_5457_1050.n2 a_5457_1050.t12 371.139
R2766 a_5457_1050.n0 a_5457_1050.t11 371.139
R2767 a_5457_1050.n3 a_5457_1050.t8 314.221
R2768 a_5457_1050.n1 a_5457_1050.t7 314.221
R2769 a_5457_1050.n9 a_5457_1050.n8 239.657
R2770 a_5457_1050.n13 a_5457_1050.n9 144.246
R2771 a_5457_1050.n3 a_5457_1050.n2 136.16
R2772 a_5457_1050.n1 a_5457_1050.n0 136.16
R2773 a_5457_1050.n4 a_5457_1050.n1 85.476
R2774 a_5457_1050.n12 a_5457_1050.n11 79.232
R2775 a_5457_1050.n9 a_5457_1050.n4 77.315
R2776 a_5457_1050.n4 a_5457_1050.n3 76
R2777 a_5457_1050.n13 a_5457_1050.n12 63.152
R2778 a_5457_1050.n8 a_5457_1050.n7 30
R2779 a_5457_1050.n6 a_5457_1050.n5 24.383
R2780 a_5457_1050.n8 a_5457_1050.n6 23.684
R2781 a_5457_1050.n12 a_5457_1050.n10 16.08
R2782 a_5457_1050.n14 a_5457_1050.n13 16.078
R2783 a_5457_1050.n10 a_5457_1050.t5 14.282
R2784 a_5457_1050.n10 a_5457_1050.t6 14.282
R2785 a_5457_1050.n11 a_5457_1050.t4 14.282
R2786 a_5457_1050.n11 a_5457_1050.t3 14.282
R2787 a_5457_1050.n14 a_5457_1050.t0 14.282
R2788 a_5457_1050.t1 a_5457_1050.n14 14.282
R2789 a_10507_187.n4 a_10507_187.t9 512.525
R2790 a_10507_187.n2 a_10507_187.t13 472.359
R2791 a_10507_187.n0 a_10507_187.t12 472.359
R2792 a_10507_187.n2 a_10507_187.t15 384.527
R2793 a_10507_187.n0 a_10507_187.t14 384.527
R2794 a_10507_187.n4 a_10507_187.t10 371.139
R2795 a_10507_187.n5 a_10507_187.t7 340.774
R2796 a_10507_187.n3 a_10507_187.t11 294.278
R2797 a_10507_187.n1 a_10507_187.t8 294.278
R2798 a_10507_187.n12 a_10507_187.n11 266.21
R2799 a_10507_187.n16 a_10507_187.n12 117.693
R2800 a_10507_187.n5 a_10507_187.n4 109.607
R2801 a_10507_187.n6 a_10507_187.n5 83.572
R2802 a_10507_187.n7 a_10507_187.n1 81.396
R2803 a_10507_187.n15 a_10507_187.n14 79.232
R2804 a_10507_187.n6 a_10507_187.n3 76
R2805 a_10507_187.n12 a_10507_187.n7 76
R2806 a_10507_187.n16 a_10507_187.n15 63.152
R2807 a_10507_187.n3 a_10507_187.n2 56.954
R2808 a_10507_187.n1 a_10507_187.n0 56.954
R2809 a_10507_187.n11 a_10507_187.n10 30
R2810 a_10507_187.n9 a_10507_187.n8 24.383
R2811 a_10507_187.n11 a_10507_187.n9 23.684
R2812 a_10507_187.n15 a_10507_187.n13 16.08
R2813 a_10507_187.n17 a_10507_187.n16 16.078
R2814 a_10507_187.n13 a_10507_187.t6 14.282
R2815 a_10507_187.n13 a_10507_187.t5 14.282
R2816 a_10507_187.n14 a_10507_187.t0 14.282
R2817 a_10507_187.n14 a_10507_187.t4 14.282
R2818 a_10507_187.t3 a_10507_187.n17 14.282
R2819 a_10507_187.n17 a_10507_187.t2 14.282
R2820 a_10507_187.n7 a_10507_187.n6 4.035
R2821 a_10451_103.n4 a_10451_103.n3 19.724
R2822 a_10451_103.t0 a_10451_103.n5 11.595
R2823 a_10451_103.t0 a_10451_103.n4 9.207
R2824 a_10451_103.n2 a_10451_103.n0 8.543
R2825 a_10451_103.t0 a_10451_103.n2 3.034
R2826 a_10451_103.n2 a_10451_103.n1 0.443
R2827 a_16421_1051.n4 a_16421_1051.n3 196.002
R2828 a_16421_1051.n2 a_16421_1051.t7 89.553
R2829 a_16421_1051.n5 a_16421_1051.n4 75.27
R2830 a_16421_1051.n3 a_16421_1051.n2 75.214
R2831 a_16421_1051.n4 a_16421_1051.n0 36.52
R2832 a_16421_1051.n3 a_16421_1051.t4 14.338
R2833 a_16421_1051.n0 a_16421_1051.t5 14.282
R2834 a_16421_1051.n0 a_16421_1051.t2 14.282
R2835 a_16421_1051.n1 a_16421_1051.t3 14.282
R2836 a_16421_1051.n1 a_16421_1051.t6 14.282
R2837 a_16421_1051.t0 a_16421_1051.n5 14.282
R2838 a_16421_1051.n5 a_16421_1051.t1 14.282
R2839 a_16421_1051.n2 a_16421_1051.n1 12.119
R2840 a_15757_1051.n4 a_15757_1051.n3 195.987
R2841 a_15757_1051.n2 a_15757_1051.t6 89.553
R2842 a_15757_1051.n5 a_15757_1051.n4 75.27
R2843 a_15757_1051.n3 a_15757_1051.n2 75.214
R2844 a_15757_1051.n4 a_15757_1051.n0 36.519
R2845 a_15757_1051.n3 a_15757_1051.t2 14.338
R2846 a_15757_1051.n0 a_15757_1051.t4 14.282
R2847 a_15757_1051.n0 a_15757_1051.t7 14.282
R2848 a_15757_1051.n1 a_15757_1051.t5 14.282
R2849 a_15757_1051.n1 a_15757_1051.t3 14.282
R2850 a_15757_1051.n5 a_15757_1051.t0 14.282
R2851 a_15757_1051.t1 a_15757_1051.n5 14.282
R2852 a_15757_1051.n2 a_15757_1051.n1 12.119
R2853 a_14511_989.n1 a_14511_989.t7 475.572
R2854 a_14511_989.n0 a_14511_989.t9 469.145
R2855 a_14511_989.n5 a_14511_989.t11 454.685
R2856 a_14511_989.n5 a_14511_989.t5 428.979
R2857 a_14511_989.n1 a_14511_989.t13 384.527
R2858 a_14511_989.n0 a_14511_989.t12 384.527
R2859 a_14511_989.n2 a_14511_989.t8 294.278
R2860 a_14511_989.n4 a_14511_989.t6 241.172
R2861 a_14511_989.n6 a_14511_989.t10 237.959
R2862 a_14511_989.n12 a_14511_989.n11 210.592
R2863 a_14511_989.n3 a_14511_989.n2 156.851
R2864 a_14511_989.n14 a_14511_989.n12 152.499
R2865 a_14511_989.n6 a_14511_989.n5 98.447
R2866 a_14511_989.n7 a_14511_989.n6 78.947
R2867 a_14511_989.n7 a_14511_989.n4 77.859
R2868 a_14511_989.n14 a_14511_989.n13 76.002
R2869 a_14511_989.n12 a_14511_989.n7 76
R2870 a_14511_989.n2 a_14511_989.n1 57.842
R2871 a_14511_989.n3 a_14511_989.n0 56.833
R2872 a_14511_989.n4 a_14511_989.n3 53.105
R2873 a_14511_989.n11 a_14511_989.n10 30
R2874 a_14511_989.n9 a_14511_989.n8 24.383
R2875 a_14511_989.n11 a_14511_989.n9 23.684
R2876 a_14511_989.n13 a_14511_989.t4 14.282
R2877 a_14511_989.n13 a_14511_989.t0 14.282
R2878 a_14511_989.t2 a_14511_989.n15 14.282
R2879 a_14511_989.n15 a_14511_989.t1 14.282
R2880 a_14511_989.n15 a_14511_989.n14 12.848
R2881 a_14189_1050.n1 a_14189_1050.t8 480.392
R2882 a_14189_1050.n1 a_14189_1050.t7 403.272
R2883 a_14189_1050.n2 a_14189_1050.t9 310.033
R2884 a_14189_1050.n7 a_14189_1050.n6 239.657
R2885 a_14189_1050.n7 a_14189_1050.n2 153.315
R2886 a_14189_1050.n8 a_14189_1050.n7 144.246
R2887 a_14189_1050.n10 a_14189_1050.n9 79.232
R2888 a_14189_1050.n2 a_14189_1050.n1 71.894
R2889 a_14189_1050.n10 a_14189_1050.n8 63.152
R2890 a_14189_1050.n6 a_14189_1050.n5 30
R2891 a_14189_1050.n4 a_14189_1050.n3 24.383
R2892 a_14189_1050.n6 a_14189_1050.n4 23.684
R2893 a_14189_1050.n8 a_14189_1050.n0 16.08
R2894 a_14189_1050.n11 a_14189_1050.n10 16.078
R2895 a_14189_1050.n0 a_14189_1050.t5 14.282
R2896 a_14189_1050.n0 a_14189_1050.t4 14.282
R2897 a_14189_1050.n9 a_14189_1050.t0 14.282
R2898 a_14189_1050.n9 a_14189_1050.t6 14.282
R2899 a_14189_1050.n11 a_14189_1050.t1 14.282
R2900 a_14189_1050.t2 a_14189_1050.n11 14.282
R2901 a_15652_101.n13 a_15652_101.n12 26.811
R2902 a_15652_101.n6 a_15652_101.n5 24.977
R2903 a_15652_101.n2 a_15652_101.n1 24.877
R2904 a_15652_101.t0 a_15652_101.n2 12.677
R2905 a_15652_101.t0 a_15652_101.n3 11.595
R2906 a_15652_101.n11 a_15652_101.n10 8.561
R2907 a_15652_101.t0 a_15652_101.n4 7.273
R2908 a_15652_101.n9 a_15652_101.n8 7.066
R2909 a_15652_101.t0 a_15652_101.n0 6.109
R2910 a_15652_101.t1 a_15652_101.n7 4.864
R2911 a_15652_101.t0 a_15652_101.n13 2.074
R2912 a_15652_101.n7 a_15652_101.n6 1.13
R2913 a_15652_101.t1 a_15652_101.n11 0.958
R2914 a_15652_101.n13 a_15652_101.t1 0.937
R2915 a_15652_101.t1 a_15652_101.n9 0.86
R2916 a_6514_210.n8 a_6514_210.n6 96.467
R2917 a_6514_210.n3 a_6514_210.n1 44.628
R2918 a_6514_210.t0 a_6514_210.n8 32.417
R2919 a_6514_210.n3 a_6514_210.n2 23.284
R2920 a_6514_210.n6 a_6514_210.n5 22.349
R2921 a_6514_210.t0 a_6514_210.n10 20.241
R2922 a_6514_210.n10 a_6514_210.n9 13.494
R2923 a_6514_210.n6 a_6514_210.n4 8.443
R2924 a_6514_210.t0 a_6514_210.n0 8.137
R2925 a_6514_210.t0 a_6514_210.n3 5.727
R2926 a_6514_210.n8 a_6514_210.n7 1.435
R2927 a_4151_989.n1 a_4151_989.t5 512.525
R2928 a_4151_989.n0 a_4151_989.t11 512.525
R2929 a_4151_989.n5 a_4151_989.t7 454.685
R2930 a_4151_989.n5 a_4151_989.t12 428.979
R2931 a_4151_989.n1 a_4151_989.t9 371.139
R2932 a_4151_989.n0 a_4151_989.t6 371.139
R2933 a_4151_989.n2 a_4151_989.n1 265.439
R2934 a_4151_989.n4 a_4151_989.n0 212.333
R2935 a_4151_989.n14 a_4151_989.n12 205.605
R2936 a_4151_989.n2 a_4151_989.t13 176.995
R2937 a_4151_989.n6 a_4151_989.t8 173.606
R2938 a_4151_989.n3 a_4151_989.t10 170.569
R2939 a_4151_989.n12 a_4151_989.n11 157.486
R2940 a_4151_989.n3 a_4151_989.n2 153.043
R2941 a_4151_989.n6 a_4151_989.n5 151.553
R2942 a_4151_989.n7 a_4151_989.n4 118.94
R2943 a_4151_989.n7 a_4151_989.n6 78.947
R2944 a_4151_989.n14 a_4151_989.n13 76.002
R2945 a_4151_989.n12 a_4151_989.n7 76
R2946 a_4151_989.n4 a_4151_989.n3 53.105
R2947 a_4151_989.n11 a_4151_989.n10 30
R2948 a_4151_989.n9 a_4151_989.n8 24.383
R2949 a_4151_989.n11 a_4151_989.n9 23.684
R2950 a_4151_989.n13 a_4151_989.t4 14.282
R2951 a_4151_989.n13 a_4151_989.t0 14.282
R2952 a_4151_989.t3 a_4151_989.n15 14.282
R2953 a_4151_989.n15 a_4151_989.t2 14.282
R2954 a_4151_989.n15 a_4151_989.n14 12.848
R2955 a_5327_187.n4 a_5327_187.t11 512.525
R2956 a_5327_187.n2 a_5327_187.t7 472.359
R2957 a_5327_187.n0 a_5327_187.t15 472.359
R2958 a_5327_187.n2 a_5327_187.t12 384.527
R2959 a_5327_187.n0 a_5327_187.t8 384.527
R2960 a_5327_187.n4 a_5327_187.t14 371.139
R2961 a_5327_187.n5 a_5327_187.t9 340.774
R2962 a_5327_187.n3 a_5327_187.t13 294.278
R2963 a_5327_187.n1 a_5327_187.t10 294.278
R2964 a_5327_187.n12 a_5327_187.n11 266.21
R2965 a_5327_187.n16 a_5327_187.n12 117.693
R2966 a_5327_187.n5 a_5327_187.n4 109.607
R2967 a_5327_187.n6 a_5327_187.n5 83.572
R2968 a_5327_187.n7 a_5327_187.n1 81.396
R2969 a_5327_187.n15 a_5327_187.n14 79.232
R2970 a_5327_187.n6 a_5327_187.n3 76
R2971 a_5327_187.n12 a_5327_187.n7 76
R2972 a_5327_187.n16 a_5327_187.n15 63.152
R2973 a_5327_187.n3 a_5327_187.n2 56.954
R2974 a_5327_187.n1 a_5327_187.n0 56.954
R2975 a_5327_187.n11 a_5327_187.n10 30
R2976 a_5327_187.n9 a_5327_187.n8 24.383
R2977 a_5327_187.n11 a_5327_187.n9 23.684
R2978 a_5327_187.n15 a_5327_187.n13 16.08
R2979 a_5327_187.n17 a_5327_187.n16 16.078
R2980 a_5327_187.n13 a_5327_187.t4 14.282
R2981 a_5327_187.n13 a_5327_187.t5 14.282
R2982 a_5327_187.n14 a_5327_187.t3 14.282
R2983 a_5327_187.n14 a_5327_187.t6 14.282
R2984 a_5327_187.n17 a_5327_187.t0 14.282
R2985 a_5327_187.t1 a_5327_187.n17 14.282
R2986 a_5327_187.n7 a_5327_187.n6 4.035
R2987 a_7321_1050.n0 a_7321_1050.t6 512.525
R2988 a_7321_1050.n0 a_7321_1050.t7 371.139
R2989 a_7321_1050.n1 a_7321_1050.t5 287.668
R2990 a_7321_1050.n6 a_7321_1050.n5 210.592
R2991 a_7321_1050.n1 a_7321_1050.n0 162.713
R2992 a_7321_1050.n6 a_7321_1050.n1 153.315
R2993 a_7321_1050.n8 a_7321_1050.n6 152.499
R2994 a_7321_1050.n8 a_7321_1050.n7 76.002
R2995 a_7321_1050.n5 a_7321_1050.n4 30
R2996 a_7321_1050.n3 a_7321_1050.n2 24.383
R2997 a_7321_1050.n5 a_7321_1050.n3 23.684
R2998 a_7321_1050.n7 a_7321_1050.t3 14.282
R2999 a_7321_1050.n7 a_7321_1050.t4 14.282
R3000 a_7321_1050.t1 a_7321_1050.n9 14.282
R3001 a_7321_1050.n9 a_7321_1050.t0 14.282
R3002 a_7321_1050.n9 a_7321_1050.n8 12.848
R3003 D.n5 D.t5 479.223
R3004 D.n2 D.t4 479.223
R3005 D.n0 D.t7 479.223
R3006 D.n5 D.t1 375.52
R3007 D.n2 D.t6 375.52
R3008 D.n0 D.t2 375.52
R3009 D.n6 D.n5 201.982
R3010 D.n3 D.n2 201.982
R3011 D.n1 D.n0 201.982
R3012 D.n6 D.t8 141.649
R3013 D.n3 D.t3 141.649
R3014 D.n1 D.t0 141.649
R3015 D.n4 D.n1 94.999
R3016 D.n4 D.n3 76
R3017 D.n7 D.n6 76
R3018 D.n7 D.n4 18.999
R3019 D.n7 D 0.046
R3020 a_11413_103.n1 a_11413_103.n0 25.576
R3021 a_11413_103.n3 a_11413_103.n2 9.111
R3022 a_11413_103.n7 a_11413_103.n5 7.859
R3023 a_11413_103.t0 a_11413_103.n7 3.034
R3024 a_11413_103.n5 a_11413_103.n3 1.964
R3025 a_11413_103.n5 a_11413_103.n4 1.964
R3026 a_11413_103.t0 a_11413_103.n1 1.871
R3027 a_11413_103.n7 a_11413_103.n6 0.443
R3028 a_11694_210.n8 a_11694_210.n6 96.467
R3029 a_11694_210.n3 a_11694_210.n1 44.628
R3030 a_11694_210.t0 a_11694_210.n8 32.417
R3031 a_11694_210.n3 a_11694_210.n2 23.284
R3032 a_11694_210.n6 a_11694_210.n5 22.349
R3033 a_11694_210.t0 a_11694_210.n10 20.241
R3034 a_11694_210.n10 a_11694_210.n9 13.494
R3035 a_11694_210.n6 a_11694_210.n4 8.443
R3036 a_11694_210.t0 a_11694_210.n0 8.137
R3037 a_11694_210.t0 a_11694_210.n3 5.727
R3038 a_11694_210.n8 a_11694_210.n7 1.435
R3039 a_14986_101.t0 a_14986_101.n1 34.62
R3040 a_14986_101.t0 a_14986_101.n0 8.137
R3041 a_14986_101.t0 a_14986_101.n2 4.69
R3042 a_12501_1050.n1 a_12501_1050.t5 512.525
R3043 a_12501_1050.n1 a_12501_1050.t7 371.139
R3044 a_12501_1050.n2 a_12501_1050.t6 287.668
R3045 a_12501_1050.n4 a_12501_1050.n3 232.331
R3046 a_12501_1050.n2 a_12501_1050.n1 162.713
R3047 a_12501_1050.n4 a_12501_1050.n2 153.315
R3048 a_12501_1050.n5 a_12501_1050.n4 152.499
R3049 a_12501_1050.n6 a_12501_1050.n5 76.001
R3050 a_12501_1050.n0 a_12501_1050.t4 14.282
R3051 a_12501_1050.n0 a_12501_1050.t3 14.282
R3052 a_12501_1050.n6 a_12501_1050.t0 14.282
R3053 a_12501_1050.t1 a_12501_1050.n6 14.282
R3054 a_12501_1050.n5 a_12501_1050.n0 12.85
R3055 a_8823_103.n4 a_8823_103.n3 19.724
R3056 a_8823_103.t0 a_8823_103.n5 11.595
R3057 a_8823_103.t0 a_8823_103.n4 9.207
R3058 a_8823_103.n2 a_8823_103.n0 8.543
R3059 a_8823_103.t0 a_8823_103.n2 3.034
R3060 a_8823_103.n2 a_8823_103.n1 0.443
R3061 a_9104_210.n8 a_9104_210.n6 96.467
R3062 a_9104_210.n3 a_9104_210.n1 44.628
R3063 a_9104_210.t0 a_9104_210.n8 32.417
R3064 a_9104_210.n3 a_9104_210.n2 23.284
R3065 a_9104_210.n6 a_9104_210.n5 22.349
R3066 a_9104_210.t0 a_9104_210.n10 20.241
R3067 a_9104_210.n10 a_9104_210.n9 13.494
R3068 a_9104_210.n6 a_9104_210.n4 8.443
R3069 a_9104_210.t0 a_9104_210.n0 8.137
R3070 a_9104_210.t0 a_9104_210.n3 5.727
R3071 a_9104_210.n8 a_9104_210.n7 1.435
R3072 a_277_1050.n4 a_277_1050.t9 512.525
R3073 a_277_1050.n2 a_277_1050.t7 512.525
R3074 a_277_1050.n4 a_277_1050.t12 371.139
R3075 a_277_1050.n2 a_277_1050.t10 371.139
R3076 a_277_1050.n5 a_277_1050.t11 314.221
R3077 a_277_1050.n3 a_277_1050.t8 314.221
R3078 a_277_1050.n8 a_277_1050.n7 261.396
R3079 a_277_1050.n9 a_277_1050.n8 144.246
R3080 a_277_1050.n5 a_277_1050.n4 136.16
R3081 a_277_1050.n3 a_277_1050.n2 136.16
R3082 a_277_1050.n6 a_277_1050.n3 85.476
R3083 a_277_1050.n11 a_277_1050.n10 79.231
R3084 a_277_1050.n8 a_277_1050.n6 77.315
R3085 a_277_1050.n6 a_277_1050.n5 76
R3086 a_277_1050.n10 a_277_1050.n9 63.152
R3087 a_277_1050.n9 a_277_1050.n1 16.08
R3088 a_277_1050.n10 a_277_1050.n0 16.08
R3089 a_277_1050.n1 a_277_1050.t4 14.282
R3090 a_277_1050.n1 a_277_1050.t3 14.282
R3091 a_277_1050.n0 a_277_1050.t6 14.282
R3092 a_277_1050.n0 a_277_1050.t5 14.282
R3093 a_277_1050.t2 a_277_1050.n11 14.282
R3094 a_277_1050.n11 a_277_1050.t1 14.282
R3095 a_16318_101.t0 a_16318_101.n0 34.602
R3096 a_16318_101.t0 a_16318_101.n1 2.138
R3097 a_10637_1050.n2 a_10637_1050.t11 512.525
R3098 a_10637_1050.n0 a_10637_1050.t10 512.525
R3099 a_10637_1050.n2 a_10637_1050.t8 371.139
R3100 a_10637_1050.n0 a_10637_1050.t7 371.139
R3101 a_10637_1050.n3 a_10637_1050.t12 314.221
R3102 a_10637_1050.n1 a_10637_1050.t9 314.221
R3103 a_10637_1050.n9 a_10637_1050.n8 239.657
R3104 a_10637_1050.n13 a_10637_1050.n9 144.246
R3105 a_10637_1050.n3 a_10637_1050.n2 136.16
R3106 a_10637_1050.n1 a_10637_1050.n0 136.16
R3107 a_10637_1050.n4 a_10637_1050.n1 85.476
R3108 a_10637_1050.n12 a_10637_1050.n11 79.232
R3109 a_10637_1050.n9 a_10637_1050.n4 77.315
R3110 a_10637_1050.n4 a_10637_1050.n3 76
R3111 a_10637_1050.n13 a_10637_1050.n12 63.152
R3112 a_10637_1050.n8 a_10637_1050.n7 30
R3113 a_10637_1050.n6 a_10637_1050.n5 24.383
R3114 a_10637_1050.n8 a_10637_1050.n6 23.684
R3115 a_10637_1050.n12 a_10637_1050.n10 16.08
R3116 a_10637_1050.n14 a_10637_1050.n13 16.078
R3117 a_10637_1050.n10 a_10637_1050.t6 14.282
R3118 a_10637_1050.n10 a_10637_1050.t5 14.282
R3119 a_10637_1050.n11 a_10637_1050.t4 14.282
R3120 a_10637_1050.n11 a_10637_1050.t3 14.282
R3121 a_10637_1050.t2 a_10637_1050.n14 14.282
R3122 a_10637_1050.n14 a_10637_1050.t1 14.282
R3123 a_599_989.n0 a_599_989.t8 480.392
R3124 a_599_989.n2 a_599_989.t12 454.685
R3125 a_599_989.n2 a_599_989.t9 428.979
R3126 a_599_989.n0 a_599_989.t11 403.272
R3127 a_599_989.n1 a_599_989.t10 283.48
R3128 a_599_989.n3 a_599_989.t7 237.959
R3129 a_599_989.n9 a_599_989.n8 213.104
R3130 a_599_989.n13 a_599_989.n9 170.799
R3131 a_599_989.n3 a_599_989.n2 98.447
R3132 a_599_989.n1 a_599_989.n0 98.447
R3133 a_599_989.n4 a_599_989.n3 80.035
R3134 a_599_989.n12 a_599_989.n11 79.232
R3135 a_599_989.n4 a_599_989.n1 77.315
R3136 a_599_989.n9 a_599_989.n4 76
R3137 a_599_989.n13 a_599_989.n12 63.152
R3138 a_599_989.n8 a_599_989.n7 30
R3139 a_599_989.n6 a_599_989.n5 24.383
R3140 a_599_989.n8 a_599_989.n6 23.684
R3141 a_599_989.n12 a_599_989.n10 16.08
R3142 a_599_989.n14 a_599_989.n13 16.078
R3143 a_599_989.n10 a_599_989.t3 14.282
R3144 a_599_989.n10 a_599_989.t4 14.282
R3145 a_599_989.n11 a_599_989.t6 14.282
R3146 a_599_989.n11 a_599_989.t5 14.282
R3147 a_599_989.n14 a_599_989.t0 14.282
R3148 a_599_989.t1 a_599_989.n14 14.282
R3149 a_372_210.n9 a_372_210.n7 82.852
R3150 a_372_210.n3 a_372_210.n1 44.628
R3151 a_372_210.t0 a_372_210.n9 32.417
R3152 a_372_210.n7 a_372_210.n6 27.2
R3153 a_372_210.n5 a_372_210.n4 23.498
R3154 a_372_210.n3 a_372_210.n2 23.284
R3155 a_372_210.n7 a_372_210.n5 22.4
R3156 a_372_210.t0 a_372_210.n11 20.241
R3157 a_372_210.n11 a_372_210.n10 13.494
R3158 a_372_210.t0 a_372_210.n0 8.137
R3159 a_372_210.t0 a_372_210.n3 5.727
R3160 a_372_210.n9 a_372_210.n8 1.435
R3161 a_10732_210.n8 a_10732_210.n6 96.467
R3162 a_10732_210.n3 a_10732_210.n1 44.628
R3163 a_10732_210.t0 a_10732_210.n8 32.417
R3164 a_10732_210.n3 a_10732_210.n2 23.284
R3165 a_10732_210.n6 a_10732_210.n5 22.349
R3166 a_10732_210.t0 a_10732_210.n10 20.241
R3167 a_10732_210.n10 a_10732_210.n9 13.494
R3168 a_10732_210.n6 a_10732_210.n4 8.443
R3169 a_10732_210.t0 a_10732_210.n0 8.137
R3170 a_10732_210.t0 a_10732_210.n3 5.727
R3171 a_10732_210.n8 a_10732_210.n7 1.435
R3172 a_6233_103.n5 a_6233_103.n4 19.724
R3173 a_6233_103.t0 a_6233_103.n3 11.595
R3174 a_6233_103.t0 a_6233_103.n5 9.207
R3175 a_6233_103.n2 a_6233_103.n1 2.455
R3176 a_6233_103.n2 a_6233_103.n0 1.32
R3177 a_6233_103.t0 a_6233_103.n2 0.246
R3178 a_5552_210.n9 a_5552_210.n7 82.852
R3179 a_5552_210.n3 a_5552_210.n1 44.628
R3180 a_5552_210.t0 a_5552_210.n9 32.417
R3181 a_5552_210.n7 a_5552_210.n6 27.2
R3182 a_5552_210.n5 a_5552_210.n4 23.498
R3183 a_5552_210.n3 a_5552_210.n2 23.284
R3184 a_5552_210.n7 a_5552_210.n5 22.4
R3185 a_5552_210.t0 a_5552_210.n11 20.241
R3186 a_5552_210.n11 a_5552_210.n10 13.494
R3187 a_5552_210.t0 a_5552_210.n0 8.137
R3188 a_5552_210.t0 a_5552_210.n3 5.727
R3189 a_5552_210.n9 a_5552_210.n8 1.435
R3190 a_16984_101.t0 a_16984_101.n1 34.62
R3191 a_16984_101.t0 a_16984_101.n0 8.137
R3192 a_16984_101.t0 a_16984_101.n2 4.69
R3193 a_2962_210.n9 a_2962_210.n7 82.852
R3194 a_2962_210.n3 a_2962_210.n1 44.628
R3195 a_2962_210.t0 a_2962_210.n9 32.417
R3196 a_2962_210.n7 a_2962_210.n6 27.2
R3197 a_2962_210.n5 a_2962_210.n4 23.498
R3198 a_2962_210.n3 a_2962_210.n2 23.284
R3199 a_2962_210.n7 a_2962_210.n5 22.4
R3200 a_2962_210.t0 a_2962_210.n11 20.241
R3201 a_2962_210.n11 a_2962_210.n10 13.494
R3202 a_2962_210.t0 a_2962_210.n0 8.137
R3203 a_2962_210.t0 a_2962_210.n3 5.727
R3204 a_2962_210.n9 a_2962_210.n8 1.435
R3205 a_7861_103.n4 a_7861_103.n3 19.724
R3206 a_7861_103.t0 a_7861_103.n5 11.595
R3207 a_7861_103.t0 a_7861_103.n4 9.207
R3208 a_7861_103.n2 a_7861_103.n0 8.543
R3209 a_7861_103.t0 a_7861_103.n2 3.034
R3210 a_7861_103.n2 a_7861_103.n1 0.443
R3211 a_8142_210.n8 a_8142_210.n6 96.467
R3212 a_8142_210.n3 a_8142_210.n1 44.628
R3213 a_8142_210.t0 a_8142_210.n8 32.417
R3214 a_8142_210.n3 a_8142_210.n2 23.284
R3215 a_8142_210.n6 a_8142_210.n5 22.349
R3216 a_8142_210.t0 a_8142_210.n10 20.241
R3217 a_8142_210.n10 a_8142_210.n9 13.494
R3218 a_8142_210.n6 a_8142_210.n4 8.443
R3219 a_8142_210.t0 a_8142_210.n0 8.137
R3220 a_8142_210.t0 a_8142_210.n3 5.727
R3221 a_8142_210.n8 a_8142_210.n7 1.435
R3222 a_9806_101.t0 a_9806_101.n1 34.62
R3223 a_9806_101.t0 a_9806_101.n0 8.137
R3224 a_9806_101.t0 a_9806_101.n2 4.69
R3225 a_3829_1050.n1 a_3829_1050.t9 480.392
R3226 a_3829_1050.n1 a_3829_1050.t7 403.272
R3227 a_3829_1050.n2 a_3829_1050.t8 310.033
R3228 a_3829_1050.n7 a_3829_1050.n6 239.657
R3229 a_3829_1050.n7 a_3829_1050.n2 153.315
R3230 a_3829_1050.n8 a_3829_1050.n7 144.246
R3231 a_3829_1050.n10 a_3829_1050.n9 79.232
R3232 a_3829_1050.n2 a_3829_1050.n1 71.894
R3233 a_3829_1050.n10 a_3829_1050.n8 63.152
R3234 a_3829_1050.n6 a_3829_1050.n5 30
R3235 a_3829_1050.n4 a_3829_1050.n3 24.383
R3236 a_3829_1050.n6 a_3829_1050.n4 23.684
R3237 a_3829_1050.n8 a_3829_1050.n0 16.08
R3238 a_3829_1050.n11 a_3829_1050.n10 16.078
R3239 a_3829_1050.n0 a_3829_1050.t2 14.282
R3240 a_3829_1050.n0 a_3829_1050.t3 14.282
R3241 a_3829_1050.n9 a_3829_1050.t6 14.282
R3242 a_3829_1050.n9 a_3829_1050.t5 14.282
R3243 a_3829_1050.t1 a_3829_1050.n11 14.282
R3244 a_3829_1050.n11 a_3829_1050.t0 14.282
R3245 a_7216_101.t0 a_7216_101.n1 34.62
R3246 a_7216_101.t0 a_7216_101.n0 8.137
R3247 a_7216_101.t0 a_7216_101.n2 4.69
R3248 a_91_103.n5 a_91_103.n4 19.724
R3249 a_91_103.t0 a_91_103.n3 11.595
R3250 a_91_103.t0 a_91_103.n5 9.207
R3251 a_91_103.n2 a_91_103.n1 2.455
R3252 a_91_103.n2 a_91_103.n0 1.32
R3253 a_91_103.t0 a_91_103.n2 0.246
R3254 a_5271_103.n5 a_5271_103.n4 19.724
R3255 a_5271_103.t0 a_5271_103.n3 11.595
R3256 a_5271_103.t0 a_5271_103.n5 9.207
R3257 a_5271_103.n2 a_5271_103.n1 2.455
R3258 a_5271_103.n2 a_5271_103.n0 1.32
R3259 a_5271_103.t0 a_5271_103.n2 0.246
R3260 a_3924_210.n10 a_3924_210.n8 82.852
R3261 a_3924_210.n7 a_3924_210.n6 32.833
R3262 a_3924_210.n8 a_3924_210.t1 32.416
R3263 a_3924_210.n10 a_3924_210.n9 27.2
R3264 a_3924_210.n11 a_3924_210.n0 23.498
R3265 a_3924_210.n3 a_3924_210.n2 23.284
R3266 a_3924_210.n11 a_3924_210.n10 22.4
R3267 a_3924_210.n7 a_3924_210.n4 19.017
R3268 a_3924_210.n6 a_3924_210.n5 13.494
R3269 a_3924_210.t1 a_3924_210.n1 7.04
R3270 a_3924_210.t1 a_3924_210.n3 5.727
R3271 a_3924_210.n8 a_3924_210.n7 1.435
R3272 a_13322_210.n9 a_13322_210.n7 82.852
R3273 a_13322_210.n3 a_13322_210.n1 44.628
R3274 a_13322_210.t0 a_13322_210.n9 32.417
R3275 a_13322_210.n7 a_13322_210.n6 27.2
R3276 a_13322_210.n5 a_13322_210.n4 23.498
R3277 a_13322_210.n3 a_13322_210.n2 23.284
R3278 a_13322_210.n7 a_13322_210.n5 22.4
R3279 a_13322_210.t0 a_13322_210.n11 20.241
R3280 a_13322_210.n11 a_13322_210.n10 13.494
R3281 a_13322_210.t0 a_13322_210.n0 8.137
R3282 a_13322_210.t0 a_13322_210.n3 5.727
R3283 a_13322_210.n9 a_13322_210.n8 1.435
R3284 a_14284_210.n10 a_14284_210.n8 82.852
R3285 a_14284_210.n7 a_14284_210.n6 32.833
R3286 a_14284_210.n8 a_14284_210.t1 32.416
R3287 a_14284_210.n10 a_14284_210.n9 27.2
R3288 a_14284_210.n11 a_14284_210.n0 23.498
R3289 a_14284_210.n3 a_14284_210.n2 23.284
R3290 a_14284_210.n11 a_14284_210.n10 22.4
R3291 a_14284_210.n7 a_14284_210.n4 19.017
R3292 a_14284_210.n6 a_14284_210.n5 13.494
R3293 a_14284_210.t1 a_14284_210.n1 7.04
R3294 a_14284_210.t1 a_14284_210.n3 5.727
R3295 a_14284_210.n8 a_14284_210.n7 1.435
R3296 a_13041_103.n5 a_13041_103.n4 19.724
R3297 a_13041_103.t0 a_13041_103.n3 11.595
R3298 a_13041_103.t0 a_13041_103.n5 9.207
R3299 a_13041_103.n2 a_13041_103.n1 2.455
R3300 a_13041_103.n2 a_13041_103.n0 1.32
R3301 a_13041_103.t0 a_13041_103.n2 0.246
R3302 a_3643_103.n1 a_3643_103.n0 25.576
R3303 a_3643_103.n3 a_3643_103.n2 9.111
R3304 a_3643_103.n7 a_3643_103.n6 2.455
R3305 a_3643_103.n5 a_3643_103.n3 1.964
R3306 a_3643_103.n5 a_3643_103.n4 1.964
R3307 a_3643_103.t0 a_3643_103.n1 1.871
R3308 a_3643_103.n7 a_3643_103.n5 0.636
R3309 a_3643_103.t0 a_3643_103.n7 0.246
R3310 a_4626_101.t0 a_4626_101.n1 34.62
R3311 a_4626_101.t0 a_4626_101.n0 8.137
R3312 a_4626_101.t0 a_4626_101.n2 4.69
R3313 a_14003_103.n5 a_14003_103.n4 19.724
R3314 a_14003_103.t0 a_14003_103.n3 11.595
R3315 a_14003_103.t0 a_14003_103.n5 9.207
R3316 a_14003_103.n2 a_14003_103.n1 2.455
R3317 a_14003_103.n2 a_14003_103.n0 1.32
R3318 a_14003_103.t0 a_14003_103.n2 0.246
R3319 a_2681_103.n5 a_2681_103.n4 19.724
R3320 a_2681_103.t0 a_2681_103.n3 11.595
R3321 a_2681_103.t0 a_2681_103.n5 9.207
R3322 a_2681_103.n2 a_2681_103.n1 2.455
R3323 a_2681_103.n2 a_2681_103.n0 1.32
R3324 a_2681_103.t0 a_2681_103.n2 0.246
R3325 a_1334_210.n9 a_1334_210.n7 82.852
R3326 a_1334_210.n3 a_1334_210.n1 44.628
R3327 a_1334_210.t0 a_1334_210.n9 32.417
R3328 a_1334_210.n7 a_1334_210.n6 27.2
R3329 a_1334_210.n5 a_1334_210.n4 23.498
R3330 a_1334_210.n3 a_1334_210.n2 23.284
R3331 a_1334_210.n7 a_1334_210.n5 22.4
R3332 a_1334_210.t0 a_1334_210.n11 20.241
R3333 a_1334_210.n11 a_1334_210.n10 13.494
R3334 a_1334_210.t0 a_1334_210.n0 8.137
R3335 a_1334_210.t0 a_1334_210.n3 5.727
R3336 a_1334_210.n9 a_1334_210.n8 1.435
R3337 a_1053_103.n1 a_1053_103.n0 25.576
R3338 a_1053_103.n3 a_1053_103.n2 9.111
R3339 a_1053_103.n7 a_1053_103.n6 2.455
R3340 a_1053_103.n5 a_1053_103.n3 1.964
R3341 a_1053_103.n5 a_1053_103.n4 1.964
R3342 a_1053_103.t0 a_1053_103.n1 1.871
R3343 a_1053_103.n7 a_1053_103.n5 0.636
R3344 a_1053_103.t0 a_1053_103.n7 0.246
C7 RN GND 10.14fF
C8 VDD GND 65.06fF
C9 a_1053_103.n0 GND 0.09fF
C10 a_1053_103.n1 GND 0.10fF
C11 a_1053_103.n2 GND 0.05fF
C12 a_1053_103.n3 GND 0.03fF
C13 a_1053_103.n4 GND 0.04fF
C14 a_1053_103.n5 GND 0.03fF
C15 a_1053_103.n6 GND 0.04fF
C16 a_1334_210.n0 GND 0.07fF
C17 a_1334_210.n1 GND 0.09fF
C18 a_1334_210.n2 GND 0.13fF
C19 a_1334_210.n3 GND 0.11fF
C20 a_1334_210.n4 GND 0.02fF
C21 a_1334_210.n5 GND 0.03fF
C22 a_1334_210.n6 GND 0.02fF
C23 a_1334_210.n7 GND 0.05fF
C24 a_1334_210.n8 GND 0.03fF
C25 a_1334_210.n9 GND 0.11fF
C26 a_1334_210.n10 GND 0.06fF
C27 a_1334_210.n11 GND 0.01fF
C28 a_1334_210.t0 GND 0.33fF
C29 a_2681_103.n0 GND 0.10fF
C30 a_2681_103.n1 GND 0.04fF
C31 a_2681_103.n2 GND 0.03fF
C32 a_2681_103.n3 GND 0.07fF
C33 a_2681_103.n4 GND 0.08fF
C34 a_2681_103.n5 GND 0.06fF
C35 a_14003_103.n0 GND 0.10fF
C36 a_14003_103.n1 GND 0.04fF
C37 a_14003_103.n2 GND 0.03fF
C38 a_14003_103.n3 GND 0.07fF
C39 a_14003_103.n4 GND 0.08fF
C40 a_14003_103.n5 GND 0.06fF
C41 a_4626_101.n0 GND 0.05fF
C42 a_4626_101.n1 GND 0.12fF
C43 a_4626_101.n2 GND 0.04fF
C44 a_3643_103.n0 GND 0.09fF
C45 a_3643_103.n1 GND 0.10fF
C46 a_3643_103.n2 GND 0.05fF
C47 a_3643_103.n3 GND 0.03fF
C48 a_3643_103.n4 GND 0.04fF
C49 a_3643_103.n5 GND 0.03fF
C50 a_3643_103.n6 GND 0.04fF
C51 a_13041_103.n0 GND 0.10fF
C52 a_13041_103.n1 GND 0.04fF
C53 a_13041_103.n2 GND 0.03fF
C54 a_13041_103.n3 GND 0.07fF
C55 a_13041_103.n4 GND 0.08fF
C56 a_13041_103.n5 GND 0.06fF
C57 a_14284_210.n0 GND 0.02fF
C58 a_14284_210.n1 GND 0.09fF
C59 a_14284_210.n2 GND 0.13fF
C60 a_14284_210.n3 GND 0.11fF
C61 a_14284_210.t1 GND 0.30fF
C62 a_14284_210.n4 GND 0.09fF
C63 a_14284_210.n5 GND 0.06fF
C64 a_14284_210.n6 GND 0.01fF
C65 a_14284_210.n7 GND 0.03fF
C66 a_14284_210.n8 GND 0.11fF
C67 a_14284_210.n9 GND 0.02fF
C68 a_14284_210.n10 GND 0.05fF
C69 a_14284_210.n11 GND 0.03fF
C70 a_13322_210.n0 GND 0.07fF
C71 a_13322_210.n1 GND 0.09fF
C72 a_13322_210.n2 GND 0.13fF
C73 a_13322_210.n3 GND 0.11fF
C74 a_13322_210.n4 GND 0.02fF
C75 a_13322_210.n5 GND 0.03fF
C76 a_13322_210.n6 GND 0.02fF
C77 a_13322_210.n7 GND 0.05fF
C78 a_13322_210.n8 GND 0.03fF
C79 a_13322_210.n9 GND 0.11fF
C80 a_13322_210.n10 GND 0.06fF
C81 a_13322_210.n11 GND 0.01fF
C82 a_13322_210.t0 GND 0.33fF
C83 a_3924_210.n0 GND 0.02fF
C84 a_3924_210.n1 GND 0.09fF
C85 a_3924_210.n2 GND 0.13fF
C86 a_3924_210.n3 GND 0.11fF
C87 a_3924_210.t1 GND 0.30fF
C88 a_3924_210.n4 GND 0.09fF
C89 a_3924_210.n5 GND 0.06fF
C90 a_3924_210.n6 GND 0.01fF
C91 a_3924_210.n7 GND 0.03fF
C92 a_3924_210.n8 GND 0.11fF
C93 a_3924_210.n9 GND 0.02fF
C94 a_3924_210.n10 GND 0.05fF
C95 a_3924_210.n11 GND 0.03fF
C96 a_5271_103.n0 GND 0.10fF
C97 a_5271_103.n1 GND 0.04fF
C98 a_5271_103.n2 GND 0.03fF
C99 a_5271_103.n3 GND 0.07fF
C100 a_5271_103.n4 GND 0.08fF
C101 a_5271_103.n5 GND 0.06fF
C102 a_91_103.n0 GND 0.10fF
C103 a_91_103.n1 GND 0.04fF
C104 a_91_103.n2 GND 0.03fF
C105 a_91_103.n3 GND 0.06fF
C106 a_91_103.n4 GND 0.08fF
C107 a_91_103.n5 GND 0.06fF
C108 a_7216_101.n0 GND 0.05fF
C109 a_7216_101.n1 GND 0.12fF
C110 a_7216_101.n2 GND 0.04fF
C111 a_3829_1050.n0 GND 0.50fF
C112 a_3829_1050.n1 GND 0.32fF
C113 a_3829_1050.n2 GND 0.54fF
C114 a_3829_1050.n3 GND 0.04fF
C115 a_3829_1050.n4 GND 0.05fF
C116 a_3829_1050.n5 GND 0.03fF
C117 a_3829_1050.n6 GND 0.31fF
C118 a_3829_1050.n7 GND 0.59fF
C119 a_3829_1050.n8 GND 0.26fF
C120 a_3829_1050.n9 GND 0.59fF
C121 a_3829_1050.n10 GND 0.19fF
C122 a_3829_1050.n11 GND 0.50fF
C123 a_9806_101.n0 GND 0.05fF
C124 a_9806_101.n1 GND 0.12fF
C125 a_9806_101.n2 GND 0.04fF
C126 a_8142_210.n0 GND 0.07fF
C127 a_8142_210.n1 GND 0.09fF
C128 a_8142_210.n2 GND 0.13fF
C129 a_8142_210.n3 GND 0.11fF
C130 a_8142_210.n4 GND 0.02fF
C131 a_8142_210.n5 GND 0.03fF
C132 a_8142_210.n6 GND 0.06fF
C133 a_8142_210.n7 GND 0.03fF
C134 a_8142_210.n8 GND 0.12fF
C135 a_8142_210.n9 GND 0.06fF
C136 a_8142_210.n10 GND 0.01fF
C137 a_8142_210.t0 GND 0.33fF
C138 a_7861_103.n0 GND 0.20fF
C139 a_7861_103.n1 GND 0.04fF
C140 a_7861_103.n2 GND 0.01fF
C141 a_7861_103.n3 GND 0.08fF
C142 a_7861_103.n4 GND 0.06fF
C143 a_7861_103.n5 GND 0.07fF
C144 a_2962_210.n0 GND 0.07fF
C145 a_2962_210.n1 GND 0.09fF
C146 a_2962_210.n2 GND 0.13fF
C147 a_2962_210.n3 GND 0.11fF
C148 a_2962_210.n4 GND 0.02fF
C149 a_2962_210.n5 GND 0.03fF
C150 a_2962_210.n6 GND 0.02fF
C151 a_2962_210.n7 GND 0.05fF
C152 a_2962_210.n8 GND 0.03fF
C153 a_2962_210.n9 GND 0.11fF
C154 a_2962_210.n10 GND 0.06fF
C155 a_2962_210.n11 GND 0.01fF
C156 a_2962_210.t0 GND 0.33fF
C157 a_16984_101.n0 GND 0.06fF
C158 a_16984_101.n1 GND 0.14fF
C159 a_16984_101.n2 GND 0.04fF
C160 a_5552_210.n0 GND 0.07fF
C161 a_5552_210.n1 GND 0.09fF
C162 a_5552_210.n2 GND 0.13fF
C163 a_5552_210.n3 GND 0.11fF
C164 a_5552_210.n4 GND 0.02fF
C165 a_5552_210.n5 GND 0.03fF
C166 a_5552_210.n6 GND 0.02fF
C167 a_5552_210.n7 GND 0.05fF
C168 a_5552_210.n8 GND 0.03fF
C169 a_5552_210.n9 GND 0.11fF
C170 a_5552_210.n10 GND 0.06fF
C171 a_5552_210.n11 GND 0.01fF
C172 a_5552_210.t0 GND 0.33fF
C173 a_6233_103.n0 GND 0.10fF
C174 a_6233_103.n1 GND 0.04fF
C175 a_6233_103.n2 GND 0.03fF
C176 a_6233_103.n3 GND 0.07fF
C177 a_6233_103.n4 GND 0.08fF
C178 a_6233_103.n5 GND 0.06fF
C179 a_10732_210.n0 GND 0.07fF
C180 a_10732_210.n1 GND 0.09fF
C181 a_10732_210.n2 GND 0.13fF
C182 a_10732_210.n3 GND 0.11fF
C183 a_10732_210.n4 GND 0.02fF
C184 a_10732_210.n5 GND 0.03fF
C185 a_10732_210.n6 GND 0.06fF
C186 a_10732_210.n7 GND 0.03fF
C187 a_10732_210.n8 GND 0.12fF
C188 a_10732_210.n9 GND 0.06fF
C189 a_10732_210.n10 GND 0.01fF
C190 a_10732_210.t0 GND 0.33fF
C191 a_372_210.n0 GND 0.07fF
C192 a_372_210.n1 GND 0.09fF
C193 a_372_210.n2 GND 0.13fF
C194 a_372_210.n3 GND 0.11fF
C195 a_372_210.n4 GND 0.02fF
C196 a_372_210.n5 GND 0.03fF
C197 a_372_210.n6 GND 0.02fF
C198 a_372_210.n7 GND 0.05fF
C199 a_372_210.n8 GND 0.03fF
C200 a_372_210.n9 GND 0.11fF
C201 a_372_210.n10 GND 0.06fF
C202 a_372_210.n11 GND 0.01fF
C203 a_372_210.t0 GND 0.33fF
C204 a_599_989.n0 GND 0.40fF
C205 a_599_989.n1 GND 0.43fF
C206 a_599_989.n2 GND 0.40fF
C207 a_599_989.t7 GND 0.57fF
C208 a_599_989.n3 GND 0.42fF
C209 a_599_989.n4 GND 1.34fF
C210 a_599_989.n5 GND 0.04fF
C211 a_599_989.n6 GND 0.06fF
C212 a_599_989.n7 GND 0.04fF
C213 a_599_989.n8 GND 0.32fF
C214 a_599_989.n9 GND 0.48fF
C215 a_599_989.n10 GND 0.58fF
C216 a_599_989.n11 GND 0.68fF
C217 a_599_989.n12 GND 0.21fF
C218 a_599_989.n13 GND 0.33fF
C219 a_599_989.n14 GND 0.58fF
C220 a_10637_1050.n0 GND 0.50fF
C221 a_10637_1050.n1 GND 0.98fF
C222 a_10637_1050.n2 GND 0.50fF
C223 a_10637_1050.n3 GND 0.78fF
C224 a_10637_1050.n4 GND 3.83fF
C225 a_10637_1050.n5 GND 0.07fF
C226 a_10637_1050.n6 GND 0.09fF
C227 a_10637_1050.n7 GND 0.06fF
C228 a_10637_1050.n8 GND 0.54fF
C229 a_10637_1050.n9 GND 0.74fF
C230 a_10637_1050.n10 GND 0.87fF
C231 a_10637_1050.n11 GND 1.02fF
C232 a_10637_1050.n12 GND 0.32fF
C233 a_10637_1050.n13 GND 0.45fF
C234 a_10637_1050.n14 GND 0.87fF
C235 a_16318_101.n0 GND 0.13fF
C236 a_16318_101.n1 GND 0.13fF
C237 a_277_1050.n0 GND 0.78fF
C238 a_277_1050.n1 GND 0.78fF
C239 a_277_1050.n2 GND 0.44fF
C240 a_277_1050.n3 GND 0.87fF
C241 a_277_1050.n4 GND 0.44fF
C242 a_277_1050.n5 GND 0.70fF
C243 a_277_1050.n6 GND 3.41fF
C244 a_277_1050.n7 GND 0.62fF
C245 a_277_1050.n8 GND 0.70fF
C246 a_277_1050.n9 GND 0.40fF
C247 a_277_1050.n10 GND 0.29fF
C248 a_277_1050.n11 GND 0.91fF
C249 a_9104_210.n0 GND 0.07fF
C250 a_9104_210.n1 GND 0.09fF
C251 a_9104_210.n2 GND 0.13fF
C252 a_9104_210.n3 GND 0.11fF
C253 a_9104_210.n4 GND 0.02fF
C254 a_9104_210.n5 GND 0.03fF
C255 a_9104_210.n6 GND 0.06fF
C256 a_9104_210.n7 GND 0.03fF
C257 a_9104_210.n8 GND 0.12fF
C258 a_9104_210.n9 GND 0.06fF
C259 a_9104_210.n10 GND 0.01fF
C260 a_9104_210.t0 GND 0.33fF
C261 a_8823_103.n0 GND 0.20fF
C262 a_8823_103.n1 GND 0.04fF
C263 a_8823_103.n2 GND 0.01fF
C264 a_8823_103.n3 GND 0.08fF
C265 a_8823_103.n4 GND 0.06fF
C266 a_8823_103.n5 GND 0.07fF
C267 a_12501_1050.n0 GND 0.60fF
C268 a_12501_1050.n1 GND 0.38fF
C269 a_12501_1050.n2 GND 0.75fF
C270 a_12501_1050.n3 GND 0.45fF
C271 a_12501_1050.n4 GND 0.72fF
C272 a_12501_1050.n5 GND 0.35fF
C273 a_12501_1050.n6 GND 0.71fF
C274 a_14986_101.n0 GND 0.05fF
C275 a_14986_101.n1 GND 0.12fF
C276 a_14986_101.n2 GND 0.04fF
C277 a_11694_210.n0 GND 0.07fF
C278 a_11694_210.n1 GND 0.09fF
C279 a_11694_210.n2 GND 0.13fF
C280 a_11694_210.n3 GND 0.11fF
C281 a_11694_210.n4 GND 0.02fF
C282 a_11694_210.n5 GND 0.03fF
C283 a_11694_210.n6 GND 0.06fF
C284 a_11694_210.n7 GND 0.03fF
C285 a_11694_210.n8 GND 0.12fF
C286 a_11694_210.n9 GND 0.06fF
C287 a_11694_210.n10 GND 0.01fF
C288 a_11694_210.t0 GND 0.33fF
C289 a_11413_103.n0 GND 0.09fF
C290 a_11413_103.n1 GND 0.10fF
C291 a_11413_103.n2 GND 0.05fF
C292 a_11413_103.n3 GND 0.03fF
C293 a_11413_103.n4 GND 0.04fF
C294 a_11413_103.n5 GND 0.11fF
C295 a_11413_103.n6 GND 0.04fF
C296 a_7321_1050.n0 GND 0.36fF
C297 a_7321_1050.n1 GND 0.70fF
C298 a_7321_1050.n2 GND 0.04fF
C299 a_7321_1050.n3 GND 0.06fF
C300 a_7321_1050.n4 GND 0.04fF
C301 a_7321_1050.n5 GND 0.32fF
C302 a_7321_1050.n6 GND 0.64fF
C303 a_7321_1050.n7 GND 0.67fF
C304 a_7321_1050.n8 GND 0.33fF
C305 a_7321_1050.n9 GND 0.56fF
C306 a_5327_187.n0 GND 0.46fF
C307 a_5327_187.t10 GND 0.98fF
C308 a_5327_187.n1 GND 0.70fF
C309 a_5327_187.n2 GND 0.46fF
C310 a_5327_187.t13 GND 0.98fF
C311 a_5327_187.n3 GND 0.63fF
C312 a_5327_187.n4 GND 0.45fF
C313 a_5327_187.n5 GND 0.94fF
C314 a_5327_187.n6 GND 3.49fF
C315 a_5327_187.n7 GND 2.75fF
C316 a_5327_187.n8 GND 0.07fF
C317 a_5327_187.n9 GND 0.09fF
C318 a_5327_187.n10 GND 0.06fF
C319 a_5327_187.n11 GND 0.60fF
C320 a_5327_187.n12 GND 0.75fF
C321 a_5327_187.n13 GND 0.89fF
C322 a_5327_187.n14 GND 1.05fF
C323 a_5327_187.n15 GND 0.33fF
C324 a_5327_187.n16 GND 0.41fF
C325 a_5327_187.n17 GND 0.89fF
C326 a_4151_989.n0 GND 0.92fF
C327 a_4151_989.n1 GND 1.06fF
C328 a_4151_989.n2 GND 1.30fF
C329 a_4151_989.t10 GND 0.98fF
C330 a_4151_989.n3 GND 0.74fF
C331 a_4151_989.n4 GND 4.56fF
C332 a_4151_989.n5 GND 0.98fF
C333 a_4151_989.t8 GND 1.07fF
C334 a_4151_989.n6 GND 0.83fF
C335 a_4151_989.n7 GND 19.06fF
C336 a_4151_989.n8 GND 0.09fF
C337 a_4151_989.n9 GND 0.12fF
C338 a_4151_989.n10 GND 0.08fF
C339 a_4151_989.n11 GND 0.53fF
C340 a_4151_989.n12 GND 0.96fF
C341 a_4151_989.n13 GND 1.40fF
C342 a_4151_989.n14 GND 0.82fF
C343 a_4151_989.n15 GND 1.19fF
C344 a_6514_210.n0 GND 0.07fF
C345 a_6514_210.n1 GND 0.09fF
C346 a_6514_210.n2 GND 0.13fF
C347 a_6514_210.n3 GND 0.11fF
C348 a_6514_210.n4 GND 0.02fF
C349 a_6514_210.n5 GND 0.03fF
C350 a_6514_210.n6 GND 0.06fF
C351 a_6514_210.n7 GND 0.03fF
C352 a_6514_210.n8 GND 0.12fF
C353 a_6514_210.n9 GND 0.06fF
C354 a_6514_210.n10 GND 0.01fF
C355 a_6514_210.t0 GND 0.33fF
C356 a_15652_101.n0 GND 0.02fF
C357 a_15652_101.n1 GND 0.09fF
C358 a_15652_101.n2 GND 0.05fF
C359 a_15652_101.n3 GND 0.06fF
C360 a_15652_101.n4 GND 0.00fF
C361 a_15652_101.n5 GND 0.04fF
C362 a_15652_101.n6 GND 0.05fF
C363 a_15652_101.n7 GND 0.02fF
C364 a_15652_101.n8 GND 0.05fF
C365 a_15652_101.n9 GND 0.09fF
C366 a_15652_101.n10 GND 0.21fF
C367 a_15652_101.n11 GND 0.07fF
C368 a_15652_101.t1 GND 0.14fF
C369 a_15652_101.n12 GND 0.04fF
C370 a_15652_101.n13 GND 0.00fF
C371 a_14189_1050.n0 GND 0.53fF
C372 a_14189_1050.n1 GND 0.34fF
C373 a_14189_1050.n2 GND 0.56fF
C374 a_14189_1050.n3 GND 0.04fF
C375 a_14189_1050.n4 GND 0.05fF
C376 a_14189_1050.n5 GND 0.03fF
C377 a_14189_1050.n6 GND 0.33fF
C378 a_14189_1050.n7 GND 0.61fF
C379 a_14189_1050.n8 GND 0.27fF
C380 a_14189_1050.n9 GND 0.62fF
C381 a_14189_1050.n10 GND 0.19fF
C382 a_14189_1050.n11 GND 0.53fF
C383 a_14511_989.n0 GND 0.30fF
C384 a_14511_989.n1 GND 0.34fF
C385 a_14511_989.t8 GND 0.64fF
C386 a_14511_989.n2 GND 1.07fF
C387 a_14511_989.n3 GND 0.76fF
C388 a_14511_989.t6 GND 0.58fF
C389 a_14511_989.n4 GND 0.35fF
C390 a_14511_989.n5 GND 0.41fF
C391 a_14511_989.t10 GND 0.58fF
C392 a_14511_989.n6 GND 0.42fF
C393 a_14511_989.n7 GND 1.24fF
C394 a_14511_989.n8 GND 0.04fF
C395 a_14511_989.n9 GND 0.06fF
C396 a_14511_989.n10 GND 0.04fF
C397 a_14511_989.n11 GND 0.33fF
C398 a_14511_989.n12 GND 0.46fF
C399 a_14511_989.n13 GND 0.69fF
C400 a_14511_989.n14 GND 0.34fF
C401 a_14511_989.n15 GND 0.58fF
C402 a_15757_1051.n0 GND 0.37fF
C403 a_15757_1051.n1 GND 0.33fF
C404 a_15757_1051.n2 GND 0.23fF
C405 a_15757_1051.n3 GND 0.62fF
C406 a_15757_1051.n4 GND 0.28fF
C407 a_15757_1051.n5 GND 0.41fF
C408 a_16421_1051.n0 GND 0.28fF
C409 a_16421_1051.n1 GND 0.29fF
C410 a_16421_1051.n2 GND 0.20fF
C411 a_16421_1051.n3 GND 0.57fF
C412 a_16421_1051.n4 GND 0.25fF
C413 a_16421_1051.n5 GND 0.35fF
C414 a_10451_103.n0 GND 0.20fF
C415 a_10451_103.n1 GND 0.04fF
C416 a_10451_103.n2 GND 0.01fF
C417 a_10451_103.n3 GND 0.08fF
C418 a_10451_103.n4 GND 0.06fF
C419 a_10451_103.n5 GND 0.07fF
C420 a_10507_187.n0 GND 0.44fF
C421 a_10507_187.t8 GND 0.93fF
C422 a_10507_187.n1 GND 0.67fF
C423 a_10507_187.n2 GND 0.44fF
C424 a_10507_187.t11 GND 0.93fF
C425 a_10507_187.n3 GND 0.60fF
C426 a_10507_187.n4 GND 0.43fF
C427 a_10507_187.n5 GND 0.89fF
C428 a_10507_187.n6 GND 3.31fF
C429 a_10507_187.n7 GND 2.61fF
C430 a_10507_187.n8 GND 0.06fF
C431 a_10507_187.n9 GND 0.08fF
C432 a_10507_187.n10 GND 0.05fF
C433 a_10507_187.n11 GND 0.57fF
C434 a_10507_187.n12 GND 0.71fF
C435 a_10507_187.n13 GND 0.84fF
C436 a_10507_187.n14 GND 0.99fF
C437 a_10507_187.n15 GND 0.31fF
C438 a_10507_187.n16 GND 0.38fF
C439 a_10507_187.n17 GND 0.84fF
C440 a_5457_1050.n0 GND 0.48fF
C441 a_5457_1050.n1 GND 0.94fF
C442 a_5457_1050.n2 GND 0.48fF
C443 a_5457_1050.n3 GND 0.76fF
C444 a_5457_1050.n4 GND 3.70fF
C445 a_5457_1050.n5 GND 0.06fF
C446 a_5457_1050.n6 GND 0.08fF
C447 a_5457_1050.n7 GND 0.05fF
C448 a_5457_1050.n8 GND 0.52fF
C449 a_5457_1050.n9 GND 0.71fF
C450 a_5457_1050.n10 GND 0.84fF
C451 a_5457_1050.n11 GND 0.99fF
C452 a_5457_1050.n12 GND 0.31fF
C453 a_5457_1050.n13 GND 0.43fF
C454 a_5457_1050.n14 GND 0.84fF
C455 Q.n0 GND 0.75fF
C456 Q.n1 GND 0.45fF
C457 Q.n2 GND 0.51fF
C458 Q.n3 GND 0.01fF
C459 a_15932_209.n0 GND 0.38fF
C460 a_15932_209.n1 GND 0.46fF
C461 a_15932_209.n2 GND 0.23fF
C462 a_15932_209.n3 GND 0.26fF
C463 a_15932_209.n4 GND 0.48fF
C464 a_15932_209.n5 GND 0.45fF
C465 a_15932_209.n6 GND 0.04fF
C466 a_15932_209.n7 GND 0.04fF
C467 a_15932_209.n8 GND 0.10fF
C468 a_15932_209.n9 GND 0.04fF
C469 a_15932_209.n10 GND 0.04fF
C470 a_15932_209.n11 GND 0.10fF
C471 a_15932_209.n12 GND 0.99fF
C472 a_15932_209.n13 GND 0.27fF
C473 a_15932_209.n14 GND 0.07fF
C474 a_15932_209.n15 GND 0.04fF
C475 a_15932_209.n16 GND 0.04fF
C476 a_2141_1050.n0 GND 0.34fF
C477 a_2141_1050.n1 GND 0.67fF
C478 a_2141_1050.n2 GND 0.40fF
C479 a_2141_1050.n3 GND 0.64fF
C480 a_2141_1050.n4 GND 0.64fF
C481 a_2141_1050.n5 GND 0.31fF
C482 a_2141_1050.n6 GND 0.54fF
C483 a_2036_101.n0 GND 0.05fF
C484 a_2036_101.n1 GND 0.12fF
C485 a_2036_101.n2 GND 0.04fF
C486 a_147_187.n0 GND 0.42fF
C487 a_147_187.t15 GND 0.90fF
C488 a_147_187.n1 GND 0.65fF
C489 a_147_187.n2 GND 0.42fF
C490 a_147_187.t7 GND 0.90fF
C491 a_147_187.n3 GND 0.58fF
C492 a_147_187.n4 GND 0.42fF
C493 a_147_187.n5 GND 0.87fF
C494 a_147_187.n6 GND 3.22fF
C495 a_147_187.n7 GND 2.54fF
C496 a_147_187.n8 GND 0.06fF
C497 a_147_187.n9 GND 0.08fF
C498 a_147_187.n10 GND 0.05fF
C499 a_147_187.n11 GND 0.56fF
C500 a_147_187.n12 GND 0.69fF
C501 a_147_187.n13 GND 0.82fF
C502 a_147_187.n14 GND 0.96fF
C503 a_147_187.n15 GND 0.30fF
C504 a_147_187.n16 GND 0.37fF
C505 a_147_187.n17 GND 0.82fF
C506 a_9009_1050.n0 GND 0.34fF
C507 a_9009_1050.n1 GND 0.56fF
C508 a_9009_1050.n2 GND 0.04fF
C509 a_9009_1050.n3 GND 0.05fF
C510 a_9009_1050.n4 GND 0.03fF
C511 a_9009_1050.n5 GND 0.33fF
C512 a_9009_1050.n6 GND 0.61fF
C513 a_9009_1050.n7 GND 0.53fF
C514 a_9009_1050.n8 GND 0.62fF
C515 a_9009_1050.n9 GND 0.19fF
C516 a_9009_1050.n10 GND 0.27fF
C517 a_9009_1050.n11 GND 0.53fF
C518 a_9331_989.n0 GND 1.05fF
C519 a_9331_989.n1 GND 1.25fF
C520 a_9331_989.n2 GND 0.67fF
C521 a_9331_989.n3 GND 0.55fF
C522 a_9331_989.n4 GND 1.47fF
C523 a_9331_989.n5 GND 0.49fF
C524 a_9331_989.n6 GND 1.11fF
C525 a_9331_989.n7 GND 1.66fF
C526 a_9331_989.n8 GND 0.81fF
C527 a_9331_989.t12 GND 1.00fF
C528 a_9331_989.n9 GND 0.75fF
C529 a_9331_989.n10 GND 9.37fF
C530 a_9331_989.n11 GND 0.87fF
C531 a_9331_989.n12 GND 0.17fF
C532 a_9331_989.n13 GND 0.51fF
C533 a_9331_989.n14 GND 0.09fF
C534 a_5779_989.n0 GND 0.46fF
C535 a_5779_989.n1 GND 0.48fF
C536 a_5779_989.n2 GND 0.46fF
C537 a_5779_989.t8 GND 0.65fF
C538 a_5779_989.n3 GND 0.48fF
C539 a_5779_989.n4 GND 1.51fF
C540 a_5779_989.n5 GND 0.05fF
C541 a_5779_989.n6 GND 0.07fF
C542 a_5779_989.n7 GND 0.04fF
C543 a_5779_989.n8 GND 0.37fF
C544 a_5779_989.n9 GND 0.55fF
C545 a_5779_989.n10 GND 0.65fF
C546 a_5779_989.n11 GND 0.76fF
C547 a_5779_989.n12 GND 0.24fF
C548 a_5779_989.n13 GND 0.37fF
C549 a_5779_989.n14 GND 0.65fF
C550 VDD.n0 GND 0.12fF
C551 VDD.n1 GND 0.03fF
C552 VDD.n2 GND 0.02fF
C553 VDD.n3 GND 0.05fF
C554 VDD.n4 GND 0.01fF
C555 VDD.n5 GND 0.02fF
C556 VDD.n6 GND 0.02fF
C557 VDD.n9 GND 0.02fF
C558 VDD.n10 GND 0.02fF
C559 VDD.n12 GND 0.02fF
C560 VDD.n14 GND 0.46fF
C561 VDD.n16 GND 0.03fF
C562 VDD.n17 GND 0.02fF
C563 VDD.n18 GND 0.02fF
C564 VDD.n19 GND 0.02fF
C565 VDD.n20 GND 0.04fF
C566 VDD.n21 GND 0.27fF
C567 VDD.n22 GND 0.02fF
C568 VDD.n23 GND 0.03fF
C569 VDD.n24 GND 0.06fF
C570 VDD.n25 GND 0.15fF
C571 VDD.n26 GND 0.20fF
C572 VDD.n27 GND 0.01fF
C573 VDD.n28 GND 0.01fF
C574 VDD.n29 GND 0.07fF
C575 VDD.n30 GND 0.17fF
C576 VDD.n31 GND 0.01fF
C577 VDD.n32 GND 0.02fF
C578 VDD.n33 GND 0.02fF
C579 VDD.n34 GND 0.15fF
C580 VDD.n35 GND 0.20fF
C581 VDD.n36 GND 0.01fF
C582 VDD.n37 GND 0.06fF
C583 VDD.n38 GND 0.01fF
C584 VDD.n39 GND 0.02fF
C585 VDD.n40 GND 0.27fF
C586 VDD.n41 GND 0.01fF
C587 VDD.n42 GND 0.02fF
C588 VDD.n43 GND 0.03fF
C589 VDD.n44 GND 0.02fF
C590 VDD.n45 GND 0.02fF
C591 VDD.n46 GND 0.02fF
C592 VDD.n47 GND 0.18fF
C593 VDD.n48 GND 0.04fF
C594 VDD.n49 GND 0.04fF
C595 VDD.n50 GND 0.02fF
C596 VDD.n52 GND 0.02fF
C597 VDD.n53 GND 0.02fF
C598 VDD.n54 GND 0.02fF
C599 VDD.n55 GND 0.02fF
C600 VDD.n57 GND 0.02fF
C601 VDD.n58 GND 0.02fF
C602 VDD.n59 GND 0.02fF
C603 VDD.n61 GND 0.27fF
C604 VDD.n63 GND 0.02fF
C605 VDD.n64 GND 0.02fF
C606 VDD.n65 GND 0.03fF
C607 VDD.n66 GND 0.02fF
C608 VDD.n67 GND 0.27fF
C609 VDD.n68 GND 0.01fF
C610 VDD.n69 GND 0.02fF
C611 VDD.n70 GND 0.03fF
C612 VDD.n71 GND 0.27fF
C613 VDD.n72 GND 0.01fF
C614 VDD.n73 GND 0.02fF
C615 VDD.n74 GND 0.02fF
C616 VDD.n75 GND 0.27fF
C617 VDD.n76 GND 0.01fF
C618 VDD.n77 GND 0.02fF
C619 VDD.n78 GND 0.02fF
C620 VDD.n79 GND 0.31fF
C621 VDD.n80 GND 0.01fF
C622 VDD.n81 GND 0.03fF
C623 VDD.n82 GND 0.03fF
C624 VDD.n83 GND 0.31fF
C625 VDD.n84 GND 0.01fF
C626 VDD.n85 GND 0.03fF
C627 VDD.n86 GND 0.03fF
C628 VDD.n87 GND 0.27fF
C629 VDD.n88 GND 0.01fF
C630 VDD.n89 GND 0.02fF
C631 VDD.n90 GND 0.02fF
C632 VDD.n91 GND 0.27fF
C633 VDD.n92 GND 0.01fF
C634 VDD.n93 GND 0.02fF
C635 VDD.n94 GND 0.02fF
C636 VDD.n95 GND 0.27fF
C637 VDD.n96 GND 0.01fF
C638 VDD.n97 GND 0.02fF
C639 VDD.n98 GND 0.03fF
C640 VDD.n99 GND 0.02fF
C641 VDD.n100 GND 0.02fF
C642 VDD.n101 GND 0.02fF
C643 VDD.n102 GND 0.22fF
C644 VDD.n103 GND 0.04fF
C645 VDD.n104 GND 0.03fF
C646 VDD.n105 GND 0.02fF
C647 VDD.n106 GND 0.02fF
C648 VDD.n107 GND 0.02fF
C649 VDD.n108 GND 0.03fF
C650 VDD.n109 GND 0.02fF
C651 VDD.n111 GND 0.02fF
C652 VDD.n112 GND 0.02fF
C653 VDD.n113 GND 0.02fF
C654 VDD.n115 GND 0.27fF
C655 VDD.n117 GND 0.02fF
C656 VDD.n118 GND 0.02fF
C657 VDD.n119 GND 0.03fF
C658 VDD.n120 GND 0.02fF
C659 VDD.n121 GND 0.27fF
C660 VDD.n122 GND 0.01fF
C661 VDD.n123 GND 0.02fF
C662 VDD.n124 GND 0.03fF
C663 VDD.n125 GND 0.27fF
C664 VDD.n126 GND 0.01fF
C665 VDD.n127 GND 0.02fF
C666 VDD.n128 GND 0.02fF
C667 VDD.n129 GND 0.27fF
C668 VDD.n130 GND 0.01fF
C669 VDD.n131 GND 0.02fF
C670 VDD.n132 GND 0.02fF
C671 VDD.n133 GND 0.31fF
C672 VDD.n134 GND 0.01fF
C673 VDD.n135 GND 0.03fF
C674 VDD.n136 GND 0.03fF
C675 VDD.n137 GND 0.31fF
C676 VDD.n138 GND 0.01fF
C677 VDD.n139 GND 0.03fF
C678 VDD.n140 GND 0.03fF
C679 VDD.n141 GND 0.27fF
C680 VDD.n142 GND 0.01fF
C681 VDD.n143 GND 0.02fF
C682 VDD.n144 GND 0.02fF
C683 VDD.n145 GND 0.27fF
C684 VDD.n146 GND 0.01fF
C685 VDD.n147 GND 0.02fF
C686 VDD.n148 GND 0.02fF
C687 VDD.n149 GND 0.27fF
C688 VDD.n150 GND 0.01fF
C689 VDD.n151 GND 0.02fF
C690 VDD.n152 GND 0.03fF
C691 VDD.n153 GND 0.02fF
C692 VDD.n154 GND 0.02fF
C693 VDD.n155 GND 0.02fF
C694 VDD.n156 GND 0.22fF
C695 VDD.n157 GND 0.04fF
C696 VDD.n158 GND 0.03fF
C697 VDD.n159 GND 0.02fF
C698 VDD.n160 GND 0.02fF
C699 VDD.n161 GND 0.02fF
C700 VDD.n162 GND 0.03fF
C701 VDD.n163 GND 0.02fF
C702 VDD.n165 GND 0.02fF
C703 VDD.n166 GND 0.02fF
C704 VDD.n167 GND 0.02fF
C705 VDD.n169 GND 0.27fF
C706 VDD.n171 GND 0.02fF
C707 VDD.n172 GND 0.02fF
C708 VDD.n173 GND 0.03fF
C709 VDD.n174 GND 0.02fF
C710 VDD.n175 GND 0.27fF
C711 VDD.n176 GND 0.01fF
C712 VDD.n177 GND 0.02fF
C713 VDD.n178 GND 0.03fF
C714 VDD.n179 GND 0.06fF
C715 VDD.n180 GND 0.24fF
C716 VDD.n181 GND 0.01fF
C717 VDD.n182 GND 0.01fF
C718 VDD.n183 GND 0.02fF
C719 VDD.n184 GND 0.14fF
C720 VDD.n185 GND 0.17fF
C721 VDD.n186 GND 0.01fF
C722 VDD.n187 GND 0.02fF
C723 VDD.n188 GND 0.02fF
C724 VDD.n189 GND 0.11fF
C725 VDD.n190 GND 0.03fF
C726 VDD.n191 GND 0.31fF
C727 VDD.n192 GND 0.01fF
C728 VDD.n193 GND 0.02fF
C729 VDD.n194 GND 0.03fF
C730 VDD.n195 GND 0.17fF
C731 VDD.n196 GND 0.14fF
C732 VDD.n197 GND 0.01fF
C733 VDD.n198 GND 0.02fF
C734 VDD.n199 GND 0.03fF
C735 VDD.n200 GND 0.14fF
C736 VDD.n201 GND 0.16fF
C737 VDD.n202 GND 0.01fF
C738 VDD.n203 GND 0.02fF
C739 VDD.n204 GND 0.02fF
C740 VDD.n205 GND 0.06fF
C741 VDD.n206 GND 0.25fF
C742 VDD.n207 GND 0.01fF
C743 VDD.n208 GND 0.01fF
C744 VDD.n209 GND 0.02fF
C745 VDD.n210 GND 0.27fF
C746 VDD.n211 GND 0.01fF
C747 VDD.n212 GND 0.02fF
C748 VDD.n213 GND 0.03fF
C749 VDD.n214 GND 0.02fF
C750 VDD.n215 GND 0.02fF
C751 VDD.n216 GND 0.02fF
C752 VDD.n217 GND 0.22fF
C753 VDD.n218 GND 0.04fF
C754 VDD.n219 GND 0.03fF
C755 VDD.n220 GND 0.02fF
C756 VDD.n221 GND 0.02fF
C757 VDD.n222 GND 0.02fF
C758 VDD.n223 GND 0.03fF
C759 VDD.n224 GND 0.02fF
C760 VDD.n226 GND 0.02fF
C761 VDD.n227 GND 0.02fF
C762 VDD.n228 GND 0.02fF
C763 VDD.n230 GND 0.27fF
C764 VDD.n232 GND 0.02fF
C765 VDD.n233 GND 0.02fF
C766 VDD.n234 GND 0.03fF
C767 VDD.n235 GND 0.02fF
C768 VDD.n236 GND 0.27fF
C769 VDD.n237 GND 0.01fF
C770 VDD.n238 GND 0.02fF
C771 VDD.n239 GND 0.03fF
C772 VDD.n240 GND 0.06fF
C773 VDD.n241 GND 0.24fF
C774 VDD.n242 GND 0.01fF
C775 VDD.n243 GND 0.01fF
C776 VDD.n244 GND 0.02fF
C777 VDD.n245 GND 0.14fF
C778 VDD.n246 GND 0.17fF
C779 VDD.n247 GND 0.01fF
C780 VDD.n248 GND 0.02fF
C781 VDD.n249 GND 0.02fF
C782 VDD.n250 GND 0.11fF
C783 VDD.n251 GND 0.03fF
C784 VDD.n252 GND 0.31fF
C785 VDD.n253 GND 0.01fF
C786 VDD.n254 GND 0.02fF
C787 VDD.n255 GND 0.03fF
C788 VDD.n256 GND 0.17fF
C789 VDD.n257 GND 0.14fF
C790 VDD.n258 GND 0.01fF
C791 VDD.n259 GND 0.02fF
C792 VDD.n260 GND 0.03fF
C793 VDD.n261 GND 0.14fF
C794 VDD.n262 GND 0.16fF
C795 VDD.n263 GND 0.01fF
C796 VDD.n264 GND 0.02fF
C797 VDD.n265 GND 0.02fF
C798 VDD.n266 GND 0.06fF
C799 VDD.n267 GND 0.25fF
C800 VDD.n268 GND 0.01fF
C801 VDD.n269 GND 0.01fF
C802 VDD.n270 GND 0.02fF
C803 VDD.n271 GND 0.27fF
C804 VDD.n272 GND 0.01fF
C805 VDD.n273 GND 0.02fF
C806 VDD.n274 GND 0.03fF
C807 VDD.n275 GND 0.02fF
C808 VDD.n276 GND 0.02fF
C809 VDD.n277 GND 0.02fF
C810 VDD.n278 GND 0.26fF
C811 VDD.n279 GND 0.04fF
C812 VDD.n280 GND 0.03fF
C813 VDD.n281 GND 0.02fF
C814 VDD.n282 GND 0.02fF
C815 VDD.n283 GND 0.02fF
C816 VDD.n284 GND 0.03fF
C817 VDD.n285 GND 0.02fF
C818 VDD.n287 GND 0.02fF
C819 VDD.n288 GND 0.02fF
C820 VDD.n289 GND 0.02fF
C821 VDD.n291 GND 0.27fF
C822 VDD.n293 GND 0.02fF
C823 VDD.n294 GND 0.02fF
C824 VDD.n295 GND 0.03fF
C825 VDD.n296 GND 0.02fF
C826 VDD.n297 GND 0.27fF
C827 VDD.n298 GND 0.01fF
C828 VDD.n299 GND 0.02fF
C829 VDD.n300 GND 0.03fF
C830 VDD.n301 GND 0.27fF
C831 VDD.n302 GND 0.01fF
C832 VDD.n303 GND 0.02fF
C833 VDD.n304 GND 0.02fF
C834 VDD.n305 GND 0.22fF
C835 VDD.n306 GND 0.01fF
C836 VDD.n307 GND 0.07fF
C837 VDD.n308 GND 0.02fF
C838 VDD.n309 GND 0.14fF
C839 VDD.n310 GND 0.17fF
C840 VDD.n311 GND 0.01fF
C841 VDD.n312 GND 0.02fF
C842 VDD.n313 GND 0.02fF
C843 VDD.n314 GND 0.14fF
C844 VDD.n315 GND 0.16fF
C845 VDD.n316 GND 0.01fF
C846 VDD.n317 GND 0.11fF
C847 VDD.n318 GND 0.02fF
C848 VDD.n319 GND 0.02fF
C849 VDD.n320 GND 0.02fF
C850 VDD.n321 GND 0.18fF
C851 VDD.n322 GND 0.15fF
C852 VDD.n323 GND 0.01fF
C853 VDD.n324 GND 0.02fF
C854 VDD.n325 GND 0.03fF
C855 VDD.n326 GND 0.18fF
C856 VDD.n327 GND 0.15fF
C857 VDD.n328 GND 0.01fF
C858 VDD.n329 GND 0.02fF
C859 VDD.n330 GND 0.03fF
C860 VDD.n331 GND 0.11fF
C861 VDD.n332 GND 0.02fF
C862 VDD.n333 GND 0.14fF
C863 VDD.n334 GND 0.16fF
C864 VDD.n335 GND 0.01fF
C865 VDD.n336 GND 0.02fF
C866 VDD.n337 GND 0.02fF
C867 VDD.n338 GND 0.14fF
C868 VDD.n339 GND 0.17fF
C869 VDD.n340 GND 0.01fF
C870 VDD.n341 GND 0.02fF
C871 VDD.n342 GND 0.02fF
C872 VDD.n343 GND 0.06fF
C873 VDD.n344 GND 0.23fF
C874 VDD.n345 GND 0.01fF
C875 VDD.n346 GND 0.01fF
C876 VDD.n347 GND 0.02fF
C877 VDD.n348 GND 0.27fF
C878 VDD.n349 GND 0.01fF
C879 VDD.n350 GND 0.02fF
C880 VDD.n351 GND 0.02fF
C881 VDD.n352 GND 0.27fF
C882 VDD.n353 GND 0.01fF
C883 VDD.n354 GND 0.02fF
C884 VDD.n355 GND 0.03fF
C885 VDD.n356 GND 0.02fF
C886 VDD.n357 GND 0.02fF
C887 VDD.n358 GND 0.02fF
C888 VDD.n359 GND 0.31fF
C889 VDD.n360 GND 0.04fF
C890 VDD.n361 GND 0.03fF
C891 VDD.n362 GND 0.02fF
C892 VDD.n363 GND 0.02fF
C893 VDD.n364 GND 0.02fF
C894 VDD.n365 GND 0.03fF
C895 VDD.n366 GND 0.02fF
C896 VDD.n368 GND 0.02fF
C897 VDD.n369 GND 0.02fF
C898 VDD.n370 GND 0.02fF
C899 VDD.n372 GND 0.27fF
C900 VDD.n374 GND 0.02fF
C901 VDD.n375 GND 0.02fF
C902 VDD.n376 GND 0.03fF
C903 VDD.n377 GND 0.02fF
C904 VDD.n378 GND 0.27fF
C905 VDD.n379 GND 0.01fF
C906 VDD.n380 GND 0.02fF
C907 VDD.n381 GND 0.03fF
C908 VDD.n382 GND 0.27fF
C909 VDD.n383 GND 0.01fF
C910 VDD.n384 GND 0.02fF
C911 VDD.n385 GND 0.02fF
C912 VDD.n386 GND 0.22fF
C913 VDD.n387 GND 0.01fF
C914 VDD.n388 GND 0.07fF
C915 VDD.n389 GND 0.02fF
C916 VDD.n390 GND 0.14fF
C917 VDD.n391 GND 0.17fF
C918 VDD.n392 GND 0.01fF
C919 VDD.n393 GND 0.02fF
C920 VDD.n394 GND 0.02fF
C921 VDD.n395 GND 0.14fF
C922 VDD.n396 GND 0.16fF
C923 VDD.n397 GND 0.01fF
C924 VDD.n398 GND 0.11fF
C925 VDD.n399 GND 0.02fF
C926 VDD.n400 GND 0.02fF
C927 VDD.n401 GND 0.02fF
C928 VDD.n402 GND 0.18fF
C929 VDD.n403 GND 0.15fF
C930 VDD.n404 GND 0.01fF
C931 VDD.n405 GND 0.02fF
C932 VDD.n406 GND 0.03fF
C933 VDD.n407 GND 0.18fF
C934 VDD.n408 GND 0.15fF
C935 VDD.n409 GND 0.01fF
C936 VDD.n410 GND 0.02fF
C937 VDD.n411 GND 0.03fF
C938 VDD.n412 GND 0.11fF
C939 VDD.n413 GND 0.02fF
C940 VDD.n414 GND 0.14fF
C941 VDD.n415 GND 0.16fF
C942 VDD.n416 GND 0.01fF
C943 VDD.n417 GND 0.02fF
C944 VDD.n418 GND 0.02fF
C945 VDD.n419 GND 0.14fF
C946 VDD.n420 GND 0.17fF
C947 VDD.n421 GND 0.01fF
C948 VDD.n422 GND 0.02fF
C949 VDD.n423 GND 0.02fF
C950 VDD.n424 GND 0.06fF
C951 VDD.n425 GND 0.23fF
C952 VDD.n426 GND 0.01fF
C953 VDD.n427 GND 0.01fF
C954 VDD.n428 GND 0.02fF
C955 VDD.n429 GND 0.27fF
C956 VDD.n430 GND 0.01fF
C957 VDD.n431 GND 0.02fF
C958 VDD.n432 GND 0.02fF
C959 VDD.n433 GND 0.27fF
C960 VDD.n434 GND 0.01fF
C961 VDD.n435 GND 0.02fF
C962 VDD.n436 GND 0.03fF
C963 VDD.n437 GND 0.02fF
C964 VDD.n438 GND 0.02fF
C965 VDD.n439 GND 0.02fF
C966 VDD.n440 GND 0.26fF
C967 VDD.n441 GND 0.04fF
C968 VDD.n442 GND 0.03fF
C969 VDD.n443 GND 0.02fF
C970 VDD.n444 GND 0.02fF
C971 VDD.n445 GND 0.02fF
C972 VDD.n446 GND 0.03fF
C973 VDD.n447 GND 0.02fF
C974 VDD.n449 GND 0.02fF
C975 VDD.n450 GND 0.02fF
C976 VDD.n451 GND 0.02fF
C977 VDD.n453 GND 0.27fF
C978 VDD.n455 GND 0.02fF
C979 VDD.n456 GND 0.02fF
C980 VDD.n457 GND 0.03fF
C981 VDD.n458 GND 0.02fF
C982 VDD.n459 GND 0.27fF
C983 VDD.n460 GND 0.01fF
C984 VDD.n461 GND 0.02fF
C985 VDD.n462 GND 0.03fF
C986 VDD.n463 GND 0.06fF
C987 VDD.n464 GND 0.24fF
C988 VDD.n465 GND 0.01fF
C989 VDD.n466 GND 0.01fF
C990 VDD.n467 GND 0.02fF
C991 VDD.n468 GND 0.14fF
C992 VDD.n469 GND 0.17fF
C993 VDD.n470 GND 0.01fF
C994 VDD.n471 GND 0.02fF
C995 VDD.n472 GND 0.02fF
C996 VDD.n473 GND 0.11fF
C997 VDD.n474 GND 0.03fF
C998 VDD.n475 GND 0.31fF
C999 VDD.n476 GND 0.01fF
C1000 VDD.n477 GND 0.02fF
C1001 VDD.n478 GND 0.03fF
C1002 VDD.n479 GND 0.17fF
C1003 VDD.n480 GND 0.14fF
C1004 VDD.n481 GND 0.01fF
C1005 VDD.n482 GND 0.02fF
C1006 VDD.n483 GND 0.03fF
C1007 VDD.n484 GND 0.14fF
C1008 VDD.n485 GND 0.16fF
C1009 VDD.n486 GND 0.01fF
C1010 VDD.n487 GND 0.02fF
C1011 VDD.n488 GND 0.02fF
C1012 VDD.n489 GND 0.06fF
C1013 VDD.n490 GND 0.25fF
C1014 VDD.n491 GND 0.01fF
C1015 VDD.n492 GND 0.01fF
C1016 VDD.n493 GND 0.02fF
C1017 VDD.n494 GND 0.27fF
C1018 VDD.n495 GND 0.01fF
C1019 VDD.n496 GND 0.02fF
C1020 VDD.n497 GND 0.03fF
C1021 VDD.n498 GND 0.02fF
C1022 VDD.n499 GND 0.02fF
C1023 VDD.n500 GND 0.02fF
C1024 VDD.n501 GND 0.26fF
C1025 VDD.n502 GND 0.04fF
C1026 VDD.n503 GND 0.03fF
C1027 VDD.n504 GND 0.02fF
C1028 VDD.n505 GND 0.02fF
C1029 VDD.n506 GND 0.02fF
C1030 VDD.n507 GND 0.03fF
C1031 VDD.n508 GND 0.02fF
C1032 VDD.n510 GND 0.02fF
C1033 VDD.n511 GND 0.02fF
C1034 VDD.n512 GND 0.02fF
C1035 VDD.n514 GND 0.27fF
C1036 VDD.n516 GND 0.02fF
C1037 VDD.n517 GND 0.02fF
C1038 VDD.n518 GND 0.03fF
C1039 VDD.n519 GND 0.02fF
C1040 VDD.n520 GND 0.27fF
C1041 VDD.n521 GND 0.01fF
C1042 VDD.n522 GND 0.02fF
C1043 VDD.n523 GND 0.03fF
C1044 VDD.n524 GND 0.27fF
C1045 VDD.n525 GND 0.01fF
C1046 VDD.n526 GND 0.02fF
C1047 VDD.n527 GND 0.02fF
C1048 VDD.n528 GND 0.22fF
C1049 VDD.n529 GND 0.01fF
C1050 VDD.n530 GND 0.07fF
C1051 VDD.n531 GND 0.02fF
C1052 VDD.n532 GND 0.14fF
C1053 VDD.n533 GND 0.17fF
C1054 VDD.n534 GND 0.01fF
C1055 VDD.n535 GND 0.02fF
C1056 VDD.n536 GND 0.02fF
C1057 VDD.n537 GND 0.14fF
C1058 VDD.n538 GND 0.16fF
C1059 VDD.n539 GND 0.01fF
C1060 VDD.n540 GND 0.11fF
C1061 VDD.n541 GND 0.02fF
C1062 VDD.n542 GND 0.02fF
C1063 VDD.n543 GND 0.02fF
C1064 VDD.n544 GND 0.18fF
C1065 VDD.n545 GND 0.15fF
C1066 VDD.n546 GND 0.01fF
C1067 VDD.n547 GND 0.02fF
C1068 VDD.n548 GND 0.03fF
C1069 VDD.n549 GND 0.18fF
C1070 VDD.n550 GND 0.15fF
C1071 VDD.n551 GND 0.01fF
C1072 VDD.n552 GND 0.02fF
C1073 VDD.n553 GND 0.03fF
C1074 VDD.n554 GND 0.11fF
C1075 VDD.n555 GND 0.02fF
C1076 VDD.n556 GND 0.14fF
C1077 VDD.n557 GND 0.16fF
C1078 VDD.n558 GND 0.01fF
C1079 VDD.n559 GND 0.02fF
C1080 VDD.n560 GND 0.02fF
C1081 VDD.n561 GND 0.14fF
C1082 VDD.n562 GND 0.17fF
C1083 VDD.n563 GND 0.01fF
C1084 VDD.n564 GND 0.02fF
C1085 VDD.n565 GND 0.02fF
C1086 VDD.n566 GND 0.06fF
C1087 VDD.n567 GND 0.23fF
C1088 VDD.n568 GND 0.01fF
C1089 VDD.n569 GND 0.01fF
C1090 VDD.n570 GND 0.02fF
C1091 VDD.n571 GND 0.27fF
C1092 VDD.n572 GND 0.01fF
C1093 VDD.n573 GND 0.02fF
C1094 VDD.n574 GND 0.02fF
C1095 VDD.n575 GND 0.27fF
C1096 VDD.n576 GND 0.01fF
C1097 VDD.n577 GND 0.02fF
C1098 VDD.n578 GND 0.03fF
C1099 VDD.n579 GND 0.02fF
C1100 VDD.n580 GND 0.02fF
C1101 VDD.n581 GND 0.02fF
C1102 VDD.n582 GND 0.31fF
C1103 VDD.n583 GND 0.04fF
C1104 VDD.n584 GND 0.03fF
C1105 VDD.n585 GND 0.02fF
C1106 VDD.n586 GND 0.02fF
C1107 VDD.n587 GND 0.02fF
C1108 VDD.n588 GND 0.03fF
C1109 VDD.n589 GND 0.02fF
C1110 VDD.n591 GND 0.02fF
C1111 VDD.n592 GND 0.02fF
C1112 VDD.n593 GND 0.02fF
C1113 VDD.n595 GND 0.27fF
C1114 VDD.n597 GND 0.02fF
C1115 VDD.n598 GND 0.02fF
C1116 VDD.n599 GND 0.03fF
C1117 VDD.n600 GND 0.02fF
C1118 VDD.n601 GND 0.27fF
C1119 VDD.n602 GND 0.01fF
C1120 VDD.n603 GND 0.02fF
C1121 VDD.n604 GND 0.03fF
C1122 VDD.n605 GND 0.27fF
C1123 VDD.n606 GND 0.01fF
C1124 VDD.n607 GND 0.02fF
C1125 VDD.n608 GND 0.02fF
C1126 VDD.n609 GND 0.22fF
C1127 VDD.n610 GND 0.01fF
C1128 VDD.n611 GND 0.07fF
C1129 VDD.n612 GND 0.02fF
C1130 VDD.n613 GND 0.14fF
C1131 VDD.n614 GND 0.17fF
C1132 VDD.n615 GND 0.01fF
C1133 VDD.n616 GND 0.02fF
C1134 VDD.n617 GND 0.02fF
C1135 VDD.n618 GND 0.14fF
C1136 VDD.n619 GND 0.16fF
C1137 VDD.n620 GND 0.01fF
C1138 VDD.n621 GND 0.11fF
C1139 VDD.n622 GND 0.02fF
C1140 VDD.n623 GND 0.02fF
C1141 VDD.n624 GND 0.02fF
C1142 VDD.n625 GND 0.18fF
C1143 VDD.n626 GND 0.15fF
C1144 VDD.n627 GND 0.01fF
C1145 VDD.n628 GND 0.02fF
C1146 VDD.n629 GND 0.03fF
C1147 VDD.n630 GND 0.18fF
C1148 VDD.n631 GND 0.15fF
C1149 VDD.n632 GND 0.01fF
C1150 VDD.n633 GND 0.02fF
C1151 VDD.n634 GND 0.03fF
C1152 VDD.n635 GND 0.11fF
C1153 VDD.n636 GND 0.02fF
C1154 VDD.n637 GND 0.14fF
C1155 VDD.n638 GND 0.16fF
C1156 VDD.n639 GND 0.01fF
C1157 VDD.n640 GND 0.02fF
C1158 VDD.n641 GND 0.02fF
C1159 VDD.n642 GND 0.14fF
C1160 VDD.n643 GND 0.17fF
C1161 VDD.n644 GND 0.01fF
C1162 VDD.n645 GND 0.02fF
C1163 VDD.n646 GND 0.02fF
C1164 VDD.n647 GND 0.06fF
C1165 VDD.n648 GND 0.23fF
C1166 VDD.n649 GND 0.01fF
C1167 VDD.n650 GND 0.01fF
C1168 VDD.n651 GND 0.02fF
C1169 VDD.n652 GND 0.27fF
C1170 VDD.n653 GND 0.01fF
C1171 VDD.n654 GND 0.02fF
C1172 VDD.n655 GND 0.02fF
C1173 VDD.n656 GND 0.27fF
C1174 VDD.n657 GND 0.01fF
C1175 VDD.n658 GND 0.02fF
C1176 VDD.n659 GND 0.03fF
C1177 VDD.n660 GND 0.02fF
C1178 VDD.n661 GND 0.02fF
C1179 VDD.n662 GND 0.02fF
C1180 VDD.n663 GND 0.26fF
C1181 VDD.n664 GND 0.04fF
C1182 VDD.n665 GND 0.03fF
C1183 VDD.n666 GND 0.02fF
C1184 VDD.n667 GND 0.02fF
C1185 VDD.n668 GND 0.02fF
C1186 VDD.n669 GND 0.03fF
C1187 VDD.n670 GND 0.02fF
C1188 VDD.n672 GND 0.02fF
C1189 VDD.n673 GND 0.02fF
C1190 VDD.n674 GND 0.02fF
C1191 VDD.n676 GND 0.27fF
C1192 VDD.n678 GND 0.02fF
C1193 VDD.n679 GND 0.02fF
C1194 VDD.n680 GND 0.03fF
C1195 VDD.n681 GND 0.02fF
C1196 VDD.n682 GND 0.27fF
C1197 VDD.n683 GND 0.01fF
C1198 VDD.n684 GND 0.02fF
C1199 VDD.n685 GND 0.03fF
C1200 VDD.n686 GND 0.06fF
C1201 VDD.n687 GND 0.24fF
C1202 VDD.n688 GND 0.01fF
C1203 VDD.n689 GND 0.01fF
C1204 VDD.n690 GND 0.02fF
C1205 VDD.n691 GND 0.14fF
C1206 VDD.n692 GND 0.17fF
C1207 VDD.n693 GND 0.01fF
C1208 VDD.n694 GND 0.02fF
C1209 VDD.n695 GND 0.02fF
C1210 VDD.n696 GND 0.11fF
C1211 VDD.n697 GND 0.03fF
C1212 VDD.n698 GND 0.31fF
C1213 VDD.n699 GND 0.01fF
C1214 VDD.n700 GND 0.02fF
C1215 VDD.n701 GND 0.03fF
C1216 VDD.n702 GND 0.17fF
C1217 VDD.n703 GND 0.14fF
C1218 VDD.n704 GND 0.01fF
C1219 VDD.n705 GND 0.02fF
C1220 VDD.n706 GND 0.03fF
C1221 VDD.n707 GND 0.14fF
C1222 VDD.n708 GND 0.16fF
C1223 VDD.n709 GND 0.01fF
C1224 VDD.n710 GND 0.02fF
C1225 VDD.n711 GND 0.02fF
C1226 VDD.n712 GND 0.06fF
C1227 VDD.n713 GND 0.25fF
C1228 VDD.n714 GND 0.01fF
C1229 VDD.n715 GND 0.01fF
C1230 VDD.n716 GND 0.02fF
C1231 VDD.n717 GND 0.27fF
C1232 VDD.n718 GND 0.01fF
C1233 VDD.n719 GND 0.02fF
C1234 VDD.n720 GND 0.03fF
C1235 VDD.n721 GND 0.02fF
C1236 VDD.n722 GND 0.02fF
C1237 VDD.n723 GND 0.02fF
C1238 VDD.n724 GND 0.26fF
C1239 VDD.n725 GND 0.04fF
C1240 VDD.n726 GND 0.03fF
C1241 VDD.n727 GND 0.02fF
C1242 VDD.n728 GND 0.02fF
C1243 VDD.n729 GND 0.02fF
C1244 VDD.n730 GND 0.03fF
C1245 VDD.n731 GND 0.02fF
C1246 VDD.n733 GND 0.02fF
C1247 VDD.n734 GND 0.02fF
C1248 VDD.n735 GND 0.02fF
C1249 VDD.n737 GND 0.27fF
C1250 VDD.n739 GND 0.02fF
C1251 VDD.n740 GND 0.02fF
C1252 VDD.n741 GND 0.03fF
C1253 VDD.n742 GND 0.02fF
C1254 VDD.n743 GND 0.27fF
C1255 VDD.n744 GND 0.01fF
C1256 VDD.n745 GND 0.02fF
C1257 VDD.n746 GND 0.03fF
C1258 VDD.n747 GND 0.27fF
C1259 VDD.n748 GND 0.01fF
C1260 VDD.n749 GND 0.02fF
C1261 VDD.n750 GND 0.02fF
C1262 VDD.n751 GND 0.22fF
C1263 VDD.n752 GND 0.01fF
C1264 VDD.n753 GND 0.07fF
C1265 VDD.n754 GND 0.02fF
C1266 VDD.n755 GND 0.14fF
C1267 VDD.n756 GND 0.17fF
C1268 VDD.n757 GND 0.01fF
C1269 VDD.n758 GND 0.02fF
C1270 VDD.n759 GND 0.02fF
C1271 VDD.n760 GND 0.14fF
C1272 VDD.n761 GND 0.16fF
C1273 VDD.n762 GND 0.01fF
C1274 VDD.n763 GND 0.11fF
C1275 VDD.n764 GND 0.02fF
C1276 VDD.n765 GND 0.02fF
C1277 VDD.n766 GND 0.02fF
C1278 VDD.n767 GND 0.18fF
C1279 VDD.n768 GND 0.15fF
C1280 VDD.n769 GND 0.01fF
C1281 VDD.n770 GND 0.02fF
C1282 VDD.n771 GND 0.03fF
C1283 VDD.n772 GND 0.18fF
C1284 VDD.n773 GND 0.15fF
C1285 VDD.n774 GND 0.01fF
C1286 VDD.n775 GND 0.02fF
C1287 VDD.n776 GND 0.03fF
C1288 VDD.n777 GND 0.11fF
C1289 VDD.n778 GND 0.02fF
C1290 VDD.n779 GND 0.14fF
C1291 VDD.n780 GND 0.16fF
C1292 VDD.n781 GND 0.01fF
C1293 VDD.n782 GND 0.02fF
C1294 VDD.n783 GND 0.02fF
C1295 VDD.n784 GND 0.14fF
C1296 VDD.n785 GND 0.17fF
C1297 VDD.n786 GND 0.01fF
C1298 VDD.n787 GND 0.02fF
C1299 VDD.n788 GND 0.02fF
C1300 VDD.n789 GND 0.02fF
C1301 VDD.n790 GND 0.02fF
C1302 VDD.n791 GND 0.02fF
C1303 VDD.n792 GND 0.20fF
C1304 VDD.n793 GND 0.03fF
C1305 VDD.n794 GND 0.02fF
C1306 VDD.n795 GND 0.02fF
C1307 VDD.n796 GND 0.02fF
C1308 VDD.n797 GND 0.03fF
C1309 VDD.n798 GND 0.02fF
C1310 VDD.n800 GND 0.02fF
C1311 VDD.n801 GND 0.02fF
C1312 VDD.n802 GND 0.02fF
C1313 VDD.n804 GND 0.46fF
C1314 VDD.n806 GND 0.03fF
C1315 VDD.n807 GND 0.04fF
C1316 VDD.n808 GND 0.27fF
C1317 VDD.n809 GND 0.02fF
C1318 VDD.n810 GND 0.03fF
C1319 VDD.n811 GND 0.03fF
C1320 VDD.n812 GND 0.27fF
C1321 VDD.n813 GND 0.01fF
C1322 VDD.n814 GND 0.02fF
C1323 VDD.n815 GND 0.02fF
C1324 VDD.n816 GND 0.06fF
C1325 VDD.n817 GND 0.23fF
C1326 VDD.n818 GND 0.01fF
C1327 VDD.n819 GND 0.01fF
C1328 VDD.n820 GND 0.02fF
C1329 VDD.n821 GND 0.14fF
C1330 VDD.n822 GND 0.17fF
C1331 VDD.n823 GND 0.01fF
C1332 VDD.n824 GND 0.02fF
C1333 VDD.n825 GND 0.02fF
C1334 VDD.n826 GND 0.11fF
C1335 VDD.n827 GND 0.02fF
C1336 VDD.n828 GND 0.14fF
C1337 VDD.n829 GND 0.16fF
C1338 VDD.n830 GND 0.01fF
C1339 VDD.n831 GND 0.02fF
C1340 VDD.n832 GND 0.02fF
C1341 VDD.n833 GND 0.18fF
C1342 VDD.n834 GND 0.15fF
C1343 VDD.n835 GND 0.01fF
C1344 VDD.n836 GND 0.02fF
C1345 VDD.n837 GND 0.03fF
C1346 VDD.n838 GND 0.18fF
C1347 VDD.n839 GND 0.15fF
C1348 VDD.n840 GND 0.01fF
C1349 VDD.n841 GND 0.02fF
C1350 VDD.n842 GND 0.03fF
C1351 VDD.n843 GND 0.14fF
C1352 VDD.n844 GND 0.16fF
C1353 VDD.n845 GND 0.01fF
C1354 VDD.n846 GND 0.11fF
C1355 VDD.n847 GND 0.02fF
C1356 VDD.n848 GND 0.02fF
C1357 VDD.n849 GND 0.02fF
C1358 VDD.n850 GND 0.14fF
C1359 VDD.n851 GND 0.17fF
C1360 VDD.n852 GND 0.01fF
C1361 VDD.n853 GND 0.02fF
C1362 VDD.n854 GND 0.02fF
C1363 VDD.n855 GND 0.22fF
C1364 VDD.n856 GND 0.01fF
C1365 VDD.n857 GND 0.07fF
C1366 VDD.n858 GND 0.02fF
C1367 VDD.n859 GND 0.27fF
C1368 VDD.n860 GND 0.01fF
C1369 VDD.n861 GND 0.02fF
C1370 VDD.n862 GND 0.02fF
C1371 VDD.n863 GND 0.27fF
C1372 VDD.n864 GND 0.01fF
C1373 VDD.n865 GND 0.02fF
C1374 VDD.n866 GND 0.03fF
C1375 VDD.n867 GND 0.02fF
C1376 VDD.n868 GND 0.02fF
C1377 VDD.n869 GND 0.02fF
C1378 VDD.n870 GND 0.02fF
C1379 VDD.n871 GND 0.02fF
C1380 VDD.n872 GND 0.02fF
C1381 VDD.n874 GND 0.02fF
C1382 VDD.n875 GND 0.02fF
C1383 VDD.n876 GND 0.02fF
C1384 VDD.n877 GND 0.02fF
C1385 VDD.n879 GND 0.04fF
C1386 VDD.n880 GND 0.02fF
C1387 VDD.n881 GND 0.31fF
C1388 VDD.n882 GND 0.04fF
C1389 VDD.n884 GND 0.27fF
C1390 VDD.n886 GND 0.02fF
C1391 VDD.n887 GND 0.02fF
C1392 VDD.n888 GND 0.03fF
C1393 VDD.n889 GND 0.02fF
C1394 VDD.n890 GND 0.27fF
C1395 VDD.n891 GND 0.01fF
C1396 VDD.n892 GND 0.02fF
C1397 VDD.n893 GND 0.03fF
C1398 VDD.n894 GND 0.27fF
C1399 VDD.n895 GND 0.01fF
C1400 VDD.n896 GND 0.02fF
C1401 VDD.n897 GND 0.02fF
C1402 VDD.n898 GND 0.06fF
C1403 VDD.n899 GND 0.23fF
C1404 VDD.n900 GND 0.01fF
C1405 VDD.n901 GND 0.01fF
C1406 VDD.n902 GND 0.02fF
C1407 VDD.n903 GND 0.14fF
C1408 VDD.n904 GND 0.17fF
C1409 VDD.n905 GND 0.01fF
C1410 VDD.n906 GND 0.02fF
C1411 VDD.n907 GND 0.02fF
C1412 VDD.n908 GND 0.11fF
C1413 VDD.n909 GND 0.02fF
C1414 VDD.n910 GND 0.14fF
C1415 VDD.n911 GND 0.16fF
C1416 VDD.n912 GND 0.01fF
C1417 VDD.n913 GND 0.02fF
C1418 VDD.n914 GND 0.02fF
C1419 VDD.n915 GND 0.18fF
C1420 VDD.n916 GND 0.15fF
C1421 VDD.n917 GND 0.01fF
C1422 VDD.n918 GND 0.02fF
C1423 VDD.n919 GND 0.03fF
C1424 VDD.n920 GND 0.18fF
C1425 VDD.n921 GND 0.15fF
C1426 VDD.n922 GND 0.01fF
C1427 VDD.n923 GND 0.02fF
C1428 VDD.n924 GND 0.03fF
C1429 VDD.n925 GND 0.14fF
C1430 VDD.n926 GND 0.16fF
C1431 VDD.n927 GND 0.01fF
C1432 VDD.n928 GND 0.11fF
C1433 VDD.n929 GND 0.02fF
C1434 VDD.n930 GND 0.02fF
C1435 VDD.n931 GND 0.02fF
C1436 VDD.n932 GND 0.14fF
C1437 VDD.n933 GND 0.17fF
C1438 VDD.n934 GND 0.01fF
C1439 VDD.n935 GND 0.02fF
C1440 VDD.n936 GND 0.02fF
C1441 VDD.n937 GND 0.22fF
C1442 VDD.n938 GND 0.01fF
C1443 VDD.n939 GND 0.07fF
C1444 VDD.n940 GND 0.02fF
C1445 VDD.n941 GND 0.27fF
C1446 VDD.n942 GND 0.01fF
C1447 VDD.n943 GND 0.02fF
C1448 VDD.n944 GND 0.02fF
C1449 VDD.n945 GND 0.27fF
C1450 VDD.n946 GND 0.01fF
C1451 VDD.n947 GND 0.02fF
C1452 VDD.n948 GND 0.03fF
C1453 VDD.n949 GND 0.02fF
C1454 VDD.n950 GND 0.02fF
C1455 VDD.n951 GND 0.02fF
C1456 VDD.n952 GND 0.26fF
C1457 VDD.n953 GND 0.04fF
C1458 VDD.n954 GND 0.03fF
C1459 VDD.n955 GND 0.02fF
C1460 VDD.n956 GND 0.02fF
C1461 VDD.n957 GND 0.02fF
C1462 VDD.n958 GND 0.03fF
C1463 VDD.n959 GND 0.02fF
C1464 VDD.n961 GND 0.02fF
C1465 VDD.n962 GND 0.02fF
C1466 VDD.n963 GND 0.02fF
C1467 VDD.n965 GND 0.27fF
C1468 VDD.n967 GND 0.02fF
C1469 VDD.n968 GND 0.02fF
C1470 VDD.n969 GND 0.03fF
C1471 VDD.n970 GND 0.02fF
C1472 VDD.n971 GND 0.27fF
C1473 VDD.n972 GND 0.01fF
C1474 VDD.n973 GND 0.02fF
C1475 VDD.n974 GND 0.03fF
C1476 VDD.n975 GND 0.06fF
C1477 VDD.n976 GND 0.25fF
C1478 VDD.n977 GND 0.01fF
C1479 VDD.n978 GND 0.01fF
C1480 VDD.n979 GND 0.02fF
C1481 VDD.n980 GND 0.14fF
C1482 VDD.n981 GND 0.16fF
C1483 VDD.n982 GND 0.01fF
C1484 VDD.n983 GND 0.02fF
C1485 VDD.n984 GND 0.02fF
C1486 VDD.n985 GND 0.17fF
C1487 VDD.n986 GND 0.14fF
C1488 VDD.n987 GND 0.01fF
C1489 VDD.n988 GND 0.02fF
C1490 VDD.n989 GND 0.03fF
C1491 VDD.n990 GND 0.11fF
C1492 VDD.n991 GND 0.03fF
C1493 VDD.n992 GND 0.31fF
C1494 VDD.n993 GND 0.01fF
C1495 VDD.n994 GND 0.02fF
C1496 VDD.n995 GND 0.03fF
C1497 VDD.n996 GND 0.14fF
C1498 VDD.n997 GND 0.17fF
C1499 VDD.n998 GND 0.01fF
C1500 VDD.n999 GND 0.02fF
C1501 VDD.n1000 GND 0.02fF
C1502 VDD.n1001 GND 0.06fF
C1503 VDD.n1002 GND 0.24fF
C1504 VDD.n1003 GND 0.01fF
C1505 VDD.n1004 GND 0.01fF
C1506 VDD.n1005 GND 0.02fF
C1507 VDD.n1006 GND 0.27fF
C1508 VDD.n1007 GND 0.01fF
C1509 VDD.n1008 GND 0.02fF
C1510 VDD.n1009 GND 0.03fF
C1511 VDD.n1010 GND 0.02fF
C1512 VDD.n1011 GND 0.02fF
C1513 VDD.n1012 GND 0.02fF
C1514 VDD.n1013 GND 0.26fF
C1515 VDD.n1014 GND 0.04fF
C1516 VDD.n1015 GND 0.03fF
C1517 VDD.n1016 GND 0.02fF
C1518 VDD.n1017 GND 0.02fF
C1519 VDD.n1018 GND 0.02fF
C1520 VDD.n1019 GND 0.03fF
C1521 VDD.n1020 GND 0.02fF
C1522 VDD.n1022 GND 0.02fF
C1523 VDD.n1023 GND 0.02fF
C1524 VDD.n1024 GND 0.02fF
C1525 VDD.n1026 GND 0.27fF
C1526 VDD.n1028 GND 0.02fF
C1527 VDD.n1029 GND 0.02fF
C1528 VDD.n1030 GND 0.03fF
C1529 VDD.n1031 GND 0.02fF
C1530 VDD.n1032 GND 0.27fF
C1531 VDD.n1033 GND 0.01fF
C1532 VDD.n1034 GND 0.02fF
C1533 VDD.n1035 GND 0.03fF
C1534 VDD.n1036 GND 0.27fF
C1535 VDD.n1037 GND 0.01fF
C1536 VDD.n1038 GND 0.02fF
C1537 VDD.n1039 GND 0.02fF
C1538 VDD.n1040 GND 0.06fF
C1539 VDD.n1041 GND 0.23fF
C1540 VDD.n1042 GND 0.01fF
C1541 VDD.n1043 GND 0.01fF
C1542 VDD.n1044 GND 0.02fF
C1543 VDD.n1045 GND 0.14fF
C1544 VDD.n1046 GND 0.17fF
C1545 VDD.n1047 GND 0.01fF
C1546 VDD.n1048 GND 0.02fF
C1547 VDD.n1049 GND 0.02fF
C1548 VDD.n1050 GND 0.11fF
C1549 VDD.n1051 GND 0.02fF
C1550 VDD.n1052 GND 0.14fF
C1551 VDD.n1053 GND 0.16fF
C1552 VDD.n1054 GND 0.01fF
C1553 VDD.n1055 GND 0.02fF
C1554 VDD.n1056 GND 0.02fF
C1555 VDD.n1057 GND 0.18fF
C1556 VDD.n1058 GND 0.15fF
C1557 VDD.n1059 GND 0.01fF
C1558 VDD.n1060 GND 0.02fF
C1559 VDD.n1061 GND 0.03fF
C1560 VDD.n1062 GND 0.18fF
C1561 VDD.n1063 GND 0.15fF
C1562 VDD.n1064 GND 0.01fF
C1563 VDD.n1065 GND 0.02fF
C1564 VDD.n1066 GND 0.03fF
C1565 VDD.n1067 GND 0.14fF
C1566 VDD.n1068 GND 0.16fF
C1567 VDD.n1069 GND 0.01fF
C1568 VDD.n1070 GND 0.11fF
C1569 VDD.n1071 GND 0.02fF
C1570 VDD.n1072 GND 0.02fF
C1571 VDD.n1073 GND 0.02fF
C1572 VDD.n1074 GND 0.14fF
C1573 VDD.n1075 GND 0.17fF
C1574 VDD.n1076 GND 0.01fF
C1575 VDD.n1077 GND 0.02fF
C1576 VDD.n1078 GND 0.02fF
C1577 VDD.n1079 GND 0.22fF
C1578 VDD.n1080 GND 0.01fF
C1579 VDD.n1081 GND 0.07fF
C1580 VDD.n1082 GND 0.02fF
C1581 VDD.n1083 GND 0.27fF
C1582 VDD.n1084 GND 0.01fF
C1583 VDD.n1085 GND 0.02fF
C1584 VDD.n1086 GND 0.02fF
C1585 VDD.n1087 GND 0.27fF
C1586 VDD.n1088 GND 0.01fF
C1587 VDD.n1089 GND 0.02fF
C1588 VDD.n1090 GND 0.03fF
C1589 VDD.n1091 GND 0.02fF
C1590 VDD.n1092 GND 0.02fF
C1591 VDD.n1093 GND 0.02fF
C1592 VDD.n1094 GND 0.31fF
C1593 VDD.n1095 GND 0.04fF
C1594 VDD.n1096 GND 0.03fF
C1595 VDD.n1097 GND 0.02fF
C1596 VDD.n1098 GND 0.02fF
C1597 VDD.n1099 GND 0.02fF
C1598 VDD.n1100 GND 0.03fF
C1599 VDD.n1101 GND 0.02fF
C1600 VDD.n1103 GND 0.02fF
C1601 VDD.n1104 GND 0.02fF
C1602 VDD.n1105 GND 0.02fF
C1603 VDD.n1107 GND 0.27fF
C1604 VDD.n1109 GND 0.02fF
C1605 VDD.n1110 GND 0.02fF
C1606 VDD.n1111 GND 0.03fF
C1607 VDD.n1112 GND 0.02fF
C1608 VDD.n1113 GND 0.27fF
C1609 VDD.n1114 GND 0.01fF
C1610 VDD.n1115 GND 0.02fF
C1611 VDD.n1116 GND 0.03fF
C1612 VDD.n1117 GND 0.27fF
C1613 VDD.n1118 GND 0.01fF
C1614 VDD.n1119 GND 0.02fF
C1615 VDD.n1120 GND 0.02fF
C1616 VDD.n1121 GND 0.06fF
C1617 VDD.n1122 GND 0.23fF
C1618 VDD.n1123 GND 0.01fF
C1619 VDD.n1124 GND 0.01fF
C1620 VDD.n1125 GND 0.02fF
C1621 VDD.n1126 GND 0.14fF
C1622 VDD.n1127 GND 0.17fF
C1623 VDD.n1128 GND 0.01fF
C1624 VDD.n1129 GND 0.02fF
C1625 VDD.n1130 GND 0.02fF
C1626 VDD.n1131 GND 0.11fF
C1627 VDD.n1132 GND 0.02fF
C1628 VDD.n1133 GND 0.14fF
C1629 VDD.n1134 GND 0.16fF
C1630 VDD.n1135 GND 0.01fF
C1631 VDD.n1136 GND 0.02fF
C1632 VDD.n1137 GND 0.02fF
C1633 VDD.n1138 GND 0.18fF
C1634 VDD.n1139 GND 0.15fF
C1635 VDD.n1140 GND 0.01fF
C1636 VDD.n1141 GND 0.02fF
C1637 VDD.n1142 GND 0.03fF
C1638 VDD.n1143 GND 0.18fF
C1639 VDD.n1144 GND 0.15fF
C1640 VDD.n1145 GND 0.01fF
C1641 VDD.n1146 GND 0.02fF
C1642 VDD.n1147 GND 0.03fF
C1643 VDD.n1148 GND 0.14fF
C1644 VDD.n1149 GND 0.16fF
C1645 VDD.n1150 GND 0.01fF
C1646 VDD.n1151 GND 0.11fF
C1647 VDD.n1152 GND 0.02fF
C1648 VDD.n1153 GND 0.02fF
C1649 VDD.n1154 GND 0.02fF
C1650 VDD.n1155 GND 0.14fF
C1651 VDD.n1156 GND 0.17fF
C1652 VDD.n1157 GND 0.01fF
C1653 VDD.n1158 GND 0.02fF
C1654 VDD.n1159 GND 0.02fF
C1655 VDD.n1160 GND 0.22fF
C1656 VDD.n1161 GND 0.01fF
C1657 VDD.n1162 GND 0.07fF
C1658 VDD.n1163 GND 0.02fF
C1659 VDD.n1164 GND 0.27fF
C1660 VDD.n1165 GND 0.01fF
C1661 VDD.n1166 GND 0.02fF
C1662 VDD.n1167 GND 0.02fF
C1663 VDD.n1168 GND 0.27fF
C1664 VDD.n1169 GND 0.01fF
C1665 VDD.n1170 GND 0.02fF
C1666 VDD.n1171 GND 0.03fF
C1667 VDD.n1172 GND 0.02fF
C1668 VDD.n1173 GND 0.02fF
C1669 VDD.n1174 GND 0.02fF
C1670 VDD.n1175 GND 0.26fF
C1671 VDD.n1176 GND 0.04fF
C1672 VDD.n1177 GND 0.03fF
C1673 VDD.n1178 GND 0.02fF
C1674 VDD.n1179 GND 0.02fF
C1675 VDD.n1180 GND 0.02fF
C1676 VDD.n1181 GND 0.03fF
C1677 VDD.n1182 GND 0.02fF
C1678 VDD.n1184 GND 0.02fF
C1679 VDD.n1185 GND 0.02fF
C1680 VDD.n1186 GND 0.02fF
C1681 VDD.n1188 GND 0.27fF
C1682 VDD.n1190 GND 0.02fF
C1683 VDD.n1191 GND 0.02fF
C1684 VDD.n1192 GND 0.03fF
C1685 VDD.n1193 GND 0.02fF
C1686 VDD.n1194 GND 0.27fF
C1687 VDD.n1195 GND 0.01fF
C1688 VDD.n1196 GND 0.02fF
C1689 VDD.n1197 GND 0.03fF
C1690 VDD.n1198 GND 0.06fF
C1691 VDD.n1199 GND 0.25fF
C1692 VDD.n1200 GND 0.01fF
C1693 VDD.n1201 GND 0.01fF
C1694 VDD.n1202 GND 0.02fF
C1695 VDD.n1203 GND 0.14fF
C1696 VDD.n1204 GND 0.16fF
C1697 VDD.n1205 GND 0.01fF
C1698 VDD.n1206 GND 0.02fF
C1699 VDD.n1207 GND 0.02fF
C1700 VDD.n1208 GND 0.17fF
C1701 VDD.n1209 GND 0.14fF
C1702 VDD.n1210 GND 0.01fF
C1703 VDD.n1211 GND 0.02fF
C1704 VDD.n1212 GND 0.03fF
C1705 VDD.n1213 GND 0.11fF
C1706 VDD.n1214 GND 0.03fF
C1707 VDD.n1215 GND 0.31fF
C1708 VDD.n1216 GND 0.01fF
C1709 VDD.n1217 GND 0.02fF
C1710 VDD.n1218 GND 0.03fF
C1711 VDD.n1219 GND 0.14fF
C1712 VDD.n1220 GND 0.17fF
C1713 VDD.n1221 GND 0.01fF
C1714 VDD.n1222 GND 0.02fF
C1715 VDD.n1223 GND 0.02fF
C1716 VDD.n1224 GND 0.06fF
C1717 VDD.n1225 GND 0.24fF
C1718 VDD.n1226 GND 0.01fF
C1719 VDD.n1227 GND 0.01fF
C1720 VDD.n1228 GND 0.02fF
C1721 VDD.n1229 GND 0.27fF
C1722 VDD.n1230 GND 0.01fF
C1723 VDD.n1231 GND 0.02fF
C1724 VDD.n1232 GND 0.03fF
C1725 VDD.n1233 GND 0.02fF
C1726 VDD.n1234 GND 0.02fF
C1727 VDD.n1235 GND 0.02fF
C1728 VDD.n1236 GND 0.26fF
C1729 VDD.n1237 GND 0.04fF
C1730 VDD.n1238 GND 0.03fF
C1731 VDD.n1239 GND 0.02fF
C1732 VDD.n1240 GND 0.02fF
C1733 VDD.n1241 GND 0.02fF
C1734 VDD.n1242 GND 0.03fF
C1735 VDD.n1243 GND 0.02fF
C1736 VDD.n1245 GND 0.02fF
C1737 VDD.n1246 GND 0.02fF
C1738 VDD.n1247 GND 0.02fF
C1739 VDD.n1249 GND 0.27fF
C1740 VDD.n1251 GND 0.02fF
C1741 VDD.n1252 GND 0.02fF
C1742 VDD.n1253 GND 0.03fF
C1743 VDD.n1254 GND 0.02fF
C1744 VDD.n1255 GND 0.27fF
C1745 VDD.n1256 GND 0.01fF
C1746 VDD.n1257 GND 0.02fF
C1747 VDD.n1258 GND 0.03fF
C1748 VDD.n1259 GND 0.27fF
C1749 VDD.n1260 GND 0.01fF
C1750 VDD.n1261 GND 0.02fF
C1751 VDD.n1262 GND 0.02fF
C1752 VDD.n1263 GND 0.06fF
C1753 VDD.n1264 GND 0.23fF
C1754 VDD.n1265 GND 0.01fF
C1755 VDD.n1266 GND 0.01fF
C1756 VDD.n1267 GND 0.02fF
C1757 VDD.n1268 GND 0.14fF
C1758 VDD.n1269 GND 0.17fF
C1759 VDD.n1270 GND 0.01fF
C1760 VDD.n1271 GND 0.02fF
C1761 VDD.n1272 GND 0.02fF
C1762 VDD.n1273 GND 0.11fF
C1763 VDD.n1274 GND 0.02fF
C1764 VDD.n1275 GND 0.14fF
C1765 VDD.n1276 GND 0.16fF
C1766 VDD.n1277 GND 0.01fF
C1767 VDD.n1278 GND 0.02fF
C1768 VDD.n1279 GND 0.02fF
C1769 VDD.n1280 GND 0.18fF
C1770 VDD.n1281 GND 0.15fF
C1771 VDD.n1282 GND 0.01fF
C1772 VDD.n1283 GND 0.02fF
C1773 VDD.n1284 GND 0.03fF
C1774 VDD.n1285 GND 0.18fF
C1775 VDD.n1286 GND 0.15fF
C1776 VDD.n1287 GND 0.01fF
C1777 VDD.n1288 GND 0.02fF
C1778 VDD.n1289 GND 0.03fF
C1779 VDD.n1290 GND 0.14fF
C1780 VDD.n1291 GND 0.16fF
C1781 VDD.n1292 GND 0.01fF
C1782 VDD.n1293 GND 0.11fF
C1783 VDD.n1294 GND 0.02fF
C1784 VDD.n1295 GND 0.02fF
C1785 VDD.n1296 GND 0.02fF
C1786 VDD.n1297 GND 0.14fF
C1787 VDD.n1298 GND 0.17fF
C1788 VDD.n1299 GND 0.01fF
C1789 VDD.n1300 GND 0.02fF
C1790 VDD.n1301 GND 0.02fF
C1791 VDD.n1302 GND 0.22fF
C1792 VDD.n1303 GND 0.01fF
C1793 VDD.n1304 GND 0.07fF
C1794 VDD.n1305 GND 0.02fF
C1795 VDD.n1306 GND 0.27fF
C1796 VDD.n1307 GND 0.01fF
C1797 VDD.n1308 GND 0.02fF
C1798 VDD.n1309 GND 0.02fF
C1799 VDD.n1310 GND 0.27fF
C1800 VDD.n1311 GND 0.01fF
C1801 VDD.n1312 GND 0.02fF
C1802 VDD.n1313 GND 0.03fF
C1803 VDD.n1314 GND 0.02fF
C1804 VDD.n1315 GND 0.02fF
C1805 VDD.n1316 GND 0.02fF
C1806 VDD.n1317 GND 0.31fF
C1807 VDD.n1318 GND 0.04fF
C1808 VDD.n1319 GND 0.03fF
C1809 VDD.n1320 GND 0.02fF
C1810 VDD.n1321 GND 0.02fF
C1811 VDD.n1322 GND 0.02fF
C1812 VDD.n1323 GND 0.03fF
C1813 VDD.n1324 GND 0.02fF
C1814 VDD.n1326 GND 0.02fF
C1815 VDD.n1327 GND 0.02fF
C1816 VDD.n1328 GND 0.02fF
C1817 VDD.n1330 GND 0.27fF
C1818 VDD.n1332 GND 0.02fF
C1819 VDD.n1333 GND 0.02fF
C1820 VDD.n1334 GND 0.03fF
C1821 VDD.n1335 GND 0.02fF
C1822 VDD.n1336 GND 0.27fF
C1823 VDD.n1337 GND 0.01fF
C1824 VDD.n1338 GND 0.02fF
C1825 VDD.n1339 GND 0.03fF
C1826 VDD.n1340 GND 0.27fF
C1827 VDD.n1341 GND 0.01fF
C1828 VDD.n1342 GND 0.02fF
C1829 VDD.n1343 GND 0.02fF
C1830 VDD.n1344 GND 0.06fF
C1831 VDD.n1345 GND 0.23fF
C1832 VDD.n1346 GND 0.01fF
C1833 VDD.n1347 GND 0.01fF
C1834 VDD.n1348 GND 0.02fF
C1835 VDD.n1349 GND 0.14fF
C1836 VDD.n1350 GND 0.17fF
C1837 VDD.n1351 GND 0.01fF
C1838 VDD.n1352 GND 0.02fF
C1839 VDD.n1353 GND 0.02fF
C1840 VDD.n1354 GND 0.11fF
C1841 VDD.n1355 GND 0.02fF
C1842 VDD.n1356 GND 0.14fF
C1843 VDD.n1357 GND 0.16fF
C1844 VDD.n1358 GND 0.01fF
C1845 VDD.n1359 GND 0.02fF
C1846 VDD.n1360 GND 0.02fF
C1847 VDD.n1361 GND 0.18fF
C1848 VDD.n1362 GND 0.15fF
C1849 VDD.n1363 GND 0.01fF
C1850 VDD.n1364 GND 0.02fF
C1851 VDD.n1365 GND 0.03fF
C1852 VDD.n1366 GND 0.18fF
C1853 VDD.n1367 GND 0.15fF
C1854 VDD.n1368 GND 0.01fF
C1855 VDD.n1369 GND 0.02fF
C1856 VDD.n1370 GND 0.03fF
C1857 VDD.n1371 GND 0.14fF
C1858 VDD.n1372 GND 0.16fF
C1859 VDD.n1373 GND 0.01fF
C1860 VDD.n1374 GND 0.11fF
C1861 VDD.n1375 GND 0.02fF
C1862 VDD.n1376 GND 0.02fF
C1863 VDD.n1377 GND 0.02fF
C1864 VDD.n1378 GND 0.14fF
C1865 VDD.n1379 GND 0.17fF
C1866 VDD.n1380 GND 0.01fF
C1867 VDD.n1381 GND 0.02fF
C1868 VDD.n1382 GND 0.02fF
C1869 VDD.n1383 GND 0.22fF
C1870 VDD.n1384 GND 0.01fF
C1871 VDD.n1385 GND 0.07fF
C1872 VDD.n1386 GND 0.02fF
C1873 VDD.n1387 GND 0.27fF
C1874 VDD.n1388 GND 0.01fF
C1875 VDD.n1389 GND 0.02fF
C1876 VDD.n1390 GND 0.02fF
C1877 VDD.n1391 GND 0.27fF
C1878 VDD.n1392 GND 0.01fF
C1879 VDD.n1393 GND 0.02fF
C1880 VDD.n1394 GND 0.03fF
C1881 VDD.n1395 GND 0.02fF
C1882 VDD.n1396 GND 0.02fF
C1883 VDD.n1397 GND 0.02fF
C1884 VDD.n1398 GND 0.26fF
C1885 VDD.n1399 GND 0.04fF
C1886 VDD.n1400 GND 0.03fF
C1887 VDD.n1401 GND 0.02fF
C1888 VDD.n1402 GND 0.02fF
C1889 VDD.n1403 GND 0.02fF
C1890 VDD.n1404 GND 0.03fF
C1891 VDD.n1405 GND 0.02fF
C1892 VDD.n1407 GND 0.02fF
C1893 VDD.n1408 GND 0.02fF
C1894 VDD.n1409 GND 0.02fF
C1895 VDD.n1411 GND 0.27fF
C1896 VDD.n1413 GND 0.02fF
C1897 VDD.n1414 GND 0.02fF
C1898 VDD.n1415 GND 0.03fF
C1899 VDD.n1416 GND 0.02fF
C1900 VDD.n1417 GND 0.27fF
C1901 VDD.n1418 GND 0.01fF
C1902 VDD.n1419 GND 0.02fF
C1903 VDD.n1420 GND 0.03fF
C1904 VDD.n1421 GND 0.06fF
C1905 VDD.n1422 GND 0.25fF
C1906 VDD.n1423 GND 0.01fF
C1907 VDD.n1424 GND 0.01fF
C1908 VDD.n1425 GND 0.02fF
C1909 VDD.n1426 GND 0.14fF
C1910 VDD.n1427 GND 0.16fF
C1911 VDD.n1428 GND 0.01fF
C1912 VDD.n1429 GND 0.02fF
C1913 VDD.n1430 GND 0.02fF
C1914 VDD.n1431 GND 0.17fF
C1915 VDD.n1432 GND 0.14fF
C1916 VDD.n1433 GND 0.01fF
C1917 VDD.n1434 GND 0.02fF
C1918 VDD.n1435 GND 0.03fF
C1919 VDD.n1436 GND 0.11fF
C1920 VDD.n1437 GND 0.03fF
C1921 VDD.n1438 GND 0.31fF
C1922 VDD.n1439 GND 0.01fF
C1923 VDD.n1440 GND 0.02fF
C1924 VDD.n1441 GND 0.03fF
C1925 VDD.n1442 GND 0.14fF
C1926 VDD.n1443 GND 0.17fF
C1927 VDD.n1444 GND 0.01fF
C1928 VDD.n1445 GND 0.02fF
C1929 VDD.n1446 GND 0.02fF
C1930 VDD.n1447 GND 0.06fF
C1931 VDD.n1448 GND 0.24fF
C1932 VDD.n1449 GND 0.01fF
C1933 VDD.n1450 GND 0.01fF
C1934 VDD.n1451 GND 0.02fF
C1935 VDD.n1452 GND 0.27fF
C1936 VDD.n1453 GND 0.01fF
C1937 VDD.n1454 GND 0.02fF
C1938 VDD.n1455 GND 0.03fF
C1939 VDD.n1456 GND 0.02fF
C1940 VDD.n1457 GND 0.02fF
C1941 VDD.n1458 GND 0.02fF
C1942 VDD.n1459 GND 0.26fF
C1943 VDD.n1460 GND 0.04fF
C1944 VDD.n1461 GND 0.03fF
C1945 VDD.n1462 GND 0.02fF
C1946 VDD.n1463 GND 0.02fF
C1947 VDD.n1464 GND 0.02fF
C1948 VDD.n1465 GND 0.03fF
C1949 VDD.n1466 GND 0.02fF
C1950 VDD.n1468 GND 0.02fF
C1951 VDD.n1469 GND 0.02fF
C1952 VDD.n1470 GND 0.02fF
C1953 VDD.n1472 GND 0.27fF
C1954 VDD.n1474 GND 0.02fF
C1955 VDD.n1475 GND 0.02fF
C1956 VDD.n1476 GND 0.03fF
C1957 VDD.n1477 GND 0.02fF
C1958 VDD.n1478 GND 0.27fF
C1959 VDD.n1479 GND 0.01fF
C1960 VDD.n1480 GND 0.02fF
C1961 VDD.n1481 GND 0.03fF
C1962 VDD.n1482 GND 0.27fF
C1963 VDD.n1483 GND 0.01fF
C1964 VDD.n1484 GND 0.02fF
C1965 VDD.n1485 GND 0.02fF
C1966 VDD.n1486 GND 0.06fF
C1967 VDD.n1487 GND 0.23fF
C1968 VDD.n1488 GND 0.01fF
C1969 VDD.n1489 GND 0.01fF
C1970 VDD.n1490 GND 0.02fF
C1971 VDD.n1491 GND 0.14fF
C1972 VDD.n1492 GND 0.17fF
C1973 VDD.n1493 GND 0.01fF
C1974 VDD.n1494 GND 0.02fF
C1975 VDD.n1495 GND 0.02fF
C1976 VDD.n1496 GND 0.11fF
C1977 VDD.n1497 GND 0.02fF
C1978 VDD.n1498 GND 0.14fF
C1979 VDD.n1499 GND 0.16fF
C1980 VDD.n1500 GND 0.01fF
C1981 VDD.n1501 GND 0.02fF
C1982 VDD.n1502 GND 0.02fF
C1983 VDD.n1503 GND 0.18fF
C1984 VDD.n1504 GND 0.15fF
C1985 VDD.n1505 GND 0.01fF
C1986 VDD.n1506 GND 0.02fF
C1987 VDD.n1507 GND 0.03fF
C1988 VDD.n1508 GND 0.18fF
C1989 VDD.n1509 GND 0.15fF
C1990 VDD.n1510 GND 0.01fF
C1991 VDD.n1511 GND 0.02fF
C1992 VDD.n1512 GND 0.03fF
C1993 VDD.n1513 GND 0.14fF
C1994 VDD.n1514 GND 0.16fF
C1995 VDD.n1515 GND 0.01fF
C1996 VDD.n1516 GND 0.11fF
C1997 VDD.n1517 GND 0.02fF
C1998 VDD.n1518 GND 0.02fF
C1999 VDD.n1519 GND 0.02fF
C2000 VDD.n1520 GND 0.14fF
C2001 VDD.n1521 GND 0.17fF
C2002 VDD.n1522 GND 0.01fF
C2003 VDD.n1523 GND 0.02fF
C2004 VDD.n1524 GND 0.02fF
C2005 VDD.n1525 GND 0.22fF
C2006 VDD.n1526 GND 0.01fF
C2007 VDD.n1527 GND 0.07fF
C2008 VDD.n1528 GND 0.02fF
C2009 VDD.n1529 GND 0.27fF
C2010 VDD.n1530 GND 0.01fF
C2011 VDD.n1531 GND 0.02fF
C2012 VDD.n1532 GND 0.02fF
C2013 VDD.n1533 GND 0.27fF
C2014 VDD.n1534 GND 0.01fF
C2015 VDD.n1535 GND 0.02fF
C2016 VDD.n1536 GND 0.03fF
C2017 VDD.n1537 GND 0.02fF
C2018 VDD.n1538 GND 0.02fF
C2019 VDD.n1539 GND 0.02fF
C2020 VDD.n1540 GND 0.31fF
C2021 VDD.n1541 GND 0.04fF
C2022 VDD.n1542 GND 0.03fF
C2023 VDD.n1543 GND 0.02fF
C2024 VDD.n1544 GND 0.02fF
C2025 VDD.n1545 GND 0.02fF
C2026 VDD.n1546 GND 0.03fF
C2027 VDD.n1547 GND 0.02fF
C2028 VDD.n1549 GND 0.02fF
C2029 VDD.n1550 GND 0.02fF
C2030 VDD.n1551 GND 0.02fF
C2031 VDD.n1553 GND 0.27fF
C2032 VDD.n1555 GND 0.02fF
C2033 VDD.n1556 GND 0.02fF
C2034 VDD.n1557 GND 0.03fF
C2035 VDD.n1558 GND 0.02fF
C2036 VDD.n1559 GND 0.27fF
C2037 VDD.n1560 GND 0.01fF
C2038 VDD.n1561 GND 0.02fF
C2039 VDD.n1562 GND 0.03fF
C2040 VDD.n1563 GND 0.27fF
C2041 VDD.n1564 GND 0.01fF
C2042 VDD.n1565 GND 0.02fF
C2043 VDD.n1566 GND 0.02fF
C2044 VDD.n1567 GND 0.06fF
C2045 VDD.n1568 GND 0.23fF
C2046 VDD.n1569 GND 0.01fF
C2047 VDD.n1570 GND 0.01fF
C2048 VDD.n1571 GND 0.02fF
C2049 RN.n0 GND 0.89fF
C2050 RN.t22 GND 0.81fF
C2051 RN.n1 GND 0.68fF
C2052 RN.n2 GND 0.86fF
C2053 RN.t11 GND 0.82fF
C2054 RN.n3 GND 0.66fF
C2055 RN.n4 GND 2.38fF
C2056 RN.n5 GND 0.86fF
C2057 RN.t20 GND 0.83fF
C2058 RN.n6 GND 0.66fF
C2059 RN.n7 GND 3.35fF
C2060 RN.n8 GND 0.89fF
C2061 RN.t4 GND 0.81fF
C2062 RN.n9 GND 0.66fF
C2063 RN.n10 GND 2.69fF
C2064 RN.n11 GND 0.86fF
C2065 RN.t26 GND 0.82fF
C2066 RN.n12 GND 0.66fF
C2067 RN.n13 GND 1.80fF
C2068 RN.n14 GND 0.86fF
C2069 RN.t2 GND 0.83fF
C2070 RN.n15 GND 0.66fF
C2071 RN.n16 GND 3.35fF
C2072 RN.n17 GND 0.89fF
C2073 RN.t18 GND 0.81fF
C2074 RN.n18 GND 0.66fF
C2075 RN.n19 GND 2.69fF
C2076 RN.n20 GND 0.86fF
C2077 RN.t7 GND 0.82fF
C2078 RN.n21 GND 0.66fF
C2079 RN.n22 GND 1.80fF
C2080 RN.n23 GND 0.86fF
C2081 RN.t16 GND 0.83fF
C2082 RN.n24 GND 0.66fF
C2083 RN.n25 GND 1.25fF
C2084 a_12396_101.n0 GND 0.02fF
C2085 a_12396_101.n1 GND 0.10fF
C2086 a_12396_101.n2 GND 0.07fF
C2087 a_12396_101.n3 GND 0.05fF
C2088 a_12396_101.n4 GND 0.00fF
C2089 a_12396_101.n5 GND 0.04fF
C2090 a_12396_101.n6 GND 0.05fF
C2091 a_12396_101.n7 GND 0.02fF
C2092 a_12396_101.n8 GND 0.05fF
C2093 a_12396_101.n9 GND 0.02fF
C2094 a_12396_101.n10 GND 0.08fF
C2095 a_12396_101.n11 GND 0.17fF
C2096 a_12396_101.t1 GND 0.23fF
C2097 a_12396_101.n12 GND 0.09fF
C2098 a_12396_101.n13 GND 0.00fF
C2099 a_10959_989.n0 GND 0.75fF
C2100 a_10959_989.n1 GND 0.75fF
C2101 a_10959_989.n2 GND 0.88fF
C2102 a_10959_989.n3 GND 0.28fF
C2103 a_10959_989.n4 GND 0.43fF
C2104 a_10959_989.n5 GND 0.53fF
C2105 a_10959_989.n6 GND 0.55fF
C2106 a_10959_989.n7 GND 0.53fF
C2107 a_10959_989.t12 GND 0.75fF
C2108 a_10959_989.n8 GND 0.55fF
C2109 a_10959_989.n9 GND 1.75fF
C2110 a_10959_989.n10 GND 0.64fF
C2111 a_10959_989.n11 GND 0.12fF
C2112 a_10959_989.n12 GND 0.41fF
C2113 a_10959_989.n13 GND 0.06fF
.ends
