magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 130 582
<< pwell >>
rect 3 38 89 195
<< psubdiff >>
rect 29 145 63 169
rect 29 64 63 111
<< nsubdiff >>
rect 29 447 63 480
rect 29 363 63 413
rect 29 305 63 329
<< psubdiffcont >>
rect 29 111 63 145
<< nsubdiffcont >>
rect 29 413 63 447
rect 29 329 63 363
<< locali >>
rect 0 527 29 561
rect 63 527 92 561
rect 17 447 75 491
rect 17 413 29 447
rect 63 413 75 447
rect 17 391 75 413
rect 17 329 29 391
rect 63 329 75 391
rect 17 294 75 329
rect 17 145 75 162
rect 17 111 29 145
rect 63 111 75 145
rect 17 17 75 111
rect 0 -17 29 17
rect 63 -17 92 17
<< viali >>
rect 29 527 63 561
rect 29 363 63 391
rect 29 357 63 363
rect 29 -17 63 17
<< metal1 >>
rect 0 561 92 592
rect 0 527 29 561
rect 63 527 92 561
rect 0 496 92 527
rect 17 391 75 397
rect 17 357 29 391
rect 63 357 75 391
rect 17 351 75 357
rect 0 17 92 48
rect 0 -17 29 17
rect 63 -17 92 17
rect 0 -48 92 -17
<< labels >>
flabel locali s 32 358 61 382 0 FreeSans 250 0 0 0 VPB
port 2 nsew power bidirectional
flabel metal1 s 29 -14 61 13 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 29 533 67 552 0 FreeSans 200 0 0 0 VPWR
port 3 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 tapvgnd2_1
rlabel metal1 s 0 -48 92 48 1 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 0 496 92 592 1 VPWR
port 3 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE WELLTAP
string FIXED_BBOX 0 0 92 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 511010
string GDS_START 509202
string path 0.000 0.000 0.460 0.000 
<< end >>
