magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 1 21 1559 203
rect 30 -17 64 21
<< locali >>
rect 119 345 153 493
rect 287 345 321 493
rect 119 297 321 345
rect 119 263 153 297
rect 17 211 153 263
rect 423 211 616 263
rect 650 211 895 263
rect 931 211 1170 263
rect 1204 211 1354 263
rect 1390 211 1547 263
rect 119 177 153 211
rect 119 143 321 177
rect 119 51 153 143
rect 287 51 321 143
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 17 297 85 527
rect 187 379 253 527
rect 355 379 489 527
rect 523 345 557 493
rect 591 379 657 527
rect 691 345 725 493
rect 771 379 809 527
rect 867 459 1289 493
rect 867 379 933 459
rect 967 345 1001 425
rect 355 297 1001 345
rect 1051 297 1105 459
rect 1139 345 1189 425
rect 1223 379 1289 459
rect 1323 345 1357 425
rect 1391 379 1457 527
rect 1491 345 1547 493
rect 1139 297 1547 345
rect 355 263 389 297
rect 187 211 389 263
rect 355 177 389 211
rect 17 17 85 177
rect 355 143 609 177
rect 187 17 253 109
rect 439 135 609 143
rect 355 17 405 109
rect 643 101 677 177
rect 711 135 1547 177
rect 439 51 861 101
rect 897 51 951 135
rect 985 17 1121 101
rect 1155 51 1189 135
rect 1223 17 1289 101
rect 1323 51 1357 135
rect 1391 17 1457 101
rect 1491 51 1547 135
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
rlabel locali s 1390 211 1547 263 6 A1
port 1 nsew signal input
rlabel locali s 1204 211 1354 263 6 A2
port 2 nsew signal input
rlabel locali s 931 211 1170 263 6 A3
port 3 nsew signal input
rlabel locali s 650 211 895 263 6 B1
port 4 nsew signal input
rlabel locali s 423 211 616 263 6 C1
port 5 nsew signal input
rlabel metal1 s 0 -48 1564 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 1559 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1602 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 287 51 321 143 6 X
port 10 nsew signal output
rlabel locali s 119 51 153 143 6 X
port 10 nsew signal output
rlabel locali s 119 143 321 177 6 X
port 10 nsew signal output
rlabel locali s 119 177 153 211 6 X
port 10 nsew signal output
rlabel locali s 17 211 153 263 6 X
port 10 nsew signal output
rlabel locali s 119 263 153 297 6 X
port 10 nsew signal output
rlabel locali s 119 297 321 345 6 X
port 10 nsew signal output
rlabel locali s 287 345 321 493 6 X
port 10 nsew signal output
rlabel locali s 119 345 153 493 6 X
port 10 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1564 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 872304
string GDS_START 860012
<< end >>
