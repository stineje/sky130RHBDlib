// File: nand2x1_pcell.spi.NAND2X1_PCELL.pxi
// Created: Tue Oct 15 15:57:39 2024
// 
simulator lang=spectre
x_PM_NAND2X1_PCELL\%noxref_2 ( N_noxref_2_c_48_p N_noxref_2_c_25_p \
 N_noxref_2_c_34_p N_noxref_2_c_23_n N_noxref_2_c_24_n N_noxref_2_M2_noxref_s \
 N_noxref_2_M3_noxref_d N_noxref_2_M5_noxref_d )  PM_NAND2X1_PCELL\%noxref_2
x_PM_NAND2X1_PCELL\%noxref_3 ( N_noxref_3_c_58_n N_noxref_3_M0_noxref_g \
 N_noxref_3_M2_noxref_g N_noxref_3_M3_noxref_g N_noxref_3_c_59_n \
 N_noxref_3_c_60_n N_noxref_3_c_61_n N_noxref_3_c_62_n N_noxref_3_c_63_n \
 N_noxref_3_c_64_n N_noxref_3_c_65_n N_noxref_3_c_66_n N_noxref_3_c_73_n )  \
 PM_NAND2X1_PCELL\%noxref_3
x_PM_NAND2X1_PCELL\%noxref_4 ( N_noxref_4_c_119_n N_noxref_4_c_111_n \
 N_noxref_4_M1_noxref_g N_noxref_4_M4_noxref_g N_noxref_4_M5_noxref_g \
 N_noxref_4_c_126_n N_noxref_4_c_129_n N_noxref_4_c_131_n N_noxref_4_c_148_p \
 N_noxref_4_c_156_p N_noxref_4_c_144_p N_noxref_4_c_134_n N_noxref_4_c_135_n \
 N_noxref_4_c_136_n N_noxref_4_c_150_p N_noxref_4_c_138_n )  \
 PM_NAND2X1_PCELL\%noxref_4
x_PM_NAND2X1_PCELL\%noxref_5 ( N_noxref_5_c_175_n N_noxref_5_c_178_n \
 N_noxref_5_c_180_n N_noxref_5_c_172_n N_noxref_5_c_223_p N_noxref_5_c_173_n \
 N_noxref_5_c_212_n N_noxref_5_M1_noxref_d N_noxref_5_M2_noxref_d \
 N_noxref_5_M4_noxref_d )  PM_NAND2X1_PCELL\%noxref_5
x_PM_NAND2X1_PCELL\%noxref_6 ( N_noxref_6_c_235_n N_noxref_6_c_229_n \
 N_noxref_6_c_230_n N_noxref_6_c_231_n N_noxref_6_c_232_n N_noxref_6_c_233_n \
 N_noxref_6_M0_noxref_s )  PM_NAND2X1_PCELL\%noxref_6
cc_1 ( noxref_1 N_noxref_2_c_23_n ) capacitor c=0.00989031f //x=0.99 //y=0.865 \
 //x2=0.74 //y2=7.4
cc_2 ( noxref_1 N_noxref_2_c_24_n ) capacitor c=0.00989031f //x=0.99 //y=0.865 \
 //x2=2.59 //y2=7.4
cc_3 ( noxref_1 N_noxref_3_c_58_n ) capacitor c=0.0180518f //x=0.99 //y=0.865 \
 //x2=1.11 //y2=2.08
cc_4 ( noxref_1 N_noxref_3_c_59_n ) capacitor c=0.00355093f //x=0.99 //y=0.865 \
 //x2=0.915 //y2=0.865
cc_5 ( noxref_1 N_noxref_3_c_60_n ) capacitor c=0.00255985f //x=0.99 //y=0.865 \
 //x2=0.915 //y2=1.21
cc_6 ( noxref_1 N_noxref_3_c_61_n ) capacitor c=0.00264481f //x=0.99 //y=0.865 \
 //x2=0.915 //y2=1.52
cc_7 ( noxref_1 N_noxref_3_c_62_n ) capacitor c=0.0121947f //x=0.99 //y=0.865 \
 //x2=0.915 //y2=1.915
cc_8 ( noxref_1 N_noxref_3_c_63_n ) capacitor c=0.0131326f //x=0.99 //y=0.865 \
 //x2=1.29 //y2=0.71
cc_9 ( noxref_1 N_noxref_3_c_64_n ) capacitor c=0.00193127f //x=0.99 //y=0.865 \
 //x2=1.29 //y2=1.365
cc_10 ( noxref_1 N_noxref_3_c_65_n ) capacitor c=0.0038847f //x=0.99 //y=0.865 \
 //x2=1.445 //y2=0.865
cc_11 ( noxref_1 N_noxref_3_c_66_n ) capacitor c=0.00255985f //x=0.99 \
 //y=0.865 //x2=1.445 //y2=1.21
cc_12 ( noxref_1 N_noxref_4_c_111_n ) capacitor c=0.0018739f //x=0.99 \
 //y=0.865 //x2=1.85 //y2=2.08
cc_13 ( noxref_1 N_noxref_5_c_172_n ) capacitor c=0.0468439f //x=0.99 \
 //y=0.865 //x2=2.505 //y2=1.655
cc_14 ( noxref_1 N_noxref_5_c_173_n ) capacitor c=0.00101801f //x=0.99 \
 //y=0.865 //x2=2.59 //y2=5.115
cc_15 ( noxref_1 N_noxref_5_M1_noxref_d ) capacitor c=0.00847534f //x=0.99 \
 //y=0.865 //x2=1.96 //y2=0.905
cc_16 ( noxref_1 N_noxref_6_c_229_n ) capacitor c=0.0191305f //x=0.99 \
 //y=0.865 //x2=1.58 //y2=1.58
cc_17 ( noxref_1 N_noxref_6_c_230_n ) capacitor c=0.0571275f //x=0.99 \
 //y=0.865 //x2=1.665 //y2=0.615
cc_18 ( noxref_1 N_noxref_6_c_231_n ) capacitor c=2.91423e-19 //x=0.99 \
 //y=0.865 //x2=1.665 //y2=1.495
cc_19 ( noxref_1 N_noxref_6_c_232_n ) capacitor c=0.0599977f //x=0.99 \
 //y=0.865 //x2=2.55 //y2=0.53
cc_20 ( noxref_1 N_noxref_6_c_233_n ) capacitor c=0.0670542f //x=0.99 \
 //y=0.865 //x2=2.635 //y2=0.615
cc_21 ( noxref_1 N_noxref_6_M0_noxref_s ) capacitor c=0.118126f //x=0.99 \
 //y=0.865 //x2=0.56 //y2=0.365
cc_22 ( N_noxref_2_c_25_p N_noxref_3_c_58_n ) capacitor c=3.97183e-19 \
 //x=1.585 //y=7.4 //x2=1.11 //y2=2.08
cc_23 ( N_noxref_2_c_23_n N_noxref_3_c_58_n ) capacitor c=0.016845f //x=0.74 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_24 ( N_noxref_2_c_25_p N_noxref_3_M2_noxref_g ) capacitor c=0.00726866f \
 //x=1.585 //y=7.4 //x2=1.01 //y2=6.02
cc_25 ( N_noxref_2_M2_noxref_s N_noxref_3_M2_noxref_g ) capacitor c=0.054195f \
 //x=0.655 //y=5.02 //x2=1.01 //y2=6.02
cc_26 ( N_noxref_2_c_25_p N_noxref_3_M3_noxref_g ) capacitor c=0.00672952f \
 //x=1.585 //y=7.4 //x2=1.45 //y2=6.02
cc_27 ( N_noxref_2_M3_noxref_d N_noxref_3_M3_noxref_g ) capacitor c=0.015318f \
 //x=1.525 //y=5.02 //x2=1.45 //y2=6.02
cc_28 ( N_noxref_2_c_23_n N_noxref_3_c_73_n ) capacitor c=0.0292267f //x=0.74 \
 //y=7.4 //x2=1.11 //y2=4.7
cc_29 ( N_noxref_2_c_23_n N_noxref_4_c_111_n ) capacitor c=6.61004e-19 \
 //x=0.74 //y=7.4 //x2=1.85 //y2=2.08
cc_30 ( N_noxref_2_c_24_n N_noxref_4_c_111_n ) capacitor c=6.09526e-19 \
 //x=2.59 //y=7.4 //x2=1.85 //y2=2.08
cc_31 ( N_noxref_2_c_34_p N_noxref_4_M4_noxref_g ) capacitor c=0.00673971f \
 //x=2.465 //y=7.4 //x2=1.89 //y2=6.02
cc_32 ( N_noxref_2_M3_noxref_d N_noxref_4_M4_noxref_g ) capacitor c=0.015318f \
 //x=1.525 //y=5.02 //x2=1.89 //y2=6.02
cc_33 ( N_noxref_2_c_34_p N_noxref_4_M5_noxref_g ) capacitor c=0.00672952f \
 //x=2.465 //y=7.4 //x2=2.33 //y2=6.02
cc_34 ( N_noxref_2_c_24_n N_noxref_4_M5_noxref_g ) capacitor c=0.024326f \
 //x=2.59 //y=7.4 //x2=2.33 //y2=6.02
cc_35 ( N_noxref_2_M5_noxref_d N_noxref_4_M5_noxref_g ) capacitor c=0.0430452f \
 //x=2.405 //y=5.02 //x2=2.33 //y2=6.02
cc_36 ( N_noxref_2_c_25_p N_noxref_5_c_175_n ) capacitor c=5.76712e-19 \
 //x=1.585 //y=7.4 //x2=2.025 //y2=5.2
cc_37 ( N_noxref_2_c_34_p N_noxref_5_c_175_n ) capacitor c=5.76712e-19 \
 //x=2.465 //y=7.4 //x2=2.025 //y2=5.2
cc_38 ( N_noxref_2_M3_noxref_d N_noxref_5_c_175_n ) capacitor c=0.0132775f \
 //x=1.525 //y=5.02 //x2=2.025 //y2=5.2
cc_39 ( N_noxref_2_c_23_n N_noxref_5_c_178_n ) capacitor c=0.00989999f \
 //x=0.74 //y=7.4 //x2=1.315 //y2=5.2
cc_40 ( N_noxref_2_M2_noxref_s N_noxref_5_c_178_n ) capacitor c=0.087833f \
 //x=0.655 //y=5.02 //x2=1.315 //y2=5.2
cc_41 ( N_noxref_2_c_34_p N_noxref_5_c_180_n ) capacitor c=8.71806e-19 \
 //x=2.465 //y=7.4 //x2=2.505 //y2=5.2
cc_42 ( N_noxref_2_M5_noxref_d N_noxref_5_c_180_n ) capacitor c=0.0167784f \
 //x=2.405 //y=5.02 //x2=2.505 //y2=5.2
cc_43 ( N_noxref_2_c_23_n N_noxref_5_c_173_n ) capacitor c=0.00159771f \
 //x=0.74 //y=7.4 //x2=2.59 //y2=5.115
cc_44 ( N_noxref_2_c_24_n N_noxref_5_c_173_n ) capacitor c=0.0468798f //x=2.59 \
 //y=7.4 //x2=2.59 //y2=5.115
cc_45 ( N_noxref_2_c_48_p N_noxref_5_M2_noxref_d ) capacitor c=0.00719513f \
 //x=2.59 //y=7.4 //x2=1.085 //y2=5.02
cc_46 ( N_noxref_2_c_25_p N_noxref_5_M2_noxref_d ) capacitor c=0.0138103f \
 //x=1.585 //y=7.4 //x2=1.085 //y2=5.02
cc_47 ( N_noxref_2_c_24_n N_noxref_5_M2_noxref_d ) capacitor c=0.00204676f \
 //x=2.59 //y=7.4 //x2=1.085 //y2=5.02
cc_48 ( N_noxref_2_M3_noxref_d N_noxref_5_M2_noxref_d ) capacitor c=0.0664752f \
 //x=1.525 //y=5.02 //x2=1.085 //y2=5.02
cc_49 ( N_noxref_2_c_48_p N_noxref_5_M4_noxref_d ) capacitor c=0.00719513f \
 //x=2.59 //y=7.4 //x2=1.965 //y2=5.02
cc_50 ( N_noxref_2_c_34_p N_noxref_5_M4_noxref_d ) capacitor c=0.0138379f \
 //x=2.465 //y=7.4 //x2=1.965 //y2=5.02
cc_51 ( N_noxref_2_c_24_n N_noxref_5_M4_noxref_d ) capacitor c=0.0136712f \
 //x=2.59 //y=7.4 //x2=1.965 //y2=5.02
cc_52 ( N_noxref_2_M2_noxref_s N_noxref_5_M4_noxref_d ) capacitor \
 c=0.00111971f //x=0.655 //y=5.02 //x2=1.965 //y2=5.02
cc_53 ( N_noxref_2_M3_noxref_d N_noxref_5_M4_noxref_d ) capacitor c=0.0664752f \
 //x=1.525 //y=5.02 //x2=1.965 //y2=5.02
cc_54 ( N_noxref_2_M5_noxref_d N_noxref_5_M4_noxref_d ) capacitor c=0.0664752f \
 //x=2.405 //y=5.02 //x2=1.965 //y2=5.02
cc_55 ( N_noxref_3_c_58_n N_noxref_4_c_119_n ) capacitor c=0.00400249f \
 //x=1.11 //y=2.08 //x2=1.85 //y2=4.535
cc_56 ( N_noxref_3_c_73_n N_noxref_4_c_119_n ) capacitor c=0.00417994f \
 //x=1.11 //y=4.7 //x2=1.85 //y2=4.535
cc_57 ( N_noxref_3_c_58_n N_noxref_4_c_111_n ) capacitor c=0.0892371f //x=1.11 \
 //y=2.08 //x2=1.85 //y2=2.08
cc_58 ( N_noxref_3_c_62_n N_noxref_4_c_111_n ) capacitor c=0.00308814f \
 //x=0.915 //y=1.915 //x2=1.85 //y2=2.08
cc_59 ( N_noxref_3_M2_noxref_g N_noxref_4_M4_noxref_g ) capacitor c=0.0104611f \
 //x=1.01 //y=6.02 //x2=1.89 //y2=6.02
cc_60 ( N_noxref_3_M3_noxref_g N_noxref_4_M4_noxref_g ) capacitor c=0.106811f \
 //x=1.45 //y=6.02 //x2=1.89 //y2=6.02
cc_61 ( N_noxref_3_M3_noxref_g N_noxref_4_M5_noxref_g ) capacitor c=0.0100341f \
 //x=1.45 //y=6.02 //x2=2.33 //y2=6.02
cc_62 ( N_noxref_3_c_59_n N_noxref_4_c_126_n ) capacitor c=4.86506e-19 \
 //x=0.915 //y=0.865 //x2=1.885 //y2=0.905
cc_63 ( N_noxref_3_c_60_n N_noxref_4_c_126_n ) capacitor c=0.00152104f \
 //x=0.915 //y=1.21 //x2=1.885 //y2=0.905
cc_64 ( N_noxref_3_c_65_n N_noxref_4_c_126_n ) capacitor c=0.0151475f \
 //x=1.445 //y=0.865 //x2=1.885 //y2=0.905
cc_65 ( N_noxref_3_c_61_n N_noxref_4_c_129_n ) capacitor c=0.00109982f \
 //x=0.915 //y=1.52 //x2=1.885 //y2=1.25
cc_66 ( N_noxref_3_c_66_n N_noxref_4_c_129_n ) capacitor c=0.0111064f \
 //x=1.445 //y=1.21 //x2=1.885 //y2=1.25
cc_67 ( N_noxref_3_c_61_n N_noxref_4_c_131_n ) capacitor c=9.57794e-19 \
 //x=0.915 //y=1.52 //x2=1.885 //y2=1.56
cc_68 ( N_noxref_3_c_62_n N_noxref_4_c_131_n ) capacitor c=0.00662747f \
 //x=0.915 //y=1.915 //x2=1.885 //y2=1.56
cc_69 ( N_noxref_3_c_66_n N_noxref_4_c_131_n ) capacitor c=0.00862358f \
 //x=1.445 //y=1.21 //x2=1.885 //y2=1.56
cc_70 ( N_noxref_3_c_65_n N_noxref_4_c_134_n ) capacitor c=0.00124821f \
 //x=1.445 //y=0.865 //x2=2.415 //y2=0.905
cc_71 ( N_noxref_3_c_66_n N_noxref_4_c_135_n ) capacitor c=0.00200715f \
 //x=1.445 //y=1.21 //x2=2.415 //y2=1.25
cc_72 ( N_noxref_3_c_58_n N_noxref_4_c_136_n ) capacitor c=0.00307062f \
 //x=1.11 //y=2.08 //x2=1.85 //y2=2.08
cc_73 ( N_noxref_3_c_62_n N_noxref_4_c_136_n ) capacitor c=0.0179092f \
 //x=0.915 //y=1.915 //x2=1.85 //y2=2.08
cc_74 ( N_noxref_3_c_58_n N_noxref_4_c_138_n ) capacitor c=0.00344981f \
 //x=1.11 //y=2.08 //x2=1.88 //y2=4.7
cc_75 ( N_noxref_3_c_73_n N_noxref_4_c_138_n ) capacitor c=0.0293367f //x=1.11 \
 //y=4.7 //x2=1.88 //y2=4.7
cc_76 ( N_noxref_3_M3_noxref_g N_noxref_5_c_175_n ) capacitor c=0.0204115f \
 //x=1.45 //y=6.02 //x2=2.025 //y2=5.2
cc_77 ( N_noxref_3_c_58_n N_noxref_5_c_178_n ) capacitor c=0.0055959f //x=1.11 \
 //y=2.08 //x2=1.315 //y2=5.2
cc_78 ( N_noxref_3_M2_noxref_g N_noxref_5_c_178_n ) capacitor c=0.0177326f \
 //x=1.01 //y=6.02 //x2=1.315 //y2=5.2
cc_79 ( N_noxref_3_c_73_n N_noxref_5_c_178_n ) capacitor c=0.00605692f \
 //x=1.11 //y=4.7 //x2=1.315 //y2=5.2
cc_80 ( N_noxref_3_c_58_n N_noxref_5_c_173_n ) capacitor c=0.00396426f \
 //x=1.11 //y=2.08 //x2=2.59 //y2=5.115
cc_81 ( N_noxref_3_M3_noxref_g N_noxref_5_M2_noxref_d ) capacitor c=0.0173476f \
 //x=1.45 //y=6.02 //x2=1.085 //y2=5.02
cc_82 ( N_noxref_3_c_62_n N_noxref_6_c_235_n ) capacitor c=0.0034165f \
 //x=0.915 //y=1.915 //x2=0.695 //y2=1.495
cc_83 ( N_noxref_3_c_58_n N_noxref_6_c_229_n ) capacitor c=0.0118986f //x=1.11 \
 //y=2.08 //x2=1.58 //y2=1.58
cc_84 ( N_noxref_3_c_61_n N_noxref_6_c_229_n ) capacitor c=0.00703567f \
 //x=0.915 //y=1.52 //x2=1.58 //y2=1.58
cc_85 ( N_noxref_3_c_62_n N_noxref_6_c_229_n ) capacitor c=0.0216532f \
 //x=0.915 //y=1.915 //x2=1.58 //y2=1.58
cc_86 ( N_noxref_3_c_64_n N_noxref_6_c_229_n ) capacitor c=0.00780629f \
 //x=1.29 //y=1.365 //x2=1.58 //y2=1.58
cc_87 ( N_noxref_3_c_66_n N_noxref_6_c_229_n ) capacitor c=0.00339872f \
 //x=1.445 //y=1.21 //x2=1.58 //y2=1.58
cc_88 ( N_noxref_3_c_62_n N_noxref_6_c_231_n ) capacitor c=6.71402e-19 \
 //x=0.915 //y=1.915 //x2=1.665 //y2=1.495
cc_89 ( N_noxref_3_c_59_n N_noxref_6_M0_noxref_s ) capacitor c=0.0326577f \
 //x=0.915 //y=0.865 //x2=0.56 //y2=0.365
cc_90 ( N_noxref_3_c_61_n N_noxref_6_M0_noxref_s ) capacitor c=3.48408e-19 \
 //x=0.915 //y=1.52 //x2=0.56 //y2=0.365
cc_91 ( N_noxref_3_c_65_n N_noxref_6_M0_noxref_s ) capacitor c=0.0120759f \
 //x=1.445 //y=0.865 //x2=0.56 //y2=0.365
cc_92 ( N_noxref_4_c_119_n N_noxref_5_c_175_n ) capacitor c=0.0127867f \
 //x=1.85 //y=4.535 //x2=2.025 //y2=5.2
cc_93 ( N_noxref_4_M4_noxref_g N_noxref_5_c_175_n ) capacitor c=0.0166699f \
 //x=1.89 //y=6.02 //x2=2.025 //y2=5.2
cc_94 ( N_noxref_4_c_138_n N_noxref_5_c_175_n ) capacitor c=0.00399417f \
 //x=1.88 //y=4.7 //x2=2.025 //y2=5.2
cc_95 ( N_noxref_4_M5_noxref_g N_noxref_5_c_180_n ) capacitor c=0.0223814f \
 //x=2.33 //y=6.02 //x2=2.505 //y2=5.2
cc_96 ( N_noxref_4_c_144_p N_noxref_5_c_172_n ) capacitor c=0.00359704f \
 //x=2.26 //y=1.405 //x2=2.505 //y2=1.655
cc_97 ( N_noxref_4_c_135_n N_noxref_5_c_172_n ) capacitor c=0.00457401f \
 //x=2.415 //y=1.25 //x2=2.505 //y2=1.655
cc_98 ( N_noxref_4_c_119_n N_noxref_5_c_173_n ) capacitor c=0.0101115f \
 //x=1.85 //y=4.535 //x2=2.59 //y2=5.115
cc_99 ( N_noxref_4_c_111_n N_noxref_5_c_173_n ) capacitor c=0.0840845f \
 //x=1.85 //y=2.08 //x2=2.59 //y2=5.115
cc_100 ( N_noxref_4_c_148_p N_noxref_5_c_173_n ) capacitor c=0.0142673f \
 //x=2.255 //y=4.79 //x2=2.59 //y2=5.115
cc_101 ( N_noxref_4_c_136_n N_noxref_5_c_173_n ) capacitor c=0.00877984f \
 //x=1.85 //y=2.08 //x2=2.59 //y2=5.115
cc_102 ( N_noxref_4_c_150_p N_noxref_5_c_173_n ) capacitor c=0.00306024f \
 //x=1.85 //y=1.915 //x2=2.59 //y2=5.115
cc_103 ( N_noxref_4_c_138_n N_noxref_5_c_173_n ) capacitor c=0.00533692f \
 //x=1.88 //y=4.7 //x2=2.59 //y2=5.115
cc_104 ( N_noxref_4_c_148_p N_noxref_5_c_212_n ) capacitor c=0.00421574f \
 //x=2.255 //y=4.79 //x2=2.11 //y2=5.2
cc_105 ( N_noxref_4_c_126_n N_noxref_5_M1_noxref_d ) capacitor c=0.00217566f \
 //x=1.885 //y=0.905 //x2=1.96 //y2=0.905
cc_106 ( N_noxref_4_c_129_n N_noxref_5_M1_noxref_d ) capacitor c=0.0034598f \
 //x=1.885 //y=1.25 //x2=1.96 //y2=0.905
cc_107 ( N_noxref_4_c_131_n N_noxref_5_M1_noxref_d ) capacitor c=0.0065582f \
 //x=1.885 //y=1.56 //x2=1.96 //y2=0.905
cc_108 ( N_noxref_4_c_156_p N_noxref_5_M1_noxref_d ) capacitor c=0.00241102f \
 //x=2.26 //y=0.75 //x2=1.96 //y2=0.905
cc_109 ( N_noxref_4_c_144_p N_noxref_5_M1_noxref_d ) capacitor c=0.0138845f \
 //x=2.26 //y=1.405 //x2=1.96 //y2=0.905
cc_110 ( N_noxref_4_c_134_n N_noxref_5_M1_noxref_d ) capacitor c=0.00132245f \
 //x=2.415 //y=0.905 //x2=1.96 //y2=0.905
cc_111 ( N_noxref_4_c_135_n N_noxref_5_M1_noxref_d ) capacitor c=0.00566463f \
 //x=2.415 //y=1.25 //x2=1.96 //y2=0.905
cc_112 ( N_noxref_4_c_150_p N_noxref_5_M1_noxref_d ) capacitor c=0.00660593f \
 //x=1.85 //y=1.915 //x2=1.96 //y2=0.905
cc_113 ( N_noxref_4_M4_noxref_g N_noxref_5_M4_noxref_d ) capacitor \
 c=0.0173476f //x=1.89 //y=6.02 //x2=1.965 //y2=5.02
cc_114 ( N_noxref_4_M5_noxref_g N_noxref_5_M4_noxref_d ) capacitor \
 c=0.0179769f //x=2.33 //y=6.02 //x2=1.965 //y2=5.02
cc_115 ( N_noxref_4_c_131_n N_noxref_6_c_231_n ) capacitor c=0.00623646f \
 //x=1.885 //y=1.56 //x2=1.665 //y2=1.495
cc_116 ( N_noxref_4_c_136_n N_noxref_6_c_231_n ) capacitor c=0.00172768f \
 //x=1.85 //y=2.08 //x2=1.665 //y2=1.495
cc_117 ( N_noxref_4_c_111_n N_noxref_6_c_232_n ) capacitor c=0.00161845f \
 //x=1.85 //y=2.08 //x2=2.55 //y2=0.53
cc_118 ( N_noxref_4_c_126_n N_noxref_6_c_232_n ) capacitor c=0.0186143f \
 //x=1.885 //y=0.905 //x2=2.55 //y2=0.53
cc_119 ( N_noxref_4_c_134_n N_noxref_6_c_232_n ) capacitor c=0.00656458f \
 //x=2.415 //y=0.905 //x2=2.55 //y2=0.53
cc_120 ( N_noxref_4_c_136_n N_noxref_6_c_232_n ) capacitor c=2.1838e-19 \
 //x=1.85 //y=2.08 //x2=2.55 //y2=0.53
cc_121 ( N_noxref_4_c_126_n N_noxref_6_M0_noxref_s ) capacitor c=0.00623646f \
 //x=1.885 //y=0.905 //x2=0.56 //y2=0.365
cc_122 ( N_noxref_4_c_134_n N_noxref_6_M0_noxref_s ) capacitor c=0.0143002f \
 //x=2.415 //y=0.905 //x2=0.56 //y2=0.365
cc_123 ( N_noxref_4_c_135_n N_noxref_6_M0_noxref_s ) capacitor c=0.00290153f \
 //x=2.415 //y=1.25 //x2=0.56 //y2=0.365
cc_124 ( N_noxref_5_c_223_p N_noxref_6_c_235_n ) capacitor c=3.15806e-19 \
 //x=2.235 //y=1.655 //x2=0.695 //y2=1.495
cc_125 ( N_noxref_5_c_223_p N_noxref_6_c_231_n ) capacitor c=0.0201674f \
 //x=2.235 //y=1.655 //x2=1.665 //y2=1.495
cc_126 ( N_noxref_5_c_172_n N_noxref_6_c_232_n ) capacitor c=0.00469114f \
 //x=2.505 //y=1.655 //x2=2.55 //y2=0.53
cc_127 ( N_noxref_5_M1_noxref_d N_noxref_6_c_232_n ) capacitor c=0.0118355f \
 //x=1.96 //y=0.905 //x2=2.55 //y2=0.53
cc_128 ( N_noxref_5_c_172_n N_noxref_6_M0_noxref_s ) capacitor c=0.0144625f \
 //x=2.505 //y=1.655 //x2=0.56 //y2=0.365
cc_129 ( N_noxref_5_M1_noxref_d N_noxref_6_M0_noxref_s ) capacitor \
 c=0.0437911f //x=1.96 //y=0.905 //x2=0.56 //y2=0.365
