* SPICE3 file created from MUX2X1.ext - technology: sky130A

.subckt MUX2X1 Y A0 A1 S VPB VNB
M1000 VPB.t2 a_787_383# a_661_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VPB.t5 a_185_182.t3 a_1327_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_661_1004.t1 a_787_383# VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t12 a_1453_383# a_1327_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_661_1004.t4 S VPB.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPB.t8 S a_185_182.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VNB a_661_1004.t5 a_1888_73.t0 nshort w=-1.605u l=1.765u
+  ad=1.6781p pd=12.81u as=0p ps=0u
M1007 a_1327_1004.t0 a_185_182.t5 VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPB.t4 a_1327_1004.t5 a_1993_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VNB a_185_182.t4 a_1222_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t6 S a_661_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1327_1004.t2 a_1453_383# VPB.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB.t10 a_661_1004.t6 a_1993_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VNB S a_556_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1993_1004.t3 a_661_1004.t7 VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_185_182.t0 S VPB.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1993_1004.t0 a_1327_1004.t7 VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 S a_787_383# 0.26fF
C1 VPB a_1453_383# 0.07fF
C2 VPB S 0.20fF
C3 VPB a_787_383# 0.07fF
R0 a_556_73.t0 a_556_73.n1 93.333
R1 a_556_73.n4 a_556_73.n2 55.07
R2 a_556_73.t0 a_556_73.n0 8.137
R3 a_556_73.n4 a_556_73.n3 4.619
R4 a_556_73.t0 a_556_73.n4 0.071
R5 a_661_1004.n3 a_661_1004.t6 480.392
R6 a_661_1004.n3 a_661_1004.t7 403.272
R7 a_661_1004.n4 a_661_1004.t5 240.421
R8 a_661_1004.n5 a_661_1004.n2 189.099
R9 a_661_1004.n7 a_661_1004.n5 174.055
R10 a_661_1004.n5 a_661_1004.n4 155.763
R11 a_661_1004.n4 a_661_1004.n3 135.047
R12 a_661_1004.n2 a_661_1004.n1 76.002
R13 a_661_1004.n7 a_661_1004.n6 15.218
R14 a_661_1004.n0 a_661_1004.t0 14.282
R15 a_661_1004.n0 a_661_1004.t1 14.282
R16 a_661_1004.n1 a_661_1004.t3 14.282
R17 a_661_1004.n1 a_661_1004.t4 14.282
R18 a_661_1004.n2 a_661_1004.n0 12.85
R19 a_661_1004.n8 a_661_1004.n7 12.014
R20 VPB VPB.n251 126.832
R21 VPB.n63 VPB.n61 94.117
R22 VPB.n225 VPB.n223 94.117
R23 VPB.n118 VPB.n116 94.117
R24 VPB.n196 VPB.n193 76
R25 VPB.n200 VPB.n199 76
R26 VPB.n227 VPB.n226 76
R27 VPB.n232 VPB.n231 76
R28 VPB.n244 VPB.n243 76
R29 VPB.n74 VPB.n73 68.979
R30 VPB.n67 VPB.n66 64.528
R31 VPB.n20 VPB.n19 61.764
R32 VPB.n207 VPB.n206 61.764
R33 VPB.n85 VPB.n84 61.764
R34 VPB.n77 VPB.t9 55.106
R35 VPB.n65 VPB.t8 55.106
R36 VPB.n53 VPB.t7 55.106
R37 VPB.n141 VPB.t0 55.106
R38 VPB.n108 VPB.t11 55.106
R39 VPB.n228 VPB.t2 55.106
R40 VPB.n123 VPB.t12 55.106
R41 VPB.n176 VPB.t4 55.106
R42 VPB.n173 VPB.n172 48.952
R43 VPB.n125 VPB.n124 48.952
R44 VPB.n37 VPB.n36 48.952
R45 VPB.n105 VPB.n104 44.502
R46 VPB.n138 VPB.n137 44.502
R47 VPB.n50 VPB.n49 44.502
R48 VPB.n44 VPB.n35 40.824
R49 VPB.n132 VPB.n78 40.824
R50 VPB.n167 VPB.n166 40.824
R51 VPB.n181 VPB.n180 35.118
R52 VPB.n248 VPB.n244 20.452
R53 VPB.n165 VPB.n162 20.452
R54 VPB.n169 VPB.n168 17.801
R55 VPB.n129 VPB.n128 17.801
R56 VPB.n41 VPB.n40 17.801
R57 VPB.n35 VPB.t1 14.282
R58 VPB.n35 VPB.t6 14.282
R59 VPB.n78 VPB.t13 14.282
R60 VPB.n78 VPB.t5 14.282
R61 VPB.n166 VPB.t3 14.282
R62 VPB.n166 VPB.t10 14.282
R63 VPB.n165 VPB.n164 13.653
R64 VPB.n164 VPB.n163 13.653
R65 VPB.n179 VPB.n178 13.653
R66 VPB.n178 VPB.n177 13.653
R67 VPB.n175 VPB.n174 13.653
R68 VPB.n174 VPB.n173 13.653
R69 VPB.n171 VPB.n170 13.653
R70 VPB.n170 VPB.n169 13.653
R71 VPB.n103 VPB.n102 13.653
R72 VPB.n102 VPB.n101 13.653
R73 VPB.n107 VPB.n106 13.653
R74 VPB.n106 VPB.n105 13.653
R75 VPB.n111 VPB.n110 13.653
R76 VPB.n110 VPB.n109 13.653
R77 VPB.n114 VPB.n113 13.653
R78 VPB.n113 VPB.n112 13.653
R79 VPB.n119 VPB.n118 13.653
R80 VPB.n118 VPB.n117 13.653
R81 VPB.n122 VPB.n121 13.653
R82 VPB.n121 VPB.n120 13.653
R83 VPB.n127 VPB.n126 13.653
R84 VPB.n126 VPB.n125 13.653
R85 VPB.n131 VPB.n130 13.653
R86 VPB.n130 VPB.n129 13.653
R87 VPB.n136 VPB.n135 13.653
R88 VPB.n135 VPB.n134 13.653
R89 VPB.n140 VPB.n139 13.653
R90 VPB.n139 VPB.n138 13.653
R91 VPB.n196 VPB.n195 13.653
R92 VPB.n195 VPB.n194 13.653
R93 VPB.n199 VPB.n198 13.653
R94 VPB.n198 VPB.n197 13.653
R95 VPB.n226 VPB.n225 13.653
R96 VPB.n225 VPB.n224 13.653
R97 VPB.n231 VPB.n230 13.653
R98 VPB.n230 VPB.n229 13.653
R99 VPB.n39 VPB.n38 13.653
R100 VPB.n38 VPB.n37 13.653
R101 VPB.n43 VPB.n42 13.653
R102 VPB.n42 VPB.n41 13.653
R103 VPB.n48 VPB.n47 13.653
R104 VPB.n47 VPB.n46 13.653
R105 VPB.n52 VPB.n51 13.653
R106 VPB.n51 VPB.n50 13.653
R107 VPB.n56 VPB.n55 13.653
R108 VPB.n55 VPB.n54 13.653
R109 VPB.n59 VPB.n58 13.653
R110 VPB.n58 VPB.n57 13.653
R111 VPB.n64 VPB.n63 13.653
R112 VPB.n63 VPB.n62 13.653
R113 VPB.n69 VPB.n68 13.653
R114 VPB.n68 VPB.n67 13.653
R115 VPB.n72 VPB.n71 13.653
R116 VPB.n71 VPB.n70 13.653
R117 VPB.n76 VPB.n75 13.653
R118 VPB.n75 VPB.n74 13.653
R119 VPB.n244 VPB.n0 13.653
R120 VPB VPB.n0 13.653
R121 VPB.n101 VPB.n100 13.35
R122 VPB.n134 VPB.n133 13.35
R123 VPB.n46 VPB.n45 13.35
R124 VPB.n248 VPB.n247 13.276
R125 VPB.n247 VPB.n245 13.276
R126 VPB.n34 VPB.n16 13.276
R127 VPB.n16 VPB.n14 13.276
R128 VPB.n221 VPB.n203 13.276
R129 VPB.n203 VPB.n201 13.276
R130 VPB.n99 VPB.n81 13.276
R131 VPB.n81 VPB.n79 13.276
R132 VPB.n175 VPB.n171 13.276
R133 VPB.n107 VPB.n103 13.276
R134 VPB.n114 VPB.n111 13.276
R135 VPB.n115 VPB.n114 13.276
R136 VPB.n119 VPB.n115 13.276
R137 VPB.n122 VPB.n119 13.276
R138 VPB.n131 VPB.n127 13.276
R139 VPB.n140 VPB.n136 13.276
R140 VPB.n199 VPB.n196 13.276
R141 VPB.n226 VPB.n222 13.276
R142 VPB.n43 VPB.n39 13.276
R143 VPB.n52 VPB.n48 13.276
R144 VPB.n59 VPB.n56 13.276
R145 VPB.n60 VPB.n59 13.276
R146 VPB.n64 VPB.n60 13.276
R147 VPB.n72 VPB.n69 13.276
R148 VPB.n76 VPB.n72 13.276
R149 VPB.n162 VPB.n144 13.276
R150 VPB.n144 VPB.n142 13.276
R151 VPB.n149 VPB.n147 12.796
R152 VPB.n149 VPB.n148 12.564
R153 VPB.n155 VPB.n154 12.198
R154 VPB.n157 VPB.n156 12.198
R155 VPB.n155 VPB.n152 12.198
R156 VPB.n176 VPB.n175 11.841
R157 VPB.n127 VPB.n123 11.841
R158 VPB.n108 VPB.n107 11.482
R159 VPB.n141 VPB.n140 11.482
R160 VPB.n53 VPB.n52 11.482
R161 VPB.n244 VPB.n77 10.944
R162 VPB.n65 VPB.n64 10.585
R163 VPB.n162 VPB.n161 7.5
R164 VPB.n147 VPB.n146 7.5
R165 VPB.n154 VPB.n153 7.5
R166 VPB.n152 VPB.n151 7.5
R167 VPB.n144 VPB.n143 7.5
R168 VPB.n159 VPB.n145 7.5
R169 VPB.n81 VPB.n80 7.5
R170 VPB.n94 VPB.n93 7.5
R171 VPB.n88 VPB.n87 7.5
R172 VPB.n90 VPB.n89 7.5
R173 VPB.n83 VPB.n82 7.5
R174 VPB.n99 VPB.n98 7.5
R175 VPB.n203 VPB.n202 7.5
R176 VPB.n216 VPB.n215 7.5
R177 VPB.n210 VPB.n209 7.5
R178 VPB.n212 VPB.n211 7.5
R179 VPB.n205 VPB.n204 7.5
R180 VPB.n221 VPB.n220 7.5
R181 VPB.n16 VPB.n15 7.5
R182 VPB.n29 VPB.n28 7.5
R183 VPB.n23 VPB.n22 7.5
R184 VPB.n25 VPB.n24 7.5
R185 VPB.n18 VPB.n17 7.5
R186 VPB.n34 VPB.n33 7.5
R187 VPB.n247 VPB.n246 7.5
R188 VPB.n12 VPB.n11 7.5
R189 VPB.n6 VPB.n5 7.5
R190 VPB.n8 VPB.n7 7.5
R191 VPB.n2 VPB.n1 7.5
R192 VPB.n249 VPB.n248 7.5
R193 VPB.n60 VPB.n34 7.176
R194 VPB.n222 VPB.n221 7.176
R195 VPB.n115 VPB.n99 7.176
R196 VPB.n136 VPB.n132 6.817
R197 VPB.n48 VPB.n44 6.817
R198 VPB.n95 VPB.n92 6.729
R199 VPB.n91 VPB.n88 6.729
R200 VPB.n86 VPB.n83 6.729
R201 VPB.n217 VPB.n214 6.729
R202 VPB.n213 VPB.n210 6.729
R203 VPB.n208 VPB.n205 6.729
R204 VPB.n30 VPB.n27 6.729
R205 VPB.n26 VPB.n23 6.729
R206 VPB.n21 VPB.n18 6.729
R207 VPB.n13 VPB.n10 6.729
R208 VPB.n9 VPB.n6 6.729
R209 VPB.n4 VPB.n2 6.729
R210 VPB.n86 VPB.n85 6.728
R211 VPB.n91 VPB.n90 6.728
R212 VPB.n95 VPB.n94 6.728
R213 VPB.n98 VPB.n97 6.728
R214 VPB.n208 VPB.n207 6.728
R215 VPB.n213 VPB.n212 6.728
R216 VPB.n217 VPB.n216 6.728
R217 VPB.n220 VPB.n219 6.728
R218 VPB.n21 VPB.n20 6.728
R219 VPB.n26 VPB.n25 6.728
R220 VPB.n30 VPB.n29 6.728
R221 VPB.n33 VPB.n32 6.728
R222 VPB.n4 VPB.n3 6.728
R223 VPB.n9 VPB.n8 6.728
R224 VPB.n13 VPB.n12 6.728
R225 VPB.n250 VPB.n249 6.728
R226 VPB.n171 VPB.n167 6.458
R227 VPB.n132 VPB.n131 6.458
R228 VPB.n44 VPB.n43 6.458
R229 VPB.n161 VPB.n160 6.398
R230 VPB.n180 VPB.n165 6.112
R231 VPB.n180 VPB.n179 6.101
R232 VPB.n69 VPB.n65 2.691
R233 VPB.n77 VPB.n76 2.332
R234 VPB.n111 VPB.n108 1.794
R235 VPB.n196 VPB.n141 1.794
R236 VPB.n56 VPB.n53 1.794
R237 VPB.n179 VPB.n176 1.435
R238 VPB.n123 VPB.n122 1.435
R239 VPB.n231 VPB.n228 1.435
R240 VPB.n159 VPB.n150 1.402
R241 VPB.n159 VPB.n155 1.402
R242 VPB.n159 VPB.n157 1.402
R243 VPB.n159 VPB.n158 1.402
R244 VPB.n160 VPB.n159 0.735
R245 VPB.n159 VPB.n149 0.735
R246 VPB.n96 VPB.n95 0.387
R247 VPB.n96 VPB.n91 0.387
R248 VPB.n96 VPB.n86 0.387
R249 VPB.n97 VPB.n96 0.387
R250 VPB.n218 VPB.n217 0.387
R251 VPB.n218 VPB.n213 0.387
R252 VPB.n218 VPB.n208 0.387
R253 VPB.n219 VPB.n218 0.387
R254 VPB.n31 VPB.n30 0.387
R255 VPB.n31 VPB.n26 0.387
R256 VPB.n31 VPB.n21 0.387
R257 VPB.n32 VPB.n31 0.387
R258 VPB.n251 VPB.n13 0.387
R259 VPB.n251 VPB.n9 0.387
R260 VPB.n251 VPB.n4 0.387
R261 VPB.n251 VPB.n250 0.387
R262 VPB.n187 VPB.n186 0.272
R263 VPB.n227 VPB.n200 0.272
R264 VPB.n239 VPB.n238 0.272
R265 VPB.n243 VPB 0.198
R266 VPB.n182 VPB.n181 0.136
R267 VPB.n183 VPB.n182 0.136
R268 VPB.n184 VPB.n183 0.136
R269 VPB.n185 VPB.n184 0.136
R270 VPB.n186 VPB.n185 0.136
R271 VPB.n188 VPB.n187 0.136
R272 VPB.n189 VPB.n188 0.136
R273 VPB.n190 VPB.n189 0.136
R274 VPB.n191 VPB.n190 0.136
R275 VPB.n192 VPB.n191 0.136
R276 VPB.n193 VPB.n192 0.136
R277 VPB.n232 VPB.n227 0.136
R278 VPB.n233 VPB.n232 0.136
R279 VPB.n234 VPB.n233 0.136
R280 VPB.n235 VPB.n234 0.136
R281 VPB.n236 VPB.n235 0.136
R282 VPB.n237 VPB.n236 0.136
R283 VPB.n238 VPB.n237 0.136
R284 VPB.n240 VPB.n239 0.136
R285 VPB.n241 VPB.n240 0.136
R286 VPB.n242 VPB.n241 0.136
R287 VPB.n243 VPB.n242 0.136
R288 VPB.n193 VPB 0.068
R289 VPB.n200 VPB 0.068
R290 a_185_182.n2 a_185_182.t3 480.392
R291 a_185_182.n2 a_185_182.t5 403.272
R292 a_185_182.n3 a_185_182.t4 266.974
R293 a_185_182.n6 a_185_182.n4 188.704
R294 a_185_182.n4 a_185_182.n1 167.143
R295 a_185_182.n4 a_185_182.n3 155.763
R296 a_185_182.n3 a_185_182.n2 108.494
R297 a_185_182.n6 a_185_182.n5 30
R298 a_185_182.n7 a_185_182.n0 24.383
R299 a_185_182.n7 a_185_182.n6 23.684
R300 a_185_182.n1 a_185_182.t1 14.282
R301 a_185_182.n1 a_185_182.t0 14.282
R302 a_1327_1004.n4 a_1327_1004.t5 472.359
R303 a_1327_1004.n4 a_1327_1004.t7 384.527
R304 a_1327_1004.n5 a_1327_1004.t6 224.666
R305 a_1327_1004.n8 a_1327_1004.n6 194.086
R306 a_1327_1004.n6 a_1327_1004.n3 162.547
R307 a_1327_1004.n6 a_1327_1004.n5 153.859
R308 a_1327_1004.n5 a_1327_1004.n4 120.107
R309 a_1327_1004.n3 a_1327_1004.n2 76.002
R310 a_1327_1004.n8 a_1327_1004.n7 30
R311 a_1327_1004.n9 a_1327_1004.n0 24.383
R312 a_1327_1004.n9 a_1327_1004.n8 23.684
R313 a_1327_1004.n1 a_1327_1004.t3 14.282
R314 a_1327_1004.n1 a_1327_1004.t2 14.282
R315 a_1327_1004.n2 a_1327_1004.t1 14.282
R316 a_1327_1004.n2 a_1327_1004.t0 14.282
R317 a_1327_1004.n3 a_1327_1004.n1 12.85
R318 a_1888_73.t0 a_1888_73.n1 93.333
R319 a_1888_73.n4 a_1888_73.n2 55.07
R320 a_1888_73.t0 a_1888_73.n0 8.137
R321 a_1888_73.n4 a_1888_73.n3 4.619
R322 a_1888_73.t0 a_1888_73.n4 0.071
R323 VNB VNB.n225 300.778
R324 VNB.n82 VNB.n81 199.897
R325 VNB.n185 VNB.n184 199.897
R326 VNB.n25 VNB.n24 199.897
R327 VNB.n194 VNB.n192 154.509
R328 VNB.n105 VNB.n103 154.509
R329 VNB.n54 VNB.n52 154.509
R330 VNB.n117 VNB.n116 121.366
R331 VNB.n92 VNB.n88 84.842
R332 VNB.n41 VNB.n31 84.842
R333 VNB.n212 VNB.n211 76
R334 VNB.n200 VNB.n199 76
R335 VNB.n196 VNB.n195 76
R336 VNB.n174 VNB.n173 76
R337 VNB.n170 VNB.n167 76
R338 VNB.n121 VNB.n71 63.835
R339 VNB.n62 VNB.n61 49.896
R340 VNB.n118 VNB.n117 36.937
R341 VNB.n94 VNB.n93 36.678
R342 VNB.n43 VNB.n42 36.678
R343 VNB.n155 VNB.n154 35.118
R344 VNB.n14 VNB.n13 35.01
R345 VNB.t1 VNB.n6 32.601
R346 VNB.n71 VNB.n70 28.421
R347 VNB.n124 VNB.n123 27.855
R348 VNB.n71 VNB.n69 25.263
R349 VNB.n69 VNB.n68 24.383
R350 VNB.n144 VNB.n141 20.452
R351 VNB.n213 VNB.n212 20.452
R352 VNB.n56 VNB.n14 20.094
R353 VNB.n60 VNB.n11 20.094
R354 VNB.n67 VNB.n9 20.094
R355 VNB.n14 VNB.n12 19.017
R356 VNB.n8 VNB.t1 17.353
R357 VNB.n125 VNB.n124 16.721
R358 VNB.n153 VNB.n152 13.653
R359 VNB.n152 VNB.n151 13.653
R360 VNB.n150 VNB.n149 13.653
R361 VNB.n149 VNB.n148 13.653
R362 VNB.n147 VNB.n146 13.653
R363 VNB.n146 VNB.n145 13.653
R364 VNB.n91 VNB.n90 13.653
R365 VNB.n90 VNB.n89 13.653
R366 VNB.n95 VNB.n94 13.653
R367 VNB.n98 VNB.n97 13.653
R368 VNB.n97 VNB.n96 13.653
R369 VNB.n101 VNB.n100 13.653
R370 VNB.n100 VNB.n99 13.653
R371 VNB.n106 VNB.n105 13.653
R372 VNB.n105 VNB.n104 13.653
R373 VNB.n109 VNB.n108 13.653
R374 VNB.n108 VNB.n107 13.653
R375 VNB.n112 VNB.n111 13.653
R376 VNB.n111 VNB.n110 13.653
R377 VNB.n115 VNB.n114 13.653
R378 VNB.n114 VNB.n113 13.653
R379 VNB.n120 VNB.n119 13.653
R380 VNB.n119 VNB.n118 13.653
R381 VNB.n126 VNB.n125 13.653
R382 VNB.n170 VNB.n169 13.653
R383 VNB.n169 VNB.n168 13.653
R384 VNB.n173 VNB.n172 13.653
R385 VNB.n172 VNB.n171 13.653
R386 VNB.n195 VNB.n194 13.653
R387 VNB.n194 VNB.n193 13.653
R388 VNB.n199 VNB.n198 13.653
R389 VNB.n198 VNB.n197 13.653
R390 VNB.n34 VNB.n33 13.653
R391 VNB.n33 VNB.n32 13.653
R392 VNB.n37 VNB.n36 13.653
R393 VNB.n36 VNB.n35 13.653
R394 VNB.n40 VNB.n39 13.653
R395 VNB.n39 VNB.n38 13.653
R396 VNB.n44 VNB.n43 13.653
R397 VNB.n47 VNB.n46 13.653
R398 VNB.n46 VNB.n45 13.653
R399 VNB.n50 VNB.n49 13.653
R400 VNB.n49 VNB.n48 13.653
R401 VNB.n55 VNB.n54 13.653
R402 VNB.n54 VNB.n53 13.653
R403 VNB.n59 VNB.n58 13.653
R404 VNB.n58 VNB.n57 13.653
R405 VNB.n63 VNB.n62 13.653
R406 VNB.n66 VNB.n65 13.653
R407 VNB.n65 VNB.n64 13.653
R408 VNB.n212 VNB.n0 13.653
R409 VNB VNB.n0 13.653
R410 VNB.n144 VNB.n143 13.653
R411 VNB.n143 VNB.n142 13.653
R412 VNB.n220 VNB.n217 13.577
R413 VNB.n129 VNB.n127 13.276
R414 VNB.n141 VNB.n129 13.276
R415 VNB.n74 VNB.n72 13.276
R416 VNB.n87 VNB.n74 13.276
R417 VNB.n177 VNB.n175 13.276
R418 VNB.n190 VNB.n177 13.276
R419 VNB.n17 VNB.n15 13.276
R420 VNB.n30 VNB.n17 13.276
R421 VNB.n153 VNB.n150 13.276
R422 VNB.n150 VNB.n147 13.276
R423 VNB.n98 VNB.n95 13.276
R424 VNB.n101 VNB.n98 13.276
R425 VNB.n102 VNB.n101 13.276
R426 VNB.n106 VNB.n102 13.276
R427 VNB.n109 VNB.n106 13.276
R428 VNB.n112 VNB.n109 13.276
R429 VNB.n115 VNB.n112 13.276
R430 VNB.n120 VNB.n115 13.276
R431 VNB.n170 VNB.n126 13.276
R432 VNB.n173 VNB.n170 13.276
R433 VNB.n195 VNB.n191 13.276
R434 VNB.n37 VNB.n34 13.276
R435 VNB.n40 VNB.n37 13.276
R436 VNB.n47 VNB.n44 13.276
R437 VNB.n50 VNB.n47 13.276
R438 VNB.n51 VNB.n50 13.276
R439 VNB.n55 VNB.n51 13.276
R440 VNB.n66 VNB.n63 13.276
R441 VNB.n3 VNB.n1 13.276
R442 VNB.n213 VNB.n3 13.276
R443 VNB.n60 VNB.n59 13.097
R444 VNB.n9 VNB.n8 12.837
R445 VNB.n92 VNB.n91 10.764
R446 VNB.n121 VNB.n120 10.764
R447 VNB.n41 VNB.n40 10.764
R448 VNB.n212 VNB.n67 9.329
R449 VNB.n56 VNB.n55 8.97
R450 VNB.n8 VNB.n7 7.566
R451 VNB.n222 VNB.n221 7.5
R452 VNB.n80 VNB.n79 7.5
R453 VNB.n76 VNB.n75 7.5
R454 VNB.n74 VNB.n73 7.5
R455 VNB.n87 VNB.n86 7.5
R456 VNB.n183 VNB.n182 7.5
R457 VNB.n179 VNB.n178 7.5
R458 VNB.n177 VNB.n176 7.5
R459 VNB.n190 VNB.n189 7.5
R460 VNB.n23 VNB.n22 7.5
R461 VNB.n19 VNB.n18 7.5
R462 VNB.n17 VNB.n16 7.5
R463 VNB.n30 VNB.n29 7.5
R464 VNB.n214 VNB.n213 7.5
R465 VNB.n3 VNB.n2 7.5
R466 VNB.n219 VNB.n218 7.5
R467 VNB.n135 VNB.n134 7.5
R468 VNB.n131 VNB.n130 7.5
R469 VNB.n129 VNB.n128 7.5
R470 VNB.n141 VNB.n140 7.5
R471 VNB.n102 VNB.n87 7.176
R472 VNB.n191 VNB.n190 7.176
R473 VNB.n51 VNB.n30 7.176
R474 VNB.n224 VNB.n222 7.011
R475 VNB.n83 VNB.n80 7.011
R476 VNB.n78 VNB.n76 7.011
R477 VNB.n186 VNB.n183 7.011
R478 VNB.n181 VNB.n179 7.011
R479 VNB.n26 VNB.n23 7.011
R480 VNB.n21 VNB.n19 7.011
R481 VNB.n137 VNB.n135 7.011
R482 VNB.n133 VNB.n131 7.011
R483 VNB.n86 VNB.n85 7.01
R484 VNB.n78 VNB.n77 7.01
R485 VNB.n83 VNB.n82 7.01
R486 VNB.n189 VNB.n188 7.01
R487 VNB.n181 VNB.n180 7.01
R488 VNB.n186 VNB.n185 7.01
R489 VNB.n29 VNB.n28 7.01
R490 VNB.n21 VNB.n20 7.01
R491 VNB.n26 VNB.n25 7.01
R492 VNB.n140 VNB.n139 7.01
R493 VNB.n133 VNB.n132 7.01
R494 VNB.n137 VNB.n136 7.01
R495 VNB.n224 VNB.n223 7.01
R496 VNB.n220 VNB.n219 6.788
R497 VNB.n215 VNB.n214 6.788
R498 VNB.n154 VNB.n144 6.111
R499 VNB.n154 VNB.n153 6.1
R500 VNB.n5 VNB.n4 4.551
R501 VNB.n59 VNB.n56 4.305
R502 VNB.n67 VNB.n66 3.947
R503 VNB.n95 VNB.n92 2.511
R504 VNB.n126 VNB.n121 2.511
R505 VNB.n44 VNB.n41 2.511
R506 VNB.t1 VNB.n5 2.238
R507 VNB.n124 VNB.n122 1.99
R508 VNB.n225 VNB.n216 0.921
R509 VNB.n225 VNB.n220 0.476
R510 VNB.n225 VNB.n215 0.475
R511 VNB.n11 VNB.n10 0.358
R512 VNB.n161 VNB.n160 0.272
R513 VNB.n196 VNB.n174 0.272
R514 VNB.n207 VNB.n206 0.272
R515 VNB.n84 VNB.n78 0.246
R516 VNB.n85 VNB.n84 0.246
R517 VNB.n84 VNB.n83 0.246
R518 VNB.n187 VNB.n181 0.246
R519 VNB.n188 VNB.n187 0.246
R520 VNB.n187 VNB.n186 0.246
R521 VNB.n27 VNB.n21 0.246
R522 VNB.n28 VNB.n27 0.246
R523 VNB.n27 VNB.n26 0.246
R524 VNB.n138 VNB.n133 0.246
R525 VNB.n139 VNB.n138 0.246
R526 VNB.n138 VNB.n137 0.246
R527 VNB.n225 VNB.n224 0.246
R528 VNB.n211 VNB 0.198
R529 VNB.n63 VNB.n60 0.179
R530 VNB.n156 VNB.n155 0.136
R531 VNB.n157 VNB.n156 0.136
R532 VNB.n158 VNB.n157 0.136
R533 VNB.n159 VNB.n158 0.136
R534 VNB.n160 VNB.n159 0.136
R535 VNB.n162 VNB.n161 0.136
R536 VNB.n163 VNB.n162 0.136
R537 VNB.n164 VNB.n163 0.136
R538 VNB.n165 VNB.n164 0.136
R539 VNB.n166 VNB.n165 0.136
R540 VNB.n167 VNB.n166 0.136
R541 VNB.n200 VNB.n196 0.136
R542 VNB.n201 VNB.n200 0.136
R543 VNB.n202 VNB.n201 0.136
R544 VNB.n203 VNB.n202 0.136
R545 VNB.n204 VNB.n203 0.136
R546 VNB.n205 VNB.n204 0.136
R547 VNB.n206 VNB.n205 0.136
R548 VNB.n208 VNB.n207 0.136
R549 VNB.n209 VNB.n208 0.136
R550 VNB.n210 VNB.n209 0.136
R551 VNB.n211 VNB.n210 0.136
R552 VNB.n167 VNB 0.068
R553 VNB.n174 VNB 0.068
R554 a_1222_73.n12 a_1222_73.n11 26.811
R555 a_1222_73.n6 a_1222_73.n5 24.977
R556 a_1222_73.n2 a_1222_73.n1 24.877
R557 a_1222_73.t0 a_1222_73.n2 12.677
R558 a_1222_73.t0 a_1222_73.n3 11.595
R559 a_1222_73.t1 a_1222_73.n8 8.137
R560 a_1222_73.t0 a_1222_73.n4 7.273
R561 a_1222_73.t0 a_1222_73.n0 6.109
R562 a_1222_73.t1 a_1222_73.n7 4.864
R563 a_1222_73.t0 a_1222_73.n12 2.074
R564 a_1222_73.n7 a_1222_73.n6 1.13
R565 a_1222_73.n12 a_1222_73.t1 0.937
R566 a_1222_73.t1 a_1222_73.n10 0.804
R567 a_1222_73.n10 a_1222_73.n9 0.136
R568 a_1993_1004.n4 a_1993_1004.n2 363.155
R569 a_1993_1004.n2 a_1993_1004.n1 76.002
R570 a_1993_1004.n4 a_1993_1004.n3 15.218
R571 a_1993_1004.n0 a_1993_1004.t1 14.282
R572 a_1993_1004.n0 a_1993_1004.t0 14.282
R573 a_1993_1004.n1 a_1993_1004.t4 14.282
R574 a_1993_1004.n1 a_1993_1004.t3 14.282
R575 a_1993_1004.n2 a_1993_1004.n0 12.85
R576 a_1993_1004.n5 a_1993_1004.n4 12.014
C4 VPB VNB 10.41fF
C5 a_1993_1004.n0 VNB 0.47fF
C6 a_1993_1004.n1 VNB 0.56fF
C7 a_1993_1004.n2 VNB 0.49fF
C8 a_1993_1004.n3 VNB 0.07fF
C9 a_1993_1004.n4 VNB 0.41fF
C10 a_1993_1004.n5 VNB 0.04fF
C11 a_1222_73.n0 VNB 0.02fF
C12 a_1222_73.n1 VNB 0.10fF
C13 a_1222_73.n2 VNB 0.06fF
C14 a_1222_73.n3 VNB 0.06fF
C15 a_1222_73.n4 VNB 0.00fF
C16 a_1222_73.n5 VNB 0.04fF
C17 a_1222_73.n6 VNB 0.05fF
C18 a_1222_73.n7 VNB 0.02fF
C19 a_1222_73.n8 VNB 0.05fF
C20 a_1222_73.n9 VNB 0.08fF
C21 a_1222_73.n10 VNB 0.17fF
C22 a_1222_73.t1 VNB 0.23fF
C23 a_1222_73.n11 VNB 0.09fF
C24 a_1222_73.n12 VNB 0.00fF
C25 a_1888_73.n0 VNB 0.05fF
C26 a_1888_73.n1 VNB 0.02fF
C27 a_1888_73.n2 VNB 0.12fF
C28 a_1888_73.n3 VNB 0.04fF
C29 a_1888_73.n4 VNB 0.16fF
C30 a_1327_1004.n0 VNB 0.04fF
C31 a_1327_1004.n1 VNB 0.49fF
C32 a_1327_1004.n2 VNB 0.58fF
C33 a_1327_1004.n3 VNB 0.30fF
C34 a_1327_1004.n4 VNB 0.32fF
C35 a_1327_1004.t6 VNB 0.48fF
C36 a_1327_1004.n5 VNB 0.56fF
C37 a_1327_1004.n6 VNB 0.61fF
C38 a_1327_1004.n7 VNB 0.03fF
C39 a_1327_1004.n8 VNB 0.26fF
C40 a_1327_1004.n9 VNB 0.05fF
C41 a_185_182.n0 VNB 0.04fF
C42 a_185_182.n1 VNB 0.79fF
C43 a_185_182.n2 VNB 0.41fF
C44 a_185_182.n3 VNB 0.89fF
C45 a_185_182.n4 VNB 0.94fF
C46 a_185_182.n5 VNB 0.04fF
C47 a_185_182.n6 VNB 0.29fF
C48 a_185_182.n7 VNB 0.06fF
C49 VPB.n0 VNB 0.03fF
C50 VPB.n1 VNB 0.03fF
C51 VPB.n2 VNB 0.02fF
C52 VPB.n3 VNB 0.10fF
C53 VPB.n5 VNB 0.02fF
C54 VPB.n6 VNB 0.02fF
C55 VPB.n7 VNB 0.02fF
C56 VPB.n8 VNB 0.02fF
C57 VPB.n10 VNB 0.02fF
C58 VPB.n11 VNB 0.02fF
C59 VPB.n12 VNB 0.02fF
C60 VPB.n14 VNB 0.02fF
C61 VPB.n15 VNB 0.02fF
C62 VPB.n16 VNB 0.02fF
C63 VPB.n17 VNB 0.03fF
C64 VPB.n18 VNB 0.02fF
C65 VPB.n19 VNB 0.16fF
C66 VPB.n20 VNB 0.04fF
C67 VPB.n22 VNB 0.02fF
C68 VPB.n23 VNB 0.02fF
C69 VPB.n24 VNB 0.02fF
C70 VPB.n25 VNB 0.02fF
C71 VPB.n27 VNB 0.02fF
C72 VPB.n28 VNB 0.02fF
C73 VPB.n29 VNB 0.02fF
C74 VPB.n31 VNB 0.26fF
C75 VPB.n33 VNB 0.02fF
C76 VPB.n34 VNB 0.02fF
C77 VPB.n35 VNB 0.10fF
C78 VPB.n36 VNB 0.13fF
C79 VPB.n37 VNB 0.15fF
C80 VPB.n38 VNB 0.02fF
C81 VPB.n39 VNB 0.02fF
C82 VPB.n40 VNB 0.13fF
C83 VPB.n41 VNB 0.14fF
C84 VPB.n42 VNB 0.02fF
C85 VPB.n43 VNB 0.02fF
C86 VPB.n44 VNB 0.02fF
C87 VPB.n45 VNB 0.13fF
C88 VPB.n46 VNB 0.14fF
C89 VPB.n47 VNB 0.02fF
C90 VPB.n48 VNB 0.02fF
C91 VPB.n49 VNB 0.13fF
C92 VPB.n50 VNB 0.15fF
C93 VPB.n51 VNB 0.02fF
C94 VPB.n52 VNB 0.02fF
C95 VPB.n53 VNB 0.06fF
C96 VPB.n54 VNB 0.22fF
C97 VPB.n55 VNB 0.02fF
C98 VPB.n56 VNB 0.01fF
C99 VPB.n57 VNB 0.26fF
C100 VPB.n58 VNB 0.01fF
C101 VPB.n59 VNB 0.02fF
C102 VPB.n60 VNB 0.03fF
C103 VPB.n61 VNB 0.03fF
C104 VPB.n62 VNB 0.26fF
C105 VPB.n63 VNB 0.01fF
C106 VPB.n64 VNB 0.02fF
C107 VPB.n65 VNB 0.05fF
C108 VPB.n66 VNB 0.13fF
C109 VPB.n67 VNB 0.18fF
C110 VPB.n68 VNB 0.02fF
C111 VPB.n69 VNB 0.01fF
C112 VPB.n70 VNB 0.15fF
C113 VPB.n71 VNB 0.02fF
C114 VPB.n72 VNB 0.02fF
C115 VPB.n73 VNB 0.13fF
C116 VPB.n74 VNB 0.18fF
C117 VPB.n75 VNB 0.02fF
C118 VPB.n76 VNB 0.01fF
C119 VPB.n77 VNB 0.05fF
C120 VPB.n78 VNB 0.10fF
C121 VPB.n79 VNB 0.02fF
C122 VPB.n80 VNB 0.02fF
C123 VPB.n81 VNB 0.02fF
C124 VPB.n82 VNB 0.03fF
C125 VPB.n83 VNB 0.02fF
C126 VPB.n84 VNB 0.19fF
C127 VPB.n85 VNB 0.04fF
C128 VPB.n87 VNB 0.02fF
C129 VPB.n88 VNB 0.02fF
C130 VPB.n89 VNB 0.02fF
C131 VPB.n90 VNB 0.02fF
C132 VPB.n92 VNB 0.02fF
C133 VPB.n93 VNB 0.02fF
C134 VPB.n94 VNB 0.02fF
C135 VPB.n96 VNB 0.26fF
C136 VPB.n98 VNB 0.02fF
C137 VPB.n99 VNB 0.02fF
C138 VPB.n100 VNB 0.13fF
C139 VPB.n101 VNB 0.14fF
C140 VPB.n102 VNB 0.02fF
C141 VPB.n103 VNB 0.02fF
C142 VPB.n104 VNB 0.13fF
C143 VPB.n105 VNB 0.15fF
C144 VPB.n106 VNB 0.02fF
C145 VPB.n107 VNB 0.02fF
C146 VPB.n108 VNB 0.06fF
C147 VPB.n109 VNB 0.22fF
C148 VPB.n110 VNB 0.02fF
C149 VPB.n111 VNB 0.01fF
C150 VPB.n112 VNB 0.26fF
C151 VPB.n113 VNB 0.01fF
C152 VPB.n114 VNB 0.02fF
C153 VPB.n115 VNB 0.03fF
C154 VPB.n116 VNB 0.03fF
C155 VPB.n117 VNB 0.26fF
C156 VPB.n118 VNB 0.01fF
C157 VPB.n119 VNB 0.02fF
C158 VPB.n120 VNB 0.22fF
C159 VPB.n121 VNB 0.02fF
C160 VPB.n122 VNB 0.01fF
C161 VPB.n123 VNB 0.05fF
C162 VPB.n124 VNB 0.13fF
C163 VPB.n125 VNB 0.15fF
C164 VPB.n126 VNB 0.02fF
C165 VPB.n127 VNB 0.02fF
C166 VPB.n128 VNB 0.13fF
C167 VPB.n129 VNB 0.14fF
C168 VPB.n130 VNB 0.02fF
C169 VPB.n131 VNB 0.02fF
C170 VPB.n132 VNB 0.02fF
C171 VPB.n133 VNB 0.13fF
C172 VPB.n134 VNB 0.14fF
C173 VPB.n135 VNB 0.02fF
C174 VPB.n136 VNB 0.02fF
C175 VPB.n137 VNB 0.13fF
C176 VPB.n138 VNB 0.15fF
C177 VPB.n139 VNB 0.02fF
C178 VPB.n140 VNB 0.02fF
C179 VPB.n141 VNB 0.06fF
C180 VPB.n142 VNB 0.02fF
C181 VPB.n143 VNB 0.02fF
C182 VPB.n144 VNB 0.02fF
C183 VPB.n145 VNB 0.13fF
C184 VPB.n146 VNB 0.03fF
C185 VPB.n147 VNB 0.02fF
C186 VPB.n148 VNB 0.04fF
C187 VPB.n149 VNB 0.01fF
C188 VPB.n151 VNB 0.02fF
C189 VPB.n152 VNB 0.02fF
C190 VPB.n153 VNB 0.02fF
C191 VPB.n154 VNB 0.02fF
C192 VPB.n156 VNB 0.02fF
C193 VPB.n159 VNB 0.43fF
C194 VPB.n161 VNB 0.03fF
C195 VPB.n162 VNB 0.04fF
C196 VPB.n163 VNB 0.26fF
C197 VPB.n164 VNB 0.03fF
C198 VPB.n165 VNB 0.03fF
C199 VPB.n166 VNB 0.10fF
C200 VPB.n167 VNB 0.02fF
C201 VPB.n168 VNB 0.13fF
C202 VPB.n169 VNB 0.14fF
C203 VPB.n170 VNB 0.02fF
C204 VPB.n171 VNB 0.02fF
C205 VPB.n172 VNB 0.13fF
C206 VPB.n173 VNB 0.15fF
C207 VPB.n174 VNB 0.02fF
C208 VPB.n175 VNB 0.02fF
C209 VPB.n176 VNB 0.05fF
C210 VPB.n177 VNB 0.22fF
C211 VPB.n178 VNB 0.02fF
C212 VPB.n179 VNB 0.01fF
C213 VPB.n180 VNB 0.00fF
C214 VPB.n181 VNB 0.09fF
C215 VPB.n182 VNB 0.02fF
C216 VPB.n183 VNB 0.02fF
C217 VPB.n184 VNB 0.02fF
C218 VPB.n185 VNB 0.02fF
C219 VPB.n186 VNB 0.03fF
C220 VPB.n187 VNB 0.03fF
C221 VPB.n188 VNB 0.02fF
C222 VPB.n189 VNB 0.02fF
C223 VPB.n190 VNB 0.02fF
C224 VPB.n191 VNB 0.02fF
C225 VPB.n192 VNB 0.02fF
C226 VPB.n193 VNB 0.02fF
C227 VPB.n194 VNB 0.22fF
C228 VPB.n195 VNB 0.02fF
C229 VPB.n196 VNB 0.01fF
C230 VPB.n197 VNB 0.26fF
C231 VPB.n198 VNB 0.01fF
C232 VPB.n199 VNB 0.02fF
C233 VPB.n200 VNB 0.03fF
C234 VPB.n201 VNB 0.02fF
C235 VPB.n202 VNB 0.02fF
C236 VPB.n203 VNB 0.02fF
C237 VPB.n204 VNB 0.03fF
C238 VPB.n205 VNB 0.02fF
C239 VPB.n206 VNB 0.18fF
C240 VPB.n207 VNB 0.04fF
C241 VPB.n209 VNB 0.02fF
C242 VPB.n210 VNB 0.02fF
C243 VPB.n211 VNB 0.02fF
C244 VPB.n212 VNB 0.02fF
C245 VPB.n214 VNB 0.02fF
C246 VPB.n215 VNB 0.02fF
C247 VPB.n216 VNB 0.02fF
C248 VPB.n218 VNB 0.26fF
C249 VPB.n220 VNB 0.02fF
C250 VPB.n221 VNB 0.02fF
C251 VPB.n222 VNB 0.03fF
C252 VPB.n223 VNB 0.03fF
C253 VPB.n224 VNB 0.26fF
C254 VPB.n225 VNB 0.01fF
C255 VPB.n226 VNB 0.02fF
C256 VPB.n227 VNB 0.03fF
C257 VPB.n228 VNB 0.05fF
C258 VPB.n229 VNB 0.22fF
C259 VPB.n230 VNB 0.02fF
C260 VPB.n231 VNB 0.01fF
C261 VPB.n232 VNB 0.02fF
C262 VPB.n233 VNB 0.02fF
C263 VPB.n234 VNB 0.02fF
C264 VPB.n235 VNB 0.02fF
C265 VPB.n236 VNB 0.02fF
C266 VPB.n237 VNB 0.02fF
C267 VPB.n238 VNB 0.03fF
C268 VPB.n239 VNB 0.03fF
C269 VPB.n240 VNB 0.02fF
C270 VPB.n241 VNB 0.02fF
C271 VPB.n242 VNB 0.02fF
C272 VPB.n243 VNB 0.03fF
C273 VPB.n244 VNB 0.03fF
C274 VPB.n245 VNB 0.02fF
C275 VPB.n246 VNB 0.02fF
C276 VPB.n247 VNB 0.02fF
C277 VPB.n248 VNB 0.04fF
C278 VPB.n249 VNB 0.03fF
C279 VPB.n251 VNB 0.40fF
C280 a_661_1004.n0 VNB 0.53fF
C281 a_661_1004.n1 VNB 0.62fF
C282 a_661_1004.n2 VNB 0.35fF
C283 a_661_1004.n3 VNB 0.42fF
C284 a_661_1004.n4 VNB 0.82fF
C285 a_661_1004.n5 VNB 0.87fF
C286 a_661_1004.n6 VNB 0.08fF
C287 a_661_1004.n7 VNB 0.24fF
C288 a_661_1004.n8 VNB 0.05fF
C289 a_556_73.n0 VNB 0.05fF
C290 a_556_73.n1 VNB 0.02fF
C291 a_556_73.n2 VNB 0.12fF
C292 a_556_73.n3 VNB 0.04fF
C293 a_556_73.n4 VNB 0.17fF
.ends
