* SPICE3 file created from DFFQX1.ext - technology: sky130A

.subckt DFFQX1 Q D CLK VPB VNB
M1000 VPB.t18 a_147_159.t5 a_1845_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VPB.t15 a_147_159.t6 a_277_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPB.t25 a_1845_1004.t5 a_147_159.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_3177_1004.t4 a_277_1004.t7 VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VNB a_599_943.t5 a_1740_73.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1005 VPB.t10 CLK a_277_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPB.t9 CLK a_147_159.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_3177_1004.t2 Q VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VNB a_147_159.t13 a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPB.t12 a_599_943.t6 a_277_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t0 a_277_1004.t8 a_599_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_3177_1004.t6 VPB.t20 pshort w=2u l=0.15u
+  ad=1.16p pd=9.16u as=0p ps=0u
M1012 VNB a_3177_1004.t5 a_3738_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPB.t14 a_147_159.t7 Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1845_1004.t4 a_147_159.t8 VPB.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VNB a_277_1004.t9 a_1074_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1016 Q a_147_159.t9 VPB.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_277_1004.t4 a_147_159.t11 VPB.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPB.t1 a_1305_383# a_599_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPB.t6 a_599_943.t7 a_1845_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_277_1004.t1 CLK VPB.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 VNB a_277_1004.t10 a_3072_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_147_159.t2 CLK VPB.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPB.t22 a_277_1004.t11 a_3177_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 Q a_147_159.t12 a_3738_73.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1025 a_277_1004.t6 a_599_943.t8 VPB.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_599_943.t3 a_277_1004.t12 VPB.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_147_159.t0 a_1845_1004.t6 VPB.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPB.t4 Q a_3177_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPB.t23 a_3177_1004.t7 Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 VNB a_1845_1004.t7 a_2406_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_599_943.t1 a_1305_383# VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1845_1004.t0 a_599_943.t10 VPB.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VPB a_1305_383# 0.07fF
C1 VPB CLK 0.70fF
C2 VPB Q 1.44fF
C3 CLK a_1305_383# 0.04fF
R0 a_147_159.n8 a_147_159.t6 512.525
R1 a_147_159.n6 a_147_159.t5 472.359
R2 a_147_159.n4 a_147_159.t7 472.359
R3 a_147_159.n6 a_147_159.t8 384.527
R4 a_147_159.n4 a_147_159.t9 384.527
R5 a_147_159.n8 a_147_159.t11 371.139
R6 a_147_159.n9 a_147_159.t13 324.268
R7 a_147_159.n7 a_147_159.t10 277.772
R8 a_147_159.n5 a_147_159.t12 277.772
R9 a_147_159.n14 a_147_159.n12 247.192
R10 a_147_159.n9 a_147_159.n8 119.654
R11 a_147_159.n12 a_147_159.n3 109.441
R12 a_147_159.n10 a_147_159.n9 82.484
R13 a_147_159.n11 a_147_159.n5 80.307
R14 a_147_159.n3 a_147_159.n2 76.002
R15 a_147_159.n10 a_147_159.n7 76
R16 a_147_159.n12 a_147_159.n11 76
R17 a_147_159.n7 a_147_159.n6 67.001
R18 a_147_159.n5 a_147_159.n4 67.001
R19 a_147_159.n14 a_147_159.n13 30
R20 a_147_159.n15 a_147_159.n0 24.383
R21 a_147_159.n15 a_147_159.n14 23.684
R22 a_147_159.n1 a_147_159.t4 14.282
R23 a_147_159.n1 a_147_159.t2 14.282
R24 a_147_159.n2 a_147_159.t1 14.282
R25 a_147_159.n2 a_147_159.t0 14.282
R26 a_147_159.n3 a_147_159.n1 12.85
R27 a_147_159.n11 a_147_159.n10 2.947
R28 a_1845_1004.n4 a_1845_1004.t5 480.392
R29 a_1845_1004.n4 a_1845_1004.t6 403.272
R30 a_1845_1004.n5 a_1845_1004.t7 266.974
R31 a_1845_1004.n8 a_1845_1004.n6 194.086
R32 a_1845_1004.n6 a_1845_1004.n3 162.547
R33 a_1845_1004.n6 a_1845_1004.n5 153.315
R34 a_1845_1004.n5 a_1845_1004.n4 108.494
R35 a_1845_1004.n3 a_1845_1004.n2 76.002
R36 a_1845_1004.n8 a_1845_1004.n7 30
R37 a_1845_1004.n9 a_1845_1004.n0 24.383
R38 a_1845_1004.n9 a_1845_1004.n8 23.684
R39 a_1845_1004.n1 a_1845_1004.t2 14.282
R40 a_1845_1004.n1 a_1845_1004.t4 14.282
R41 a_1845_1004.n2 a_1845_1004.t1 14.282
R42 a_1845_1004.n2 a_1845_1004.t0 14.282
R43 a_1845_1004.n3 a_1845_1004.n1 12.85
R44 VPB VPB.n413 126.832
R45 VPB.n40 VPB.n38 94.117
R46 VPB.n355 VPB.n353 94.117
R47 VPB.n294 VPB.n292 94.117
R48 VPB.n132 VPB.n130 94.117
R49 VPB.n247 VPB.n245 94.117
R50 VPB.n50 VPB.n49 80.104
R51 VPB.n298 VPB.n82 76
R52 VPB.n208 VPB.n207 76
R53 VPB.n213 VPB.n212 76
R54 VPB.n218 VPB.n217 76
R55 VPB.n222 VPB.n221 76
R56 VPB.n249 VPB.n248 76
R57 VPB.n254 VPB.n253 76
R58 VPB.n259 VPB.n258 76
R59 VPB.n266 VPB.n265 76
R60 VPB.n271 VPB.n270 76
R61 VPB.n276 VPB.n275 76
R62 VPB.n281 VPB.n280 76
R63 VPB.n295 VPB.n291 76
R64 VPB.n304 VPB.n303 76
R65 VPB.n311 VPB.n310 76
R66 VPB.n316 VPB.n315 76
R67 VPB.n321 VPB.n320 76
R68 VPB.n326 VPB.n325 76
R69 VPB.n330 VPB.n329 76
R70 VPB.n357 VPB.n356 76
R71 VPB.n362 VPB.n361 76
R72 VPB.n367 VPB.n366 76
R73 VPB.n374 VPB.n373 76
R74 VPB.n379 VPB.n378 76
R75 VPB.n384 VPB.n383 76
R76 VPB.n389 VPB.n388 76
R77 VPB.n393 VPB.n392 76
R78 VPB.n406 VPB.n405 76
R79 VPB.n72 VPB.n71 75.654
R80 VPB.n22 VPB.n21 61.764
R81 VPB.n337 VPB.n336 61.764
R82 VPB.n89 VPB.n88 61.764
R83 VPB.n111 VPB.n110 61.764
R84 VPB.n229 VPB.n228 61.764
R85 VPB.n78 VPB.t16 55.106
R86 VPB.n385 VPB.t21 55.106
R87 VPB.n322 VPB.t5 55.106
R88 VPB.n155 VPB.t24 55.106
R89 VPB.n277 VPB.t11 55.106
R90 VPB.n214 VPB.t20 55.106
R91 VPB.n45 VPB.t12 55.106
R92 VPB.n358 VPB.t1 55.106
R93 VPB.n299 VPB.t18 55.106
R94 VPB.n137 VPB.t9 55.106
R95 VPB.n250 VPB.t4 55.106
R96 VPB.n197 VPB.t14 55.106
R97 VPB.n194 VPB.n193 48.952
R98 VPB.n256 VPB.n255 48.952
R99 VPB.n139 VPB.n138 48.952
R100 VPB.n301 VPB.n300 48.952
R101 VPB.n364 VPB.n363 48.952
R102 VPB.n54 VPB.n53 48.952
R103 VPB.n210 VPB.n209 44.502
R104 VPB.n273 VPB.n272 44.502
R105 VPB.n152 VPB.n151 44.502
R106 VPB.n318 VPB.n317 44.502
R107 VPB.n381 VPB.n380 44.502
R108 VPB.n68 VPB.n67 44.502
R109 VPB.n66 VPB.n14 40.824
R110 VPB.n57 VPB.n15 40.824
R111 VPB.n369 VPB.n368 40.824
R112 VPB.n306 VPB.n305 40.824
R113 VPB.n146 VPB.n104 40.824
R114 VPB.n261 VPB.n260 40.824
R115 VPB.n188 VPB.n187 40.824
R116 VPB.n202 VPB.n201 35.118
R117 VPB.n410 VPB.n406 20.452
R118 VPB.n186 VPB.n183 20.452
R119 VPB.n190 VPB.n189 17.801
R120 VPB.n263 VPB.n262 17.801
R121 VPB.n143 VPB.n142 17.801
R122 VPB.n308 VPB.n307 17.801
R123 VPB.n371 VPB.n370 17.801
R124 VPB.n59 VPB.n58 17.801
R125 VPB.n14 VPB.t7 14.282
R126 VPB.n14 VPB.t15 14.282
R127 VPB.n15 VPB.t19 14.282
R128 VPB.n15 VPB.t10 14.282
R129 VPB.n368 VPB.t2 14.282
R130 VPB.n368 VPB.t0 14.282
R131 VPB.n305 VPB.t17 14.282
R132 VPB.n305 VPB.t6 14.282
R133 VPB.n104 VPB.t8 14.282
R134 VPB.n104 VPB.t25 14.282
R135 VPB.n260 VPB.t3 14.282
R136 VPB.n260 VPB.t22 14.282
R137 VPB.n187 VPB.t13 14.282
R138 VPB.n187 VPB.t23 14.282
R139 VPB.n186 VPB.n185 13.653
R140 VPB.n185 VPB.n184 13.653
R141 VPB.n200 VPB.n199 13.653
R142 VPB.n199 VPB.n198 13.653
R143 VPB.n196 VPB.n195 13.653
R144 VPB.n195 VPB.n194 13.653
R145 VPB.n192 VPB.n191 13.653
R146 VPB.n191 VPB.n190 13.653
R147 VPB.n207 VPB.n206 13.653
R148 VPB.n206 VPB.n205 13.653
R149 VPB.n212 VPB.n211 13.653
R150 VPB.n211 VPB.n210 13.653
R151 VPB.n217 VPB.n216 13.653
R152 VPB.n216 VPB.n215 13.653
R153 VPB.n221 VPB.n220 13.653
R154 VPB.n220 VPB.n219 13.653
R155 VPB.n248 VPB.n247 13.653
R156 VPB.n247 VPB.n246 13.653
R157 VPB.n253 VPB.n252 13.653
R158 VPB.n252 VPB.n251 13.653
R159 VPB.n258 VPB.n257 13.653
R160 VPB.n257 VPB.n256 13.653
R161 VPB.n265 VPB.n264 13.653
R162 VPB.n264 VPB.n263 13.653
R163 VPB.n270 VPB.n269 13.653
R164 VPB.n269 VPB.n268 13.653
R165 VPB.n275 VPB.n274 13.653
R166 VPB.n274 VPB.n273 13.653
R167 VPB.n280 VPB.n279 13.653
R168 VPB.n279 VPB.n278 13.653
R169 VPB.n128 VPB.n127 13.653
R170 VPB.n127 VPB.n126 13.653
R171 VPB.n133 VPB.n132 13.653
R172 VPB.n132 VPB.n131 13.653
R173 VPB.n136 VPB.n135 13.653
R174 VPB.n135 VPB.n134 13.653
R175 VPB.n141 VPB.n140 13.653
R176 VPB.n140 VPB.n139 13.653
R177 VPB.n145 VPB.n144 13.653
R178 VPB.n144 VPB.n143 13.653
R179 VPB.n150 VPB.n149 13.653
R180 VPB.n149 VPB.n148 13.653
R181 VPB.n154 VPB.n153 13.653
R182 VPB.n153 VPB.n152 13.653
R183 VPB.n158 VPB.n157 13.653
R184 VPB.n157 VPB.n156 13.653
R185 VPB.n161 VPB.n160 13.653
R186 VPB.n160 VPB.n159 13.653
R187 VPB.n295 VPB.n294 13.653
R188 VPB.n294 VPB.n293 13.653
R189 VPB.n298 VPB.n297 13.653
R190 VPB.n297 VPB.n296 13.653
R191 VPB.n303 VPB.n302 13.653
R192 VPB.n302 VPB.n301 13.653
R193 VPB.n310 VPB.n309 13.653
R194 VPB.n309 VPB.n308 13.653
R195 VPB.n315 VPB.n314 13.653
R196 VPB.n314 VPB.n313 13.653
R197 VPB.n320 VPB.n319 13.653
R198 VPB.n319 VPB.n318 13.653
R199 VPB.n325 VPB.n324 13.653
R200 VPB.n324 VPB.n323 13.653
R201 VPB.n329 VPB.n328 13.653
R202 VPB.n328 VPB.n327 13.653
R203 VPB.n356 VPB.n355 13.653
R204 VPB.n355 VPB.n354 13.653
R205 VPB.n361 VPB.n360 13.653
R206 VPB.n360 VPB.n359 13.653
R207 VPB.n366 VPB.n365 13.653
R208 VPB.n365 VPB.n364 13.653
R209 VPB.n373 VPB.n372 13.653
R210 VPB.n372 VPB.n371 13.653
R211 VPB.n378 VPB.n377 13.653
R212 VPB.n377 VPB.n376 13.653
R213 VPB.n383 VPB.n382 13.653
R214 VPB.n382 VPB.n381 13.653
R215 VPB.n388 VPB.n387 13.653
R216 VPB.n387 VPB.n386 13.653
R217 VPB.n392 VPB.n391 13.653
R218 VPB.n391 VPB.n390 13.653
R219 VPB.n41 VPB.n40 13.653
R220 VPB.n40 VPB.n39 13.653
R221 VPB.n44 VPB.n43 13.653
R222 VPB.n43 VPB.n42 13.653
R223 VPB.n48 VPB.n47 13.653
R224 VPB.n47 VPB.n46 13.653
R225 VPB.n52 VPB.n51 13.653
R226 VPB.n51 VPB.n50 13.653
R227 VPB.n56 VPB.n55 13.653
R228 VPB.n55 VPB.n54 13.653
R229 VPB.n61 VPB.n60 13.653
R230 VPB.n60 VPB.n59 13.653
R231 VPB.n65 VPB.n64 13.653
R232 VPB.n64 VPB.n63 13.653
R233 VPB.n70 VPB.n69 13.653
R234 VPB.n69 VPB.n68 13.653
R235 VPB.n74 VPB.n73 13.653
R236 VPB.n73 VPB.n72 13.653
R237 VPB.n77 VPB.n76 13.653
R238 VPB.n76 VPB.n75 13.653
R239 VPB.n81 VPB.n80 13.653
R240 VPB.n80 VPB.n79 13.653
R241 VPB.n406 VPB.n0 13.653
R242 VPB VPB.n0 13.653
R243 VPB.n205 VPB.n204 13.35
R244 VPB.n268 VPB.n267 13.35
R245 VPB.n148 VPB.n147 13.35
R246 VPB.n313 VPB.n312 13.35
R247 VPB.n376 VPB.n375 13.35
R248 VPB.n63 VPB.n62 13.35
R249 VPB.n410 VPB.n409 13.276
R250 VPB.n409 VPB.n407 13.276
R251 VPB.n36 VPB.n18 13.276
R252 VPB.n18 VPB.n16 13.276
R253 VPB.n351 VPB.n333 13.276
R254 VPB.n333 VPB.n331 13.276
R255 VPB.n103 VPB.n85 13.276
R256 VPB.n85 VPB.n83 13.276
R257 VPB.n125 VPB.n107 13.276
R258 VPB.n107 VPB.n105 13.276
R259 VPB.n243 VPB.n225 13.276
R260 VPB.n225 VPB.n223 13.276
R261 VPB.n196 VPB.n192 13.276
R262 VPB.n248 VPB.n244 13.276
R263 VPB.n129 VPB.n128 13.276
R264 VPB.n133 VPB.n129 13.276
R265 VPB.n136 VPB.n133 13.276
R266 VPB.n145 VPB.n141 13.276
R267 VPB.n154 VPB.n150 13.276
R268 VPB.n161 VPB.n158 13.276
R269 VPB.n162 VPB.n161 13.276
R270 VPB.n295 VPB.n162 13.276
R271 VPB.n298 VPB.n295 13.276
R272 VPB.n356 VPB.n352 13.276
R273 VPB.n41 VPB.n37 13.276
R274 VPB.n44 VPB.n41 13.276
R275 VPB.n52 VPB.n48 13.276
R276 VPB.n56 VPB.n52 13.276
R277 VPB.n65 VPB.n61 13.276
R278 VPB.n74 VPB.n70 13.276
R279 VPB.n77 VPB.n74 13.276
R280 VPB.n406 VPB.n81 13.276
R281 VPB.n183 VPB.n165 13.276
R282 VPB.n165 VPB.n163 13.276
R283 VPB.n170 VPB.n168 12.796
R284 VPB.n170 VPB.n169 12.564
R285 VPB.n81 VPB.n78 12.558
R286 VPB.n45 VPB.n44 12.2
R287 VPB.n176 VPB.n175 12.198
R288 VPB.n178 VPB.n177 12.198
R289 VPB.n176 VPB.n173 12.198
R290 VPB.n197 VPB.n196 11.841
R291 VPB.n141 VPB.n137 11.841
R292 VPB.n303 VPB.n299 11.841
R293 VPB.n155 VPB.n154 11.482
R294 VPB.n61 VPB.n57 9.329
R295 VPB.n66 VPB.n65 8.97
R296 VPB.n183 VPB.n182 7.5
R297 VPB.n168 VPB.n167 7.5
R298 VPB.n175 VPB.n174 7.5
R299 VPB.n173 VPB.n172 7.5
R300 VPB.n165 VPB.n164 7.5
R301 VPB.n180 VPB.n166 7.5
R302 VPB.n225 VPB.n224 7.5
R303 VPB.n238 VPB.n237 7.5
R304 VPB.n232 VPB.n231 7.5
R305 VPB.n234 VPB.n233 7.5
R306 VPB.n227 VPB.n226 7.5
R307 VPB.n243 VPB.n242 7.5
R308 VPB.n107 VPB.n106 7.5
R309 VPB.n120 VPB.n119 7.5
R310 VPB.n114 VPB.n113 7.5
R311 VPB.n116 VPB.n115 7.5
R312 VPB.n109 VPB.n108 7.5
R313 VPB.n125 VPB.n124 7.5
R314 VPB.n85 VPB.n84 7.5
R315 VPB.n98 VPB.n97 7.5
R316 VPB.n92 VPB.n91 7.5
R317 VPB.n94 VPB.n93 7.5
R318 VPB.n87 VPB.n86 7.5
R319 VPB.n103 VPB.n102 7.5
R320 VPB.n333 VPB.n332 7.5
R321 VPB.n346 VPB.n345 7.5
R322 VPB.n340 VPB.n339 7.5
R323 VPB.n342 VPB.n341 7.5
R324 VPB.n335 VPB.n334 7.5
R325 VPB.n351 VPB.n350 7.5
R326 VPB.n18 VPB.n17 7.5
R327 VPB.n31 VPB.n30 7.5
R328 VPB.n25 VPB.n24 7.5
R329 VPB.n27 VPB.n26 7.5
R330 VPB.n20 VPB.n19 7.5
R331 VPB.n36 VPB.n35 7.5
R332 VPB.n409 VPB.n408 7.5
R333 VPB.n12 VPB.n11 7.5
R334 VPB.n6 VPB.n5 7.5
R335 VPB.n8 VPB.n7 7.5
R336 VPB.n2 VPB.n1 7.5
R337 VPB.n411 VPB.n410 7.5
R338 VPB.n37 VPB.n36 7.176
R339 VPB.n352 VPB.n351 7.176
R340 VPB.n162 VPB.n103 7.176
R341 VPB.n129 VPB.n125 7.176
R342 VPB.n244 VPB.n243 7.176
R343 VPB.n150 VPB.n146 6.817
R344 VPB.n239 VPB.n236 6.729
R345 VPB.n235 VPB.n232 6.729
R346 VPB.n230 VPB.n227 6.729
R347 VPB.n121 VPB.n118 6.729
R348 VPB.n117 VPB.n114 6.729
R349 VPB.n112 VPB.n109 6.729
R350 VPB.n99 VPB.n96 6.729
R351 VPB.n95 VPB.n92 6.729
R352 VPB.n90 VPB.n87 6.729
R353 VPB.n347 VPB.n344 6.729
R354 VPB.n343 VPB.n340 6.729
R355 VPB.n338 VPB.n335 6.729
R356 VPB.n32 VPB.n29 6.729
R357 VPB.n28 VPB.n25 6.729
R358 VPB.n23 VPB.n20 6.729
R359 VPB.n13 VPB.n10 6.729
R360 VPB.n9 VPB.n6 6.729
R361 VPB.n4 VPB.n2 6.729
R362 VPB.n230 VPB.n229 6.728
R363 VPB.n235 VPB.n234 6.728
R364 VPB.n239 VPB.n238 6.728
R365 VPB.n242 VPB.n241 6.728
R366 VPB.n112 VPB.n111 6.728
R367 VPB.n117 VPB.n116 6.728
R368 VPB.n121 VPB.n120 6.728
R369 VPB.n124 VPB.n123 6.728
R370 VPB.n90 VPB.n89 6.728
R371 VPB.n95 VPB.n94 6.728
R372 VPB.n99 VPB.n98 6.728
R373 VPB.n102 VPB.n101 6.728
R374 VPB.n338 VPB.n337 6.728
R375 VPB.n343 VPB.n342 6.728
R376 VPB.n347 VPB.n346 6.728
R377 VPB.n350 VPB.n349 6.728
R378 VPB.n23 VPB.n22 6.728
R379 VPB.n28 VPB.n27 6.728
R380 VPB.n32 VPB.n31 6.728
R381 VPB.n35 VPB.n34 6.728
R382 VPB.n4 VPB.n3 6.728
R383 VPB.n9 VPB.n8 6.728
R384 VPB.n13 VPB.n12 6.728
R385 VPB.n412 VPB.n411 6.728
R386 VPB.n192 VPB.n188 6.458
R387 VPB.n265 VPB.n261 6.458
R388 VPB.n146 VPB.n145 6.458
R389 VPB.n310 VPB.n306 6.458
R390 VPB.n373 VPB.n369 6.458
R391 VPB.n182 VPB.n181 6.398
R392 VPB.n201 VPB.n186 6.112
R393 VPB.n201 VPB.n200 6.101
R394 VPB.n70 VPB.n66 4.305
R395 VPB.n57 VPB.n56 3.947
R396 VPB.n217 VPB.n214 1.794
R397 VPB.n280 VPB.n277 1.794
R398 VPB.n158 VPB.n155 1.794
R399 VPB.n325 VPB.n322 1.794
R400 VPB.n388 VPB.n385 1.794
R401 VPB.n200 VPB.n197 1.435
R402 VPB.n253 VPB.n250 1.435
R403 VPB.n137 VPB.n136 1.435
R404 VPB.n299 VPB.n298 1.435
R405 VPB.n361 VPB.n358 1.435
R406 VPB.n180 VPB.n171 1.402
R407 VPB.n180 VPB.n176 1.402
R408 VPB.n180 VPB.n178 1.402
R409 VPB.n180 VPB.n179 1.402
R410 VPB.n48 VPB.n45 1.076
R411 VPB.n181 VPB.n180 0.735
R412 VPB.n180 VPB.n170 0.735
R413 VPB.n78 VPB.n77 0.717
R414 VPB.n240 VPB.n239 0.387
R415 VPB.n240 VPB.n235 0.387
R416 VPB.n240 VPB.n230 0.387
R417 VPB.n241 VPB.n240 0.387
R418 VPB.n122 VPB.n121 0.387
R419 VPB.n122 VPB.n117 0.387
R420 VPB.n122 VPB.n112 0.387
R421 VPB.n123 VPB.n122 0.387
R422 VPB.n100 VPB.n99 0.387
R423 VPB.n100 VPB.n95 0.387
R424 VPB.n100 VPB.n90 0.387
R425 VPB.n101 VPB.n100 0.387
R426 VPB.n348 VPB.n347 0.387
R427 VPB.n348 VPB.n343 0.387
R428 VPB.n348 VPB.n338 0.387
R429 VPB.n349 VPB.n348 0.387
R430 VPB.n33 VPB.n32 0.387
R431 VPB.n33 VPB.n28 0.387
R432 VPB.n33 VPB.n23 0.387
R433 VPB.n34 VPB.n33 0.387
R434 VPB.n413 VPB.n13 0.387
R435 VPB.n413 VPB.n9 0.387
R436 VPB.n413 VPB.n4 0.387
R437 VPB.n413 VPB.n412 0.387
R438 VPB.n249 VPB.n222 0.272
R439 VPB.n283 VPB.n282 0.272
R440 VPB.n291 VPB.n290 0.272
R441 VPB.n357 VPB.n330 0.272
R442 VPB.n394 VPB.n393 0.272
R443 VPB.n405 VPB 0.198
R444 VPB.n203 VPB.n202 0.136
R445 VPB.n208 VPB.n203 0.136
R446 VPB.n213 VPB.n208 0.136
R447 VPB.n218 VPB.n213 0.136
R448 VPB.n222 VPB.n218 0.136
R449 VPB.n254 VPB.n249 0.136
R450 VPB.n259 VPB.n254 0.136
R451 VPB.n266 VPB.n259 0.136
R452 VPB.n271 VPB.n266 0.136
R453 VPB.n276 VPB.n271 0.136
R454 VPB.n281 VPB.n276 0.136
R455 VPB.n282 VPB.n281 0.136
R456 VPB.n284 VPB.n283 0.136
R457 VPB.n285 VPB.n284 0.136
R458 VPB.n286 VPB.n285 0.136
R459 VPB.n287 VPB.n286 0.136
R460 VPB.n288 VPB.n287 0.136
R461 VPB.n289 VPB.n288 0.136
R462 VPB.n290 VPB.n289 0.136
R463 VPB.n291 VPB.n82 0.136
R464 VPB.n304 VPB.n82 0.136
R465 VPB.n311 VPB.n304 0.136
R466 VPB.n316 VPB.n311 0.136
R467 VPB.n321 VPB.n316 0.136
R468 VPB.n326 VPB.n321 0.136
R469 VPB.n330 VPB.n326 0.136
R470 VPB.n362 VPB.n357 0.136
R471 VPB.n367 VPB.n362 0.136
R472 VPB.n374 VPB.n367 0.136
R473 VPB.n379 VPB.n374 0.136
R474 VPB.n384 VPB.n379 0.136
R475 VPB.n389 VPB.n384 0.136
R476 VPB.n393 VPB.n389 0.136
R477 VPB.n395 VPB.n394 0.136
R478 VPB.n396 VPB.n395 0.136
R479 VPB.n397 VPB.n396 0.136
R480 VPB.n398 VPB.n397 0.136
R481 VPB.n399 VPB.n398 0.136
R482 VPB.n400 VPB.n399 0.136
R483 VPB.n401 VPB.n400 0.136
R484 VPB.n402 VPB.n401 0.136
R485 VPB.n403 VPB.n402 0.136
R486 VPB.n404 VPB.n403 0.136
R487 VPB.n405 VPB.n404 0.136
R488 a_277_1004.n8 a_277_1004.t8 480.392
R489 a_277_1004.n6 a_277_1004.t11 480.392
R490 a_277_1004.n8 a_277_1004.t12 403.272
R491 a_277_1004.n6 a_277_1004.t7 403.272
R492 a_277_1004.n9 a_277_1004.t9 293.527
R493 a_277_1004.n7 a_277_1004.t10 293.527
R494 a_277_1004.n13 a_277_1004.n11 223.151
R495 a_277_1004.n11 a_277_1004.n5 154.293
R496 a_277_1004.n10 a_277_1004.n7 83.3
R497 a_277_1004.n9 a_277_1004.n8 81.941
R498 a_277_1004.n7 a_277_1004.n6 81.941
R499 a_277_1004.n4 a_277_1004.n3 79.232
R500 a_277_1004.n11 a_277_1004.n10 77.315
R501 a_277_1004.n10 a_277_1004.n9 76
R502 a_277_1004.n5 a_277_1004.n4 63.152
R503 a_277_1004.n13 a_277_1004.n12 30
R504 a_277_1004.n14 a_277_1004.n0 24.383
R505 a_277_1004.n14 a_277_1004.n13 23.684
R506 a_277_1004.n5 a_277_1004.n1 16.08
R507 a_277_1004.n4 a_277_1004.n2 16.08
R508 a_277_1004.n1 a_277_1004.t3 14.282
R509 a_277_1004.n1 a_277_1004.t6 14.282
R510 a_277_1004.n2 a_277_1004.t2 14.282
R511 a_277_1004.n2 a_277_1004.t1 14.282
R512 a_277_1004.n3 a_277_1004.t5 14.282
R513 a_277_1004.n3 a_277_1004.t4 14.282
R514 a_3177_1004.n4 a_3177_1004.t7 480.392
R515 a_3177_1004.n4 a_3177_1004.t6 403.272
R516 a_3177_1004.n5 a_3177_1004.t5 266.974
R517 a_3177_1004.n8 a_3177_1004.n6 194.086
R518 a_3177_1004.n6 a_3177_1004.n3 162.547
R519 a_3177_1004.n6 a_3177_1004.n5 153.315
R520 a_3177_1004.n5 a_3177_1004.n4 108.494
R521 a_3177_1004.n3 a_3177_1004.n2 76.002
R522 a_3177_1004.n8 a_3177_1004.n7 30
R523 a_3177_1004.n9 a_3177_1004.n0 24.383
R524 a_3177_1004.n9 a_3177_1004.n8 23.684
R525 a_3177_1004.n1 a_3177_1004.t1 14.282
R526 a_3177_1004.n1 a_3177_1004.t2 14.282
R527 a_3177_1004.n2 a_3177_1004.t3 14.282
R528 a_3177_1004.n2 a_3177_1004.t4 14.282
R529 a_3177_1004.n3 a_3177_1004.n1 12.85
R530 a_91_75.t0 a_91_75.n0 117.777
R531 a_91_75.n2 a_91_75.n1 55.228
R532 a_91_75.n4 a_91_75.n3 9.111
R533 a_91_75.n8 a_91_75.n6 7.859
R534 a_91_75.t0 a_91_75.n2 4.04
R535 a_91_75.t0 a_91_75.n8 3.034
R536 a_91_75.n6 a_91_75.n4 1.964
R537 a_91_75.n6 a_91_75.n5 1.964
R538 a_91_75.n8 a_91_75.n7 0.443
R539 a_372_182.n8 a_372_182.n6 96.467
R540 a_372_182.n3 a_372_182.n1 44.628
R541 a_372_182.t0 a_372_182.n8 32.417
R542 a_372_182.n3 a_372_182.n2 23.284
R543 a_372_182.n6 a_372_182.n5 22.349
R544 a_372_182.t0 a_372_182.n10 20.241
R545 a_372_182.n10 a_372_182.n9 13.494
R546 a_372_182.n6 a_372_182.n4 8.443
R547 a_372_182.t0 a_372_182.n0 8.137
R548 a_372_182.t0 a_372_182.n3 5.727
R549 a_372_182.n8 a_372_182.n7 1.435
R550 a_599_943.n4 a_599_943.t7 480.392
R551 a_599_943.n6 a_599_943.t8 454.685
R552 a_599_943.n6 a_599_943.t6 428.979
R553 a_599_943.n4 a_599_943.t10 403.272
R554 a_599_943.n5 a_599_943.t5 266.974
R555 a_599_943.n7 a_599_943.t9 221.453
R556 a_599_943.n11 a_599_943.n9 194.086
R557 a_599_943.n9 a_599_943.n3 162.547
R558 a_599_943.n7 a_599_943.n6 108.494
R559 a_599_943.n5 a_599_943.n4 108.494
R560 a_599_943.n8 a_599_943.n7 78.947
R561 a_599_943.n8 a_599_943.n5 77.315
R562 a_599_943.n3 a_599_943.n2 76.002
R563 a_599_943.n9 a_599_943.n8 76
R564 a_599_943.n11 a_599_943.n10 30
R565 a_599_943.n12 a_599_943.n0 24.383
R566 a_599_943.n12 a_599_943.n11 23.684
R567 a_599_943.n1 a_599_943.t2 14.282
R568 a_599_943.n1 a_599_943.t1 14.282
R569 a_599_943.n2 a_599_943.t4 14.282
R570 a_599_943.n2 a_599_943.t3 14.282
R571 a_599_943.n3 a_599_943.n1 12.85
R572 a_1740_73.t0 a_1740_73.n1 93.333
R573 a_1740_73.n4 a_1740_73.n2 55.07
R574 a_1740_73.t0 a_1740_73.n0 8.137
R575 a_1740_73.n4 a_1740_73.n3 4.619
R576 a_1740_73.t0 a_1740_73.n4 0.071
R577 VNB VNB.n366 300.778
R578 VNB.n194 VNB.n193 199.897
R579 VNB.n88 VNB.n87 199.897
R580 VNB.n68 VNB.n67 199.897
R581 VNB.n292 VNB.n291 199.897
R582 VNB.n15 VNB.n14 199.897
R583 VNB.n100 VNB.n98 154.509
R584 VNB.n203 VNB.n201 154.509
R585 VNB.n301 VNB.n299 154.509
R586 VNB.n251 VNB.n249 154.509
R587 VNB.n24 VNB.n22 154.509
R588 VNB.n160 VNB.n159 121.366
R589 VNB.n219 VNB.n218 121.366
R590 VNB.n112 VNB.n111 121.366
R591 VNB.n317 VNB.n316 121.366
R592 VNB.n53 VNB.n4 85.559
R593 VNB.n269 VNB.n268 84.842
R594 VNB.n255 VNB.n57 76
R595 VNB.n353 VNB.n352 76
R596 VNB.n340 VNB.n339 76
R597 VNB.n336 VNB.n335 76
R598 VNB.n332 VNB.n331 76
R599 VNB.n321 VNB.n320 76
R600 VNB.n315 VNB.n314 76
R601 VNB.n311 VNB.n310 76
R602 VNB.n307 VNB.n306 76
R603 VNB.n303 VNB.n302 76
R604 VNB.n281 VNB.n280 76
R605 VNB.n277 VNB.n276 76
R606 VNB.n273 VNB.n272 76
R607 VNB.n267 VNB.n266 76
R608 VNB.n263 VNB.n262 76
R609 VNB.n259 VNB.n258 76
R610 VNB.n252 VNB.n248 76
R611 VNB.n238 VNB.n237 76
R612 VNB.n234 VNB.n233 76
R613 VNB.n223 VNB.n222 76
R614 VNB.n217 VNB.n216 76
R615 VNB.n213 VNB.n212 76
R616 VNB.n209 VNB.n208 76
R617 VNB.n205 VNB.n204 76
R618 VNB.n183 VNB.n182 76
R619 VNB.n179 VNB.n178 76
R620 VNB.n175 VNB.n174 76
R621 VNB.n164 VNB.n163 76
R622 VNB.n169 VNB.n168 63.835
R623 VNB.n228 VNB.n227 63.835
R624 VNB.n116 VNB.n77 63.835
R625 VNB.n326 VNB.n325 63.835
R626 VNB.n51 VNB.n50 41.971
R627 VNB.n161 VNB.n160 36.937
R628 VNB.n220 VNB.n219 36.937
R629 VNB.n113 VNB.n112 36.937
R630 VNB.n318 VNB.n317 36.937
R631 VNB.n271 VNB.n270 36.678
R632 VNB.n157 VNB.n156 35.118
R633 VNB.n168 VNB.n167 28.421
R634 VNB.n227 VNB.n226 28.421
R635 VNB.n77 VNB.n76 28.421
R636 VNB.n325 VNB.n324 28.421
R637 VNB.n172 VNB.n171 27.855
R638 VNB.n231 VNB.n230 27.855
R639 VNB.n119 VNB.n118 27.855
R640 VNB.n329 VNB.n328 27.855
R641 VNB.n168 VNB.n166 25.263
R642 VNB.n227 VNB.n225 25.263
R643 VNB.n77 VNB.n75 25.263
R644 VNB.n325 VNB.n323 25.263
R645 VNB.n166 VNB.n165 24.383
R646 VNB.n225 VNB.n224 24.383
R647 VNB.n75 VNB.n74 24.383
R648 VNB.n323 VNB.n322 24.383
R649 VNB.n146 VNB.n143 20.452
R650 VNB.n354 VNB.n353 20.452
R651 VNB.n173 VNB.n172 16.721
R652 VNB.n232 VNB.n231 16.721
R653 VNB.n120 VNB.n119 16.721
R654 VNB.n330 VNB.n329 16.721
R655 VNB.n155 VNB.n154 13.653
R656 VNB.n154 VNB.n153 13.653
R657 VNB.n152 VNB.n151 13.653
R658 VNB.n151 VNB.n150 13.653
R659 VNB.n149 VNB.n148 13.653
R660 VNB.n148 VNB.n147 13.653
R661 VNB.n163 VNB.n162 13.653
R662 VNB.n162 VNB.n161 13.653
R663 VNB.n174 VNB.n173 13.653
R664 VNB.n178 VNB.n177 13.653
R665 VNB.n177 VNB.n176 13.653
R666 VNB.n182 VNB.n181 13.653
R667 VNB.n181 VNB.n180 13.653
R668 VNB.n204 VNB.n203 13.653
R669 VNB.n203 VNB.n202 13.653
R670 VNB.n208 VNB.n207 13.653
R671 VNB.n207 VNB.n206 13.653
R672 VNB.n212 VNB.n211 13.653
R673 VNB.n211 VNB.n210 13.653
R674 VNB.n216 VNB.n215 13.653
R675 VNB.n215 VNB.n214 13.653
R676 VNB.n222 VNB.n221 13.653
R677 VNB.n221 VNB.n220 13.653
R678 VNB.n233 VNB.n232 13.653
R679 VNB.n237 VNB.n236 13.653
R680 VNB.n236 VNB.n235 13.653
R681 VNB.n96 VNB.n95 13.653
R682 VNB.n95 VNB.n94 13.653
R683 VNB.n101 VNB.n100 13.653
R684 VNB.n100 VNB.n99 13.653
R685 VNB.n104 VNB.n103 13.653
R686 VNB.n103 VNB.n102 13.653
R687 VNB.n107 VNB.n106 13.653
R688 VNB.n106 VNB.n105 13.653
R689 VNB.n110 VNB.n109 13.653
R690 VNB.n109 VNB.n108 13.653
R691 VNB.n115 VNB.n114 13.653
R692 VNB.n114 VNB.n113 13.653
R693 VNB.n121 VNB.n120 13.653
R694 VNB.n124 VNB.n123 13.653
R695 VNB.n123 VNB.n122 13.653
R696 VNB.n127 VNB.n126 13.653
R697 VNB.n126 VNB.n125 13.653
R698 VNB.n252 VNB.n251 13.653
R699 VNB.n251 VNB.n250 13.653
R700 VNB.n255 VNB.n254 13.653
R701 VNB.n254 VNB.n253 13.653
R702 VNB.n258 VNB.n257 13.653
R703 VNB.n257 VNB.n256 13.653
R704 VNB.n262 VNB.n261 13.653
R705 VNB.n261 VNB.n260 13.653
R706 VNB.n266 VNB.n265 13.653
R707 VNB.n265 VNB.n264 13.653
R708 VNB.n272 VNB.n271 13.653
R709 VNB.n276 VNB.n275 13.653
R710 VNB.n275 VNB.n274 13.653
R711 VNB.n280 VNB.n279 13.653
R712 VNB.n279 VNB.n278 13.653
R713 VNB.n302 VNB.n301 13.653
R714 VNB.n301 VNB.n300 13.653
R715 VNB.n306 VNB.n305 13.653
R716 VNB.n305 VNB.n304 13.653
R717 VNB.n310 VNB.n309 13.653
R718 VNB.n309 VNB.n308 13.653
R719 VNB.n314 VNB.n313 13.653
R720 VNB.n313 VNB.n312 13.653
R721 VNB.n320 VNB.n319 13.653
R722 VNB.n319 VNB.n318 13.653
R723 VNB.n331 VNB.n330 13.653
R724 VNB.n335 VNB.n334 13.653
R725 VNB.n334 VNB.n333 13.653
R726 VNB.n339 VNB.n338 13.653
R727 VNB.n338 VNB.n337 13.653
R728 VNB.n25 VNB.n24 13.653
R729 VNB.n24 VNB.n23 13.653
R730 VNB.n28 VNB.n27 13.653
R731 VNB.n27 VNB.n26 13.653
R732 VNB.n31 VNB.n30 13.653
R733 VNB.n30 VNB.n29 13.653
R734 VNB.n34 VNB.n33 13.653
R735 VNB.n33 VNB.n32 13.653
R736 VNB.n37 VNB.n36 13.653
R737 VNB.n36 VNB.n35 13.653
R738 VNB.n40 VNB.n39 13.653
R739 VNB.n39 VNB.n38 13.653
R740 VNB.n43 VNB.n42 13.653
R741 VNB.n42 VNB.n41 13.653
R742 VNB.n46 VNB.n45 13.653
R743 VNB.n45 VNB.n44 13.653
R744 VNB.n49 VNB.n48 13.653
R745 VNB.n48 VNB.n47 13.653
R746 VNB.n52 VNB.n51 13.653
R747 VNB.n56 VNB.n55 13.653
R748 VNB.n55 VNB.n54 13.653
R749 VNB.n353 VNB.n0 13.653
R750 VNB VNB.n0 13.653
R751 VNB.n146 VNB.n145 13.653
R752 VNB.n145 VNB.n144 13.653
R753 VNB.n361 VNB.n358 13.577
R754 VNB.n131 VNB.n129 13.276
R755 VNB.n143 VNB.n131 13.276
R756 VNB.n186 VNB.n184 13.276
R757 VNB.n199 VNB.n186 13.276
R758 VNB.n80 VNB.n78 13.276
R759 VNB.n93 VNB.n80 13.276
R760 VNB.n60 VNB.n58 13.276
R761 VNB.n73 VNB.n60 13.276
R762 VNB.n284 VNB.n282 13.276
R763 VNB.n297 VNB.n284 13.276
R764 VNB.n7 VNB.n5 13.276
R765 VNB.n20 VNB.n7 13.276
R766 VNB.n155 VNB.n152 13.276
R767 VNB.n152 VNB.n149 13.276
R768 VNB.n204 VNB.n200 13.276
R769 VNB.n97 VNB.n96 13.276
R770 VNB.n101 VNB.n97 13.276
R771 VNB.n104 VNB.n101 13.276
R772 VNB.n107 VNB.n104 13.276
R773 VNB.n110 VNB.n107 13.276
R774 VNB.n115 VNB.n110 13.276
R775 VNB.n124 VNB.n121 13.276
R776 VNB.n127 VNB.n124 13.276
R777 VNB.n128 VNB.n127 13.276
R778 VNB.n252 VNB.n128 13.276
R779 VNB.n255 VNB.n252 13.276
R780 VNB.n258 VNB.n255 13.276
R781 VNB.n302 VNB.n298 13.276
R782 VNB.n25 VNB.n21 13.276
R783 VNB.n28 VNB.n25 13.276
R784 VNB.n31 VNB.n28 13.276
R785 VNB.n34 VNB.n31 13.276
R786 VNB.n37 VNB.n34 13.276
R787 VNB.n40 VNB.n37 13.276
R788 VNB.n43 VNB.n40 13.276
R789 VNB.n46 VNB.n43 13.276
R790 VNB.n49 VNB.n46 13.276
R791 VNB.n52 VNB.n49 13.276
R792 VNB.n353 VNB.n56 13.276
R793 VNB.n3 VNB.n1 13.276
R794 VNB.n354 VNB.n3 13.276
R795 VNB.n56 VNB.n53 12.02
R796 VNB.n116 VNB.n115 10.764
R797 VNB.n363 VNB.n362 7.5
R798 VNB.n192 VNB.n191 7.5
R799 VNB.n188 VNB.n187 7.5
R800 VNB.n186 VNB.n185 7.5
R801 VNB.n199 VNB.n198 7.5
R802 VNB.n86 VNB.n85 7.5
R803 VNB.n82 VNB.n81 7.5
R804 VNB.n80 VNB.n79 7.5
R805 VNB.n93 VNB.n92 7.5
R806 VNB.n66 VNB.n65 7.5
R807 VNB.n62 VNB.n61 7.5
R808 VNB.n60 VNB.n59 7.5
R809 VNB.n73 VNB.n72 7.5
R810 VNB.n290 VNB.n289 7.5
R811 VNB.n286 VNB.n285 7.5
R812 VNB.n284 VNB.n283 7.5
R813 VNB.n297 VNB.n296 7.5
R814 VNB.n13 VNB.n12 7.5
R815 VNB.n9 VNB.n8 7.5
R816 VNB.n7 VNB.n6 7.5
R817 VNB.n20 VNB.n19 7.5
R818 VNB.n355 VNB.n354 7.5
R819 VNB.n3 VNB.n2 7.5
R820 VNB.n360 VNB.n359 7.5
R821 VNB.n137 VNB.n136 7.5
R822 VNB.n133 VNB.n132 7.5
R823 VNB.n131 VNB.n130 7.5
R824 VNB.n143 VNB.n142 7.5
R825 VNB.n200 VNB.n199 7.176
R826 VNB.n97 VNB.n93 7.176
R827 VNB.n128 VNB.n73 7.176
R828 VNB.n298 VNB.n297 7.176
R829 VNB.n21 VNB.n20 7.176
R830 VNB.n365 VNB.n363 7.011
R831 VNB.n195 VNB.n192 7.011
R832 VNB.n190 VNB.n188 7.011
R833 VNB.n89 VNB.n86 7.011
R834 VNB.n84 VNB.n82 7.011
R835 VNB.n69 VNB.n66 7.011
R836 VNB.n64 VNB.n62 7.011
R837 VNB.n293 VNB.n290 7.011
R838 VNB.n288 VNB.n286 7.011
R839 VNB.n16 VNB.n13 7.011
R840 VNB.n11 VNB.n9 7.011
R841 VNB.n139 VNB.n137 7.011
R842 VNB.n135 VNB.n133 7.011
R843 VNB.n198 VNB.n197 7.01
R844 VNB.n190 VNB.n189 7.01
R845 VNB.n195 VNB.n194 7.01
R846 VNB.n92 VNB.n91 7.01
R847 VNB.n84 VNB.n83 7.01
R848 VNB.n89 VNB.n88 7.01
R849 VNB.n72 VNB.n71 7.01
R850 VNB.n64 VNB.n63 7.01
R851 VNB.n69 VNB.n68 7.01
R852 VNB.n296 VNB.n295 7.01
R853 VNB.n288 VNB.n287 7.01
R854 VNB.n293 VNB.n292 7.01
R855 VNB.n19 VNB.n18 7.01
R856 VNB.n11 VNB.n10 7.01
R857 VNB.n16 VNB.n15 7.01
R858 VNB.n142 VNB.n141 7.01
R859 VNB.n135 VNB.n134 7.01
R860 VNB.n139 VNB.n138 7.01
R861 VNB.n365 VNB.n364 7.01
R862 VNB.n361 VNB.n360 6.788
R863 VNB.n356 VNB.n355 6.788
R864 VNB.n156 VNB.n146 6.111
R865 VNB.n156 VNB.n155 6.1
R866 VNB.n174 VNB.n169 2.511
R867 VNB.n233 VNB.n228 2.511
R868 VNB.n121 VNB.n116 2.511
R869 VNB.n272 VNB.n269 2.511
R870 VNB.n331 VNB.n326 2.511
R871 VNB.n172 VNB.n170 1.99
R872 VNB.n231 VNB.n229 1.99
R873 VNB.n119 VNB.n117 1.99
R874 VNB.n329 VNB.n327 1.99
R875 VNB.n53 VNB.n52 1.255
R876 VNB.n366 VNB.n357 0.921
R877 VNB.n366 VNB.n361 0.476
R878 VNB.n366 VNB.n356 0.475
R879 VNB.n205 VNB.n183 0.272
R880 VNB.n240 VNB.n239 0.272
R881 VNB.n248 VNB.n247 0.272
R882 VNB.n303 VNB.n281 0.272
R883 VNB.n341 VNB.n340 0.272
R884 VNB.n196 VNB.n190 0.246
R885 VNB.n197 VNB.n196 0.246
R886 VNB.n196 VNB.n195 0.246
R887 VNB.n90 VNB.n84 0.246
R888 VNB.n91 VNB.n90 0.246
R889 VNB.n90 VNB.n89 0.246
R890 VNB.n70 VNB.n64 0.246
R891 VNB.n71 VNB.n70 0.246
R892 VNB.n70 VNB.n69 0.246
R893 VNB.n294 VNB.n288 0.246
R894 VNB.n295 VNB.n294 0.246
R895 VNB.n294 VNB.n293 0.246
R896 VNB.n17 VNB.n11 0.246
R897 VNB.n18 VNB.n17 0.246
R898 VNB.n17 VNB.n16 0.246
R899 VNB.n140 VNB.n135 0.246
R900 VNB.n141 VNB.n140 0.246
R901 VNB.n140 VNB.n139 0.246
R902 VNB.n366 VNB.n365 0.246
R903 VNB.n352 VNB 0.198
R904 VNB.n158 VNB.n157 0.136
R905 VNB.n164 VNB.n158 0.136
R906 VNB.n175 VNB.n164 0.136
R907 VNB.n179 VNB.n175 0.136
R908 VNB.n183 VNB.n179 0.136
R909 VNB.n209 VNB.n205 0.136
R910 VNB.n213 VNB.n209 0.136
R911 VNB.n217 VNB.n213 0.136
R912 VNB.n223 VNB.n217 0.136
R913 VNB.n234 VNB.n223 0.136
R914 VNB.n238 VNB.n234 0.136
R915 VNB.n239 VNB.n238 0.136
R916 VNB.n241 VNB.n240 0.136
R917 VNB.n242 VNB.n241 0.136
R918 VNB.n243 VNB.n242 0.136
R919 VNB.n244 VNB.n243 0.136
R920 VNB.n245 VNB.n244 0.136
R921 VNB.n246 VNB.n245 0.136
R922 VNB.n247 VNB.n246 0.136
R923 VNB.n248 VNB.n57 0.136
R924 VNB.n259 VNB.n57 0.136
R925 VNB.n263 VNB.n259 0.136
R926 VNB.n267 VNB.n263 0.136
R927 VNB.n273 VNB.n267 0.136
R928 VNB.n277 VNB.n273 0.136
R929 VNB.n281 VNB.n277 0.136
R930 VNB.n307 VNB.n303 0.136
R931 VNB.n311 VNB.n307 0.136
R932 VNB.n315 VNB.n311 0.136
R933 VNB.n321 VNB.n315 0.136
R934 VNB.n332 VNB.n321 0.136
R935 VNB.n336 VNB.n332 0.136
R936 VNB.n340 VNB.n336 0.136
R937 VNB.n342 VNB.n341 0.136
R938 VNB.n343 VNB.n342 0.136
R939 VNB.n344 VNB.n343 0.136
R940 VNB.n345 VNB.n344 0.136
R941 VNB.n346 VNB.n345 0.136
R942 VNB.n347 VNB.n346 0.136
R943 VNB.n348 VNB.n347 0.136
R944 VNB.n349 VNB.n348 0.136
R945 VNB.n350 VNB.n349 0.136
R946 VNB.n351 VNB.n350 0.136
R947 VNB.n352 VNB.n351 0.136
R948 a_2406_73.t0 a_2406_73.n1 34.62
R949 a_2406_73.t0 a_2406_73.n0 8.137
R950 a_2406_73.t0 a_2406_73.n2 4.69
R951 a_3738_73.n12 a_3738_73.n11 26.811
R952 a_3738_73.n6 a_3738_73.n5 24.977
R953 a_3738_73.n2 a_3738_73.n1 24.877
R954 a_3738_73.t0 a_3738_73.n2 12.677
R955 a_3738_73.t0 a_3738_73.n3 11.595
R956 a_3738_73.t1 a_3738_73.n8 8.137
R957 a_3738_73.t0 a_3738_73.n4 7.273
R958 a_3738_73.t0 a_3738_73.n0 6.109
R959 a_3738_73.t1 a_3738_73.n7 4.864
R960 a_3738_73.t0 a_3738_73.n12 2.074
R961 a_3738_73.n7 a_3738_73.n6 1.13
R962 a_3738_73.n12 a_3738_73.t1 0.937
R963 a_3738_73.t1 a_3738_73.n10 0.804
R964 a_3738_73.n10 a_3738_73.n9 0.136
R965 a_1074_73.t0 a_1074_73.n1 34.62
R966 a_1074_73.t0 a_1074_73.n0 8.137
R967 a_1074_73.t0 a_1074_73.n2 4.69
R968 a_3072_73.t0 a_3072_73.n1 34.62
R969 a_3072_73.t0 a_3072_73.n0 8.137
R970 a_3072_73.t0 a_3072_73.n2 4.69
C4 VPB VNB 17.10fF
C5 a_3072_73.n0 VNB 0.05fF
C6 a_3072_73.n1 VNB 0.12fF
C7 a_3072_73.n2 VNB 0.04fF
C8 a_1074_73.n0 VNB 0.05fF
C9 a_1074_73.n1 VNB 0.12fF
C10 a_1074_73.n2 VNB 0.04fF
C11 a_3738_73.n0 VNB 0.02fF
C12 a_3738_73.n1 VNB 0.10fF
C13 a_3738_73.n2 VNB 0.06fF
C14 a_3738_73.n3 VNB 0.06fF
C15 a_3738_73.n4 VNB 0.00fF
C16 a_3738_73.n5 VNB 0.04fF
C17 a_3738_73.n6 VNB 0.05fF
C18 a_3738_73.n7 VNB 0.02fF
C19 a_3738_73.n8 VNB 0.05fF
C20 a_3738_73.n9 VNB 0.07fF
C21 a_3738_73.n10 VNB 0.17fF
C22 a_3738_73.n11 VNB 0.09fF
C23 a_3738_73.n12 VNB 0.00fF
C24 a_2406_73.n0 VNB 0.05fF
C25 a_2406_73.n1 VNB 0.12fF
C26 a_2406_73.n2 VNB 0.04fF
C27 a_1740_73.n0 VNB 0.05fF
C28 a_1740_73.n1 VNB 0.02fF
C29 a_1740_73.n2 VNB 0.12fF
C30 a_1740_73.n3 VNB 0.04fF
C31 a_1740_73.n4 VNB 0.17fF
C32 a_599_943.n0 VNB 0.04fF
C33 a_599_943.n1 VNB 0.56fF
C34 a_599_943.n2 VNB 0.66fF
C35 a_599_943.n3 VNB 0.33fF
C36 a_599_943.n4 VNB 0.41fF
C37 a_599_943.n5 VNB 0.41fF
C38 a_599_943.n6 VNB 0.41fF
C39 a_599_943.t9 VNB 0.54fF
C40 a_599_943.n7 VNB 0.39fF
C41 a_599_943.n8 VNB 1.07fF
C42 a_599_943.n9 VNB 0.44fF
C43 a_599_943.n10 VNB 0.04fF
C44 a_599_943.n11 VNB 0.29fF
C45 a_599_943.n12 VNB 0.06fF
C46 a_372_182.n0 VNB 0.07fF
C47 a_372_182.n1 VNB 0.09fF
C48 a_372_182.n2 VNB 0.13fF
C49 a_372_182.n3 VNB 0.11fF
C50 a_372_182.n4 VNB 0.02fF
C51 a_372_182.n5 VNB 0.03fF
C52 a_372_182.n6 VNB 0.06fF
C53 a_372_182.n7 VNB 0.03fF
C54 a_372_182.n8 VNB 0.12fF
C55 a_372_182.n9 VNB 0.06fF
C56 a_372_182.n10 VNB 0.01fF
C57 a_372_182.t0 VNB 0.33fF
C58 a_91_75.n0 VNB 0.03fF
C59 a_91_75.n1 VNB 0.10fF
C60 a_91_75.n2 VNB 0.10fF
C61 a_91_75.n3 VNB 0.04fF
C62 a_91_75.n4 VNB 0.03fF
C63 a_91_75.n5 VNB 0.03fF
C64 a_91_75.n6 VNB 0.11fF
C65 a_91_75.n7 VNB 0.04fF
C66 a_3177_1004.n0 VNB 0.04fF
C67 a_3177_1004.n1 VNB 0.51fF
C68 a_3177_1004.n2 VNB 0.60fF
C69 a_3177_1004.n3 VNB 0.30fF
C70 a_3177_1004.n4 VNB 0.37fF
C71 a_3177_1004.n5 VNB 0.54fF
C72 a_3177_1004.n6 VNB 0.57fF
C73 a_3177_1004.n7 VNB 0.03fF
C74 a_3177_1004.n8 VNB 0.27fF
C75 a_3177_1004.n9 VNB 0.05fF
C76 a_277_1004.n0 VNB 0.05fF
C77 a_277_1004.n1 VNB 0.69fF
C78 a_277_1004.n2 VNB 0.69fF
C79 a_277_1004.n3 VNB 0.82fF
C80 a_277_1004.n4 VNB 0.26fF
C81 a_277_1004.n5 VNB 0.37fF
C82 a_277_1004.n6 VNB 0.46fF
C83 a_277_1004.n7 VNB 0.60fF
C84 a_277_1004.n8 VNB 0.46fF
C85 a_277_1004.n9 VNB 0.50fF
C86 a_277_1004.n10 VNB 2.48fF
C87 a_277_1004.n11 VNB 0.58fF
C88 a_277_1004.n12 VNB 0.04fF
C89 a_277_1004.n13 VNB 0.41fF
C90 a_277_1004.n14 VNB 0.07fF
C91 VPB.n0 VNB 0.03fF
C92 VPB.n1 VNB 0.04fF
C93 VPB.n2 VNB 0.02fF
C94 VPB.n3 VNB 0.19fF
C95 VPB.n5 VNB 0.02fF
C96 VPB.n6 VNB 0.02fF
C97 VPB.n7 VNB 0.02fF
C98 VPB.n8 VNB 0.02fF
C99 VPB.n10 VNB 0.02fF
C100 VPB.n11 VNB 0.02fF
C101 VPB.n12 VNB 0.02fF
C102 VPB.n14 VNB 0.10fF
C103 VPB.n15 VNB 0.10fF
C104 VPB.n16 VNB 0.02fF
C105 VPB.n17 VNB 0.02fF
C106 VPB.n18 VNB 0.02fF
C107 VPB.n19 VNB 0.04fF
C108 VPB.n20 VNB 0.02fF
C109 VPB.n21 VNB 0.25fF
C110 VPB.n22 VNB 0.04fF
C111 VPB.n24 VNB 0.02fF
C112 VPB.n25 VNB 0.02fF
C113 VPB.n26 VNB 0.02fF
C114 VPB.n27 VNB 0.02fF
C115 VPB.n29 VNB 0.02fF
C116 VPB.n30 VNB 0.02fF
C117 VPB.n31 VNB 0.02fF
C118 VPB.n33 VNB 0.27fF
C119 VPB.n35 VNB 0.03fF
C120 VPB.n36 VNB 0.02fF
C121 VPB.n37 VNB 0.03fF
C122 VPB.n38 VNB 0.03fF
C123 VPB.n39 VNB 0.27fF
C124 VPB.n40 VNB 0.01fF
C125 VPB.n41 VNB 0.02fF
C126 VPB.n42 VNB 0.27fF
C127 VPB.n43 VNB 0.02fF
C128 VPB.n44 VNB 0.02fF
C129 VPB.n45 VNB 0.05fF
C130 VPB.n46 VNB 0.21fF
C131 VPB.n47 VNB 0.02fF
C132 VPB.n48 VNB 0.01fF
C133 VPB.n49 VNB 0.14fF
C134 VPB.n50 VNB 0.16fF
C135 VPB.n51 VNB 0.02fF
C136 VPB.n52 VNB 0.02fF
C137 VPB.n53 VNB 0.14fF
C138 VPB.n54 VNB 0.16fF
C139 VPB.n55 VNB 0.02fF
C140 VPB.n56 VNB 0.02fF
C141 VPB.n57 VNB 0.02fF
C142 VPB.n58 VNB 0.14fF
C143 VPB.n59 VNB 0.15fF
C144 VPB.n60 VNB 0.02fF
C145 VPB.n61 VNB 0.02fF
C146 VPB.n62 VNB 0.14fF
C147 VPB.n63 VNB 0.15fF
C148 VPB.n64 VNB 0.02fF
C149 VPB.n65 VNB 0.02fF
C150 VPB.n66 VNB 0.02fF
C151 VPB.n67 VNB 0.14fF
C152 VPB.n68 VNB 0.16fF
C153 VPB.n69 VNB 0.02fF
C154 VPB.n70 VNB 0.02fF
C155 VPB.n71 VNB 0.14fF
C156 VPB.n72 VNB 0.16fF
C157 VPB.n73 VNB 0.02fF
C158 VPB.n74 VNB 0.02fF
C159 VPB.n75 VNB 0.21fF
C160 VPB.n76 VNB 0.02fF
C161 VPB.n77 VNB 0.01fF
C162 VPB.n78 VNB 0.06fF
C163 VPB.n79 VNB 0.27fF
C164 VPB.n80 VNB 0.02fF
C165 VPB.n81 VNB 0.02fF
C166 VPB.n82 VNB 0.02fF
C167 VPB.n83 VNB 0.02fF
C168 VPB.n84 VNB 0.02fF
C169 VPB.n85 VNB 0.02fF
C170 VPB.n86 VNB 0.04fF
C171 VPB.n87 VNB 0.02fF
C172 VPB.n88 VNB 0.20fF
C173 VPB.n89 VNB 0.04fF
C174 VPB.n91 VNB 0.02fF
C175 VPB.n92 VNB 0.02fF
C176 VPB.n93 VNB 0.02fF
C177 VPB.n94 VNB 0.02fF
C178 VPB.n96 VNB 0.02fF
C179 VPB.n97 VNB 0.02fF
C180 VPB.n98 VNB 0.02fF
C181 VPB.n100 VNB 0.27fF
C182 VPB.n102 VNB 0.03fF
C183 VPB.n103 VNB 0.02fF
C184 VPB.n104 VNB 0.10fF
C185 VPB.n105 VNB 0.02fF
C186 VPB.n106 VNB 0.02fF
C187 VPB.n107 VNB 0.02fF
C188 VPB.n108 VNB 0.04fF
C189 VPB.n109 VNB 0.02fF
C190 VPB.n110 VNB 0.20fF
C191 VPB.n111 VNB 0.04fF
C192 VPB.n113 VNB 0.02fF
C193 VPB.n114 VNB 0.02fF
C194 VPB.n115 VNB 0.02fF
C195 VPB.n116 VNB 0.02fF
C196 VPB.n118 VNB 0.02fF
C197 VPB.n119 VNB 0.02fF
C198 VPB.n120 VNB 0.02fF
C199 VPB.n122 VNB 0.27fF
C200 VPB.n124 VNB 0.03fF
C201 VPB.n125 VNB 0.02fF
C202 VPB.n126 VNB 0.27fF
C203 VPB.n127 VNB 0.01fF
C204 VPB.n128 VNB 0.02fF
C205 VPB.n129 VNB 0.03fF
C206 VPB.n130 VNB 0.03fF
C207 VPB.n131 VNB 0.27fF
C208 VPB.n132 VNB 0.01fF
C209 VPB.n133 VNB 0.02fF
C210 VPB.n134 VNB 0.23fF
C211 VPB.n135 VNB 0.02fF
C212 VPB.n136 VNB 0.01fF
C213 VPB.n137 VNB 0.05fF
C214 VPB.n138 VNB 0.14fF
C215 VPB.n139 VNB 0.16fF
C216 VPB.n140 VNB 0.02fF
C217 VPB.n141 VNB 0.02fF
C218 VPB.n142 VNB 0.14fF
C219 VPB.n143 VNB 0.15fF
C220 VPB.n144 VNB 0.02fF
C221 VPB.n145 VNB 0.02fF
C222 VPB.n146 VNB 0.02fF
C223 VPB.n147 VNB 0.14fF
C224 VPB.n148 VNB 0.15fF
C225 VPB.n149 VNB 0.02fF
C226 VPB.n150 VNB 0.02fF
C227 VPB.n151 VNB 0.14fF
C228 VPB.n152 VNB 0.16fF
C229 VPB.n153 VNB 0.02fF
C230 VPB.n154 VNB 0.02fF
C231 VPB.n155 VNB 0.06fF
C232 VPB.n156 VNB 0.24fF
C233 VPB.n157 VNB 0.02fF
C234 VPB.n158 VNB 0.01fF
C235 VPB.n159 VNB 0.27fF
C236 VPB.n160 VNB 0.01fF
C237 VPB.n161 VNB 0.02fF
C238 VPB.n162 VNB 0.03fF
C239 VPB.n163 VNB 0.02fF
C240 VPB.n164 VNB 0.02fF
C241 VPB.n165 VNB 0.02fF
C242 VPB.n166 VNB 0.14fF
C243 VPB.n167 VNB 0.03fF
C244 VPB.n168 VNB 0.02fF
C245 VPB.n169 VNB 0.05fF
C246 VPB.n170 VNB 0.01fF
C247 VPB.n172 VNB 0.02fF
C248 VPB.n173 VNB 0.02fF
C249 VPB.n174 VNB 0.02fF
C250 VPB.n175 VNB 0.02fF
C251 VPB.n177 VNB 0.02fF
C252 VPB.n180 VNB 0.46fF
C253 VPB.n182 VNB 0.04fF
C254 VPB.n183 VNB 0.04fF
C255 VPB.n184 VNB 0.27fF
C256 VPB.n185 VNB 0.03fF
C257 VPB.n186 VNB 0.04fF
C258 VPB.n187 VNB 0.10fF
C259 VPB.n188 VNB 0.02fF
C260 VPB.n189 VNB 0.14fF
C261 VPB.n190 VNB 0.15fF
C262 VPB.n191 VNB 0.02fF
C263 VPB.n192 VNB 0.02fF
C264 VPB.n193 VNB 0.14fF
C265 VPB.n194 VNB 0.16fF
C266 VPB.n195 VNB 0.02fF
C267 VPB.n196 VNB 0.02fF
C268 VPB.n197 VNB 0.05fF
C269 VPB.n198 VNB 0.23fF
C270 VPB.n199 VNB 0.02fF
C271 VPB.n200 VNB 0.01fF
C272 VPB.n201 VNB 0.00fF
C273 VPB.n202 VNB 0.10fF
C274 VPB.n203 VNB 0.02fF
C275 VPB.n204 VNB 0.14fF
C276 VPB.n205 VNB 0.15fF
C277 VPB.n206 VNB 0.02fF
C278 VPB.n207 VNB 0.02fF
C279 VPB.n208 VNB 0.02fF
C280 VPB.n209 VNB 0.14fF
C281 VPB.n210 VNB 0.16fF
C282 VPB.n211 VNB 0.02fF
C283 VPB.n212 VNB 0.02fF
C284 VPB.n213 VNB 0.02fF
C285 VPB.n214 VNB 0.06fF
C286 VPB.n215 VNB 0.24fF
C287 VPB.n216 VNB 0.02fF
C288 VPB.n217 VNB 0.01fF
C289 VPB.n218 VNB 0.02fF
C290 VPB.n219 VNB 0.27fF
C291 VPB.n220 VNB 0.01fF
C292 VPB.n221 VNB 0.02fF
C293 VPB.n222 VNB 0.04fF
C294 VPB.n223 VNB 0.02fF
C295 VPB.n224 VNB 0.02fF
C296 VPB.n225 VNB 0.02fF
C297 VPB.n226 VNB 0.04fF
C298 VPB.n227 VNB 0.02fF
C299 VPB.n228 VNB 0.20fF
C300 VPB.n229 VNB 0.04fF
C301 VPB.n231 VNB 0.02fF
C302 VPB.n232 VNB 0.02fF
C303 VPB.n233 VNB 0.02fF
C304 VPB.n234 VNB 0.02fF
C305 VPB.n236 VNB 0.02fF
C306 VPB.n237 VNB 0.02fF
C307 VPB.n238 VNB 0.02fF
C308 VPB.n240 VNB 0.27fF
C309 VPB.n242 VNB 0.03fF
C310 VPB.n243 VNB 0.02fF
C311 VPB.n244 VNB 0.03fF
C312 VPB.n245 VNB 0.03fF
C313 VPB.n246 VNB 0.27fF
C314 VPB.n247 VNB 0.01fF
C315 VPB.n248 VNB 0.02fF
C316 VPB.n249 VNB 0.04fF
C317 VPB.n250 VNB 0.05fF
C318 VPB.n251 VNB 0.23fF
C319 VPB.n252 VNB 0.02fF
C320 VPB.n253 VNB 0.01fF
C321 VPB.n254 VNB 0.02fF
C322 VPB.n255 VNB 0.14fF
C323 VPB.n256 VNB 0.16fF
C324 VPB.n257 VNB 0.02fF
C325 VPB.n258 VNB 0.02fF
C326 VPB.n259 VNB 0.02fF
C327 VPB.n260 VNB 0.10fF
C328 VPB.n261 VNB 0.02fF
C329 VPB.n262 VNB 0.14fF
C330 VPB.n263 VNB 0.15fF
C331 VPB.n264 VNB 0.02fF
C332 VPB.n265 VNB 0.02fF
C333 VPB.n266 VNB 0.02fF
C334 VPB.n267 VNB 0.14fF
C335 VPB.n268 VNB 0.15fF
C336 VPB.n269 VNB 0.02fF
C337 VPB.n270 VNB 0.02fF
C338 VPB.n271 VNB 0.02fF
C339 VPB.n272 VNB 0.14fF
C340 VPB.n273 VNB 0.16fF
C341 VPB.n274 VNB 0.02fF
C342 VPB.n275 VNB 0.02fF
C343 VPB.n276 VNB 0.02fF
C344 VPB.n277 VNB 0.06fF
C345 VPB.n278 VNB 0.24fF
C346 VPB.n279 VNB 0.02fF
C347 VPB.n280 VNB 0.01fF
C348 VPB.n281 VNB 0.02fF
C349 VPB.n282 VNB 0.04fF
C350 VPB.n283 VNB 0.04fF
C351 VPB.n284 VNB 0.02fF
C352 VPB.n285 VNB 0.02fF
C353 VPB.n286 VNB 0.02fF
C354 VPB.n287 VNB 0.02fF
C355 VPB.n288 VNB 0.02fF
C356 VPB.n289 VNB 0.02fF
C357 VPB.n290 VNB 0.04fF
C358 VPB.n291 VNB 0.04fF
C359 VPB.n292 VNB 0.03fF
C360 VPB.n293 VNB 0.27fF
C361 VPB.n294 VNB 0.01fF
C362 VPB.n295 VNB 0.02fF
C363 VPB.n296 VNB 0.23fF
C364 VPB.n297 VNB 0.02fF
C365 VPB.n298 VNB 0.01fF
C366 VPB.n299 VNB 0.05fF
C367 VPB.n300 VNB 0.14fF
C368 VPB.n301 VNB 0.16fF
C369 VPB.n302 VNB 0.02fF
C370 VPB.n303 VNB 0.02fF
C371 VPB.n304 VNB 0.02fF
C372 VPB.n305 VNB 0.10fF
C373 VPB.n306 VNB 0.02fF
C374 VPB.n307 VNB 0.14fF
C375 VPB.n308 VNB 0.15fF
C376 VPB.n309 VNB 0.02fF
C377 VPB.n310 VNB 0.02fF
C378 VPB.n311 VNB 0.02fF
C379 VPB.n312 VNB 0.14fF
C380 VPB.n313 VNB 0.15fF
C381 VPB.n314 VNB 0.02fF
C382 VPB.n315 VNB 0.02fF
C383 VPB.n316 VNB 0.02fF
C384 VPB.n317 VNB 0.14fF
C385 VPB.n318 VNB 0.16fF
C386 VPB.n319 VNB 0.02fF
C387 VPB.n320 VNB 0.02fF
C388 VPB.n321 VNB 0.02fF
C389 VPB.n322 VNB 0.06fF
C390 VPB.n323 VNB 0.24fF
C391 VPB.n324 VNB 0.02fF
C392 VPB.n325 VNB 0.01fF
C393 VPB.n326 VNB 0.02fF
C394 VPB.n327 VNB 0.27fF
C395 VPB.n328 VNB 0.01fF
C396 VPB.n329 VNB 0.02fF
C397 VPB.n330 VNB 0.04fF
C398 VPB.n331 VNB 0.02fF
C399 VPB.n332 VNB 0.02fF
C400 VPB.n333 VNB 0.02fF
C401 VPB.n334 VNB 0.04fF
C402 VPB.n335 VNB 0.02fF
C403 VPB.n336 VNB 0.20fF
C404 VPB.n337 VNB 0.04fF
C405 VPB.n339 VNB 0.02fF
C406 VPB.n340 VNB 0.02fF
C407 VPB.n341 VNB 0.02fF
C408 VPB.n342 VNB 0.02fF
C409 VPB.n344 VNB 0.02fF
C410 VPB.n345 VNB 0.02fF
C411 VPB.n346 VNB 0.02fF
C412 VPB.n348 VNB 0.27fF
C413 VPB.n350 VNB 0.03fF
C414 VPB.n351 VNB 0.02fF
C415 VPB.n352 VNB 0.03fF
C416 VPB.n353 VNB 0.03fF
C417 VPB.n354 VNB 0.27fF
C418 VPB.n355 VNB 0.01fF
C419 VPB.n356 VNB 0.02fF
C420 VPB.n357 VNB 0.04fF
C421 VPB.n358 VNB 0.05fF
C422 VPB.n359 VNB 0.23fF
C423 VPB.n360 VNB 0.02fF
C424 VPB.n361 VNB 0.01fF
C425 VPB.n362 VNB 0.02fF
C426 VPB.n363 VNB 0.14fF
C427 VPB.n364 VNB 0.16fF
C428 VPB.n365 VNB 0.02fF
C429 VPB.n366 VNB 0.02fF
C430 VPB.n367 VNB 0.02fF
C431 VPB.n368 VNB 0.10fF
C432 VPB.n369 VNB 0.02fF
C433 VPB.n370 VNB 0.14fF
C434 VPB.n371 VNB 0.15fF
C435 VPB.n372 VNB 0.02fF
C436 VPB.n373 VNB 0.02fF
C437 VPB.n374 VNB 0.02fF
C438 VPB.n375 VNB 0.14fF
C439 VPB.n376 VNB 0.15fF
C440 VPB.n377 VNB 0.02fF
C441 VPB.n378 VNB 0.02fF
C442 VPB.n379 VNB 0.02fF
C443 VPB.n380 VNB 0.14fF
C444 VPB.n381 VNB 0.16fF
C445 VPB.n382 VNB 0.02fF
C446 VPB.n383 VNB 0.02fF
C447 VPB.n384 VNB 0.02fF
C448 VPB.n385 VNB 0.06fF
C449 VPB.n386 VNB 0.24fF
C450 VPB.n387 VNB 0.02fF
C451 VPB.n388 VNB 0.01fF
C452 VPB.n389 VNB 0.02fF
C453 VPB.n390 VNB 0.27fF
C454 VPB.n391 VNB 0.01fF
C455 VPB.n392 VNB 0.02fF
C456 VPB.n393 VNB 0.04fF
C457 VPB.n394 VNB 0.04fF
C458 VPB.n395 VNB 0.02fF
C459 VPB.n396 VNB 0.02fF
C460 VPB.n397 VNB 0.02fF
C461 VPB.n398 VNB 0.02fF
C462 VPB.n399 VNB 0.02fF
C463 VPB.n400 VNB 0.02fF
C464 VPB.n401 VNB 0.02fF
C465 VPB.n402 VNB 0.02fF
C466 VPB.n403 VNB 0.02fF
C467 VPB.n404 VNB 0.02fF
C468 VPB.n405 VNB 0.03fF
C469 VPB.n406 VNB 0.04fF
C470 VPB.n407 VNB 0.02fF
C471 VPB.n408 VNB 0.02fF
C472 VPB.n409 VNB 0.02fF
C473 VPB.n410 VNB 0.04fF
C474 VPB.n411 VNB 0.04fF
C475 VPB.n413 VNB 0.43fF
C476 a_1845_1004.n0 VNB 0.04fF
C477 a_1845_1004.n1 VNB 0.53fF
C478 a_1845_1004.n2 VNB 0.62fF
C479 a_1845_1004.n3 VNB 0.32fF
C480 a_1845_1004.n4 VNB 0.38fF
C481 a_1845_1004.n5 VNB 0.56fF
C482 a_1845_1004.n6 VNB 0.59fF
C483 a_1845_1004.n7 VNB 0.03fF
C484 a_1845_1004.n8 VNB 0.28fF
C485 a_1845_1004.n9 VNB 0.05fF
C486 a_147_159.n0 VNB 0.06fF
C487 a_147_159.n1 VNB 0.73fF
C488 a_147_159.n2 VNB 0.86fF
C489 a_147_159.n3 VNB 0.35fF
C490 a_147_159.n4 VNB 0.39fF
C491 a_147_159.n5 VNB 0.55fF
C492 a_147_159.n6 VNB 0.39fF
C493 a_147_159.t10 VNB 0.78fF
C494 a_147_159.n7 VNB 0.51fF
C495 a_147_159.n8 VNB 0.39fF
C496 a_147_159.n9 VNB 0.73fF
C497 a_147_159.n10 VNB 2.41fF
C498 a_147_159.n11 VNB 1.79fF
C499 a_147_159.n12 VNB 0.57fF
C500 a_147_159.n13 VNB 0.05fF
C501 a_147_159.n14 VNB 0.47fF
C502 a_147_159.n15 VNB 0.07fF
.ends
