* SPICE3 file created from NAND2X1.ext - technology: sky130A

.subckt NAND2X1 Y A B VDD GND
M1000 GND A.t1 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1001 VDD.t3 A.t0 Y.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t0 B.t0 Y.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B.t1 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1004 Y.t4 A.t2 VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y.t1 B.t2 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 Y VDD 1.33fF
C1 A B 0.27fF
C2 Y A 0.10fF
C3 A VDD 0.08fF
C4 Y B 0.26fF
C5 B VDD 0.07fF
R0 A.n0 A.t0 480.392
R1 A.n0 A.t2 403.272
R2 A.n1 A.t1 310.033
R3 A A.n1 76
R4 A.n1 A.n0 71.894
R5 Y.n7 Y.n6 184.039
R6 Y.n7 Y.n2 179.052
R7 Y.n2 Y.n1 76.002
R8 Y Y.n7 76
R9 Y.n6 Y.n5 30
R10 Y.n4 Y.n3 24.383
R11 Y.n6 Y.n4 23.684
R12 Y.n0 Y.t0 14.282
R13 Y.n0 Y.t1 14.282
R14 Y.n1 Y.t3 14.282
R15 Y.n1 Y.t4 14.282
R16 Y.n2 Y.n0 12.85
R17 VDD.n78 VDD.n77 76
R18 VDD.n73 VDD.n72 76
R19 VDD.n68 VDD.n67 76
R20 VDD.n63 VDD.n62 76
R21 VDD.n64 VDD.t2 55.106
R22 VDD.n33 VDD.t0 55.106
R23 VDD.n28 VDD.n27 40.824
R24 VDD.n25 VDD.n24 36.608
R25 VDD.n38 VDD.n37 34.942
R26 VDD.n70 VDD.n69 32.032
R27 VDD.n62 VDD.n59 21.841
R28 VDD.n23 VDD.n20 21.841
R29 VDD.n27 VDD.t1 14.282
R30 VDD.n27 VDD.t3 14.282
R31 VDD.n59 VDD.n41 14.167
R32 VDD.n41 VDD.n40 14.167
R33 VDD.n20 VDD.n19 14.167
R34 VDD.n19 VDD.n17 14.167
R35 VDD.n32 VDD.n31 14.167
R36 VDD.n23 VDD.n22 13.653
R37 VDD.n22 VDD.n21 13.653
R38 VDD.n36 VDD.n35 13.653
R39 VDD.n35 VDD.n34 13.653
R40 VDD.n32 VDD.n26 13.653
R41 VDD.n26 VDD.n25 13.653
R42 VDD.n31 VDD.n30 13.653
R43 VDD.n30 VDD.n29 13.653
R44 VDD.n77 VDD.n76 13.653
R45 VDD.n76 VDD.n75 13.653
R46 VDD.n72 VDD.n71 13.653
R47 VDD.n71 VDD.n70 13.653
R48 VDD.n67 VDD.n66 13.653
R49 VDD.n66 VDD.n65 13.653
R50 VDD.n62 VDD.n61 13.653
R51 VDD.n61 VDD.n60 13.653
R52 VDD.n4 VDD.n2 12.915
R53 VDD.n4 VDD.n3 12.66
R54 VDD.n10 VDD.n9 12.343
R55 VDD.n12 VDD.n11 12.343
R56 VDD.n10 VDD.n7 12.343
R57 VDD.n33 VDD.n32 11.806
R58 VDD.n31 VDD.n28 8.658
R59 VDD.n45 VDD.n44 7.5
R60 VDD.n48 VDD.n47 7.5
R61 VDD.n50 VDD.n49 7.5
R62 VDD.n53 VDD.n52 7.5
R63 VDD.n59 VDD.n58 7.5
R64 VDD.n20 VDD.n16 7.5
R65 VDD.n2 VDD.n1 7.5
R66 VDD.n9 VDD.n8 7.5
R67 VDD.n7 VDD.n6 7.5
R68 VDD.n19 VDD.n18 7.5
R69 VDD.n14 VDD.n0 7.5
R70 VDD.n58 VDD.n57 6.772
R71 VDD.n46 VDD.n43 6.772
R72 VDD.n51 VDD.n48 6.772
R73 VDD.n55 VDD.n53 6.772
R74 VDD.n55 VDD.n54 6.772
R75 VDD.n51 VDD.n50 6.772
R76 VDD.n46 VDD.n45 6.772
R77 VDD.n57 VDD.n42 6.772
R78 VDD.n37 VDD.n23 6.487
R79 VDD.n37 VDD.n36 6.475
R80 VDD.n16 VDD.n15 6.458
R81 VDD.n75 VDD.n74 4.576
R82 VDD.n67 VDD.n64 2.754
R83 VDD.n36 VDD.n33 2.361
R84 VDD.n14 VDD.n5 1.329
R85 VDD.n14 VDD.n10 1.329
R86 VDD.n14 VDD.n12 1.329
R87 VDD.n14 VDD.n13 1.329
R88 VDD.n15 VDD.n14 0.696
R89 VDD.n14 VDD.n4 0.696
R90 VDD.n56 VDD.n55 0.365
R91 VDD.n56 VDD.n51 0.365
R92 VDD.n56 VDD.n46 0.365
R93 VDD.n57 VDD.n56 0.365
R94 VDD.n63 VDD 0.207
R95 VDD.n39 VDD.n38 0.145
R96 VDD.n78 VDD.n73 0.145
R97 VDD.n73 VDD.n68 0.145
R98 VDD.n68 VDD.n63 0.145
R99 VDD VDD.n39 0.09
R100 VDD VDD.n78 0.09
R101 a_112_101.t0 a_112_101.n1 93.333
R102 a_112_101.n4 a_112_101.n2 55.07
R103 a_112_101.t0 a_112_101.n0 8.137
R104 a_112_101.n4 a_112_101.n3 4.619
R105 a_112_101.t0 a_112_101.n4 0.071
R106 GND.n17 GND.n16 84.842
R107 GND.n12 GND.n11 76
R108 GND.n23 GND.n22 76
R109 GND.n20 GND.n19 76
R110 GND.n15 GND.n14 76
R111 GND.n8 GND.n7 34.942
R112 GND.n6 GND.n5 14.167
R113 GND.n5 GND.n4 14.167
R114 GND.n14 GND.n13 13.653
R115 GND.n19 GND.n18 13.653
R116 GND.n22 GND.n21 13.653
R117 GND.n4 GND.n3 13.653
R118 GND.n5 GND.n2 13.653
R119 GND.n6 GND.n1 13.653
R120 GND.n7 GND.n0 7.083
R121 GND.n7 GND.n6 6.474
R122 GND.n19 GND.n17 3.935
R123 GND.n11 GND.n10 0.596
R124 GND.n12 GND 0.207
R125 GND.n9 GND.n8 0.145
R126 GND.n23 GND.n20 0.145
R127 GND.n20 GND.n15 0.145
R128 GND.n15 GND.n12 0.145
R129 GND GND.n9 0.09
R130 GND GND.n23 0.09
R131 B.n0 B.t0 472.359
R132 B.n0 B.t2 384.527
R133 B.n1 B.t1 241.172
R134 B.n1 B.n0 110.06
R135 B B.n1 76
C6 VDD GND 3.28fF
C7 a_112_101.n0 GND 0.05fF
C8 a_112_101.n1 GND 0.02fF
C9 a_112_101.n2 GND 0.11fF
C10 a_112_101.n3 GND 0.04fF
C11 a_112_101.n4 GND 0.15fF
C12 VDD.n0 GND 0.14fF
C13 VDD.n1 GND 0.02fF
C14 VDD.n2 GND 0.02fF
C15 VDD.n3 GND 0.04fF
C16 VDD.n4 GND 0.01fF
C17 VDD.n6 GND 0.02fF
C18 VDD.n7 GND 0.02fF
C19 VDD.n8 GND 0.02fF
C20 VDD.n9 GND 0.02fF
C21 VDD.n11 GND 0.02fF
C22 VDD.n14 GND 0.41fF
C23 VDD.n16 GND 0.03fF
C24 VDD.n17 GND 0.02fF
C25 VDD.n18 GND 0.02fF
C26 VDD.n19 GND 0.02fF
C27 VDD.n20 GND 0.03fF
C28 VDD.n21 GND 0.25fF
C29 VDD.n22 GND 0.02fF
C30 VDD.n23 GND 0.03fF
C31 VDD.n24 GND 0.12fF
C32 VDD.n25 GND 0.15fF
C33 VDD.n26 GND 0.01fF
C34 VDD.n27 GND 0.10fF
C35 VDD.n28 GND 0.02fF
C36 VDD.n29 GND 0.27fF
C37 VDD.n30 GND 0.01fF
C38 VDD.n31 GND 0.02fF
C39 VDD.n32 GND 0.02fF
C40 VDD.n33 GND 0.05fF
C41 VDD.n34 GND 0.22fF
C42 VDD.n35 GND 0.01fF
C43 VDD.n36 GND 0.01fF
C44 VDD.n37 GND 0.00fF
C45 VDD.n38 GND 0.08fF
C46 VDD.n39 GND 0.02fF
C47 VDD.n40 GND 0.02fF
C48 VDD.n41 GND 0.02fF
C49 VDD.n42 GND 0.02fF
C50 VDD.n43 GND 0.02fF
C51 VDD.n44 GND 0.02fF
C52 VDD.n45 GND 0.02fF
C53 VDD.n47 GND 0.02fF
C54 VDD.n48 GND 0.02fF
C55 VDD.n49 GND 0.02fF
C56 VDD.n50 GND 0.02fF
C57 VDD.n52 GND 0.03fF
C58 VDD.n53 GND 0.02fF
C59 VDD.n54 GND 0.14fF
C60 VDD.n56 GND 0.41fF
C61 VDD.n58 GND 0.03fF
C62 VDD.n59 GND 0.03fF
C63 VDD.n60 GND 0.25fF
C64 VDD.n61 GND 0.02fF
C65 VDD.n62 GND 0.03fF
C66 VDD.n63 GND 0.02fF
C67 VDD.n64 GND 0.05fF
C68 VDD.n65 GND 0.22fF
C69 VDD.n66 GND 0.01fF
C70 VDD.n67 GND 0.01fF
C71 VDD.n68 GND 0.02fF
C72 VDD.n69 GND 0.12fF
C73 VDD.n70 GND 0.15fF
C74 VDD.n71 GND 0.01fF
C75 VDD.n72 GND 0.02fF
C76 VDD.n73 GND 0.02fF
C77 VDD.n74 GND 0.15fF
C78 VDD.n75 GND 0.13fF
C79 VDD.n76 GND 0.01fF
C80 VDD.n77 GND 0.02fF
C81 VDD.n78 GND 0.02fF
C82 Y.n0 GND 0.47fF
C83 Y.n1 GND 0.56fF
C84 Y.n2 GND 0.30fF
C85 Y.n3 GND 0.04fF
C86 Y.n4 GND 0.05fF
C87 Y.n5 GND 0.03fF
C88 Y.n6 GND 0.24fF
C89 Y.n7 GND 0.38fF
.ends
