magic
tech sky130A
magscale 1 2
timestamp 1652395942
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 3461 945 3495 979
rect 4127 945 4161 979
rect 427 871 461 905
rect 2647 871 2681 905
rect 3313 871 3347 905
rect 3461 871 3495 905
rect 3831 871 3865 905
rect 4127 871 4161 905
rect 4127 797 4161 831
rect 427 723 461 757
rect 3313 723 3347 757
rect 4127 723 4161 757
rect 427 649 461 683
rect 2647 649 2681 683
rect 3313 649 3347 683
rect 3461 649 3495 683
rect 3831 649 3865 683
rect 4127 649 4161 683
rect 427 575 461 609
rect 1315 575 1349 609
rect 2647 575 2681 609
rect 3313 575 3347 609
rect 3461 575 3495 609
rect 3831 575 3865 609
rect 4127 575 4161 609
rect 427 501 461 535
rect 1315 501 1349 535
rect 2647 501 2681 535
rect 3313 501 3347 535
rect 3461 501 3495 535
rect 3831 501 3865 535
rect 4127 501 4161 535
rect 427 427 461 461
rect 1315 427 1349 461
rect 2647 427 2681 461
rect 3313 427 3347 461
rect 3461 427 3495 461
rect 3831 427 3865 461
rect 4127 427 4161 461
<< metal1 >>
rect -34 1445 4326 1514
rect 3349 723 4115 757
rect 3497 649 3807 683
rect -34 -34 4326 34
use dffx1_pcell  dffx1_pcell_0 pcells
timestamp 1652395794
transform 1 0 0 0 1 0
box -87 -34 4379 1550
use li1_M1_contact  li1_M1_contact_15 pcells
timestamp 1648061256
transform 1 0 4144 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform -1 0 3330 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 3478 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 3848 0 1 666
box -53 -33 29 33
<< labels >>
rlabel locali 4127 723 4161 757 1 Q
port 1 nsew signal output
rlabel locali 4127 797 4161 831 1 Q
port 1 nsew signal output
rlabel locali 4127 871 4161 905 1 Q
port 1 nsew signal output
rlabel locali 4127 945 4161 979 1 Q
port 1 nsew signal output
rlabel locali 4127 649 4161 683 1 Q
port 1 nsew signal output
rlabel locali 4127 575 4161 609 1 Q
port 1 nsew signal output
rlabel locali 4127 501 4161 535 1 Q
port 1 nsew signal output
rlabel locali 4127 427 4161 461 1 Q
port 1 nsew signal output
rlabel locali 3313 871 3347 905 1 Q
port 1 nsew signal output
rlabel locali 3313 723 3347 757 1 Q
port 1 nsew signal output
rlabel locali 3313 649 3347 683 1 Q
port 1 nsew signal output
rlabel locali 3313 575 3347 609 1 Q
port 1 nsew signal output
rlabel locali 3313 501 3347 535 1 Q
port 1 nsew signal output
rlabel locali 3313 427 3347 461 1 Q
port 1 nsew signal output
rlabel locali 3831 649 3865 683 1 QN
port 2 nsew signal output
rlabel locali 3831 871 3865 905 1 QN
port 2 nsew signal output
rlabel locali 3831 575 3865 609 1 QN
port 2 nsew signal output
rlabel locali 3831 501 3865 535 1 QN
port 2 nsew signal output
rlabel locali 3831 427 3865 461 1 QN
port 2 nsew signal output
rlabel locali 3461 427 3495 461 1 QN
port 2 nsew signal output
rlabel locali 3461 501 3495 535 1 QN
port 2 nsew signal output
rlabel locali 3461 575 3495 609 1 QN
port 2 nsew signal output
rlabel locali 3461 649 3495 683 1 QN
port 2 nsew signal output
rlabel locali 3461 871 3495 905 1 QN
port 2 nsew signal output
rlabel locali 3461 945 3495 979 1 QN
port 2 nsew signal output
rlabel locali 1315 575 1349 609 1 D
port 3 nsew signal input
rlabel locali 1315 501 1349 535 1 D
port 3 nsew signal input
rlabel locali 1315 427 1349 461 1 D
port 3 nsew signal input
rlabel locali 427 871 461 905 1 CLK
port 4 nsew signal input
rlabel locali 427 723 461 757 1 CLK
port 4 nsew signal input
rlabel locali 427 649 461 683 1 CLK
port 4 nsew signal input
rlabel locali 427 575 461 609 1 CLK
port 4 nsew signal input
rlabel locali 427 501 461 535 1 CLK
port 4 nsew signal input
rlabel locali 427 427 461 461 1 CLK
port 4 nsew signal input
rlabel locali 2647 427 2681 461 1 CLK
port 4 nsew signal input
rlabel locali 2647 501 2681 535 1 CLK
port 4 nsew signal input
rlabel locali 2647 575 2681 609 1 CLK
port 4 nsew signal input
rlabel locali 2647 649 2681 683 1 CLK
port 4 nsew signal input
rlabel locali 2647 871 2681 905 1 CLK
port 4 nsew signal input
rlabel metal1 -34 1445 4326 1514 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 -34 -34 4326 34 1 GND
port 6 nsew ground bidirectional abutment


<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 4292 1480
string LEFsymmetry X Y R90
<< end >>
