* SPICE3 file created from TMRDFFSNQNX1.ext - technology: sky130A

.subckt TMRDFFSNQNX1 QN D CLK SN VDD GND
M1000 a_8357_1050.t2 a_8483_411.t7 VDD.t34 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_3599_411.t1 a_3473_1050.t5 VDD.t40 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VDD.t86 CLK.t0 a_6149_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD.t32 a_8483_411.t8 a_14869_1051.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 GND a_11673_1050.t7 a_12470_101.t0 nshort w=-1.605u l=1.765u
+  ad=3.7611p pd=32.97u as=0p ps=0u
M1005 a_343_411.t5 a_1265_989.t5 VDD.t56 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_13367_411.t2 a_11033_989.t5 VDD.t39 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VDD.t46 a_343_411.t7 a_3473_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_5227_411.t4 a_5101_1050.t5 VDD.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 VDD.t10 SN.t2 a_8483_411.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1265_989.t3 CLK.t1 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 GND a_8483_411.t9 a_15430_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1012 VDD.t63 SN.t3 a_1905_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_11673_1050.t3 a_9985_1050.t6 VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t42 CLK.t2 a_5227_411.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_15533_1051.t3 a_3599_411.t7 QN.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_3599_411.t3 SN.t4 VDD.t65 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 GND a_217_1050.t5 a_757_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1018 QN a_13367_411.t9 a_16096_101.t0 nshort w=-1.83u l=2.06u
+  ad=0.5373p pd=4.72u as=0p ps=0u
M1019 VDD.t5 CLK.t4 a_11033_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 GND D.t2 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1021 VDD.t64 a_8357_1050.t5 a_8483_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_5227_411.t5 CLK.t5 VDD.t92 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 GND a_343_411.t8 a_3368_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1024 VDD.t9 D.t0 a_5101_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_14869_1051.t1 a_3599_411.t8 a_15533_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VDD.t22 D.t1 a_217_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VDD.t14 a_1265_989.t7 a_1905_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_9985_1050.t4 a_10111_411.t7 VDD.t87 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 GND a_8357_1050.t6 a_8897_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1030 VDD.t24 a_5101_1050.t6 a_6789_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_15533_1051.t5 a_13367_411.t8 QN.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 VDD.t7 a_11033_989.t7 a_11673_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_3599_411.t5 a_1265_989.t9 VDD.t55 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_6789_1050.t2 a_6149_989.t5 VDD.t82 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_13241_1050.t1 a_10111_411.t8 VDD.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1905_1050.t2 a_217_1050.t6 VDD.t53 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VDD.t29 a_11673_1050.t8 a_11033_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_14869_1051.t3 a_8483_411.t10 a_15533_1051.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 VDD.t89 a_343_411.t9 a_217_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 VDD.t47 a_5227_411.t8 a_5101_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 GND D.t3 a_9880_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1042 VDD.t37 a_217_1050.t7 a_343_411.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_11673_1050.t4 a_11033_989.t8 VDD.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1044 VDD.t77 a_13241_1050.t5 a_13367_411.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1045 GND a_217_1050.t8 a_1719_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_3473_1050.t2 a_3599_411.t9 VDD.t50 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_10111_411.t3 CLK.t7 VDD.t61 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 QN a_3599_411.t10 a_15430_101.t0 nshort w=-1.235u l=1.535u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_5227_411.t2 a_6149_989.t8 VDD.t81 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_13241_1050.t4 a_13367_411.t10 VDD.t74 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1051 VDD.t36 a_11033_989.t9 a_10111_411.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 VDD.t59 a_5227_411.t9 a_8357_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 a_6149_989.t1 CLK.t8 VDD.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_14869_1051.t4 a_8483_411.t11 VDD.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 a_13367_411.t3 a_13241_1050.t6 VDD.t76 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 VDD.t73 a_6149_989.t9 a_8483_411.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 VDD.t85 a_13367_411.t11 a_14869_1051.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 VDD.t41 CLK.t9 a_343_411.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1059 GND a_10111_411.t11 a_13136_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1060 GND a_1905_1050.t8 a_2702_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1061 a_3473_1050.t0 a_343_411.t10 VDD.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 VDD.t60 a_1905_1050.t7 a_1265_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 a_8483_411.t3 SN.t7 VDD.t72 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1064 VDD.t68 SN.t8 a_13367_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 a_10111_411.t1 a_9985_1050.t7 VDD.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 GND a_13241_1050.t7 a_13781_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1067 GND a_5227_411.t10 a_8252_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_15533_1051.t6 a_8483_411.t12 a_14869_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 VDD.t52 a_10111_411.t9 a_9985_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 VDD.t70 SN.t9 a_11673_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 GND a_5101_1050.t9 a_5641_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1072 a_6149_989.t0 a_6789_1050.t7 VDD.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1073 VDD.t43 a_3473_1050.t6 a_3599_411.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1074 VDD.t88 a_1265_989.t10 a_3599_411.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 GND a_8483_411.t13 a_14764_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1076 VDD.t13 a_1265_989.t11 a_343_411.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 a_8483_411.t2 a_8357_1050.t7 VDD.t69 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1078 VDD.t90 a_11033_989.t11 a_13367_411.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 VDD.t48 a_5101_1050.t7 a_5227_411.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 a_15533_1051.t0 a_3599_411.t11 a_14869_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 a_8483_411.t6 a_6149_989.t10 VDD.t80 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1082 a_217_1050.t3 D.t4 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 VDD.t11 D.t5 a_9985_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 a_1905_1050.t5 a_1265_989.t12 VDD.t45 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 a_6789_1050.t5 a_5101_1050.t8 VDD.t51 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 VDD.t38 a_9985_1050.t8 a_11673_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 GND a_5101_1050.t10 a_6603_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1088 QN.t5 a_13367_411.t12 a_15533_1051.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 GND a_3473_1050.t7 a_4013_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1090 VDD.t66 SN.t12 a_3599_411.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 VDD.t27 SN.t13 a_6789_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1092 QN a_13367_411.t13 a_14764_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1093 a_11033_989.t0 a_11673_1050.t9 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 GND a_6789_1050.t9 a_7586_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1095 a_1905_1050.t0 SN.t14 VDD.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1096 a_217_1050.t0 a_343_411.t12 VDD.t57 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 a_5101_1050.t1 a_5227_411.t11 VDD.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 GND a_9985_1050.t10 a_10525_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1099 GND a_3599_411.t14 a_16096_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1100 GND D.t7 a_4996_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1101 a_6789_1050.t3 SN.t15 VDD.t35 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 QN.t0 a_3599_411.t13 a_15533_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 VDD.t44 a_9985_1050.t9 a_10111_411.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 a_343_411.t0 a_217_1050.t9 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 VDD.t33 a_8483_411.t14 a_8357_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 VDD.t79 a_6149_989.t11 a_6789_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 a_10111_411.t5 a_11033_989.t13 VDD.t58 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 VDD.t19 a_10111_411.t12 a_13241_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 VDD.t62 a_217_1050.t10 a_1905_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 a_8357_1050.t3 a_5227_411.t12 VDD.t49 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 VDD.t54 a_6789_1050.t8 a_6149_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1112 a_11033_989.t3 CLK.t13 VDD.t83 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1113 a_5101_1050.t4 D.t6 VDD.t84 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1114 a_14869_1051.t6 a_13367_411.t14 VDD.t67 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1115 a_343_411.t1 CLK.t14 VDD.t93 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1116 GND a_9985_1050.t5 a_11487_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1117 a_9985_1050.t1 D.t8 VDD.t23 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1118 a_13367_411.t0 SN.t16 VDD.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1119 a_1265_989.t0 a_1905_1050.t9 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1120 VDD.t91 a_3599_411.t15 a_3473_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1121 VDD.t75 CLK.t15 a_10111_411.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1122 a_11673_1050.t0 SN.t17 VDD.t71 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1123 VDD.t4 CLK.t17 a_1265_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1124 VDD.t78 a_6149_989.t13 a_5227_411.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1125 VDD.t26 a_13367_411.t15 a_13241_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VDD D 0.24fF
C1 VDD CLK 1.68fF
C2 QN VDD 0.29fF
C3 D CLK 0.39fF
C4 VDD SN 0.30fF
C5 D SN 9.38fF
C6 CLK SN 0.46fF
R0 a_8483_411.n8 a_8483_411.t8 512.525
R1 a_8483_411.n6 a_8483_411.t10 477.179
R2 a_8483_411.n11 a_8483_411.t14 472.359
R3 a_8483_411.n6 a_8483_411.t12 406.485
R4 a_8483_411.n11 a_8483_411.t7 384.527
R5 a_8483_411.n8 a_8483_411.t11 371.139
R6 a_8483_411.n7 a_8483_411.t9 363.924
R7 a_8483_411.n10 a_8483_411.t13 277.053
R8 a_8483_411.n12 a_8483_411.t15 241.172
R9 a_8483_411.n16 a_8483_411.n14 213.104
R10 a_8483_411.n14 a_8483_411.n5 170.799
R11 a_8483_411.n12 a_8483_411.n11 110.06
R12 a_8483_411.n9 a_8483_411.n7 101.359
R13 a_8483_411.n13 a_8483_411.n10 94.999
R14 a_8483_411.n10 a_8483_411.n9 80.444
R15 a_8483_411.n13 a_8483_411.n12 80.035
R16 a_8483_411.n4 a_8483_411.n3 79.232
R17 a_8483_411.n14 a_8483_411.n13 76
R18 a_8483_411.n9 a_8483_411.n8 71.88
R19 a_8483_411.n5 a_8483_411.n4 63.152
R20 a_8483_411.n17 a_8483_411.n0 55.263
R21 a_8483_411.n16 a_8483_411.n15 30
R22 a_8483_411.n17 a_8483_411.n16 23.684
R23 a_8483_411.n5 a_8483_411.n1 16.08
R24 a_8483_411.n4 a_8483_411.n2 16.08
R25 a_8483_411.n7 a_8483_411.n6 15.776
R26 a_8483_411.n1 a_8483_411.t4 14.282
R27 a_8483_411.n1 a_8483_411.t6 14.282
R28 a_8483_411.n2 a_8483_411.t0 14.282
R29 a_8483_411.n2 a_8483_411.t3 14.282
R30 a_8483_411.n3 a_8483_411.t1 14.282
R31 a_8483_411.n3 a_8483_411.t2 14.282
R32 VDD.n809 VDD.n807 144.705
R33 VDD.n890 VDD.n888 144.705
R34 VDD.n971 VDD.n969 144.705
R35 VDD.n1032 VDD.n1030 144.705
R36 VDD.n1093 VDD.n1091 144.705
R37 VDD.n1174 VDD.n1172 144.705
R38 VDD.n1235 VDD.n1233 144.705
R39 VDD.n1316 VDD.n1314 144.705
R40 VDD.n1397 VDD.n1395 144.705
R41 VDD.n698 VDD.n696 144.705
R42 VDD.n1458 VDD.n1456 144.705
R43 VDD.n617 VDD.n615 144.705
R44 VDD.n556 VDD.n554 144.705
R45 VDD.n475 VDD.n473 144.705
R46 VDD.n394 VDD.n392 144.705
R47 VDD.n333 VDD.n331 144.705
R48 VDD.n272 VDD.n270 144.705
R49 VDD.n191 VDD.n189 144.705
R50 VDD.n130 VDD.n128 144.705
R51 VDD.n76 VDD.n74 144.705
R52 VDD.n39 VDD.n38 76
R53 VDD.n43 VDD.n42 76
R54 VDD.n47 VDD.n46 76
R55 VDD.n51 VDD.n50 76
R56 VDD.n78 VDD.n77 76
R57 VDD.n82 VDD.n81 76
R58 VDD.n86 VDD.n85 76
R59 VDD.n90 VDD.n89 76
R60 VDD.n94 VDD.n93 76
R61 VDD.n98 VDD.n97 76
R62 VDD.n102 VDD.n101 76
R63 VDD.n106 VDD.n105 76
R64 VDD.n132 VDD.n131 76
R65 VDD.n137 VDD.n136 76
R66 VDD.n142 VDD.n141 76
R67 VDD.n148 VDD.n147 76
R68 VDD.n153 VDD.n152 76
R69 VDD.n158 VDD.n157 76
R70 VDD.n163 VDD.n162 76
R71 VDD.n167 VDD.n166 76
R72 VDD.n193 VDD.n192 76
R73 VDD.n197 VDD.n196 76
R74 VDD.n201 VDD.n200 76
R75 VDD.n206 VDD.n205 76
R76 VDD.n213 VDD.n212 76
R77 VDD.n218 VDD.n217 76
R78 VDD.n223 VDD.n222 76
R79 VDD.n230 VDD.n229 76
R80 VDD.n235 VDD.n234 76
R81 VDD.n240 VDD.n239 76
R82 VDD.n244 VDD.n243 76
R83 VDD.n248 VDD.n247 76
R84 VDD.n274 VDD.n273 76
R85 VDD.n279 VDD.n278 76
R86 VDD.n284 VDD.n283 76
R87 VDD.n290 VDD.n289 76
R88 VDD.n295 VDD.n294 76
R89 VDD.n300 VDD.n299 76
R90 VDD.n305 VDD.n304 76
R91 VDD.n309 VDD.n308 76
R92 VDD.n335 VDD.n334 76
R93 VDD.n340 VDD.n339 76
R94 VDD.n345 VDD.n344 76
R95 VDD.n351 VDD.n350 76
R96 VDD.n356 VDD.n355 76
R97 VDD.n361 VDD.n360 76
R98 VDD.n366 VDD.n365 76
R99 VDD.n370 VDD.n369 76
R100 VDD.n396 VDD.n395 76
R101 VDD.n400 VDD.n399 76
R102 VDD.n404 VDD.n403 76
R103 VDD.n409 VDD.n408 76
R104 VDD.n416 VDD.n415 76
R105 VDD.n421 VDD.n420 76
R106 VDD.n426 VDD.n425 76
R107 VDD.n433 VDD.n432 76
R108 VDD.n438 VDD.n437 76
R109 VDD.n443 VDD.n442 76
R110 VDD.n447 VDD.n446 76
R111 VDD.n451 VDD.n450 76
R112 VDD.n477 VDD.n476 76
R113 VDD.n481 VDD.n480 76
R114 VDD.n485 VDD.n484 76
R115 VDD.n490 VDD.n489 76
R116 VDD.n497 VDD.n496 76
R117 VDD.n502 VDD.n501 76
R118 VDD.n507 VDD.n506 76
R119 VDD.n514 VDD.n513 76
R120 VDD.n519 VDD.n518 76
R121 VDD.n524 VDD.n523 76
R122 VDD.n528 VDD.n527 76
R123 VDD.n532 VDD.n531 76
R124 VDD.n558 VDD.n557 76
R125 VDD.n563 VDD.n562 76
R126 VDD.n568 VDD.n567 76
R127 VDD.n574 VDD.n573 76
R128 VDD.n579 VDD.n578 76
R129 VDD.n584 VDD.n583 76
R130 VDD.n589 VDD.n588 76
R131 VDD.n593 VDD.n592 76
R132 VDD.n619 VDD.n618 76
R133 VDD.n623 VDD.n622 76
R134 VDD.n627 VDD.n626 76
R135 VDD.n632 VDD.n631 76
R136 VDD.n639 VDD.n638 76
R137 VDD.n644 VDD.n643 76
R138 VDD.n649 VDD.n648 76
R139 VDD.n656 VDD.n655 76
R140 VDD.n661 VDD.n660 76
R141 VDD.n666 VDD.n665 76
R142 VDD.n670 VDD.n669 76
R143 VDD.n674 VDD.n673 76
R144 VDD.n700 VDD.n699 76
R145 VDD.n705 VDD.n704 76
R146 VDD.n710 VDD.n709 76
R147 VDD.n716 VDD.n715 76
R148 VDD.n721 VDD.n720 76
R149 VDD.n726 VDD.n725 76
R150 VDD.n1465 VDD.n1464 76
R151 VDD.n1460 VDD.n1459 76
R152 VDD.n1434 VDD.n1433 76
R153 VDD.n1430 VDD.n1429 76
R154 VDD.n1425 VDD.n1424 76
R155 VDD.n1420 VDD.n1419 76
R156 VDD.n1414 VDD.n1413 76
R157 VDD.n1409 VDD.n1408 76
R158 VDD.n1404 VDD.n1403 76
R159 VDD.n1399 VDD.n1398 76
R160 VDD.n1373 VDD.n1372 76
R161 VDD.n1369 VDD.n1368 76
R162 VDD.n1365 VDD.n1364 76
R163 VDD.n1361 VDD.n1360 76
R164 VDD.n1356 VDD.n1355 76
R165 VDD.n1349 VDD.n1348 76
R166 VDD.n1344 VDD.n1343 76
R167 VDD.n1339 VDD.n1338 76
R168 VDD.n1332 VDD.n1331 76
R169 VDD.n1327 VDD.n1326 76
R170 VDD.n1322 VDD.n1321 76
R171 VDD.n1318 VDD.n1317 76
R172 VDD.n1292 VDD.n1291 76
R173 VDD.n1288 VDD.n1287 76
R174 VDD.n1284 VDD.n1283 76
R175 VDD.n1280 VDD.n1279 76
R176 VDD.n1275 VDD.n1274 76
R177 VDD.n1268 VDD.n1267 76
R178 VDD.n1263 VDD.n1262 76
R179 VDD.n1258 VDD.n1257 76
R180 VDD.n1251 VDD.n1250 76
R181 VDD.n1246 VDD.n1245 76
R182 VDD.n1241 VDD.n1240 76
R183 VDD.n1237 VDD.n1236 76
R184 VDD.n1211 VDD.n1210 76
R185 VDD.n1207 VDD.n1206 76
R186 VDD.n1202 VDD.n1201 76
R187 VDD.n1197 VDD.n1196 76
R188 VDD.n1191 VDD.n1190 76
R189 VDD.n1186 VDD.n1185 76
R190 VDD.n1181 VDD.n1180 76
R191 VDD.n1176 VDD.n1175 76
R192 VDD.n1150 VDD.n1149 76
R193 VDD.n1146 VDD.n1145 76
R194 VDD.n1142 VDD.n1141 76
R195 VDD.n1138 VDD.n1137 76
R196 VDD.n1133 VDD.n1132 76
R197 VDD.n1126 VDD.n1125 76
R198 VDD.n1121 VDD.n1120 76
R199 VDD.n1116 VDD.n1115 76
R200 VDD.n1109 VDD.n1108 76
R201 VDD.n1104 VDD.n1103 76
R202 VDD.n1099 VDD.n1098 76
R203 VDD.n1095 VDD.n1094 76
R204 VDD.n1069 VDD.n1068 76
R205 VDD.n1065 VDD.n1064 76
R206 VDD.n1060 VDD.n1059 76
R207 VDD.n1055 VDD.n1054 76
R208 VDD.n1049 VDD.n1048 76
R209 VDD.n1044 VDD.n1043 76
R210 VDD.n1039 VDD.n1038 76
R211 VDD.n1034 VDD.n1033 76
R212 VDD.n1008 VDD.n1007 76
R213 VDD.n1004 VDD.n1003 76
R214 VDD.n999 VDD.n998 76
R215 VDD.n994 VDD.n993 76
R216 VDD.n988 VDD.n987 76
R217 VDD.n983 VDD.n982 76
R218 VDD.n978 VDD.n977 76
R219 VDD.n973 VDD.n972 76
R220 VDD.n947 VDD.n946 76
R221 VDD.n943 VDD.n942 76
R222 VDD.n939 VDD.n938 76
R223 VDD.n935 VDD.n934 76
R224 VDD.n930 VDD.n929 76
R225 VDD.n923 VDD.n922 76
R226 VDD.n918 VDD.n917 76
R227 VDD.n913 VDD.n912 76
R228 VDD.n906 VDD.n905 76
R229 VDD.n901 VDD.n900 76
R230 VDD.n896 VDD.n895 76
R231 VDD.n892 VDD.n891 76
R232 VDD.n866 VDD.n865 76
R233 VDD.n862 VDD.n861 76
R234 VDD.n858 VDD.n857 76
R235 VDD.n854 VDD.n853 76
R236 VDD.n849 VDD.n848 76
R237 VDD.n842 VDD.n841 76
R238 VDD.n837 VDD.n836 76
R239 VDD.n832 VDD.n831 76
R240 VDD.n825 VDD.n824 76
R241 VDD.n820 VDD.n819 76
R242 VDD.n815 VDD.n814 76
R243 VDD.n811 VDD.n810 76
R244 VDD.n784 VDD.n783 76
R245 VDD.n780 VDD.n779 76
R246 VDD.n775 VDD.n774 76
R247 VDD.n770 VDD.n769 76
R248 VDD.n764 VDD.n763 76
R249 VDD.n759 VDD.n758 76
R250 VDD.n754 VDD.n753 76
R251 VDD.n749 VDD.n748 76
R252 VDD.n203 VDD.n202 64.064
R253 VDD.n406 VDD.n405 64.064
R254 VDD.n487 VDD.n486 64.064
R255 VDD.n629 VDD.n628 64.064
R256 VDD.n1358 VDD.n1357 64.064
R257 VDD.n1277 VDD.n1276 64.064
R258 VDD.n1135 VDD.n1134 64.064
R259 VDD.n932 VDD.n931 64.064
R260 VDD.n851 VDD.n850 64.064
R261 VDD.n232 VDD.n231 59.488
R262 VDD.n435 VDD.n434 59.488
R263 VDD.n516 VDD.n515 59.488
R264 VDD.n658 VDD.n657 59.488
R265 VDD.n1329 VDD.n1328 59.488
R266 VDD.n1248 VDD.n1247 59.488
R267 VDD.n1106 VDD.n1105 59.488
R268 VDD.n903 VDD.n902 59.488
R269 VDD.n822 VDD.n821 59.488
R270 VDD.n159 VDD.t31 55.465
R271 VDD.n133 VDD.t85 55.465
R272 VDD.n750 VDD.t1 55.106
R273 VDD.n816 VDD.t8 55.106
R274 VDD.n897 VDD.t53 55.106
R275 VDD.n974 VDD.t18 55.106
R276 VDD.n1035 VDD.t15 55.106
R277 VDD.n1100 VDD.t40 55.106
R278 VDD.n1177 VDD.t84 55.106
R279 VDD.n1242 VDD.t28 55.106
R280 VDD.n1323 VDD.t51 55.106
R281 VDD.n1400 VDD.t21 55.106
R282 VDD.n1461 VDD.t49 55.106
R283 VDD.n662 VDD.t69 55.106
R284 VDD.n585 VDD.t23 55.106
R285 VDD.n520 VDD.t30 55.106
R286 VDD.n439 VDD.t2 55.106
R287 VDD.n362 VDD.t0 55.106
R288 VDD.n301 VDD.t20 55.106
R289 VDD.n236 VDD.t76 55.106
R290 VDD.n857 VDD.t13 55.106
R291 VDD.n938 VDD.t14 55.106
R292 VDD.n1141 VDD.t88 55.106
R293 VDD.n1283 VDD.t78 55.106
R294 VDD.n1364 VDD.t79 55.106
R295 VDD.n626 VDD.t73 55.106
R296 VDD.n484 VDD.t36 55.106
R297 VDD.n403 VDD.t7 55.106
R298 VDD.n200 VDD.t90 55.106
R299 VDD.n776 VDD.t89 55.106
R300 VDD.n1000 VDD.t4 55.106
R301 VDD.n1061 VDD.t91 55.106
R302 VDD.n1203 VDD.t47 55.106
R303 VDD.n1426 VDD.t86 55.106
R304 VDD.n701 VDD.t33 55.106
R305 VDD.n559 VDD.t52 55.106
R306 VDD.n336 VDD.t5 55.106
R307 VDD.n275 VDD.t26 55.106
R308 VDD.n144 VDD.n143 41.183
R309 VDD.n766 VDD.n765 40.824
R310 VDD.n827 VDD.n826 40.824
R311 VDD.n847 VDD.n846 40.824
R312 VDD.n908 VDD.n907 40.824
R313 VDD.n928 VDD.n927 40.824
R314 VDD.n990 VDD.n989 40.824
R315 VDD.n1051 VDD.n1050 40.824
R316 VDD.n1111 VDD.n1110 40.824
R317 VDD.n1131 VDD.n1130 40.824
R318 VDD.n1193 VDD.n1192 40.824
R319 VDD.n1253 VDD.n1252 40.824
R320 VDD.n1273 VDD.n1272 40.824
R321 VDD.n1334 VDD.n1333 40.824
R322 VDD.n1354 VDD.n1353 40.824
R323 VDD.n1416 VDD.n1415 40.824
R324 VDD.n712 VDD.n711 40.824
R325 VDD.n651 VDD.n650 40.824
R326 VDD.n637 VDD.n636 40.824
R327 VDD.n570 VDD.n569 40.824
R328 VDD.n509 VDD.n508 40.824
R329 VDD.n495 VDD.n494 40.824
R330 VDD.n428 VDD.n427 40.824
R331 VDD.n414 VDD.n413 40.824
R332 VDD.n347 VDD.n346 40.824
R333 VDD.n286 VDD.n285 40.824
R334 VDD.n225 VDD.n224 40.824
R335 VDD.n211 VDD.n210 40.824
R336 VDD.n871 VDD.n870 36.774
R337 VDD.n952 VDD.n951 36.774
R338 VDD.n1013 VDD.n1012 36.774
R339 VDD.n1074 VDD.n1073 36.774
R340 VDD.n1155 VDD.n1154 36.774
R341 VDD.n1216 VDD.n1215 36.774
R342 VDD.n1297 VDD.n1296 36.774
R343 VDD.n1378 VDD.n1377 36.774
R344 VDD.n1439 VDD.n1438 36.774
R345 VDD.n679 VDD.n678 36.774
R346 VDD.n598 VDD.n597 36.774
R347 VDD.n537 VDD.n536 36.774
R348 VDD.n456 VDD.n455 36.774
R349 VDD.n375 VDD.n374 36.774
R350 VDD.n314 VDD.n313 36.774
R351 VDD.n253 VDD.n252 36.774
R352 VDD.n172 VDD.n171 36.774
R353 VDD.n111 VDD.n110 36.774
R354 VDD.n56 VDD.n55 36.774
R355 VDD.n800 VDD.n799 36.774
R356 VDD.n139 VDD.n138 36.608
R357 VDD.n281 VDD.n280 36.608
R358 VDD.n342 VDD.n341 36.608
R359 VDD.n565 VDD.n564 36.608
R360 VDD.n707 VDD.n706 36.608
R361 VDD.n1422 VDD.n1421 36.608
R362 VDD.n1199 VDD.n1198 36.608
R363 VDD.n1057 VDD.n1056 36.608
R364 VDD.n996 VDD.n995 36.608
R365 VDD.n772 VDD.n771 36.608
R366 VDD.n34 VDD.n33 34.942
R367 VDD.n155 VDD.n154 32.032
R368 VDD.n297 VDD.n296 32.032
R369 VDD.n358 VDD.n357 32.032
R370 VDD.n581 VDD.n580 32.032
R371 VDD.n723 VDD.n722 32.032
R372 VDD.n1406 VDD.n1405 32.032
R373 VDD.n1183 VDD.n1182 32.032
R374 VDD.n1041 VDD.n1040 32.032
R375 VDD.n980 VDD.n979 32.032
R376 VDD.n756 VDD.n755 32.032
R377 VDD.n208 VDD.n207 27.456
R378 VDD.n411 VDD.n410 27.456
R379 VDD.n492 VDD.n491 27.456
R380 VDD.n634 VDD.n633 27.456
R381 VDD.n1351 VDD.n1350 27.456
R382 VDD.n1270 VDD.n1269 27.456
R383 VDD.n1128 VDD.n1127 27.456
R384 VDD.n925 VDD.n924 27.456
R385 VDD.n844 VDD.n843 27.456
R386 VDD.n227 VDD.n226 22.88
R387 VDD.n430 VDD.n429 22.88
R388 VDD.n511 VDD.n510 22.88
R389 VDD.n653 VDD.n652 22.88
R390 VDD.n1336 VDD.n1335 22.88
R391 VDD.n1255 VDD.n1254 22.88
R392 VDD.n1113 VDD.n1112 22.88
R393 VDD.n910 VDD.n909 22.88
R394 VDD.n829 VDD.n828 22.88
R395 VDD.n748 VDD.n745 21.841
R396 VDD.n23 VDD.n20 21.841
R397 VDD.n765 VDD.t57 14.282
R398 VDD.n765 VDD.t22 14.282
R399 VDD.n826 VDD.t93 14.282
R400 VDD.n826 VDD.t37 14.282
R401 VDD.n846 VDD.t56 14.282
R402 VDD.n846 VDD.t41 14.282
R403 VDD.n907 VDD.t12 14.282
R404 VDD.n907 VDD.t62 14.282
R405 VDD.n927 VDD.t45 14.282
R406 VDD.n927 VDD.t63 14.282
R407 VDD.n989 VDD.t3 14.282
R408 VDD.n989 VDD.t60 14.282
R409 VDD.n1050 VDD.t50 14.282
R410 VDD.n1050 VDD.t46 14.282
R411 VDD.n1110 VDD.t65 14.282
R412 VDD.n1110 VDD.t43 14.282
R413 VDD.n1130 VDD.t55 14.282
R414 VDD.n1130 VDD.t66 14.282
R415 VDD.n1192 VDD.t17 14.282
R416 VDD.n1192 VDD.t9 14.282
R417 VDD.n1252 VDD.t92 14.282
R418 VDD.n1252 VDD.t48 14.282
R419 VDD.n1272 VDD.t81 14.282
R420 VDD.n1272 VDD.t42 14.282
R421 VDD.n1333 VDD.t35 14.282
R422 VDD.n1333 VDD.t24 14.282
R423 VDD.n1353 VDD.t82 14.282
R424 VDD.n1353 VDD.t27 14.282
R425 VDD.n1415 VDD.t6 14.282
R426 VDD.n1415 VDD.t54 14.282
R427 VDD.n711 VDD.t34 14.282
R428 VDD.n711 VDD.t59 14.282
R429 VDD.n650 VDD.t72 14.282
R430 VDD.n650 VDD.t64 14.282
R431 VDD.n636 VDD.t80 14.282
R432 VDD.n636 VDD.t10 14.282
R433 VDD.n569 VDD.t87 14.282
R434 VDD.n569 VDD.t11 14.282
R435 VDD.n508 VDD.t61 14.282
R436 VDD.n508 VDD.t44 14.282
R437 VDD.n494 VDD.t58 14.282
R438 VDD.n494 VDD.t75 14.282
R439 VDD.n427 VDD.t71 14.282
R440 VDD.n427 VDD.t38 14.282
R441 VDD.n413 VDD.t16 14.282
R442 VDD.n413 VDD.t70 14.282
R443 VDD.n346 VDD.t83 14.282
R444 VDD.n346 VDD.t29 14.282
R445 VDD.n285 VDD.t74 14.282
R446 VDD.n285 VDD.t19 14.282
R447 VDD.n224 VDD.t25 14.282
R448 VDD.n224 VDD.t77 14.282
R449 VDD.n210 VDD.t39 14.282
R450 VDD.n210 VDD.t68 14.282
R451 VDD.n143 VDD.t67 14.282
R452 VDD.n143 VDD.t32 14.282
R453 VDD.n745 VDD.n728 14.167
R454 VDD.n728 VDD.n727 14.167
R455 VDD.n886 VDD.n868 14.167
R456 VDD.n868 VDD.n867 14.167
R457 VDD.n967 VDD.n949 14.167
R458 VDD.n949 VDD.n948 14.167
R459 VDD.n1028 VDD.n1010 14.167
R460 VDD.n1010 VDD.n1009 14.167
R461 VDD.n1089 VDD.n1071 14.167
R462 VDD.n1071 VDD.n1070 14.167
R463 VDD.n1170 VDD.n1152 14.167
R464 VDD.n1152 VDD.n1151 14.167
R465 VDD.n1231 VDD.n1213 14.167
R466 VDD.n1213 VDD.n1212 14.167
R467 VDD.n1312 VDD.n1294 14.167
R468 VDD.n1294 VDD.n1293 14.167
R469 VDD.n1393 VDD.n1375 14.167
R470 VDD.n1375 VDD.n1374 14.167
R471 VDD.n1454 VDD.n1436 14.167
R472 VDD.n1436 VDD.n1435 14.167
R473 VDD.n694 VDD.n676 14.167
R474 VDD.n676 VDD.n675 14.167
R475 VDD.n613 VDD.n595 14.167
R476 VDD.n595 VDD.n594 14.167
R477 VDD.n552 VDD.n534 14.167
R478 VDD.n534 VDD.n533 14.167
R479 VDD.n471 VDD.n453 14.167
R480 VDD.n453 VDD.n452 14.167
R481 VDD.n390 VDD.n372 14.167
R482 VDD.n372 VDD.n371 14.167
R483 VDD.n329 VDD.n311 14.167
R484 VDD.n311 VDD.n310 14.167
R485 VDD.n268 VDD.n250 14.167
R486 VDD.n250 VDD.n249 14.167
R487 VDD.n187 VDD.n169 14.167
R488 VDD.n169 VDD.n168 14.167
R489 VDD.n126 VDD.n108 14.167
R490 VDD.n108 VDD.n107 14.167
R491 VDD.n72 VDD.n53 14.167
R492 VDD.n53 VDD.n52 14.167
R493 VDD.n805 VDD.n786 14.167
R494 VDD.n786 VDD.n785 14.167
R495 VDD.n20 VDD.n19 14.167
R496 VDD.n19 VDD.n17 14.167
R497 VDD.n32 VDD.n29 14.167
R498 VDD.n29 VDD.n28 14.167
R499 VDD.n77 VDD.n73 14.167
R500 VDD.n131 VDD.n127 14.167
R501 VDD.n192 VDD.n188 14.167
R502 VDD.n273 VDD.n269 14.167
R503 VDD.n334 VDD.n330 14.167
R504 VDD.n395 VDD.n391 14.167
R505 VDD.n476 VDD.n472 14.167
R506 VDD.n557 VDD.n553 14.167
R507 VDD.n618 VDD.n614 14.167
R508 VDD.n699 VDD.n695 14.167
R509 VDD.n1459 VDD.n1455 14.167
R510 VDD.n1398 VDD.n1394 14.167
R511 VDD.n1317 VDD.n1313 14.167
R512 VDD.n1236 VDD.n1232 14.167
R513 VDD.n1175 VDD.n1171 14.167
R514 VDD.n1094 VDD.n1090 14.167
R515 VDD.n1033 VDD.n1029 14.167
R516 VDD.n972 VDD.n968 14.167
R517 VDD.n891 VDD.n887 14.167
R518 VDD.n810 VDD.n806 14.167
R519 VDD.n220 VDD.n219 13.728
R520 VDD.n423 VDD.n422 13.728
R521 VDD.n504 VDD.n503 13.728
R522 VDD.n646 VDD.n645 13.728
R523 VDD.n1341 VDD.n1340 13.728
R524 VDD.n1260 VDD.n1259 13.728
R525 VDD.n1118 VDD.n1117 13.728
R526 VDD.n915 VDD.n914 13.728
R527 VDD.n834 VDD.n833 13.728
R528 VDD.n23 VDD.n22 13.653
R529 VDD.n22 VDD.n21 13.653
R530 VDD.n32 VDD.n31 13.653
R531 VDD.n31 VDD.n30 13.653
R532 VDD.n29 VDD.n25 13.653
R533 VDD.n25 VDD.n24 13.653
R534 VDD.n28 VDD.n27 13.653
R535 VDD.n27 VDD.n26 13.653
R536 VDD.n38 VDD.n37 13.653
R537 VDD.n37 VDD.n36 13.653
R538 VDD.n42 VDD.n41 13.653
R539 VDD.n41 VDD.n40 13.653
R540 VDD.n46 VDD.n45 13.653
R541 VDD.n45 VDD.n44 13.653
R542 VDD.n50 VDD.n49 13.653
R543 VDD.n49 VDD.n48 13.653
R544 VDD.n77 VDD.n76 13.653
R545 VDD.n76 VDD.n75 13.653
R546 VDD.n81 VDD.n80 13.653
R547 VDD.n80 VDD.n79 13.653
R548 VDD.n85 VDD.n84 13.653
R549 VDD.n84 VDD.n83 13.653
R550 VDD.n89 VDD.n88 13.653
R551 VDD.n88 VDD.n87 13.653
R552 VDD.n93 VDD.n92 13.653
R553 VDD.n92 VDD.n91 13.653
R554 VDD.n97 VDD.n96 13.653
R555 VDD.n96 VDD.n95 13.653
R556 VDD.n101 VDD.n100 13.653
R557 VDD.n100 VDD.n99 13.653
R558 VDD.n105 VDD.n104 13.653
R559 VDD.n104 VDD.n103 13.653
R560 VDD.n131 VDD.n130 13.653
R561 VDD.n130 VDD.n129 13.653
R562 VDD.n136 VDD.n135 13.653
R563 VDD.n135 VDD.n134 13.653
R564 VDD.n141 VDD.n140 13.653
R565 VDD.n140 VDD.n139 13.653
R566 VDD.n147 VDD.n146 13.653
R567 VDD.n146 VDD.n145 13.653
R568 VDD.n152 VDD.n151 13.653
R569 VDD.n151 VDD.n150 13.653
R570 VDD.n157 VDD.n156 13.653
R571 VDD.n156 VDD.n155 13.653
R572 VDD.n162 VDD.n161 13.653
R573 VDD.n161 VDD.n160 13.653
R574 VDD.n166 VDD.n165 13.653
R575 VDD.n165 VDD.n164 13.653
R576 VDD.n192 VDD.n191 13.653
R577 VDD.n191 VDD.n190 13.653
R578 VDD.n196 VDD.n195 13.653
R579 VDD.n195 VDD.n194 13.653
R580 VDD.n200 VDD.n199 13.653
R581 VDD.n199 VDD.n198 13.653
R582 VDD.n205 VDD.n204 13.653
R583 VDD.n204 VDD.n203 13.653
R584 VDD.n212 VDD.n209 13.653
R585 VDD.n209 VDD.n208 13.653
R586 VDD.n217 VDD.n216 13.653
R587 VDD.n216 VDD.n215 13.653
R588 VDD.n222 VDD.n221 13.653
R589 VDD.n221 VDD.n220 13.653
R590 VDD.n229 VDD.n228 13.653
R591 VDD.n228 VDD.n227 13.653
R592 VDD.n234 VDD.n233 13.653
R593 VDD.n233 VDD.n232 13.653
R594 VDD.n239 VDD.n238 13.653
R595 VDD.n238 VDD.n237 13.653
R596 VDD.n243 VDD.n242 13.653
R597 VDD.n242 VDD.n241 13.653
R598 VDD.n247 VDD.n246 13.653
R599 VDD.n246 VDD.n245 13.653
R600 VDD.n273 VDD.n272 13.653
R601 VDD.n272 VDD.n271 13.653
R602 VDD.n278 VDD.n277 13.653
R603 VDD.n277 VDD.n276 13.653
R604 VDD.n283 VDD.n282 13.653
R605 VDD.n282 VDD.n281 13.653
R606 VDD.n289 VDD.n288 13.653
R607 VDD.n288 VDD.n287 13.653
R608 VDD.n294 VDD.n293 13.653
R609 VDD.n293 VDD.n292 13.653
R610 VDD.n299 VDD.n298 13.653
R611 VDD.n298 VDD.n297 13.653
R612 VDD.n304 VDD.n303 13.653
R613 VDD.n303 VDD.n302 13.653
R614 VDD.n308 VDD.n307 13.653
R615 VDD.n307 VDD.n306 13.653
R616 VDD.n334 VDD.n333 13.653
R617 VDD.n333 VDD.n332 13.653
R618 VDD.n339 VDD.n338 13.653
R619 VDD.n338 VDD.n337 13.653
R620 VDD.n344 VDD.n343 13.653
R621 VDD.n343 VDD.n342 13.653
R622 VDD.n350 VDD.n349 13.653
R623 VDD.n349 VDD.n348 13.653
R624 VDD.n355 VDD.n354 13.653
R625 VDD.n354 VDD.n353 13.653
R626 VDD.n360 VDD.n359 13.653
R627 VDD.n359 VDD.n358 13.653
R628 VDD.n365 VDD.n364 13.653
R629 VDD.n364 VDD.n363 13.653
R630 VDD.n369 VDD.n368 13.653
R631 VDD.n368 VDD.n367 13.653
R632 VDD.n395 VDD.n394 13.653
R633 VDD.n394 VDD.n393 13.653
R634 VDD.n399 VDD.n398 13.653
R635 VDD.n398 VDD.n397 13.653
R636 VDD.n403 VDD.n402 13.653
R637 VDD.n402 VDD.n401 13.653
R638 VDD.n408 VDD.n407 13.653
R639 VDD.n407 VDD.n406 13.653
R640 VDD.n415 VDD.n412 13.653
R641 VDD.n412 VDD.n411 13.653
R642 VDD.n420 VDD.n419 13.653
R643 VDD.n419 VDD.n418 13.653
R644 VDD.n425 VDD.n424 13.653
R645 VDD.n424 VDD.n423 13.653
R646 VDD.n432 VDD.n431 13.653
R647 VDD.n431 VDD.n430 13.653
R648 VDD.n437 VDD.n436 13.653
R649 VDD.n436 VDD.n435 13.653
R650 VDD.n442 VDD.n441 13.653
R651 VDD.n441 VDD.n440 13.653
R652 VDD.n446 VDD.n445 13.653
R653 VDD.n445 VDD.n444 13.653
R654 VDD.n450 VDD.n449 13.653
R655 VDD.n449 VDD.n448 13.653
R656 VDD.n476 VDD.n475 13.653
R657 VDD.n475 VDD.n474 13.653
R658 VDD.n480 VDD.n479 13.653
R659 VDD.n479 VDD.n478 13.653
R660 VDD.n484 VDD.n483 13.653
R661 VDD.n483 VDD.n482 13.653
R662 VDD.n489 VDD.n488 13.653
R663 VDD.n488 VDD.n487 13.653
R664 VDD.n496 VDD.n493 13.653
R665 VDD.n493 VDD.n492 13.653
R666 VDD.n501 VDD.n500 13.653
R667 VDD.n500 VDD.n499 13.653
R668 VDD.n506 VDD.n505 13.653
R669 VDD.n505 VDD.n504 13.653
R670 VDD.n513 VDD.n512 13.653
R671 VDD.n512 VDD.n511 13.653
R672 VDD.n518 VDD.n517 13.653
R673 VDD.n517 VDD.n516 13.653
R674 VDD.n523 VDD.n522 13.653
R675 VDD.n522 VDD.n521 13.653
R676 VDD.n527 VDD.n526 13.653
R677 VDD.n526 VDD.n525 13.653
R678 VDD.n531 VDD.n530 13.653
R679 VDD.n530 VDD.n529 13.653
R680 VDD.n557 VDD.n556 13.653
R681 VDD.n556 VDD.n555 13.653
R682 VDD.n562 VDD.n561 13.653
R683 VDD.n561 VDD.n560 13.653
R684 VDD.n567 VDD.n566 13.653
R685 VDD.n566 VDD.n565 13.653
R686 VDD.n573 VDD.n572 13.653
R687 VDD.n572 VDD.n571 13.653
R688 VDD.n578 VDD.n577 13.653
R689 VDD.n577 VDD.n576 13.653
R690 VDD.n583 VDD.n582 13.653
R691 VDD.n582 VDD.n581 13.653
R692 VDD.n588 VDD.n587 13.653
R693 VDD.n587 VDD.n586 13.653
R694 VDD.n592 VDD.n591 13.653
R695 VDD.n591 VDD.n590 13.653
R696 VDD.n618 VDD.n617 13.653
R697 VDD.n617 VDD.n616 13.653
R698 VDD.n622 VDD.n621 13.653
R699 VDD.n621 VDD.n620 13.653
R700 VDD.n626 VDD.n625 13.653
R701 VDD.n625 VDD.n624 13.653
R702 VDD.n631 VDD.n630 13.653
R703 VDD.n630 VDD.n629 13.653
R704 VDD.n638 VDD.n635 13.653
R705 VDD.n635 VDD.n634 13.653
R706 VDD.n643 VDD.n642 13.653
R707 VDD.n642 VDD.n641 13.653
R708 VDD.n648 VDD.n647 13.653
R709 VDD.n647 VDD.n646 13.653
R710 VDD.n655 VDD.n654 13.653
R711 VDD.n654 VDD.n653 13.653
R712 VDD.n660 VDD.n659 13.653
R713 VDD.n659 VDD.n658 13.653
R714 VDD.n665 VDD.n664 13.653
R715 VDD.n664 VDD.n663 13.653
R716 VDD.n669 VDD.n668 13.653
R717 VDD.n668 VDD.n667 13.653
R718 VDD.n673 VDD.n672 13.653
R719 VDD.n672 VDD.n671 13.653
R720 VDD.n699 VDD.n698 13.653
R721 VDD.n698 VDD.n697 13.653
R722 VDD.n704 VDD.n703 13.653
R723 VDD.n703 VDD.n702 13.653
R724 VDD.n709 VDD.n708 13.653
R725 VDD.n708 VDD.n707 13.653
R726 VDD.n715 VDD.n714 13.653
R727 VDD.n714 VDD.n713 13.653
R728 VDD.n720 VDD.n719 13.653
R729 VDD.n719 VDD.n718 13.653
R730 VDD.n725 VDD.n724 13.653
R731 VDD.n724 VDD.n723 13.653
R732 VDD.n1464 VDD.n1463 13.653
R733 VDD.n1463 VDD.n1462 13.653
R734 VDD.n1459 VDD.n1458 13.653
R735 VDD.n1458 VDD.n1457 13.653
R736 VDD.n1433 VDD.n1432 13.653
R737 VDD.n1432 VDD.n1431 13.653
R738 VDD.n1429 VDD.n1428 13.653
R739 VDD.n1428 VDD.n1427 13.653
R740 VDD.n1424 VDD.n1423 13.653
R741 VDD.n1423 VDD.n1422 13.653
R742 VDD.n1419 VDD.n1418 13.653
R743 VDD.n1418 VDD.n1417 13.653
R744 VDD.n1413 VDD.n1412 13.653
R745 VDD.n1412 VDD.n1411 13.653
R746 VDD.n1408 VDD.n1407 13.653
R747 VDD.n1407 VDD.n1406 13.653
R748 VDD.n1403 VDD.n1402 13.653
R749 VDD.n1402 VDD.n1401 13.653
R750 VDD.n1398 VDD.n1397 13.653
R751 VDD.n1397 VDD.n1396 13.653
R752 VDD.n1372 VDD.n1371 13.653
R753 VDD.n1371 VDD.n1370 13.653
R754 VDD.n1368 VDD.n1367 13.653
R755 VDD.n1367 VDD.n1366 13.653
R756 VDD.n1364 VDD.n1363 13.653
R757 VDD.n1363 VDD.n1362 13.653
R758 VDD.n1360 VDD.n1359 13.653
R759 VDD.n1359 VDD.n1358 13.653
R760 VDD.n1355 VDD.n1352 13.653
R761 VDD.n1352 VDD.n1351 13.653
R762 VDD.n1348 VDD.n1347 13.653
R763 VDD.n1347 VDD.n1346 13.653
R764 VDD.n1343 VDD.n1342 13.653
R765 VDD.n1342 VDD.n1341 13.653
R766 VDD.n1338 VDD.n1337 13.653
R767 VDD.n1337 VDD.n1336 13.653
R768 VDD.n1331 VDD.n1330 13.653
R769 VDD.n1330 VDD.n1329 13.653
R770 VDD.n1326 VDD.n1325 13.653
R771 VDD.n1325 VDD.n1324 13.653
R772 VDD.n1321 VDD.n1320 13.653
R773 VDD.n1320 VDD.n1319 13.653
R774 VDD.n1317 VDD.n1316 13.653
R775 VDD.n1316 VDD.n1315 13.653
R776 VDD.n1291 VDD.n1290 13.653
R777 VDD.n1290 VDD.n1289 13.653
R778 VDD.n1287 VDD.n1286 13.653
R779 VDD.n1286 VDD.n1285 13.653
R780 VDD.n1283 VDD.n1282 13.653
R781 VDD.n1282 VDD.n1281 13.653
R782 VDD.n1279 VDD.n1278 13.653
R783 VDD.n1278 VDD.n1277 13.653
R784 VDD.n1274 VDD.n1271 13.653
R785 VDD.n1271 VDD.n1270 13.653
R786 VDD.n1267 VDD.n1266 13.653
R787 VDD.n1266 VDD.n1265 13.653
R788 VDD.n1262 VDD.n1261 13.653
R789 VDD.n1261 VDD.n1260 13.653
R790 VDD.n1257 VDD.n1256 13.653
R791 VDD.n1256 VDD.n1255 13.653
R792 VDD.n1250 VDD.n1249 13.653
R793 VDD.n1249 VDD.n1248 13.653
R794 VDD.n1245 VDD.n1244 13.653
R795 VDD.n1244 VDD.n1243 13.653
R796 VDD.n1240 VDD.n1239 13.653
R797 VDD.n1239 VDD.n1238 13.653
R798 VDD.n1236 VDD.n1235 13.653
R799 VDD.n1235 VDD.n1234 13.653
R800 VDD.n1210 VDD.n1209 13.653
R801 VDD.n1209 VDD.n1208 13.653
R802 VDD.n1206 VDD.n1205 13.653
R803 VDD.n1205 VDD.n1204 13.653
R804 VDD.n1201 VDD.n1200 13.653
R805 VDD.n1200 VDD.n1199 13.653
R806 VDD.n1196 VDD.n1195 13.653
R807 VDD.n1195 VDD.n1194 13.653
R808 VDD.n1190 VDD.n1189 13.653
R809 VDD.n1189 VDD.n1188 13.653
R810 VDD.n1185 VDD.n1184 13.653
R811 VDD.n1184 VDD.n1183 13.653
R812 VDD.n1180 VDD.n1179 13.653
R813 VDD.n1179 VDD.n1178 13.653
R814 VDD.n1175 VDD.n1174 13.653
R815 VDD.n1174 VDD.n1173 13.653
R816 VDD.n1149 VDD.n1148 13.653
R817 VDD.n1148 VDD.n1147 13.653
R818 VDD.n1145 VDD.n1144 13.653
R819 VDD.n1144 VDD.n1143 13.653
R820 VDD.n1141 VDD.n1140 13.653
R821 VDD.n1140 VDD.n1139 13.653
R822 VDD.n1137 VDD.n1136 13.653
R823 VDD.n1136 VDD.n1135 13.653
R824 VDD.n1132 VDD.n1129 13.653
R825 VDD.n1129 VDD.n1128 13.653
R826 VDD.n1125 VDD.n1124 13.653
R827 VDD.n1124 VDD.n1123 13.653
R828 VDD.n1120 VDD.n1119 13.653
R829 VDD.n1119 VDD.n1118 13.653
R830 VDD.n1115 VDD.n1114 13.653
R831 VDD.n1114 VDD.n1113 13.653
R832 VDD.n1108 VDD.n1107 13.653
R833 VDD.n1107 VDD.n1106 13.653
R834 VDD.n1103 VDD.n1102 13.653
R835 VDD.n1102 VDD.n1101 13.653
R836 VDD.n1098 VDD.n1097 13.653
R837 VDD.n1097 VDD.n1096 13.653
R838 VDD.n1094 VDD.n1093 13.653
R839 VDD.n1093 VDD.n1092 13.653
R840 VDD.n1068 VDD.n1067 13.653
R841 VDD.n1067 VDD.n1066 13.653
R842 VDD.n1064 VDD.n1063 13.653
R843 VDD.n1063 VDD.n1062 13.653
R844 VDD.n1059 VDD.n1058 13.653
R845 VDD.n1058 VDD.n1057 13.653
R846 VDD.n1054 VDD.n1053 13.653
R847 VDD.n1053 VDD.n1052 13.653
R848 VDD.n1048 VDD.n1047 13.653
R849 VDD.n1047 VDD.n1046 13.653
R850 VDD.n1043 VDD.n1042 13.653
R851 VDD.n1042 VDD.n1041 13.653
R852 VDD.n1038 VDD.n1037 13.653
R853 VDD.n1037 VDD.n1036 13.653
R854 VDD.n1033 VDD.n1032 13.653
R855 VDD.n1032 VDD.n1031 13.653
R856 VDD.n1007 VDD.n1006 13.653
R857 VDD.n1006 VDD.n1005 13.653
R858 VDD.n1003 VDD.n1002 13.653
R859 VDD.n1002 VDD.n1001 13.653
R860 VDD.n998 VDD.n997 13.653
R861 VDD.n997 VDD.n996 13.653
R862 VDD.n993 VDD.n992 13.653
R863 VDD.n992 VDD.n991 13.653
R864 VDD.n987 VDD.n986 13.653
R865 VDD.n986 VDD.n985 13.653
R866 VDD.n982 VDD.n981 13.653
R867 VDD.n981 VDD.n980 13.653
R868 VDD.n977 VDD.n976 13.653
R869 VDD.n976 VDD.n975 13.653
R870 VDD.n972 VDD.n971 13.653
R871 VDD.n971 VDD.n970 13.653
R872 VDD.n946 VDD.n945 13.653
R873 VDD.n945 VDD.n944 13.653
R874 VDD.n942 VDD.n941 13.653
R875 VDD.n941 VDD.n940 13.653
R876 VDD.n938 VDD.n937 13.653
R877 VDD.n937 VDD.n936 13.653
R878 VDD.n934 VDD.n933 13.653
R879 VDD.n933 VDD.n932 13.653
R880 VDD.n929 VDD.n926 13.653
R881 VDD.n926 VDD.n925 13.653
R882 VDD.n922 VDD.n921 13.653
R883 VDD.n921 VDD.n920 13.653
R884 VDD.n917 VDD.n916 13.653
R885 VDD.n916 VDD.n915 13.653
R886 VDD.n912 VDD.n911 13.653
R887 VDD.n911 VDD.n910 13.653
R888 VDD.n905 VDD.n904 13.653
R889 VDD.n904 VDD.n903 13.653
R890 VDD.n900 VDD.n899 13.653
R891 VDD.n899 VDD.n898 13.653
R892 VDD.n895 VDD.n894 13.653
R893 VDD.n894 VDD.n893 13.653
R894 VDD.n891 VDD.n890 13.653
R895 VDD.n890 VDD.n889 13.653
R896 VDD.n865 VDD.n864 13.653
R897 VDD.n864 VDD.n863 13.653
R898 VDD.n861 VDD.n860 13.653
R899 VDD.n860 VDD.n859 13.653
R900 VDD.n857 VDD.n856 13.653
R901 VDD.n856 VDD.n855 13.653
R902 VDD.n853 VDD.n852 13.653
R903 VDD.n852 VDD.n851 13.653
R904 VDD.n848 VDD.n845 13.653
R905 VDD.n845 VDD.n844 13.653
R906 VDD.n841 VDD.n840 13.653
R907 VDD.n840 VDD.n839 13.653
R908 VDD.n836 VDD.n835 13.653
R909 VDD.n835 VDD.n834 13.653
R910 VDD.n831 VDD.n830 13.653
R911 VDD.n830 VDD.n829 13.653
R912 VDD.n824 VDD.n823 13.653
R913 VDD.n823 VDD.n822 13.653
R914 VDD.n819 VDD.n818 13.653
R915 VDD.n818 VDD.n817 13.653
R916 VDD.n814 VDD.n813 13.653
R917 VDD.n813 VDD.n812 13.653
R918 VDD.n810 VDD.n809 13.653
R919 VDD.n809 VDD.n808 13.653
R920 VDD.n783 VDD.n782 13.653
R921 VDD.n782 VDD.n781 13.653
R922 VDD.n779 VDD.n778 13.653
R923 VDD.n778 VDD.n777 13.653
R924 VDD.n774 VDD.n773 13.653
R925 VDD.n773 VDD.n772 13.653
R926 VDD.n769 VDD.n768 13.653
R927 VDD.n768 VDD.n767 13.653
R928 VDD.n763 VDD.n762 13.653
R929 VDD.n762 VDD.n761 13.653
R930 VDD.n758 VDD.n757 13.653
R931 VDD.n757 VDD.n756 13.653
R932 VDD.n753 VDD.n752 13.653
R933 VDD.n752 VDD.n751 13.653
R934 VDD.n748 VDD.n747 13.653
R935 VDD.n747 VDD.n746 13.653
R936 VDD.n4 VDD.n2 12.915
R937 VDD.n4 VDD.n3 12.66
R938 VDD.n13 VDD.n12 12.343
R939 VDD.n11 VDD.n10 12.343
R940 VDD.n7 VDD.n6 12.343
R941 VDD.n215 VDD.n214 9.152
R942 VDD.n418 VDD.n417 9.152
R943 VDD.n499 VDD.n498 9.152
R944 VDD.n641 VDD.n640 9.152
R945 VDD.n1346 VDD.n1345 9.152
R946 VDD.n1265 VDD.n1264 9.152
R947 VDD.n1123 VDD.n1122 9.152
R948 VDD.n920 VDD.n919 9.152
R949 VDD.n839 VDD.n838 9.152
R950 VDD.n147 VDD.n144 8.658
R951 VDD.n289 VDD.n286 8.658
R952 VDD.n350 VDD.n347 8.658
R953 VDD.n573 VDD.n570 8.658
R954 VDD.n715 VDD.n712 8.658
R955 VDD.n1419 VDD.n1416 8.658
R956 VDD.n1196 VDD.n1193 8.658
R957 VDD.n1054 VDD.n1051 8.658
R958 VDD.n993 VDD.n990 8.658
R959 VDD.n769 VDD.n766 8.658
R960 VDD.n887 VDD.n886 7.674
R961 VDD.n968 VDD.n967 7.674
R962 VDD.n1029 VDD.n1028 7.674
R963 VDD.n1090 VDD.n1089 7.674
R964 VDD.n1171 VDD.n1170 7.674
R965 VDD.n1232 VDD.n1231 7.674
R966 VDD.n1313 VDD.n1312 7.674
R967 VDD.n1394 VDD.n1393 7.674
R968 VDD.n1455 VDD.n1454 7.674
R969 VDD.n695 VDD.n694 7.674
R970 VDD.n614 VDD.n613 7.674
R971 VDD.n553 VDD.n552 7.674
R972 VDD.n472 VDD.n471 7.674
R973 VDD.n391 VDD.n390 7.674
R974 VDD.n330 VDD.n329 7.674
R975 VDD.n269 VDD.n268 7.674
R976 VDD.n188 VDD.n187 7.674
R977 VDD.n127 VDD.n126 7.674
R978 VDD.n73 VDD.n72 7.674
R979 VDD.n806 VDD.n805 7.674
R980 VDD.n67 VDD.n66 7.5
R981 VDD.n61 VDD.n60 7.5
R982 VDD.n63 VDD.n62 7.5
R983 VDD.n58 VDD.n57 7.5
R984 VDD.n72 VDD.n71 7.5
R985 VDD.n121 VDD.n120 7.5
R986 VDD.n115 VDD.n114 7.5
R987 VDD.n117 VDD.n116 7.5
R988 VDD.n123 VDD.n113 7.5
R989 VDD.n123 VDD.n111 7.5
R990 VDD.n126 VDD.n125 7.5
R991 VDD.n182 VDD.n181 7.5
R992 VDD.n176 VDD.n175 7.5
R993 VDD.n178 VDD.n177 7.5
R994 VDD.n184 VDD.n174 7.5
R995 VDD.n184 VDD.n172 7.5
R996 VDD.n187 VDD.n186 7.5
R997 VDD.n263 VDD.n262 7.5
R998 VDD.n257 VDD.n256 7.5
R999 VDD.n259 VDD.n258 7.5
R1000 VDD.n265 VDD.n255 7.5
R1001 VDD.n265 VDD.n253 7.5
R1002 VDD.n268 VDD.n267 7.5
R1003 VDD.n324 VDD.n323 7.5
R1004 VDD.n318 VDD.n317 7.5
R1005 VDD.n320 VDD.n319 7.5
R1006 VDD.n326 VDD.n316 7.5
R1007 VDD.n326 VDD.n314 7.5
R1008 VDD.n329 VDD.n328 7.5
R1009 VDD.n385 VDD.n384 7.5
R1010 VDD.n379 VDD.n378 7.5
R1011 VDD.n381 VDD.n380 7.5
R1012 VDD.n387 VDD.n377 7.5
R1013 VDD.n387 VDD.n375 7.5
R1014 VDD.n390 VDD.n389 7.5
R1015 VDD.n466 VDD.n465 7.5
R1016 VDD.n460 VDD.n459 7.5
R1017 VDD.n462 VDD.n461 7.5
R1018 VDD.n468 VDD.n458 7.5
R1019 VDD.n468 VDD.n456 7.5
R1020 VDD.n471 VDD.n470 7.5
R1021 VDD.n547 VDD.n546 7.5
R1022 VDD.n541 VDD.n540 7.5
R1023 VDD.n543 VDD.n542 7.5
R1024 VDD.n549 VDD.n539 7.5
R1025 VDD.n549 VDD.n537 7.5
R1026 VDD.n552 VDD.n551 7.5
R1027 VDD.n608 VDD.n607 7.5
R1028 VDD.n602 VDD.n601 7.5
R1029 VDD.n604 VDD.n603 7.5
R1030 VDD.n610 VDD.n600 7.5
R1031 VDD.n610 VDD.n598 7.5
R1032 VDD.n613 VDD.n612 7.5
R1033 VDD.n689 VDD.n688 7.5
R1034 VDD.n683 VDD.n682 7.5
R1035 VDD.n685 VDD.n684 7.5
R1036 VDD.n691 VDD.n681 7.5
R1037 VDD.n691 VDD.n679 7.5
R1038 VDD.n694 VDD.n693 7.5
R1039 VDD.n1449 VDD.n1448 7.5
R1040 VDD.n1443 VDD.n1442 7.5
R1041 VDD.n1445 VDD.n1444 7.5
R1042 VDD.n1451 VDD.n1441 7.5
R1043 VDD.n1451 VDD.n1439 7.5
R1044 VDD.n1454 VDD.n1453 7.5
R1045 VDD.n1388 VDD.n1387 7.5
R1046 VDD.n1382 VDD.n1381 7.5
R1047 VDD.n1384 VDD.n1383 7.5
R1048 VDD.n1390 VDD.n1380 7.5
R1049 VDD.n1390 VDD.n1378 7.5
R1050 VDD.n1393 VDD.n1392 7.5
R1051 VDD.n1307 VDD.n1306 7.5
R1052 VDD.n1301 VDD.n1300 7.5
R1053 VDD.n1303 VDD.n1302 7.5
R1054 VDD.n1309 VDD.n1299 7.5
R1055 VDD.n1309 VDD.n1297 7.5
R1056 VDD.n1312 VDD.n1311 7.5
R1057 VDD.n1226 VDD.n1225 7.5
R1058 VDD.n1220 VDD.n1219 7.5
R1059 VDD.n1222 VDD.n1221 7.5
R1060 VDD.n1228 VDD.n1218 7.5
R1061 VDD.n1228 VDD.n1216 7.5
R1062 VDD.n1231 VDD.n1230 7.5
R1063 VDD.n1165 VDD.n1164 7.5
R1064 VDD.n1159 VDD.n1158 7.5
R1065 VDD.n1161 VDD.n1160 7.5
R1066 VDD.n1167 VDD.n1157 7.5
R1067 VDD.n1167 VDD.n1155 7.5
R1068 VDD.n1170 VDD.n1169 7.5
R1069 VDD.n1084 VDD.n1083 7.5
R1070 VDD.n1078 VDD.n1077 7.5
R1071 VDD.n1080 VDD.n1079 7.5
R1072 VDD.n1086 VDD.n1076 7.5
R1073 VDD.n1086 VDD.n1074 7.5
R1074 VDD.n1089 VDD.n1088 7.5
R1075 VDD.n1023 VDD.n1022 7.5
R1076 VDD.n1017 VDD.n1016 7.5
R1077 VDD.n1019 VDD.n1018 7.5
R1078 VDD.n1025 VDD.n1015 7.5
R1079 VDD.n1025 VDD.n1013 7.5
R1080 VDD.n1028 VDD.n1027 7.5
R1081 VDD.n962 VDD.n961 7.5
R1082 VDD.n956 VDD.n955 7.5
R1083 VDD.n958 VDD.n957 7.5
R1084 VDD.n964 VDD.n954 7.5
R1085 VDD.n964 VDD.n952 7.5
R1086 VDD.n967 VDD.n966 7.5
R1087 VDD.n881 VDD.n880 7.5
R1088 VDD.n875 VDD.n874 7.5
R1089 VDD.n877 VDD.n876 7.5
R1090 VDD.n883 VDD.n873 7.5
R1091 VDD.n883 VDD.n871 7.5
R1092 VDD.n886 VDD.n885 7.5
R1093 VDD.n790 VDD.n789 7.5
R1094 VDD.n793 VDD.n792 7.5
R1095 VDD.n795 VDD.n794 7.5
R1096 VDD.n798 VDD.n797 7.5
R1097 VDD.n805 VDD.n804 7.5
R1098 VDD.n740 VDD.n739 7.5
R1099 VDD.n734 VDD.n733 7.5
R1100 VDD.n736 VDD.n735 7.5
R1101 VDD.n742 VDD.n732 7.5
R1102 VDD.n742 VDD.n730 7.5
R1103 VDD.n745 VDD.n744 7.5
R1104 VDD.n20 VDD.n16 7.5
R1105 VDD.n2 VDD.n1 7.5
R1106 VDD.n6 VDD.n5 7.5
R1107 VDD.n10 VDD.n9 7.5
R1108 VDD.n19 VDD.n18 7.5
R1109 VDD.n14 VDD.n0 7.5
R1110 VDD.n59 VDD.n56 6.772
R1111 VDD.n70 VDD.n54 6.772
R1112 VDD.n68 VDD.n65 6.772
R1113 VDD.n64 VDD.n61 6.772
R1114 VDD.n124 VDD.n109 6.772
R1115 VDD.n122 VDD.n119 6.772
R1116 VDD.n118 VDD.n115 6.772
R1117 VDD.n185 VDD.n170 6.772
R1118 VDD.n183 VDD.n180 6.772
R1119 VDD.n179 VDD.n176 6.772
R1120 VDD.n266 VDD.n251 6.772
R1121 VDD.n264 VDD.n261 6.772
R1122 VDD.n260 VDD.n257 6.772
R1123 VDD.n327 VDD.n312 6.772
R1124 VDD.n325 VDD.n322 6.772
R1125 VDD.n321 VDD.n318 6.772
R1126 VDD.n388 VDD.n373 6.772
R1127 VDD.n386 VDD.n383 6.772
R1128 VDD.n382 VDD.n379 6.772
R1129 VDD.n469 VDD.n454 6.772
R1130 VDD.n467 VDD.n464 6.772
R1131 VDD.n463 VDD.n460 6.772
R1132 VDD.n550 VDD.n535 6.772
R1133 VDD.n548 VDD.n545 6.772
R1134 VDD.n544 VDD.n541 6.772
R1135 VDD.n611 VDD.n596 6.772
R1136 VDD.n609 VDD.n606 6.772
R1137 VDD.n605 VDD.n602 6.772
R1138 VDD.n692 VDD.n677 6.772
R1139 VDD.n690 VDD.n687 6.772
R1140 VDD.n686 VDD.n683 6.772
R1141 VDD.n1452 VDD.n1437 6.772
R1142 VDD.n1450 VDD.n1447 6.772
R1143 VDD.n1446 VDD.n1443 6.772
R1144 VDD.n1391 VDD.n1376 6.772
R1145 VDD.n1389 VDD.n1386 6.772
R1146 VDD.n1385 VDD.n1382 6.772
R1147 VDD.n1310 VDD.n1295 6.772
R1148 VDD.n1308 VDD.n1305 6.772
R1149 VDD.n1304 VDD.n1301 6.772
R1150 VDD.n1229 VDD.n1214 6.772
R1151 VDD.n1227 VDD.n1224 6.772
R1152 VDD.n1223 VDD.n1220 6.772
R1153 VDD.n1168 VDD.n1153 6.772
R1154 VDD.n1166 VDD.n1163 6.772
R1155 VDD.n1162 VDD.n1159 6.772
R1156 VDD.n1087 VDD.n1072 6.772
R1157 VDD.n1085 VDD.n1082 6.772
R1158 VDD.n1081 VDD.n1078 6.772
R1159 VDD.n1026 VDD.n1011 6.772
R1160 VDD.n1024 VDD.n1021 6.772
R1161 VDD.n1020 VDD.n1017 6.772
R1162 VDD.n965 VDD.n950 6.772
R1163 VDD.n963 VDD.n960 6.772
R1164 VDD.n959 VDD.n956 6.772
R1165 VDD.n884 VDD.n869 6.772
R1166 VDD.n882 VDD.n879 6.772
R1167 VDD.n878 VDD.n875 6.772
R1168 VDD.n743 VDD.n729 6.772
R1169 VDD.n741 VDD.n738 6.772
R1170 VDD.n737 VDD.n734 6.772
R1171 VDD.n59 VDD.n58 6.772
R1172 VDD.n64 VDD.n63 6.772
R1173 VDD.n68 VDD.n67 6.772
R1174 VDD.n71 VDD.n70 6.772
R1175 VDD.n118 VDD.n117 6.772
R1176 VDD.n122 VDD.n121 6.772
R1177 VDD.n125 VDD.n124 6.772
R1178 VDD.n179 VDD.n178 6.772
R1179 VDD.n183 VDD.n182 6.772
R1180 VDD.n186 VDD.n185 6.772
R1181 VDD.n260 VDD.n259 6.772
R1182 VDD.n264 VDD.n263 6.772
R1183 VDD.n267 VDD.n266 6.772
R1184 VDD.n321 VDD.n320 6.772
R1185 VDD.n325 VDD.n324 6.772
R1186 VDD.n328 VDD.n327 6.772
R1187 VDD.n382 VDD.n381 6.772
R1188 VDD.n386 VDD.n385 6.772
R1189 VDD.n389 VDD.n388 6.772
R1190 VDD.n463 VDD.n462 6.772
R1191 VDD.n467 VDD.n466 6.772
R1192 VDD.n470 VDD.n469 6.772
R1193 VDD.n544 VDD.n543 6.772
R1194 VDD.n548 VDD.n547 6.772
R1195 VDD.n551 VDD.n550 6.772
R1196 VDD.n605 VDD.n604 6.772
R1197 VDD.n609 VDD.n608 6.772
R1198 VDD.n612 VDD.n611 6.772
R1199 VDD.n686 VDD.n685 6.772
R1200 VDD.n690 VDD.n689 6.772
R1201 VDD.n693 VDD.n692 6.772
R1202 VDD.n1446 VDD.n1445 6.772
R1203 VDD.n1450 VDD.n1449 6.772
R1204 VDD.n1453 VDD.n1452 6.772
R1205 VDD.n1385 VDD.n1384 6.772
R1206 VDD.n1389 VDD.n1388 6.772
R1207 VDD.n1392 VDD.n1391 6.772
R1208 VDD.n1304 VDD.n1303 6.772
R1209 VDD.n1308 VDD.n1307 6.772
R1210 VDD.n1311 VDD.n1310 6.772
R1211 VDD.n1223 VDD.n1222 6.772
R1212 VDD.n1227 VDD.n1226 6.772
R1213 VDD.n1230 VDD.n1229 6.772
R1214 VDD.n1162 VDD.n1161 6.772
R1215 VDD.n1166 VDD.n1165 6.772
R1216 VDD.n1169 VDD.n1168 6.772
R1217 VDD.n1081 VDD.n1080 6.772
R1218 VDD.n1085 VDD.n1084 6.772
R1219 VDD.n1088 VDD.n1087 6.772
R1220 VDD.n1020 VDD.n1019 6.772
R1221 VDD.n1024 VDD.n1023 6.772
R1222 VDD.n1027 VDD.n1026 6.772
R1223 VDD.n959 VDD.n958 6.772
R1224 VDD.n963 VDD.n962 6.772
R1225 VDD.n966 VDD.n965 6.772
R1226 VDD.n878 VDD.n877 6.772
R1227 VDD.n882 VDD.n881 6.772
R1228 VDD.n885 VDD.n884 6.772
R1229 VDD.n737 VDD.n736 6.772
R1230 VDD.n741 VDD.n740 6.772
R1231 VDD.n744 VDD.n743 6.772
R1232 VDD.n804 VDD.n803 6.772
R1233 VDD.n791 VDD.n788 6.772
R1234 VDD.n796 VDD.n793 6.772
R1235 VDD.n801 VDD.n798 6.772
R1236 VDD.n801 VDD.n800 6.772
R1237 VDD.n796 VDD.n795 6.772
R1238 VDD.n791 VDD.n790 6.772
R1239 VDD.n803 VDD.n787 6.772
R1240 VDD.n229 VDD.n225 6.69
R1241 VDD.n432 VDD.n428 6.69
R1242 VDD.n513 VDD.n509 6.69
R1243 VDD.n655 VDD.n651 6.69
R1244 VDD.n1338 VDD.n1334 6.69
R1245 VDD.n1257 VDD.n1253 6.69
R1246 VDD.n1115 VDD.n1111 6.69
R1247 VDD.n912 VDD.n908 6.69
R1248 VDD.n831 VDD.n827 6.69
R1249 VDD.n33 VDD.n23 6.487
R1250 VDD.n33 VDD.n32 6.475
R1251 VDD.n16 VDD.n15 6.458
R1252 VDD.n212 VDD.n211 6.296
R1253 VDD.n415 VDD.n414 6.296
R1254 VDD.n496 VDD.n495 6.296
R1255 VDD.n638 VDD.n637 6.296
R1256 VDD.n1355 VDD.n1354 6.296
R1257 VDD.n1274 VDD.n1273 6.296
R1258 VDD.n1132 VDD.n1131 6.296
R1259 VDD.n929 VDD.n928 6.296
R1260 VDD.n848 VDD.n847 6.296
R1261 VDD.n113 VDD.n112 6.202
R1262 VDD.n174 VDD.n173 6.202
R1263 VDD.n255 VDD.n254 6.202
R1264 VDD.n316 VDD.n315 6.202
R1265 VDD.n377 VDD.n376 6.202
R1266 VDD.n458 VDD.n457 6.202
R1267 VDD.n539 VDD.n538 6.202
R1268 VDD.n600 VDD.n599 6.202
R1269 VDD.n681 VDD.n680 6.202
R1270 VDD.n1441 VDD.n1440 6.202
R1271 VDD.n1380 VDD.n1379 6.202
R1272 VDD.n1299 VDD.n1298 6.202
R1273 VDD.n1218 VDD.n1217 6.202
R1274 VDD.n1157 VDD.n1156 6.202
R1275 VDD.n1076 VDD.n1075 6.202
R1276 VDD.n1015 VDD.n1014 6.202
R1277 VDD.n954 VDD.n953 6.202
R1278 VDD.n873 VDD.n872 6.202
R1279 VDD.n732 VDD.n731 6.202
R1280 VDD.n150 VDD.n149 4.576
R1281 VDD.n292 VDD.n291 4.576
R1282 VDD.n353 VDD.n352 4.576
R1283 VDD.n576 VDD.n575 4.576
R1284 VDD.n718 VDD.n717 4.576
R1285 VDD.n1411 VDD.n1410 4.576
R1286 VDD.n1188 VDD.n1187 4.576
R1287 VDD.n1046 VDD.n1045 4.576
R1288 VDD.n985 VDD.n984 4.576
R1289 VDD.n761 VDD.n760 4.576
R1290 VDD.n162 VDD.n159 2.754
R1291 VDD.n304 VDD.n301 2.754
R1292 VDD.n365 VDD.n362 2.754
R1293 VDD.n588 VDD.n585 2.754
R1294 VDD.n1464 VDD.n1461 2.754
R1295 VDD.n1403 VDD.n1400 2.754
R1296 VDD.n1180 VDD.n1177 2.754
R1297 VDD.n1038 VDD.n1035 2.754
R1298 VDD.n977 VDD.n974 2.754
R1299 VDD.n753 VDD.n750 2.754
R1300 VDD.n136 VDD.n133 2.361
R1301 VDD.n278 VDD.n275 2.361
R1302 VDD.n339 VDD.n336 2.361
R1303 VDD.n562 VDD.n559 2.361
R1304 VDD.n704 VDD.n701 2.361
R1305 VDD.n1429 VDD.n1426 2.361
R1306 VDD.n1206 VDD.n1203 2.361
R1307 VDD.n1064 VDD.n1061 2.361
R1308 VDD.n1003 VDD.n1000 2.361
R1309 VDD.n779 VDD.n776 2.361
R1310 VDD.n14 VDD.n7 1.329
R1311 VDD.n14 VDD.n8 1.329
R1312 VDD.n14 VDD.n11 1.329
R1313 VDD.n14 VDD.n13 1.329
R1314 VDD.n15 VDD.n14 0.696
R1315 VDD.n14 VDD.n4 0.696
R1316 VDD.n239 VDD.n236 0.393
R1317 VDD.n442 VDD.n439 0.393
R1318 VDD.n523 VDD.n520 0.393
R1319 VDD.n665 VDD.n662 0.393
R1320 VDD.n1326 VDD.n1323 0.393
R1321 VDD.n1245 VDD.n1242 0.393
R1322 VDD.n1103 VDD.n1100 0.393
R1323 VDD.n900 VDD.n897 0.393
R1324 VDD.n819 VDD.n816 0.393
R1325 VDD.n69 VDD.n68 0.365
R1326 VDD.n69 VDD.n64 0.365
R1327 VDD.n69 VDD.n59 0.365
R1328 VDD.n70 VDD.n69 0.365
R1329 VDD.n123 VDD.n122 0.365
R1330 VDD.n123 VDD.n118 0.365
R1331 VDD.n124 VDD.n123 0.365
R1332 VDD.n184 VDD.n183 0.365
R1333 VDD.n184 VDD.n179 0.365
R1334 VDD.n185 VDD.n184 0.365
R1335 VDD.n265 VDD.n264 0.365
R1336 VDD.n265 VDD.n260 0.365
R1337 VDD.n266 VDD.n265 0.365
R1338 VDD.n326 VDD.n325 0.365
R1339 VDD.n326 VDD.n321 0.365
R1340 VDD.n327 VDD.n326 0.365
R1341 VDD.n387 VDD.n386 0.365
R1342 VDD.n387 VDD.n382 0.365
R1343 VDD.n388 VDD.n387 0.365
R1344 VDD.n468 VDD.n467 0.365
R1345 VDD.n468 VDD.n463 0.365
R1346 VDD.n469 VDD.n468 0.365
R1347 VDD.n549 VDD.n548 0.365
R1348 VDD.n549 VDD.n544 0.365
R1349 VDD.n550 VDD.n549 0.365
R1350 VDD.n610 VDD.n609 0.365
R1351 VDD.n610 VDD.n605 0.365
R1352 VDD.n611 VDD.n610 0.365
R1353 VDD.n691 VDD.n690 0.365
R1354 VDD.n691 VDD.n686 0.365
R1355 VDD.n692 VDD.n691 0.365
R1356 VDD.n1451 VDD.n1450 0.365
R1357 VDD.n1451 VDD.n1446 0.365
R1358 VDD.n1452 VDD.n1451 0.365
R1359 VDD.n1390 VDD.n1389 0.365
R1360 VDD.n1390 VDD.n1385 0.365
R1361 VDD.n1391 VDD.n1390 0.365
R1362 VDD.n1309 VDD.n1308 0.365
R1363 VDD.n1309 VDD.n1304 0.365
R1364 VDD.n1310 VDD.n1309 0.365
R1365 VDD.n1228 VDD.n1227 0.365
R1366 VDD.n1228 VDD.n1223 0.365
R1367 VDD.n1229 VDD.n1228 0.365
R1368 VDD.n1167 VDD.n1166 0.365
R1369 VDD.n1167 VDD.n1162 0.365
R1370 VDD.n1168 VDD.n1167 0.365
R1371 VDD.n1086 VDD.n1085 0.365
R1372 VDD.n1086 VDD.n1081 0.365
R1373 VDD.n1087 VDD.n1086 0.365
R1374 VDD.n1025 VDD.n1024 0.365
R1375 VDD.n1025 VDD.n1020 0.365
R1376 VDD.n1026 VDD.n1025 0.365
R1377 VDD.n964 VDD.n963 0.365
R1378 VDD.n964 VDD.n959 0.365
R1379 VDD.n965 VDD.n964 0.365
R1380 VDD.n883 VDD.n882 0.365
R1381 VDD.n883 VDD.n878 0.365
R1382 VDD.n884 VDD.n883 0.365
R1383 VDD.n742 VDD.n741 0.365
R1384 VDD.n742 VDD.n737 0.365
R1385 VDD.n743 VDD.n742 0.365
R1386 VDD.n802 VDD.n801 0.365
R1387 VDD.n802 VDD.n796 0.365
R1388 VDD.n802 VDD.n791 0.365
R1389 VDD.n803 VDD.n802 0.365
R1390 VDD.n78 VDD.n51 0.29
R1391 VDD.n132 VDD.n106 0.29
R1392 VDD.n193 VDD.n167 0.29
R1393 VDD.n274 VDD.n248 0.29
R1394 VDD.n335 VDD.n309 0.29
R1395 VDD.n396 VDD.n370 0.29
R1396 VDD.n477 VDD.n451 0.29
R1397 VDD.n558 VDD.n532 0.29
R1398 VDD.n619 VDD.n593 0.29
R1399 VDD.n700 VDD.n674 0.29
R1400 VDD.n1460 VDD.n1434 0.29
R1401 VDD.n1399 VDD.n1373 0.29
R1402 VDD.n1318 VDD.n1292 0.29
R1403 VDD.n1237 VDD.n1211 0.29
R1404 VDD.n1176 VDD.n1150 0.29
R1405 VDD.n1095 VDD.n1069 0.29
R1406 VDD.n1034 VDD.n1008 0.29
R1407 VDD.n973 VDD.n947 0.29
R1408 VDD.n892 VDD.n866 0.29
R1409 VDD.n811 VDD.n784 0.29
R1410 VDD.n749 VDD 0.207
R1411 VDD.n223 VDD.n218 0.197
R1412 VDD.n426 VDD.n421 0.197
R1413 VDD.n507 VDD.n502 0.197
R1414 VDD.n649 VDD.n644 0.197
R1415 VDD.n1349 VDD.n1344 0.197
R1416 VDD.n1268 VDD.n1263 0.197
R1417 VDD.n1126 VDD.n1121 0.197
R1418 VDD.n923 VDD.n918 0.197
R1419 VDD.n842 VDD.n837 0.197
R1420 VDD.n39 VDD.n35 0.181
R1421 VDD.n94 VDD.n90 0.181
R1422 VDD.n153 VDD.n148 0.181
R1423 VDD.n295 VDD.n290 0.181
R1424 VDD.n356 VDD.n351 0.181
R1425 VDD.n579 VDD.n574 0.181
R1426 VDD.n721 VDD.n716 0.181
R1427 VDD.n1420 VDD.n1414 0.181
R1428 VDD.n1197 VDD.n1191 0.181
R1429 VDD.n1055 VDD.n1049 0.181
R1430 VDD.n994 VDD.n988 0.181
R1431 VDD.n770 VDD.n764 0.181
R1432 VDD.n35 VDD.n34 0.145
R1433 VDD.n43 VDD.n39 0.145
R1434 VDD.n47 VDD.n43 0.145
R1435 VDD.n51 VDD.n47 0.145
R1436 VDD.n82 VDD.n78 0.145
R1437 VDD.n86 VDD.n82 0.145
R1438 VDD.n90 VDD.n86 0.145
R1439 VDD.n98 VDD.n94 0.145
R1440 VDD.n102 VDD.n98 0.145
R1441 VDD.n106 VDD.n102 0.145
R1442 VDD.n137 VDD.n132 0.145
R1443 VDD.n142 VDD.n137 0.145
R1444 VDD.n148 VDD.n142 0.145
R1445 VDD.n158 VDD.n153 0.145
R1446 VDD.n163 VDD.n158 0.145
R1447 VDD.n167 VDD.n163 0.145
R1448 VDD.n197 VDD.n193 0.145
R1449 VDD.n201 VDD.n197 0.145
R1450 VDD.n206 VDD.n201 0.145
R1451 VDD.n213 VDD.n206 0.145
R1452 VDD.n218 VDD.n213 0.145
R1453 VDD.n230 VDD.n223 0.145
R1454 VDD.n235 VDD.n230 0.145
R1455 VDD.n240 VDD.n235 0.145
R1456 VDD.n244 VDD.n240 0.145
R1457 VDD.n248 VDD.n244 0.145
R1458 VDD.n279 VDD.n274 0.145
R1459 VDD.n284 VDD.n279 0.145
R1460 VDD.n290 VDD.n284 0.145
R1461 VDD.n300 VDD.n295 0.145
R1462 VDD.n305 VDD.n300 0.145
R1463 VDD.n309 VDD.n305 0.145
R1464 VDD.n340 VDD.n335 0.145
R1465 VDD.n345 VDD.n340 0.145
R1466 VDD.n351 VDD.n345 0.145
R1467 VDD.n361 VDD.n356 0.145
R1468 VDD.n366 VDD.n361 0.145
R1469 VDD.n370 VDD.n366 0.145
R1470 VDD.n400 VDD.n396 0.145
R1471 VDD.n404 VDD.n400 0.145
R1472 VDD.n409 VDD.n404 0.145
R1473 VDD.n416 VDD.n409 0.145
R1474 VDD.n421 VDD.n416 0.145
R1475 VDD.n433 VDD.n426 0.145
R1476 VDD.n438 VDD.n433 0.145
R1477 VDD.n443 VDD.n438 0.145
R1478 VDD.n447 VDD.n443 0.145
R1479 VDD.n451 VDD.n447 0.145
R1480 VDD.n481 VDD.n477 0.145
R1481 VDD.n485 VDD.n481 0.145
R1482 VDD.n490 VDD.n485 0.145
R1483 VDD.n497 VDD.n490 0.145
R1484 VDD.n502 VDD.n497 0.145
R1485 VDD.n514 VDD.n507 0.145
R1486 VDD.n519 VDD.n514 0.145
R1487 VDD.n524 VDD.n519 0.145
R1488 VDD.n528 VDD.n524 0.145
R1489 VDD.n532 VDD.n528 0.145
R1490 VDD.n563 VDD.n558 0.145
R1491 VDD.n568 VDD.n563 0.145
R1492 VDD.n574 VDD.n568 0.145
R1493 VDD.n584 VDD.n579 0.145
R1494 VDD.n589 VDD.n584 0.145
R1495 VDD.n593 VDD.n589 0.145
R1496 VDD.n623 VDD.n619 0.145
R1497 VDD.n627 VDD.n623 0.145
R1498 VDD.n632 VDD.n627 0.145
R1499 VDD.n639 VDD.n632 0.145
R1500 VDD.n644 VDD.n639 0.145
R1501 VDD.n656 VDD.n649 0.145
R1502 VDD.n661 VDD.n656 0.145
R1503 VDD.n666 VDD.n661 0.145
R1504 VDD.n670 VDD.n666 0.145
R1505 VDD.n674 VDD.n670 0.145
R1506 VDD.n705 VDD.n700 0.145
R1507 VDD.n710 VDD.n705 0.145
R1508 VDD.n716 VDD.n710 0.145
R1509 VDD.n726 VDD.n721 0.145
R1510 VDD.n1465 VDD.n1460 0.145
R1511 VDD.n1434 VDD.n1430 0.145
R1512 VDD.n1430 VDD.n1425 0.145
R1513 VDD.n1425 VDD.n1420 0.145
R1514 VDD.n1414 VDD.n1409 0.145
R1515 VDD.n1409 VDD.n1404 0.145
R1516 VDD.n1404 VDD.n1399 0.145
R1517 VDD.n1373 VDD.n1369 0.145
R1518 VDD.n1369 VDD.n1365 0.145
R1519 VDD.n1365 VDD.n1361 0.145
R1520 VDD.n1361 VDD.n1356 0.145
R1521 VDD.n1356 VDD.n1349 0.145
R1522 VDD.n1344 VDD.n1339 0.145
R1523 VDD.n1339 VDD.n1332 0.145
R1524 VDD.n1332 VDD.n1327 0.145
R1525 VDD.n1327 VDD.n1322 0.145
R1526 VDD.n1322 VDD.n1318 0.145
R1527 VDD.n1292 VDD.n1288 0.145
R1528 VDD.n1288 VDD.n1284 0.145
R1529 VDD.n1284 VDD.n1280 0.145
R1530 VDD.n1280 VDD.n1275 0.145
R1531 VDD.n1275 VDD.n1268 0.145
R1532 VDD.n1263 VDD.n1258 0.145
R1533 VDD.n1258 VDD.n1251 0.145
R1534 VDD.n1251 VDD.n1246 0.145
R1535 VDD.n1246 VDD.n1241 0.145
R1536 VDD.n1241 VDD.n1237 0.145
R1537 VDD.n1211 VDD.n1207 0.145
R1538 VDD.n1207 VDD.n1202 0.145
R1539 VDD.n1202 VDD.n1197 0.145
R1540 VDD.n1191 VDD.n1186 0.145
R1541 VDD.n1186 VDD.n1181 0.145
R1542 VDD.n1181 VDD.n1176 0.145
R1543 VDD.n1150 VDD.n1146 0.145
R1544 VDD.n1146 VDD.n1142 0.145
R1545 VDD.n1142 VDD.n1138 0.145
R1546 VDD.n1138 VDD.n1133 0.145
R1547 VDD.n1133 VDD.n1126 0.145
R1548 VDD.n1121 VDD.n1116 0.145
R1549 VDD.n1116 VDD.n1109 0.145
R1550 VDD.n1109 VDD.n1104 0.145
R1551 VDD.n1104 VDD.n1099 0.145
R1552 VDD.n1099 VDD.n1095 0.145
R1553 VDD.n1069 VDD.n1065 0.145
R1554 VDD.n1065 VDD.n1060 0.145
R1555 VDD.n1060 VDD.n1055 0.145
R1556 VDD.n1049 VDD.n1044 0.145
R1557 VDD.n1044 VDD.n1039 0.145
R1558 VDD.n1039 VDD.n1034 0.145
R1559 VDD.n1008 VDD.n1004 0.145
R1560 VDD.n1004 VDD.n999 0.145
R1561 VDD.n999 VDD.n994 0.145
R1562 VDD.n988 VDD.n983 0.145
R1563 VDD.n983 VDD.n978 0.145
R1564 VDD.n978 VDD.n973 0.145
R1565 VDD.n947 VDD.n943 0.145
R1566 VDD.n943 VDD.n939 0.145
R1567 VDD.n939 VDD.n935 0.145
R1568 VDD.n935 VDD.n930 0.145
R1569 VDD.n930 VDD.n923 0.145
R1570 VDD.n918 VDD.n913 0.145
R1571 VDD.n913 VDD.n906 0.145
R1572 VDD.n906 VDD.n901 0.145
R1573 VDD.n901 VDD.n896 0.145
R1574 VDD.n896 VDD.n892 0.145
R1575 VDD.n866 VDD.n862 0.145
R1576 VDD.n862 VDD.n858 0.145
R1577 VDD.n858 VDD.n854 0.145
R1578 VDD.n854 VDD.n849 0.145
R1579 VDD.n849 VDD.n842 0.145
R1580 VDD.n837 VDD.n832 0.145
R1581 VDD.n832 VDD.n825 0.145
R1582 VDD.n825 VDD.n820 0.145
R1583 VDD.n820 VDD.n815 0.145
R1584 VDD.n815 VDD.n811 0.145
R1585 VDD.n784 VDD.n780 0.145
R1586 VDD.n780 VDD.n775 0.145
R1587 VDD.n775 VDD.n770 0.145
R1588 VDD.n764 VDD.n759 0.145
R1589 VDD.n759 VDD.n754 0.145
R1590 VDD.n754 VDD.n749 0.145
R1591 VDD VDD.n1465 0.082
R1592 VDD VDD.n726 0.062
R1593 a_8357_1050.n0 a_8357_1050.t5 512.525
R1594 a_8357_1050.n0 a_8357_1050.t7 371.139
R1595 a_8357_1050.n1 a_8357_1050.t6 340.774
R1596 a_8357_1050.n6 a_8357_1050.n5 263.698
R1597 a_8357_1050.n6 a_8357_1050.n1 153.315
R1598 a_8357_1050.n1 a_8357_1050.n0 109.607
R1599 a_8357_1050.n8 a_8357_1050.n6 99.394
R1600 a_8357_1050.n8 a_8357_1050.n7 76.002
R1601 a_8357_1050.n5 a_8357_1050.n4 30
R1602 a_8357_1050.n3 a_8357_1050.n2 24.383
R1603 a_8357_1050.n5 a_8357_1050.n3 23.684
R1604 a_8357_1050.n7 a_8357_1050.t4 14.282
R1605 a_8357_1050.n7 a_8357_1050.t3 14.282
R1606 a_8357_1050.n9 a_8357_1050.t1 14.282
R1607 a_8357_1050.t2 a_8357_1050.n9 14.282
R1608 a_8357_1050.n9 a_8357_1050.n8 12.848
R1609 SN.n14 SN.t3 479.223
R1610 SN.n11 SN.t12 479.223
R1611 SN.n8 SN.t13 479.223
R1612 SN.n5 SN.t2 479.223
R1613 SN.n2 SN.t9 479.223
R1614 SN.n0 SN.t8 479.223
R1615 SN.n14 SN.t14 375.52
R1616 SN.n11 SN.t4 375.52
R1617 SN.n8 SN.t15 375.52
R1618 SN.n5 SN.t7 375.52
R1619 SN.n2 SN.t17 375.52
R1620 SN.n0 SN.t16 375.52
R1621 SN.n15 SN.n14 175.429
R1622 SN.n12 SN.n11 175.429
R1623 SN.n9 SN.n8 175.429
R1624 SN.n6 SN.n5 175.429
R1625 SN.n3 SN.n2 175.429
R1626 SN.n1 SN.n0 175.429
R1627 SN.n15 SN.t11 162.048
R1628 SN.n12 SN.t1 162.048
R1629 SN.n9 SN.t0 162.048
R1630 SN.n6 SN.t6 162.048
R1631 SN.n3 SN.t5 162.048
R1632 SN.n1 SN.t10 162.048
R1633 SN.n4 SN.n1 84.388
R1634 SN.n4 SN.n3 76
R1635 SN.n7 SN.n6 76
R1636 SN.n10 SN.n9 76
R1637 SN.n13 SN.n12 76
R1638 SN.n16 SN.n15 76
R1639 SN.n7 SN.n4 9.476
R1640 SN.n13 SN.n10 9.476
R1641 SN.n10 SN.n7 8.388
R1642 SN.n16 SN.n13 8.388
R1643 SN.n16 SN 0.046
R1644 a_6603_103.t0 a_6603_103.n0 117.777
R1645 a_6603_103.n2 a_6603_103.n1 55.228
R1646 a_6603_103.n4 a_6603_103.n3 9.111
R1647 a_6603_103.n8 a_6603_103.n6 7.859
R1648 a_6603_103.t0 a_6603_103.n2 4.04
R1649 a_6603_103.t0 a_6603_103.n8 3.034
R1650 a_6603_103.n6 a_6603_103.n4 1.964
R1651 a_6603_103.n6 a_6603_103.n5 1.964
R1652 a_6603_103.n8 a_6603_103.n7 0.443
R1653 a_6884_210.n10 a_6884_210.n8 82.852
R1654 a_6884_210.n11 a_6884_210.n0 49.6
R1655 a_6884_210.n7 a_6884_210.n6 32.833
R1656 a_6884_210.n8 a_6884_210.t1 32.416
R1657 a_6884_210.n10 a_6884_210.n9 27.2
R1658 a_6884_210.n3 a_6884_210.n2 23.284
R1659 a_6884_210.n11 a_6884_210.n10 22.4
R1660 a_6884_210.n7 a_6884_210.n4 19.017
R1661 a_6884_210.n6 a_6884_210.n5 13.494
R1662 a_6884_210.t1 a_6884_210.n1 7.04
R1663 a_6884_210.t1 a_6884_210.n3 5.727
R1664 a_6884_210.n8 a_6884_210.n7 1.435
R1665 a_3473_1050.n3 a_3473_1050.t6 512.525
R1666 a_3473_1050.n3 a_3473_1050.t5 371.139
R1667 a_3473_1050.n4 a_3473_1050.t7 340.774
R1668 a_3473_1050.n7 a_3473_1050.n5 270.22
R1669 a_3473_1050.n5 a_3473_1050.n4 153.315
R1670 a_3473_1050.n4 a_3473_1050.n3 109.607
R1671 a_3473_1050.n5 a_3473_1050.n2 99.394
R1672 a_3473_1050.n2 a_3473_1050.n1 76.002
R1673 a_3473_1050.n7 a_3473_1050.n6 15.218
R1674 a_3473_1050.n0 a_3473_1050.t4 14.282
R1675 a_3473_1050.n0 a_3473_1050.t2 14.282
R1676 a_3473_1050.n1 a_3473_1050.t1 14.282
R1677 a_3473_1050.n1 a_3473_1050.t0 14.282
R1678 a_3473_1050.n2 a_3473_1050.n0 12.85
R1679 a_3473_1050.n8 a_3473_1050.n7 12.014
R1680 a_3599_411.n3 a_3599_411.t7 512.525
R1681 a_3599_411.n2 a_3599_411.t11 512.525
R1682 a_3599_411.n7 a_3599_411.t15 472.359
R1683 a_3599_411.n7 a_3599_411.t9 384.527
R1684 a_3599_411.n3 a_3599_411.t13 371.139
R1685 a_3599_411.n2 a_3599_411.t8 371.139
R1686 a_3599_411.n4 a_3599_411.n3 265.439
R1687 a_3599_411.n8 a_3599_411.t12 214.619
R1688 a_3599_411.n15 a_3599_411.n14 197.352
R1689 a_3599_411.n14 a_3599_411.n13 186.551
R1690 a_3599_411.n6 a_3599_411.n2 185.78
R1691 a_3599_411.n4 a_3599_411.t14 176.995
R1692 a_3599_411.n5 a_3599_411.t10 170.569
R1693 a_3599_411.n5 a_3599_411.n4 153.043
R1694 a_3599_411.n8 a_3599_411.n7 136.613
R1695 a_3599_411.n9 a_3599_411.n6 116.763
R1696 a_3599_411.n9 a_3599_411.n8 80.035
R1697 a_3599_411.n6 a_3599_411.n5 79.658
R1698 a_3599_411.n17 a_3599_411.n16 79.231
R1699 a_3599_411.n14 a_3599_411.n9 76
R1700 a_3599_411.n16 a_3599_411.n15 63.152
R1701 a_3599_411.n13 a_3599_411.n12 30
R1702 a_3599_411.n11 a_3599_411.n10 24.383
R1703 a_3599_411.n13 a_3599_411.n11 23.684
R1704 a_3599_411.n15 a_3599_411.n1 16.08
R1705 a_3599_411.n16 a_3599_411.n0 16.08
R1706 a_3599_411.n1 a_3599_411.t6 14.282
R1707 a_3599_411.n1 a_3599_411.t5 14.282
R1708 a_3599_411.n0 a_3599_411.t2 14.282
R1709 a_3599_411.n0 a_3599_411.t3 14.282
R1710 a_3599_411.n17 a_3599_411.t0 14.282
R1711 a_3599_411.t1 a_3599_411.n17 14.282
R1712 CLK.n15 CLK.t17 472.359
R1713 CLK.n6 CLK.t0 472.359
R1714 CLK.n0 CLK.t4 472.359
R1715 CLK.n20 CLK.t9 459.505
R1716 CLK.n11 CLK.t2 459.505
R1717 CLK.n2 CLK.t15 459.505
R1718 CLK.n20 CLK.t14 384.527
R1719 CLK.n15 CLK.t1 384.527
R1720 CLK.n11 CLK.t5 384.527
R1721 CLK.n6 CLK.t8 384.527
R1722 CLK.n2 CLK.t7 384.527
R1723 CLK.n0 CLK.t13 384.527
R1724 CLK.n21 CLK.t11 322.152
R1725 CLK.n12 CLK.t12 322.151
R1726 CLK.n3 CLK.t3 322.151
R1727 CLK.n1 CLK.t10 321.724
R1728 CLK.n17 CLK.t16 319.581
R1729 CLK.n8 CLK.t6 319.581
R1730 CLK.n9 CLK.n8 75.621
R1731 CLK.n18 CLK.n17 75.621
R1732 CLK.n22 CLK.n21 49.342
R1733 CLK.n4 CLK.n3 49.342
R1734 CLK.n13 CLK.n12 49.342
R1735 CLK.n4 CLK.n1 43.573
R1736 CLK.n21 CLK.n20 27.599
R1737 CLK.n3 CLK.n2 27.599
R1738 CLK.n12 CLK.n11 27.599
R1739 CLK.n1 CLK.n0 23.329
R1740 CLK.n16 CLK.n15 21.176
R1741 CLK.n7 CLK.n6 21.176
R1742 CLK.n5 CLK.n4 11.101
R1743 CLK.n14 CLK.n13 11.101
R1744 CLK.n13 CLK.n10 6.718
R1745 CLK.n22 CLK.n19 6.718
R1746 CLK.n17 CLK.n16 4.419
R1747 CLK.n8 CLK.n7 4.419
R1748 CLK.n22 CLK 0.046
R1749 CLK.n10 CLK.n9 0.038
R1750 CLK.n19 CLK.n18 0.038
R1751 CLK.n9 CLK.n5 0.008
R1752 CLK.n18 CLK.n14 0.008
R1753 a_6149_989.n2 a_6149_989.t5 454.685
R1754 a_6149_989.n4 a_6149_989.t8 454.685
R1755 a_6149_989.n0 a_6149_989.t10 454.685
R1756 a_6149_989.n2 a_6149_989.t11 428.979
R1757 a_6149_989.n4 a_6149_989.t13 428.979
R1758 a_6149_989.n0 a_6149_989.t9 428.979
R1759 a_6149_989.n3 a_6149_989.t7 264.512
R1760 a_6149_989.n5 a_6149_989.t6 264.512
R1761 a_6149_989.n1 a_6149_989.t12 264.512
R1762 a_6149_989.n12 a_6149_989.n11 237.145
R1763 a_6149_989.n14 a_6149_989.n12 125.947
R1764 a_6149_989.n7 a_6149_989.n1 81.396
R1765 a_6149_989.n6 a_6149_989.n5 79.491
R1766 a_6149_989.n14 a_6149_989.n13 76.002
R1767 a_6149_989.n6 a_6149_989.n3 76
R1768 a_6149_989.n12 a_6149_989.n7 76
R1769 a_6149_989.n3 a_6149_989.n2 71.894
R1770 a_6149_989.n5 a_6149_989.n4 71.894
R1771 a_6149_989.n1 a_6149_989.n0 71.894
R1772 a_6149_989.n11 a_6149_989.n10 30
R1773 a_6149_989.n9 a_6149_989.n8 24.383
R1774 a_6149_989.n11 a_6149_989.n9 23.684
R1775 a_6149_989.n13 a_6149_989.t4 14.282
R1776 a_6149_989.n13 a_6149_989.t0 14.282
R1777 a_6149_989.t2 a_6149_989.n15 14.282
R1778 a_6149_989.n15 a_6149_989.t1 14.282
R1779 a_6149_989.n15 a_6149_989.n14 12.848
R1780 a_6149_989.n7 a_6149_989.n6 2.947
R1781 a_14869_1051.n4 a_14869_1051.n3 195.987
R1782 a_14869_1051.n2 a_14869_1051.t1 89.553
R1783 a_14869_1051.n5 a_14869_1051.n4 75.27
R1784 a_14869_1051.n3 a_14869_1051.n2 75.214
R1785 a_14869_1051.n4 a_14869_1051.n0 36.519
R1786 a_14869_1051.n3 a_14869_1051.t2 14.338
R1787 a_14869_1051.n0 a_14869_1051.t7 14.282
R1788 a_14869_1051.n0 a_14869_1051.t6 14.282
R1789 a_14869_1051.n1 a_14869_1051.t0 14.282
R1790 a_14869_1051.n1 a_14869_1051.t3 14.282
R1791 a_14869_1051.t5 a_14869_1051.n5 14.282
R1792 a_14869_1051.n5 a_14869_1051.t4 14.282
R1793 a_14869_1051.n2 a_14869_1051.n1 12.119
R1794 a_13367_411.n1 a_13367_411.t8 475.572
R1795 a_13367_411.n6 a_13367_411.t15 472.359
R1796 a_13367_411.n3 a_13367_411.t11 469.145
R1797 a_13367_411.n6 a_13367_411.t10 384.527
R1798 a_13367_411.n3 a_13367_411.t14 384.527
R1799 a_13367_411.n1 a_13367_411.t12 384.527
R1800 a_13367_411.n7 a_13367_411.t7 294.278
R1801 a_13367_411.n4 a_13367_411.t13 294.278
R1802 a_13367_411.n2 a_13367_411.t9 294.278
R1803 a_13367_411.n12 a_13367_411.n11 281.733
R1804 a_13367_411.n13 a_13367_411.n12 117.693
R1805 a_13367_411.n5 a_13367_411.n2 80.851
R1806 a_13367_411.n8 a_13367_411.n7 80.035
R1807 a_13367_411.n15 a_13367_411.n14 79.232
R1808 a_13367_411.n5 a_13367_411.n4 76
R1809 a_13367_411.n12 a_13367_411.n8 76
R1810 a_13367_411.n15 a_13367_411.n13 63.152
R1811 a_13367_411.n2 a_13367_411.n1 57.842
R1812 a_13367_411.n7 a_13367_411.n6 56.954
R1813 a_13367_411.n4 a_13367_411.n3 56.833
R1814 a_13367_411.n11 a_13367_411.n10 22.578
R1815 a_13367_411.n13 a_13367_411.n0 16.08
R1816 a_13367_411.n16 a_13367_411.n15 16.078
R1817 a_13367_411.n0 a_13367_411.t5 14.282
R1818 a_13367_411.n0 a_13367_411.t2 14.282
R1819 a_13367_411.n14 a_13367_411.t4 14.282
R1820 a_13367_411.n14 a_13367_411.t3 14.282
R1821 a_13367_411.t1 a_13367_411.n16 14.282
R1822 a_13367_411.n16 a_13367_411.t0 14.282
R1823 a_13367_411.n11 a_13367_411.n9 8.58
R1824 a_13367_411.n8 a_13367_411.n5 1.859
R1825 a_13136_101.t0 a_13136_101.n1 93.333
R1826 a_13136_101.n4 a_13136_101.n2 55.07
R1827 a_13136_101.t0 a_13136_101.n0 8.137
R1828 a_13136_101.n4 a_13136_101.n3 4.619
R1829 a_13136_101.t0 a_13136_101.n4 0.071
R1830 a_13241_1050.n0 a_13241_1050.t5 512.525
R1831 a_13241_1050.n0 a_13241_1050.t6 371.139
R1832 a_13241_1050.n1 a_13241_1050.t7 368.112
R1833 a_13241_1050.n3 a_13241_1050.n2 311.99
R1834 a_13241_1050.n3 a_13241_1050.n1 126.657
R1835 a_13241_1050.n1 a_13241_1050.n0 79.811
R1836 a_13241_1050.n5 a_13241_1050.n4 76.002
R1837 a_13241_1050.n5 a_13241_1050.n3 72.841
R1838 a_13241_1050.n4 a_13241_1050.t0 14.282
R1839 a_13241_1050.n4 a_13241_1050.t1 14.282
R1840 a_13241_1050.n6 a_13241_1050.t3 14.282
R1841 a_13241_1050.t4 a_13241_1050.n6 14.282
R1842 a_13241_1050.n6 a_13241_1050.n5 12.848
R1843 a_4013_103.t0 a_4013_103.n3 117.777
R1844 a_4013_103.n6 a_4013_103.n5 45.444
R1845 a_4013_103.t0 a_4013_103.n6 21.213
R1846 a_4013_103.t0 a_4013_103.n4 11.595
R1847 a_4013_103.n2 a_4013_103.n0 8.543
R1848 a_4013_103.t0 a_4013_103.n2 3.034
R1849 a_4013_103.n2 a_4013_103.n1 0.443
R1850 a_4294_210.n10 a_4294_210.n8 82.852
R1851 a_4294_210.n11 a_4294_210.n0 49.6
R1852 a_4294_210.n7 a_4294_210.n6 32.833
R1853 a_4294_210.n8 a_4294_210.t1 32.416
R1854 a_4294_210.n10 a_4294_210.n9 27.2
R1855 a_4294_210.n3 a_4294_210.n2 23.284
R1856 a_4294_210.n11 a_4294_210.n10 22.4
R1857 a_4294_210.n7 a_4294_210.n4 19.017
R1858 a_4294_210.n6 a_4294_210.n5 13.494
R1859 a_4294_210.t1 a_4294_210.n1 7.04
R1860 a_4294_210.t1 a_4294_210.n3 5.727
R1861 a_4294_210.n8 a_4294_210.n7 1.435
R1862 a_9985_1050.n5 a_9985_1050.t9 512.525
R1863 a_9985_1050.n3 a_9985_1050.t8 512.525
R1864 a_9985_1050.n5 a_9985_1050.t7 371.139
R1865 a_9985_1050.n3 a_9985_1050.t6 371.139
R1866 a_9985_1050.n4 a_9985_1050.t5 234.562
R1867 a_9985_1050.n6 a_9985_1050.t10 234.204
R1868 a_9985_1050.n6 a_9985_1050.n5 216.178
R1869 a_9985_1050.n4 a_9985_1050.n3 215.819
R1870 a_9985_1050.n8 a_9985_1050.n2 205.605
R1871 a_9985_1050.n10 a_9985_1050.n8 164.008
R1872 a_9985_1050.n7 a_9985_1050.n4 79.488
R1873 a_9985_1050.n8 a_9985_1050.n7 77.314
R1874 a_9985_1050.n2 a_9985_1050.n1 76.002
R1875 a_9985_1050.n7 a_9985_1050.n6 76
R1876 a_9985_1050.n10 a_9985_1050.n9 15.218
R1877 a_9985_1050.n0 a_9985_1050.t3 14.282
R1878 a_9985_1050.n0 a_9985_1050.t4 14.282
R1879 a_9985_1050.n1 a_9985_1050.t0 14.282
R1880 a_9985_1050.n1 a_9985_1050.t1 14.282
R1881 a_9985_1050.n2 a_9985_1050.n0 12.85
R1882 a_9985_1050.n11 a_9985_1050.n10 12.014
R1883 a_11487_103.t0 a_11487_103.n0 117.777
R1884 a_11487_103.n2 a_11487_103.n1 55.228
R1885 a_11487_103.n4 a_11487_103.n3 9.111
R1886 a_11487_103.n8 a_11487_103.n6 7.859
R1887 a_11487_103.t0 a_11487_103.n2 4.04
R1888 a_11487_103.t0 a_11487_103.n8 3.034
R1889 a_11487_103.n6 a_11487_103.n4 1.964
R1890 a_11487_103.n6 a_11487_103.n5 1.964
R1891 a_11487_103.n8 a_11487_103.n7 0.443
R1892 GND.n29 GND.n27 219.745
R1893 GND.n62 GND.n60 219.745
R1894 GND.n413 GND.n412 219.745
R1895 GND.n455 GND.n453 219.745
R1896 GND.n497 GND.n495 219.745
R1897 GND.n527 GND.n525 219.745
R1898 GND.n557 GND.n555 219.745
R1899 GND.n599 GND.n597 219.745
R1900 GND.n629 GND.n627 219.745
R1901 GND.n671 GND.n669 219.745
R1902 GND.n713 GND.n711 219.745
R1903 GND.n743 GND.n741 219.745
R1904 GND.n362 GND.n360 219.745
R1905 GND.n317 GND.n315 219.745
R1906 GND.n287 GND.n285 219.745
R1907 GND.n242 GND.n240 219.745
R1908 GND.n200 GND.n198 219.745
R1909 GND.n170 GND.n168 219.745
R1910 GND.n140 GND.n138 219.745
R1911 GND.n95 GND.n94 219.745
R1912 GND.n231 GND.n230 85.559
R1913 GND.n680 GND.n679 85.559
R1914 GND.n638 GND.n637 85.559
R1915 GND.n566 GND.n565 85.559
R1916 GND.n464 GND.n463 85.559
R1917 GND.n422 GND.n421 85.559
R1918 GND.n29 GND.n28 85.529
R1919 GND.n62 GND.n61 85.529
R1920 GND.n413 GND.n411 85.529
R1921 GND.n455 GND.n454 85.529
R1922 GND.n497 GND.n496 85.529
R1923 GND.n527 GND.n526 85.529
R1924 GND.n557 GND.n556 85.529
R1925 GND.n599 GND.n598 85.529
R1926 GND.n629 GND.n628 85.529
R1927 GND.n671 GND.n670 85.529
R1928 GND.n713 GND.n712 85.529
R1929 GND.n743 GND.n742 85.529
R1930 GND.n362 GND.n361 85.529
R1931 GND.n317 GND.n316 85.529
R1932 GND.n287 GND.n286 85.529
R1933 GND.n242 GND.n241 85.529
R1934 GND.n200 GND.n199 85.529
R1935 GND.n170 GND.n169 85.529
R1936 GND.n140 GND.n139 85.529
R1937 GND.n95 GND.n93 85.529
R1938 GND.n158 GND.n157 84.842
R1939 GND.n188 GND.n187 84.842
R1940 GND.n305 GND.n304 84.842
R1941 GND.n380 GND.n379 84.842
R1942 GND.n721 GND.n720 84.842
R1943 GND.n607 GND.n606 84.842
R1944 GND.n535 GND.n534 84.842
R1945 GND.n505 GND.n504 84.842
R1946 GND.n391 GND.n390 84.842
R1947 GND.n386 GND.n385 76
R1948 GND.n42 GND.n41 76
R1949 GND.n45 GND.n44 76
R1950 GND.n53 GND.n52 76
R1951 GND.n56 GND.n55 76
R1952 GND.n59 GND.n58 76
R1953 GND.n66 GND.n65 76
R1954 GND.n69 GND.n68 76
R1955 GND.n72 GND.n71 76
R1956 GND.n75 GND.n74 76
R1957 GND.n78 GND.n77 76
R1958 GND.n86 GND.n85 76
R1959 GND.n89 GND.n88 76
R1960 GND.n92 GND.n91 76
R1961 GND.n99 GND.n98 76
R1962 GND.n102 GND.n101 76
R1963 GND.n105 GND.n104 76
R1964 GND.n108 GND.n107 76
R1965 GND.n111 GND.n110 76
R1966 GND.n114 GND.n113 76
R1967 GND.n117 GND.n116 76
R1968 GND.n120 GND.n119 76
R1969 GND.n123 GND.n122 76
R1970 GND.n131 GND.n130 76
R1971 GND.n134 GND.n133 76
R1972 GND.n137 GND.n136 76
R1973 GND.n144 GND.n143 76
R1974 GND.n147 GND.n146 76
R1975 GND.n150 GND.n149 76
R1976 GND.n153 GND.n152 76
R1977 GND.n156 GND.n155 76
R1978 GND.n161 GND.n160 76
R1979 GND.n164 GND.n163 76
R1980 GND.n167 GND.n166 76
R1981 GND.n174 GND.n173 76
R1982 GND.n177 GND.n176 76
R1983 GND.n180 GND.n179 76
R1984 GND.n183 GND.n182 76
R1985 GND.n186 GND.n185 76
R1986 GND.n191 GND.n190 76
R1987 GND.n194 GND.n193 76
R1988 GND.n197 GND.n196 76
R1989 GND.n204 GND.n203 76
R1990 GND.n207 GND.n206 76
R1991 GND.n210 GND.n209 76
R1992 GND.n213 GND.n212 76
R1993 GND.n216 GND.n215 76
R1994 GND.n219 GND.n218 76
R1995 GND.n222 GND.n221 76
R1996 GND.n225 GND.n224 76
R1997 GND.n228 GND.n227 76
R1998 GND.n233 GND.n232 76
R1999 GND.n236 GND.n235 76
R2000 GND.n239 GND.n238 76
R2001 GND.n246 GND.n245 76
R2002 GND.n249 GND.n248 76
R2003 GND.n252 GND.n251 76
R2004 GND.n255 GND.n254 76
R2005 GND.n258 GND.n257 76
R2006 GND.n261 GND.n260 76
R2007 GND.n264 GND.n263 76
R2008 GND.n267 GND.n266 76
R2009 GND.n270 GND.n269 76
R2010 GND.n278 GND.n277 76
R2011 GND.n281 GND.n280 76
R2012 GND.n284 GND.n283 76
R2013 GND.n291 GND.n290 76
R2014 GND.n294 GND.n293 76
R2015 GND.n297 GND.n296 76
R2016 GND.n300 GND.n299 76
R2017 GND.n303 GND.n302 76
R2018 GND.n308 GND.n307 76
R2019 GND.n311 GND.n310 76
R2020 GND.n314 GND.n313 76
R2021 GND.n321 GND.n320 76
R2022 GND.n324 GND.n323 76
R2023 GND.n327 GND.n326 76
R2024 GND.n330 GND.n329 76
R2025 GND.n333 GND.n332 76
R2026 GND.n336 GND.n335 76
R2027 GND.n339 GND.n338 76
R2028 GND.n342 GND.n341 76
R2029 GND.n345 GND.n344 76
R2030 GND.n353 GND.n352 76
R2031 GND.n356 GND.n355 76
R2032 GND.n359 GND.n358 76
R2033 GND.n366 GND.n365 76
R2034 GND.n369 GND.n368 76
R2035 GND.n372 GND.n371 76
R2036 GND.n375 GND.n374 76
R2037 GND.n378 GND.n377 76
R2038 GND.n383 GND.n382 76
R2039 GND.n749 GND.n748 76
R2040 GND.n746 GND.n745 76
R2041 GND.n739 GND.n738 76
R2042 GND.n736 GND.n735 76
R2043 GND.n733 GND.n732 76
R2044 GND.n730 GND.n729 76
R2045 GND.n727 GND.n726 76
R2046 GND.n724 GND.n723 76
R2047 GND.n719 GND.n718 76
R2048 GND.n716 GND.n715 76
R2049 GND.n709 GND.n708 76
R2050 GND.n706 GND.n705 76
R2051 GND.n703 GND.n702 76
R2052 GND.n700 GND.n699 76
R2053 GND.n697 GND.n696 76
R2054 GND.n694 GND.n693 76
R2055 GND.n691 GND.n690 76
R2056 GND.n688 GND.n687 76
R2057 GND.n685 GND.n684 76
R2058 GND.n682 GND.n681 76
R2059 GND.n677 GND.n676 76
R2060 GND.n674 GND.n673 76
R2061 GND.n667 GND.n666 76
R2062 GND.n664 GND.n663 76
R2063 GND.n661 GND.n660 76
R2064 GND.n658 GND.n657 76
R2065 GND.n655 GND.n654 76
R2066 GND.n652 GND.n651 76
R2067 GND.n649 GND.n648 76
R2068 GND.n646 GND.n645 76
R2069 GND.n643 GND.n642 76
R2070 GND.n640 GND.n639 76
R2071 GND.n635 GND.n634 76
R2072 GND.n632 GND.n631 76
R2073 GND.n625 GND.n624 76
R2074 GND.n622 GND.n621 76
R2075 GND.n619 GND.n618 76
R2076 GND.n616 GND.n615 76
R2077 GND.n613 GND.n612 76
R2078 GND.n610 GND.n609 76
R2079 GND.n605 GND.n604 76
R2080 GND.n602 GND.n601 76
R2081 GND.n595 GND.n594 76
R2082 GND.n592 GND.n591 76
R2083 GND.n589 GND.n588 76
R2084 GND.n586 GND.n585 76
R2085 GND.n583 GND.n582 76
R2086 GND.n580 GND.n579 76
R2087 GND.n577 GND.n576 76
R2088 GND.n574 GND.n573 76
R2089 GND.n571 GND.n570 76
R2090 GND.n568 GND.n567 76
R2091 GND.n563 GND.n562 76
R2092 GND.n560 GND.n559 76
R2093 GND.n553 GND.n552 76
R2094 GND.n550 GND.n549 76
R2095 GND.n547 GND.n546 76
R2096 GND.n544 GND.n543 76
R2097 GND.n541 GND.n540 76
R2098 GND.n538 GND.n537 76
R2099 GND.n533 GND.n532 76
R2100 GND.n530 GND.n529 76
R2101 GND.n523 GND.n522 76
R2102 GND.n520 GND.n519 76
R2103 GND.n517 GND.n516 76
R2104 GND.n514 GND.n513 76
R2105 GND.n511 GND.n510 76
R2106 GND.n508 GND.n507 76
R2107 GND.n503 GND.n502 76
R2108 GND.n500 GND.n499 76
R2109 GND.n493 GND.n492 76
R2110 GND.n490 GND.n489 76
R2111 GND.n487 GND.n486 76
R2112 GND.n484 GND.n483 76
R2113 GND.n481 GND.n480 76
R2114 GND.n478 GND.n477 76
R2115 GND.n475 GND.n474 76
R2116 GND.n472 GND.n471 76
R2117 GND.n469 GND.n468 76
R2118 GND.n466 GND.n465 76
R2119 GND.n461 GND.n460 76
R2120 GND.n458 GND.n457 76
R2121 GND.n451 GND.n450 76
R2122 GND.n448 GND.n447 76
R2123 GND.n445 GND.n444 76
R2124 GND.n442 GND.n441 76
R2125 GND.n439 GND.n438 76
R2126 GND.n436 GND.n435 76
R2127 GND.n433 GND.n432 76
R2128 GND.n430 GND.n429 76
R2129 GND.n427 GND.n426 76
R2130 GND.n424 GND.n423 76
R2131 GND.n419 GND.n418 76
R2132 GND.n416 GND.n415 76
R2133 GND.n409 GND.n408 76
R2134 GND.n406 GND.n405 76
R2135 GND.n403 GND.n402 76
R2136 GND.n400 GND.n399 76
R2137 GND.n397 GND.n396 76
R2138 GND.n394 GND.n393 76
R2139 GND.n389 GND.n388 76
R2140 GND.n12 GND.n11 76
R2141 GND.n20 GND.n19 76
R2142 GND.n23 GND.n22 76
R2143 GND.n26 GND.n25 76
R2144 GND.n33 GND.n32 76
R2145 GND.n36 GND.n35 76
R2146 GND.n39 GND.n38 76
R2147 GND.n129 GND.n128 64.552
R2148 GND.n276 GND.n275 64.552
R2149 GND.n351 GND.n350 64.552
R2150 GND.n50 GND.n49 63.835
R2151 GND.n83 GND.n82 63.835
R2152 GND.n17 GND.n16 63.835
R2153 GND.n8 GND.n7 34.942
R2154 GND.n49 GND.n48 28.421
R2155 GND.n82 GND.n81 28.421
R2156 GND.n128 GND.n127 28.421
R2157 GND.n275 GND.n274 28.421
R2158 GND.n350 GND.n349 28.421
R2159 GND.n16 GND.n15 28.421
R2160 GND.n49 GND.n47 25.263
R2161 GND.n82 GND.n80 25.263
R2162 GND.n128 GND.n126 25.263
R2163 GND.n275 GND.n273 25.263
R2164 GND.n350 GND.n348 25.263
R2165 GND.n16 GND.n14 25.263
R2166 GND.n47 GND.n46 24.383
R2167 GND.n80 GND.n79 24.383
R2168 GND.n126 GND.n125 24.383
R2169 GND.n273 GND.n272 24.383
R2170 GND.n348 GND.n347 24.383
R2171 GND.n14 GND.n13 24.383
R2172 GND.n5 GND.n4 14.167
R2173 GND.n4 GND.n2 14.167
R2174 GND.n32 GND.n30 14.167
R2175 GND.n65 GND.n63 14.167
R2176 GND.n98 GND.n96 14.167
R2177 GND.n143 GND.n141 14.167
R2178 GND.n173 GND.n171 14.167
R2179 GND.n203 GND.n201 14.167
R2180 GND.n245 GND.n243 14.167
R2181 GND.n290 GND.n288 14.167
R2182 GND.n320 GND.n318 14.167
R2183 GND.n365 GND.n363 14.167
R2184 GND.n745 GND.n744 14.167
R2185 GND.n715 GND.n714 14.167
R2186 GND.n673 GND.n672 14.167
R2187 GND.n631 GND.n630 14.167
R2188 GND.n601 GND.n600 14.167
R2189 GND.n559 GND.n558 14.167
R2190 GND.n529 GND.n528 14.167
R2191 GND.n499 GND.n498 14.167
R2192 GND.n457 GND.n456 14.167
R2193 GND.n415 GND.n414 14.167
R2194 GND.n388 GND.n387 13.653
R2195 GND.n393 GND.n392 13.653
R2196 GND.n396 GND.n395 13.653
R2197 GND.n399 GND.n398 13.653
R2198 GND.n402 GND.n401 13.653
R2199 GND.n405 GND.n404 13.653
R2200 GND.n408 GND.n407 13.653
R2201 GND.n415 GND.n410 13.653
R2202 GND.n418 GND.n417 13.653
R2203 GND.n423 GND.n420 13.653
R2204 GND.n426 GND.n425 13.653
R2205 GND.n429 GND.n428 13.653
R2206 GND.n432 GND.n431 13.653
R2207 GND.n435 GND.n434 13.653
R2208 GND.n438 GND.n437 13.653
R2209 GND.n441 GND.n440 13.653
R2210 GND.n444 GND.n443 13.653
R2211 GND.n447 GND.n446 13.653
R2212 GND.n450 GND.n449 13.653
R2213 GND.n457 GND.n452 13.653
R2214 GND.n460 GND.n459 13.653
R2215 GND.n465 GND.n462 13.653
R2216 GND.n468 GND.n467 13.653
R2217 GND.n471 GND.n470 13.653
R2218 GND.n474 GND.n473 13.653
R2219 GND.n477 GND.n476 13.653
R2220 GND.n480 GND.n479 13.653
R2221 GND.n483 GND.n482 13.653
R2222 GND.n486 GND.n485 13.653
R2223 GND.n489 GND.n488 13.653
R2224 GND.n492 GND.n491 13.653
R2225 GND.n499 GND.n494 13.653
R2226 GND.n502 GND.n501 13.653
R2227 GND.n507 GND.n506 13.653
R2228 GND.n510 GND.n509 13.653
R2229 GND.n513 GND.n512 13.653
R2230 GND.n516 GND.n515 13.653
R2231 GND.n519 GND.n518 13.653
R2232 GND.n522 GND.n521 13.653
R2233 GND.n529 GND.n524 13.653
R2234 GND.n532 GND.n531 13.653
R2235 GND.n537 GND.n536 13.653
R2236 GND.n540 GND.n539 13.653
R2237 GND.n543 GND.n542 13.653
R2238 GND.n546 GND.n545 13.653
R2239 GND.n549 GND.n548 13.653
R2240 GND.n552 GND.n551 13.653
R2241 GND.n559 GND.n554 13.653
R2242 GND.n562 GND.n561 13.653
R2243 GND.n567 GND.n564 13.653
R2244 GND.n570 GND.n569 13.653
R2245 GND.n573 GND.n572 13.653
R2246 GND.n576 GND.n575 13.653
R2247 GND.n579 GND.n578 13.653
R2248 GND.n582 GND.n581 13.653
R2249 GND.n585 GND.n584 13.653
R2250 GND.n588 GND.n587 13.653
R2251 GND.n591 GND.n590 13.653
R2252 GND.n594 GND.n593 13.653
R2253 GND.n601 GND.n596 13.653
R2254 GND.n604 GND.n603 13.653
R2255 GND.n609 GND.n608 13.653
R2256 GND.n612 GND.n611 13.653
R2257 GND.n615 GND.n614 13.653
R2258 GND.n618 GND.n617 13.653
R2259 GND.n621 GND.n620 13.653
R2260 GND.n624 GND.n623 13.653
R2261 GND.n631 GND.n626 13.653
R2262 GND.n634 GND.n633 13.653
R2263 GND.n639 GND.n636 13.653
R2264 GND.n642 GND.n641 13.653
R2265 GND.n645 GND.n644 13.653
R2266 GND.n648 GND.n647 13.653
R2267 GND.n651 GND.n650 13.653
R2268 GND.n654 GND.n653 13.653
R2269 GND.n657 GND.n656 13.653
R2270 GND.n660 GND.n659 13.653
R2271 GND.n663 GND.n662 13.653
R2272 GND.n666 GND.n665 13.653
R2273 GND.n673 GND.n668 13.653
R2274 GND.n676 GND.n675 13.653
R2275 GND.n681 GND.n678 13.653
R2276 GND.n684 GND.n683 13.653
R2277 GND.n687 GND.n686 13.653
R2278 GND.n690 GND.n689 13.653
R2279 GND.n693 GND.n692 13.653
R2280 GND.n696 GND.n695 13.653
R2281 GND.n699 GND.n698 13.653
R2282 GND.n702 GND.n701 13.653
R2283 GND.n705 GND.n704 13.653
R2284 GND.n708 GND.n707 13.653
R2285 GND.n715 GND.n710 13.653
R2286 GND.n718 GND.n717 13.653
R2287 GND.n723 GND.n722 13.653
R2288 GND.n726 GND.n725 13.653
R2289 GND.n729 GND.n728 13.653
R2290 GND.n732 GND.n731 13.653
R2291 GND.n735 GND.n734 13.653
R2292 GND.n738 GND.n737 13.653
R2293 GND.n745 GND.n740 13.653
R2294 GND.n748 GND.n747 13.653
R2295 GND.n382 GND.n381 13.653
R2296 GND.n377 GND.n376 13.653
R2297 GND.n374 GND.n373 13.653
R2298 GND.n371 GND.n370 13.653
R2299 GND.n368 GND.n367 13.653
R2300 GND.n365 GND.n364 13.653
R2301 GND.n358 GND.n357 13.653
R2302 GND.n355 GND.n354 13.653
R2303 GND.n352 GND.n346 13.653
R2304 GND.n344 GND.n343 13.653
R2305 GND.n341 GND.n340 13.653
R2306 GND.n338 GND.n337 13.653
R2307 GND.n335 GND.n334 13.653
R2308 GND.n332 GND.n331 13.653
R2309 GND.n329 GND.n328 13.653
R2310 GND.n326 GND.n325 13.653
R2311 GND.n323 GND.n322 13.653
R2312 GND.n320 GND.n319 13.653
R2313 GND.n313 GND.n312 13.653
R2314 GND.n310 GND.n309 13.653
R2315 GND.n307 GND.n306 13.653
R2316 GND.n302 GND.n301 13.653
R2317 GND.n299 GND.n298 13.653
R2318 GND.n296 GND.n295 13.653
R2319 GND.n293 GND.n292 13.653
R2320 GND.n290 GND.n289 13.653
R2321 GND.n283 GND.n282 13.653
R2322 GND.n280 GND.n279 13.653
R2323 GND.n277 GND.n271 13.653
R2324 GND.n269 GND.n268 13.653
R2325 GND.n266 GND.n265 13.653
R2326 GND.n263 GND.n262 13.653
R2327 GND.n260 GND.n259 13.653
R2328 GND.n257 GND.n256 13.653
R2329 GND.n254 GND.n253 13.653
R2330 GND.n251 GND.n250 13.653
R2331 GND.n248 GND.n247 13.653
R2332 GND.n245 GND.n244 13.653
R2333 GND.n238 GND.n237 13.653
R2334 GND.n235 GND.n234 13.653
R2335 GND.n232 GND.n229 13.653
R2336 GND.n227 GND.n226 13.653
R2337 GND.n224 GND.n223 13.653
R2338 GND.n221 GND.n220 13.653
R2339 GND.n218 GND.n217 13.653
R2340 GND.n215 GND.n214 13.653
R2341 GND.n212 GND.n211 13.653
R2342 GND.n209 GND.n208 13.653
R2343 GND.n206 GND.n205 13.653
R2344 GND.n203 GND.n202 13.653
R2345 GND.n196 GND.n195 13.653
R2346 GND.n193 GND.n192 13.653
R2347 GND.n190 GND.n189 13.653
R2348 GND.n185 GND.n184 13.653
R2349 GND.n182 GND.n181 13.653
R2350 GND.n179 GND.n178 13.653
R2351 GND.n176 GND.n175 13.653
R2352 GND.n173 GND.n172 13.653
R2353 GND.n166 GND.n165 13.653
R2354 GND.n163 GND.n162 13.653
R2355 GND.n160 GND.n159 13.653
R2356 GND.n155 GND.n154 13.653
R2357 GND.n152 GND.n151 13.653
R2358 GND.n149 GND.n148 13.653
R2359 GND.n146 GND.n145 13.653
R2360 GND.n143 GND.n142 13.653
R2361 GND.n136 GND.n135 13.653
R2362 GND.n133 GND.n132 13.653
R2363 GND.n130 GND.n124 13.653
R2364 GND.n122 GND.n121 13.653
R2365 GND.n119 GND.n118 13.653
R2366 GND.n116 GND.n115 13.653
R2367 GND.n113 GND.n112 13.653
R2368 GND.n110 GND.n109 13.653
R2369 GND.n107 GND.n106 13.653
R2370 GND.n104 GND.n103 13.653
R2371 GND.n101 GND.n100 13.653
R2372 GND.n98 GND.n97 13.653
R2373 GND.n91 GND.n90 13.653
R2374 GND.n88 GND.n87 13.653
R2375 GND.n85 GND.n84 13.653
R2376 GND.n77 GND.n76 13.653
R2377 GND.n74 GND.n73 13.653
R2378 GND.n71 GND.n70 13.653
R2379 GND.n68 GND.n67 13.653
R2380 GND.n65 GND.n64 13.653
R2381 GND.n58 GND.n57 13.653
R2382 GND.n55 GND.n54 13.653
R2383 GND.n52 GND.n51 13.653
R2384 GND.n44 GND.n43 13.653
R2385 GND.n41 GND.n40 13.653
R2386 GND.n5 GND.n0 13.653
R2387 GND.n4 GND.n3 13.653
R2388 GND.n2 GND.n1 13.653
R2389 GND.n11 GND.n10 13.653
R2390 GND.n19 GND.n18 13.653
R2391 GND.n22 GND.n21 13.653
R2392 GND.n25 GND.n24 13.653
R2393 GND.n32 GND.n31 13.653
R2394 GND.n35 GND.n34 13.653
R2395 GND.n38 GND.n37 13.653
R2396 GND.n30 GND.n29 7.312
R2397 GND.n63 GND.n62 7.312
R2398 GND.n414 GND.n413 7.312
R2399 GND.n456 GND.n455 7.312
R2400 GND.n498 GND.n497 7.312
R2401 GND.n528 GND.n527 7.312
R2402 GND.n558 GND.n557 7.312
R2403 GND.n600 GND.n599 7.312
R2404 GND.n630 GND.n629 7.312
R2405 GND.n672 GND.n671 7.312
R2406 GND.n714 GND.n713 7.312
R2407 GND.n744 GND.n743 7.312
R2408 GND.n363 GND.n362 7.312
R2409 GND.n318 GND.n317 7.312
R2410 GND.n288 GND.n287 7.312
R2411 GND.n243 GND.n242 7.312
R2412 GND.n201 GND.n200 7.312
R2413 GND.n171 GND.n170 7.312
R2414 GND.n141 GND.n140 7.312
R2415 GND.n96 GND.n95 7.312
R2416 GND.n7 GND.n6 7.084
R2417 GND.n7 GND.n5 6.475
R2418 GND.n19 GND.n17 3.935
R2419 GND.n52 GND.n50 3.935
R2420 GND.n85 GND.n83 3.935
R2421 GND.n160 GND.n158 3.935
R2422 GND.n190 GND.n188 3.935
R2423 GND.n307 GND.n305 3.935
R2424 GND.n382 GND.n380 3.935
R2425 GND.n723 GND.n721 3.935
R2426 GND.n609 GND.n607 3.935
R2427 GND.n537 GND.n535 3.935
R2428 GND.n507 GND.n505 3.935
R2429 GND.n393 GND.n391 3.935
R2430 GND.n385 GND.n384 0.596
R2431 GND.n33 GND.n26 0.29
R2432 GND.n66 GND.n59 0.29
R2433 GND.n99 GND.n92 0.29
R2434 GND.n144 GND.n137 0.29
R2435 GND.n174 GND.n167 0.29
R2436 GND.n204 GND.n197 0.29
R2437 GND.n246 GND.n239 0.29
R2438 GND.n291 GND.n284 0.29
R2439 GND.n321 GND.n314 0.29
R2440 GND.n366 GND.n359 0.29
R2441 GND.n746 GND.n739 0.29
R2442 GND.n716 GND.n709 0.29
R2443 GND.n674 GND.n667 0.29
R2444 GND.n632 GND.n625 0.29
R2445 GND.n602 GND.n595 0.29
R2446 GND.n560 GND.n553 0.29
R2447 GND.n530 GND.n523 0.29
R2448 GND.n500 GND.n493 0.29
R2449 GND.n458 GND.n451 0.29
R2450 GND.n416 GND.n409 0.29
R2451 GND.n386 GND 0.207
R2452 GND.n117 GND.n114 0.197
R2453 GND.n222 GND.n219 0.197
R2454 GND.n264 GND.n261 0.197
R2455 GND.n339 GND.n336 0.197
R2456 GND.n694 GND.n691 0.197
R2457 GND.n652 GND.n649 0.197
R2458 GND.n580 GND.n577 0.197
R2459 GND.n478 GND.n475 0.197
R2460 GND.n436 GND.n433 0.197
R2461 GND.n130 GND.n129 0.196
R2462 GND.n232 GND.n231 0.196
R2463 GND.n277 GND.n276 0.196
R2464 GND.n352 GND.n351 0.196
R2465 GND.n681 GND.n680 0.196
R2466 GND.n639 GND.n638 0.196
R2467 GND.n567 GND.n566 0.196
R2468 GND.n465 GND.n464 0.196
R2469 GND.n423 GND.n422 0.196
R2470 GND.n12 GND.n9 0.181
R2471 GND.n45 GND.n42 0.181
R2472 GND.n78 GND.n75 0.181
R2473 GND.n156 GND.n153 0.181
R2474 GND.n186 GND.n183 0.181
R2475 GND.n303 GND.n300 0.181
R2476 GND.n378 GND.n375 0.181
R2477 GND.n730 GND.n727 0.181
R2478 GND.n616 GND.n613 0.181
R2479 GND.n544 GND.n541 0.181
R2480 GND.n514 GND.n511 0.181
R2481 GND.n400 GND.n397 0.181
R2482 GND.n9 GND.n8 0.145
R2483 GND.n20 GND.n12 0.145
R2484 GND.n23 GND.n20 0.145
R2485 GND.n26 GND.n23 0.145
R2486 GND.n36 GND.n33 0.145
R2487 GND.n39 GND.n36 0.145
R2488 GND.n42 GND.n39 0.145
R2489 GND.n53 GND.n45 0.145
R2490 GND.n56 GND.n53 0.145
R2491 GND.n59 GND.n56 0.145
R2492 GND.n69 GND.n66 0.145
R2493 GND.n72 GND.n69 0.145
R2494 GND.n75 GND.n72 0.145
R2495 GND.n86 GND.n78 0.145
R2496 GND.n89 GND.n86 0.145
R2497 GND.n92 GND.n89 0.145
R2498 GND.n102 GND.n99 0.145
R2499 GND.n105 GND.n102 0.145
R2500 GND.n108 GND.n105 0.145
R2501 GND.n111 GND.n108 0.145
R2502 GND.n114 GND.n111 0.145
R2503 GND.n120 GND.n117 0.145
R2504 GND.n123 GND.n120 0.145
R2505 GND.n131 GND.n123 0.145
R2506 GND.n134 GND.n131 0.145
R2507 GND.n137 GND.n134 0.145
R2508 GND.n147 GND.n144 0.145
R2509 GND.n150 GND.n147 0.145
R2510 GND.n153 GND.n150 0.145
R2511 GND.n161 GND.n156 0.145
R2512 GND.n164 GND.n161 0.145
R2513 GND.n167 GND.n164 0.145
R2514 GND.n177 GND.n174 0.145
R2515 GND.n180 GND.n177 0.145
R2516 GND.n183 GND.n180 0.145
R2517 GND.n191 GND.n186 0.145
R2518 GND.n194 GND.n191 0.145
R2519 GND.n197 GND.n194 0.145
R2520 GND.n207 GND.n204 0.145
R2521 GND.n210 GND.n207 0.145
R2522 GND.n213 GND.n210 0.145
R2523 GND.n216 GND.n213 0.145
R2524 GND.n219 GND.n216 0.145
R2525 GND.n225 GND.n222 0.145
R2526 GND.n228 GND.n225 0.145
R2527 GND.n233 GND.n228 0.145
R2528 GND.n236 GND.n233 0.145
R2529 GND.n239 GND.n236 0.145
R2530 GND.n249 GND.n246 0.145
R2531 GND.n252 GND.n249 0.145
R2532 GND.n255 GND.n252 0.145
R2533 GND.n258 GND.n255 0.145
R2534 GND.n261 GND.n258 0.145
R2535 GND.n267 GND.n264 0.145
R2536 GND.n270 GND.n267 0.145
R2537 GND.n278 GND.n270 0.145
R2538 GND.n281 GND.n278 0.145
R2539 GND.n284 GND.n281 0.145
R2540 GND.n294 GND.n291 0.145
R2541 GND.n297 GND.n294 0.145
R2542 GND.n300 GND.n297 0.145
R2543 GND.n308 GND.n303 0.145
R2544 GND.n311 GND.n308 0.145
R2545 GND.n314 GND.n311 0.145
R2546 GND.n324 GND.n321 0.145
R2547 GND.n327 GND.n324 0.145
R2548 GND.n330 GND.n327 0.145
R2549 GND.n333 GND.n330 0.145
R2550 GND.n336 GND.n333 0.145
R2551 GND.n342 GND.n339 0.145
R2552 GND.n345 GND.n342 0.145
R2553 GND.n353 GND.n345 0.145
R2554 GND.n356 GND.n353 0.145
R2555 GND.n359 GND.n356 0.145
R2556 GND.n369 GND.n366 0.145
R2557 GND.n372 GND.n369 0.145
R2558 GND.n375 GND.n372 0.145
R2559 GND.n383 GND.n378 0.145
R2560 GND.n749 GND.n746 0.145
R2561 GND.n739 GND.n736 0.145
R2562 GND.n736 GND.n733 0.145
R2563 GND.n733 GND.n730 0.145
R2564 GND.n727 GND.n724 0.145
R2565 GND.n724 GND.n719 0.145
R2566 GND.n719 GND.n716 0.145
R2567 GND.n709 GND.n706 0.145
R2568 GND.n706 GND.n703 0.145
R2569 GND.n703 GND.n700 0.145
R2570 GND.n700 GND.n697 0.145
R2571 GND.n697 GND.n694 0.145
R2572 GND.n691 GND.n688 0.145
R2573 GND.n688 GND.n685 0.145
R2574 GND.n685 GND.n682 0.145
R2575 GND.n682 GND.n677 0.145
R2576 GND.n677 GND.n674 0.145
R2577 GND.n667 GND.n664 0.145
R2578 GND.n664 GND.n661 0.145
R2579 GND.n661 GND.n658 0.145
R2580 GND.n658 GND.n655 0.145
R2581 GND.n655 GND.n652 0.145
R2582 GND.n649 GND.n646 0.145
R2583 GND.n646 GND.n643 0.145
R2584 GND.n643 GND.n640 0.145
R2585 GND.n640 GND.n635 0.145
R2586 GND.n635 GND.n632 0.145
R2587 GND.n625 GND.n622 0.145
R2588 GND.n622 GND.n619 0.145
R2589 GND.n619 GND.n616 0.145
R2590 GND.n613 GND.n610 0.145
R2591 GND.n610 GND.n605 0.145
R2592 GND.n605 GND.n602 0.145
R2593 GND.n595 GND.n592 0.145
R2594 GND.n592 GND.n589 0.145
R2595 GND.n589 GND.n586 0.145
R2596 GND.n586 GND.n583 0.145
R2597 GND.n583 GND.n580 0.145
R2598 GND.n577 GND.n574 0.145
R2599 GND.n574 GND.n571 0.145
R2600 GND.n571 GND.n568 0.145
R2601 GND.n568 GND.n563 0.145
R2602 GND.n563 GND.n560 0.145
R2603 GND.n553 GND.n550 0.145
R2604 GND.n550 GND.n547 0.145
R2605 GND.n547 GND.n544 0.145
R2606 GND.n541 GND.n538 0.145
R2607 GND.n538 GND.n533 0.145
R2608 GND.n533 GND.n530 0.145
R2609 GND.n523 GND.n520 0.145
R2610 GND.n520 GND.n517 0.145
R2611 GND.n517 GND.n514 0.145
R2612 GND.n511 GND.n508 0.145
R2613 GND.n508 GND.n503 0.145
R2614 GND.n503 GND.n500 0.145
R2615 GND.n493 GND.n490 0.145
R2616 GND.n490 GND.n487 0.145
R2617 GND.n487 GND.n484 0.145
R2618 GND.n484 GND.n481 0.145
R2619 GND.n481 GND.n478 0.145
R2620 GND.n475 GND.n472 0.145
R2621 GND.n472 GND.n469 0.145
R2622 GND.n469 GND.n466 0.145
R2623 GND.n466 GND.n461 0.145
R2624 GND.n461 GND.n458 0.145
R2625 GND.n451 GND.n448 0.145
R2626 GND.n448 GND.n445 0.145
R2627 GND.n445 GND.n442 0.145
R2628 GND.n442 GND.n439 0.145
R2629 GND.n439 GND.n436 0.145
R2630 GND.n433 GND.n430 0.145
R2631 GND.n430 GND.n427 0.145
R2632 GND.n427 GND.n424 0.145
R2633 GND.n424 GND.n419 0.145
R2634 GND.n419 GND.n416 0.145
R2635 GND.n409 GND.n406 0.145
R2636 GND.n406 GND.n403 0.145
R2637 GND.n403 GND.n400 0.145
R2638 GND.n397 GND.n394 0.145
R2639 GND.n394 GND.n389 0.145
R2640 GND.n389 GND.n386 0.145
R2641 GND GND.n749 0.082
R2642 GND GND.n383 0.062
R2643 a_1265_989.n2 a_1265_989.t12 454.685
R2644 a_1265_989.n4 a_1265_989.t5 454.685
R2645 a_1265_989.n0 a_1265_989.t9 454.685
R2646 a_1265_989.n2 a_1265_989.t7 428.979
R2647 a_1265_989.n4 a_1265_989.t11 428.979
R2648 a_1265_989.n0 a_1265_989.t10 428.979
R2649 a_1265_989.n3 a_1265_989.t6 264.512
R2650 a_1265_989.n5 a_1265_989.t8 264.512
R2651 a_1265_989.n1 a_1265_989.t13 264.512
R2652 a_1265_989.n12 a_1265_989.n11 237.145
R2653 a_1265_989.n14 a_1265_989.n12 125.947
R2654 a_1265_989.n7 a_1265_989.n1 81.396
R2655 a_1265_989.n6 a_1265_989.n5 79.491
R2656 a_1265_989.n14 a_1265_989.n13 76.002
R2657 a_1265_989.n6 a_1265_989.n3 76
R2658 a_1265_989.n12 a_1265_989.n7 76
R2659 a_1265_989.n3 a_1265_989.n2 71.894
R2660 a_1265_989.n5 a_1265_989.n4 71.894
R2661 a_1265_989.n1 a_1265_989.n0 71.894
R2662 a_1265_989.n11 a_1265_989.n10 30
R2663 a_1265_989.n9 a_1265_989.n8 24.383
R2664 a_1265_989.n11 a_1265_989.n9 23.684
R2665 a_1265_989.n13 a_1265_989.t4 14.282
R2666 a_1265_989.n13 a_1265_989.t0 14.282
R2667 a_1265_989.n15 a_1265_989.t2 14.282
R2668 a_1265_989.t3 a_1265_989.n15 14.282
R2669 a_1265_989.n15 a_1265_989.n14 12.848
R2670 a_1265_989.n7 a_1265_989.n6 2.947
R2671 a_343_411.n1 a_343_411.t7 480.392
R2672 a_343_411.n3 a_343_411.t9 472.359
R2673 a_343_411.n1 a_343_411.t10 403.272
R2674 a_343_411.n3 a_343_411.t12 384.527
R2675 a_343_411.n2 a_343_411.t8 336.586
R2676 a_343_411.n4 a_343_411.t11 294.278
R2677 a_343_411.n10 a_343_411.n9 265.87
R2678 a_343_411.n11 a_343_411.n10 117.354
R2679 a_343_411.n5 a_343_411.n2 83.304
R2680 a_343_411.n5 a_343_411.n4 80.032
R2681 a_343_411.n13 a_343_411.n12 79.232
R2682 a_343_411.n10 a_343_411.n5 76
R2683 a_343_411.n13 a_343_411.n11 63.152
R2684 a_343_411.n4 a_343_411.n3 56.954
R2685 a_343_411.n2 a_343_411.n1 45.341
R2686 a_343_411.n9 a_343_411.n8 30
R2687 a_343_411.n7 a_343_411.n6 24.383
R2688 a_343_411.n9 a_343_411.n7 23.684
R2689 a_343_411.n11 a_343_411.n0 16.08
R2690 a_343_411.n14 a_343_411.n13 16.078
R2691 a_343_411.n0 a_343_411.t4 14.282
R2692 a_343_411.n0 a_343_411.t5 14.282
R2693 a_343_411.n12 a_343_411.t3 14.282
R2694 a_343_411.n12 a_343_411.t0 14.282
R2695 a_343_411.t2 a_343_411.n14 14.282
R2696 a_343_411.n14 a_343_411.t1 14.282
R2697 a_11033_989.n2 a_11033_989.t8 454.685
R2698 a_11033_989.n4 a_11033_989.t13 454.685
R2699 a_11033_989.n0 a_11033_989.t5 454.685
R2700 a_11033_989.n2 a_11033_989.t7 428.979
R2701 a_11033_989.n4 a_11033_989.t9 428.979
R2702 a_11033_989.n0 a_11033_989.t11 428.979
R2703 a_11033_989.n3 a_11033_989.t12 264.512
R2704 a_11033_989.n5 a_11033_989.t10 264.512
R2705 a_11033_989.n1 a_11033_989.t6 264.512
R2706 a_11033_989.n12 a_11033_989.n11 237.145
R2707 a_11033_989.n14 a_11033_989.n12 125.947
R2708 a_11033_989.n7 a_11033_989.n1 81.396
R2709 a_11033_989.n6 a_11033_989.n5 79.491
R2710 a_11033_989.n14 a_11033_989.n13 76.002
R2711 a_11033_989.n6 a_11033_989.n3 76
R2712 a_11033_989.n12 a_11033_989.n7 76
R2713 a_11033_989.n3 a_11033_989.n2 71.894
R2714 a_11033_989.n5 a_11033_989.n4 71.894
R2715 a_11033_989.n1 a_11033_989.n0 71.894
R2716 a_11033_989.n11 a_11033_989.n10 30
R2717 a_11033_989.n9 a_11033_989.n8 24.383
R2718 a_11033_989.n11 a_11033_989.n9 23.684
R2719 a_11033_989.n13 a_11033_989.t1 14.282
R2720 a_11033_989.n13 a_11033_989.t0 14.282
R2721 a_11033_989.t4 a_11033_989.n15 14.282
R2722 a_11033_989.n15 a_11033_989.t3 14.282
R2723 a_11033_989.n15 a_11033_989.n14 12.848
R2724 a_11033_989.n7 a_11033_989.n6 2.947
R2725 a_5101_1050.n5 a_5101_1050.t7 512.525
R2726 a_5101_1050.n3 a_5101_1050.t6 512.525
R2727 a_5101_1050.n5 a_5101_1050.t5 371.139
R2728 a_5101_1050.n3 a_5101_1050.t8 371.139
R2729 a_5101_1050.n4 a_5101_1050.t10 234.562
R2730 a_5101_1050.n6 a_5101_1050.t9 234.204
R2731 a_5101_1050.n6 a_5101_1050.n5 216.178
R2732 a_5101_1050.n4 a_5101_1050.n3 215.819
R2733 a_5101_1050.n8 a_5101_1050.n2 205.605
R2734 a_5101_1050.n10 a_5101_1050.n8 164.008
R2735 a_5101_1050.n7 a_5101_1050.n4 79.488
R2736 a_5101_1050.n8 a_5101_1050.n7 77.314
R2737 a_5101_1050.n2 a_5101_1050.n1 76.002
R2738 a_5101_1050.n7 a_5101_1050.n6 76
R2739 a_5101_1050.n10 a_5101_1050.n9 15.218
R2740 a_5101_1050.n0 a_5101_1050.t2 14.282
R2741 a_5101_1050.n0 a_5101_1050.t1 14.282
R2742 a_5101_1050.n1 a_5101_1050.t0 14.282
R2743 a_5101_1050.n1 a_5101_1050.t4 14.282
R2744 a_5101_1050.n2 a_5101_1050.n0 12.85
R2745 a_5101_1050.n11 a_5101_1050.n10 12.014
R2746 a_5227_411.n0 a_5227_411.t9 480.392
R2747 a_5227_411.n2 a_5227_411.t8 472.359
R2748 a_5227_411.n0 a_5227_411.t12 403.272
R2749 a_5227_411.n2 a_5227_411.t11 384.527
R2750 a_5227_411.n1 a_5227_411.t10 336.586
R2751 a_5227_411.n3 a_5227_411.t7 294.278
R2752 a_5227_411.n9 a_5227_411.n8 265.87
R2753 a_5227_411.n13 a_5227_411.n9 117.354
R2754 a_5227_411.n4 a_5227_411.n1 83.304
R2755 a_5227_411.n4 a_5227_411.n3 80.032
R2756 a_5227_411.n12 a_5227_411.n11 79.232
R2757 a_5227_411.n9 a_5227_411.n4 76
R2758 a_5227_411.n13 a_5227_411.n12 63.152
R2759 a_5227_411.n3 a_5227_411.n2 56.954
R2760 a_5227_411.n1 a_5227_411.n0 45.341
R2761 a_5227_411.n8 a_5227_411.n7 30
R2762 a_5227_411.n6 a_5227_411.n5 24.383
R2763 a_5227_411.n8 a_5227_411.n6 23.684
R2764 a_5227_411.n12 a_5227_411.n10 16.08
R2765 a_5227_411.n14 a_5227_411.n13 16.078
R2766 a_5227_411.n10 a_5227_411.t6 14.282
R2767 a_5227_411.n10 a_5227_411.t5 14.282
R2768 a_5227_411.n11 a_5227_411.t3 14.282
R2769 a_5227_411.n11 a_5227_411.t4 14.282
R2770 a_5227_411.n14 a_5227_411.t1 14.282
R2771 a_5227_411.t2 a_5227_411.n14 14.282
R2772 a_1905_1050.n1 a_1905_1050.t7 480.392
R2773 a_1905_1050.n1 a_1905_1050.t9 403.272
R2774 a_1905_1050.n2 a_1905_1050.t8 230.374
R2775 a_1905_1050.n8 a_1905_1050.n7 223.905
R2776 a_1905_1050.n7 a_1905_1050.n6 159.998
R2777 a_1905_1050.n7 a_1905_1050.n2 153.315
R2778 a_1905_1050.n2 a_1905_1050.n1 151.553
R2779 a_1905_1050.n10 a_1905_1050.n9 79.232
R2780 a_1905_1050.n10 a_1905_1050.n8 63.152
R2781 a_1905_1050.n6 a_1905_1050.n5 30
R2782 a_1905_1050.n4 a_1905_1050.n3 24.383
R2783 a_1905_1050.n6 a_1905_1050.n4 23.684
R2784 a_1905_1050.n8 a_1905_1050.n0 16.08
R2785 a_1905_1050.n11 a_1905_1050.n10 16.078
R2786 a_1905_1050.n0 a_1905_1050.t6 14.282
R2787 a_1905_1050.n0 a_1905_1050.t5 14.282
R2788 a_1905_1050.n9 a_1905_1050.t3 14.282
R2789 a_1905_1050.n9 a_1905_1050.t2 14.282
R2790 a_1905_1050.t1 a_1905_1050.n11 14.282
R2791 a_1905_1050.n11 a_1905_1050.t0 14.282
R2792 a_11673_1050.n1 a_11673_1050.t8 480.392
R2793 a_11673_1050.n1 a_11673_1050.t9 403.272
R2794 a_11673_1050.n2 a_11673_1050.t7 230.374
R2795 a_11673_1050.n8 a_11673_1050.n7 223.905
R2796 a_11673_1050.n7 a_11673_1050.n6 159.998
R2797 a_11673_1050.n7 a_11673_1050.n2 153.315
R2798 a_11673_1050.n2 a_11673_1050.n1 151.553
R2799 a_11673_1050.n10 a_11673_1050.n9 79.232
R2800 a_11673_1050.n10 a_11673_1050.n8 63.152
R2801 a_11673_1050.n6 a_11673_1050.n5 30
R2802 a_11673_1050.n4 a_11673_1050.n3 24.383
R2803 a_11673_1050.n6 a_11673_1050.n4 23.684
R2804 a_11673_1050.n8 a_11673_1050.n0 16.08
R2805 a_11673_1050.n11 a_11673_1050.n10 16.078
R2806 a_11673_1050.n0 a_11673_1050.t5 14.282
R2807 a_11673_1050.n0 a_11673_1050.t4 14.282
R2808 a_11673_1050.n9 a_11673_1050.t2 14.282
R2809 a_11673_1050.n9 a_11673_1050.t3 14.282
R2810 a_11673_1050.t1 a_11673_1050.n11 14.282
R2811 a_11673_1050.n11 a_11673_1050.t0 14.282
R2812 QN.n16 QN.n15 216.728
R2813 QN.n16 QN.n2 126.664
R2814 QN.n11 QN.n10 98.501
R2815 QN.n11 QN.n6 96.417
R2816 QN.n14 QN.n12 80.526
R2817 QN.n15 QN.n11 78.403
R2818 QN.n17 QN.n16 76
R2819 QN.n2 QN.n1 75.271
R2820 QN.n6 QN.n5 30
R2821 QN.n10 QN.n9 30
R2822 QN.n14 QN.n13 30
R2823 QN.n4 QN.n3 24.383
R2824 QN.n8 QN.n7 24.383
R2825 QN.n6 QN.n4 23.684
R2826 QN.n10 QN.n8 23.684
R2827 QN.n15 QN.n14 20.417
R2828 QN.n0 QN.t4 14.282
R2829 QN.n0 QN.t5 14.282
R2830 QN.n1 QN.t1 14.282
R2831 QN.n1 QN.t0 14.282
R2832 QN.n2 QN.n0 12.119
R2833 QN.n17 QN 0.046
R2834 a_15533_1051.n4 a_15533_1051.n3 196.002
R2835 a_15533_1051.n2 a_15533_1051.t5 89.553
R2836 a_15533_1051.n4 a_15533_1051.n0 75.271
R2837 a_15533_1051.n3 a_15533_1051.n2 75.214
R2838 a_15533_1051.n5 a_15533_1051.n4 36.519
R2839 a_15533_1051.n3 a_15533_1051.t2 14.338
R2840 a_15533_1051.n1 a_15533_1051.t4 14.282
R2841 a_15533_1051.n1 a_15533_1051.t3 14.282
R2842 a_15533_1051.n0 a_15533_1051.t7 14.282
R2843 a_15533_1051.n0 a_15533_1051.t6 14.282
R2844 a_15533_1051.t1 a_15533_1051.n5 14.282
R2845 a_15533_1051.n5 a_15533_1051.t0 14.282
R2846 a_15533_1051.n2 a_15533_1051.n1 12.119
R2847 a_2000_210.n10 a_2000_210.n8 82.852
R2848 a_2000_210.n7 a_2000_210.n6 32.833
R2849 a_2000_210.n8 a_2000_210.t1 32.416
R2850 a_2000_210.n10 a_2000_210.n9 27.2
R2851 a_2000_210.n11 a_2000_210.n0 23.498
R2852 a_2000_210.n3 a_2000_210.n2 23.284
R2853 a_2000_210.n11 a_2000_210.n10 22.4
R2854 a_2000_210.n7 a_2000_210.n4 19.017
R2855 a_2000_210.n6 a_2000_210.n5 13.494
R2856 a_2000_210.t1 a_2000_210.n1 7.04
R2857 a_2000_210.t1 a_2000_210.n3 5.727
R2858 a_2000_210.n8 a_2000_210.n7 1.435
R2859 a_10525_103.n4 a_10525_103.n3 19.724
R2860 a_10525_103.t0 a_10525_103.n5 11.595
R2861 a_10525_103.t0 a_10525_103.n4 9.207
R2862 a_10525_103.n2 a_10525_103.n0 8.543
R2863 a_10525_103.t0 a_10525_103.n2 3.034
R2864 a_10525_103.n2 a_10525_103.n1 0.443
R2865 a_10806_210.n12 a_10806_210.n10 82.852
R2866 a_10806_210.n13 a_10806_210.n0 49.6
R2867 a_10806_210.t1 a_10806_210.n2 46.91
R2868 a_10806_210.n7 a_10806_210.n5 34.805
R2869 a_10806_210.n7 a_10806_210.n6 32.622
R2870 a_10806_210.n10 a_10806_210.t1 32.416
R2871 a_10806_210.n12 a_10806_210.n11 27.2
R2872 a_10806_210.n13 a_10806_210.n12 22.4
R2873 a_10806_210.n9 a_10806_210.n7 19.017
R2874 a_10806_210.n2 a_10806_210.n1 17.006
R2875 a_10806_210.n5 a_10806_210.n4 7.5
R2876 a_10806_210.n9 a_10806_210.n8 7.5
R2877 a_10806_210.t1 a_10806_210.n3 7.04
R2878 a_10806_210.n10 a_10806_210.n9 1.435
R2879 a_12470_101.n12 a_12470_101.n11 26.811
R2880 a_12470_101.n6 a_12470_101.n5 24.977
R2881 a_12470_101.n2 a_12470_101.n1 24.877
R2882 a_12470_101.t0 a_12470_101.n2 12.677
R2883 a_12470_101.t0 a_12470_101.n3 11.595
R2884 a_12470_101.t1 a_12470_101.n8 8.137
R2885 a_12470_101.t0 a_12470_101.n4 7.273
R2886 a_12470_101.t0 a_12470_101.n0 6.109
R2887 a_12470_101.t1 a_12470_101.n7 4.864
R2888 a_12470_101.t0 a_12470_101.n12 2.074
R2889 a_12470_101.n7 a_12470_101.n6 1.13
R2890 a_12470_101.n12 a_12470_101.t1 0.937
R2891 a_12470_101.t1 a_12470_101.n10 0.804
R2892 a_12470_101.n10 a_12470_101.n9 0.136
R2893 D.n5 D.t1 480.392
R2894 D.n2 D.t0 480.392
R2895 D.n0 D.t5 480.392
R2896 D.n5 D.t4 403.272
R2897 D.n2 D.t6 403.272
R2898 D.n0 D.t8 403.272
R2899 D.n6 D.n5 204.659
R2900 D.n3 D.n2 204.659
R2901 D.n1 D.n0 204.659
R2902 D.n6 D.t2 183.422
R2903 D.n3 D.t7 183.422
R2904 D.n1 D.t3 183.422
R2905 D.n4 D.n1 93.91
R2906 D.n4 D.n3 76
R2907 D.n7 D.n6 76
R2908 D.n7 D.n4 17.91
R2909 D.n7 D 0.046
R2910 a_217_1050.n2 a_217_1050.t7 512.525
R2911 a_217_1050.n0 a_217_1050.t10 512.525
R2912 a_217_1050.n2 a_217_1050.t9 371.139
R2913 a_217_1050.n0 a_217_1050.t6 371.139
R2914 a_217_1050.n1 a_217_1050.t8 234.562
R2915 a_217_1050.n3 a_217_1050.t5 234.204
R2916 a_217_1050.n3 a_217_1050.n2 216.178
R2917 a_217_1050.n1 a_217_1050.n0 215.819
R2918 a_217_1050.n11 a_217_1050.n9 205.605
R2919 a_217_1050.n9 a_217_1050.n8 157.486
R2920 a_217_1050.n4 a_217_1050.n1 79.488
R2921 a_217_1050.n9 a_217_1050.n4 77.314
R2922 a_217_1050.n11 a_217_1050.n10 76.002
R2923 a_217_1050.n4 a_217_1050.n3 76
R2924 a_217_1050.n8 a_217_1050.n7 30
R2925 a_217_1050.n6 a_217_1050.n5 24.383
R2926 a_217_1050.n8 a_217_1050.n6 23.684
R2927 a_217_1050.n10 a_217_1050.t4 14.282
R2928 a_217_1050.n10 a_217_1050.t3 14.282
R2929 a_217_1050.t1 a_217_1050.n12 14.282
R2930 a_217_1050.n12 a_217_1050.t0 14.282
R2931 a_217_1050.n12 a_217_1050.n11 12.848
R2932 a_15430_101.t0 a_15430_101.n0 34.602
R2933 a_15430_101.t0 a_15430_101.n1 2.138
R2934 a_10111_411.n2 a_10111_411.t12 480.392
R2935 a_10111_411.n4 a_10111_411.t9 472.359
R2936 a_10111_411.n2 a_10111_411.t8 403.272
R2937 a_10111_411.n4 a_10111_411.t7 384.527
R2938 a_10111_411.n3 a_10111_411.t11 336.586
R2939 a_10111_411.n5 a_10111_411.t10 294.278
R2940 a_10111_411.n10 a_10111_411.n9 281.393
R2941 a_10111_411.n11 a_10111_411.n10 117.354
R2942 a_10111_411.n6 a_10111_411.n3 83.304
R2943 a_10111_411.n6 a_10111_411.n5 80.032
R2944 a_10111_411.n13 a_10111_411.n12 79.231
R2945 a_10111_411.n10 a_10111_411.n6 76
R2946 a_10111_411.n12 a_10111_411.n11 63.152
R2947 a_10111_411.n5 a_10111_411.n4 56.954
R2948 a_10111_411.n3 a_10111_411.n2 45.341
R2949 a_10111_411.n9 a_10111_411.n8 22.578
R2950 a_10111_411.n11 a_10111_411.n1 16.08
R2951 a_10111_411.n12 a_10111_411.n0 16.08
R2952 a_10111_411.n1 a_10111_411.t6 14.282
R2953 a_10111_411.n1 a_10111_411.t5 14.282
R2954 a_10111_411.n0 a_10111_411.t2 14.282
R2955 a_10111_411.n0 a_10111_411.t3 14.282
R2956 a_10111_411.n13 a_10111_411.t0 14.282
R2957 a_10111_411.t1 a_10111_411.n13 14.282
R2958 a_10111_411.n9 a_10111_411.n7 8.58
R2959 a_6789_1050.n0 a_6789_1050.t8 480.392
R2960 a_6789_1050.n0 a_6789_1050.t7 403.272
R2961 a_6789_1050.n1 a_6789_1050.t9 230.374
R2962 a_6789_1050.n7 a_6789_1050.n3 223.905
R2963 a_6789_1050.n3 a_6789_1050.n2 181.737
R2964 a_6789_1050.n3 a_6789_1050.n1 153.315
R2965 a_6789_1050.n1 a_6789_1050.n0 151.553
R2966 a_6789_1050.n6 a_6789_1050.n5 79.232
R2967 a_6789_1050.n7 a_6789_1050.n6 63.152
R2968 a_6789_1050.n6 a_6789_1050.n4 16.08
R2969 a_6789_1050.n8 a_6789_1050.n7 16.078
R2970 a_6789_1050.n4 a_6789_1050.t4 14.282
R2971 a_6789_1050.n4 a_6789_1050.t3 14.282
R2972 a_6789_1050.n5 a_6789_1050.t6 14.282
R2973 a_6789_1050.n5 a_6789_1050.t5 14.282
R2974 a_6789_1050.n8 a_6789_1050.t1 14.282
R2975 a_6789_1050.t2 a_6789_1050.n8 14.282
R2976 a_1038_210.n10 a_1038_210.n8 82.852
R2977 a_1038_210.n7 a_1038_210.n6 32.833
R2978 a_1038_210.n8 a_1038_210.t1 32.416
R2979 a_1038_210.n10 a_1038_210.n9 27.2
R2980 a_1038_210.n11 a_1038_210.n0 23.498
R2981 a_1038_210.n3 a_1038_210.n2 23.284
R2982 a_1038_210.n11 a_1038_210.n10 22.4
R2983 a_1038_210.n7 a_1038_210.n4 19.017
R2984 a_1038_210.n6 a_1038_210.n5 13.494
R2985 a_1038_210.t1 a_1038_210.n1 7.04
R2986 a_1038_210.t1 a_1038_210.n3 5.727
R2987 a_1038_210.n8 a_1038_210.n7 1.435
R2988 a_14062_210.n10 a_14062_210.n8 82.852
R2989 a_14062_210.n7 a_14062_210.n6 32.833
R2990 a_14062_210.n8 a_14062_210.t1 32.416
R2991 a_14062_210.n10 a_14062_210.n9 27.2
R2992 a_14062_210.n11 a_14062_210.n0 23.498
R2993 a_14062_210.n3 a_14062_210.n2 23.284
R2994 a_14062_210.n11 a_14062_210.n10 22.4
R2995 a_14062_210.n7 a_14062_210.n4 19.017
R2996 a_14062_210.n6 a_14062_210.n5 13.494
R2997 a_14062_210.t1 a_14062_210.n1 7.04
R2998 a_14062_210.t1 a_14062_210.n3 5.727
R2999 a_14062_210.n8 a_14062_210.n7 1.435
R3000 a_11768_210.n10 a_11768_210.n8 82.852
R3001 a_11768_210.n11 a_11768_210.n0 49.6
R3002 a_11768_210.n7 a_11768_210.n6 32.833
R3003 a_11768_210.n8 a_11768_210.t1 32.416
R3004 a_11768_210.n10 a_11768_210.n9 27.2
R3005 a_11768_210.n3 a_11768_210.n2 23.284
R3006 a_11768_210.n11 a_11768_210.n10 22.4
R3007 a_11768_210.n7 a_11768_210.n4 19.017
R3008 a_11768_210.n6 a_11768_210.n5 13.494
R3009 a_11768_210.t1 a_11768_210.n1 7.04
R3010 a_11768_210.t1 a_11768_210.n3 5.727
R3011 a_11768_210.n8 a_11768_210.n7 1.435
R3012 a_7586_101.n12 a_7586_101.n11 26.811
R3013 a_7586_101.n6 a_7586_101.n5 24.977
R3014 a_7586_101.n2 a_7586_101.n1 24.877
R3015 a_7586_101.t0 a_7586_101.n2 12.677
R3016 a_7586_101.t0 a_7586_101.n3 11.595
R3017 a_7586_101.t1 a_7586_101.n8 8.137
R3018 a_7586_101.t0 a_7586_101.n4 7.273
R3019 a_7586_101.t0 a_7586_101.n0 6.109
R3020 a_7586_101.t1 a_7586_101.n7 4.864
R3021 a_7586_101.t0 a_7586_101.n12 2.074
R3022 a_7586_101.n7 a_7586_101.n6 1.13
R3023 a_7586_101.n12 a_7586_101.t1 0.937
R3024 a_7586_101.t1 a_7586_101.n10 0.804
R3025 a_7586_101.n10 a_7586_101.n9 0.136
R3026 a_757_103.n5 a_757_103.n4 19.724
R3027 a_757_103.t0 a_757_103.n3 11.595
R3028 a_757_103.t0 a_757_103.n5 9.207
R3029 a_757_103.n2 a_757_103.n1 2.455
R3030 a_757_103.n2 a_757_103.n0 1.32
R3031 a_757_103.t0 a_757_103.n2 0.246
R3032 a_5922_210.n9 a_5922_210.n7 82.852
R3033 a_5922_210.n3 a_5922_210.n1 44.628
R3034 a_5922_210.t0 a_5922_210.n9 32.417
R3035 a_5922_210.n7 a_5922_210.n6 27.2
R3036 a_5922_210.n5 a_5922_210.n4 23.498
R3037 a_5922_210.n3 a_5922_210.n2 23.284
R3038 a_5922_210.n7 a_5922_210.n5 22.4
R3039 a_5922_210.t0 a_5922_210.n11 20.241
R3040 a_5922_210.n11 a_5922_210.n10 13.494
R3041 a_5922_210.t0 a_5922_210.n0 8.137
R3042 a_5922_210.t0 a_5922_210.n3 5.727
R3043 a_5922_210.n9 a_5922_210.n8 1.435
R3044 a_16096_101.t0 a_16096_101.n1 34.62
R3045 a_16096_101.t0 a_16096_101.n0 8.137
R3046 a_16096_101.t0 a_16096_101.n2 4.69
R3047 a_4996_101.t0 a_4996_101.n1 34.62
R3048 a_4996_101.t0 a_4996_101.n0 8.137
R3049 a_4996_101.t0 a_4996_101.n2 4.69
R3050 a_112_101.t0 a_112_101.n1 34.62
R3051 a_112_101.t0 a_112_101.n0 8.137
R3052 a_112_101.t0 a_112_101.n2 4.69
R3053 a_8897_103.n1 a_8897_103.n0 25.576
R3054 a_8897_103.n3 a_8897_103.n2 9.111
R3055 a_8897_103.n7 a_8897_103.n5 7.859
R3056 a_8897_103.t0 a_8897_103.n7 3.034
R3057 a_8897_103.n5 a_8897_103.n3 1.964
R3058 a_8897_103.n5 a_8897_103.n4 1.964
R3059 a_8897_103.t0 a_8897_103.n1 1.871
R3060 a_8897_103.n7 a_8897_103.n6 0.443
R3061 a_9178_210.n8 a_9178_210.n6 96.467
R3062 a_9178_210.n3 a_9178_210.n1 44.628
R3063 a_9178_210.t0 a_9178_210.n8 32.417
R3064 a_9178_210.n3 a_9178_210.n2 23.284
R3065 a_9178_210.n6 a_9178_210.n5 22.349
R3066 a_9178_210.t0 a_9178_210.n10 20.241
R3067 a_9178_210.n10 a_9178_210.n9 13.494
R3068 a_9178_210.n6 a_9178_210.n4 8.443
R3069 a_9178_210.t0 a_9178_210.n0 8.137
R3070 a_9178_210.t0 a_9178_210.n3 5.727
R3071 a_9178_210.n8 a_9178_210.n7 1.435
R3072 a_3368_101.t0 a_3368_101.n1 34.62
R3073 a_3368_101.t0 a_3368_101.n0 8.137
R3074 a_3368_101.t0 a_3368_101.n2 4.69
R3075 a_9880_101.n12 a_9880_101.n11 26.811
R3076 a_9880_101.n6 a_9880_101.n5 24.977
R3077 a_9880_101.n2 a_9880_101.n1 24.877
R3078 a_9880_101.t0 a_9880_101.n2 12.677
R3079 a_9880_101.t0 a_9880_101.n3 11.595
R3080 a_9880_101.t1 a_9880_101.n8 8.137
R3081 a_9880_101.t0 a_9880_101.n4 7.273
R3082 a_9880_101.t0 a_9880_101.n0 6.109
R3083 a_9880_101.t1 a_9880_101.n7 4.864
R3084 a_9880_101.t0 a_9880_101.n12 2.074
R3085 a_9880_101.n7 a_9880_101.n6 1.13
R3086 a_9880_101.n12 a_9880_101.t1 0.937
R3087 a_9880_101.t1 a_9880_101.n10 0.804
R3088 a_9880_101.n10 a_9880_101.n9 0.136
R3089 a_1719_103.n1 a_1719_103.n0 25.576
R3090 a_1719_103.n3 a_1719_103.n2 9.111
R3091 a_1719_103.n7 a_1719_103.n6 2.455
R3092 a_1719_103.n5 a_1719_103.n3 1.964
R3093 a_1719_103.n5 a_1719_103.n4 1.964
R3094 a_1719_103.t0 a_1719_103.n1 1.871
R3095 a_1719_103.n7 a_1719_103.n5 0.636
R3096 a_1719_103.t0 a_1719_103.n7 0.246
R3097 a_13781_103.n5 a_13781_103.n4 19.724
R3098 a_13781_103.t0 a_13781_103.n3 11.595
R3099 a_13781_103.t0 a_13781_103.n5 9.207
R3100 a_13781_103.n2 a_13781_103.n1 2.455
R3101 a_13781_103.n2 a_13781_103.n0 1.32
R3102 a_13781_103.t0 a_13781_103.n2 0.246
R3103 a_2702_101.n12 a_2702_101.n11 26.811
R3104 a_2702_101.n6 a_2702_101.n5 24.977
R3105 a_2702_101.n2 a_2702_101.n1 24.877
R3106 a_2702_101.t0 a_2702_101.n2 12.677
R3107 a_2702_101.t0 a_2702_101.n3 11.595
R3108 a_2702_101.t1 a_2702_101.n8 8.137
R3109 a_2702_101.t0 a_2702_101.n4 7.273
R3110 a_2702_101.t0 a_2702_101.n0 6.109
R3111 a_2702_101.t1 a_2702_101.n7 4.864
R3112 a_2702_101.t0 a_2702_101.n12 2.074
R3113 a_2702_101.n7 a_2702_101.n6 1.13
R3114 a_2702_101.n12 a_2702_101.t1 0.937
R3115 a_2702_101.t1 a_2702_101.n10 0.804
R3116 a_2702_101.n10 a_2702_101.n9 0.136
R3117 a_8252_101.n12 a_8252_101.n11 26.811
R3118 a_8252_101.n6 a_8252_101.n5 24.977
R3119 a_8252_101.n2 a_8252_101.n1 24.877
R3120 a_8252_101.t0 a_8252_101.n2 12.677
R3121 a_8252_101.t0 a_8252_101.n3 11.595
R3122 a_8252_101.t1 a_8252_101.n8 8.137
R3123 a_8252_101.t0 a_8252_101.n4 7.273
R3124 a_8252_101.t0 a_8252_101.n0 6.109
R3125 a_8252_101.t1 a_8252_101.n7 4.864
R3126 a_8252_101.t0 a_8252_101.n12 2.074
R3127 a_8252_101.n7 a_8252_101.n6 1.13
R3128 a_8252_101.n12 a_8252_101.t1 0.937
R3129 a_8252_101.t1 a_8252_101.n10 0.804
R3130 a_8252_101.n10 a_8252_101.n9 0.136
R3131 a_5641_103.n5 a_5641_103.n4 19.724
R3132 a_5641_103.t0 a_5641_103.n3 11.595
R3133 a_5641_103.t0 a_5641_103.n5 9.207
R3134 a_5641_103.n2 a_5641_103.n1 2.455
R3135 a_5641_103.n2 a_5641_103.n0 1.32
R3136 a_5641_103.t0 a_5641_103.n2 0.246
R3137 a_14764_101.n1 a_14764_101.n0 32.249
R3138 a_14764_101.t0 a_14764_101.n5 7.911
R3139 a_14764_101.n4 a_14764_101.n2 4.032
R3140 a_14764_101.n4 a_14764_101.n3 3.644
R3141 a_14764_101.t0 a_14764_101.n1 2.534
R3142 a_14764_101.t0 a_14764_101.n4 1.099
C7 SN GND 8.21fF
C8 VDD GND 60.49fF
C9 a_14764_101.n0 GND 0.11fF
C10 a_14764_101.n1 GND 0.09fF
C11 a_14764_101.n2 GND 0.08fF
C12 a_14764_101.n3 GND 0.02fF
C13 a_14764_101.n4 GND 0.01fF
C14 a_14764_101.n5 GND 0.06fF
C15 a_5641_103.n0 GND 0.10fF
C16 a_5641_103.n1 GND 0.04fF
C17 a_5641_103.n2 GND 0.03fF
C18 a_5641_103.n3 GND 0.07fF
C19 a_5641_103.n4 GND 0.08fF
C20 a_5641_103.n5 GND 0.06fF
C21 a_8252_101.n0 GND 0.02fF
C22 a_8252_101.n1 GND 0.10fF
C23 a_8252_101.n2 GND 0.06fF
C24 a_8252_101.n3 GND 0.06fF
C25 a_8252_101.n4 GND 0.00fF
C26 a_8252_101.n5 GND 0.04fF
C27 a_8252_101.n6 GND 0.05fF
C28 a_8252_101.n7 GND 0.02fF
C29 a_8252_101.n8 GND 0.05fF
C30 a_8252_101.n9 GND 0.08fF
C31 a_8252_101.n10 GND 0.17fF
C32 a_8252_101.t1 GND 0.23fF
C33 a_8252_101.n11 GND 0.09fF
C34 a_8252_101.n12 GND 0.00fF
C35 a_2702_101.n0 GND 0.02fF
C36 a_2702_101.n1 GND 0.10fF
C37 a_2702_101.n2 GND 0.06fF
C38 a_2702_101.n3 GND 0.06fF
C39 a_2702_101.n4 GND 0.00fF
C40 a_2702_101.n5 GND 0.04fF
C41 a_2702_101.n6 GND 0.05fF
C42 a_2702_101.n7 GND 0.02fF
C43 a_2702_101.n8 GND 0.05fF
C44 a_2702_101.n9 GND 0.08fF
C45 a_2702_101.n10 GND 0.17fF
C46 a_2702_101.t1 GND 0.23fF
C47 a_2702_101.n11 GND 0.09fF
C48 a_2702_101.n12 GND 0.00fF
C49 a_13781_103.n0 GND 0.10fF
C50 a_13781_103.n1 GND 0.04fF
C51 a_13781_103.n2 GND 0.03fF
C52 a_13781_103.n3 GND 0.07fF
C53 a_13781_103.n4 GND 0.08fF
C54 a_13781_103.n5 GND 0.06fF
C55 a_1719_103.n0 GND 0.09fF
C56 a_1719_103.n1 GND 0.10fF
C57 a_1719_103.n2 GND 0.05fF
C58 a_1719_103.n3 GND 0.03fF
C59 a_1719_103.n4 GND 0.04fF
C60 a_1719_103.n5 GND 0.03fF
C61 a_1719_103.n6 GND 0.04fF
C62 a_9880_101.n0 GND 0.02fF
C63 a_9880_101.n1 GND 0.10fF
C64 a_9880_101.n2 GND 0.06fF
C65 a_9880_101.n3 GND 0.06fF
C66 a_9880_101.n4 GND 0.00fF
C67 a_9880_101.n5 GND 0.04fF
C68 a_9880_101.n6 GND 0.05fF
C69 a_9880_101.n7 GND 0.02fF
C70 a_9880_101.n8 GND 0.05fF
C71 a_9880_101.n9 GND 0.08fF
C72 a_9880_101.n10 GND 0.17fF
C73 a_9880_101.t1 GND 0.23fF
C74 a_9880_101.n11 GND 0.09fF
C75 a_9880_101.n12 GND 0.00fF
C76 a_3368_101.n0 GND 0.05fF
C77 a_3368_101.n1 GND 0.12fF
C78 a_3368_101.n2 GND 0.04fF
C79 a_9178_210.n0 GND 0.07fF
C80 a_9178_210.n1 GND 0.09fF
C81 a_9178_210.n2 GND 0.13fF
C82 a_9178_210.n3 GND 0.11fF
C83 a_9178_210.n4 GND 0.02fF
C84 a_9178_210.n5 GND 0.03fF
C85 a_9178_210.n6 GND 0.06fF
C86 a_9178_210.n7 GND 0.03fF
C87 a_9178_210.n8 GND 0.12fF
C88 a_9178_210.n9 GND 0.06fF
C89 a_9178_210.n10 GND 0.01fF
C90 a_9178_210.t0 GND 0.33fF
C91 a_8897_103.n0 GND 0.09fF
C92 a_8897_103.n1 GND 0.10fF
C93 a_8897_103.n2 GND 0.05fF
C94 a_8897_103.n3 GND 0.03fF
C95 a_8897_103.n4 GND 0.04fF
C96 a_8897_103.n5 GND 0.11fF
C97 a_8897_103.n6 GND 0.04fF
C98 a_112_101.n0 GND 0.05fF
C99 a_112_101.n1 GND 0.12fF
C100 a_112_101.n2 GND 0.04fF
C101 a_4996_101.n0 GND 0.05fF
C102 a_4996_101.n1 GND 0.12fF
C103 a_4996_101.n2 GND 0.04fF
C104 a_16096_101.n0 GND 0.06fF
C105 a_16096_101.n1 GND 0.13fF
C106 a_16096_101.n2 GND 0.04fF
C107 a_5922_210.n0 GND 0.07fF
C108 a_5922_210.n1 GND 0.09fF
C109 a_5922_210.n2 GND 0.13fF
C110 a_5922_210.n3 GND 0.11fF
C111 a_5922_210.n4 GND 0.02fF
C112 a_5922_210.n5 GND 0.03fF
C113 a_5922_210.n6 GND 0.02fF
C114 a_5922_210.n7 GND 0.05fF
C115 a_5922_210.n8 GND 0.03fF
C116 a_5922_210.n9 GND 0.11fF
C117 a_5922_210.n10 GND 0.06fF
C118 a_5922_210.n11 GND 0.01fF
C119 a_5922_210.t0 GND 0.33fF
C120 a_757_103.n0 GND 0.10fF
C121 a_757_103.n1 GND 0.04fF
C122 a_757_103.n2 GND 0.03fF
C123 a_757_103.n3 GND 0.07fF
C124 a_757_103.n4 GND 0.08fF
C125 a_757_103.n5 GND 0.06fF
C126 a_7586_101.n0 GND 0.02fF
C127 a_7586_101.n1 GND 0.10fF
C128 a_7586_101.n2 GND 0.06fF
C129 a_7586_101.n3 GND 0.06fF
C130 a_7586_101.n4 GND 0.00fF
C131 a_7586_101.n5 GND 0.04fF
C132 a_7586_101.n6 GND 0.05fF
C133 a_7586_101.n7 GND 0.02fF
C134 a_7586_101.n8 GND 0.05fF
C135 a_7586_101.n9 GND 0.08fF
C136 a_7586_101.n10 GND 0.17fF
C137 a_7586_101.t1 GND 0.23fF
C138 a_7586_101.n11 GND 0.09fF
C139 a_7586_101.n12 GND 0.00fF
C140 a_11768_210.n0 GND 0.02fF
C141 a_11768_210.n1 GND 0.09fF
C142 a_11768_210.n2 GND 0.13fF
C143 a_11768_210.n3 GND 0.11fF
C144 a_11768_210.t1 GND 0.30fF
C145 a_11768_210.n4 GND 0.09fF
C146 a_11768_210.n5 GND 0.06fF
C147 a_11768_210.n6 GND 0.01fF
C148 a_11768_210.n7 GND 0.03fF
C149 a_11768_210.n8 GND 0.11fF
C150 a_11768_210.n9 GND 0.02fF
C151 a_11768_210.n10 GND 0.05fF
C152 a_11768_210.n11 GND 0.02fF
C153 a_14062_210.n0 GND 0.02fF
C154 a_14062_210.n1 GND 0.09fF
C155 a_14062_210.n2 GND 0.13fF
C156 a_14062_210.n3 GND 0.11fF
C157 a_14062_210.t1 GND 0.30fF
C158 a_14062_210.n4 GND 0.09fF
C159 a_14062_210.n5 GND 0.06fF
C160 a_14062_210.n6 GND 0.01fF
C161 a_14062_210.n7 GND 0.03fF
C162 a_14062_210.n8 GND 0.11fF
C163 a_14062_210.n9 GND 0.02fF
C164 a_14062_210.n10 GND 0.05fF
C165 a_14062_210.n11 GND 0.03fF
C166 a_1038_210.n0 GND 0.02fF
C167 a_1038_210.n1 GND 0.09fF
C168 a_1038_210.n2 GND 0.13fF
C169 a_1038_210.n3 GND 0.11fF
C170 a_1038_210.t1 GND 0.30fF
C171 a_1038_210.n4 GND 0.09fF
C172 a_1038_210.n5 GND 0.06fF
C173 a_1038_210.n6 GND 0.01fF
C174 a_1038_210.n7 GND 0.03fF
C175 a_1038_210.n8 GND 0.11fF
C176 a_1038_210.n9 GND 0.02fF
C177 a_1038_210.n10 GND 0.05fF
C178 a_1038_210.n11 GND 0.03fF
C179 a_6789_1050.n0 GND 0.45fF
C180 a_6789_1050.n1 GND 0.58fF
C181 a_6789_1050.n2 GND 0.35fF
C182 a_6789_1050.n3 GND 0.68fF
C183 a_6789_1050.n4 GND 0.55fF
C184 a_6789_1050.n5 GND 0.65fF
C185 a_6789_1050.n6 GND 0.21fF
C186 a_6789_1050.n7 GND 0.38fF
C187 a_6789_1050.n8 GND 0.55fF
C188 a_10111_411.n0 GND 0.86fF
C189 a_10111_411.n1 GND 0.86fF
C190 a_10111_411.n2 GND 0.50fF
C191 a_10111_411.n3 GND 0.76fF
C192 a_10111_411.n4 GND 0.44fF
C193 a_10111_411.t10 GND 0.94fF
C194 a_10111_411.n5 GND 0.65fF
C195 a_10111_411.n6 GND 4.01fF
C196 a_10111_411.n7 GND 0.07fF
C197 a_10111_411.n8 GND 0.09fF
C198 a_10111_411.n9 GND 0.60fF
C199 a_10111_411.n10 GND 0.76fF
C200 a_10111_411.n11 GND 0.39fF
C201 a_10111_411.n12 GND 0.32fF
C202 a_10111_411.n13 GND 1.01fF
C203 a_15430_101.n0 GND 0.13fF
C204 a_15430_101.n1 GND 0.13fF
C205 a_217_1050.n0 GND 0.35fF
C206 a_217_1050.n1 GND 0.42fF
C207 a_217_1050.n2 GND 0.35fF
C208 a_217_1050.n3 GND 0.41fF
C209 a_217_1050.n4 GND 0.99fF
C210 a_217_1050.n5 GND 0.04fF
C211 a_217_1050.n6 GND 0.05fF
C212 a_217_1050.n7 GND 0.03fF
C213 a_217_1050.n8 GND 0.21fF
C214 a_217_1050.n9 GND 0.38fF
C215 a_217_1050.n10 GND 0.55fF
C216 a_217_1050.n11 GND 0.32fF
C217 a_217_1050.n12 GND 0.46fF
C218 a_12470_101.n0 GND 0.02fF
C219 a_12470_101.n1 GND 0.10fF
C220 a_12470_101.n2 GND 0.06fF
C221 a_12470_101.n3 GND 0.06fF
C222 a_12470_101.n4 GND 0.00fF
C223 a_12470_101.n5 GND 0.04fF
C224 a_12470_101.n6 GND 0.05fF
C225 a_12470_101.n7 GND 0.02fF
C226 a_12470_101.n8 GND 0.05fF
C227 a_12470_101.n9 GND 0.08fF
C228 a_12470_101.n10 GND 0.17fF
C229 a_12470_101.t1 GND 0.23fF
C230 a_12470_101.n11 GND 0.09fF
C231 a_12470_101.n12 GND 0.00fF
C232 a_10806_210.n0 GND 0.02fF
C233 a_10806_210.n1 GND 0.07fF
C234 a_10806_210.n2 GND 0.13fF
C235 a_10806_210.n3 GND 0.09fF
C236 a_10806_210.t1 GND 0.25fF
C237 a_10806_210.n4 GND 0.05fF
C238 a_10806_210.n5 GND 0.06fF
C239 a_10806_210.n6 GND 0.07fF
C240 a_10806_210.n7 GND 0.07fF
C241 a_10806_210.n8 GND 0.03fF
C242 a_10806_210.n9 GND 0.01fF
C243 a_10806_210.n10 GND 0.11fF
C244 a_10806_210.n11 GND 0.02fF
C245 a_10806_210.n12 GND 0.05fF
C246 a_10806_210.n13 GND 0.02fF
C247 a_10525_103.n0 GND 0.20fF
C248 a_10525_103.n1 GND 0.04fF
C249 a_10525_103.n2 GND 0.01fF
C250 a_10525_103.n3 GND 0.08fF
C251 a_10525_103.n4 GND 0.06fF
C252 a_10525_103.n5 GND 0.07fF
C253 a_2000_210.n0 GND 0.02fF
C254 a_2000_210.n1 GND 0.09fF
C255 a_2000_210.n2 GND 0.13fF
C256 a_2000_210.n3 GND 0.11fF
C257 a_2000_210.t1 GND 0.30fF
C258 a_2000_210.n4 GND 0.09fF
C259 a_2000_210.n5 GND 0.06fF
C260 a_2000_210.n6 GND 0.01fF
C261 a_2000_210.n7 GND 0.03fF
C262 a_2000_210.n8 GND 0.11fF
C263 a_2000_210.n9 GND 0.02fF
C264 a_2000_210.n10 GND 0.05fF
C265 a_2000_210.n11 GND 0.03fF
C266 a_15533_1051.n0 GND 0.35fF
C267 a_15533_1051.n1 GND 0.29fF
C268 a_15533_1051.n2 GND 0.20fF
C269 a_15533_1051.n3 GND 0.56fF
C270 a_15533_1051.n4 GND 0.25fF
C271 a_15533_1051.n5 GND 0.28fF
C272 QN.n0 GND 0.42fF
C273 QN.n1 GND 0.51fF
C274 QN.n2 GND 0.25fF
C275 QN.n3 GND 0.04fF
C276 QN.n4 GND 0.05fF
C277 QN.n5 GND 0.03fF
C278 QN.n6 GND 0.09fF
C279 QN.n7 GND 0.04fF
C280 QN.n8 GND 0.05fF
C281 QN.n9 GND 0.03fF
C282 QN.n10 GND 0.10fF
C283 QN.n11 GND 1.06fF
C284 QN.n12 GND 0.06fF
C285 QN.n13 GND 0.03fF
C286 QN.n14 GND 0.08fF
C287 QN.n15 GND 0.28fF
C288 QN.n16 GND 0.37fF
C289 QN.n17 GND 0.01fF
C290 a_11673_1050.n0 GND 0.55fF
C291 a_11673_1050.n1 GND 0.45fF
C292 a_11673_1050.n2 GND 0.57fF
C293 a_11673_1050.n3 GND 0.04fF
C294 a_11673_1050.n4 GND 0.06fF
C295 a_11673_1050.n5 GND 0.04fF
C296 a_11673_1050.n6 GND 0.24fF
C297 a_11673_1050.n7 GND 0.65fF
C298 a_11673_1050.n8 GND 0.38fF
C299 a_11673_1050.n9 GND 0.65fF
C300 a_11673_1050.n10 GND 0.20fF
C301 a_11673_1050.n11 GND 0.55fF
C302 a_1905_1050.n0 GND 0.50fF
C303 a_1905_1050.n1 GND 0.41fF
C304 a_1905_1050.n2 GND 0.53fF
C305 a_1905_1050.n3 GND 0.04fF
C306 a_1905_1050.n4 GND 0.05fF
C307 a_1905_1050.n5 GND 0.03fF
C308 a_1905_1050.n6 GND 0.22fF
C309 a_1905_1050.n7 GND 0.59fF
C310 a_1905_1050.n8 GND 0.35fF
C311 a_1905_1050.n9 GND 0.59fF
C312 a_1905_1050.n10 GND 0.19fF
C313 a_1905_1050.n11 GND 0.50fF
C314 a_5227_411.n0 GND 0.48fF
C315 a_5227_411.n1 GND 0.74fF
C316 a_5227_411.n2 GND 0.43fF
C317 a_5227_411.t7 GND 0.91fF
C318 a_5227_411.n3 GND 0.63fF
C319 a_5227_411.n4 GND 3.88fF
C320 a_5227_411.n5 GND 0.06fF
C321 a_5227_411.n6 GND 0.08fF
C322 a_5227_411.n7 GND 0.05fF
C323 a_5227_411.n8 GND 0.56fF
C324 a_5227_411.n9 GND 0.70fF
C325 a_5227_411.n10 GND 0.83fF
C326 a_5227_411.n11 GND 0.98fF
C327 a_5227_411.n12 GND 0.31fF
C328 a_5227_411.n13 GND 0.38fF
C329 a_5227_411.n14 GND 0.83fF
C330 a_5101_1050.n0 GND 0.71fF
C331 a_5101_1050.n1 GND 0.84fF
C332 a_5101_1050.n2 GND 0.49fF
C333 a_5101_1050.n3 GND 0.54fF
C334 a_5101_1050.n4 GND 0.65fF
C335 a_5101_1050.n5 GND 0.54fF
C336 a_5101_1050.n6 GND 0.63fF
C337 a_5101_1050.n7 GND 1.52fF
C338 a_5101_1050.n8 GND 0.59fF
C339 a_5101_1050.n9 GND 0.11fF
C340 a_5101_1050.n10 GND 0.30fF
C341 a_5101_1050.n11 GND 0.06fF
C342 a_11033_989.n0 GND 0.59fF
C343 a_11033_989.t6 GND 0.97fF
C344 a_11033_989.n1 GND 0.71fF
C345 a_11033_989.n2 GND 0.59fF
C346 a_11033_989.t12 GND 0.96fF
C347 a_11033_989.n3 GND 0.64fF
C348 a_11033_989.n4 GND 0.59fF
C349 a_11033_989.t10 GND 0.97fF
C350 a_11033_989.n5 GND 0.67fF
C351 a_11033_989.n6 GND 1.96fF
C352 a_11033_989.n7 GND 2.64fF
C353 a_11033_989.n8 GND 0.07fF
C354 a_11033_989.n9 GND 0.09fF
C355 a_11033_989.n10 GND 0.06fF
C356 a_11033_989.n11 GND 0.57fF
C357 a_11033_989.n12 GND 0.73fF
C358 a_11033_989.n13 GND 1.08fF
C359 a_11033_989.n14 GND 0.47fF
C360 a_11033_989.n15 GND 0.91fF
C361 a_343_411.n0 GND 0.72fF
C362 a_343_411.n1 GND 0.42fF
C363 a_343_411.n2 GND 0.64fF
C364 a_343_411.n3 GND 0.37fF
C365 a_343_411.t11 GND 0.79fF
C366 a_343_411.n4 GND 0.55fF
C367 a_343_411.n5 GND 3.36fF
C368 a_343_411.n6 GND 0.05fF
C369 a_343_411.n7 GND 0.07fF
C370 a_343_411.n8 GND 0.05fF
C371 a_343_411.n9 GND 0.49fF
C372 a_343_411.n10 GND 0.61fF
C373 a_343_411.n11 GND 0.33fF
C374 a_343_411.n12 GND 0.85fF
C375 a_343_411.n13 GND 0.27fF
C376 a_343_411.n14 GND 0.72fF
C377 a_1265_989.n0 GND 0.45fF
C378 a_1265_989.t13 GND 0.73fF
C379 a_1265_989.n1 GND 0.54fF
C380 a_1265_989.n2 GND 0.45fF
C381 a_1265_989.t6 GND 0.73fF
C382 a_1265_989.n3 GND 0.48fF
C383 a_1265_989.n4 GND 0.45fF
C384 a_1265_989.t8 GND 0.73fF
C385 a_1265_989.n5 GND 0.51fF
C386 a_1265_989.n6 GND 1.49fF
C387 a_1265_989.n7 GND 2.01fF
C388 a_1265_989.n8 GND 0.05fF
C389 a_1265_989.n9 GND 0.07fF
C390 a_1265_989.n10 GND 0.04fF
C391 a_1265_989.n11 GND 0.43fF
C392 a_1265_989.n12 GND 0.55fF
C393 a_1265_989.n13 GND 0.82fF
C394 a_1265_989.n14 GND 0.36fF
C395 a_1265_989.n15 GND 0.69fF
C396 a_11487_103.n0 GND 0.03fF
C397 a_11487_103.n1 GND 0.10fF
C398 a_11487_103.n2 GND 0.10fF
C399 a_11487_103.n3 GND 0.05fF
C400 a_11487_103.n4 GND 0.03fF
C401 a_11487_103.n5 GND 0.04fF
C402 a_11487_103.n6 GND 0.11fF
C403 a_11487_103.n7 GND 0.04fF
C404 a_9985_1050.n0 GND 0.71fF
C405 a_9985_1050.n1 GND 0.83fF
C406 a_9985_1050.n2 GND 0.49fF
C407 a_9985_1050.n3 GND 0.53fF
C408 a_9985_1050.n4 GND 0.65fF
C409 a_9985_1050.n5 GND 0.53fF
C410 a_9985_1050.n6 GND 0.62fF
C411 a_9985_1050.n7 GND 1.51fF
C412 a_9985_1050.n8 GND 0.58fF
C413 a_9985_1050.n9 GND 0.11fF
C414 a_9985_1050.n10 GND 0.30fF
C415 a_9985_1050.n11 GND 0.06fF
C416 a_4294_210.n0 GND 0.02fF
C417 a_4294_210.n1 GND 0.09fF
C418 a_4294_210.n2 GND 0.13fF
C419 a_4294_210.n3 GND 0.11fF
C420 a_4294_210.t1 GND 0.30fF
C421 a_4294_210.n4 GND 0.09fF
C422 a_4294_210.n5 GND 0.06fF
C423 a_4294_210.n6 GND 0.01fF
C424 a_4294_210.n7 GND 0.03fF
C425 a_4294_210.n8 GND 0.11fF
C426 a_4294_210.n9 GND 0.02fF
C427 a_4294_210.n10 GND 0.05fF
C428 a_4294_210.n11 GND 0.02fF
C429 a_4013_103.n0 GND 0.20fF
C430 a_4013_103.n1 GND 0.04fF
C431 a_4013_103.n2 GND 0.01fF
C432 a_4013_103.n3 GND 0.03fF
C433 a_4013_103.n4 GND 0.05fF
C434 a_4013_103.n5 GND 0.09fF
C435 a_4013_103.n6 GND 0.07fF
C436 a_13241_1050.n0 GND 0.24fF
C437 a_13241_1050.n1 GND 0.70fF
C438 a_13241_1050.n2 GND 0.48fF
C439 a_13241_1050.n3 GND 0.59fF
C440 a_13241_1050.n4 GND 0.62fF
C441 a_13241_1050.n5 GND 0.21fF
C442 a_13241_1050.n6 GND 0.52fF
C443 a_13136_101.n0 GND 0.05fF
C444 a_13136_101.n1 GND 0.02fF
C445 a_13136_101.n2 GND 0.12fF
C446 a_13136_101.n3 GND 0.04fF
C447 a_13136_101.n4 GND 0.17fF
C448 a_13367_411.n0 GND 0.58fF
C449 a_13367_411.n1 GND 0.33fF
C450 a_13367_411.n2 GND 0.47fF
C451 a_13367_411.n3 GND 0.30fF
C452 a_13367_411.n4 GND 0.41fF
C453 a_13367_411.n5 GND 1.40fF
C454 a_13367_411.n6 GND 0.30fF
C455 a_13367_411.t7 GND 0.63fF
C456 a_13367_411.n7 GND 0.44fF
C457 a_13367_411.n8 GND 1.22fF
C458 a_13367_411.n9 GND 0.05fF
C459 a_13367_411.n10 GND 0.06fF
C460 a_13367_411.n11 GND 0.40fF
C461 a_13367_411.n12 GND 0.51fF
C462 a_13367_411.n13 GND 0.26fF
C463 a_13367_411.n14 GND 0.68fF
C464 a_13367_411.n15 GND 0.21fF
C465 a_13367_411.n16 GND 0.58fF
C466 a_14869_1051.n0 GND 0.37fF
C467 a_14869_1051.n1 GND 0.33fF
C468 a_14869_1051.n2 GND 0.23fF
C469 a_14869_1051.n3 GND 0.63fF
C470 a_14869_1051.n4 GND 0.28fF
C471 a_14869_1051.n5 GND 0.41fF
C472 a_6149_989.n0 GND 0.53fF
C473 a_6149_989.t12 GND 0.86fF
C474 a_6149_989.n1 GND 0.63fF
C475 a_6149_989.n2 GND 0.53fF
C476 a_6149_989.t7 GND 0.85fF
C477 a_6149_989.n3 GND 0.56fF
C478 a_6149_989.n4 GND 0.53fF
C479 a_6149_989.t6 GND 0.86fF
C480 a_6149_989.n5 GND 0.59fF
C481 a_6149_989.n6 GND 1.74fF
C482 a_6149_989.n7 GND 2.34fF
C483 a_6149_989.n8 GND 0.06fF
C484 a_6149_989.n9 GND 0.08fF
C485 a_6149_989.n10 GND 0.05fF
C486 a_6149_989.n11 GND 0.50fF
C487 a_6149_989.n12 GND 0.65fF
C488 a_6149_989.n13 GND 0.96fF
C489 a_6149_989.n14 GND 0.42fF
C490 a_6149_989.n15 GND 0.81fF
C491 a_3599_411.n0 GND 1.04fF
C492 a_3599_411.n1 GND 1.04fF
C493 a_3599_411.n2 GND 0.73fF
C494 a_3599_411.n3 GND 0.91fF
C495 a_3599_411.n4 GND 1.13fF
C496 a_3599_411.n5 GND 0.70fF
C497 a_3599_411.n6 GND 3.68fF
C498 a_3599_411.n7 GND 0.71fF
C499 a_3599_411.t12 GND 0.98fF
C500 a_3599_411.n8 GND 0.78fF
C501 a_3599_411.n9 GND 16.28fF
C502 a_3599_411.n10 GND 0.08fF
C503 a_3599_411.n11 GND 0.10fF
C504 a_3599_411.n12 GND 0.07fF
C505 a_3599_411.n13 GND 0.52fF
C506 a_3599_411.n14 GND 0.87fF
C507 a_3599_411.n15 GND 0.65fF
C508 a_3599_411.n16 GND 0.38fF
C509 a_3599_411.n17 GND 1.22fF
C510 a_3473_1050.n0 GND 0.57fF
C511 a_3473_1050.n1 GND 0.67fF
C512 a_3473_1050.n2 GND 0.26fF
C513 a_3473_1050.n3 GND 0.29fF
C514 a_3473_1050.n4 GND 0.71fF
C515 a_3473_1050.n5 GND 0.65fF
C516 a_3473_1050.n6 GND 0.09fF
C517 a_3473_1050.n7 GND 0.38fF
C518 a_3473_1050.n8 GND 0.05fF
C519 a_6884_210.n0 GND 0.02fF
C520 a_6884_210.n1 GND 0.09fF
C521 a_6884_210.n2 GND 0.13fF
C522 a_6884_210.n3 GND 0.11fF
C523 a_6884_210.t1 GND 0.30fF
C524 a_6884_210.n4 GND 0.09fF
C525 a_6884_210.n5 GND 0.06fF
C526 a_6884_210.n6 GND 0.01fF
C527 a_6884_210.n7 GND 0.03fF
C528 a_6884_210.n8 GND 0.11fF
C529 a_6884_210.n9 GND 0.02fF
C530 a_6884_210.n10 GND 0.05fF
C531 a_6884_210.n11 GND 0.02fF
C532 a_6603_103.n0 GND 0.03fF
C533 a_6603_103.n1 GND 0.10fF
C534 a_6603_103.n2 GND 0.10fF
C535 a_6603_103.n3 GND 0.05fF
C536 a_6603_103.n4 GND 0.03fF
C537 a_6603_103.n5 GND 0.04fF
C538 a_6603_103.n6 GND 0.11fF
C539 a_6603_103.n7 GND 0.04fF
C540 SN.n0 GND 0.87fF
C541 SN.t10 GND 0.80fF
C542 SN.n1 GND 0.83fF
C543 SN.n2 GND 0.87fF
C544 SN.t5 GND 0.80fF
C545 SN.n3 GND 0.65fF
C546 SN.n4 GND 5.21fF
C547 SN.n5 GND 0.87fF
C548 SN.t6 GND 0.80fF
C549 SN.n6 GND 0.65fF
C550 SN.n7 GND 3.64fF
C551 SN.n8 GND 0.87fF
C552 SN.t0 GND 0.80fF
C553 SN.n9 GND 0.65fF
C554 SN.n10 GND 3.64fF
C555 SN.n11 GND 0.87fF
C556 SN.t1 GND 0.80fF
C557 SN.n12 GND 0.65fF
C558 SN.n13 GND 3.64fF
C559 SN.n14 GND 0.87fF
C560 SN.t11 GND 0.80fF
C561 SN.n15 GND 0.65fF
C562 SN.n16 GND 1.73fF
C563 a_8357_1050.n0 GND 0.31fF
C564 a_8357_1050.n1 GND 0.74fF
C565 a_8357_1050.n2 GND 0.05fF
C566 a_8357_1050.n3 GND 0.06fF
C567 a_8357_1050.n4 GND 0.04fF
C568 a_8357_1050.n5 GND 0.40fF
C569 a_8357_1050.n6 GND 0.67fF
C570 a_8357_1050.n7 GND 0.70fF
C571 a_8357_1050.n8 GND 0.27fF
C572 a_8357_1050.n9 GND 0.59fF
C573 VDD.n0 GND 0.15fF
C574 VDD.n1 GND 0.03fF
C575 VDD.n2 GND 0.02fF
C576 VDD.n3 GND 0.05fF
C577 VDD.n4 GND 0.01fF
C578 VDD.n5 GND 0.02fF
C579 VDD.n6 GND 0.02fF
C580 VDD.n9 GND 0.02fF
C581 VDD.n10 GND 0.02fF
C582 VDD.n12 GND 0.02fF
C583 VDD.n14 GND 0.46fF
C584 VDD.n16 GND 0.03fF
C585 VDD.n17 GND 0.02fF
C586 VDD.n18 GND 0.02fF
C587 VDD.n19 GND 0.02fF
C588 VDD.n20 GND 0.04fF
C589 VDD.n21 GND 0.28fF
C590 VDD.n22 GND 0.02fF
C591 VDD.n23 GND 0.03fF
C592 VDD.n24 GND 0.28fF
C593 VDD.n25 GND 0.01fF
C594 VDD.n26 GND 0.31fF
C595 VDD.n27 GND 0.01fF
C596 VDD.n28 GND 0.03fF
C597 VDD.n29 GND 0.02fF
C598 VDD.n30 GND 0.28fF
C599 VDD.n31 GND 0.01fF
C600 VDD.n32 GND 0.02fF
C601 VDD.n33 GND 0.00fF
C602 VDD.n34 GND 0.09fF
C603 VDD.n35 GND 0.03fF
C604 VDD.n36 GND 0.31fF
C605 VDD.n37 GND 0.01fF
C606 VDD.n38 GND 0.03fF
C607 VDD.n39 GND 0.03fF
C608 VDD.n40 GND 0.28fF
C609 VDD.n41 GND 0.01fF
C610 VDD.n42 GND 0.02fF
C611 VDD.n43 GND 0.02fF
C612 VDD.n44 GND 0.28fF
C613 VDD.n45 GND 0.01fF
C614 VDD.n46 GND 0.02fF
C615 VDD.n47 GND 0.02fF
C616 VDD.n48 GND 0.28fF
C617 VDD.n49 GND 0.01fF
C618 VDD.n50 GND 0.02fF
C619 VDD.n51 GND 0.03fF
C620 VDD.n52 GND 0.02fF
C621 VDD.n53 GND 0.02fF
C622 VDD.n54 GND 0.02fF
C623 VDD.n55 GND 0.22fF
C624 VDD.n56 GND 0.04fF
C625 VDD.n57 GND 0.04fF
C626 VDD.n58 GND 0.02fF
C627 VDD.n60 GND 0.02fF
C628 VDD.n61 GND 0.02fF
C629 VDD.n62 GND 0.02fF
C630 VDD.n63 GND 0.02fF
C631 VDD.n65 GND 0.02fF
C632 VDD.n66 GND 0.02fF
C633 VDD.n67 GND 0.02fF
C634 VDD.n69 GND 0.28fF
C635 VDD.n71 GND 0.02fF
C636 VDD.n72 GND 0.02fF
C637 VDD.n73 GND 0.03fF
C638 VDD.n74 GND 0.02fF
C639 VDD.n75 GND 0.28fF
C640 VDD.n76 GND 0.01fF
C641 VDD.n77 GND 0.02fF
C642 VDD.n78 GND 0.03fF
C643 VDD.n79 GND 0.28fF
C644 VDD.n80 GND 0.01fF
C645 VDD.n81 GND 0.02fF
C646 VDD.n82 GND 0.02fF
C647 VDD.n83 GND 0.28fF
C648 VDD.n84 GND 0.01fF
C649 VDD.n85 GND 0.02fF
C650 VDD.n86 GND 0.02fF
C651 VDD.n87 GND 0.31fF
C652 VDD.n88 GND 0.01fF
C653 VDD.n89 GND 0.03fF
C654 VDD.n90 GND 0.03fF
C655 VDD.n91 GND 0.31fF
C656 VDD.n92 GND 0.01fF
C657 VDD.n93 GND 0.03fF
C658 VDD.n94 GND 0.03fF
C659 VDD.n95 GND 0.28fF
C660 VDD.n96 GND 0.01fF
C661 VDD.n97 GND 0.02fF
C662 VDD.n98 GND 0.02fF
C663 VDD.n99 GND 0.28fF
C664 VDD.n100 GND 0.01fF
C665 VDD.n101 GND 0.02fF
C666 VDD.n102 GND 0.02fF
C667 VDD.n103 GND 0.28fF
C668 VDD.n104 GND 0.01fF
C669 VDD.n105 GND 0.02fF
C670 VDD.n106 GND 0.03fF
C671 VDD.n107 GND 0.02fF
C672 VDD.n108 GND 0.02fF
C673 VDD.n109 GND 0.02fF
C674 VDD.n110 GND 0.22fF
C675 VDD.n111 GND 0.04fF
C676 VDD.n112 GND 0.03fF
C677 VDD.n113 GND 0.02fF
C678 VDD.n114 GND 0.02fF
C679 VDD.n115 GND 0.02fF
C680 VDD.n116 GND 0.03fF
C681 VDD.n117 GND 0.02fF
C682 VDD.n119 GND 0.02fF
C683 VDD.n120 GND 0.02fF
C684 VDD.n121 GND 0.02fF
C685 VDD.n123 GND 0.28fF
C686 VDD.n125 GND 0.02fF
C687 VDD.n126 GND 0.02fF
C688 VDD.n127 GND 0.03fF
C689 VDD.n128 GND 0.02fF
C690 VDD.n129 GND 0.28fF
C691 VDD.n130 GND 0.01fF
C692 VDD.n131 GND 0.02fF
C693 VDD.n132 GND 0.03fF
C694 VDD.n133 GND 0.06fF
C695 VDD.n134 GND 0.24fF
C696 VDD.n135 GND 0.01fF
C697 VDD.n136 GND 0.01fF
C698 VDD.n137 GND 0.02fF
C699 VDD.n138 GND 0.14fF
C700 VDD.n139 GND 0.17fF
C701 VDD.n140 GND 0.01fF
C702 VDD.n141 GND 0.02fF
C703 VDD.n142 GND 0.02fF
C704 VDD.n143 GND 0.11fF
C705 VDD.n144 GND 0.03fF
C706 VDD.n145 GND 0.31fF
C707 VDD.n146 GND 0.01fF
C708 VDD.n147 GND 0.02fF
C709 VDD.n148 GND 0.03fF
C710 VDD.n149 GND 0.17fF
C711 VDD.n150 GND 0.14fF
C712 VDD.n151 GND 0.01fF
C713 VDD.n152 GND 0.02fF
C714 VDD.n153 GND 0.03fF
C715 VDD.n154 GND 0.14fF
C716 VDD.n155 GND 0.16fF
C717 VDD.n156 GND 0.01fF
C718 VDD.n157 GND 0.02fF
C719 VDD.n158 GND 0.02fF
C720 VDD.n159 GND 0.06fF
C721 VDD.n160 GND 0.25fF
C722 VDD.n161 GND 0.01fF
C723 VDD.n162 GND 0.01fF
C724 VDD.n163 GND 0.02fF
C725 VDD.n164 GND 0.28fF
C726 VDD.n165 GND 0.01fF
C727 VDD.n166 GND 0.02fF
C728 VDD.n167 GND 0.03fF
C729 VDD.n168 GND 0.02fF
C730 VDD.n169 GND 0.02fF
C731 VDD.n170 GND 0.02fF
C732 VDD.n171 GND 0.26fF
C733 VDD.n172 GND 0.04fF
C734 VDD.n173 GND 0.03fF
C735 VDD.n174 GND 0.02fF
C736 VDD.n175 GND 0.02fF
C737 VDD.n176 GND 0.02fF
C738 VDD.n177 GND 0.03fF
C739 VDD.n178 GND 0.02fF
C740 VDD.n180 GND 0.02fF
C741 VDD.n181 GND 0.02fF
C742 VDD.n182 GND 0.02fF
C743 VDD.n184 GND 0.28fF
C744 VDD.n186 GND 0.02fF
C745 VDD.n187 GND 0.02fF
C746 VDD.n188 GND 0.03fF
C747 VDD.n189 GND 0.02fF
C748 VDD.n190 GND 0.28fF
C749 VDD.n191 GND 0.01fF
C750 VDD.n192 GND 0.02fF
C751 VDD.n193 GND 0.03fF
C752 VDD.n194 GND 0.28fF
C753 VDD.n195 GND 0.01fF
C754 VDD.n196 GND 0.02fF
C755 VDD.n197 GND 0.02fF
C756 VDD.n198 GND 0.22fF
C757 VDD.n199 GND 0.01fF
C758 VDD.n200 GND 0.07fF
C759 VDD.n201 GND 0.02fF
C760 VDD.n202 GND 0.14fF
C761 VDD.n203 GND 0.17fF
C762 VDD.n204 GND 0.01fF
C763 VDD.n205 GND 0.02fF
C764 VDD.n206 GND 0.02fF
C765 VDD.n207 GND 0.14fF
C766 VDD.n208 GND 0.16fF
C767 VDD.n209 GND 0.01fF
C768 VDD.n210 GND 0.11fF
C769 VDD.n211 GND 0.02fF
C770 VDD.n212 GND 0.02fF
C771 VDD.n213 GND 0.02fF
C772 VDD.n214 GND 0.18fF
C773 VDD.n215 GND 0.15fF
C774 VDD.n216 GND 0.01fF
C775 VDD.n217 GND 0.02fF
C776 VDD.n218 GND 0.03fF
C777 VDD.n219 GND 0.18fF
C778 VDD.n220 GND 0.15fF
C779 VDD.n221 GND 0.01fF
C780 VDD.n222 GND 0.02fF
C781 VDD.n223 GND 0.03fF
C782 VDD.n224 GND 0.11fF
C783 VDD.n225 GND 0.02fF
C784 VDD.n226 GND 0.14fF
C785 VDD.n227 GND 0.16fF
C786 VDD.n228 GND 0.01fF
C787 VDD.n229 GND 0.02fF
C788 VDD.n230 GND 0.02fF
C789 VDD.n231 GND 0.14fF
C790 VDD.n232 GND 0.17fF
C791 VDD.n233 GND 0.01fF
C792 VDD.n234 GND 0.02fF
C793 VDD.n235 GND 0.02fF
C794 VDD.n236 GND 0.06fF
C795 VDD.n237 GND 0.23fF
C796 VDD.n238 GND 0.01fF
C797 VDD.n239 GND 0.01fF
C798 VDD.n240 GND 0.02fF
C799 VDD.n241 GND 0.28fF
C800 VDD.n242 GND 0.01fF
C801 VDD.n243 GND 0.02fF
C802 VDD.n244 GND 0.02fF
C803 VDD.n245 GND 0.28fF
C804 VDD.n246 GND 0.01fF
C805 VDD.n247 GND 0.02fF
C806 VDD.n248 GND 0.03fF
C807 VDD.n249 GND 0.02fF
C808 VDD.n250 GND 0.02fF
C809 VDD.n251 GND 0.02fF
C810 VDD.n252 GND 0.26fF
C811 VDD.n253 GND 0.04fF
C812 VDD.n254 GND 0.03fF
C813 VDD.n255 GND 0.02fF
C814 VDD.n256 GND 0.02fF
C815 VDD.n257 GND 0.02fF
C816 VDD.n258 GND 0.03fF
C817 VDD.n259 GND 0.02fF
C818 VDD.n261 GND 0.02fF
C819 VDD.n262 GND 0.02fF
C820 VDD.n263 GND 0.02fF
C821 VDD.n265 GND 0.28fF
C822 VDD.n267 GND 0.02fF
C823 VDD.n268 GND 0.02fF
C824 VDD.n269 GND 0.03fF
C825 VDD.n270 GND 0.02fF
C826 VDD.n271 GND 0.28fF
C827 VDD.n272 GND 0.01fF
C828 VDD.n273 GND 0.02fF
C829 VDD.n274 GND 0.03fF
C830 VDD.n275 GND 0.06fF
C831 VDD.n276 GND 0.24fF
C832 VDD.n277 GND 0.01fF
C833 VDD.n278 GND 0.01fF
C834 VDD.n279 GND 0.02fF
C835 VDD.n280 GND 0.14fF
C836 VDD.n281 GND 0.17fF
C837 VDD.n282 GND 0.01fF
C838 VDD.n283 GND 0.02fF
C839 VDD.n284 GND 0.02fF
C840 VDD.n285 GND 0.11fF
C841 VDD.n286 GND 0.03fF
C842 VDD.n287 GND 0.31fF
C843 VDD.n288 GND 0.01fF
C844 VDD.n289 GND 0.02fF
C845 VDD.n290 GND 0.03fF
C846 VDD.n291 GND 0.17fF
C847 VDD.n292 GND 0.14fF
C848 VDD.n293 GND 0.01fF
C849 VDD.n294 GND 0.02fF
C850 VDD.n295 GND 0.03fF
C851 VDD.n296 GND 0.14fF
C852 VDD.n297 GND 0.16fF
C853 VDD.n298 GND 0.01fF
C854 VDD.n299 GND 0.02fF
C855 VDD.n300 GND 0.02fF
C856 VDD.n301 GND 0.06fF
C857 VDD.n302 GND 0.25fF
C858 VDD.n303 GND 0.01fF
C859 VDD.n304 GND 0.01fF
C860 VDD.n305 GND 0.02fF
C861 VDD.n306 GND 0.28fF
C862 VDD.n307 GND 0.01fF
C863 VDD.n308 GND 0.02fF
C864 VDD.n309 GND 0.03fF
C865 VDD.n310 GND 0.02fF
C866 VDD.n311 GND 0.02fF
C867 VDD.n312 GND 0.02fF
C868 VDD.n313 GND 0.22fF
C869 VDD.n314 GND 0.04fF
C870 VDD.n315 GND 0.03fF
C871 VDD.n316 GND 0.02fF
C872 VDD.n317 GND 0.02fF
C873 VDD.n318 GND 0.02fF
C874 VDD.n319 GND 0.03fF
C875 VDD.n320 GND 0.02fF
C876 VDD.n322 GND 0.02fF
C877 VDD.n323 GND 0.02fF
C878 VDD.n324 GND 0.02fF
C879 VDD.n326 GND 0.28fF
C880 VDD.n328 GND 0.02fF
C881 VDD.n329 GND 0.02fF
C882 VDD.n330 GND 0.03fF
C883 VDD.n331 GND 0.02fF
C884 VDD.n332 GND 0.28fF
C885 VDD.n333 GND 0.01fF
C886 VDD.n334 GND 0.02fF
C887 VDD.n335 GND 0.03fF
C888 VDD.n336 GND 0.06fF
C889 VDD.n337 GND 0.24fF
C890 VDD.n338 GND 0.01fF
C891 VDD.n339 GND 0.01fF
C892 VDD.n340 GND 0.02fF
C893 VDD.n341 GND 0.14fF
C894 VDD.n342 GND 0.17fF
C895 VDD.n343 GND 0.01fF
C896 VDD.n344 GND 0.02fF
C897 VDD.n345 GND 0.02fF
C898 VDD.n346 GND 0.11fF
C899 VDD.n347 GND 0.03fF
C900 VDD.n348 GND 0.31fF
C901 VDD.n349 GND 0.01fF
C902 VDD.n350 GND 0.02fF
C903 VDD.n351 GND 0.03fF
C904 VDD.n352 GND 0.17fF
C905 VDD.n353 GND 0.14fF
C906 VDD.n354 GND 0.01fF
C907 VDD.n355 GND 0.02fF
C908 VDD.n356 GND 0.03fF
C909 VDD.n357 GND 0.14fF
C910 VDD.n358 GND 0.16fF
C911 VDD.n359 GND 0.01fF
C912 VDD.n360 GND 0.02fF
C913 VDD.n361 GND 0.02fF
C914 VDD.n362 GND 0.06fF
C915 VDD.n363 GND 0.25fF
C916 VDD.n364 GND 0.01fF
C917 VDD.n365 GND 0.01fF
C918 VDD.n366 GND 0.02fF
C919 VDD.n367 GND 0.28fF
C920 VDD.n368 GND 0.01fF
C921 VDD.n369 GND 0.02fF
C922 VDD.n370 GND 0.03fF
C923 VDD.n371 GND 0.02fF
C924 VDD.n372 GND 0.02fF
C925 VDD.n373 GND 0.02fF
C926 VDD.n374 GND 0.26fF
C927 VDD.n375 GND 0.04fF
C928 VDD.n376 GND 0.03fF
C929 VDD.n377 GND 0.02fF
C930 VDD.n378 GND 0.02fF
C931 VDD.n379 GND 0.02fF
C932 VDD.n380 GND 0.03fF
C933 VDD.n381 GND 0.02fF
C934 VDD.n383 GND 0.02fF
C935 VDD.n384 GND 0.02fF
C936 VDD.n385 GND 0.02fF
C937 VDD.n387 GND 0.28fF
C938 VDD.n389 GND 0.02fF
C939 VDD.n390 GND 0.02fF
C940 VDD.n391 GND 0.03fF
C941 VDD.n392 GND 0.02fF
C942 VDD.n393 GND 0.28fF
C943 VDD.n394 GND 0.01fF
C944 VDD.n395 GND 0.02fF
C945 VDD.n396 GND 0.03fF
C946 VDD.n397 GND 0.28fF
C947 VDD.n398 GND 0.01fF
C948 VDD.n399 GND 0.02fF
C949 VDD.n400 GND 0.02fF
C950 VDD.n401 GND 0.22fF
C951 VDD.n402 GND 0.01fF
C952 VDD.n403 GND 0.07fF
C953 VDD.n404 GND 0.02fF
C954 VDD.n405 GND 0.14fF
C955 VDD.n406 GND 0.17fF
C956 VDD.n407 GND 0.01fF
C957 VDD.n408 GND 0.02fF
C958 VDD.n409 GND 0.02fF
C959 VDD.n410 GND 0.14fF
C960 VDD.n411 GND 0.16fF
C961 VDD.n412 GND 0.01fF
C962 VDD.n413 GND 0.11fF
C963 VDD.n414 GND 0.02fF
C964 VDD.n415 GND 0.02fF
C965 VDD.n416 GND 0.02fF
C966 VDD.n417 GND 0.18fF
C967 VDD.n418 GND 0.15fF
C968 VDD.n419 GND 0.01fF
C969 VDD.n420 GND 0.02fF
C970 VDD.n421 GND 0.03fF
C971 VDD.n422 GND 0.18fF
C972 VDD.n423 GND 0.15fF
C973 VDD.n424 GND 0.01fF
C974 VDD.n425 GND 0.02fF
C975 VDD.n426 GND 0.03fF
C976 VDD.n427 GND 0.11fF
C977 VDD.n428 GND 0.02fF
C978 VDD.n429 GND 0.14fF
C979 VDD.n430 GND 0.16fF
C980 VDD.n431 GND 0.01fF
C981 VDD.n432 GND 0.02fF
C982 VDD.n433 GND 0.02fF
C983 VDD.n434 GND 0.14fF
C984 VDD.n435 GND 0.17fF
C985 VDD.n436 GND 0.01fF
C986 VDD.n437 GND 0.02fF
C987 VDD.n438 GND 0.02fF
C988 VDD.n439 GND 0.06fF
C989 VDD.n440 GND 0.23fF
C990 VDD.n441 GND 0.01fF
C991 VDD.n442 GND 0.01fF
C992 VDD.n443 GND 0.02fF
C993 VDD.n444 GND 0.28fF
C994 VDD.n445 GND 0.01fF
C995 VDD.n446 GND 0.02fF
C996 VDD.n447 GND 0.02fF
C997 VDD.n448 GND 0.28fF
C998 VDD.n449 GND 0.01fF
C999 VDD.n450 GND 0.02fF
C1000 VDD.n451 GND 0.03fF
C1001 VDD.n452 GND 0.02fF
C1002 VDD.n453 GND 0.02fF
C1003 VDD.n454 GND 0.02fF
C1004 VDD.n455 GND 0.31fF
C1005 VDD.n456 GND 0.04fF
C1006 VDD.n457 GND 0.03fF
C1007 VDD.n458 GND 0.02fF
C1008 VDD.n459 GND 0.02fF
C1009 VDD.n460 GND 0.02fF
C1010 VDD.n461 GND 0.03fF
C1011 VDD.n462 GND 0.02fF
C1012 VDD.n464 GND 0.02fF
C1013 VDD.n465 GND 0.02fF
C1014 VDD.n466 GND 0.02fF
C1015 VDD.n468 GND 0.28fF
C1016 VDD.n470 GND 0.02fF
C1017 VDD.n471 GND 0.02fF
C1018 VDD.n472 GND 0.03fF
C1019 VDD.n473 GND 0.02fF
C1020 VDD.n474 GND 0.28fF
C1021 VDD.n475 GND 0.01fF
C1022 VDD.n476 GND 0.02fF
C1023 VDD.n477 GND 0.03fF
C1024 VDD.n478 GND 0.28fF
C1025 VDD.n479 GND 0.01fF
C1026 VDD.n480 GND 0.02fF
C1027 VDD.n481 GND 0.02fF
C1028 VDD.n482 GND 0.22fF
C1029 VDD.n483 GND 0.01fF
C1030 VDD.n484 GND 0.07fF
C1031 VDD.n485 GND 0.02fF
C1032 VDD.n486 GND 0.14fF
C1033 VDD.n487 GND 0.17fF
C1034 VDD.n488 GND 0.01fF
C1035 VDD.n489 GND 0.02fF
C1036 VDD.n490 GND 0.02fF
C1037 VDD.n491 GND 0.14fF
C1038 VDD.n492 GND 0.16fF
C1039 VDD.n493 GND 0.01fF
C1040 VDD.n494 GND 0.11fF
C1041 VDD.n495 GND 0.02fF
C1042 VDD.n496 GND 0.02fF
C1043 VDD.n497 GND 0.02fF
C1044 VDD.n498 GND 0.18fF
C1045 VDD.n499 GND 0.15fF
C1046 VDD.n500 GND 0.01fF
C1047 VDD.n501 GND 0.02fF
C1048 VDD.n502 GND 0.03fF
C1049 VDD.n503 GND 0.18fF
C1050 VDD.n504 GND 0.15fF
C1051 VDD.n505 GND 0.01fF
C1052 VDD.n506 GND 0.02fF
C1053 VDD.n507 GND 0.03fF
C1054 VDD.n508 GND 0.11fF
C1055 VDD.n509 GND 0.02fF
C1056 VDD.n510 GND 0.14fF
C1057 VDD.n511 GND 0.16fF
C1058 VDD.n512 GND 0.01fF
C1059 VDD.n513 GND 0.02fF
C1060 VDD.n514 GND 0.02fF
C1061 VDD.n515 GND 0.14fF
C1062 VDD.n516 GND 0.17fF
C1063 VDD.n517 GND 0.01fF
C1064 VDD.n518 GND 0.02fF
C1065 VDD.n519 GND 0.02fF
C1066 VDD.n520 GND 0.06fF
C1067 VDD.n521 GND 0.23fF
C1068 VDD.n522 GND 0.01fF
C1069 VDD.n523 GND 0.01fF
C1070 VDD.n524 GND 0.02fF
C1071 VDD.n525 GND 0.28fF
C1072 VDD.n526 GND 0.01fF
C1073 VDD.n527 GND 0.02fF
C1074 VDD.n528 GND 0.02fF
C1075 VDD.n529 GND 0.28fF
C1076 VDD.n530 GND 0.01fF
C1077 VDD.n531 GND 0.02fF
C1078 VDD.n532 GND 0.03fF
C1079 VDD.n533 GND 0.02fF
C1080 VDD.n534 GND 0.02fF
C1081 VDD.n535 GND 0.02fF
C1082 VDD.n536 GND 0.26fF
C1083 VDD.n537 GND 0.04fF
C1084 VDD.n538 GND 0.03fF
C1085 VDD.n539 GND 0.02fF
C1086 VDD.n540 GND 0.02fF
C1087 VDD.n541 GND 0.02fF
C1088 VDD.n542 GND 0.03fF
C1089 VDD.n543 GND 0.02fF
C1090 VDD.n545 GND 0.02fF
C1091 VDD.n546 GND 0.02fF
C1092 VDD.n547 GND 0.02fF
C1093 VDD.n549 GND 0.28fF
C1094 VDD.n551 GND 0.02fF
C1095 VDD.n552 GND 0.02fF
C1096 VDD.n553 GND 0.03fF
C1097 VDD.n554 GND 0.02fF
C1098 VDD.n555 GND 0.28fF
C1099 VDD.n556 GND 0.01fF
C1100 VDD.n557 GND 0.02fF
C1101 VDD.n558 GND 0.03fF
C1102 VDD.n559 GND 0.06fF
C1103 VDD.n560 GND 0.24fF
C1104 VDD.n561 GND 0.01fF
C1105 VDD.n562 GND 0.01fF
C1106 VDD.n563 GND 0.02fF
C1107 VDD.n564 GND 0.14fF
C1108 VDD.n565 GND 0.17fF
C1109 VDD.n566 GND 0.01fF
C1110 VDD.n567 GND 0.02fF
C1111 VDD.n568 GND 0.02fF
C1112 VDD.n569 GND 0.11fF
C1113 VDD.n570 GND 0.03fF
C1114 VDD.n571 GND 0.31fF
C1115 VDD.n572 GND 0.01fF
C1116 VDD.n573 GND 0.02fF
C1117 VDD.n574 GND 0.03fF
C1118 VDD.n575 GND 0.17fF
C1119 VDD.n576 GND 0.14fF
C1120 VDD.n577 GND 0.01fF
C1121 VDD.n578 GND 0.02fF
C1122 VDD.n579 GND 0.03fF
C1123 VDD.n580 GND 0.14fF
C1124 VDD.n581 GND 0.16fF
C1125 VDD.n582 GND 0.01fF
C1126 VDD.n583 GND 0.02fF
C1127 VDD.n584 GND 0.02fF
C1128 VDD.n585 GND 0.06fF
C1129 VDD.n586 GND 0.25fF
C1130 VDD.n587 GND 0.01fF
C1131 VDD.n588 GND 0.01fF
C1132 VDD.n589 GND 0.02fF
C1133 VDD.n590 GND 0.28fF
C1134 VDD.n591 GND 0.01fF
C1135 VDD.n592 GND 0.02fF
C1136 VDD.n593 GND 0.03fF
C1137 VDD.n594 GND 0.02fF
C1138 VDD.n595 GND 0.02fF
C1139 VDD.n596 GND 0.02fF
C1140 VDD.n597 GND 0.26fF
C1141 VDD.n598 GND 0.04fF
C1142 VDD.n599 GND 0.03fF
C1143 VDD.n600 GND 0.02fF
C1144 VDD.n601 GND 0.02fF
C1145 VDD.n602 GND 0.02fF
C1146 VDD.n603 GND 0.03fF
C1147 VDD.n604 GND 0.02fF
C1148 VDD.n606 GND 0.02fF
C1149 VDD.n607 GND 0.02fF
C1150 VDD.n608 GND 0.02fF
C1151 VDD.n610 GND 0.28fF
C1152 VDD.n612 GND 0.02fF
C1153 VDD.n613 GND 0.02fF
C1154 VDD.n614 GND 0.03fF
C1155 VDD.n615 GND 0.02fF
C1156 VDD.n616 GND 0.28fF
C1157 VDD.n617 GND 0.01fF
C1158 VDD.n618 GND 0.02fF
C1159 VDD.n619 GND 0.03fF
C1160 VDD.n620 GND 0.28fF
C1161 VDD.n621 GND 0.01fF
C1162 VDD.n622 GND 0.02fF
C1163 VDD.n623 GND 0.02fF
C1164 VDD.n624 GND 0.22fF
C1165 VDD.n625 GND 0.01fF
C1166 VDD.n626 GND 0.07fF
C1167 VDD.n627 GND 0.02fF
C1168 VDD.n628 GND 0.14fF
C1169 VDD.n629 GND 0.17fF
C1170 VDD.n630 GND 0.01fF
C1171 VDD.n631 GND 0.02fF
C1172 VDD.n632 GND 0.02fF
C1173 VDD.n633 GND 0.14fF
C1174 VDD.n634 GND 0.16fF
C1175 VDD.n635 GND 0.01fF
C1176 VDD.n636 GND 0.11fF
C1177 VDD.n637 GND 0.02fF
C1178 VDD.n638 GND 0.02fF
C1179 VDD.n639 GND 0.02fF
C1180 VDD.n640 GND 0.18fF
C1181 VDD.n641 GND 0.15fF
C1182 VDD.n642 GND 0.01fF
C1183 VDD.n643 GND 0.02fF
C1184 VDD.n644 GND 0.03fF
C1185 VDD.n645 GND 0.18fF
C1186 VDD.n646 GND 0.15fF
C1187 VDD.n647 GND 0.01fF
C1188 VDD.n648 GND 0.02fF
C1189 VDD.n649 GND 0.03fF
C1190 VDD.n650 GND 0.11fF
C1191 VDD.n651 GND 0.02fF
C1192 VDD.n652 GND 0.14fF
C1193 VDD.n653 GND 0.16fF
C1194 VDD.n654 GND 0.01fF
C1195 VDD.n655 GND 0.02fF
C1196 VDD.n656 GND 0.02fF
C1197 VDD.n657 GND 0.14fF
C1198 VDD.n658 GND 0.17fF
C1199 VDD.n659 GND 0.01fF
C1200 VDD.n660 GND 0.02fF
C1201 VDD.n661 GND 0.02fF
C1202 VDD.n662 GND 0.06fF
C1203 VDD.n663 GND 0.23fF
C1204 VDD.n664 GND 0.01fF
C1205 VDD.n665 GND 0.01fF
C1206 VDD.n666 GND 0.02fF
C1207 VDD.n667 GND 0.28fF
C1208 VDD.n668 GND 0.01fF
C1209 VDD.n669 GND 0.02fF
C1210 VDD.n670 GND 0.02fF
C1211 VDD.n671 GND 0.28fF
C1212 VDD.n672 GND 0.01fF
C1213 VDD.n673 GND 0.02fF
C1214 VDD.n674 GND 0.03fF
C1215 VDD.n675 GND 0.02fF
C1216 VDD.n676 GND 0.02fF
C1217 VDD.n677 GND 0.02fF
C1218 VDD.n678 GND 0.26fF
C1219 VDD.n679 GND 0.04fF
C1220 VDD.n680 GND 0.03fF
C1221 VDD.n681 GND 0.02fF
C1222 VDD.n682 GND 0.02fF
C1223 VDD.n683 GND 0.02fF
C1224 VDD.n684 GND 0.03fF
C1225 VDD.n685 GND 0.02fF
C1226 VDD.n687 GND 0.02fF
C1227 VDD.n688 GND 0.02fF
C1228 VDD.n689 GND 0.02fF
C1229 VDD.n691 GND 0.28fF
C1230 VDD.n693 GND 0.02fF
C1231 VDD.n694 GND 0.02fF
C1232 VDD.n695 GND 0.03fF
C1233 VDD.n696 GND 0.02fF
C1234 VDD.n697 GND 0.28fF
C1235 VDD.n698 GND 0.01fF
C1236 VDD.n699 GND 0.02fF
C1237 VDD.n700 GND 0.03fF
C1238 VDD.n701 GND 0.06fF
C1239 VDD.n702 GND 0.24fF
C1240 VDD.n703 GND 0.01fF
C1241 VDD.n704 GND 0.01fF
C1242 VDD.n705 GND 0.02fF
C1243 VDD.n706 GND 0.14fF
C1244 VDD.n707 GND 0.17fF
C1245 VDD.n708 GND 0.01fF
C1246 VDD.n709 GND 0.02fF
C1247 VDD.n710 GND 0.02fF
C1248 VDD.n711 GND 0.11fF
C1249 VDD.n712 GND 0.03fF
C1250 VDD.n713 GND 0.31fF
C1251 VDD.n714 GND 0.01fF
C1252 VDD.n715 GND 0.02fF
C1253 VDD.n716 GND 0.03fF
C1254 VDD.n717 GND 0.17fF
C1255 VDD.n718 GND 0.14fF
C1256 VDD.n719 GND 0.01fF
C1257 VDD.n720 GND 0.02fF
C1258 VDD.n721 GND 0.03fF
C1259 VDD.n722 GND 0.14fF
C1260 VDD.n723 GND 0.16fF
C1261 VDD.n724 GND 0.01fF
C1262 VDD.n725 GND 0.02fF
C1263 VDD.n726 GND 0.02fF
C1264 VDD.n727 GND 0.02fF
C1265 VDD.n728 GND 0.02fF
C1266 VDD.n729 GND 0.02fF
C1267 VDD.n730 GND 0.15fF
C1268 VDD.n731 GND 0.03fF
C1269 VDD.n732 GND 0.02fF
C1270 VDD.n733 GND 0.02fF
C1271 VDD.n734 GND 0.02fF
C1272 VDD.n735 GND 0.03fF
C1273 VDD.n736 GND 0.02fF
C1274 VDD.n738 GND 0.02fF
C1275 VDD.n739 GND 0.02fF
C1276 VDD.n740 GND 0.02fF
C1277 VDD.n742 GND 0.46fF
C1278 VDD.n744 GND 0.03fF
C1279 VDD.n745 GND 0.04fF
C1280 VDD.n746 GND 0.28fF
C1281 VDD.n747 GND 0.02fF
C1282 VDD.n748 GND 0.03fF
C1283 VDD.n749 GND 0.03fF
C1284 VDD.n750 GND 0.06fF
C1285 VDD.n751 GND 0.25fF
C1286 VDD.n752 GND 0.01fF
C1287 VDD.n753 GND 0.01fF
C1288 VDD.n754 GND 0.02fF
C1289 VDD.n755 GND 0.14fF
C1290 VDD.n756 GND 0.16fF
C1291 VDD.n757 GND 0.01fF
C1292 VDD.n758 GND 0.02fF
C1293 VDD.n759 GND 0.02fF
C1294 VDD.n760 GND 0.17fF
C1295 VDD.n761 GND 0.14fF
C1296 VDD.n762 GND 0.01fF
C1297 VDD.n763 GND 0.02fF
C1298 VDD.n764 GND 0.03fF
C1299 VDD.n765 GND 0.11fF
C1300 VDD.n766 GND 0.03fF
C1301 VDD.n767 GND 0.31fF
C1302 VDD.n768 GND 0.01fF
C1303 VDD.n769 GND 0.02fF
C1304 VDD.n770 GND 0.03fF
C1305 VDD.n771 GND 0.14fF
C1306 VDD.n772 GND 0.17fF
C1307 VDD.n773 GND 0.01fF
C1308 VDD.n774 GND 0.02fF
C1309 VDD.n775 GND 0.02fF
C1310 VDD.n776 GND 0.06fF
C1311 VDD.n777 GND 0.24fF
C1312 VDD.n778 GND 0.01fF
C1313 VDD.n779 GND 0.01fF
C1314 VDD.n780 GND 0.02fF
C1315 VDD.n781 GND 0.28fF
C1316 VDD.n782 GND 0.01fF
C1317 VDD.n783 GND 0.02fF
C1318 VDD.n784 GND 0.03fF
C1319 VDD.n785 GND 0.02fF
C1320 VDD.n786 GND 0.02fF
C1321 VDD.n787 GND 0.02fF
C1322 VDD.n788 GND 0.02fF
C1323 VDD.n789 GND 0.02fF
C1324 VDD.n790 GND 0.02fF
C1325 VDD.n792 GND 0.02fF
C1326 VDD.n793 GND 0.02fF
C1327 VDD.n794 GND 0.02fF
C1328 VDD.n795 GND 0.02fF
C1329 VDD.n797 GND 0.04fF
C1330 VDD.n798 GND 0.02fF
C1331 VDD.n799 GND 0.27fF
C1332 VDD.n800 GND 0.04fF
C1333 VDD.n802 GND 0.28fF
C1334 VDD.n804 GND 0.02fF
C1335 VDD.n805 GND 0.02fF
C1336 VDD.n806 GND 0.03fF
C1337 VDD.n807 GND 0.02fF
C1338 VDD.n808 GND 0.28fF
C1339 VDD.n809 GND 0.01fF
C1340 VDD.n810 GND 0.02fF
C1341 VDD.n811 GND 0.03fF
C1342 VDD.n812 GND 0.28fF
C1343 VDD.n813 GND 0.01fF
C1344 VDD.n814 GND 0.02fF
C1345 VDD.n815 GND 0.02fF
C1346 VDD.n816 GND 0.06fF
C1347 VDD.n817 GND 0.23fF
C1348 VDD.n818 GND 0.01fF
C1349 VDD.n819 GND 0.01fF
C1350 VDD.n820 GND 0.02fF
C1351 VDD.n821 GND 0.14fF
C1352 VDD.n822 GND 0.17fF
C1353 VDD.n823 GND 0.01fF
C1354 VDD.n824 GND 0.02fF
C1355 VDD.n825 GND 0.02fF
C1356 VDD.n826 GND 0.11fF
C1357 VDD.n827 GND 0.02fF
C1358 VDD.n828 GND 0.14fF
C1359 VDD.n829 GND 0.16fF
C1360 VDD.n830 GND 0.01fF
C1361 VDD.n831 GND 0.02fF
C1362 VDD.n832 GND 0.02fF
C1363 VDD.n833 GND 0.18fF
C1364 VDD.n834 GND 0.15fF
C1365 VDD.n835 GND 0.01fF
C1366 VDD.n836 GND 0.02fF
C1367 VDD.n837 GND 0.03fF
C1368 VDD.n838 GND 0.18fF
C1369 VDD.n839 GND 0.15fF
C1370 VDD.n840 GND 0.01fF
C1371 VDD.n841 GND 0.02fF
C1372 VDD.n842 GND 0.03fF
C1373 VDD.n843 GND 0.14fF
C1374 VDD.n844 GND 0.16fF
C1375 VDD.n845 GND 0.01fF
C1376 VDD.n846 GND 0.11fF
C1377 VDD.n847 GND 0.02fF
C1378 VDD.n848 GND 0.02fF
C1379 VDD.n849 GND 0.02fF
C1380 VDD.n850 GND 0.14fF
C1381 VDD.n851 GND 0.17fF
C1382 VDD.n852 GND 0.01fF
C1383 VDD.n853 GND 0.02fF
C1384 VDD.n854 GND 0.02fF
C1385 VDD.n855 GND 0.22fF
C1386 VDD.n856 GND 0.01fF
C1387 VDD.n857 GND 0.07fF
C1388 VDD.n858 GND 0.02fF
C1389 VDD.n859 GND 0.28fF
C1390 VDD.n860 GND 0.01fF
C1391 VDD.n861 GND 0.02fF
C1392 VDD.n862 GND 0.02fF
C1393 VDD.n863 GND 0.28fF
C1394 VDD.n864 GND 0.01fF
C1395 VDD.n865 GND 0.02fF
C1396 VDD.n866 GND 0.03fF
C1397 VDD.n867 GND 0.02fF
C1398 VDD.n868 GND 0.02fF
C1399 VDD.n869 GND 0.02fF
C1400 VDD.n870 GND 0.31fF
C1401 VDD.n871 GND 0.04fF
C1402 VDD.n872 GND 0.03fF
C1403 VDD.n873 GND 0.02fF
C1404 VDD.n874 GND 0.02fF
C1405 VDD.n875 GND 0.02fF
C1406 VDD.n876 GND 0.03fF
C1407 VDD.n877 GND 0.02fF
C1408 VDD.n879 GND 0.02fF
C1409 VDD.n880 GND 0.02fF
C1410 VDD.n881 GND 0.02fF
C1411 VDD.n883 GND 0.28fF
C1412 VDD.n885 GND 0.02fF
C1413 VDD.n886 GND 0.02fF
C1414 VDD.n887 GND 0.03fF
C1415 VDD.n888 GND 0.02fF
C1416 VDD.n889 GND 0.28fF
C1417 VDD.n890 GND 0.01fF
C1418 VDD.n891 GND 0.02fF
C1419 VDD.n892 GND 0.03fF
C1420 VDD.n893 GND 0.28fF
C1421 VDD.n894 GND 0.01fF
C1422 VDD.n895 GND 0.02fF
C1423 VDD.n896 GND 0.02fF
C1424 VDD.n897 GND 0.06fF
C1425 VDD.n898 GND 0.23fF
C1426 VDD.n899 GND 0.01fF
C1427 VDD.n900 GND 0.01fF
C1428 VDD.n901 GND 0.02fF
C1429 VDD.n902 GND 0.14fF
C1430 VDD.n903 GND 0.17fF
C1431 VDD.n904 GND 0.01fF
C1432 VDD.n905 GND 0.02fF
C1433 VDD.n906 GND 0.02fF
C1434 VDD.n907 GND 0.11fF
C1435 VDD.n908 GND 0.02fF
C1436 VDD.n909 GND 0.14fF
C1437 VDD.n910 GND 0.16fF
C1438 VDD.n911 GND 0.01fF
C1439 VDD.n912 GND 0.02fF
C1440 VDD.n913 GND 0.02fF
C1441 VDD.n914 GND 0.18fF
C1442 VDD.n915 GND 0.15fF
C1443 VDD.n916 GND 0.01fF
C1444 VDD.n917 GND 0.02fF
C1445 VDD.n918 GND 0.03fF
C1446 VDD.n919 GND 0.18fF
C1447 VDD.n920 GND 0.15fF
C1448 VDD.n921 GND 0.01fF
C1449 VDD.n922 GND 0.02fF
C1450 VDD.n923 GND 0.03fF
C1451 VDD.n924 GND 0.14fF
C1452 VDD.n925 GND 0.16fF
C1453 VDD.n926 GND 0.01fF
C1454 VDD.n927 GND 0.11fF
C1455 VDD.n928 GND 0.02fF
C1456 VDD.n929 GND 0.02fF
C1457 VDD.n930 GND 0.02fF
C1458 VDD.n931 GND 0.14fF
C1459 VDD.n932 GND 0.17fF
C1460 VDD.n933 GND 0.01fF
C1461 VDD.n934 GND 0.02fF
C1462 VDD.n935 GND 0.02fF
C1463 VDD.n936 GND 0.22fF
C1464 VDD.n937 GND 0.01fF
C1465 VDD.n938 GND 0.07fF
C1466 VDD.n939 GND 0.02fF
C1467 VDD.n940 GND 0.28fF
C1468 VDD.n941 GND 0.01fF
C1469 VDD.n942 GND 0.02fF
C1470 VDD.n943 GND 0.02fF
C1471 VDD.n944 GND 0.28fF
C1472 VDD.n945 GND 0.01fF
C1473 VDD.n946 GND 0.02fF
C1474 VDD.n947 GND 0.03fF
C1475 VDD.n948 GND 0.02fF
C1476 VDD.n949 GND 0.02fF
C1477 VDD.n950 GND 0.02fF
C1478 VDD.n951 GND 0.26fF
C1479 VDD.n952 GND 0.04fF
C1480 VDD.n953 GND 0.03fF
C1481 VDD.n954 GND 0.02fF
C1482 VDD.n955 GND 0.02fF
C1483 VDD.n956 GND 0.02fF
C1484 VDD.n957 GND 0.03fF
C1485 VDD.n958 GND 0.02fF
C1486 VDD.n960 GND 0.02fF
C1487 VDD.n961 GND 0.02fF
C1488 VDD.n962 GND 0.02fF
C1489 VDD.n964 GND 0.28fF
C1490 VDD.n966 GND 0.02fF
C1491 VDD.n967 GND 0.02fF
C1492 VDD.n968 GND 0.03fF
C1493 VDD.n969 GND 0.02fF
C1494 VDD.n970 GND 0.28fF
C1495 VDD.n971 GND 0.01fF
C1496 VDD.n972 GND 0.02fF
C1497 VDD.n973 GND 0.03fF
C1498 VDD.n974 GND 0.06fF
C1499 VDD.n975 GND 0.25fF
C1500 VDD.n976 GND 0.01fF
C1501 VDD.n977 GND 0.01fF
C1502 VDD.n978 GND 0.02fF
C1503 VDD.n979 GND 0.14fF
C1504 VDD.n980 GND 0.16fF
C1505 VDD.n981 GND 0.01fF
C1506 VDD.n982 GND 0.02fF
C1507 VDD.n983 GND 0.02fF
C1508 VDD.n984 GND 0.17fF
C1509 VDD.n985 GND 0.14fF
C1510 VDD.n986 GND 0.01fF
C1511 VDD.n987 GND 0.02fF
C1512 VDD.n988 GND 0.03fF
C1513 VDD.n989 GND 0.11fF
C1514 VDD.n990 GND 0.03fF
C1515 VDD.n991 GND 0.31fF
C1516 VDD.n992 GND 0.01fF
C1517 VDD.n993 GND 0.02fF
C1518 VDD.n994 GND 0.03fF
C1519 VDD.n995 GND 0.14fF
C1520 VDD.n996 GND 0.17fF
C1521 VDD.n997 GND 0.01fF
C1522 VDD.n998 GND 0.02fF
C1523 VDD.n999 GND 0.02fF
C1524 VDD.n1000 GND 0.06fF
C1525 VDD.n1001 GND 0.24fF
C1526 VDD.n1002 GND 0.01fF
C1527 VDD.n1003 GND 0.01fF
C1528 VDD.n1004 GND 0.02fF
C1529 VDD.n1005 GND 0.28fF
C1530 VDD.n1006 GND 0.01fF
C1531 VDD.n1007 GND 0.02fF
C1532 VDD.n1008 GND 0.03fF
C1533 VDD.n1009 GND 0.02fF
C1534 VDD.n1010 GND 0.02fF
C1535 VDD.n1011 GND 0.02fF
C1536 VDD.n1012 GND 0.22fF
C1537 VDD.n1013 GND 0.04fF
C1538 VDD.n1014 GND 0.03fF
C1539 VDD.n1015 GND 0.02fF
C1540 VDD.n1016 GND 0.02fF
C1541 VDD.n1017 GND 0.02fF
C1542 VDD.n1018 GND 0.03fF
C1543 VDD.n1019 GND 0.02fF
C1544 VDD.n1021 GND 0.02fF
C1545 VDD.n1022 GND 0.02fF
C1546 VDD.n1023 GND 0.02fF
C1547 VDD.n1025 GND 0.28fF
C1548 VDD.n1027 GND 0.02fF
C1549 VDD.n1028 GND 0.02fF
C1550 VDD.n1029 GND 0.03fF
C1551 VDD.n1030 GND 0.02fF
C1552 VDD.n1031 GND 0.28fF
C1553 VDD.n1032 GND 0.01fF
C1554 VDD.n1033 GND 0.02fF
C1555 VDD.n1034 GND 0.03fF
C1556 VDD.n1035 GND 0.06fF
C1557 VDD.n1036 GND 0.25fF
C1558 VDD.n1037 GND 0.01fF
C1559 VDD.n1038 GND 0.01fF
C1560 VDD.n1039 GND 0.02fF
C1561 VDD.n1040 GND 0.14fF
C1562 VDD.n1041 GND 0.16fF
C1563 VDD.n1042 GND 0.01fF
C1564 VDD.n1043 GND 0.02fF
C1565 VDD.n1044 GND 0.02fF
C1566 VDD.n1045 GND 0.17fF
C1567 VDD.n1046 GND 0.14fF
C1568 VDD.n1047 GND 0.01fF
C1569 VDD.n1048 GND 0.02fF
C1570 VDD.n1049 GND 0.03fF
C1571 VDD.n1050 GND 0.11fF
C1572 VDD.n1051 GND 0.03fF
C1573 VDD.n1052 GND 0.31fF
C1574 VDD.n1053 GND 0.01fF
C1575 VDD.n1054 GND 0.02fF
C1576 VDD.n1055 GND 0.03fF
C1577 VDD.n1056 GND 0.14fF
C1578 VDD.n1057 GND 0.17fF
C1579 VDD.n1058 GND 0.01fF
C1580 VDD.n1059 GND 0.02fF
C1581 VDD.n1060 GND 0.02fF
C1582 VDD.n1061 GND 0.06fF
C1583 VDD.n1062 GND 0.24fF
C1584 VDD.n1063 GND 0.01fF
C1585 VDD.n1064 GND 0.01fF
C1586 VDD.n1065 GND 0.02fF
C1587 VDD.n1066 GND 0.28fF
C1588 VDD.n1067 GND 0.01fF
C1589 VDD.n1068 GND 0.02fF
C1590 VDD.n1069 GND 0.03fF
C1591 VDD.n1070 GND 0.02fF
C1592 VDD.n1071 GND 0.02fF
C1593 VDD.n1072 GND 0.02fF
C1594 VDD.n1073 GND 0.26fF
C1595 VDD.n1074 GND 0.04fF
C1596 VDD.n1075 GND 0.03fF
C1597 VDD.n1076 GND 0.02fF
C1598 VDD.n1077 GND 0.02fF
C1599 VDD.n1078 GND 0.02fF
C1600 VDD.n1079 GND 0.03fF
C1601 VDD.n1080 GND 0.02fF
C1602 VDD.n1082 GND 0.02fF
C1603 VDD.n1083 GND 0.02fF
C1604 VDD.n1084 GND 0.02fF
C1605 VDD.n1086 GND 0.28fF
C1606 VDD.n1088 GND 0.02fF
C1607 VDD.n1089 GND 0.02fF
C1608 VDD.n1090 GND 0.03fF
C1609 VDD.n1091 GND 0.02fF
C1610 VDD.n1092 GND 0.28fF
C1611 VDD.n1093 GND 0.01fF
C1612 VDD.n1094 GND 0.02fF
C1613 VDD.n1095 GND 0.03fF
C1614 VDD.n1096 GND 0.28fF
C1615 VDD.n1097 GND 0.01fF
C1616 VDD.n1098 GND 0.02fF
C1617 VDD.n1099 GND 0.02fF
C1618 VDD.n1100 GND 0.06fF
C1619 VDD.n1101 GND 0.23fF
C1620 VDD.n1102 GND 0.01fF
C1621 VDD.n1103 GND 0.01fF
C1622 VDD.n1104 GND 0.02fF
C1623 VDD.n1105 GND 0.14fF
C1624 VDD.n1106 GND 0.17fF
C1625 VDD.n1107 GND 0.01fF
C1626 VDD.n1108 GND 0.02fF
C1627 VDD.n1109 GND 0.02fF
C1628 VDD.n1110 GND 0.11fF
C1629 VDD.n1111 GND 0.02fF
C1630 VDD.n1112 GND 0.14fF
C1631 VDD.n1113 GND 0.16fF
C1632 VDD.n1114 GND 0.01fF
C1633 VDD.n1115 GND 0.02fF
C1634 VDD.n1116 GND 0.02fF
C1635 VDD.n1117 GND 0.18fF
C1636 VDD.n1118 GND 0.15fF
C1637 VDD.n1119 GND 0.01fF
C1638 VDD.n1120 GND 0.02fF
C1639 VDD.n1121 GND 0.03fF
C1640 VDD.n1122 GND 0.18fF
C1641 VDD.n1123 GND 0.15fF
C1642 VDD.n1124 GND 0.01fF
C1643 VDD.n1125 GND 0.02fF
C1644 VDD.n1126 GND 0.03fF
C1645 VDD.n1127 GND 0.14fF
C1646 VDD.n1128 GND 0.16fF
C1647 VDD.n1129 GND 0.01fF
C1648 VDD.n1130 GND 0.11fF
C1649 VDD.n1131 GND 0.02fF
C1650 VDD.n1132 GND 0.02fF
C1651 VDD.n1133 GND 0.02fF
C1652 VDD.n1134 GND 0.14fF
C1653 VDD.n1135 GND 0.17fF
C1654 VDD.n1136 GND 0.01fF
C1655 VDD.n1137 GND 0.02fF
C1656 VDD.n1138 GND 0.02fF
C1657 VDD.n1139 GND 0.22fF
C1658 VDD.n1140 GND 0.01fF
C1659 VDD.n1141 GND 0.07fF
C1660 VDD.n1142 GND 0.02fF
C1661 VDD.n1143 GND 0.28fF
C1662 VDD.n1144 GND 0.01fF
C1663 VDD.n1145 GND 0.02fF
C1664 VDD.n1146 GND 0.02fF
C1665 VDD.n1147 GND 0.28fF
C1666 VDD.n1148 GND 0.01fF
C1667 VDD.n1149 GND 0.02fF
C1668 VDD.n1150 GND 0.03fF
C1669 VDD.n1151 GND 0.02fF
C1670 VDD.n1152 GND 0.02fF
C1671 VDD.n1153 GND 0.02fF
C1672 VDD.n1154 GND 0.26fF
C1673 VDD.n1155 GND 0.04fF
C1674 VDD.n1156 GND 0.03fF
C1675 VDD.n1157 GND 0.02fF
C1676 VDD.n1158 GND 0.02fF
C1677 VDD.n1159 GND 0.02fF
C1678 VDD.n1160 GND 0.03fF
C1679 VDD.n1161 GND 0.02fF
C1680 VDD.n1163 GND 0.02fF
C1681 VDD.n1164 GND 0.02fF
C1682 VDD.n1165 GND 0.02fF
C1683 VDD.n1167 GND 0.28fF
C1684 VDD.n1169 GND 0.02fF
C1685 VDD.n1170 GND 0.02fF
C1686 VDD.n1171 GND 0.03fF
C1687 VDD.n1172 GND 0.02fF
C1688 VDD.n1173 GND 0.28fF
C1689 VDD.n1174 GND 0.01fF
C1690 VDD.n1175 GND 0.02fF
C1691 VDD.n1176 GND 0.03fF
C1692 VDD.n1177 GND 0.06fF
C1693 VDD.n1178 GND 0.25fF
C1694 VDD.n1179 GND 0.01fF
C1695 VDD.n1180 GND 0.01fF
C1696 VDD.n1181 GND 0.02fF
C1697 VDD.n1182 GND 0.14fF
C1698 VDD.n1183 GND 0.16fF
C1699 VDD.n1184 GND 0.01fF
C1700 VDD.n1185 GND 0.02fF
C1701 VDD.n1186 GND 0.02fF
C1702 VDD.n1187 GND 0.17fF
C1703 VDD.n1188 GND 0.14fF
C1704 VDD.n1189 GND 0.01fF
C1705 VDD.n1190 GND 0.02fF
C1706 VDD.n1191 GND 0.03fF
C1707 VDD.n1192 GND 0.11fF
C1708 VDD.n1193 GND 0.03fF
C1709 VDD.n1194 GND 0.31fF
C1710 VDD.n1195 GND 0.01fF
C1711 VDD.n1196 GND 0.02fF
C1712 VDD.n1197 GND 0.03fF
C1713 VDD.n1198 GND 0.14fF
C1714 VDD.n1199 GND 0.17fF
C1715 VDD.n1200 GND 0.01fF
C1716 VDD.n1201 GND 0.02fF
C1717 VDD.n1202 GND 0.02fF
C1718 VDD.n1203 GND 0.06fF
C1719 VDD.n1204 GND 0.24fF
C1720 VDD.n1205 GND 0.01fF
C1721 VDD.n1206 GND 0.01fF
C1722 VDD.n1207 GND 0.02fF
C1723 VDD.n1208 GND 0.28fF
C1724 VDD.n1209 GND 0.01fF
C1725 VDD.n1210 GND 0.02fF
C1726 VDD.n1211 GND 0.03fF
C1727 VDD.n1212 GND 0.02fF
C1728 VDD.n1213 GND 0.02fF
C1729 VDD.n1214 GND 0.02fF
C1730 VDD.n1215 GND 0.26fF
C1731 VDD.n1216 GND 0.04fF
C1732 VDD.n1217 GND 0.03fF
C1733 VDD.n1218 GND 0.02fF
C1734 VDD.n1219 GND 0.02fF
C1735 VDD.n1220 GND 0.02fF
C1736 VDD.n1221 GND 0.03fF
C1737 VDD.n1222 GND 0.02fF
C1738 VDD.n1224 GND 0.02fF
C1739 VDD.n1225 GND 0.02fF
C1740 VDD.n1226 GND 0.02fF
C1741 VDD.n1228 GND 0.28fF
C1742 VDD.n1230 GND 0.02fF
C1743 VDD.n1231 GND 0.02fF
C1744 VDD.n1232 GND 0.03fF
C1745 VDD.n1233 GND 0.02fF
C1746 VDD.n1234 GND 0.28fF
C1747 VDD.n1235 GND 0.01fF
C1748 VDD.n1236 GND 0.02fF
C1749 VDD.n1237 GND 0.03fF
C1750 VDD.n1238 GND 0.28fF
C1751 VDD.n1239 GND 0.01fF
C1752 VDD.n1240 GND 0.02fF
C1753 VDD.n1241 GND 0.02fF
C1754 VDD.n1242 GND 0.06fF
C1755 VDD.n1243 GND 0.23fF
C1756 VDD.n1244 GND 0.01fF
C1757 VDD.n1245 GND 0.01fF
C1758 VDD.n1246 GND 0.02fF
C1759 VDD.n1247 GND 0.14fF
C1760 VDD.n1248 GND 0.17fF
C1761 VDD.n1249 GND 0.01fF
C1762 VDD.n1250 GND 0.02fF
C1763 VDD.n1251 GND 0.02fF
C1764 VDD.n1252 GND 0.11fF
C1765 VDD.n1253 GND 0.02fF
C1766 VDD.n1254 GND 0.14fF
C1767 VDD.n1255 GND 0.16fF
C1768 VDD.n1256 GND 0.01fF
C1769 VDD.n1257 GND 0.02fF
C1770 VDD.n1258 GND 0.02fF
C1771 VDD.n1259 GND 0.18fF
C1772 VDD.n1260 GND 0.15fF
C1773 VDD.n1261 GND 0.01fF
C1774 VDD.n1262 GND 0.02fF
C1775 VDD.n1263 GND 0.03fF
C1776 VDD.n1264 GND 0.18fF
C1777 VDD.n1265 GND 0.15fF
C1778 VDD.n1266 GND 0.01fF
C1779 VDD.n1267 GND 0.02fF
C1780 VDD.n1268 GND 0.03fF
C1781 VDD.n1269 GND 0.14fF
C1782 VDD.n1270 GND 0.16fF
C1783 VDD.n1271 GND 0.01fF
C1784 VDD.n1272 GND 0.11fF
C1785 VDD.n1273 GND 0.02fF
C1786 VDD.n1274 GND 0.02fF
C1787 VDD.n1275 GND 0.02fF
C1788 VDD.n1276 GND 0.14fF
C1789 VDD.n1277 GND 0.17fF
C1790 VDD.n1278 GND 0.01fF
C1791 VDD.n1279 GND 0.02fF
C1792 VDD.n1280 GND 0.02fF
C1793 VDD.n1281 GND 0.22fF
C1794 VDD.n1282 GND 0.01fF
C1795 VDD.n1283 GND 0.07fF
C1796 VDD.n1284 GND 0.02fF
C1797 VDD.n1285 GND 0.28fF
C1798 VDD.n1286 GND 0.01fF
C1799 VDD.n1287 GND 0.02fF
C1800 VDD.n1288 GND 0.02fF
C1801 VDD.n1289 GND 0.28fF
C1802 VDD.n1290 GND 0.01fF
C1803 VDD.n1291 GND 0.02fF
C1804 VDD.n1292 GND 0.03fF
C1805 VDD.n1293 GND 0.02fF
C1806 VDD.n1294 GND 0.02fF
C1807 VDD.n1295 GND 0.02fF
C1808 VDD.n1296 GND 0.31fF
C1809 VDD.n1297 GND 0.04fF
C1810 VDD.n1298 GND 0.03fF
C1811 VDD.n1299 GND 0.02fF
C1812 VDD.n1300 GND 0.02fF
C1813 VDD.n1301 GND 0.02fF
C1814 VDD.n1302 GND 0.03fF
C1815 VDD.n1303 GND 0.02fF
C1816 VDD.n1305 GND 0.02fF
C1817 VDD.n1306 GND 0.02fF
C1818 VDD.n1307 GND 0.02fF
C1819 VDD.n1309 GND 0.28fF
C1820 VDD.n1311 GND 0.02fF
C1821 VDD.n1312 GND 0.02fF
C1822 VDD.n1313 GND 0.03fF
C1823 VDD.n1314 GND 0.02fF
C1824 VDD.n1315 GND 0.28fF
C1825 VDD.n1316 GND 0.01fF
C1826 VDD.n1317 GND 0.02fF
C1827 VDD.n1318 GND 0.03fF
C1828 VDD.n1319 GND 0.28fF
C1829 VDD.n1320 GND 0.01fF
C1830 VDD.n1321 GND 0.02fF
C1831 VDD.n1322 GND 0.02fF
C1832 VDD.n1323 GND 0.06fF
C1833 VDD.n1324 GND 0.23fF
C1834 VDD.n1325 GND 0.01fF
C1835 VDD.n1326 GND 0.01fF
C1836 VDD.n1327 GND 0.02fF
C1837 VDD.n1328 GND 0.14fF
C1838 VDD.n1329 GND 0.17fF
C1839 VDD.n1330 GND 0.01fF
C1840 VDD.n1331 GND 0.02fF
C1841 VDD.n1332 GND 0.02fF
C1842 VDD.n1333 GND 0.11fF
C1843 VDD.n1334 GND 0.02fF
C1844 VDD.n1335 GND 0.14fF
C1845 VDD.n1336 GND 0.16fF
C1846 VDD.n1337 GND 0.01fF
C1847 VDD.n1338 GND 0.02fF
C1848 VDD.n1339 GND 0.02fF
C1849 VDD.n1340 GND 0.18fF
C1850 VDD.n1341 GND 0.15fF
C1851 VDD.n1342 GND 0.01fF
C1852 VDD.n1343 GND 0.02fF
C1853 VDD.n1344 GND 0.03fF
C1854 VDD.n1345 GND 0.18fF
C1855 VDD.n1346 GND 0.15fF
C1856 VDD.n1347 GND 0.01fF
C1857 VDD.n1348 GND 0.02fF
C1858 VDD.n1349 GND 0.03fF
C1859 VDD.n1350 GND 0.14fF
C1860 VDD.n1351 GND 0.16fF
C1861 VDD.n1352 GND 0.01fF
C1862 VDD.n1353 GND 0.11fF
C1863 VDD.n1354 GND 0.02fF
C1864 VDD.n1355 GND 0.02fF
C1865 VDD.n1356 GND 0.02fF
C1866 VDD.n1357 GND 0.14fF
C1867 VDD.n1358 GND 0.17fF
C1868 VDD.n1359 GND 0.01fF
C1869 VDD.n1360 GND 0.02fF
C1870 VDD.n1361 GND 0.02fF
C1871 VDD.n1362 GND 0.22fF
C1872 VDD.n1363 GND 0.01fF
C1873 VDD.n1364 GND 0.07fF
C1874 VDD.n1365 GND 0.02fF
C1875 VDD.n1366 GND 0.28fF
C1876 VDD.n1367 GND 0.01fF
C1877 VDD.n1368 GND 0.02fF
C1878 VDD.n1369 GND 0.02fF
C1879 VDD.n1370 GND 0.28fF
C1880 VDD.n1371 GND 0.01fF
C1881 VDD.n1372 GND 0.02fF
C1882 VDD.n1373 GND 0.03fF
C1883 VDD.n1374 GND 0.02fF
C1884 VDD.n1375 GND 0.02fF
C1885 VDD.n1376 GND 0.02fF
C1886 VDD.n1377 GND 0.26fF
C1887 VDD.n1378 GND 0.04fF
C1888 VDD.n1379 GND 0.03fF
C1889 VDD.n1380 GND 0.02fF
C1890 VDD.n1381 GND 0.02fF
C1891 VDD.n1382 GND 0.02fF
C1892 VDD.n1383 GND 0.03fF
C1893 VDD.n1384 GND 0.02fF
C1894 VDD.n1386 GND 0.02fF
C1895 VDD.n1387 GND 0.02fF
C1896 VDD.n1388 GND 0.02fF
C1897 VDD.n1390 GND 0.28fF
C1898 VDD.n1392 GND 0.02fF
C1899 VDD.n1393 GND 0.02fF
C1900 VDD.n1394 GND 0.03fF
C1901 VDD.n1395 GND 0.02fF
C1902 VDD.n1396 GND 0.28fF
C1903 VDD.n1397 GND 0.01fF
C1904 VDD.n1398 GND 0.02fF
C1905 VDD.n1399 GND 0.03fF
C1906 VDD.n1400 GND 0.06fF
C1907 VDD.n1401 GND 0.25fF
C1908 VDD.n1402 GND 0.01fF
C1909 VDD.n1403 GND 0.01fF
C1910 VDD.n1404 GND 0.02fF
C1911 VDD.n1405 GND 0.14fF
C1912 VDD.n1406 GND 0.16fF
C1913 VDD.n1407 GND 0.01fF
C1914 VDD.n1408 GND 0.02fF
C1915 VDD.n1409 GND 0.02fF
C1916 VDD.n1410 GND 0.17fF
C1917 VDD.n1411 GND 0.14fF
C1918 VDD.n1412 GND 0.01fF
C1919 VDD.n1413 GND 0.02fF
C1920 VDD.n1414 GND 0.03fF
C1921 VDD.n1415 GND 0.11fF
C1922 VDD.n1416 GND 0.03fF
C1923 VDD.n1417 GND 0.31fF
C1924 VDD.n1418 GND 0.01fF
C1925 VDD.n1419 GND 0.02fF
C1926 VDD.n1420 GND 0.03fF
C1927 VDD.n1421 GND 0.14fF
C1928 VDD.n1422 GND 0.17fF
C1929 VDD.n1423 GND 0.01fF
C1930 VDD.n1424 GND 0.02fF
C1931 VDD.n1425 GND 0.02fF
C1932 VDD.n1426 GND 0.06fF
C1933 VDD.n1427 GND 0.24fF
C1934 VDD.n1428 GND 0.01fF
C1935 VDD.n1429 GND 0.01fF
C1936 VDD.n1430 GND 0.02fF
C1937 VDD.n1431 GND 0.28fF
C1938 VDD.n1432 GND 0.01fF
C1939 VDD.n1433 GND 0.02fF
C1940 VDD.n1434 GND 0.03fF
C1941 VDD.n1435 GND 0.02fF
C1942 VDD.n1436 GND 0.02fF
C1943 VDD.n1437 GND 0.02fF
C1944 VDD.n1438 GND 0.22fF
C1945 VDD.n1439 GND 0.04fF
C1946 VDD.n1440 GND 0.03fF
C1947 VDD.n1441 GND 0.02fF
C1948 VDD.n1442 GND 0.02fF
C1949 VDD.n1443 GND 0.02fF
C1950 VDD.n1444 GND 0.03fF
C1951 VDD.n1445 GND 0.02fF
C1952 VDD.n1447 GND 0.02fF
C1953 VDD.n1448 GND 0.02fF
C1954 VDD.n1449 GND 0.02fF
C1955 VDD.n1451 GND 0.28fF
C1956 VDD.n1453 GND 0.02fF
C1957 VDD.n1454 GND 0.02fF
C1958 VDD.n1455 GND 0.03fF
C1959 VDD.n1456 GND 0.02fF
C1960 VDD.n1457 GND 0.28fF
C1961 VDD.n1458 GND 0.01fF
C1962 VDD.n1459 GND 0.02fF
C1963 VDD.n1460 GND 0.03fF
C1964 VDD.n1461 GND 0.06fF
C1965 VDD.n1462 GND 0.25fF
C1966 VDD.n1463 GND 0.01fF
C1967 VDD.n1464 GND 0.01fF
C1968 VDD.n1465 GND 0.02fF
C1969 a_8483_411.n0 GND 0.08fF
C1970 a_8483_411.n1 GND 1.05fF
C1971 a_8483_411.n2 GND 1.05fF
C1972 a_8483_411.n3 GND 1.23fF
C1973 a_8483_411.n4 GND 0.39fF
C1974 a_8483_411.n5 GND 0.60fF
C1975 a_8483_411.n6 GND 0.54fF
C1976 a_8483_411.n7 GND 1.45fF
C1977 a_8483_411.n8 GND 0.48fF
C1978 a_8483_411.n9 GND 1.04fF
C1979 a_8483_411.n10 GND 1.55fF
C1980 a_8483_411.n11 GND 0.66fF
C1981 a_8483_411.t15 GND 1.04fF
C1982 a_8483_411.n12 GND 0.79fF
C1983 a_8483_411.n13 GND 9.28fF
C1984 a_8483_411.n14 GND 0.88fF
C1985 a_8483_411.n15 GND 0.08fF
C1986 a_8483_411.n16 GND 0.59fF
C1987 a_8483_411.n17 GND 0.09fF
.ends
