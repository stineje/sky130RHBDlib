// File: INVX1.spi.pex
// Created: Tue Oct 15 15:49:25 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_INVX1\%GND ( 1 7 19 23 35 41 48 )
c26 ( 48 0 ) capacitor c=0.061451f //x=0.495 //y=0.37
c27 ( 41 0 ) capacitor c=0.234259f //x=1.6 //y=0
c28 ( 35 0 ) capacitor c=0.192978f //x=0.63 //y=0
c29 ( 26 0 ) capacitor c=0.00587411f //x=1.6 //y=0.45
c30 ( 23 0 ) capacitor c=0.00542558f //x=1.515 //y=0.535
c31 ( 22 0 ) capacitor c=0.00479856f //x=1.115 //y=0.45
c32 ( 19 0 ) capacitor c=0.00707849f //x=1.03 //y=0.535
c33 ( 14 0 ) capacitor c=0.00592191f //x=0.63 //y=0.45
c34 ( 7 0 ) capacitor c=0.11013f //x=1.48 //y=0
r35 (  40 41 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=1.48 //y=0 //x2=1.6 //y2=0
r36 (  38 40 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=1.115 //y=0 //x2=1.48 //y2=0
r37 (  37 38 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.115 //y2=0
r38 (  35 37 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=0.63 //y=0 //x2=0.74 //y2=0
r39 (  27 48 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.6 //y=0.62 //x2=1.6 //y2=0.535
r40 (  27 48 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.62 //x2=1.6 //y2=1.225
r41 (  26 48 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.6 //y=0.45 //x2=1.6 //y2=0.535
r42 (  25 41 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.6 //y=0.17 //x2=1.6 //y2=0
r43 (  25 26 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.6 //y=0.17 //x2=1.6 //y2=0.45
r44 (  24 48 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.2 //y=0.535 //x2=1.115 //y2=0.535
r45 (  23 48 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.6 //y2=0.535
r46 (  23 24 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.515 //y=0.535 //x2=1.2 //y2=0.535
r47 (  22 48 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.45 //x2=1.115 //y2=0.535
r48 (  21 38 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.115 //y=0.17 //x2=1.115 //y2=0
r49 (  21 22 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=1.115 //y=0.17 //x2=1.115 //y2=0.45
r50 (  20 48 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.715 //y=0.535 //x2=0.63 //y2=0.535
r51 (  19 48 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.03 //y=0.535 //x2=1.115 //y2=0.535
r52 (  19 20 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.03 //y=0.535 //x2=0.715 //y2=0.535
r53 (  15 48 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=0.63 //y=0.62 //x2=0.63 //y2=0.535
r54 (  15 48 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.62 //x2=0.63 //y2=1.225
r55 (  14 48 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=0.63 //y=0.45 //x2=0.63 //y2=0.535
r56 (  13 35 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=0.63 //y=0.17 //x2=0.63 //y2=0
r57 (  13 14 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=0.63 //y=0.17 //x2=0.63 //y2=0.45
r58 (  7 40 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=1.48 //y=0 //x2=1.48 //y2=0
r59 (  3 37 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=0.74 \
 //y=0 //x2=0.74 //y2=0
r60 (  1 7 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=1.11 //y=0 //x2=1.48 //y2=0
r61 (  1 3 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=1.11 //y=0 //x2=0.74 //y2=0
ends PM_INVX1\%GND

subckt PM_INVX1\%VDD ( 1 7 19 32 34 35 36 )
c23 ( 36 0 ) capacitor c=0.0451925f //x=1.41 //y=5.02
c24 ( 35 0 ) capacitor c=0.0427416f //x=0.54 //y=5.02
c25 ( 34 0 ) capacitor c=0.234796f //x=1.48 //y=7.4
c26 ( 32 0 ) capacitor c=0.233263f //x=0.74 //y=7.4
c27 ( 19 0 ) capacitor c=0.028745f //x=1.47 //y=7.4
c28 ( 7 0 ) capacitor c=0.110692f //x=1.48 //y=7.4
r29 (  21 34 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.555 //y=7.23 //x2=1.555 //y2=7.4
r30 (  21 36 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.555 //y=7.23 //x2=1.555 //y2=6.405
r31 (  20 32 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.76 //y=7.4 //x2=0.675 //y2=7.4
r32 (  19 34 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=1.555 //y2=7.4
r33 (  19 20 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.47 //y=7.4 //x2=0.76 //y2=7.4
r34 (  13 32 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=0.675 //y=7.23 //x2=0.675 //y2=7.4
r35 (  13 35 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.675 //y=7.23 //x2=0.675 //y2=6.405
r36 (  7 34 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=1.48 //y=7.4 //x2=1.48 //y2=7.4
r37 (  3 32 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=0.74 \
 //y=7.4 //x2=0.74 //y2=7.4
r38 (  1 7 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=1.11 //y=7.4 //x2=1.48 //y2=7.4
r39 (  1 3 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=1.11 //y=7.4 //x2=0.74 //y2=7.4
ends PM_INVX1\%VDD

subckt PM_INVX1\%A ( 1 2 3 4 5 6 7 9 21 22 23 24 25 26 27 31 32 33 35 41 42 44 )
c46 ( 44 0 ) capacitor c=0.0537799f //x=0.74 //y=2.085
c47 ( 42 0 ) capacitor c=0.0435629f //x=1.38 //y=1.255
c48 ( 41 0 ) capacitor c=0.0200386f //x=1.38 //y=0.91
c49 ( 35 0 ) capacitor c=0.0152946f //x=1.225 //y=1.41
c50 ( 33 0 ) capacitor c=0.0157804f //x=1.225 //y=0.755
c51 ( 32 0 ) capacitor c=0.0524167f //x=0.97 //y=4.79
c52 ( 31 0 ) capacitor c=0.0322983f //x=1.26 //y=4.79
c53 ( 27 0 ) capacitor c=0.0290017f //x=0.85 //y=1.92
c54 ( 26 0 ) capacitor c=0.0250027f //x=0.85 //y=1.565
c55 ( 25 0 ) capacitor c=0.0234316f //x=0.85 //y=1.255
c56 ( 24 0 ) capacitor c=0.0200596f //x=0.85 //y=0.91
c57 ( 23 0 ) capacitor c=0.154218f //x=1.335 //y=6.02
c58 ( 22 0 ) capacitor c=0.154243f //x=0.895 //y=6.02
c59 ( 9 0 ) capacitor c=0.115492f //x=0.74 //y=2.085
r60 (  44 45 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=0.74 //y=2.085 //x2=0.85 //y2=2.085
r61 (  42 51 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=1.255 //x2=1.34 //y2=1.41
r62 (  41 50 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.34 //y2=0.755
r63 (  41 42 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.38 //y=0.91 //x2=1.38 //y2=1.255
r64 (  36 49 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=1.41 //x2=0.89 //y2=1.41
r65 (  35 51 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=1.41 //x2=1.34 //y2=1.41
r66 (  34 48 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.005 //y=0.755 //x2=0.89 //y2=0.755
r67 (  33 50 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.34 //y2=0.755
r68 (  33 34 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.225 //y=0.755 //x2=1.005 //y2=0.755
r69 (  31 38 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=1.335 //y2=4.865
r70 (  31 32 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.26 //y=4.79 //x2=0.97 //y2=4.79
r71 (  28 32 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.97 //y2=4.79
r72 (  28 47 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=0.895 //y=4.865 //x2=0.74 //y2=4.7
r73 (  27 45 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.92 //x2=0.85 //y2=2.085
r74 (  26 49 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.89 //y2=1.41
r75 (  26 27 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.565 //x2=0.85 //y2=1.92
r76 (  25 49 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=1.255 //x2=0.89 //y2=1.41
r77 (  24 48 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.89 //y2=0.755
r78 (  24 25 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.85 //y=0.91 //x2=0.85 //y2=1.255
r79 (  23 38 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.335 //y=6.02 //x2=1.335 //y2=4.865
r80 (  22 28 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=0.895 //y=6.02 //x2=0.895 //y2=4.865
r81 (  21 35 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.225 //y2=1.41
r82 (  21 36 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.115 //y=1.41 //x2=1.005 //y2=1.41
r83 (  19 47 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=4.7 //x2=0.74 //y2=4.7
r84 (  9 44 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.74 //y=2.085 //x2=0.74 //y2=2.085
r85 (  7 19 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li //thickness=0.1 \
 //x=0.74 //y=4.44 //x2=0.74 //y2=4.7
r86 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=4.07 //x2=0.74 //y2=4.44
r87 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=3.7 //x2=0.74 //y2=4.07
r88 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=3.33 //x2=0.74 //y2=3.7
r89 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.96 //x2=0.74 //y2=3.33
r90 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.59 //x2=0.74 //y2=2.96
r91 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.22 //x2=0.74 //y2=2.59
r92 (  1 9 ) resistor r=9.24064 //w=0.187 //l=0.135 //layer=li //thickness=0.1 \
 //x=0.74 //y=2.22 //x2=0.74 //y2=2.085
ends PM_INVX1\%A

subckt PM_INVX1\%Y ( 1 2 3 4 5 6 7 18 19 20 21 31 33 )
c39 ( 33 0 ) capacitor c=0.028734f //x=0.97 //y=5.02
c40 ( 31 0 ) capacitor c=0.0173218f //x=0.925 //y=0.91
c41 ( 21 0 ) capacitor c=0.00575887f //x=1.2 //y=4.58
c42 ( 20 0 ) capacitor c=0.0146395f //x=1.395 //y=4.58
c43 ( 19 0 ) capacitor c=0.00636159f //x=1.195 //y=2.08
c44 ( 18 0 ) capacitor c=0.0141837f //x=1.395 //y=2.08
c45 ( 1 0 ) capacitor c=0.10647f //x=1.48 //y=2.22
r46 (  20 23 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.48 //y2=4.495
r47 (  20 21 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=1.395 //y=4.58 //x2=1.2 //y2=4.58
r48 (  18 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.395 //y=2.08 //x2=1.48 //y2=2.165
r49 (  18 19 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=1.395 //y=2.08 //x2=1.195 //y2=2.08
r50 (  12 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.2 //y2=4.58
r51 (  12 33 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=1.115 //y=4.665 //x2=1.115 //y2=5.725
r52 (  8 19 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.11 //y=1.995 //x2=1.195 //y2=2.08
r53 (  8 31 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=1.11 //y=1.995 //x2=1.11 //y2=1.005
r54 (  7 23 ) resistor r=3.76471 //w=0.187 //l=0.055 //layer=li \
 //thickness=0.1 //x=1.48 //y=4.44 //x2=1.48 //y2=4.495
r55 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.48 //y=4.07 //x2=1.48 //y2=4.44
r56 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.48 //y=3.7 //x2=1.48 //y2=4.07
r57 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.48 //y=3.33 //x2=1.48 //y2=3.7
r58 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.48 //y=2.96 //x2=1.48 //y2=3.33
r59 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.48 //y=2.59 //x2=1.48 //y2=2.96
r60 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.48 //y=2.22 //x2=1.48 //y2=2.59
r61 (  1 22 ) resistor r=3.76471 //w=0.187 //l=0.055 //layer=li \
 //thickness=0.1 //x=1.48 //y=2.22 //x2=1.48 //y2=2.165
ends PM_INVX1\%Y

