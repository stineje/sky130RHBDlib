* SPICE3 file created from OR2X1.ext - technology: sky130A

.subckt OR2X1 Y A B VPB VNB
M1000 a_198_181.t2 a_343_383# a_131_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_851_182.t1 a_198_181.t4 VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_131_1005.t2 a_164_908# VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t0 a_198_181.t5 a_851_182.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_131_1005.t0 a_343_383# a_198_181.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPB.t2 a_164_908# a_131_1005.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 a_343_383# VPB 0.07fF
C1 a_343_383# a_164_908# 0.26fF
C2 VPB a_164_908# 0.08fF
R0 a_131_1005.t0 a_131_1005.n0 101.663
R1 a_131_1005.n0 a_131_1005.t3 101.661
R2 a_131_1005.n0 a_131_1005.t1 14.294
R3 a_131_1005.n0 a_131_1005.t2 14.282
R4 a_198_181.n2 a_198_181.t5 512.525
R5 a_198_181.n2 a_198_181.t4 371.139
R6 a_198_181.n3 a_198_181.t6 220.263
R7 a_198_181.n4 a_198_181.n1 175.383
R8 a_198_181.n3 a_198_181.n2 158.3
R9 a_198_181.n4 a_198_181.n3 153.043
R10 a_198_181.n9 a_198_181.n4 145.681
R11 a_198_181.n9 a_198_181.n8 118.016
R12 a_198_181.n12 a_198_181.n0 55.263
R13 a_198_181.n11 a_198_181.n9 48.405
R14 a_198_181.n8 a_198_181.n7 30
R15 a_198_181.n11 a_198_181.n10 30
R16 a_198_181.n12 a_198_181.n11 25.263
R17 a_198_181.n6 a_198_181.n5 24.383
R18 a_198_181.n8 a_198_181.n6 23.684
R19 a_198_181.n1 a_198_181.t1 14.282
R20 a_198_181.n1 a_198_181.t2 14.282
R21 VPB VPB.n121 126.832
R22 VPB.n104 VPB.n102 94.117
R23 VPB.n106 VPB.n105 76
R24 VPB.n114 VPB.n113 76
R25 VPB.n75 VPB.n74 68.979
R26 VPB.n68 VPB.n67 64.528
R27 VPB.n27 VPB.n26 61.764
R28 VPB.n78 VPB.t1 55.106
R29 VPB.n66 VPB.t0 55.106
R30 VPB.n85 VPB.n84 44.502
R31 VPB.n88 VPB.n83 41.183
R32 VPB.n118 VPB.n114 20.452
R33 VPB.n65 VPB.n62 20.452
R34 VPB.n83 VPB.t3 14.282
R35 VPB.n83 VPB.t2 14.282
R36 VPB.n65 VPB.n64 13.653
R37 VPB.n64 VPB.n63 13.653
R38 VPB.n70 VPB.n69 13.653
R39 VPB.n69 VPB.n68 13.653
R40 VPB.n73 VPB.n72 13.653
R41 VPB.n72 VPB.n71 13.653
R42 VPB.n77 VPB.n76 13.653
R43 VPB.n76 VPB.n75 13.653
R44 VPB.n81 VPB.n80 13.653
R45 VPB.n80 VPB.n79 13.653
R46 VPB.n105 VPB.n104 13.653
R47 VPB.n104 VPB.n103 13.653
R48 VPB.n101 VPB.n100 13.653
R49 VPB.n100 VPB.n99 13.653
R50 VPB.n98 VPB.n97 13.653
R51 VPB.n97 VPB.n96 13.653
R52 VPB.n95 VPB.n94 13.653
R53 VPB.n94 VPB.n93 13.653
R54 VPB.n92 VPB.n91 13.653
R55 VPB.n91 VPB.n90 13.653
R56 VPB.n87 VPB.n86 13.653
R57 VPB.n86 VPB.n85 13.653
R58 VPB.n16 VPB.n15 13.653
R59 VPB.n15 VPB.n14 13.653
R60 VPB.n114 VPB.n0 13.653
R61 VPB VPB.n0 13.653
R62 VPB.n90 VPB.n89 13.35
R63 VPB.n118 VPB.n117 13.276
R64 VPB.n117 VPB.n115 13.276
R65 VPB.n41 VPB.n23 13.276
R66 VPB.n23 VPB.n21 13.276
R67 VPB.n73 VPB.n70 13.276
R68 VPB.n77 VPB.n73 13.276
R69 VPB.n82 VPB.n81 13.276
R70 VPB.n105 VPB.n82 13.276
R71 VPB.n105 VPB.n101 13.276
R72 VPB.n101 VPB.n98 13.276
R73 VPB.n98 VPB.n95 13.276
R74 VPB.n95 VPB.n92 13.276
R75 VPB.n87 VPB.n16 13.276
R76 VPB.n114 VPB.n16 13.276
R77 VPB.n62 VPB.n44 13.276
R78 VPB.n44 VPB.n42 13.276
R79 VPB.n49 VPB.n47 12.796
R80 VPB.n49 VPB.n48 12.564
R81 VPB.n55 VPB.n54 12.198
R82 VPB.n57 VPB.n56 12.198
R83 VPB.n55 VPB.n52 12.198
R84 VPB.n81 VPB.n78 10.944
R85 VPB.n66 VPB.n65 10.585
R86 VPB.n92 VPB.n88 8.97
R87 VPB.n62 VPB.n61 7.5
R88 VPB.n47 VPB.n46 7.5
R89 VPB.n54 VPB.n53 7.5
R90 VPB.n52 VPB.n51 7.5
R91 VPB.n44 VPB.n43 7.5
R92 VPB.n59 VPB.n45 7.5
R93 VPB.n23 VPB.n22 7.5
R94 VPB.n36 VPB.n35 7.5
R95 VPB.n30 VPB.n29 7.5
R96 VPB.n32 VPB.n31 7.5
R97 VPB.n25 VPB.n24 7.5
R98 VPB.n41 VPB.n40 7.5
R99 VPB.n117 VPB.n116 7.5
R100 VPB.n12 VPB.n11 7.5
R101 VPB.n6 VPB.n5 7.5
R102 VPB.n8 VPB.n7 7.5
R103 VPB.n2 VPB.n1 7.5
R104 VPB.n119 VPB.n118 7.5
R105 VPB.n82 VPB.n41 7.176
R106 VPB.n37 VPB.n34 6.729
R107 VPB.n33 VPB.n30 6.729
R108 VPB.n28 VPB.n25 6.729
R109 VPB.n13 VPB.n10 6.729
R110 VPB.n9 VPB.n6 6.729
R111 VPB.n4 VPB.n2 6.729
R112 VPB.n28 VPB.n27 6.728
R113 VPB.n33 VPB.n32 6.728
R114 VPB.n37 VPB.n36 6.728
R115 VPB.n40 VPB.n39 6.728
R116 VPB.n4 VPB.n3 6.728
R117 VPB.n9 VPB.n8 6.728
R118 VPB.n13 VPB.n12 6.728
R119 VPB.n120 VPB.n119 6.728
R120 VPB.n61 VPB.n60 6.398
R121 VPB.n88 VPB.n87 4.305
R122 VPB.n70 VPB.n66 2.691
R123 VPB.n78 VPB.n77 2.332
R124 VPB.n59 VPB.n50 1.402
R125 VPB.n59 VPB.n55 1.402
R126 VPB.n59 VPB.n57 1.402
R127 VPB.n59 VPB.n58 1.402
R128 VPB.n60 VPB.n59 0.735
R129 VPB.n59 VPB.n49 0.735
R130 VPB.n38 VPB.n37 0.387
R131 VPB.n38 VPB.n33 0.387
R132 VPB.n38 VPB.n28 0.387
R133 VPB.n39 VPB.n38 0.387
R134 VPB.n121 VPB.n13 0.387
R135 VPB.n121 VPB.n9 0.387
R136 VPB.n121 VPB.n4 0.387
R137 VPB.n121 VPB.n120 0.387
R138 VPB.n106 VPB.n20 0.272
R139 VPB.n113 VPB 0.198
R140 VPB.n18 VPB.n17 0.136
R141 VPB.n19 VPB.n18 0.136
R142 VPB.n20 VPB.n19 0.136
R143 VPB.n108 VPB.n107 0.136
R144 VPB.n109 VPB.n108 0.136
R145 VPB.n110 VPB.n109 0.136
R146 VPB.n111 VPB.n110 0.136
R147 VPB.n112 VPB.n111 0.136
R148 VPB.n113 VPB.n112 0.136
R149 VPB VPB.n106 0.068
R150 VPB.n107 VPB 0.068
R151 a_851_182.n3 a_851_182.n1 355.848
R152 a_851_182.n3 a_851_182.n2 30
R153 a_851_182.n4 a_851_182.n0 24.383
R154 a_851_182.n4 a_851_182.n3 23.684
R155 a_851_182.n1 a_851_182.t0 14.282
R156 a_851_182.n1 a_851_182.t1 14.282
R157 VNB VNB.n128 300.778
R158 VNB.n22 VNB.n21 199.897
R159 VNB.n105 VNB.n103 154.509
R160 VNB.n115 VNB.n114 76
R161 VNB.n107 VNB.n106 76
R162 VNB.n85 VNB.n84 62.533
R163 VNB.n63 VNB.n62 49.896
R164 VNB.n97 VNB.n96 36.267
R165 VNB.n38 VNB.n37 35.01
R166 VNB.t1 VNB.n30 32.601
R167 VNB.n56 VNB.n53 20.452
R168 VNB.n116 VNB.n115 20.452
R169 VNB.n57 VNB.n38 20.094
R170 VNB.n61 VNB.n35 20.094
R171 VNB.n68 VNB.n33 20.094
R172 VNB.n87 VNB.n80 19.735
R173 VNB.n91 VNB.n79 19.735
R174 VNB.n95 VNB.n76 19.735
R175 VNB.n102 VNB.n75 19.735
R176 VNB.n7 VNB.n6 19.735
R177 VNB.n38 VNB.n36 19.017
R178 VNB.n32 VNB.t1 17.353
R179 VNB.n5 VNB.t2 17.353
R180 VNB.n78 VNB.t0 13.654
R181 VNB.n60 VNB.n59 13.653
R182 VNB.n59 VNB.n58 13.653
R183 VNB.n64 VNB.n63 13.653
R184 VNB.n67 VNB.n66 13.653
R185 VNB.n66 VNB.n65 13.653
R186 VNB.n71 VNB.n70 13.653
R187 VNB.n70 VNB.n69 13.653
R188 VNB.n106 VNB.n105 13.653
R189 VNB.n105 VNB.n104 13.653
R190 VNB.n101 VNB.n100 13.653
R191 VNB.n100 VNB.n99 13.653
R192 VNB.n98 VNB.n97 13.653
R193 VNB.n94 VNB.n93 13.653
R194 VNB.n93 VNB.n92 13.653
R195 VNB.n90 VNB.n89 13.653
R196 VNB.n89 VNB.n88 13.653
R197 VNB.n86 VNB.n85 13.653
R198 VNB.n83 VNB.n82 13.653
R199 VNB.n82 VNB.n81 13.653
R200 VNB.n115 VNB.n0 13.653
R201 VNB VNB.n0 13.653
R202 VNB.n56 VNB.n55 13.653
R203 VNB.n55 VNB.n54 13.653
R204 VNB.n123 VNB.n120 13.577
R205 VNB.n41 VNB.n39 13.276
R206 VNB.n53 VNB.n41 13.276
R207 VNB.n14 VNB.n12 13.276
R208 VNB.n27 VNB.n14 13.276
R209 VNB.n67 VNB.n64 13.276
R210 VNB.n72 VNB.n71 13.276
R211 VNB.n106 VNB.n72 13.276
R212 VNB.n101 VNB.n98 13.276
R213 VNB.n86 VNB.n83 13.276
R214 VNB.n3 VNB.n1 13.276
R215 VNB.n116 VNB.n3 13.276
R216 VNB.n61 VNB.n60 13.097
R217 VNB.n33 VNB.n32 12.837
R218 VNB.n6 VNB.n5 12.837
R219 VNB.n106 VNB.n102 11.661
R220 VNB.n115 VNB.n7 11.661
R221 VNB.n75 VNB.n74 11.605
R222 VNB.n95 VNB.n94 10.764
R223 VNB.n90 VNB.n87 10.764
R224 VNB.n74 VNB.n73 9.809
R225 VNB.n71 VNB.n68 9.329
R226 VNB.n57 VNB.n56 8.97
R227 VNB.n32 VNB.n31 7.566
R228 VNB.n5 VNB.n4 7.566
R229 VNB.n125 VNB.n124 7.5
R230 VNB.n20 VNB.n19 7.5
R231 VNB.n16 VNB.n15 7.5
R232 VNB.n14 VNB.n13 7.5
R233 VNB.n27 VNB.n26 7.5
R234 VNB.n117 VNB.n116 7.5
R235 VNB.n3 VNB.n2 7.5
R236 VNB.n122 VNB.n121 7.5
R237 VNB.n47 VNB.n46 7.5
R238 VNB.n43 VNB.n42 7.5
R239 VNB.n41 VNB.n40 7.5
R240 VNB.n53 VNB.n52 7.5
R241 VNB.n72 VNB.n27 7.176
R242 VNB.t0 VNB.n77 7.04
R243 VNB.n127 VNB.n125 7.011
R244 VNB.n23 VNB.n20 7.011
R245 VNB.n18 VNB.n16 7.011
R246 VNB.n49 VNB.n47 7.011
R247 VNB.n45 VNB.n43 7.011
R248 VNB.n26 VNB.n25 7.01
R249 VNB.n18 VNB.n17 7.01
R250 VNB.n23 VNB.n22 7.01
R251 VNB.n52 VNB.n51 7.01
R252 VNB.n45 VNB.n44 7.01
R253 VNB.n49 VNB.n48 7.01
R254 VNB.n127 VNB.n126 7.01
R255 VNB.n123 VNB.n122 6.788
R256 VNB.n118 VNB.n117 6.788
R257 VNB.n94 VNB.n91 6.638
R258 VNB.n91 VNB.n90 6.638
R259 VNB.n79 VNB.n78 5.774
R260 VNB.n29 VNB.n28 4.551
R261 VNB.n60 VNB.n57 4.305
R262 VNB.n68 VNB.n67 3.947
R263 VNB.n98 VNB.n95 2.511
R264 VNB.n87 VNB.n86 2.511
R265 VNB.t1 VNB.n29 2.238
R266 VNB.n102 VNB.n101 1.614
R267 VNB.n83 VNB.n7 1.614
R268 VNB.n128 VNB.n119 0.921
R269 VNB.n128 VNB.n123 0.476
R270 VNB.n128 VNB.n118 0.475
R271 VNB.n35 VNB.n34 0.358
R272 VNB.n107 VNB.n11 0.272
R273 VNB.n24 VNB.n18 0.246
R274 VNB.n25 VNB.n24 0.246
R275 VNB.n24 VNB.n23 0.246
R276 VNB.n50 VNB.n45 0.246
R277 VNB.n51 VNB.n50 0.246
R278 VNB.n50 VNB.n49 0.246
R279 VNB.n128 VNB.n127 0.246
R280 VNB.n114 VNB 0.198
R281 VNB.n64 VNB.n61 0.179
R282 VNB.n9 VNB.n8 0.136
R283 VNB.n10 VNB.n9 0.136
R284 VNB.n11 VNB.n10 0.136
R285 VNB.n109 VNB.n108 0.136
R286 VNB.n110 VNB.n109 0.136
R287 VNB.n111 VNB.n110 0.136
R288 VNB.n112 VNB.n111 0.136
R289 VNB.n113 VNB.n112 0.136
R290 VNB.n114 VNB.n113 0.136
R291 VNB VNB.n107 0.068
R292 VNB.n108 VNB 0.068
C3 VPB VNB 5.42fF
C4 a_851_182.n0 VNB 0.04fF
C5 a_851_182.n1 VNB 1.02fF
C6 a_851_182.n2 VNB 0.04fF
C7 a_851_182.n3 VNB 0.50fF
C8 a_851_182.n4 VNB 0.06fF
C9 VPB.n0 VNB 0.03fF
C10 VPB.n1 VNB 0.03fF
C11 VPB.n2 VNB 0.02fF
C12 VPB.n3 VNB 0.13fF
C13 VPB.n5 VNB 0.02fF
C14 VPB.n6 VNB 0.02fF
C15 VPB.n7 VNB 0.02fF
C16 VPB.n8 VNB 0.02fF
C17 VPB.n10 VNB 0.02fF
C18 VPB.n11 VNB 0.02fF
C19 VPB.n12 VNB 0.02fF
C20 VPB.n14 VNB 0.22fF
C21 VPB.n15 VNB 0.02fF
C22 VPB.n16 VNB 0.02fF
C23 VPB.n17 VNB 0.07fF
C24 VPB.n18 VNB 0.02fF
C25 VPB.n19 VNB 0.02fF
C26 VPB.n20 VNB 0.03fF
C27 VPB.n21 VNB 0.02fF
C28 VPB.n22 VNB 0.02fF
C29 VPB.n23 VNB 0.02fF
C30 VPB.n24 VNB 0.03fF
C31 VPB.n25 VNB 0.02fF
C32 VPB.n26 VNB 0.16fF
C33 VPB.n27 VNB 0.04fF
C34 VPB.n29 VNB 0.02fF
C35 VPB.n30 VNB 0.02fF
C36 VPB.n31 VNB 0.02fF
C37 VPB.n32 VNB 0.02fF
C38 VPB.n34 VNB 0.02fF
C39 VPB.n35 VNB 0.02fF
C40 VPB.n36 VNB 0.02fF
C41 VPB.n38 VNB 0.26fF
C42 VPB.n40 VNB 0.02fF
C43 VPB.n41 VNB 0.02fF
C44 VPB.n42 VNB 0.02fF
C45 VPB.n43 VNB 0.02fF
C46 VPB.n44 VNB 0.02fF
C47 VPB.n45 VNB 0.10fF
C48 VPB.n46 VNB 0.03fF
C49 VPB.n47 VNB 0.02fF
C50 VPB.n48 VNB 0.04fF
C51 VPB.n49 VNB 0.01fF
C52 VPB.n51 VNB 0.02fF
C53 VPB.n52 VNB 0.02fF
C54 VPB.n53 VNB 0.02fF
C55 VPB.n54 VNB 0.02fF
C56 VPB.n56 VNB 0.02fF
C57 VPB.n59 VNB 0.43fF
C58 VPB.n61 VNB 0.03fF
C59 VPB.n62 VNB 0.04fF
C60 VPB.n63 VNB 0.26fF
C61 VPB.n64 VNB 0.03fF
C62 VPB.n65 VNB 0.03fF
C63 VPB.n66 VNB 0.05fF
C64 VPB.n67 VNB 0.13fF
C65 VPB.n68 VNB 0.18fF
C66 VPB.n69 VNB 0.02fF
C67 VPB.n70 VNB 0.01fF
C68 VPB.n71 VNB 0.15fF
C69 VPB.n72 VNB 0.02fF
C70 VPB.n73 VNB 0.02fF
C71 VPB.n74 VNB 0.13fF
C72 VPB.n75 VNB 0.18fF
C73 VPB.n76 VNB 0.02fF
C74 VPB.n77 VNB 0.01fF
C75 VPB.n78 VNB 0.05fF
C76 VPB.n79 VNB 0.26fF
C77 VPB.n80 VNB 0.01fF
C78 VPB.n81 VNB 0.02fF
C79 VPB.n82 VNB 0.03fF
C80 VPB.n83 VNB 0.09fF
C81 VPB.n84 VNB 0.13fF
C82 VPB.n85 VNB 0.15fF
C83 VPB.n86 VNB 0.02fF
C84 VPB.n87 VNB 0.02fF
C85 VPB.n88 VNB 0.02fF
C86 VPB.n89 VNB 0.13fF
C87 VPB.n90 VNB 0.14fF
C88 VPB.n91 VNB 0.02fF
C89 VPB.n92 VNB 0.02fF
C90 VPB.n93 VNB 0.26fF
C91 VPB.n94 VNB 0.02fF
C92 VPB.n95 VNB 0.02fF
C93 VPB.n96 VNB 0.26fF
C94 VPB.n97 VNB 0.02fF
C95 VPB.n98 VNB 0.02fF
C96 VPB.n99 VNB 0.26fF
C97 VPB.n100 VNB 0.02fF
C98 VPB.n101 VNB 0.02fF
C99 VPB.n102 VNB 0.03fF
C100 VPB.n103 VNB 0.26fF
C101 VPB.n104 VNB 0.01fF
C102 VPB.n105 VNB 0.02fF
C103 VPB.n106 VNB 0.03fF
C104 VPB.n107 VNB 0.02fF
C105 VPB.n108 VNB 0.02fF
C106 VPB.n109 VNB 0.02fF
C107 VPB.n110 VNB 0.02fF
C108 VPB.n111 VNB 0.02fF
C109 VPB.n112 VNB 0.02fF
C110 VPB.n113 VNB 0.03fF
C111 VPB.n114 VNB 0.03fF
C112 VPB.n115 VNB 0.02fF
C113 VPB.n116 VNB 0.02fF
C114 VPB.n117 VNB 0.02fF
C115 VPB.n118 VNB 0.04fF
C116 VPB.n119 VNB 0.03fF
C117 VPB.n121 VNB 0.40fF
C118 a_198_181.n0 VNB 0.04fF
C119 a_198_181.n1 VNB 0.56fF
C120 a_198_181.n2 VNB 0.29fF
C121 a_198_181.t6 VNB 0.43fF
C122 a_198_181.n3 VNB 0.48fF
C123 a_198_181.n4 VNB 0.43fF
C124 a_198_181.n5 VNB 0.03fF
C125 a_198_181.n6 VNB 0.04fF
C126 a_198_181.n7 VNB 0.03fF
C127 a_198_181.n8 VNB 0.15fF
C128 a_198_181.n9 VNB 0.31fF
C129 a_198_181.n10 VNB 0.03fF
C130 a_198_181.n11 VNB 0.08fF
C131 a_198_181.n12 VNB 0.04fF
C132 a_131_1005.n0 VNB 0.52fF
.ends
