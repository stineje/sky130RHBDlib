* SPICE3 file created from NAND2X1.ext - technology: sky130A

.subckt NAND2X1 Y A B VPB VNB
X0 VPB a_343_383# a_217_1004# VPB sky130_fd_pr__pfet_01v8 ad=1.68e+12p pd=1.368e+07u as=0p ps=0u w=2e+06u l=150000u M=2
X1 VNB a_168_157# a_112_73# VNB sky130_fd_pr__nfet_01v8 ad=1.791e+11p pd=1.57e+06u as=0p ps=0u w=3e+06u l=150000u
X2 a_217_1004# a_168_157# VPB VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u M=2
X3 a_217_1004# a_343_383# a_112_73# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
.ends
