magic
tech sky130A
magscale 1 2
timestamp 1652491038
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 3757 945 3791 979
rect 205 871 239 905
rect 1093 871 1127 905
rect 2943 871 2977 905
rect 3757 871 3791 905
rect 4127 871 4161 905
rect 4349 871 4383 905
rect 205 797 239 831
rect 3757 797 3791 831
rect 4127 797 4161 831
rect 4349 797 4383 831
rect 205 723 239 757
rect 1093 723 1127 757
rect 205 649 239 683
rect 1093 649 1127 683
rect 2055 649 2089 683
rect 2943 649 2977 683
rect 205 575 239 609
rect 1093 575 1127 609
rect 2055 575 2089 609
rect 2943 575 2977 609
rect 3757 575 3791 609
rect 4127 575 4161 609
rect 4349 575 4383 609
rect 205 501 239 535
rect 2055 501 2089 535
rect 2943 501 2977 535
rect 3757 501 3791 535
rect 4127 501 4161 535
rect 4349 501 4383 535
rect 205 427 239 461
rect 2055 427 2089 461
rect 4349 427 4383 461
<< metal1 >>
rect -34 1446 4918 1514
rect 3679 649 4683 683
rect 3827 575 4091 609
rect -34 -34 4918 34
use dffsnx1_pcell  dffsnx1_pcell_0 pcells
timestamp 1652396184
transform 1 0 0 0 1 0
box -87 -34 4971 1550
use li1_M1_contact  li1_M1_contact_2 pcells
timestamp 1648061256
transform -1 0 3626 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 3774 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 4144 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform 1 0 4736 0 1 666
box -53 -33 29 33
<< labels >>
rlabel locali 4127 575 4161 609 1 QN
port 1 nsew signal output
rlabel locali 4127 797 4161 831 1 QN
port 1 nsew signal output
rlabel locali 4127 871 4161 905 1 QN
port 1 nsew signal output
rlabel locali 4127 501 4161 535 1 QN
port 1 nsew signal output
rlabel locali 3757 501 3791 535 1 QN
port 1 nsew signal output
rlabel locali 3757 575 3791 609 1 QN
port 1 nsew signal output
rlabel locali 3757 797 3791 831 1 QN
port 1 nsew signal output
rlabel locali 3757 871 3791 905 1 QN
port 1 nsew signal output
rlabel locali 3757 945 3791 979 1 QN
port 1 nsew signal output
rlabel locali 205 723 239 757 1 D
port 2 nsew signal input
rlabel locali 205 649 239 683 1 D
port 2 nsew signal input
rlabel locali 205 575 239 609 1 D
port 2 nsew signal input
rlabel locali 205 501 239 535 1 D
port 2 nsew signal input
rlabel locali 205 427 239 461 1 D
port 2 nsew signal input
rlabel locali 205 797 239 831 1 D
port 2 nsew signal input
rlabel locali 205 871 239 905 1 D
port 2 nsew signal input
rlabel locali 1093 871 1127 905 1 CLK
port 3 nsew signal input
rlabel locali 1093 723 1127 757 1 CLK
port 3 nsew signal input
rlabel locali 1093 649 1127 683 1 CLK
port 3 nsew signal input
rlabel locali 1093 575 1127 609 1 CLK
port 3 nsew signal input
rlabel locali 2943 575 2977 609 1 CLK
port 3 nsew signal input
rlabel locali 2943 649 2977 683 1 CLK
port 3 nsew signal input
rlabel locali 2943 871 2977 905 1 CLK
port 3 nsew signal input
rlabel locali 2943 501 2977 535 1 CLK
port 3 nsew signal input
rlabel locali 2055 427 2089 461 1 SN
port 4 nsew signal input
rlabel locali 2055 501 2089 535 1 SN
port 4 nsew signal input
rlabel locali 2055 575 2089 609 1 SN
port 4 nsew signal input
rlabel locali 2055 649 2089 683 1 SN
port 4 nsew signal input
rlabel locali 4349 427 4383 461 1 SN
port 4 nsew signal input
rlabel locali 4349 501 4383 535 1 SN
port 4 nsew signal input
rlabel locali 4349 575 4383 609 1 SN
port 4 nsew signal input
rlabel locali 4349 797 4383 831 1 SN
port 4 nsew signal input
rlabel locali 4349 871 4383 905 1 SN
port 4 nsew signal input
rlabel metal1 -34 1446 4918 1514 1 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 -34 -34 4918 34 1 VGND
port 6 nsew ground bidirectional abutment
rlabel nwell 57 1463 91 1497 1 VPB
rlabel pwell 57 -17 91 17 1 VNB
<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 4884 1480
string LEFsymmetry X Y R90
<< end >>
