// File: nor2x1_pcell.spi.pex
// Created: Tue Oct 15 15:59:23 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_NOR2X1_PCELL\%noxref_1 ( 7 19 23 31 35 47 57 68 )
c37 ( 68 0 ) capacitor c=0.0747013f //x=0.56 //y=0.365
c38 ( 57 0 ) capacitor c=0.270467f //x=2.635 //y=0
c39 ( 47 0 ) capacitor c=0.202778f //x=0.695 //y=0
c40 ( 38 0 ) capacitor c=0.00609805f //x=2.635 //y=0.445
c41 ( 35 0 ) capacitor c=0.00510317f //x=2.55 //y=0.53
c42 ( 34 0 ) capacitor c=0.00468234f //x=2.15 //y=0.445
c43 ( 31 0 ) capacitor c=0.00556167f //x=2.065 //y=0.53
c44 ( 26 0 ) capacitor c=0.00468234f //x=1.665 //y=0.445
c45 ( 23 0 ) capacitor c=0.00556167f //x=1.58 //y=0.53
c46 ( 22 0 ) capacitor c=0.00468234f //x=1.18 //y=0.445
c47 ( 19 0 ) capacitor c=0.00709092f //x=1.095 //y=0.53
c48 ( 14 0 ) capacitor c=0.00609805f //x=0.695 //y=0.445
c49 ( 7 0 ) capacitor c=0.149169f //x=2.59 //y=0
r50 (  56 57 ) resistor r=1.61345 //w=0.357 //l=0.045 //layer=li \
 //thickness=0.1 //x=2.59 //y=0 //x2=2.635 //y2=0
r51 (  54 56 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=2.15 //y=0 //x2=2.59 //y2=0
r52 (  53 54 ) resistor r=10.7563 //w=0.357 //l=0.3 //layer=li //thickness=0.1 \
 //x=1.85 //y=0 //x2=2.15 //y2=0
r53 (  51 53 ) resistor r=6.63305 //w=0.357 //l=0.185 //layer=li \
 //thickness=0.1 //x=1.665 //y=0 //x2=1.85 //y2=0
r54 (  50 51 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.18 //y=0 //x2=1.665 //y2=0
r55 (  49 50 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.18 //y2=0
r56 (  47 49 ) resistor r=1.61345 //w=0.357 //l=0.045 //layer=li \
 //thickness=0.1 //x=0.695 //y=0 //x2=0.74 //y2=0
r57 (  39 68 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.635 //y=0.615 //x2=2.635 //y2=0.53
r58 (  39 68 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r59 (  38 68 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.635 //y=0.445 //x2=2.635 //y2=0.53
r60 (  37 57 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.635 //y=0.17 //x2=2.635 //y2=0
r61 (  37 38 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.17 //x2=2.635 //y2=0.445
r62 (  36 68 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.235 //y=0.53 //x2=2.15 //y2=0.53
r63 (  35 68 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.53
r64 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.235 //y2=0.53
r65 (  34 68 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.445 //x2=2.15 //y2=0.53
r66 (  33 54 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.15 //y=0.17 //x2=2.15 //y2=0
r67 (  33 34 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.17 //x2=2.15 //y2=0.445
r68 (  32 68 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=1.665 //y2=0.53
r69 (  31 68 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.065 //y=0.53 //x2=2.15 //y2=0.53
r70 (  31 32 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=2.065 //y=0.53 //x2=1.75 //y2=0.53
r71 (  27 68 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.53
r72 (  27 68 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r73 (  26 68 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.445 //x2=1.665 //y2=0.53
r74 (  25 51 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.17 //x2=1.665 //y2=0
r75 (  25 26 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.17 //x2=1.665 //y2=0.445
r76 (  24 68 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.265 //y=0.53 //x2=1.18 //y2=0.53
r77 (  23 68 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.58 //y=0.53 //x2=1.665 //y2=0.53
r78 (  23 24 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.58 //y=0.53 //x2=1.265 //y2=0.53
r79 (  22 68 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.445 //x2=1.18 //y2=0.53
r80 (  21 50 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r81 (  21 22 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.445
r82 (  20 68 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.78 //y=0.53 //x2=0.695 //y2=0.53
r83 (  19 68 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.095 //y=0.53 //x2=1.18 //y2=0.53
r84 (  19 20 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.095 //y=0.53 //x2=0.78 //y2=0.53
r85 (  15 68 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=0.695 //y=0.615 //x2=0.695 //y2=0.53
r86 (  15 68 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.615 //x2=0.695 //y2=1.22
r87 (  14 68 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=0.695 //y=0.445 //x2=0.695 //y2=0.53
r88 (  13 47 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=0.695 //y=0.17 //x2=0.695 //y2=0
r89 (  13 14 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.17 //x2=0.695 //y2=0.445
r90 (  7 56 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=2.59 //y=0 //x2=2.59 //y2=0
r91 (  5 53 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=1.85 \
 //y=0 //x2=1.85 //y2=0
r92 (  5 7 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.59 //y2=0
r93 (  2 49 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=0.74 \
 //y=0 //x2=0.74 //y2=0
r94 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
ends PM_NOR2X1_PCELL\%noxref_1

subckt PM_NOR2X1_PCELL\%noxref_2 ( 7 11 14 26 30 )
c36 ( 30 0 ) capacitor c=0.0256796f //x=1.085 //y=5.025
c37 ( 29 0 ) capacitor c=0.00591168f //x=1.23 //y=7.4
c38 ( 26 0 ) capacitor c=0.287106f //x=2.59 //y=7.4
c39 ( 14 0 ) capacitor c=0.210107f //x=0.74 //y=7.4
c40 ( 11 0 ) capacitor c=0.0465804f //x=1.145 //y=7.4
c41 ( 7 0 ) capacitor c=0.151267f //x=2.59 //y=7.4
r42 (  24 26 ) resistor r=26.5322 //w=0.357 //l=0.74 //layer=li \
 //thickness=0.1 //x=1.85 //y=7.4 //x2=2.59 //y2=7.4
r43 (  22 29 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.315 //y=7.4 //x2=1.23 //y2=7.4
r44 (  22 24 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=1.315 //y=7.4 //x2=1.85 //y2=7.4
r45 (  15 29 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.23 //y=7.23 //x2=1.23 //y2=7.4
r46 (  15 30 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=1.23 //y=7.23 //x2=1.23 //y2=6.74
r47 (  11 29 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.145 //y=7.4 //x2=1.23 //y2=7.4
r48 (  11 14 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=1.145 //y=7.4 //x2=0.74 //y2=7.4
r49 (  7 26 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=2.59 //y=7.4 //x2=2.59 //y2=7.4
r50 (  5 24 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=1.85 \
 //y=7.4 //x2=1.85 //y2=7.4
r51 (  5 7 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.59 //y2=7.4
r52 (  2 14 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=0.74 \
 //y=7.4 //x2=0.74 //y2=7.4
r53 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_NOR2X1_PCELL\%noxref_2

subckt PM_NOR2X1_PCELL\%noxref_3 ( 3 6 8 9 10 11 12 13 14 18 20 23 25 26 31 )
c65 ( 31 0 ) capacitor c=0.04214f //x=0.955 //y=4.705
c66 ( 26 0 ) capacitor c=0.0321911f //x=1.445 //y=1.25
c67 ( 25 0 ) capacitor c=0.0185201f //x=1.445 //y=0.905
c68 ( 23 0 ) capacitor c=0.0344254f //x=1.375 //y=4.795
c69 ( 20 0 ) capacitor c=0.0133656f //x=1.29 //y=1.405
c70 ( 18 0 ) capacitor c=0.0157804f //x=1.29 //y=0.75
c71 ( 14 0 ) capacitor c=0.0828832f //x=0.915 //y=1.915
c72 ( 13 0 ) capacitor c=0.022867f //x=0.915 //y=1.56
c73 ( 12 0 ) capacitor c=0.0234318f //x=0.915 //y=1.25
c74 ( 11 0 ) capacitor c=0.0192004f //x=0.915 //y=0.905
c75 ( 10 0 ) capacitor c=0.110795f //x=1.45 //y=6.025
c76 ( 9 0 ) capacitor c=0.153847f //x=1.01 //y=6.025
c77 ( 6 0 ) capacitor c=0.00995068f //x=0.955 //y=4.705
c78 ( 3 0 ) capacitor c=0.112895f //x=1.11 //y=2.08
r79 (  33 34 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=0.955 //y=4.795 //x2=0.955 //y2=4.87
r80 (  31 33 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=0.955 //y=4.705 //x2=0.955 //y2=4.795
r81 (  26 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.25 //x2=1.405 //y2=1.405
r82 (  25 39 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.905 //x2=1.405 //y2=0.75
r83 (  25 26 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.905 //x2=1.445 //y2=1.25
r84 (  24 33 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=1.09 //y=4.795 //x2=0.955 //y2=4.795
r85 (  23 27 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.375 //y=4.795 //x2=1.45 //y2=4.87
r86 (  23 24 ) resistor r=146.138 //w=0.094 //l=0.285 //layer=ply \
 //thickness=0.18 //x=1.375 //y=4.795 //x2=1.09 //y2=4.795
r87 (  21 38 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.405 //x2=0.955 //y2=1.405
r88 (  20 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.405 //x2=1.405 //y2=1.405
r89 (  19 37 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.75 //x2=0.955 //y2=0.75
r90 (  18 39 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.75 //x2=1.405 //y2=0.75
r91 (  18 19 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.75 //x2=1.07 //y2=0.75
r92 (  14 36 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r93 (  13 38 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.56 //x2=0.955 //y2=1.405
r94 (  13 14 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.56 //x2=0.915 //y2=1.915
r95 (  12 38 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.25 //x2=0.955 //y2=1.405
r96 (  11 37 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.905 //x2=0.955 //y2=0.75
r97 (  11 12 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.905 //x2=0.915 //y2=1.25
r98 (  10 27 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.025 //x2=1.45 //y2=4.87
r99 (  9 34 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.025 //x2=1.01 //y2=4.87
r100 (  8 20 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.405 //x2=1.29 //y2=1.405
r101 (  8 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.405 //x2=1.07 //y2=1.405
r102 (  6 31 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.955 //y=4.705 //x2=0.955 //y2=4.705
r103 (  6 7 ) resistor r=7.81102 //w=0.254 //l=0.155 //layer=li \
 //thickness=0.1 //x=0.955 //y=4.705 //x2=1.11 //y2=4.705
r104 (  3 36 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r105 (  1 7 ) resistor r=3.23951 //w=0.254 //l=0.165 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.54 //x2=1.11 //y2=4.705
r106 (  1 3 ) resistor r=168.385 //w=0.187 //l=2.46 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.54 //x2=1.11 //y2=2.08
ends PM_NOR2X1_PCELL\%noxref_3

subckt PM_NOR2X1_PCELL\%noxref_4 ( 1 3 7 8 9 10 11 12 17 19 21 27 28 30 31 34 )
c66 ( 34 0 ) capacitor c=0.0369822f //x=1.885 //y=4.705
c67 ( 31 0 ) capacitor c=0.0279572f //x=1.85 //y=1.915
c68 ( 30 0 ) capacitor c=0.0422144f //x=1.85 //y=2.08
c69 ( 28 0 ) capacitor c=0.0237734f //x=2.415 //y=1.255
c70 ( 27 0 ) capacitor c=0.0191782f //x=2.415 //y=0.905
c71 ( 21 0 ) capacitor c=0.0346941f //x=2.26 //y=1.405
c72 ( 19 0 ) capacitor c=0.0157803f //x=2.26 //y=0.75
c73 ( 17 0 ) capacitor c=0.0359964f //x=2.255 //y=4.795
c74 ( 12 0 ) capacitor c=0.0199921f //x=1.885 //y=1.56
c75 ( 11 0 ) capacitor c=0.0169608f //x=1.885 //y=1.255
c76 ( 10 0 ) capacitor c=0.0185462f //x=1.885 //y=0.905
c77 ( 9 0 ) capacitor c=0.15325f //x=2.33 //y=6.025
c78 ( 8 0 ) capacitor c=0.110232f //x=1.89 //y=6.025
c79 ( 3 0 ) capacitor c=0.0818408f //x=1.85 //y=2.08
c80 ( 1 0 ) capacitor c=0.00521267f //x=1.85 //y=4.54
r81 (  36 37 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.885 //y=4.795 //x2=1.885 //y2=4.87
r82 (  34 36 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.885 //y=4.705 //x2=1.885 //y2=4.795
r83 (  30 31 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r84 (  28 41 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.255 //x2=2.415 //y2=1.367
r85 (  27 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r86 (  27 28 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.255
r87 (  22 39 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r88 (  21 41 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.415 //y2=1.367
r89 (  20 38 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r90 (  19 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r91 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r92 (  18 36 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.02 //y=4.795 //x2=1.885 //y2=4.795
r93 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.795 //x2=2.33 //y2=4.87
r94 (  17 18 ) resistor r=120.5 //w=0.094 //l=0.235 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.795 //x2=2.02 //y2=4.795
r95 (  12 39 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r96 (  12 31 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r97 (  11 39 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.255 //x2=1.925 //y2=1.405
r98 (  10 38 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r99 (  10 11 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.255
r100 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.025 //x2=2.33 //y2=4.87
r101 (  8 37 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.025 //x2=1.89 //y2=4.87
r102 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r103 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r104 (  6 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.885 //y=4.705 //x2=1.885 //y2=4.705
r105 (  3 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r106 (  1 6 ) resistor r=11.332 //w=0.189 //l=0.173292 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.54 //x2=1.867 //y2=4.705
r107 (  1 3 ) resistor r=168.385 //w=0.187 //l=2.46 //layer=li //thickness=0.1 \
 //x=1.85 //y=4.54 //x2=1.85 //y2=2.08
ends PM_NOR2X1_PCELL\%noxref_4

subckt PM_NOR2X1_PCELL\%noxref_5 ( 5 6 17 18 19 22 24 25 28 )
c65 ( 28 0 ) capacitor c=0.0159573f //x=1.965 //y=5.025
c66 ( 25 0 ) capacitor c=0.00905936f //x=1.96 //y=0.905
c67 ( 24 0 ) capacitor c=0.007684f //x=0.99 //y=0.905
c68 ( 23 0 ) capacitor c=0.00710337f //x=2.15 //y=1.655
c69 ( 22 0 ) capacitor c=0.133888f //x=2.59 //y=5.125
c70 ( 19 0 ) capacitor c=0.0169019f //x=2.505 //y=1.655
c71 ( 18 0 ) capacitor c=0.00499395f //x=2.195 //y=5.21
c72 ( 17 0 ) capacitor c=0.0164583f //x=2.505 //y=5.21
c73 ( 6 0 ) capacitor c=0.00277607f //x=1.265 //y=1.655
c74 ( 5 0 ) capacitor c=0.0280953f //x=2.065 //y=1.655
r75 (  21 22 ) resistor r=231.701 //w=0.187 //l=3.385 //layer=li \
 //thickness=0.1 //x=2.59 //y=1.74 //x2=2.59 //y2=5.125
r76 (  20 23 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.235 //y=1.655 //x2=2.15 //y2=1.655
r77 (  19 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.59 //y2=1.74
r78 (  19 20 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.235 //y2=1.655
r79 (  17 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.21 //x2=2.59 //y2=5.125
r80 (  17 18 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.21 //x2=2.195 //y2=5.21
r81 (  13 23 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1.655
r82 (  13 25 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r83 (  7 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.295 //x2=2.195 //y2=5.21
r84 (  7 28 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.295 //x2=2.11 //y2=5.72
r85 (  5 23 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.065 //y=1.655 //x2=2.15 //y2=1.655
r86 (  5 6 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li //thickness=0.1 \
 //x=2.065 //y=1.655 //x2=1.265 //y2=1.655
r87 (  1 6 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.18 //y=1.57 //x2=1.265 //y2=1.655
r88 (  1 24 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=1.18 //y=1.57 //x2=1.18 //y2=1
ends PM_NOR2X1_PCELL\%noxref_5

subckt PM_NOR2X1_PCELL\%noxref_6 ( 7 8 15 16 23 24 25 )
c37 ( 25 0 ) capacitor c=0.0308836f //x=2.405 //y=5.025
c38 ( 24 0 ) capacitor c=0.0185379f //x=1.525 //y=5.025
c39 ( 23 0 ) capacitor c=0.0409962f //x=0.655 //y=5.025
c40 ( 16 0 ) capacitor c=0.00193672f //x=1.755 //y=6.91
c41 ( 15 0 ) capacitor c=0.01354f //x=2.465 //y=6.91
c42 ( 8 0 ) capacitor c=0.00844339f //x=0.875 //y=5.21
c43 ( 7 0 ) capacitor c=0.0252644f //x=1.585 //y=5.21
r44 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.55 //y=6.825 //x2=2.55 //y2=6.74
r45 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.465 //y=6.91 //x2=2.55 //y2=6.825
r46 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.465 //y=6.91 //x2=1.755 //y2=6.91
r47 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.67 //y=6.825 //x2=1.755 //y2=6.91
r48 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.67 //y=6.825 //x2=1.67 //y2=6.4
r49 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.67 //y=5.295 //x2=1.67 //y2=5.72
r50 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.585 //y=5.21 //x2=1.67 //y2=5.295
r51 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=1.585 //y=5.21 //x2=0.875 //y2=5.21
r52 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=0.79 //y=5.295 //x2=0.875 //y2=5.21
r53 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=0.79 //y=5.295 //x2=0.79 //y2=5.72
ends PM_NOR2X1_PCELL\%noxref_6

