// File: pmos2_1.spi.pex
// Created: Tue Oct 15 16:00:29 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_PMOS2_1\%noxref_4 ( 1 2 6 )
c5 ( 7 0 ) capacitor c=0.0190444f //x=0.87 //y=-2.225
c6 ( 6 0 ) capacitor c=0.0437142f //x=1.16 //y=-2.225
c7 ( 2 0 ) capacitor c=0.177708f //x=1.235 //y=-0.995
c8 ( 1 0 ) capacitor c=0.177708f //x=0.795 //y=-0.995
r9 (  6 8 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.16 //y=-2.225 //x2=1.235 //y2=-2.15
r10 (  6 7 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.16 //y=-2.225 //x2=0.87 //y2=-2.225
r11 (  3 7 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=0.795 //y=-2.15 //x2=0.87 //y2=-2.225
r12 (  2 8 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.235 //y=-0.995 //x2=1.235 //y2=-2.15
r13 (  1 3 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=0.795 //y=-0.995 //x2=0.795 //y2=-2.15
ends PM_PMOS2_1\%noxref_4

