// File: aoa4x1_pcell.spi.pex
// Created: Tue Oct 15 15:54:59 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_AOA4X1_PCELL\%noxref_1 ( 21 25 28 33 44 49 53 61 65 68 77 85 96 101 \
 105 118 138 140 147 154 155 156 157 )
c169 ( 157 0 ) capacitor c=0.0597349f //x=10.485 //y=0.37
c170 ( 156 0 ) capacitor c=0.0207703f //x=7.65 //y=0.865
c171 ( 155 0 ) capacitor c=0.0698863f //x=3.89 //y=0.365
c172 ( 154 0 ) capacitor c=0.0208404f //x=0.99 //y=0.865
c173 ( 147 0 ) capacitor c=0.233789f //x=11.59 //y=0
c174 ( 140 0 ) capacitor c=0.101261f //x=9.99 //y=0
c175 ( 139 0 ) capacitor c=0.00440095f //x=7.84 //y=0
c176 ( 138 0 ) capacitor c=0.10428f //x=6.66 //y=0
c177 ( 118 0 ) capacitor c=0.107062f //x=3.33 //y=0
c178 ( 117 0 ) capacitor c=0.00440095f //x=1.18 //y=0
c179 ( 108 0 ) capacitor c=0.00583665f //x=11.59 //y=0.45
c180 ( 105 0 ) capacitor c=0.00542558f //x=11.505 //y=0.535
c181 ( 104 0 ) capacitor c=0.00479856f //x=11.105 //y=0.45
c182 ( 101 0 ) capacitor c=0.00690112f //x=11.02 //y=0.535
c183 ( 96 0 ) capacitor c=0.00588377f //x=10.62 //y=0.45
c184 ( 93 0 ) capacitor c=0.0190475f //x=10.535 //y=0
c185 ( 85 0 ) capacitor c=0.0751168f //x=9.82 //y=0
c186 ( 77 0 ) capacitor c=0.0426751f //x=7.755 //y=0
c187 ( 74 0 ) capacitor c=0.0659312f //x=6.05 //y=0
c188 ( 73 0 ) capacitor c=0.0227441f //x=6.49 //y=0
c189 ( 68 0 ) capacitor c=0.00609805f //x=5.965 //y=0.445
c190 ( 65 0 ) capacitor c=0.00508073f //x=5.88 //y=0.53
c191 ( 64 0 ) capacitor c=0.00468234f //x=5.48 //y=0.445
c192 ( 61 0 ) capacitor c=0.00556167f //x=5.395 //y=0.53
c193 ( 56 0 ) capacitor c=0.00468234f //x=4.995 //y=0.445
c194 ( 53 0 ) capacitor c=0.00556167f //x=4.91 //y=0.53
c195 ( 52 0 ) capacitor c=0.00468234f //x=4.51 //y=0.445
c196 ( 49 0 ) capacitor c=0.00692577f //x=4.425 //y=0.53
c197 ( 44 0 ) capacitor c=0.00609805f //x=4.025 //y=0.445
c198 ( 41 0 ) capacitor c=0.0227441f //x=3.94 //y=0
c199 ( 33 0 ) capacitor c=0.0751168f //x=3.16 //y=0
c200 ( 28 0 ) capacitor c=0.179504f //x=0.74 //y=0
c201 ( 25 0 ) capacitor c=0.0426751f //x=1.095 //y=0
c202 ( 21 0 ) capacitor c=0.458606f //x=11.47 //y=0
r203 (  146 147 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=11.47 //y=0 //x2=11.59 //y2=0
r204 (  144 146 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=11.105 //y=0 //x2=11.47 //y2=0
r205 (  143 144 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=10.73 //y=0 //x2=11.105 //y2=0
r206 (  141 143 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=10.62 //y=0 //x2=10.73 //y2=0
r207 (  126 127 ) resistor r=14.8796 //w=0.357 //l=0.415 //layer=li \
 //thickness=0.1 //x=5.55 //y=0 //x2=5.965 //y2=0
r208 (  124 126 ) resistor r=2.5098 //w=0.357 //l=0.07 //layer=li \
 //thickness=0.1 //x=5.48 //y=0 //x2=5.55 //y2=0
r209 (  123 124 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.995 //y=0 //x2=5.48 //y2=0
r210 (  122 123 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.51 //y=0 //x2=4.995 //y2=0
r211 (  121 122 ) resistor r=2.5098 //w=0.357 //l=0.07 //layer=li \
 //thickness=0.1 //x=4.44 //y=0 //x2=4.51 //y2=0
r212 (  119 121 ) resistor r=14.8796 //w=0.357 //l=0.415 //layer=li \
 //thickness=0.1 //x=4.025 //y=0 //x2=4.44 //y2=0
r213 (  109 157 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.59 //y=0.62 //x2=11.59 //y2=0.535
r214 (  109 157 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=11.59 //y=0.62 //x2=11.59 //y2=1.225
r215 (  108 157 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.59 //y=0.45 //x2=11.59 //y2=0.535
r216 (  107 147 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.59 //y=0.17 //x2=11.59 //y2=0
r217 (  107 108 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=11.59 //y=0.17 //x2=11.59 //y2=0.45
r218 (  106 157 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.19 //y=0.535 //x2=11.105 //y2=0.535
r219 (  105 157 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.505 //y=0.535 //x2=11.59 //y2=0.535
r220 (  105 106 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=11.505 //y=0.535 //x2=11.19 //y2=0.535
r221 (  104 157 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.105 //y=0.45 //x2=11.105 //y2=0.535
r222 (  103 144 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.105 //y=0.17 //x2=11.105 //y2=0
r223 (  103 104 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=11.105 //y=0.17 //x2=11.105 //y2=0.45
r224 (  102 157 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.705 //y=0.535 //x2=10.62 //y2=0.535
r225 (  101 157 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.02 //y=0.535 //x2=11.105 //y2=0.535
r226 (  101 102 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=11.02 //y=0.535 //x2=10.705 //y2=0.535
r227 (  97 157 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.62 //y=0.62 //x2=10.62 //y2=0.535
r228 (  97 157 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=10.62 //y=0.62 //x2=10.62 //y2=1.225
r229 (  96 157 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.62 //y=0.45 //x2=10.62 //y2=0.535
r230 (  95 141 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.62 //y=0.17 //x2=10.62 //y2=0
r231 (  95 96 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=10.62 //y=0.17 //x2=10.62 //y2=0.45
r232 (  94 140 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.16 //y=0 //x2=9.99 //y2=0
r233 (  93 141 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.535 //y=0 //x2=10.62 //y2=0
r234 (  93 94 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=10.535 //y=0 //x2=10.16 //y2=0
r235 (  88 90 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=8.14 //y=0 //x2=9.25 //y2=0
r236 (  86 139 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.925 //y=0 //x2=7.84 //y2=0
r237 (  86 88 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=7.925 //y=0 //x2=8.14 //y2=0
r238 (  85 140 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.82 //y=0 //x2=9.99 //y2=0
r239 (  85 90 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.82 //y=0 //x2=9.25 //y2=0
r240 (  81 139 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.84 //y=0.17 //x2=7.84 //y2=0
r241 (  81 156 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=7.84 //y=0.17 //x2=7.84 //y2=0.955
r242 (  78 138 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.83 //y=0 //x2=6.66 //y2=0
r243 (  78 80 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=6.83 //y=0 //x2=7.03 //y2=0
r244 (  77 139 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.755 //y=0 //x2=7.84 //y2=0
r245 (  77 80 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=7.755 //y=0 //x2=7.03 //y2=0
r246 (  74 127 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.05 //y=0 //x2=5.965 //y2=0
r247 (  73 138 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.49 //y=0 //x2=6.66 //y2=0
r248 (  73 74 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=6.49 //y=0 //x2=6.05 //y2=0
r249 (  69 155 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.965 //y=0.615 //x2=5.965 //y2=0.53
r250 (  69 155 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=5.965 //y=0.615 //x2=5.965 //y2=0.88
r251 (  68 155 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.965 //y=0.445 //x2=5.965 //y2=0.53
r252 (  67 127 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.965 //y=0.17 //x2=5.965 //y2=0
r253 (  67 68 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=5.965 //y=0.17 //x2=5.965 //y2=0.445
r254 (  66 155 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.565 //y=0.53 //x2=5.48 //y2=0.53
r255 (  65 155 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.88 //y=0.53 //x2=5.965 //y2=0.53
r256 (  65 66 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=5.88 //y=0.53 //x2=5.565 //y2=0.53
r257 (  64 155 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.48 //y=0.445 //x2=5.48 //y2=0.53
r258 (  63 124 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.48 //y=0.17 //x2=5.48 //y2=0
r259 (  63 64 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=5.48 //y=0.17 //x2=5.48 //y2=0.445
r260 (  62 155 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=5.08 //y=0.53 //x2=4.995 //y2=0.53
r261 (  61 155 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.395 //y=0.53 //x2=5.48 //y2=0.53
r262 (  61 62 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=5.395 //y=0.53 //x2=5.08 //y2=0.53
r263 (  57 155 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=4.995 //y=0.615 //x2=4.995 //y2=0.53
r264 (  57 155 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.995 //y=0.615 //x2=4.995 //y2=0.88
r265 (  56 155 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=4.995 //y=0.445 //x2=4.995 //y2=0.53
r266 (  55 123 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.995 //y=0.17 //x2=4.995 //y2=0
r267 (  55 56 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=4.995 //y=0.17 //x2=4.995 //y2=0.445
r268 (  54 155 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.595 //y=0.53 //x2=4.51 //y2=0.53
r269 (  53 155 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=4.91 //y=0.53 //x2=4.995 //y2=0.53
r270 (  53 54 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=4.91 //y=0.53 //x2=4.595 //y2=0.53
r271 (  52 155 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.51 //y=0.445 //x2=4.51 //y2=0.53
r272 (  51 122 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.51 //y=0.17 //x2=4.51 //y2=0
r273 (  51 52 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=4.51 //y=0.17 //x2=4.51 //y2=0.445
r274 (  50 155 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.11 //y=0.53 //x2=4.025 //y2=0.53
r275 (  49 155 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.425 //y=0.53 //x2=4.51 //y2=0.53
r276 (  49 50 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=4.425 //y=0.53 //x2=4.11 //y2=0.53
r277 (  45 155 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.025 //y=0.615 //x2=4.025 //y2=0.53
r278 (  45 155 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=4.025 //y=0.615 //x2=4.025 //y2=1.22
r279 (  44 155 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.025 //y=0.445 //x2=4.025 //y2=0.53
r280 (  43 119 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.025 //y=0.17 //x2=4.025 //y2=0
r281 (  43 44 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=4.025 //y=0.17 //x2=4.025 //y2=0.445
r282 (  42 118 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=0 //x2=3.33 //y2=0
r283 (  41 119 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.94 //y=0 //x2=4.025 //y2=0
r284 (  41 42 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=3.94 //y=0 //x2=3.5 //y2=0
r285 (  36 38 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r286 (  34 117 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.18 //y2=0
r287 (  34 36 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.85 //y2=0
r288 (  33 118 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=3.33 //y2=0
r289 (  33 38 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=2.96 //y2=0
r290 (  29 117 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r291 (  29 154 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.955
r292 (  25 117 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=1.18 //y2=0
r293 (  25 28 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=0.74 //y2=0
r294 (  21 146 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=11.47 //y=0 //x2=11.47 //y2=0
r295 (  19 143 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.73 //y=0 //x2=10.73 //y2=0
r296 (  19 21 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=0 //x2=11.47 //y2=0
r297 (  17 90 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=0 //x2=9.25 //y2=0
r298 (  17 19 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=0 //x2=10.73 //y2=0
r299 (  15 88 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.14 //y=0 //x2=8.14 //y2=0
r300 (  15 17 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=8.14 //y=0 //x2=9.25 //y2=0
r301 (  13 80 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=0 //x2=7.03 //y2=0
r302 (  13 15 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=0 //x2=8.14 //y2=0
r303 (  11 126 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r304 (  11 13 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=7.03 //y2=0
r305 (  9 121 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r306 (  9 11 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.55 //y2=0
r307 (  7 38 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r308 (  7 9 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.44 //y2=0
r309 (  5 36 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r310 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r311 (  2 28 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r312 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
ends PM_AOA4X1_PCELL\%noxref_1

subckt PM_AOA4X1_PCELL\%noxref_2 ( 21 33 41 57 67 83 93 113 126 129 131 136 \
 140 141 142 143 144 145 146 147 148 149 )
c141 ( 149 0 ) capacitor c=0.0451925f //x=11.4 //y=5.02
c142 ( 148 0 ) capacitor c=0.0429269f //x=10.53 //y=5.02
c143 ( 147 0 ) capacitor c=0.0383753f //x=9.065 //y=5.02
c144 ( 146 0 ) capacitor c=0.0243052f //x=8.185 //y=5.02
c145 ( 145 0 ) capacitor c=0.053196f //x=7.315 //y=5.02
c146 ( 144 0 ) capacitor c=0.0256796f //x=4.415 //y=5.025
c147 ( 143 0 ) capacitor c=0.0383753f //x=2.405 //y=5.02
c148 ( 142 0 ) capacitor c=0.0243052f //x=1.525 //y=5.02
c149 ( 141 0 ) capacitor c=0.053196f //x=0.655 //y=5.02
c150 ( 140 0 ) capacitor c=0.234796f //x=11.47 //y=7.4
c151 ( 138 0 ) capacitor c=0.00591168f //x=10.73 //y=7.4
c152 ( 136 0 ) capacitor c=0.111641f //x=9.99 //y=7.4
c153 ( 135 0 ) capacitor c=0.00591168f //x=9.25 //y=7.4
c154 ( 133 0 ) capacitor c=0.00591168f //x=8.33 //y=7.4
c155 ( 132 0 ) capacitor c=0.00591168f //x=7.45 //y=7.4
c156 ( 131 0 ) capacitor c=0.119284f //x=6.66 //y=7.4
c157 ( 130 0 ) capacitor c=0.00591168f //x=4.56 //y=7.4
c158 ( 129 0 ) capacitor c=0.116004f //x=3.33 //y=7.4
c159 ( 128 0 ) capacitor c=0.00591168f //x=2.55 //y=7.4
c160 ( 127 0 ) capacitor c=0.00591168f //x=1.67 //y=7.4
c161 ( 126 0 ) capacitor c=0.24846f //x=0.74 //y=7.4
c162 ( 113 0 ) capacitor c=0.028745f //x=11.46 //y=7.4
c163 ( 105 0 ) capacitor c=0.0216067f //x=10.58 //y=7.4
c164 ( 101 0 ) capacitor c=0.0275781f //x=9.82 //y=7.4
c165 ( 93 0 ) capacitor c=0.0285035f //x=9.125 //y=7.4
c166 ( 83 0 ) capacitor c=0.0286367f //x=8.245 //y=7.4
c167 ( 73 0 ) capacitor c=0.0281468f //x=7.365 //y=7.4
c168 ( 67 0 ) capacitor c=0.0778183f //x=6.49 //y=7.4
c169 ( 57 0 ) capacitor c=0.0465804f //x=4.475 //y=7.4
c170 ( 51 0 ) capacitor c=0.0275781f //x=3.16 //y=7.4
c171 ( 41 0 ) capacitor c=0.0285035f //x=2.465 //y=7.4
c172 ( 33 0 ) capacitor c=0.0286367f //x=1.585 //y=7.4
c173 ( 21 0 ) capacitor c=0.476129f //x=11.47 //y=7.4
r174 (  115 140 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.545 //y=7.23 //x2=11.545 //y2=7.4
r175 (  115 149 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=11.545 //y=7.23 //x2=11.545 //y2=6.405
r176 (  114 138 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.75 //y=7.4 //x2=10.665 //y2=7.4
r177 (  113 140 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.46 //y=7.4 //x2=11.545 //y2=7.4
r178 (  113 114 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.46 //y=7.4 //x2=10.75 //y2=7.4
r179 (  107 138 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.665 //y=7.23 //x2=10.665 //y2=7.4
r180 (  107 148 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=10.665 //y=7.23 //x2=10.665 //y2=6.405
r181 (  106 136 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.16 //y=7.4 //x2=9.99 //y2=7.4
r182 (  105 138 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.58 //y=7.4 //x2=10.665 //y2=7.4
r183 (  105 106 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=10.58 //y=7.4 //x2=10.16 //y2=7.4
r184 (  102 135 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.295 //y=7.4 //x2=9.21 //y2=7.4
r185 (  101 136 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.82 //y=7.4 //x2=9.99 //y2=7.4
r186 (  101 102 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=9.82 //y=7.4 //x2=9.295 //y2=7.4
r187 (  95 135 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.21 //y=7.23 //x2=9.21 //y2=7.4
r188 (  95 147 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=9.21 //y=7.23 //x2=9.21 //y2=6.745
r189 (  94 133 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.415 //y=7.4 //x2=8.33 //y2=7.4
r190 (  93 135 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.125 //y=7.4 //x2=9.21 //y2=7.4
r191 (  93 94 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=9.125 //y=7.4 //x2=8.415 //y2=7.4
r192 (  87 133 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.33 //y=7.23 //x2=8.33 //y2=7.4
r193 (  87 146 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.33 //y=7.23 //x2=8.33 //y2=6.745
r194 (  84 132 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.535 //y=7.4 //x2=7.45 //y2=7.4
r195 (  84 86 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=7.535 //y=7.4 //x2=8.14 //y2=7.4
r196 (  83 133 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.245 //y=7.4 //x2=8.33 //y2=7.4
r197 (  83 86 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=8.245 //y=7.4 //x2=8.14 //y2=7.4
r198 (  77 132 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.45 //y=7.23 //x2=7.45 //y2=7.4
r199 (  77 145 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=7.45 //y=7.23 //x2=7.45 //y2=6.405
r200 (  74 131 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.83 //y=7.4 //x2=6.66 //y2=7.4
r201 (  74 76 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=6.83 //y=7.4 //x2=7.03 //y2=7.4
r202 (  73 132 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.365 //y=7.4 //x2=7.45 //y2=7.4
r203 (  73 76 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=7.365 //y=7.4 //x2=7.03 //y2=7.4
r204 (  68 130 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.645 //y=7.4 //x2=4.56 //y2=7.4
r205 (  68 70 ) resistor r=32.4482 //w=0.357 //l=0.905 //layer=li \
 //thickness=0.1 //x=4.645 //y=7.4 //x2=5.55 //y2=7.4
r206 (  67 131 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.49 //y=7.4 //x2=6.66 //y2=7.4
r207 (  67 70 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=6.49 //y=7.4 //x2=5.55 //y2=7.4
r208 (  61 130 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.56 //y=7.23 //x2=4.56 //y2=7.4
r209 (  61 144 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=4.56 //y=7.23 //x2=4.56 //y2=6.74
r210 (  58 129 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=7.4 //x2=3.33 //y2=7.4
r211 (  58 60 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=3.5 //y=7.4 //x2=4.44 //y2=7.4
r212 (  57 130 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.475 //y=7.4 //x2=4.56 //y2=7.4
r213 (  57 60 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=4.475 //y=7.4 //x2=4.44 //y2=7.4
r214 (  52 128 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.55 //y2=7.4
r215 (  52 54 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.96 //y2=7.4
r216 (  51 129 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=3.33 //y2=7.4
r217 (  51 54 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=2.96 //y2=7.4
r218 (  45 128 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=7.4
r219 (  45 143 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=6.745
r220 (  42 127 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.67 //y2=7.4
r221 (  42 44 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.85 //y2=7.4
r222 (  41 128 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=2.55 //y2=7.4
r223 (  41 44 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=1.85 //y2=7.4
r224 (  35 127 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=7.4
r225 (  35 142 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=6.745
r226 (  34 126 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.875 //y=7.4 //x2=0.79 //y2=7.4
r227 (  33 127 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=1.67 //y2=7.4
r228 (  33 34 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=0.875 //y2=7.4
r229 (  27 126 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=7.4
r230 (  27 141 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=6.405
r231 (  21 140 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=11.47 //y=7.4 //x2=11.47 //y2=7.4
r232 (  19 138 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.73 //y=7.4 //x2=10.73 //y2=7.4
r233 (  19 21 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=10.73 //y=7.4 //x2=11.47 //y2=7.4
r234 (  17 135 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=7.4 //x2=9.25 //y2=7.4
r235 (  17 19 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=7.4 //x2=10.73 //y2=7.4
r236 (  15 86 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.14 //y=7.4 //x2=8.14 //y2=7.4
r237 (  15 17 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=8.14 //y=7.4 //x2=9.25 //y2=7.4
r238 (  13 76 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.03 //y=7.4 //x2=7.03 //y2=7.4
r239 (  13 15 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.03 //y=7.4 //x2=8.14 //y2=7.4
r240 (  11 70 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r241 (  11 13 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=7.03 //y2=7.4
r242 (  9 60 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r243 (  9 11 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.55 //y2=7.4
r244 (  7 54 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r245 (  7 9 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.44 //y2=7.4
r246 (  5 44 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r247 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r248 (  2 126 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r249 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_AOA4X1_PCELL\%noxref_2

subckt PM_AOA4X1_PCELL\%noxref_3 ( 1 2 13 14 25 27 28 32 35 39 41 43 44 45 46 \
 47 48 49 53 55 58 60 61 66 76 78 79 )
c144 ( 79 0 ) capacitor c=0.0220291f //x=1.965 //y=5.02
c145 ( 78 0 ) capacitor c=0.0217503f //x=1.085 //y=5.02
c146 ( 76 0 ) capacitor c=0.00865153f //x=1.96 //y=0.905
c147 ( 66 0 ) capacitor c=0.04214f //x=4.285 //y=4.705
c148 ( 61 0 ) capacitor c=0.0321911f //x=4.775 //y=1.25
c149 ( 60 0 ) capacitor c=0.0185201f //x=4.775 //y=0.905
c150 ( 58 0 ) capacitor c=0.0344254f //x=4.705 //y=4.795
c151 ( 55 0 ) capacitor c=0.0133656f //x=4.62 //y=1.405
c152 ( 53 0 ) capacitor c=0.0157804f //x=4.62 //y=0.75
c153 ( 49 0 ) capacitor c=0.0785055f //x=4.245 //y=1.915
c154 ( 48 0 ) capacitor c=0.022867f //x=4.245 //y=1.56
c155 ( 47 0 ) capacitor c=0.0234318f //x=4.245 //y=1.25
c156 ( 46 0 ) capacitor c=0.0192004f //x=4.245 //y=0.905
c157 ( 45 0 ) capacitor c=0.110795f //x=4.78 //y=6.025
c158 ( 44 0 ) capacitor c=0.153847f //x=4.34 //y=6.025
c159 ( 41 0 ) capacitor c=0.00995068f //x=4.285 //y=4.705
c160 ( 39 0 ) capacitor c=0.00427536f //x=2.11 //y=5.2
c161 ( 35 0 ) capacitor c=0.0968481f //x=4.44 //y=2.08
c162 ( 32 0 ) capacitor c=0.117241f //x=2.59 //y=2.59
c163 ( 28 0 ) capacitor c=0.00781917f //x=2.235 //y=1.655
c164 ( 27 0 ) capacitor c=0.0159132f //x=2.505 //y=1.655
c165 ( 25 0 ) capacitor c=0.017841f //x=2.505 //y=5.2
c166 ( 14 0 ) capacitor c=0.00387264f //x=1.315 //y=5.2
c167 ( 13 0 ) capacitor c=0.0222171f //x=2.025 //y=5.2
c168 ( 2 0 ) capacitor c=0.0173935f //x=2.705 //y=2.59
c169 ( 1 0 ) capacitor c=0.111807f //x=4.325 //y=2.59
r170 (  68 69 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=4.285 //y=4.795 //x2=4.285 //y2=4.87
r171 (  66 68 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=4.285 //y=4.705 //x2=4.285 //y2=4.795
r172 (  61 75 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.775 //y=1.25 //x2=4.735 //y2=1.405
r173 (  60 74 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.775 //y=0.905 //x2=4.735 //y2=0.75
r174 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.775 //y=0.905 //x2=4.775 //y2=1.25
r175 (  59 68 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=4.42 //y=4.795 //x2=4.285 //y2=4.795
r176 (  58 62 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.705 //y=4.795 //x2=4.78 //y2=4.87
r177 (  58 59 ) resistor r=146.138 //w=0.094 //l=0.285 //layer=ply \
 //thickness=0.18 //x=4.705 //y=4.795 //x2=4.42 //y2=4.795
r178 (  56 73 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.4 //y=1.405 //x2=4.285 //y2=1.405
r179 (  55 75 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.62 //y=1.405 //x2=4.735 //y2=1.405
r180 (  54 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.4 //y=0.75 //x2=4.285 //y2=0.75
r181 (  53 74 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.62 //y=0.75 //x2=4.735 //y2=0.75
r182 (  53 54 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.62 //y=0.75 //x2=4.4 //y2=0.75
r183 (  49 71 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=4.245 //y=1.915 //x2=4.44 //y2=2.08
r184 (  48 73 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.245 //y=1.56 //x2=4.285 //y2=1.405
r185 (  48 49 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=4.245 //y=1.56 //x2=4.245 //y2=1.915
r186 (  47 73 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.245 //y=1.25 //x2=4.285 //y2=1.405
r187 (  46 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.245 //y=0.905 //x2=4.285 //y2=0.75
r188 (  46 47 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.245 //y=0.905 //x2=4.245 //y2=1.25
r189 (  45 62 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.78 //y=6.025 //x2=4.78 //y2=4.87
r190 (  44 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.34 //y=6.025 //x2=4.34 //y2=4.87
r191 (  43 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.51 //y=1.405 //x2=4.62 //y2=1.405
r192 (  43 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.51 //y=1.405 //x2=4.4 //y2=1.405
r193 (  41 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.285 //y=4.705 //x2=4.285 //y2=4.705
r194 (  41 42 ) resistor r=7.81102 //w=0.254 //l=0.155 //layer=li \
 //thickness=0.1 //x=4.285 //y=4.705 //x2=4.44 //y2=4.705
r195 (  35 71 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=2.08 //x2=4.44 //y2=2.08
r196 (  35 38 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.08 //x2=4.44 //y2=2.59
r197 (  33 42 ) resistor r=3.23951 //w=0.254 //l=0.165 //layer=li \
 //thickness=0.1 //x=4.44 //y=4.54 //x2=4.44 //y2=4.705
r198 (  33 38 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=4.44 //y=4.54 //x2=4.44 //y2=2.59
r199 (  30 32 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=2.59 //y=5.115 //x2=2.59 //y2=2.59
r200 (  29 32 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=2.59 //y=1.74 //x2=2.59 //y2=2.59
r201 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.59 //y2=1.74
r202 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.235 //y2=1.655
r203 (  26 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.195 //y=5.2 //x2=2.11 //y2=5.2
r204 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.59 //y2=5.115
r205 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.195 //y2=5.2
r206 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.235 //y2=1.655
r207 (  21 76 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r208 (  15 39 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.2
r209 (  15 79 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.725
r210 (  13 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=2.11 //y2=5.2
r211 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=1.315 //y2=5.2
r212 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.315 //y2=5.2
r213 (  7 78 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.23 //y2=5.725
r214 (  6 38 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.44 //y=2.59 //x2=4.44 //y2=2.59
r215 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.59 //y=2.59 //x2=2.59 //y2=2.59
r216 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.705 //y=2.59 //x2=2.59 //y2=2.59
r217 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.325 //y=2.59 //x2=4.44 //y2=2.59
r218 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=4.325 //y=2.59 //x2=2.705 //y2=2.59
ends PM_AOA4X1_PCELL\%noxref_3

subckt PM_AOA4X1_PCELL\%noxref_4 ( 1 2 11 12 23 24 25 30 32 40 41 42 43 44 45 \
 46 50 52 55 56 66 69 70 73 )
c142 ( 73 0 ) capacitor c=0.0159573f //x=5.295 //y=5.025
c143 ( 70 0 ) capacitor c=0.00925154f //x=5.29 //y=0.905
c144 ( 69 0 ) capacitor c=0.007684f //x=4.32 //y=0.905
c145 ( 66 0 ) capacitor c=0.0667949f //x=7.77 //y=4.7
c146 ( 56 0 ) capacitor c=0.0318948f //x=8.105 //y=1.21
c147 ( 55 0 ) capacitor c=0.0187384f //x=8.105 //y=0.865
c148 ( 52 0 ) capacitor c=0.0141798f //x=7.95 //y=1.365
c149 ( 50 0 ) capacitor c=0.0149844f //x=7.95 //y=0.71
c150 ( 46 0 ) capacitor c=0.0816272f //x=7.575 //y=1.915
c151 ( 45 0 ) capacitor c=0.0229531f //x=7.575 //y=1.52
c152 ( 44 0 ) capacitor c=0.0234352f //x=7.575 //y=1.21
c153 ( 43 0 ) capacitor c=0.0199343f //x=7.575 //y=0.865
c154 ( 42 0 ) capacitor c=0.110275f //x=8.11 //y=6.02
c155 ( 41 0 ) capacitor c=0.154305f //x=7.67 //y=6.02
c156 ( 39 0 ) capacitor c=0.00710337f //x=5.48 //y=1.655
c157 ( 32 0 ) capacitor c=0.101048f //x=7.77 //y=2.08
c158 ( 30 0 ) capacitor c=0.117944f //x=5.92 //y=2.59
c159 ( 25 0 ) capacitor c=0.0160526f //x=5.835 //y=1.655
c160 ( 24 0 ) capacitor c=0.00499395f //x=5.525 //y=5.21
c161 ( 23 0 ) capacitor c=0.0164583f //x=5.835 //y=5.21
c162 ( 12 0 ) capacitor c=0.00220849f //x=4.595 //y=1.655
c163 ( 11 0 ) capacitor c=0.0280953f //x=5.395 //y=1.655
c164 ( 2 0 ) capacitor c=0.0120303f //x=6.035 //y=2.59
c165 ( 1 0 ) capacitor c=0.112452f //x=7.655 //y=2.59
r166 (  64 66 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=7.67 //y=4.7 //x2=7.77 //y2=4.7
r167 (  57 66 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=8.11 //y=4.865 //x2=7.77 //y2=4.7
r168 (  56 68 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.105 //y=1.21 //x2=8.065 //y2=1.365
r169 (  55 67 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.105 //y=0.865 //x2=8.065 //y2=0.71
r170 (  55 56 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.105 //y=0.865 //x2=8.105 //y2=1.21
r171 (  53 63 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.73 //y=1.365 //x2=7.615 //y2=1.365
r172 (  52 68 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.95 //y=1.365 //x2=8.065 //y2=1.365
r173 (  51 62 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.73 //y=0.71 //x2=7.615 //y2=0.71
r174 (  50 67 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.95 //y=0.71 //x2=8.065 //y2=0.71
r175 (  50 51 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.95 //y=0.71 //x2=7.73 //y2=0.71
r176 (  47 64 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=7.67 //y=4.865 //x2=7.67 //y2=4.7
r177 (  46 61 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=7.575 //y=1.915 //x2=7.77 //y2=2.08
r178 (  45 63 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.575 //y=1.52 //x2=7.615 //y2=1.365
r179 (  45 46 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=7.575 //y=1.52 //x2=7.575 //y2=1.915
r180 (  44 63 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.575 //y=1.21 //x2=7.615 //y2=1.365
r181 (  43 62 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.575 //y=0.865 //x2=7.615 //y2=0.71
r182 (  43 44 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.575 //y=0.865 //x2=7.575 //y2=1.21
r183 (  42 57 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.11 //y=6.02 //x2=8.11 //y2=4.865
r184 (  41 47 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.67 //y=6.02 //x2=7.67 //y2=4.865
r185 (  40 52 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.84 //y=1.365 //x2=7.95 //y2=1.365
r186 (  40 53 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=7.84 //y=1.365 //x2=7.73 //y2=1.365
r187 (  37 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.77 //y=4.7 //x2=7.77 //y2=4.7
r188 (  35 37 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=7.77 //y=2.59 //x2=7.77 //y2=4.7
r189 (  32 61 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.77 //y=2.08 //x2=7.77 //y2=2.08
r190 (  32 35 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=7.77 //y=2.08 //x2=7.77 //y2=2.59
r191 (  28 30 ) resistor r=173.519 //w=0.187 //l=2.535 //layer=li \
 //thickness=0.1 //x=5.92 //y=5.125 //x2=5.92 //y2=2.59
r192 (  27 30 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=5.92 //y=1.74 //x2=5.92 //y2=2.59
r193 (  26 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.565 //y=1.655 //x2=5.48 //y2=1.655
r194 (  25 27 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5.835 //y=1.655 //x2=5.92 //y2=1.74
r195 (  25 26 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=5.835 //y=1.655 //x2=5.565 //y2=1.655
r196 (  23 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5.835 //y=5.21 //x2=5.92 //y2=5.125
r197 (  23 24 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=5.835 //y=5.21 //x2=5.525 //y2=5.21
r198 (  19 39 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.48 //y=1.57 //x2=5.48 //y2=1.655
r199 (  19 70 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=5.48 //y=1.57 //x2=5.48 //y2=1
r200 (  13 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5.44 //y=5.295 //x2=5.525 //y2=5.21
r201 (  13 73 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=5.44 //y=5.295 //x2=5.44 //y2=5.72
r202 (  11 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.395 //y=1.655 //x2=5.48 //y2=1.655
r203 (  11 12 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li \
 //thickness=0.1 //x=5.395 //y=1.655 //x2=4.595 //y2=1.655
r204 (  7 12 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.51 //y=1.57 //x2=4.595 //y2=1.655
r205 (  7 69 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=4.51 //y=1.57 //x2=4.51 //y2=1
r206 (  6 35 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.77 //y=2.59 //x2=7.77 //y2=2.59
r207 (  4 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.92 //y=2.59 //x2=5.92 //y2=2.59
r208 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.035 //y=2.59 //x2=5.92 //y2=2.59
r209 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.655 //y=2.59 //x2=7.77 //y2=2.59
r210 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=7.655 //y=2.59 //x2=6.035 //y2=2.59
ends PM_AOA4X1_PCELL\%noxref_4

subckt PM_AOA4X1_PCELL\%noxref_5 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 \
 47 48 52 53 54 56 62 63 65 73 75 76 )
c126 ( 76 0 ) capacitor c=0.0220291f //x=8.625 //y=5.02
c127 ( 75 0 ) capacitor c=0.0217503f //x=7.745 //y=5.02
c128 ( 73 0 ) capacitor c=0.0084702f //x=8.62 //y=0.905
c129 ( 65 0 ) capacitor c=0.0517753f //x=10.73 //y=2.085
c130 ( 63 0 ) capacitor c=0.0435629f //x=11.37 //y=1.255
c131 ( 62 0 ) capacitor c=0.0200386f //x=11.37 //y=0.91
c132 ( 56 0 ) capacitor c=0.0152946f //x=11.215 //y=1.41
c133 ( 54 0 ) capacitor c=0.0157804f //x=11.215 //y=0.755
c134 ( 53 0 ) capacitor c=0.0524991f //x=10.96 //y=4.79
c135 ( 52 0 ) capacitor c=0.0322983f //x=11.25 //y=4.79
c136 ( 48 0 ) capacitor c=0.0290017f //x=10.84 //y=1.92
c137 ( 47 0 ) capacitor c=0.0250027f //x=10.84 //y=1.565
c138 ( 46 0 ) capacitor c=0.0234316f //x=10.84 //y=1.255
c139 ( 45 0 ) capacitor c=0.0200596f //x=10.84 //y=0.91
c140 ( 44 0 ) capacitor c=0.154218f //x=11.325 //y=6.02
c141 ( 43 0 ) capacitor c=0.154243f //x=10.885 //y=6.02
c142 ( 41 0 ) capacitor c=0.00427536f //x=8.77 //y=5.2
c143 ( 34 0 ) capacitor c=0.0948753f //x=10.73 //y=2.085
c144 ( 32 0 ) capacitor c=0.113415f //x=9.25 //y=2.59
c145 ( 28 0 ) capacitor c=0.00781917f //x=8.895 //y=1.655
c146 ( 27 0 ) capacitor c=0.0159132f //x=9.165 //y=1.655
c147 ( 25 0 ) capacitor c=0.0180264f //x=9.165 //y=5.2
c148 ( 14 0 ) capacitor c=0.00391676f //x=7.975 //y=5.2
c149 ( 13 0 ) capacitor c=0.0222171f //x=8.685 //y=5.2
c150 ( 2 0 ) capacitor c=0.0119586f //x=9.365 //y=2.59
c151 ( 1 0 ) capacitor c=0.0934424f //x=10.615 //y=2.59
r152 (  65 66 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.73 //y=2.085 //x2=10.84 //y2=2.085
r153 (  63 72 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.37 //y=1.255 //x2=11.33 //y2=1.41
r154 (  62 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.37 //y=0.91 //x2=11.33 //y2=0.755
r155 (  62 63 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.37 //y=0.91 //x2=11.37 //y2=1.255
r156 (  57 70 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.995 //y=1.41 //x2=10.88 //y2=1.41
r157 (  56 72 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.215 //y=1.41 //x2=11.33 //y2=1.41
r158 (  55 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.995 //y=0.755 //x2=10.88 //y2=0.755
r159 (  54 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.215 //y=0.755 //x2=11.33 //y2=0.755
r160 (  54 55 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=11.215 //y=0.755 //x2=10.995 //y2=0.755
r161 (  52 59 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=11.25 //y=4.79 //x2=11.325 //y2=4.865
r162 (  52 53 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=11.25 //y=4.79 //x2=10.96 //y2=4.79
r163 (  49 53 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.885 //y=4.865 //x2=10.96 //y2=4.79
r164 (  49 68 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=10.885 //y=4.865 //x2=10.73 //y2=4.7
r165 (  48 66 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=10.84 //y=1.92 //x2=10.84 //y2=2.085
r166 (  47 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.84 //y=1.565 //x2=10.88 //y2=1.41
r167 (  47 48 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=10.84 //y=1.565 //x2=10.84 //y2=1.92
r168 (  46 70 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.84 //y=1.255 //x2=10.88 //y2=1.41
r169 (  45 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.84 //y=0.91 //x2=10.88 //y2=0.755
r170 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.84 //y=0.91 //x2=10.84 //y2=1.255
r171 (  44 59 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.325 //y=6.02 //x2=11.325 //y2=4.865
r172 (  43 49 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.885 //y=6.02 //x2=10.885 //y2=4.865
r173 (  42 56 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.105 //y=1.41 //x2=11.215 //y2=1.41
r174 (  42 57 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.105 //y=1.41 //x2=10.995 //y2=1.41
r175 (  39 68 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=4.7 //x2=10.73 //y2=4.7
r176 (  37 39 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.59 //x2=10.73 //y2=4.7
r177 (  34 65 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=2.085 //x2=10.73 //y2=2.085
r178 (  34 37 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.085 //x2=10.73 //y2=2.59
r179 (  30 32 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=9.25 //y=5.115 //x2=9.25 //y2=2.59
r180 (  29 32 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=9.25 //y=1.74 //x2=9.25 //y2=2.59
r181 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.165 //y=1.655 //x2=9.25 //y2=1.74
r182 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=9.165 //y=1.655 //x2=8.895 //y2=1.655
r183 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.855 //y=5.2 //x2=8.77 //y2=5.2
r184 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.165 //y=5.2 //x2=9.25 //y2=5.115
r185 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=9.165 //y=5.2 //x2=8.855 //y2=5.2
r186 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.81 //y=1.57 //x2=8.895 //y2=1.655
r187 (  21 73 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=8.81 //y=1.57 //x2=8.81 //y2=1
r188 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.77 //y=5.285 //x2=8.77 //y2=5.2
r189 (  15 76 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=8.77 //y=5.285 //x2=8.77 //y2=5.725
r190 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.685 //y=5.2 //x2=8.77 //y2=5.2
r191 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.685 //y=5.2 //x2=7.975 //y2=5.2
r192 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.89 //y=5.285 //x2=7.975 //y2=5.2
r193 (  7 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=7.89 //y=5.285 //x2=7.89 //y2=5.725
r194 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.73 //y=2.59 //x2=10.73 //y2=2.59
r195 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.25 //y=2.59 //x2=9.25 //y2=2.59
r196 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.365 //y=2.59 //x2=9.25 //y2=2.59
r197 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=2.59 //x2=10.73 //y2=2.59
r198 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=2.59 //x2=9.365 //y2=2.59
ends PM_AOA4X1_PCELL\%noxref_5

subckt PM_AOA4X1_PCELL\%noxref_6 ( 2 7 8 9 10 11 12 13 17 19 22 23 33 )
c55 ( 33 0 ) capacitor c=0.0667949f //x=1.11 //y=4.7
c56 ( 23 0 ) capacitor c=0.0318948f //x=1.445 //y=1.21
c57 ( 22 0 ) capacitor c=0.0187384f //x=1.445 //y=0.865
c58 ( 19 0 ) capacitor c=0.0141798f //x=1.29 //y=1.365
c59 ( 17 0 ) capacitor c=0.0149844f //x=1.29 //y=0.71
c60 ( 13 0 ) capacitor c=0.0860049f //x=0.915 //y=1.915
c61 ( 12 0 ) capacitor c=0.0229722f //x=0.915 //y=1.52
c62 ( 11 0 ) capacitor c=0.0234352f //x=0.915 //y=1.21
c63 ( 10 0 ) capacitor c=0.0199343f //x=0.915 //y=0.865
c64 ( 9 0 ) capacitor c=0.110275f //x=1.45 //y=6.02
c65 ( 8 0 ) capacitor c=0.154305f //x=1.01 //y=6.02
c66 ( 2 0 ) capacitor c=0.116498f //x=1.11 //y=2.08
r67 (  31 33 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.7 //x2=1.11 //y2=4.7
r68 (  24 33 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=1.45 //y=4.865 //x2=1.11 //y2=4.7
r69 (  23 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.21 //x2=1.405 //y2=1.365
r70 (  22 34 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.405 //y2=0.71
r71 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.445 //y2=1.21
r72 (  20 30 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.365 //x2=0.955 //y2=1.365
r73 (  19 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.365 //x2=1.405 //y2=1.365
r74 (  18 29 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.71 //x2=0.955 //y2=0.71
r75 (  17 34 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.405 //y2=0.71
r76 (  17 18 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.07 //y2=0.71
r77 (  14 31 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.865 //x2=1.01 //y2=4.7
r78 (  13 28 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r79 (  12 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.955 //y2=1.365
r80 (  12 13 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.915 //y2=1.915
r81 (  11 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.21 //x2=0.955 //y2=1.365
r82 (  10 29 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.955 //y2=0.71
r83 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.915 //y2=1.21
r84 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.02 //x2=1.45 //y2=4.865
r85 (  8 14 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.02 //x2=1.01 //y2=4.865
r86 (  7 19 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.29 //y2=1.365
r87 (  7 20 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.07 //y2=1.365
r88 (  5 33 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r89 (  2 28 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r90 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=4.7
ends PM_AOA4X1_PCELL\%noxref_6

subckt PM_AOA4X1_PCELL\%noxref_7 ( 1 3 7 8 9 10 11 12 17 19 21 27 28 30 31 34 )
c64 ( 34 0 ) capacitor c=0.034715f //x=1.88 //y=4.7
c65 ( 31 0 ) capacitor c=0.0279499f //x=1.85 //y=1.915
c66 ( 30 0 ) capacitor c=0.0437302f //x=1.85 //y=2.08
c67 ( 28 0 ) capacitor c=0.0429696f //x=2.415 //y=1.25
c68 ( 27 0 ) capacitor c=0.0192208f //x=2.415 //y=0.905
c69 ( 21 0 ) capacitor c=0.0158629f //x=2.26 //y=1.405
c70 ( 19 0 ) capacitor c=0.0157803f //x=2.26 //y=0.75
c71 ( 17 0 ) capacitor c=0.0366192f //x=2.255 //y=4.79
c72 ( 12 0 ) capacitor c=0.0205163f //x=1.885 //y=1.56
c73 ( 11 0 ) capacitor c=0.0168481f //x=1.885 //y=1.25
c74 ( 10 0 ) capacitor c=0.0174783f //x=1.885 //y=0.905
c75 ( 9 0 ) capacitor c=0.15358f //x=2.33 //y=6.02
c76 ( 8 0 ) capacitor c=0.110281f //x=1.89 //y=6.02
c77 ( 3 0 ) capacitor c=0.0813556f //x=1.85 //y=2.08
c78 ( 1 0 ) capacitor c=0.00453889f //x=1.85 //y=4.535
r79 (  36 37 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.79 //x2=1.88 //y2=4.865
r80 (  34 36 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.7 //x2=1.88 //y2=4.79
r81 (  30 31 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r82 (  28 41 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.25 //x2=2.375 //y2=1.405
r83 (  27 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r84 (  27 28 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.25
r85 (  22 39 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r86 (  21 41 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.375 //y2=1.405
r87 (  20 38 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r88 (  19 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r89 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r90 (  18 36 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.015 //y=4.79 //x2=1.88 //y2=4.79
r91 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.33 //y2=4.865
r92 (  17 18 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.015 //y2=4.79
r93 (  12 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r94 (  12 31 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r95 (  11 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.25 //x2=1.925 //y2=1.405
r96 (  10 38 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r97 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.25
r98 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.02 //x2=2.33 //y2=4.865
r99 (  8 37 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.02 //x2=1.89 //y2=4.865
r100 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r101 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r102 (  6 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.88 //y=4.7 //x2=1.88 //y2=4.7
r103 (  3 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r104 (  1 6 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.865 //y2=4.7
r105 (  1 3 ) resistor r=168.043 //w=0.187 //l=2.455 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.85 //y2=2.08
ends PM_AOA4X1_PCELL\%noxref_7

subckt PM_AOA4X1_PCELL\%noxref_8 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632971f //x=0.56 //y=0.365
c52 ( 17 0 ) capacitor c=0.00722223f //x=2.635 //y=0.615
c53 ( 13 0 ) capacitor c=0.0154397f //x=2.55 //y=0.53
c54 ( 10 0 ) capacitor c=0.0092508f //x=1.665 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=1.665 //y=0.615
c56 ( 5 0 ) capacitor c=0.0255599f //x=1.58 //y=1.58
c57 ( 1 0 ) capacitor c=0.0113547f //x=0.695 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.75 //y=0.53 //x2=1.665 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=2.15 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.55 //y=0.53 //x2=2.15 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.78 //y=1.58 //x2=0.695 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.78 //y=1.58 //x2=1.18 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.58 //y=1.58 //x2=1.665 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.58 //y=1.58 //x2=1.18 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.695 //y=1.495 //x2=0.695 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.695 //y=1.495 //x2=0.695 //y2=0.88
ends PM_AOA4X1_PCELL\%noxref_8

subckt PM_AOA4X1_PCELL\%noxref_9 ( 1 3 7 8 9 10 11 12 17 19 21 27 28 30 31 34 )
c71 ( 34 0 ) capacitor c=0.0369822f //x=5.215 //y=4.705
c72 ( 31 0 ) capacitor c=0.0279572f //x=5.18 //y=1.915
c73 ( 30 0 ) capacitor c=0.0422144f //x=5.18 //y=2.08
c74 ( 28 0 ) capacitor c=0.0237734f //x=5.745 //y=1.255
c75 ( 27 0 ) capacitor c=0.0191782f //x=5.745 //y=0.905
c76 ( 21 0 ) capacitor c=0.0346941f //x=5.59 //y=1.405
c77 ( 19 0 ) capacitor c=0.0157803f //x=5.59 //y=0.75
c78 ( 17 0 ) capacitor c=0.0359964f //x=5.585 //y=4.795
c79 ( 12 0 ) capacitor c=0.0199921f //x=5.215 //y=1.56
c80 ( 11 0 ) capacitor c=0.0169608f //x=5.215 //y=1.255
c81 ( 10 0 ) capacitor c=0.0185462f //x=5.215 //y=0.905
c82 ( 9 0 ) capacitor c=0.15325f //x=5.66 //y=6.025
c83 ( 8 0 ) capacitor c=0.110232f //x=5.22 //y=6.025
c84 ( 3 0 ) capacitor c=0.0800125f //x=5.18 //y=2.08
c85 ( 1 0 ) capacitor c=0.00521267f //x=5.18 //y=4.54
r86 (  36 37 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=5.215 //y=4.795 //x2=5.215 //y2=4.87
r87 (  34 36 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=5.215 //y=4.705 //x2=5.215 //y2=4.795
r88 (  30 31 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=5.18 //y=2.08 //x2=5.18 //y2=1.915
r89 (  28 41 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=5.745 //y=1.255 //x2=5.745 //y2=1.367
r90 (  27 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.745 //y=0.905 //x2=5.705 //y2=0.75
r91 (  27 28 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=5.745 //y=0.905 //x2=5.745 //y2=1.255
r92 (  22 39 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.37 //y=1.405 //x2=5.255 //y2=1.405
r93 (  21 41 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=5.59 //y=1.405 //x2=5.745 //y2=1.367
r94 (  20 38 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.37 //y=0.75 //x2=5.255 //y2=0.75
r95 (  19 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.59 //y=0.75 //x2=5.705 //y2=0.75
r96 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=5.59 //y=0.75 //x2=5.37 //y2=0.75
r97 (  18 36 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=5.35 //y=4.795 //x2=5.215 //y2=4.795
r98 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.585 //y=4.795 //x2=5.66 //y2=4.87
r99 (  17 18 ) resistor r=120.5 //w=0.094 //l=0.235 //layer=ply \
 //thickness=0.18 //x=5.585 //y=4.795 //x2=5.35 //y2=4.795
r100 (  12 39 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.215 //y=1.56 //x2=5.255 //y2=1.405
r101 (  12 31 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=5.215 //y=1.56 //x2=5.215 //y2=1.915
r102 (  11 39 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=5.215 //y=1.255 //x2=5.255 //y2=1.405
r103 (  10 38 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.215 //y=0.905 //x2=5.255 //y2=0.75
r104 (  10 11 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=5.215 //y=0.905 //x2=5.215 //y2=1.255
r105 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.66 //y=6.025 //x2=5.66 //y2=4.87
r106 (  8 37 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.22 //y=6.025 //x2=5.22 //y2=4.87
r107 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.48 //y=1.405 //x2=5.59 //y2=1.405
r108 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.48 //y=1.405 //x2=5.37 //y2=1.405
r109 (  6 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.215 //y=4.705 //x2=5.215 //y2=4.705
r110 (  3 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.18 //y=2.08 //x2=5.18 //y2=2.08
r111 (  1 6 ) resistor r=11.332 //w=0.189 //l=0.173292 //layer=li \
 //thickness=0.1 //x=5.18 //y=4.54 //x2=5.197 //y2=4.705
r112 (  1 3 ) resistor r=168.385 //w=0.187 //l=2.46 //layer=li //thickness=0.1 \
 //x=5.18 //y=4.54 //x2=5.18 //y2=2.08
ends PM_AOA4X1_PCELL\%noxref_9

subckt PM_AOA4X1_PCELL\%noxref_10 ( 7 8 15 16 23 24 25 )
c43 ( 25 0 ) capacitor c=0.0308836f //x=5.735 //y=5.025
c44 ( 24 0 ) capacitor c=0.0185379f //x=4.855 //y=5.025
c45 ( 23 0 ) capacitor c=0.0409962f //x=3.985 //y=5.025
c46 ( 16 0 ) capacitor c=0.00193672f //x=5.085 //y=6.91
c47 ( 15 0 ) capacitor c=0.01354f //x=5.795 //y=6.91
c48 ( 8 0 ) capacitor c=0.00844339f //x=4.205 //y=5.21
c49 ( 7 0 ) capacitor c=0.0252644f //x=4.915 //y=5.21
r50 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.88 //y=6.825 //x2=5.88 //y2=6.74
r51 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5.795 //y=6.91 //x2=5.88 //y2=6.825
r52 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=5.795 //y=6.91 //x2=5.085 //y2=6.91
r53 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5 //y=6.825 //x2=5.085 //y2=6.91
r54 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=5 //y=6.825 //x2=5 //y2=6.4
r55 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=5 //y=5.295 //x2=5 //y2=5.72
r56 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.915 //y=5.21 //x2=5 //y2=5.295
r57 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=4.915 //y=5.21 //x2=4.205 //y2=5.21
r58 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.12 //y=5.295 //x2=4.205 //y2=5.21
r59 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=4.12 //y=5.295 //x2=4.12 //y2=5.72
ends PM_AOA4X1_PCELL\%noxref_10

subckt PM_AOA4X1_PCELL\%noxref_11 ( 1 3 7 8 9 10 11 12 17 19 21 27 28 30 31 34 )
c66 ( 34 0 ) capacitor c=0.034715f //x=8.54 //y=4.7
c67 ( 31 0 ) capacitor c=0.0279499f //x=8.51 //y=1.915
c68 ( 30 0 ) capacitor c=0.0437302f //x=8.51 //y=2.08
c69 ( 28 0 ) capacitor c=0.0429696f //x=9.075 //y=1.25
c70 ( 27 0 ) capacitor c=0.0192208f //x=9.075 //y=0.905
c71 ( 21 0 ) capacitor c=0.0158629f //x=8.92 //y=1.405
c72 ( 19 0 ) capacitor c=0.0157803f //x=8.92 //y=0.75
c73 ( 17 0 ) capacitor c=0.0367015f //x=8.915 //y=4.79
c74 ( 12 0 ) capacitor c=0.0205163f //x=8.545 //y=1.56
c75 ( 11 0 ) capacitor c=0.0168481f //x=8.545 //y=1.25
c76 ( 10 0 ) capacitor c=0.0174783f //x=8.545 //y=0.905
c77 ( 9 0 ) capacitor c=0.15358f //x=8.99 //y=6.02
c78 ( 8 0 ) capacitor c=0.110281f //x=8.55 //y=6.02
c79 ( 3 0 ) capacitor c=0.0804986f //x=8.51 //y=2.08
c80 ( 1 0 ) capacitor c=0.00453889f //x=8.51 //y=4.535
r81 (  36 37 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=8.54 //y=4.79 //x2=8.54 //y2=4.865
r82 (  34 36 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=8.54 //y=4.7 //x2=8.54 //y2=4.79
r83 (  30 31 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=8.51 //y=2.08 //x2=8.51 //y2=1.915
r84 (  28 41 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.075 //y=1.25 //x2=9.035 //y2=1.405
r85 (  27 40 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.075 //y=0.905 //x2=9.035 //y2=0.75
r86 (  27 28 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.075 //y=0.905 //x2=9.075 //y2=1.25
r87 (  22 39 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.7 //y=1.405 //x2=8.585 //y2=1.405
r88 (  21 41 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.92 //y=1.405 //x2=9.035 //y2=1.405
r89 (  20 38 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.7 //y=0.75 //x2=8.585 //y2=0.75
r90 (  19 40 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.92 //y=0.75 //x2=9.035 //y2=0.75
r91 (  19 20 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=8.92 //y=0.75 //x2=8.7 //y2=0.75
r92 (  18 36 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=8.675 //y=4.79 //x2=8.54 //y2=4.79
r93 (  17 24 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=8.915 //y=4.79 //x2=8.99 //y2=4.865
r94 (  17 18 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=8.915 //y=4.79 //x2=8.675 //y2=4.79
r95 (  12 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.545 //y=1.56 //x2=8.585 //y2=1.405
r96 (  12 31 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=8.545 //y=1.56 //x2=8.545 //y2=1.915
r97 (  11 39 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.545 //y=1.25 //x2=8.585 //y2=1.405
r98 (  10 38 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.545 //y=0.905 //x2=8.585 //y2=0.75
r99 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.545 //y=0.905 //x2=8.545 //y2=1.25
r100 (  9 24 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.99 //y=6.02 //x2=8.99 //y2=4.865
r101 (  8 37 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.55 //y=6.02 //x2=8.55 //y2=4.865
r102 (  7 21 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.81 //y=1.405 //x2=8.92 //y2=1.405
r103 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.81 //y=1.405 //x2=8.7 //y2=1.405
r104 (  6 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.54 //y=4.7 //x2=8.54 //y2=4.7
r105 (  3 30 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.51 //y=2.08 //x2=8.51 //y2=2.08
r106 (  1 6 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=8.51 //y=4.535 //x2=8.525 //y2=4.7
r107 (  1 3 ) resistor r=168.043 //w=0.187 //l=2.455 //layer=li \
 //thickness=0.1 //x=8.51 //y=4.535 //x2=8.51 //y2=2.08
ends PM_AOA4X1_PCELL\%noxref_11

subckt PM_AOA4X1_PCELL\%noxref_12 ( 1 5 9 10 13 17 29 )
c55 ( 29 0 ) capacitor c=0.0632684f //x=7.22 //y=0.365
c56 ( 17 0 ) capacitor c=0.00722223f //x=9.295 //y=0.615
c57 ( 13 0 ) capacitor c=0.0154397f //x=9.21 //y=0.53
c58 ( 10 0 ) capacitor c=0.0092508f //x=8.325 //y=1.495
c59 ( 9 0 ) capacitor c=0.006761f //x=8.325 //y=0.615
c60 ( 5 0 ) capacitor c=0.0235093f //x=8.24 //y=1.58
c61 ( 1 0 ) capacitor c=0.00765941f //x=7.355 //y=1.495
r62 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=9.295 //y=0.615 //x2=9.295 //y2=0.49
r63 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=9.295 //y=0.615 //x2=9.295 //y2=0.88
r64 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.41 //y=0.53 //x2=8.325 //y2=0.49
r65 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.41 //y=0.53 //x2=8.81 //y2=0.53
r66 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.21 //y=0.53 //x2=9.295 //y2=0.49
r67 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.21 //y=0.53 //x2=8.81 //y2=0.53
r68 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=8.325 //y=1.495 //x2=8.325 //y2=1.62
r69 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=8.325 //y=1.495 //x2=8.325 //y2=0.88
r70 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=8.325 //y=0.615 //x2=8.325 //y2=0.49
r71 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=8.325 //y=0.615 //x2=8.325 //y2=0.88
r72 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.44 //y=1.58 //x2=7.355 //y2=1.62
r73 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.44 //y=1.58 //x2=7.84 //y2=1.58
r74 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.24 //y=1.58 //x2=8.325 //y2=1.62
r75 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.24 //y=1.58 //x2=7.84 //y2=1.58
r76 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=7.355 //y=1.495 //x2=7.355 //y2=1.62
r77 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=7.355 //y=1.495 //x2=7.355 //y2=0.88
ends PM_AOA4X1_PCELL\%noxref_12

subckt PM_AOA4X1_PCELL\%noxref_13 ( 11 12 13 14 16 17 19 )
c43 ( 19 0 ) capacitor c=0.028734f //x=10.96 //y=5.02
c44 ( 17 0 ) capacitor c=0.0173218f //x=10.915 //y=0.91
c45 ( 16 0 ) capacitor c=0.105613f //x=11.47 //y=4.495
c46 ( 14 0 ) capacitor c=0.00575887f //x=11.19 //y=4.58
c47 ( 13 0 ) capacitor c=0.0146395f //x=11.385 //y=4.58
c48 ( 12 0 ) capacitor c=0.00636159f //x=11.185 //y=2.08
c49 ( 11 0 ) capacitor c=0.0141837f //x=11.385 //y=2.08
r50 (  15 16 ) resistor r=159.487 //w=0.187 //l=2.33 //layer=li \
 //thickness=0.1 //x=11.47 //y=2.165 //x2=11.47 //y2=4.495
r51 (  13 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.385 //y=4.58 //x2=11.47 //y2=4.495
r52 (  13 14 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=11.385 //y=4.58 //x2=11.19 //y2=4.58
r53 (  11 15 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.385 //y=2.08 //x2=11.47 //y2=2.165
r54 (  11 12 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=11.385 //y=2.08 //x2=11.185 //y2=2.08
r55 (  5 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.105 //y=4.665 //x2=11.19 //y2=4.58
r56 (  5 19 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li //thickness=0.1 \
 //x=11.105 //y=4.665 //x2=11.105 //y2=5.725
r57 (  1 12 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.1 //y=1.995 //x2=11.185 //y2=2.08
r58 (  1 17 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=11.1 //y=1.995 //x2=11.1 //y2=1.005
ends PM_AOA4X1_PCELL\%noxref_13

