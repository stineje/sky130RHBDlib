* SPICE3 file created from DFFSNQNX1.ext - technology: sky130A

.subckt DFFSNQNX1 QN D CLK SN VPB VNB
M1000 VNB a_168_157# a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1001 VNB a_343_383.t12 a_3368_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_3599_383.t6 SN VPB.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t6 a_168_157# a_217_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPB.t22 a_1265_943.t5 a_1905_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_3599_383.t3 a_1265_943.t6 VPB.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_1905_1004.t6 a_217_1004.t6 VPB.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPB.t4 a_343_383.t7 a_217_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPB.t9 a_217_1004.t7 a_343_383.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 QN a_3599_383.t7 VPB.t23 pshort w=2u l=0.15u
+  ad=1.16p pd=9.16u as=0p ps=0u
M1010 VNB a_217_1004.t10 a_757_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1011 VNB a_1905_1004.t7 a_2702_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPB.t3 CLK a_343_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPB.t19 a_1905_1004.t8 a_1265_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 QN a_343_383.t9 VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 QN a_3599_383.t8 a_3368_73.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1016 VPB.t10 QN a_3599_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPB.t17 a_1265_943.t8 a_3599_383.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 VNB a_217_1004.t5 a_1719_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPB.t21 a_1265_943.t9 a_343_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_217_1004.t1 a_168_157# VPB.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1905_1004.t0 a_1265_943.t10 VPB.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t26 SN a_3599_383.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_217_1004.t3 a_343_383.t10 VPB.t15 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1905_1004.t4 SN VPB.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_343_383.t5 a_217_1004.t8 VPB.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPB.t16 a_217_1004.t9 a_1905_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_343_383.t0 CLK VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1265_943.t4 a_1905_1004.t9 VPB.t29 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPB.t5 a_3599_383.t9 QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 VNB QN a_4013_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPB.t2 CLK a_1265_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_3599_383.t0 QN VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_343_383.t2 a_1265_943.t13 VPB.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPB.t13 a_343_383.t11 QN pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPB.t27 SN a_1905_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1265_943.t0 CLK VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 CLK SN 0.08fF
C1 CLK VPB 0.59fF
C2 a_168_157# VPB 0.08fF
C3 SN QN 0.43fF
C4 SN VPB 0.10fF
C5 VPB QN 1.45fF
R0 VPB VPB.n453 126.832
R1 VPB.n49 VPB.n47 94.117
R2 VPB.n389 VPB.n387 94.117
R3 VPB.n308 VPB.n306 94.117
R4 VPB.n126 VPB.n124 94.117
R5 VPB.n261 VPB.n259 94.117
R6 VPB.n185 VPB.n184 84.554
R7 VPB.n319 VPB.n318 80.104
R8 VPB.n402 VPB.n401 80.104
R9 VPB.n312 VPB.n76 76
R10 VPB.n201 VPB.n200 76
R11 VPB.n206 VPB.n205 76
R12 VPB.n211 VPB.n210 76
R13 VPB.n218 VPB.n217 76
R14 VPB.n223 VPB.n222 76
R15 VPB.n228 VPB.n227 76
R16 VPB.n232 VPB.n231 76
R17 VPB.n236 VPB.n235 76
R18 VPB.n263 VPB.n262 76
R19 VPB.n268 VPB.n267 76
R20 VPB.n273 VPB.n272 76
R21 VPB.n280 VPB.n279 76
R22 VPB.n285 VPB.n284 76
R23 VPB.n290 VPB.n289 76
R24 VPB.n295 VPB.n294 76
R25 VPB.n309 VPB.n305 76
R26 VPB.n317 VPB.n316 76
R27 VPB.n322 VPB.n321 76
R28 VPB.n329 VPB.n328 76
R29 VPB.n334 VPB.n333 76
R30 VPB.n339 VPB.n338 76
R31 VPB.n346 VPB.n345 76
R32 VPB.n351 VPB.n350 76
R33 VPB.n356 VPB.n355 76
R34 VPB.n360 VPB.n359 76
R35 VPB.n364 VPB.n363 76
R36 VPB.n391 VPB.n390 76
R37 VPB.n395 VPB.n394 76
R38 VPB.n400 VPB.n399 76
R39 VPB.n405 VPB.n404 76
R40 VPB.n412 VPB.n411 76
R41 VPB.n417 VPB.n416 76
R42 VPB.n422 VPB.n421 76
R43 VPB.n429 VPB.n428 76
R44 VPB.n434 VPB.n433 76
R45 VPB.n446 VPB.n445 76
R46 VPB.n220 VPB.n219 75.654
R47 VPB.n348 VPB.n347 75.654
R48 VPB.n431 VPB.n430 75.654
R49 VPB.n21 VPB.n20 61.764
R50 VPB.n371 VPB.n370 61.764
R51 VPB.n83 VPB.n82 61.764
R52 VPB.n105 VPB.n104 61.764
R53 VPB.n243 VPB.n242 61.764
R54 VPB.n72 VPB.t7 55.106
R55 VPB.n39 VPB.t14 55.106
R56 VPB.n352 VPB.t20 55.106
R57 VPB.n149 VPB.t29 55.106
R58 VPB.n291 VPB.t12 55.106
R59 VPB.n224 VPB.t11 55.106
R60 VPB.n54 VPB.t4 55.106
R61 VPB.n396 VPB.t21 55.106
R62 VPB.n313 VPB.t22 55.106
R63 VPB.n131 VPB.t2 55.106
R64 VPB.n264 VPB.t5 55.106
R65 VPB.n188 VPB.t17 55.106
R66 VPB.n198 VPB.n197 48.952
R67 VPB.n270 VPB.n269 48.952
R68 VPB.n133 VPB.n132 48.952
R69 VPB.n326 VPB.n325 48.952
R70 VPB.n409 VPB.n408 48.952
R71 VPB.n56 VPB.n55 48.952
R72 VPB.n215 VPB.n214 44.502
R73 VPB.n287 VPB.n286 44.502
R74 VPB.n146 VPB.n145 44.502
R75 VPB.n343 VPB.n342 44.502
R76 VPB.n426 VPB.n425 44.502
R77 VPB.n69 VPB.n68 44.502
R78 VPB.n63 VPB.n14 40.824
R79 VPB.n424 VPB.n423 40.824
R80 VPB.n407 VPB.n406 40.824
R81 VPB.n341 VPB.n340 40.824
R82 VPB.n324 VPB.n323 40.824
R83 VPB.n140 VPB.n98 40.824
R84 VPB.n275 VPB.n274 40.824
R85 VPB.n213 VPB.n212 40.824
R86 VPB.n196 VPB.n195 40.824
R87 VPB.n193 VPB.n192 35.118
R88 VPB.n450 VPB.n446 20.452
R89 VPB.n180 VPB.n177 20.452
R90 VPB.n203 VPB.n202 17.801
R91 VPB.n277 VPB.n276 17.801
R92 VPB.n137 VPB.n136 17.801
R93 VPB.n331 VPB.n330 17.801
R94 VPB.n414 VPB.n413 17.801
R95 VPB.n60 VPB.n59 17.801
R96 VPB.n14 VPB.t15 14.282
R97 VPB.n14 VPB.t6 14.282
R98 VPB.n423 VPB.t0 14.282
R99 VPB.n423 VPB.t9 14.282
R100 VPB.n406 VPB.t28 14.282
R101 VPB.n406 VPB.t3 14.282
R102 VPB.n340 VPB.t25 14.282
R103 VPB.n340 VPB.t16 14.282
R104 VPB.n323 VPB.t8 14.282
R105 VPB.n323 VPB.t27 14.282
R106 VPB.n98 VPB.t1 14.282
R107 VPB.n98 VPB.t19 14.282
R108 VPB.n274 VPB.t23 14.282
R109 VPB.n274 VPB.t13 14.282
R110 VPB.n212 VPB.t24 14.282
R111 VPB.n212 VPB.t10 14.282
R112 VPB.n195 VPB.t18 14.282
R113 VPB.n195 VPB.t26 14.282
R114 VPB.n180 VPB.n179 13.653
R115 VPB.n179 VPB.n178 13.653
R116 VPB.n191 VPB.n190 13.653
R117 VPB.n190 VPB.n189 13.653
R118 VPB.n187 VPB.n186 13.653
R119 VPB.n186 VPB.n185 13.653
R120 VPB.n183 VPB.n182 13.653
R121 VPB.n182 VPB.n181 13.653
R122 VPB.n200 VPB.n199 13.653
R123 VPB.n199 VPB.n198 13.653
R124 VPB.n205 VPB.n204 13.653
R125 VPB.n204 VPB.n203 13.653
R126 VPB.n210 VPB.n209 13.653
R127 VPB.n209 VPB.n208 13.653
R128 VPB.n217 VPB.n216 13.653
R129 VPB.n216 VPB.n215 13.653
R130 VPB.n222 VPB.n221 13.653
R131 VPB.n221 VPB.n220 13.653
R132 VPB.n227 VPB.n226 13.653
R133 VPB.n226 VPB.n225 13.653
R134 VPB.n231 VPB.n230 13.653
R135 VPB.n230 VPB.n229 13.653
R136 VPB.n235 VPB.n234 13.653
R137 VPB.n234 VPB.n233 13.653
R138 VPB.n262 VPB.n261 13.653
R139 VPB.n261 VPB.n260 13.653
R140 VPB.n267 VPB.n266 13.653
R141 VPB.n266 VPB.n265 13.653
R142 VPB.n272 VPB.n271 13.653
R143 VPB.n271 VPB.n270 13.653
R144 VPB.n279 VPB.n278 13.653
R145 VPB.n278 VPB.n277 13.653
R146 VPB.n284 VPB.n283 13.653
R147 VPB.n283 VPB.n282 13.653
R148 VPB.n289 VPB.n288 13.653
R149 VPB.n288 VPB.n287 13.653
R150 VPB.n294 VPB.n293 13.653
R151 VPB.n293 VPB.n292 13.653
R152 VPB.n122 VPB.n121 13.653
R153 VPB.n121 VPB.n120 13.653
R154 VPB.n127 VPB.n126 13.653
R155 VPB.n126 VPB.n125 13.653
R156 VPB.n130 VPB.n129 13.653
R157 VPB.n129 VPB.n128 13.653
R158 VPB.n135 VPB.n134 13.653
R159 VPB.n134 VPB.n133 13.653
R160 VPB.n139 VPB.n138 13.653
R161 VPB.n138 VPB.n137 13.653
R162 VPB.n144 VPB.n143 13.653
R163 VPB.n143 VPB.n142 13.653
R164 VPB.n148 VPB.n147 13.653
R165 VPB.n147 VPB.n146 13.653
R166 VPB.n152 VPB.n151 13.653
R167 VPB.n151 VPB.n150 13.653
R168 VPB.n155 VPB.n154 13.653
R169 VPB.n154 VPB.n153 13.653
R170 VPB.n309 VPB.n308 13.653
R171 VPB.n308 VPB.n307 13.653
R172 VPB.n312 VPB.n311 13.653
R173 VPB.n311 VPB.n310 13.653
R174 VPB.n316 VPB.n315 13.653
R175 VPB.n315 VPB.n314 13.653
R176 VPB.n321 VPB.n320 13.653
R177 VPB.n320 VPB.n319 13.653
R178 VPB.n328 VPB.n327 13.653
R179 VPB.n327 VPB.n326 13.653
R180 VPB.n333 VPB.n332 13.653
R181 VPB.n332 VPB.n331 13.653
R182 VPB.n338 VPB.n337 13.653
R183 VPB.n337 VPB.n336 13.653
R184 VPB.n345 VPB.n344 13.653
R185 VPB.n344 VPB.n343 13.653
R186 VPB.n350 VPB.n349 13.653
R187 VPB.n349 VPB.n348 13.653
R188 VPB.n355 VPB.n354 13.653
R189 VPB.n354 VPB.n353 13.653
R190 VPB.n359 VPB.n358 13.653
R191 VPB.n358 VPB.n357 13.653
R192 VPB.n363 VPB.n362 13.653
R193 VPB.n362 VPB.n361 13.653
R194 VPB.n390 VPB.n389 13.653
R195 VPB.n389 VPB.n388 13.653
R196 VPB.n394 VPB.n393 13.653
R197 VPB.n393 VPB.n392 13.653
R198 VPB.n399 VPB.n398 13.653
R199 VPB.n398 VPB.n397 13.653
R200 VPB.n404 VPB.n403 13.653
R201 VPB.n403 VPB.n402 13.653
R202 VPB.n411 VPB.n410 13.653
R203 VPB.n410 VPB.n409 13.653
R204 VPB.n416 VPB.n415 13.653
R205 VPB.n415 VPB.n414 13.653
R206 VPB.n421 VPB.n420 13.653
R207 VPB.n420 VPB.n419 13.653
R208 VPB.n428 VPB.n427 13.653
R209 VPB.n427 VPB.n426 13.653
R210 VPB.n433 VPB.n432 13.653
R211 VPB.n432 VPB.n431 13.653
R212 VPB.n38 VPB.n37 13.653
R213 VPB.n37 VPB.n36 13.653
R214 VPB.n42 VPB.n41 13.653
R215 VPB.n41 VPB.n40 13.653
R216 VPB.n45 VPB.n44 13.653
R217 VPB.n44 VPB.n43 13.653
R218 VPB.n50 VPB.n49 13.653
R219 VPB.n49 VPB.n48 13.653
R220 VPB.n53 VPB.n52 13.653
R221 VPB.n52 VPB.n51 13.653
R222 VPB.n58 VPB.n57 13.653
R223 VPB.n57 VPB.n56 13.653
R224 VPB.n62 VPB.n61 13.653
R225 VPB.n61 VPB.n60 13.653
R226 VPB.n67 VPB.n66 13.653
R227 VPB.n66 VPB.n65 13.653
R228 VPB.n71 VPB.n70 13.653
R229 VPB.n70 VPB.n69 13.653
R230 VPB.n75 VPB.n74 13.653
R231 VPB.n74 VPB.n73 13.653
R232 VPB.n446 VPB.n0 13.653
R233 VPB VPB.n0 13.653
R234 VPB.n208 VPB.n207 13.35
R235 VPB.n282 VPB.n281 13.35
R236 VPB.n142 VPB.n141 13.35
R237 VPB.n336 VPB.n335 13.35
R238 VPB.n419 VPB.n418 13.35
R239 VPB.n65 VPB.n64 13.35
R240 VPB.n450 VPB.n449 13.276
R241 VPB.n449 VPB.n447 13.276
R242 VPB.n35 VPB.n17 13.276
R243 VPB.n17 VPB.n15 13.276
R244 VPB.n385 VPB.n367 13.276
R245 VPB.n367 VPB.n365 13.276
R246 VPB.n97 VPB.n79 13.276
R247 VPB.n79 VPB.n77 13.276
R248 VPB.n119 VPB.n101 13.276
R249 VPB.n101 VPB.n99 13.276
R250 VPB.n257 VPB.n239 13.276
R251 VPB.n239 VPB.n237 13.276
R252 VPB.n187 VPB.n183 13.276
R253 VPB.n262 VPB.n258 13.276
R254 VPB.n123 VPB.n122 13.276
R255 VPB.n127 VPB.n123 13.276
R256 VPB.n130 VPB.n127 13.276
R257 VPB.n139 VPB.n135 13.276
R258 VPB.n148 VPB.n144 13.276
R259 VPB.n155 VPB.n152 13.276
R260 VPB.n156 VPB.n155 13.276
R261 VPB.n309 VPB.n156 13.276
R262 VPB.n312 VPB.n309 13.276
R263 VPB.n390 VPB.n386 13.276
R264 VPB.n45 VPB.n42 13.276
R265 VPB.n46 VPB.n45 13.276
R266 VPB.n50 VPB.n46 13.276
R267 VPB.n53 VPB.n50 13.276
R268 VPB.n62 VPB.n58 13.276
R269 VPB.n71 VPB.n67 13.276
R270 VPB.n446 VPB.n75 13.276
R271 VPB.n177 VPB.n159 13.276
R272 VPB.n159 VPB.n157 13.276
R273 VPB.n164 VPB.n162 12.796
R274 VPB.n164 VPB.n163 12.564
R275 VPB.n42 VPB.n39 12.558
R276 VPB.n191 VPB.n188 12.2
R277 VPB.n313 VPB.n312 12.2
R278 VPB.n173 VPB.n172 12.198
R279 VPB.n170 VPB.n169 12.198
R280 VPB.n167 VPB.n166 12.198
R281 VPB.n135 VPB.n131 11.841
R282 VPB.n58 VPB.n54 11.841
R283 VPB.n149 VPB.n148 11.482
R284 VPB.n72 VPB.n71 11.482
R285 VPB.n177 VPB.n176 7.5
R286 VPB.n162 VPB.n161 7.5
R287 VPB.n166 VPB.n165 7.5
R288 VPB.n169 VPB.n168 7.5
R289 VPB.n159 VPB.n158 7.5
R290 VPB.n174 VPB.n160 7.5
R291 VPB.n239 VPB.n238 7.5
R292 VPB.n252 VPB.n251 7.5
R293 VPB.n246 VPB.n245 7.5
R294 VPB.n248 VPB.n247 7.5
R295 VPB.n241 VPB.n240 7.5
R296 VPB.n257 VPB.n256 7.5
R297 VPB.n101 VPB.n100 7.5
R298 VPB.n114 VPB.n113 7.5
R299 VPB.n108 VPB.n107 7.5
R300 VPB.n110 VPB.n109 7.5
R301 VPB.n103 VPB.n102 7.5
R302 VPB.n119 VPB.n118 7.5
R303 VPB.n79 VPB.n78 7.5
R304 VPB.n92 VPB.n91 7.5
R305 VPB.n86 VPB.n85 7.5
R306 VPB.n88 VPB.n87 7.5
R307 VPB.n81 VPB.n80 7.5
R308 VPB.n97 VPB.n96 7.5
R309 VPB.n367 VPB.n366 7.5
R310 VPB.n380 VPB.n379 7.5
R311 VPB.n374 VPB.n373 7.5
R312 VPB.n376 VPB.n375 7.5
R313 VPB.n369 VPB.n368 7.5
R314 VPB.n385 VPB.n384 7.5
R315 VPB.n17 VPB.n16 7.5
R316 VPB.n30 VPB.n29 7.5
R317 VPB.n24 VPB.n23 7.5
R318 VPB.n26 VPB.n25 7.5
R319 VPB.n19 VPB.n18 7.5
R320 VPB.n35 VPB.n34 7.5
R321 VPB.n449 VPB.n448 7.5
R322 VPB.n12 VPB.n11 7.5
R323 VPB.n6 VPB.n5 7.5
R324 VPB.n8 VPB.n7 7.5
R325 VPB.n2 VPB.n1 7.5
R326 VPB.n451 VPB.n450 7.5
R327 VPB.n46 VPB.n35 7.176
R328 VPB.n386 VPB.n385 7.176
R329 VPB.n156 VPB.n97 7.176
R330 VPB.n123 VPB.n119 7.176
R331 VPB.n258 VPB.n257 7.176
R332 VPB.n144 VPB.n140 6.817
R333 VPB.n67 VPB.n63 6.817
R334 VPB.n253 VPB.n250 6.729
R335 VPB.n249 VPB.n246 6.729
R336 VPB.n244 VPB.n241 6.729
R337 VPB.n115 VPB.n112 6.729
R338 VPB.n111 VPB.n108 6.729
R339 VPB.n106 VPB.n103 6.729
R340 VPB.n93 VPB.n90 6.729
R341 VPB.n89 VPB.n86 6.729
R342 VPB.n84 VPB.n81 6.729
R343 VPB.n381 VPB.n378 6.729
R344 VPB.n377 VPB.n374 6.729
R345 VPB.n372 VPB.n369 6.729
R346 VPB.n31 VPB.n28 6.729
R347 VPB.n27 VPB.n24 6.729
R348 VPB.n22 VPB.n19 6.729
R349 VPB.n13 VPB.n10 6.729
R350 VPB.n9 VPB.n6 6.729
R351 VPB.n4 VPB.n2 6.729
R352 VPB.n244 VPB.n243 6.728
R353 VPB.n249 VPB.n248 6.728
R354 VPB.n253 VPB.n252 6.728
R355 VPB.n256 VPB.n255 6.728
R356 VPB.n106 VPB.n105 6.728
R357 VPB.n111 VPB.n110 6.728
R358 VPB.n115 VPB.n114 6.728
R359 VPB.n118 VPB.n117 6.728
R360 VPB.n84 VPB.n83 6.728
R361 VPB.n89 VPB.n88 6.728
R362 VPB.n93 VPB.n92 6.728
R363 VPB.n96 VPB.n95 6.728
R364 VPB.n372 VPB.n371 6.728
R365 VPB.n377 VPB.n376 6.728
R366 VPB.n381 VPB.n380 6.728
R367 VPB.n384 VPB.n383 6.728
R368 VPB.n22 VPB.n21 6.728
R369 VPB.n27 VPB.n26 6.728
R370 VPB.n31 VPB.n30 6.728
R371 VPB.n34 VPB.n33 6.728
R372 VPB.n4 VPB.n3 6.728
R373 VPB.n9 VPB.n8 6.728
R374 VPB.n13 VPB.n12 6.728
R375 VPB.n452 VPB.n451 6.728
R376 VPB.n279 VPB.n275 6.458
R377 VPB.n140 VPB.n139 6.458
R378 VPB.n63 VPB.n62 6.458
R379 VPB.n176 VPB.n175 6.398
R380 VPB.n192 VPB.n180 6.112
R381 VPB.n192 VPB.n191 6.101
R382 VPB.n217 VPB.n213 4.305
R383 VPB.n345 VPB.n341 4.305
R384 VPB.n428 VPB.n424 4.305
R385 VPB.n200 VPB.n196 3.947
R386 VPB.n328 VPB.n324 3.947
R387 VPB.n411 VPB.n407 3.947
R388 VPB.n294 VPB.n291 1.794
R389 VPB.n152 VPB.n149 1.794
R390 VPB.n75 VPB.n72 1.794
R391 VPB.n267 VPB.n264 1.435
R392 VPB.n131 VPB.n130 1.435
R393 VPB.n54 VPB.n53 1.435
R394 VPB.n174 VPB.n167 1.402
R395 VPB.n174 VPB.n170 1.402
R396 VPB.n174 VPB.n171 1.402
R397 VPB.n174 VPB.n173 1.402
R398 VPB.n188 VPB.n187 1.076
R399 VPB.n316 VPB.n313 1.076
R400 VPB.n399 VPB.n396 1.076
R401 VPB.n175 VPB.n174 0.735
R402 VPB.n174 VPB.n164 0.735
R403 VPB.n227 VPB.n224 0.717
R404 VPB.n355 VPB.n352 0.717
R405 VPB.n39 VPB.n38 0.717
R406 VPB.n254 VPB.n253 0.387
R407 VPB.n254 VPB.n249 0.387
R408 VPB.n254 VPB.n244 0.387
R409 VPB.n255 VPB.n254 0.387
R410 VPB.n116 VPB.n115 0.387
R411 VPB.n116 VPB.n111 0.387
R412 VPB.n116 VPB.n106 0.387
R413 VPB.n117 VPB.n116 0.387
R414 VPB.n94 VPB.n93 0.387
R415 VPB.n94 VPB.n89 0.387
R416 VPB.n94 VPB.n84 0.387
R417 VPB.n95 VPB.n94 0.387
R418 VPB.n382 VPB.n381 0.387
R419 VPB.n382 VPB.n377 0.387
R420 VPB.n382 VPB.n372 0.387
R421 VPB.n383 VPB.n382 0.387
R422 VPB.n32 VPB.n31 0.387
R423 VPB.n32 VPB.n27 0.387
R424 VPB.n32 VPB.n22 0.387
R425 VPB.n33 VPB.n32 0.387
R426 VPB.n453 VPB.n13 0.387
R427 VPB.n453 VPB.n9 0.387
R428 VPB.n453 VPB.n4 0.387
R429 VPB.n453 VPB.n452 0.387
R430 VPB.n263 VPB.n236 0.272
R431 VPB.n297 VPB.n296 0.272
R432 VPB.n305 VPB.n304 0.272
R433 VPB.n391 VPB.n364 0.272
R434 VPB.n438 VPB.n437 0.272
R435 VPB.n445 VPB 0.198
R436 VPB.n194 VPB.n193 0.136
R437 VPB.n201 VPB.n194 0.136
R438 VPB.n206 VPB.n201 0.136
R439 VPB.n211 VPB.n206 0.136
R440 VPB.n218 VPB.n211 0.136
R441 VPB.n223 VPB.n218 0.136
R442 VPB.n228 VPB.n223 0.136
R443 VPB.n232 VPB.n228 0.136
R444 VPB.n236 VPB.n232 0.136
R445 VPB.n268 VPB.n263 0.136
R446 VPB.n273 VPB.n268 0.136
R447 VPB.n280 VPB.n273 0.136
R448 VPB.n285 VPB.n280 0.136
R449 VPB.n290 VPB.n285 0.136
R450 VPB.n295 VPB.n290 0.136
R451 VPB.n296 VPB.n295 0.136
R452 VPB.n298 VPB.n297 0.136
R453 VPB.n299 VPB.n298 0.136
R454 VPB.n300 VPB.n299 0.136
R455 VPB.n301 VPB.n300 0.136
R456 VPB.n302 VPB.n301 0.136
R457 VPB.n303 VPB.n302 0.136
R458 VPB.n304 VPB.n303 0.136
R459 VPB.n305 VPB.n76 0.136
R460 VPB.n317 VPB.n76 0.136
R461 VPB.n322 VPB.n317 0.136
R462 VPB.n329 VPB.n322 0.136
R463 VPB.n334 VPB.n329 0.136
R464 VPB.n339 VPB.n334 0.136
R465 VPB.n346 VPB.n339 0.136
R466 VPB.n351 VPB.n346 0.136
R467 VPB.n356 VPB.n351 0.136
R468 VPB.n360 VPB.n356 0.136
R469 VPB.n364 VPB.n360 0.136
R470 VPB.n395 VPB.n391 0.136
R471 VPB.n400 VPB.n395 0.136
R472 VPB.n405 VPB.n400 0.136
R473 VPB.n412 VPB.n405 0.136
R474 VPB.n417 VPB.n412 0.136
R475 VPB.n422 VPB.n417 0.136
R476 VPB.n429 VPB.n422 0.136
R477 VPB.n434 VPB.n429 0.136
R478 VPB.n435 VPB.n434 0.136
R479 VPB.n436 VPB.n435 0.136
R480 VPB.n437 VPB.n436 0.136
R481 VPB.n439 VPB.n438 0.136
R482 VPB.n440 VPB.n439 0.136
R483 VPB.n441 VPB.n440 0.136
R484 VPB.n442 VPB.n441 0.136
R485 VPB.n443 VPB.n442 0.136
R486 VPB.n444 VPB.n443 0.136
R487 VPB.n445 VPB.n444 0.136
R488 a_3599_383.n6 a_3599_383.t9 472.359
R489 a_3599_383.n6 a_3599_383.t7 384.527
R490 a_3599_383.n7 a_3599_383.t8 224.666
R491 a_3599_383.n10 a_3599_383.n8 196.598
R492 a_3599_383.n8 a_3599_383.n5 180.846
R493 a_3599_383.n8 a_3599_383.n7 156.035
R494 a_3599_383.n7 a_3599_383.n6 120.107
R495 a_3599_383.n4 a_3599_383.n3 79.232
R496 a_3599_383.n5 a_3599_383.n4 63.152
R497 a_3599_383.n11 a_3599_383.n0 55.263
R498 a_3599_383.n10 a_3599_383.n9 30
R499 a_3599_383.n11 a_3599_383.n10 23.684
R500 a_3599_383.n5 a_3599_383.n1 16.08
R501 a_3599_383.n4 a_3599_383.n2 16.08
R502 a_3599_383.n1 a_3599_383.t2 14.282
R503 a_3599_383.n1 a_3599_383.t3 14.282
R504 a_3599_383.n2 a_3599_383.t5 14.282
R505 a_3599_383.n2 a_3599_383.t6 14.282
R506 a_3599_383.n3 a_3599_383.t1 14.282
R507 a_3599_383.n3 a_3599_383.t0 14.282
R508 a_217_1004.n5 a_217_1004.t7 512.525
R509 a_217_1004.n3 a_217_1004.t9 512.525
R510 a_217_1004.n5 a_217_1004.t8 371.139
R511 a_217_1004.n3 a_217_1004.t6 371.139
R512 a_217_1004.n6 a_217_1004.n5 226.225
R513 a_217_1004.n4 a_217_1004.n3 225.866
R514 a_217_1004.n4 a_217_1004.t5 218.057
R515 a_217_1004.n6 a_217_1004.t10 217.698
R516 a_217_1004.n8 a_217_1004.n2 215.652
R517 a_217_1004.n10 a_217_1004.n8 147.503
R518 a_217_1004.n7 a_217_1004.n4 79.488
R519 a_217_1004.n8 a_217_1004.n7 77.314
R520 a_217_1004.n2 a_217_1004.n1 76.002
R521 a_217_1004.n7 a_217_1004.n6 76
R522 a_217_1004.n10 a_217_1004.n9 15.218
R523 a_217_1004.n0 a_217_1004.t0 14.282
R524 a_217_1004.n0 a_217_1004.t3 14.282
R525 a_217_1004.n1 a_217_1004.t2 14.282
R526 a_217_1004.n1 a_217_1004.t1 14.282
R527 a_217_1004.n2 a_217_1004.n0 12.85
R528 a_217_1004.n11 a_217_1004.n10 12.014
R529 a_1265_943.n6 a_1265_943.t10 454.685
R530 a_1265_943.n8 a_1265_943.t13 454.685
R531 a_1265_943.n4 a_1265_943.t6 454.685
R532 a_1265_943.n6 a_1265_943.t5 428.979
R533 a_1265_943.n8 a_1265_943.t9 428.979
R534 a_1265_943.n4 a_1265_943.t8 428.979
R535 a_1265_943.n7 a_1265_943.t11 248.006
R536 a_1265_943.n9 a_1265_943.t12 248.006
R537 a_1265_943.n5 a_1265_943.t7 248.006
R538 a_1265_943.n14 a_1265_943.n12 220.639
R539 a_1265_943.n12 a_1265_943.n3 135.994
R540 a_1265_943.n7 a_1265_943.n6 81.941
R541 a_1265_943.n9 a_1265_943.n8 81.941
R542 a_1265_943.n5 a_1265_943.n4 81.941
R543 a_1265_943.n11 a_1265_943.n5 81.396
R544 a_1265_943.n10 a_1265_943.n9 79.491
R545 a_1265_943.n3 a_1265_943.n2 76.002
R546 a_1265_943.n10 a_1265_943.n7 76
R547 a_1265_943.n12 a_1265_943.n11 76
R548 a_1265_943.n14 a_1265_943.n13 30
R549 a_1265_943.n15 a_1265_943.n0 24.383
R550 a_1265_943.n15 a_1265_943.n14 23.684
R551 a_1265_943.n1 a_1265_943.t1 14.282
R552 a_1265_943.n1 a_1265_943.t0 14.282
R553 a_1265_943.n2 a_1265_943.t3 14.282
R554 a_1265_943.n2 a_1265_943.t4 14.282
R555 a_1265_943.n3 a_1265_943.n1 12.85
R556 a_1265_943.n11 a_1265_943.n10 2.947
R557 a_1905_1004.n6 a_1905_1004.t8 480.392
R558 a_1905_1004.n6 a_1905_1004.t9 403.272
R559 a_1905_1004.n8 a_1905_1004.n5 233.952
R560 a_1905_1004.n7 a_1905_1004.t7 213.869
R561 a_1905_1004.n7 a_1905_1004.n6 161.6
R562 a_1905_1004.n8 a_1905_1004.n7 153.315
R563 a_1905_1004.n10 a_1905_1004.n8 143.492
R564 a_1905_1004.n4 a_1905_1004.n3 79.232
R565 a_1905_1004.n5 a_1905_1004.n4 63.152
R566 a_1905_1004.n10 a_1905_1004.n9 30
R567 a_1905_1004.n11 a_1905_1004.n0 24.383
R568 a_1905_1004.n11 a_1905_1004.n10 23.684
R569 a_1905_1004.n5 a_1905_1004.n1 16.08
R570 a_1905_1004.n4 a_1905_1004.n2 16.08
R571 a_1905_1004.n1 a_1905_1004.t1 14.282
R572 a_1905_1004.n1 a_1905_1004.t0 14.282
R573 a_1905_1004.n2 a_1905_1004.t3 14.282
R574 a_1905_1004.n2 a_1905_1004.t4 14.282
R575 a_1905_1004.n3 a_1905_1004.t5 14.282
R576 a_1905_1004.n3 a_1905_1004.t6 14.282
R577 a_1719_75.t0 a_1719_75.n0 117.777
R578 a_1719_75.n2 a_1719_75.n1 55.228
R579 a_1719_75.n4 a_1719_75.n3 9.111
R580 a_1719_75.n8 a_1719_75.n6 7.859
R581 a_1719_75.t0 a_1719_75.n2 4.04
R582 a_1719_75.t0 a_1719_75.n8 3.034
R583 a_1719_75.n6 a_1719_75.n4 1.964
R584 a_1719_75.n6 a_1719_75.n5 1.964
R585 a_1719_75.n8 a_1719_75.n7 0.443
R586 VNB VNB.n398 300.778
R587 VNB.n222 VNB.n221 199.897
R588 VNB.n100 VNB.n99 199.897
R589 VNB.n80 VNB.n79 199.897
R590 VNB.n329 VNB.n328 199.897
R591 VNB.n18 VNB.n17 199.897
R592 VNB.n112 VNB.n110 154.509
R593 VNB.n231 VNB.n229 154.509
R594 VNB.n338 VNB.n336 154.509
R595 VNB.n272 VNB.n270 154.509
R596 VNB.n44 VNB.n42 154.509
R597 VNB.n188 VNB.n187 147.75
R598 VNB.n370 VNB.n369 147.75
R599 VNB.n200 VNB.n197 121.366
R600 VNB.n124 VNB.n123 121.366
R601 VNB.n30 VNB.n28 121.366
R602 VNB.n56 VNB.n55 121.366
R603 VNB.n306 VNB.n305 85.559
R604 VNB.n251 VNB.n250 84.842
R605 VNB.n276 VNB.n69 76
R606 VNB.n385 VNB.n384 76
R607 VNB.n373 VNB.n372 76
R608 VNB.n368 VNB.n367 76
R609 VNB.n364 VNB.n363 76
R610 VNB.n360 VNB.n359 76
R611 VNB.n356 VNB.n355 76
R612 VNB.n352 VNB.n351 76
R613 VNB.n348 VNB.n347 76
R614 VNB.n344 VNB.n343 76
R615 VNB.n340 VNB.n339 76
R616 VNB.n318 VNB.n317 76
R617 VNB.n314 VNB.n313 76
R618 VNB.n310 VNB.n309 76
R619 VNB.n304 VNB.n303 76
R620 VNB.n300 VNB.n299 76
R621 VNB.n296 VNB.n295 76
R622 VNB.n292 VNB.n291 76
R623 VNB.n288 VNB.n287 76
R624 VNB.n284 VNB.n283 76
R625 VNB.n280 VNB.n279 76
R626 VNB.n273 VNB.n269 76
R627 VNB.n259 VNB.n258 76
R628 VNB.n255 VNB.n254 76
R629 VNB.n249 VNB.n248 76
R630 VNB.n245 VNB.n244 76
R631 VNB.n241 VNB.n240 76
R632 VNB.n237 VNB.n236 76
R633 VNB.n233 VNB.n232 76
R634 VNB.n211 VNB.n210 76
R635 VNB.n207 VNB.n206 76
R636 VNB.n203 VNB.n202 76
R637 VNB.n191 VNB.n190 76
R638 VNB.n186 VNB.n185 76
R639 VNB.n182 VNB.n181 76
R640 VNB.n178 VNB.n177 76
R641 VNB.n174 VNB.n173 76
R642 VNB.n35 VNB.n34 73.875
R643 VNB.n196 VNB.n195 64.552
R644 VNB.n33 VNB.n27 64.552
R645 VNB.n128 VNB.n89 63.835
R646 VNB.n60 VNB.n7 63.835
R647 VNB.n308 VNB.n307 41.971
R648 VNB.n200 VNB.n199 36.937
R649 VNB.n125 VNB.n124 36.937
R650 VNB.n30 VNB.n29 36.937
R651 VNB.n57 VNB.n56 36.937
R652 VNB.n253 VNB.n252 36.678
R653 VNB.n169 VNB.n168 35.118
R654 VNB.n199 VNB.n198 29.844
R655 VNB.n195 VNB.n194 28.421
R656 VNB.n89 VNB.n88 28.421
R657 VNB.n27 VNB.n26 28.421
R658 VNB.n7 VNB.n6 28.421
R659 VNB.n131 VNB.n130 27.855
R660 VNB.n63 VNB.n62 27.855
R661 VNB.n195 VNB.n193 25.263
R662 VNB.n89 VNB.n87 25.263
R663 VNB.n27 VNB.n25 25.263
R664 VNB.n7 VNB.n5 25.263
R665 VNB.n193 VNB.n192 24.383
R666 VNB.n87 VNB.n86 24.383
R667 VNB.n25 VNB.n24 24.383
R668 VNB.n5 VNB.n4 24.383
R669 VNB.n158 VNB.n155 20.452
R670 VNB.n386 VNB.n385 20.452
R671 VNB.n132 VNB.n131 16.721
R672 VNB.n64 VNB.n63 16.721
R673 VNB.n167 VNB.n166 13.653
R674 VNB.n166 VNB.n165 13.653
R675 VNB.n164 VNB.n163 13.653
R676 VNB.n163 VNB.n162 13.653
R677 VNB.n161 VNB.n160 13.653
R678 VNB.n160 VNB.n159 13.653
R679 VNB.n173 VNB.n172 13.653
R680 VNB.n172 VNB.n171 13.653
R681 VNB.n177 VNB.n176 13.653
R682 VNB.n176 VNB.n175 13.653
R683 VNB.n181 VNB.n180 13.653
R684 VNB.n180 VNB.n179 13.653
R685 VNB.n185 VNB.n184 13.653
R686 VNB.n184 VNB.n183 13.653
R687 VNB.n190 VNB.n189 13.653
R688 VNB.n189 VNB.n188 13.653
R689 VNB.n202 VNB.n201 13.653
R690 VNB.n201 VNB.n200 13.653
R691 VNB.n206 VNB.n205 13.653
R692 VNB.n205 VNB.n204 13.653
R693 VNB.n210 VNB.n209 13.653
R694 VNB.n209 VNB.n208 13.653
R695 VNB.n232 VNB.n231 13.653
R696 VNB.n231 VNB.n230 13.653
R697 VNB.n236 VNB.n235 13.653
R698 VNB.n235 VNB.n234 13.653
R699 VNB.n240 VNB.n239 13.653
R700 VNB.n239 VNB.n238 13.653
R701 VNB.n244 VNB.n243 13.653
R702 VNB.n243 VNB.n242 13.653
R703 VNB.n248 VNB.n247 13.653
R704 VNB.n247 VNB.n246 13.653
R705 VNB.n254 VNB.n253 13.653
R706 VNB.n258 VNB.n257 13.653
R707 VNB.n257 VNB.n256 13.653
R708 VNB.n108 VNB.n107 13.653
R709 VNB.n107 VNB.n106 13.653
R710 VNB.n113 VNB.n112 13.653
R711 VNB.n112 VNB.n111 13.653
R712 VNB.n116 VNB.n115 13.653
R713 VNB.n115 VNB.n114 13.653
R714 VNB.n119 VNB.n118 13.653
R715 VNB.n118 VNB.n117 13.653
R716 VNB.n122 VNB.n121 13.653
R717 VNB.n121 VNB.n120 13.653
R718 VNB.n127 VNB.n126 13.653
R719 VNB.n126 VNB.n125 13.653
R720 VNB.n133 VNB.n132 13.653
R721 VNB.n136 VNB.n135 13.653
R722 VNB.n135 VNB.n134 13.653
R723 VNB.n139 VNB.n138 13.653
R724 VNB.n138 VNB.n137 13.653
R725 VNB.n273 VNB.n272 13.653
R726 VNB.n272 VNB.n271 13.653
R727 VNB.n276 VNB.n275 13.653
R728 VNB.n275 VNB.n274 13.653
R729 VNB.n279 VNB.n278 13.653
R730 VNB.n278 VNB.n277 13.653
R731 VNB.n283 VNB.n282 13.653
R732 VNB.n282 VNB.n281 13.653
R733 VNB.n287 VNB.n286 13.653
R734 VNB.n286 VNB.n285 13.653
R735 VNB.n291 VNB.n290 13.653
R736 VNB.n290 VNB.n289 13.653
R737 VNB.n295 VNB.n294 13.653
R738 VNB.n294 VNB.n293 13.653
R739 VNB.n299 VNB.n298 13.653
R740 VNB.n298 VNB.n297 13.653
R741 VNB.n303 VNB.n302 13.653
R742 VNB.n302 VNB.n301 13.653
R743 VNB.n309 VNB.n308 13.653
R744 VNB.n313 VNB.n312 13.653
R745 VNB.n312 VNB.n311 13.653
R746 VNB.n317 VNB.n316 13.653
R747 VNB.n316 VNB.n315 13.653
R748 VNB.n339 VNB.n338 13.653
R749 VNB.n338 VNB.n337 13.653
R750 VNB.n343 VNB.n342 13.653
R751 VNB.n342 VNB.n341 13.653
R752 VNB.n347 VNB.n346 13.653
R753 VNB.n346 VNB.n345 13.653
R754 VNB.n351 VNB.n350 13.653
R755 VNB.n350 VNB.n349 13.653
R756 VNB.n355 VNB.n354 13.653
R757 VNB.n354 VNB.n353 13.653
R758 VNB.n359 VNB.n358 13.653
R759 VNB.n358 VNB.n357 13.653
R760 VNB.n363 VNB.n362 13.653
R761 VNB.n362 VNB.n361 13.653
R762 VNB.n367 VNB.n366 13.653
R763 VNB.n366 VNB.n365 13.653
R764 VNB.n372 VNB.n371 13.653
R765 VNB.n371 VNB.n370 13.653
R766 VNB.n32 VNB.n31 13.653
R767 VNB.n31 VNB.n30 13.653
R768 VNB.n37 VNB.n36 13.653
R769 VNB.n36 VNB.n35 13.653
R770 VNB.n40 VNB.n39 13.653
R771 VNB.n39 VNB.n38 13.653
R772 VNB.n45 VNB.n44 13.653
R773 VNB.n44 VNB.n43 13.653
R774 VNB.n48 VNB.n47 13.653
R775 VNB.n47 VNB.n46 13.653
R776 VNB.n51 VNB.n50 13.653
R777 VNB.n50 VNB.n49 13.653
R778 VNB.n54 VNB.n53 13.653
R779 VNB.n53 VNB.n52 13.653
R780 VNB.n59 VNB.n58 13.653
R781 VNB.n58 VNB.n57 13.653
R782 VNB.n65 VNB.n64 13.653
R783 VNB.n68 VNB.n67 13.653
R784 VNB.n67 VNB.n66 13.653
R785 VNB.n385 VNB.n0 13.653
R786 VNB VNB.n0 13.653
R787 VNB.n158 VNB.n157 13.653
R788 VNB.n157 VNB.n156 13.653
R789 VNB.n393 VNB.n390 13.577
R790 VNB.n143 VNB.n141 13.276
R791 VNB.n155 VNB.n143 13.276
R792 VNB.n214 VNB.n212 13.276
R793 VNB.n227 VNB.n214 13.276
R794 VNB.n92 VNB.n90 13.276
R795 VNB.n105 VNB.n92 13.276
R796 VNB.n72 VNB.n70 13.276
R797 VNB.n85 VNB.n72 13.276
R798 VNB.n321 VNB.n319 13.276
R799 VNB.n334 VNB.n321 13.276
R800 VNB.n10 VNB.n8 13.276
R801 VNB.n23 VNB.n10 13.276
R802 VNB.n167 VNB.n164 13.276
R803 VNB.n164 VNB.n161 13.276
R804 VNB.n232 VNB.n228 13.276
R805 VNB.n109 VNB.n108 13.276
R806 VNB.n113 VNB.n109 13.276
R807 VNB.n116 VNB.n113 13.276
R808 VNB.n119 VNB.n116 13.276
R809 VNB.n122 VNB.n119 13.276
R810 VNB.n127 VNB.n122 13.276
R811 VNB.n136 VNB.n133 13.276
R812 VNB.n139 VNB.n136 13.276
R813 VNB.n140 VNB.n139 13.276
R814 VNB.n273 VNB.n140 13.276
R815 VNB.n276 VNB.n273 13.276
R816 VNB.n279 VNB.n276 13.276
R817 VNB.n339 VNB.n335 13.276
R818 VNB.n40 VNB.n37 13.276
R819 VNB.n41 VNB.n40 13.276
R820 VNB.n45 VNB.n41 13.276
R821 VNB.n48 VNB.n45 13.276
R822 VNB.n51 VNB.n48 13.276
R823 VNB.n54 VNB.n51 13.276
R824 VNB.n59 VNB.n54 13.276
R825 VNB.n68 VNB.n65 13.276
R826 VNB.n385 VNB.n68 13.276
R827 VNB.n3 VNB.n1 13.276
R828 VNB.n386 VNB.n3 13.276
R829 VNB.n37 VNB.n33 12.02
R830 VNB.n128 VNB.n127 10.764
R831 VNB.n60 VNB.n59 10.764
R832 VNB.n395 VNB.n394 7.5
R833 VNB.n220 VNB.n219 7.5
R834 VNB.n216 VNB.n215 7.5
R835 VNB.n214 VNB.n213 7.5
R836 VNB.n227 VNB.n226 7.5
R837 VNB.n98 VNB.n97 7.5
R838 VNB.n94 VNB.n93 7.5
R839 VNB.n92 VNB.n91 7.5
R840 VNB.n105 VNB.n104 7.5
R841 VNB.n78 VNB.n77 7.5
R842 VNB.n74 VNB.n73 7.5
R843 VNB.n72 VNB.n71 7.5
R844 VNB.n85 VNB.n84 7.5
R845 VNB.n327 VNB.n326 7.5
R846 VNB.n323 VNB.n322 7.5
R847 VNB.n321 VNB.n320 7.5
R848 VNB.n334 VNB.n333 7.5
R849 VNB.n16 VNB.n15 7.5
R850 VNB.n12 VNB.n11 7.5
R851 VNB.n10 VNB.n9 7.5
R852 VNB.n23 VNB.n22 7.5
R853 VNB.n387 VNB.n386 7.5
R854 VNB.n3 VNB.n2 7.5
R855 VNB.n392 VNB.n391 7.5
R856 VNB.n149 VNB.n148 7.5
R857 VNB.n145 VNB.n144 7.5
R858 VNB.n143 VNB.n142 7.5
R859 VNB.n155 VNB.n154 7.5
R860 VNB.n228 VNB.n227 7.176
R861 VNB.n109 VNB.n105 7.176
R862 VNB.n140 VNB.n85 7.176
R863 VNB.n335 VNB.n334 7.176
R864 VNB.n41 VNB.n23 7.176
R865 VNB.n397 VNB.n395 7.011
R866 VNB.n223 VNB.n220 7.011
R867 VNB.n218 VNB.n216 7.011
R868 VNB.n101 VNB.n98 7.011
R869 VNB.n96 VNB.n94 7.011
R870 VNB.n81 VNB.n78 7.011
R871 VNB.n76 VNB.n74 7.011
R872 VNB.n330 VNB.n327 7.011
R873 VNB.n325 VNB.n323 7.011
R874 VNB.n19 VNB.n16 7.011
R875 VNB.n14 VNB.n12 7.011
R876 VNB.n151 VNB.n149 7.011
R877 VNB.n147 VNB.n145 7.011
R878 VNB.n226 VNB.n225 7.01
R879 VNB.n218 VNB.n217 7.01
R880 VNB.n223 VNB.n222 7.01
R881 VNB.n104 VNB.n103 7.01
R882 VNB.n96 VNB.n95 7.01
R883 VNB.n101 VNB.n100 7.01
R884 VNB.n84 VNB.n83 7.01
R885 VNB.n76 VNB.n75 7.01
R886 VNB.n81 VNB.n80 7.01
R887 VNB.n333 VNB.n332 7.01
R888 VNB.n325 VNB.n324 7.01
R889 VNB.n330 VNB.n329 7.01
R890 VNB.n22 VNB.n21 7.01
R891 VNB.n14 VNB.n13 7.01
R892 VNB.n19 VNB.n18 7.01
R893 VNB.n154 VNB.n153 7.01
R894 VNB.n147 VNB.n146 7.01
R895 VNB.n151 VNB.n150 7.01
R896 VNB.n397 VNB.n396 7.01
R897 VNB.n393 VNB.n392 6.788
R898 VNB.n388 VNB.n387 6.788
R899 VNB.n168 VNB.n158 6.111
R900 VNB.n168 VNB.n167 6.1
R901 VNB.n254 VNB.n251 2.511
R902 VNB.n133 VNB.n128 2.511
R903 VNB.n65 VNB.n60 2.511
R904 VNB.n131 VNB.n129 1.99
R905 VNB.n63 VNB.n61 1.99
R906 VNB.n202 VNB.n196 1.255
R907 VNB.n309 VNB.n306 1.255
R908 VNB.n33 VNB.n32 1.255
R909 VNB.n398 VNB.n389 0.921
R910 VNB.n398 VNB.n393 0.476
R911 VNB.n398 VNB.n388 0.475
R912 VNB.n233 VNB.n211 0.272
R913 VNB.n261 VNB.n260 0.272
R914 VNB.n269 VNB.n268 0.272
R915 VNB.n340 VNB.n318 0.272
R916 VNB.n377 VNB.n376 0.272
R917 VNB.n224 VNB.n218 0.246
R918 VNB.n225 VNB.n224 0.246
R919 VNB.n224 VNB.n223 0.246
R920 VNB.n102 VNB.n96 0.246
R921 VNB.n103 VNB.n102 0.246
R922 VNB.n102 VNB.n101 0.246
R923 VNB.n82 VNB.n76 0.246
R924 VNB.n83 VNB.n82 0.246
R925 VNB.n82 VNB.n81 0.246
R926 VNB.n331 VNB.n325 0.246
R927 VNB.n332 VNB.n331 0.246
R928 VNB.n331 VNB.n330 0.246
R929 VNB.n20 VNB.n14 0.246
R930 VNB.n21 VNB.n20 0.246
R931 VNB.n20 VNB.n19 0.246
R932 VNB.n152 VNB.n147 0.246
R933 VNB.n153 VNB.n152 0.246
R934 VNB.n152 VNB.n151 0.246
R935 VNB.n398 VNB.n397 0.246
R936 VNB.n384 VNB 0.198
R937 VNB.n170 VNB.n169 0.136
R938 VNB.n174 VNB.n170 0.136
R939 VNB.n178 VNB.n174 0.136
R940 VNB.n182 VNB.n178 0.136
R941 VNB.n186 VNB.n182 0.136
R942 VNB.n191 VNB.n186 0.136
R943 VNB.n203 VNB.n191 0.136
R944 VNB.n207 VNB.n203 0.136
R945 VNB.n211 VNB.n207 0.136
R946 VNB.n237 VNB.n233 0.136
R947 VNB.n241 VNB.n237 0.136
R948 VNB.n245 VNB.n241 0.136
R949 VNB.n249 VNB.n245 0.136
R950 VNB.n255 VNB.n249 0.136
R951 VNB.n259 VNB.n255 0.136
R952 VNB.n260 VNB.n259 0.136
R953 VNB.n262 VNB.n261 0.136
R954 VNB.n263 VNB.n262 0.136
R955 VNB.n264 VNB.n263 0.136
R956 VNB.n265 VNB.n264 0.136
R957 VNB.n266 VNB.n265 0.136
R958 VNB.n267 VNB.n266 0.136
R959 VNB.n268 VNB.n267 0.136
R960 VNB.n269 VNB.n69 0.136
R961 VNB.n280 VNB.n69 0.136
R962 VNB.n284 VNB.n280 0.136
R963 VNB.n288 VNB.n284 0.136
R964 VNB.n292 VNB.n288 0.136
R965 VNB.n296 VNB.n292 0.136
R966 VNB.n300 VNB.n296 0.136
R967 VNB.n304 VNB.n300 0.136
R968 VNB.n310 VNB.n304 0.136
R969 VNB.n314 VNB.n310 0.136
R970 VNB.n318 VNB.n314 0.136
R971 VNB.n344 VNB.n340 0.136
R972 VNB.n348 VNB.n344 0.136
R973 VNB.n352 VNB.n348 0.136
R974 VNB.n356 VNB.n352 0.136
R975 VNB.n360 VNB.n356 0.136
R976 VNB.n364 VNB.n360 0.136
R977 VNB.n368 VNB.n364 0.136
R978 VNB.n373 VNB.n368 0.136
R979 VNB.n374 VNB.n373 0.136
R980 VNB.n375 VNB.n374 0.136
R981 VNB.n376 VNB.n375 0.136
R982 VNB.n378 VNB.n377 0.136
R983 VNB.n379 VNB.n378 0.136
R984 VNB.n380 VNB.n379 0.136
R985 VNB.n381 VNB.n380 0.136
R986 VNB.n382 VNB.n381 0.136
R987 VNB.n383 VNB.n382 0.136
R988 VNB.n384 VNB.n383 0.136
R989 a_757_75.n1 a_757_75.n0 25.576
R990 a_757_75.n3 a_757_75.n2 9.111
R991 a_757_75.n7 a_757_75.n5 7.859
R992 a_757_75.t0 a_757_75.n7 3.034
R993 a_757_75.n5 a_757_75.n3 1.964
R994 a_757_75.n5 a_757_75.n4 1.964
R995 a_757_75.t0 a_757_75.n1 1.871
R996 a_757_75.n7 a_757_75.n6 0.443
R997 a_1038_182.n12 a_1038_182.n10 82.852
R998 a_1038_182.n13 a_1038_182.n0 49.6
R999 a_1038_182.t1 a_1038_182.n2 46.91
R1000 a_1038_182.n7 a_1038_182.n5 34.805
R1001 a_1038_182.n7 a_1038_182.n6 32.622
R1002 a_1038_182.n10 a_1038_182.t1 32.416
R1003 a_1038_182.n12 a_1038_182.n11 27.2
R1004 a_1038_182.n13 a_1038_182.n12 22.4
R1005 a_1038_182.n9 a_1038_182.n7 19.017
R1006 a_1038_182.n2 a_1038_182.n1 17.006
R1007 a_1038_182.n5 a_1038_182.n4 7.5
R1008 a_1038_182.n9 a_1038_182.n8 7.5
R1009 a_1038_182.t1 a_1038_182.n3 7.04
R1010 a_1038_182.n10 a_1038_182.n9 1.435
R1011 a_343_383.n6 a_343_383.t11 480.392
R1012 a_343_383.n8 a_343_383.t7 472.359
R1013 a_343_383.n6 a_343_383.t9 403.272
R1014 a_343_383.n8 a_343_383.t10 384.527
R1015 a_343_383.n7 a_343_383.t12 320.08
R1016 a_343_383.n9 a_343_383.t8 277.772
R1017 a_343_383.n13 a_343_383.n11 249.364
R1018 a_343_383.n11 a_343_383.n5 127.401
R1019 a_343_383.n10 a_343_383.n7 83.304
R1020 a_343_383.n10 a_343_383.n9 80.032
R1021 a_343_383.n4 a_343_383.n3 79.232
R1022 a_343_383.n11 a_343_383.n10 76
R1023 a_343_383.n9 a_343_383.n8 67.001
R1024 a_343_383.n5 a_343_383.n4 63.152
R1025 a_343_383.n7 a_343_383.n6 55.388
R1026 a_343_383.n14 a_343_383.n0 55.263
R1027 a_343_383.n13 a_343_383.n12 30
R1028 a_343_383.n14 a_343_383.n13 23.684
R1029 a_343_383.n5 a_343_383.n1 16.08
R1030 a_343_383.n4 a_343_383.n2 16.08
R1031 a_343_383.n1 a_343_383.t3 14.282
R1032 a_343_383.n1 a_343_383.t2 14.282
R1033 a_343_383.n2 a_343_383.t1 14.282
R1034 a_343_383.n2 a_343_383.t0 14.282
R1035 a_343_383.n3 a_343_383.t6 14.282
R1036 a_343_383.n3 a_343_383.t5 14.282
R1037 a_2702_73.t0 a_2702_73.n1 34.62
R1038 a_2702_73.t0 a_2702_73.n0 8.137
R1039 a_2702_73.t0 a_2702_73.n2 4.69
R1040 a_112_73.n12 a_112_73.n11 26.811
R1041 a_112_73.n6 a_112_73.n5 24.977
R1042 a_112_73.n2 a_112_73.n1 24.877
R1043 a_112_73.t0 a_112_73.n2 12.677
R1044 a_112_73.t0 a_112_73.n3 11.595
R1045 a_112_73.t1 a_112_73.n8 8.137
R1046 a_112_73.t0 a_112_73.n4 7.273
R1047 a_112_73.t0 a_112_73.n0 6.109
R1048 a_112_73.t1 a_112_73.n7 4.864
R1049 a_112_73.t0 a_112_73.n12 2.074
R1050 a_112_73.n7 a_112_73.n6 1.13
R1051 a_112_73.n12 a_112_73.t1 0.937
R1052 a_112_73.t1 a_112_73.n10 0.804
R1053 a_112_73.n10 a_112_73.n9 0.136
R1054 a_4294_182.n9 a_4294_182.n7 82.852
R1055 a_4294_182.n3 a_4294_182.n1 44.628
R1056 a_4294_182.t0 a_4294_182.n9 32.417
R1057 a_4294_182.n7 a_4294_182.n6 27.2
R1058 a_4294_182.n5 a_4294_182.n4 23.498
R1059 a_4294_182.n3 a_4294_182.n2 23.284
R1060 a_4294_182.n7 a_4294_182.n5 22.4
R1061 a_4294_182.t0 a_4294_182.n11 20.241
R1062 a_4294_182.n11 a_4294_182.n10 13.494
R1063 a_4294_182.t0 a_4294_182.n0 8.137
R1064 a_4294_182.t0 a_4294_182.n3 5.727
R1065 a_4294_182.n9 a_4294_182.n8 1.435
R1066 a_2000_182.n8 a_2000_182.n6 96.467
R1067 a_2000_182.n3 a_2000_182.n1 44.628
R1068 a_2000_182.t0 a_2000_182.n8 32.417
R1069 a_2000_182.n3 a_2000_182.n2 23.284
R1070 a_2000_182.n6 a_2000_182.n5 22.349
R1071 a_2000_182.t0 a_2000_182.n10 20.241
R1072 a_2000_182.n10 a_2000_182.n9 13.494
R1073 a_2000_182.n6 a_2000_182.n4 8.443
R1074 a_2000_182.t0 a_2000_182.n0 8.137
R1075 a_2000_182.t0 a_2000_182.n3 5.727
R1076 a_2000_182.n8 a_2000_182.n7 1.435
R1077 a_3368_73.t0 a_3368_73.n1 34.62
R1078 a_3368_73.t0 a_3368_73.n0 8.137
R1079 a_3368_73.t0 a_3368_73.n2 4.69
R1080 a_4013_75.n5 a_4013_75.n4 19.724
R1081 a_4013_75.t0 a_4013_75.n3 11.595
R1082 a_4013_75.t0 a_4013_75.n5 9.207
R1083 a_4013_75.n2 a_4013_75.n1 2.455
R1084 a_4013_75.n2 a_4013_75.n0 1.32
R1085 a_4013_75.t0 a_4013_75.n2 0.246
C6 VPB VNB 19.03fF
C7 a_4013_75.n0 VNB 0.10fF
C8 a_4013_75.n1 VNB 0.04fF
C9 a_4013_75.n2 VNB 0.03fF
C10 a_4013_75.n3 VNB 0.07fF
C11 a_4013_75.n4 VNB 0.08fF
C12 a_4013_75.n5 VNB 0.06fF
C13 a_3368_73.n0 VNB 0.05fF
C14 a_3368_73.n1 VNB 0.12fF
C15 a_3368_73.n2 VNB 0.04fF
C16 a_2000_182.n0 VNB 0.07fF
C17 a_2000_182.n1 VNB 0.09fF
C18 a_2000_182.n2 VNB 0.13fF
C19 a_2000_182.n3 VNB 0.11fF
C20 a_2000_182.n4 VNB 0.02fF
C21 a_2000_182.n5 VNB 0.03fF
C22 a_2000_182.n6 VNB 0.06fF
C23 a_2000_182.n7 VNB 0.03fF
C24 a_2000_182.n8 VNB 0.12fF
C25 a_2000_182.n9 VNB 0.06fF
C26 a_2000_182.n10 VNB 0.01fF
C27 a_2000_182.t0 VNB 0.33fF
C28 a_4294_182.n0 VNB 0.07fF
C29 a_4294_182.n1 VNB 0.09fF
C30 a_4294_182.n2 VNB 0.13fF
C31 a_4294_182.n3 VNB 0.11fF
C32 a_4294_182.n4 VNB 0.02fF
C33 a_4294_182.n5 VNB 0.03fF
C34 a_4294_182.n6 VNB 0.02fF
C35 a_4294_182.n7 VNB 0.05fF
C36 a_4294_182.n8 VNB 0.03fF
C37 a_4294_182.n9 VNB 0.11fF
C38 a_4294_182.n10 VNB 0.05fF
C39 a_4294_182.n11 VNB 0.01fF
C40 a_4294_182.t0 VNB 0.32fF
C41 a_112_73.n0 VNB 0.02fF
C42 a_112_73.n1 VNB 0.10fF
C43 a_112_73.n2 VNB 0.06fF
C44 a_112_73.n3 VNB 0.06fF
C45 a_112_73.n4 VNB 0.00fF
C46 a_112_73.n5 VNB 0.04fF
C47 a_112_73.n6 VNB 0.05fF
C48 a_112_73.n7 VNB 0.02fF
C49 a_112_73.n8 VNB 0.05fF
C50 a_112_73.n9 VNB 0.07fF
C51 a_112_73.n10 VNB 0.17fF
C52 a_112_73.t1 VNB 0.22fF
C53 a_112_73.n11 VNB 0.09fF
C54 a_112_73.n12 VNB 0.00fF
C55 a_2702_73.n0 VNB 0.05fF
C56 a_2702_73.n1 VNB 0.12fF
C57 a_2702_73.n2 VNB 0.04fF
C58 a_343_383.n0 VNB 0.05fF
C59 a_343_383.n1 VNB 0.68fF
C60 a_343_383.n2 VNB 0.68fF
C61 a_343_383.n3 VNB 0.80fF
C62 a_343_383.n4 VNB 0.25fF
C63 a_343_383.n5 VNB 0.32fF
C64 a_343_383.n6 VNB 0.41fF
C65 a_343_383.n7 VNB 0.59fF
C66 a_343_383.n8 VNB 0.36fF
C67 a_343_383.t8 VNB 0.72fF
C68 a_343_383.n9 VNB 0.50fF
C69 a_343_383.n10 VNB 3.16fF
C70 a_343_383.n11 VNB 0.56fF
C71 a_343_383.n12 VNB 0.05fF
C72 a_343_383.n13 VNB 0.43fF
C73 a_343_383.n14 VNB 0.06fF
C74 a_1038_182.n0 VNB 0.02fF
C75 a_1038_182.n1 VNB 0.07fF
C76 a_1038_182.n2 VNB 0.13fF
C77 a_1038_182.n3 VNB 0.09fF
C78 a_1038_182.t1 VNB 0.25fF
C79 a_1038_182.n4 VNB 0.05fF
C80 a_1038_182.n5 VNB 0.06fF
C81 a_1038_182.n6 VNB 0.07fF
C82 a_1038_182.n7 VNB 0.07fF
C83 a_1038_182.n8 VNB 0.03fF
C84 a_1038_182.n9 VNB 0.01fF
C85 a_1038_182.n10 VNB 0.11fF
C86 a_1038_182.n11 VNB 0.02fF
C87 a_1038_182.n12 VNB 0.05fF
C88 a_1038_182.n13 VNB 0.02fF
C89 a_757_75.n0 VNB 0.09fF
C90 a_757_75.n1 VNB 0.10fF
C91 a_757_75.n2 VNB 0.05fF
C92 a_757_75.n3 VNB 0.03fF
C93 a_757_75.n4 VNB 0.04fF
C94 a_757_75.n5 VNB 0.11fF
C95 a_757_75.n6 VNB 0.04fF
C96 a_1719_75.n0 VNB 0.03fF
C97 a_1719_75.n1 VNB 0.10fF
C98 a_1719_75.n2 VNB 0.10fF
C99 a_1719_75.n3 VNB 0.05fF
C100 a_1719_75.n4 VNB 0.03fF
C101 a_1719_75.n5 VNB 0.04fF
C102 a_1719_75.n6 VNB 0.11fF
C103 a_1719_75.n7 VNB 0.04fF
C104 a_1905_1004.n0 VNB 0.04fF
C105 a_1905_1004.n1 VNB 0.48fF
C106 a_1905_1004.n2 VNB 0.48fF
C107 a_1905_1004.n3 VNB 0.57fF
C108 a_1905_1004.n4 VNB 0.18fF
C109 a_1905_1004.n5 VNB 0.34fF
C110 a_1905_1004.n6 VNB 0.40fF
C111 a_1905_1004.n7 VNB 0.49fF
C112 a_1905_1004.n8 VNB 0.56fF
C113 a_1905_1004.n9 VNB 0.03fF
C114 a_1905_1004.n10 VNB 0.20fF
C115 a_1905_1004.n11 VNB 0.05fF
C116 a_1265_943.n0 VNB 0.05fF
C117 a_1265_943.n1 VNB 0.65fF
C118 a_1265_943.n2 VNB 0.76fF
C119 a_1265_943.n3 VNB 0.35fF
C120 a_1265_943.n4 VNB 0.43fF
C121 a_1265_943.t7 VNB 0.66fF
C122 a_1265_943.n5 VNB 0.49fF
C123 a_1265_943.n6 VNB 0.43fF
C124 a_1265_943.t11 VNB 0.66fF
C125 a_1265_943.n7 VNB 0.44fF
C126 a_1265_943.n8 VNB 0.43fF
C127 a_1265_943.t12 VNB 0.66fF
C128 a_1265_943.n9 VNB 0.46fF
C129 a_1265_943.n10 VNB 1.39fF
C130 a_1265_943.n11 VNB 1.87fF
C131 a_1265_943.n12 VNB 0.51fF
C132 a_1265_943.n13 VNB 0.04fF
C133 a_1265_943.n14 VNB 0.38fF
C134 a_1265_943.n15 VNB 0.07fF
C135 a_217_1004.n0 VNB 0.42fF
C136 a_217_1004.n1 VNB 0.50fF
C137 a_217_1004.n2 VNB 0.30fF
C138 a_217_1004.n3 VNB 0.33fF
C139 a_217_1004.n4 VNB 0.38fF
C140 a_217_1004.n5 VNB 0.33fF
C141 a_217_1004.n6 VNB 0.36fF
C142 a_217_1004.n7 VNB 0.90fF
C143 a_217_1004.n8 VNB 0.34fF
C144 a_217_1004.n9 VNB 0.07fF
C145 a_217_1004.n10 VNB 0.16fF
C146 a_217_1004.n11 VNB 0.04fF
C147 a_3599_383.n0 VNB 0.04fF
C148 a_3599_383.n1 VNB 0.55fF
C149 a_3599_383.n2 VNB 0.55fF
C150 a_3599_383.n3 VNB 0.65fF
C151 a_3599_383.n4 VNB 0.20fF
C152 a_3599_383.n5 VNB 0.33fF
C153 a_3599_383.n6 VNB 0.36fF
C154 a_3599_383.n7 VNB 0.87fF
C155 a_3599_383.n8 VNB 0.95fF
C156 a_3599_383.n9 VNB 0.04fF
C157 a_3599_383.n10 VNB 0.29fF
C158 a_3599_383.n11 VNB 0.05fF
C159 VPB.n0 VNB 0.03fF
C160 VPB.n1 VNB 0.04fF
C161 VPB.n2 VNB 0.02fF
C162 VPB.n3 VNB 0.14fF
C163 VPB.n5 VNB 0.02fF
C164 VPB.n6 VNB 0.02fF
C165 VPB.n7 VNB 0.02fF
C166 VPB.n8 VNB 0.02fF
C167 VPB.n10 VNB 0.02fF
C168 VPB.n11 VNB 0.02fF
C169 VPB.n12 VNB 0.02fF
C170 VPB.n14 VNB 0.10fF
C171 VPB.n15 VNB 0.02fF
C172 VPB.n16 VNB 0.02fF
C173 VPB.n17 VNB 0.02fF
C174 VPB.n18 VNB 0.04fF
C175 VPB.n19 VNB 0.02fF
C176 VPB.n20 VNB 0.24fF
C177 VPB.n21 VNB 0.04fF
C178 VPB.n23 VNB 0.02fF
C179 VPB.n24 VNB 0.02fF
C180 VPB.n25 VNB 0.02fF
C181 VPB.n26 VNB 0.02fF
C182 VPB.n28 VNB 0.02fF
C183 VPB.n29 VNB 0.02fF
C184 VPB.n30 VNB 0.02fF
C185 VPB.n32 VNB 0.27fF
C186 VPB.n34 VNB 0.03fF
C187 VPB.n35 VNB 0.02fF
C188 VPB.n36 VNB 0.21fF
C189 VPB.n37 VNB 0.02fF
C190 VPB.n38 VNB 0.01fF
C191 VPB.n39 VNB 0.06fF
C192 VPB.n40 VNB 0.27fF
C193 VPB.n41 VNB 0.02fF
C194 VPB.n42 VNB 0.02fF
C195 VPB.n43 VNB 0.27fF
C196 VPB.n44 VNB 0.01fF
C197 VPB.n45 VNB 0.02fF
C198 VPB.n46 VNB 0.03fF
C199 VPB.n47 VNB 0.03fF
C200 VPB.n48 VNB 0.27fF
C201 VPB.n49 VNB 0.01fF
C202 VPB.n50 VNB 0.02fF
C203 VPB.n51 VNB 0.23fF
C204 VPB.n52 VNB 0.02fF
C205 VPB.n53 VNB 0.01fF
C206 VPB.n54 VNB 0.05fF
C207 VPB.n55 VNB 0.13fF
C208 VPB.n56 VNB 0.16fF
C209 VPB.n57 VNB 0.02fF
C210 VPB.n58 VNB 0.02fF
C211 VPB.n59 VNB 0.13fF
C212 VPB.n60 VNB 0.15fF
C213 VPB.n61 VNB 0.02fF
C214 VPB.n62 VNB 0.02fF
C215 VPB.n63 VNB 0.02fF
C216 VPB.n64 VNB 0.13fF
C217 VPB.n65 VNB 0.14fF
C218 VPB.n66 VNB 0.02fF
C219 VPB.n67 VNB 0.02fF
C220 VPB.n68 VNB 0.13fF
C221 VPB.n69 VNB 0.16fF
C222 VPB.n70 VNB 0.02fF
C223 VPB.n71 VNB 0.02fF
C224 VPB.n72 VNB 0.06fF
C225 VPB.n73 VNB 0.23fF
C226 VPB.n74 VNB 0.02fF
C227 VPB.n75 VNB 0.01fF
C228 VPB.n76 VNB 0.02fF
C229 VPB.n77 VNB 0.02fF
C230 VPB.n78 VNB 0.02fF
C231 VPB.n79 VNB 0.02fF
C232 VPB.n80 VNB 0.04fF
C233 VPB.n81 VNB 0.02fF
C234 VPB.n82 VNB 0.23fF
C235 VPB.n83 VNB 0.04fF
C236 VPB.n85 VNB 0.02fF
C237 VPB.n86 VNB 0.02fF
C238 VPB.n87 VNB 0.02fF
C239 VPB.n88 VNB 0.02fF
C240 VPB.n90 VNB 0.02fF
C241 VPB.n91 VNB 0.02fF
C242 VPB.n92 VNB 0.02fF
C243 VPB.n94 VNB 0.27fF
C244 VPB.n96 VNB 0.03fF
C245 VPB.n97 VNB 0.02fF
C246 VPB.n98 VNB 0.10fF
C247 VPB.n99 VNB 0.02fF
C248 VPB.n100 VNB 0.02fF
C249 VPB.n101 VNB 0.02fF
C250 VPB.n102 VNB 0.04fF
C251 VPB.n103 VNB 0.02fF
C252 VPB.n104 VNB 0.19fF
C253 VPB.n105 VNB 0.04fF
C254 VPB.n107 VNB 0.02fF
C255 VPB.n108 VNB 0.02fF
C256 VPB.n109 VNB 0.02fF
C257 VPB.n110 VNB 0.02fF
C258 VPB.n112 VNB 0.02fF
C259 VPB.n113 VNB 0.02fF
C260 VPB.n114 VNB 0.02fF
C261 VPB.n116 VNB 0.27fF
C262 VPB.n118 VNB 0.03fF
C263 VPB.n119 VNB 0.02fF
C264 VPB.n120 VNB 0.27fF
C265 VPB.n121 VNB 0.01fF
C266 VPB.n122 VNB 0.02fF
C267 VPB.n123 VNB 0.03fF
C268 VPB.n124 VNB 0.03fF
C269 VPB.n125 VNB 0.27fF
C270 VPB.n126 VNB 0.01fF
C271 VPB.n127 VNB 0.02fF
C272 VPB.n128 VNB 0.23fF
C273 VPB.n129 VNB 0.02fF
C274 VPB.n130 VNB 0.01fF
C275 VPB.n131 VNB 0.05fF
C276 VPB.n132 VNB 0.13fF
C277 VPB.n133 VNB 0.16fF
C278 VPB.n134 VNB 0.02fF
C279 VPB.n135 VNB 0.02fF
C280 VPB.n136 VNB 0.13fF
C281 VPB.n137 VNB 0.15fF
C282 VPB.n138 VNB 0.02fF
C283 VPB.n139 VNB 0.02fF
C284 VPB.n140 VNB 0.02fF
C285 VPB.n141 VNB 0.13fF
C286 VPB.n142 VNB 0.14fF
C287 VPB.n143 VNB 0.02fF
C288 VPB.n144 VNB 0.02fF
C289 VPB.n145 VNB 0.13fF
C290 VPB.n146 VNB 0.16fF
C291 VPB.n147 VNB 0.02fF
C292 VPB.n148 VNB 0.02fF
C293 VPB.n149 VNB 0.06fF
C294 VPB.n150 VNB 0.23fF
C295 VPB.n151 VNB 0.02fF
C296 VPB.n152 VNB 0.01fF
C297 VPB.n153 VNB 0.27fF
C298 VPB.n154 VNB 0.01fF
C299 VPB.n155 VNB 0.02fF
C300 VPB.n156 VNB 0.03fF
C301 VPB.n157 VNB 0.02fF
C302 VPB.n158 VNB 0.02fF
C303 VPB.n159 VNB 0.02fF
C304 VPB.n160 VNB 0.18fF
C305 VPB.n161 VNB 0.03fF
C306 VPB.n162 VNB 0.02fF
C307 VPB.n163 VNB 0.05fF
C308 VPB.n164 VNB 0.01fF
C309 VPB.n165 VNB 0.02fF
C310 VPB.n166 VNB 0.02fF
C311 VPB.n168 VNB 0.02fF
C312 VPB.n169 VNB 0.02fF
C313 VPB.n172 VNB 0.02fF
C314 VPB.n174 VNB 0.45fF
C315 VPB.n176 VNB 0.04fF
C316 VPB.n177 VNB 0.04fF
C317 VPB.n178 VNB 0.27fF
C318 VPB.n179 VNB 0.03fF
C319 VPB.n180 VNB 0.03fF
C320 VPB.n181 VNB 0.16fF
C321 VPB.n182 VNB 0.02fF
C322 VPB.n183 VNB 0.02fF
C323 VPB.n184 VNB 0.13fF
C324 VPB.n185 VNB 0.20fF
C325 VPB.n186 VNB 0.02fF
C326 VPB.n187 VNB 0.01fF
C327 VPB.n188 VNB 0.05fF
C328 VPB.n189 VNB 0.27fF
C329 VPB.n190 VNB 0.02fF
C330 VPB.n191 VNB 0.02fF
C331 VPB.n192 VNB 0.00fF
C332 VPB.n193 VNB 0.09fF
C333 VPB.n194 VNB 0.02fF
C334 VPB.n195 VNB 0.10fF
C335 VPB.n196 VNB 0.02fF
C336 VPB.n197 VNB 0.13fF
C337 VPB.n198 VNB 0.16fF
C338 VPB.n199 VNB 0.02fF
C339 VPB.n200 VNB 0.02fF
C340 VPB.n201 VNB 0.02fF
C341 VPB.n202 VNB 0.13fF
C342 VPB.n203 VNB 0.15fF
C343 VPB.n204 VNB 0.02fF
C344 VPB.n205 VNB 0.02fF
C345 VPB.n206 VNB 0.02fF
C346 VPB.n207 VNB 0.13fF
C347 VPB.n208 VNB 0.14fF
C348 VPB.n209 VNB 0.02fF
C349 VPB.n210 VNB 0.02fF
C350 VPB.n211 VNB 0.02fF
C351 VPB.n212 VNB 0.10fF
C352 VPB.n213 VNB 0.02fF
C353 VPB.n214 VNB 0.13fF
C354 VPB.n215 VNB 0.16fF
C355 VPB.n216 VNB 0.02fF
C356 VPB.n217 VNB 0.02fF
C357 VPB.n218 VNB 0.02fF
C358 VPB.n219 VNB 0.13fF
C359 VPB.n220 VNB 0.16fF
C360 VPB.n221 VNB 0.02fF
C361 VPB.n222 VNB 0.02fF
C362 VPB.n223 VNB 0.02fF
C363 VPB.n224 VNB 0.06fF
C364 VPB.n225 VNB 0.21fF
C365 VPB.n226 VNB 0.02fF
C366 VPB.n227 VNB 0.01fF
C367 VPB.n228 VNB 0.02fF
C368 VPB.n229 VNB 0.27fF
C369 VPB.n230 VNB 0.02fF
C370 VPB.n231 VNB 0.02fF
C371 VPB.n232 VNB 0.02fF
C372 VPB.n233 VNB 0.27fF
C373 VPB.n234 VNB 0.01fF
C374 VPB.n235 VNB 0.02fF
C375 VPB.n236 VNB 0.04fF
C376 VPB.n237 VNB 0.02fF
C377 VPB.n238 VNB 0.02fF
C378 VPB.n239 VNB 0.02fF
C379 VPB.n240 VNB 0.04fF
C380 VPB.n241 VNB 0.02fF
C381 VPB.n242 VNB 0.24fF
C382 VPB.n243 VNB 0.04fF
C383 VPB.n245 VNB 0.02fF
C384 VPB.n246 VNB 0.02fF
C385 VPB.n247 VNB 0.02fF
C386 VPB.n248 VNB 0.02fF
C387 VPB.n250 VNB 0.02fF
C388 VPB.n251 VNB 0.02fF
C389 VPB.n252 VNB 0.02fF
C390 VPB.n254 VNB 0.27fF
C391 VPB.n256 VNB 0.03fF
C392 VPB.n257 VNB 0.02fF
C393 VPB.n258 VNB 0.03fF
C394 VPB.n259 VNB 0.03fF
C395 VPB.n260 VNB 0.27fF
C396 VPB.n261 VNB 0.01fF
C397 VPB.n262 VNB 0.02fF
C398 VPB.n263 VNB 0.04fF
C399 VPB.n264 VNB 0.05fF
C400 VPB.n265 VNB 0.23fF
C401 VPB.n266 VNB 0.02fF
C402 VPB.n267 VNB 0.01fF
C403 VPB.n268 VNB 0.02fF
C404 VPB.n269 VNB 0.13fF
C405 VPB.n270 VNB 0.16fF
C406 VPB.n271 VNB 0.02fF
C407 VPB.n272 VNB 0.02fF
C408 VPB.n273 VNB 0.02fF
C409 VPB.n274 VNB 0.10fF
C410 VPB.n275 VNB 0.02fF
C411 VPB.n276 VNB 0.13fF
C412 VPB.n277 VNB 0.15fF
C413 VPB.n278 VNB 0.02fF
C414 VPB.n279 VNB 0.02fF
C415 VPB.n280 VNB 0.02fF
C416 VPB.n281 VNB 0.13fF
C417 VPB.n282 VNB 0.14fF
C418 VPB.n283 VNB 0.02fF
C419 VPB.n284 VNB 0.02fF
C420 VPB.n285 VNB 0.02fF
C421 VPB.n286 VNB 0.13fF
C422 VPB.n287 VNB 0.16fF
C423 VPB.n288 VNB 0.02fF
C424 VPB.n289 VNB 0.02fF
C425 VPB.n290 VNB 0.02fF
C426 VPB.n291 VNB 0.06fF
C427 VPB.n292 VNB 0.23fF
C428 VPB.n293 VNB 0.02fF
C429 VPB.n294 VNB 0.01fF
C430 VPB.n295 VNB 0.02fF
C431 VPB.n296 VNB 0.04fF
C432 VPB.n297 VNB 0.04fF
C433 VPB.n298 VNB 0.02fF
C434 VPB.n299 VNB 0.02fF
C435 VPB.n300 VNB 0.02fF
C436 VPB.n301 VNB 0.02fF
C437 VPB.n302 VNB 0.02fF
C438 VPB.n303 VNB 0.02fF
C439 VPB.n304 VNB 0.04fF
C440 VPB.n305 VNB 0.04fF
C441 VPB.n306 VNB 0.03fF
C442 VPB.n307 VNB 0.27fF
C443 VPB.n308 VNB 0.01fF
C444 VPB.n309 VNB 0.02fF
C445 VPB.n310 VNB 0.27fF
C446 VPB.n311 VNB 0.02fF
C447 VPB.n312 VNB 0.02fF
C448 VPB.n313 VNB 0.05fF
C449 VPB.n314 VNB 0.20fF
C450 VPB.n315 VNB 0.02fF
C451 VPB.n316 VNB 0.01fF
C452 VPB.n317 VNB 0.02fF
C453 VPB.n318 VNB 0.13fF
C454 VPB.n319 VNB 0.16fF
C455 VPB.n320 VNB 0.02fF
C456 VPB.n321 VNB 0.02fF
C457 VPB.n322 VNB 0.02fF
C458 VPB.n323 VNB 0.10fF
C459 VPB.n324 VNB 0.02fF
C460 VPB.n325 VNB 0.13fF
C461 VPB.n326 VNB 0.16fF
C462 VPB.n327 VNB 0.02fF
C463 VPB.n328 VNB 0.02fF
C464 VPB.n329 VNB 0.02fF
C465 VPB.n330 VNB 0.13fF
C466 VPB.n331 VNB 0.15fF
C467 VPB.n332 VNB 0.02fF
C468 VPB.n333 VNB 0.02fF
C469 VPB.n334 VNB 0.02fF
C470 VPB.n335 VNB 0.13fF
C471 VPB.n336 VNB 0.14fF
C472 VPB.n337 VNB 0.02fF
C473 VPB.n338 VNB 0.02fF
C474 VPB.n339 VNB 0.02fF
C475 VPB.n340 VNB 0.10fF
C476 VPB.n341 VNB 0.02fF
C477 VPB.n342 VNB 0.13fF
C478 VPB.n343 VNB 0.16fF
C479 VPB.n344 VNB 0.02fF
C480 VPB.n345 VNB 0.02fF
C481 VPB.n346 VNB 0.02fF
C482 VPB.n347 VNB 0.13fF
C483 VPB.n348 VNB 0.16fF
C484 VPB.n349 VNB 0.02fF
C485 VPB.n350 VNB 0.02fF
C486 VPB.n351 VNB 0.02fF
C487 VPB.n352 VNB 0.06fF
C488 VPB.n353 VNB 0.21fF
C489 VPB.n354 VNB 0.02fF
C490 VPB.n355 VNB 0.01fF
C491 VPB.n356 VNB 0.02fF
C492 VPB.n357 VNB 0.27fF
C493 VPB.n358 VNB 0.02fF
C494 VPB.n359 VNB 0.02fF
C495 VPB.n360 VNB 0.02fF
C496 VPB.n361 VNB 0.27fF
C497 VPB.n362 VNB 0.01fF
C498 VPB.n363 VNB 0.02fF
C499 VPB.n364 VNB 0.04fF
C500 VPB.n365 VNB 0.02fF
C501 VPB.n366 VNB 0.02fF
C502 VPB.n367 VNB 0.02fF
C503 VPB.n368 VNB 0.04fF
C504 VPB.n369 VNB 0.02fF
C505 VPB.n370 VNB 0.28fF
C506 VPB.n371 VNB 0.04fF
C507 VPB.n373 VNB 0.02fF
C508 VPB.n374 VNB 0.02fF
C509 VPB.n375 VNB 0.02fF
C510 VPB.n376 VNB 0.02fF
C511 VPB.n378 VNB 0.02fF
C512 VPB.n379 VNB 0.02fF
C513 VPB.n380 VNB 0.02fF
C514 VPB.n382 VNB 0.27fF
C515 VPB.n384 VNB 0.03fF
C516 VPB.n385 VNB 0.02fF
C517 VPB.n386 VNB 0.03fF
C518 VPB.n387 VNB 0.03fF
C519 VPB.n388 VNB 0.27fF
C520 VPB.n389 VNB 0.01fF
C521 VPB.n390 VNB 0.02fF
C522 VPB.n391 VNB 0.04fF
C523 VPB.n392 VNB 0.27fF
C524 VPB.n393 VNB 0.02fF
C525 VPB.n394 VNB 0.02fF
C526 VPB.n395 VNB 0.02fF
C527 VPB.n396 VNB 0.05fF
C528 VPB.n397 VNB 0.20fF
C529 VPB.n398 VNB 0.02fF
C530 VPB.n399 VNB 0.01fF
C531 VPB.n400 VNB 0.02fF
C532 VPB.n401 VNB 0.13fF
C533 VPB.n402 VNB 0.16fF
C534 VPB.n403 VNB 0.02fF
C535 VPB.n404 VNB 0.02fF
C536 VPB.n405 VNB 0.02fF
C537 VPB.n406 VNB 0.10fF
C538 VPB.n407 VNB 0.02fF
C539 VPB.n408 VNB 0.13fF
C540 VPB.n409 VNB 0.16fF
C541 VPB.n410 VNB 0.02fF
C542 VPB.n411 VNB 0.02fF
C543 VPB.n412 VNB 0.02fF
C544 VPB.n413 VNB 0.13fF
C545 VPB.n414 VNB 0.15fF
C546 VPB.n415 VNB 0.02fF
C547 VPB.n416 VNB 0.02fF
C548 VPB.n417 VNB 0.02fF
C549 VPB.n418 VNB 0.13fF
C550 VPB.n419 VNB 0.14fF
C551 VPB.n420 VNB 0.02fF
C552 VPB.n421 VNB 0.02fF
C553 VPB.n422 VNB 0.02fF
C554 VPB.n423 VNB 0.10fF
C555 VPB.n424 VNB 0.02fF
C556 VPB.n425 VNB 0.13fF
C557 VPB.n426 VNB 0.16fF
C558 VPB.n427 VNB 0.02fF
C559 VPB.n428 VNB 0.02fF
C560 VPB.n429 VNB 0.02fF
C561 VPB.n430 VNB 0.13fF
C562 VPB.n431 VNB 0.16fF
C563 VPB.n432 VNB 0.02fF
C564 VPB.n433 VNB 0.02fF
C565 VPB.n434 VNB 0.02fF
C566 VPB.n435 VNB 0.02fF
C567 VPB.n436 VNB 0.02fF
C568 VPB.n437 VNB 0.04fF
C569 VPB.n438 VNB 0.04fF
C570 VPB.n439 VNB 0.02fF
C571 VPB.n440 VNB 0.02fF
C572 VPB.n441 VNB 0.02fF
C573 VPB.n442 VNB 0.02fF
C574 VPB.n443 VNB 0.02fF
C575 VPB.n444 VNB 0.02fF
C576 VPB.n445 VNB 0.03fF
C577 VPB.n446 VNB 0.03fF
C578 VPB.n447 VNB 0.02fF
C579 VPB.n448 VNB 0.02fF
C580 VPB.n449 VNB 0.02fF
C581 VPB.n450 VNB 0.04fF
C582 VPB.n451 VNB 0.04fF
C583 VPB.n453 VNB 0.42fF
.ends
