* SPICE3 file created from TMRDFFSNQX1.ext - technology: sky130A

.subckt TMRDFFSNQX1 Q D CLK SN VDD GND
X0 a_1905_1004 a_217_1004 VDD VDD pshort w=2 l=0.15 M=2
X1 GND a_217_1004 a_757_75 GND nshort w=3 l=0.15
X2 a_5227_383 a_6149_943 a_5922_182 GND nshort w=3 l=0.15
X3 VDD a_11673_1004 a_11033_943 VDD pshort w=2 l=0.15 M=2
X4 a_15044_181 a_8483_383 a_16096_73 GND nshort w=3 l=0.15
X5 a_5101_1004 a_5227_383 a_4996_73 GND nshort w=3 l=0.15
X6 GND D a_112_73 GND nshort w=3 l=0.15
X7 a_14869_1005 a_13367_383 a_15533_1005 VDD pshort w=2 l=0.15 M=2
X8 VDD a_343_383 a_217_1004 VDD pshort w=2 l=0.15 M=2
X9 VDD a_5227_383 a_5101_1004 VDD pshort w=2 l=0.15 M=2
X10 a_9178_182 SN a_8897_75 GND nshort w=3 l=0.15
X11 GND a_343_383 a_3368_73 GND nshort w=3 l=0.15
X12 VDD a_217_1004 a_343_383 VDD pshort w=2 l=0.15 M=2
X13 VDD a_15044_181 Q VDD pshort w=2 l=0.15 M=2
X14 a_11673_1004 a_11033_943 VDD VDD pshort w=2 l=0.15 M=2
X15 GND a_8357_1004 a_8897_75 GND nshort w=3 l=0.15
X16 VDD a_13241_1004 a_13367_383 VDD pshort w=2 l=0.15 M=2
X17 a_3473_1004 a_3599_383 VDD VDD pshort w=2 l=0.15 M=2
X18 a_10111_383 CLK VDD VDD pshort w=2 l=0.15 M=2
X19 a_6789_1004 a_6149_943 a_6884_182 GND nshort w=3 l=0.15
X20 a_5227_383 a_6149_943 VDD VDD pshort w=2 l=0.15 M=2
X21 a_13241_1004 a_13367_383 VDD VDD pshort w=2 l=0.15 M=2
X22 VDD a_11033_943 a_10111_383 VDD pshort w=2 l=0.15 M=2
X23 VDD a_5227_383 a_8357_1004 VDD pshort w=2 l=0.15 M=2
X24 a_6149_943 CLK VDD VDD pshort w=2 l=0.15 M=2
X25 a_14869_1005 a_13367_383 VDD VDD pshort w=2 l=0.15 M=2
X26 VDD a_6149_943 a_8483_383 VDD pshort w=2 l=0.15 M=2
X27 VDD CLK a_343_383 VDD pshort w=2 l=0.15 M=2
X28 VDD a_8483_383 a_14869_1005 VDD pshort w=2 l=0.15 M=2
X29 a_3473_1004 a_343_383 VDD VDD pshort w=2 l=0.15 M=2
X30 GND D a_9880_73 GND nshort w=3 l=0.15
X31 a_8483_383 SN VDD VDD pshort w=2 l=0.15 M=2
X32 VDD SN a_13367_383 VDD pshort w=2 l=0.15 M=2
X33 a_10111_383 a_9985_1004 VDD VDD pshort w=2 l=0.15 M=2
X34 VDD a_1905_1004 a_1265_943 VDD pshort w=2 l=0.15 M=2
X35 GND a_217_1004 a_1719_75 GND nshort w=3 l=0.15
X36 VDD a_10111_383 a_9985_1004 VDD pshort w=2 l=0.15 M=2
X37 a_11033_943 CLK a_12470_73 GND nshort w=3 l=0.15
X38 VDD SN a_11673_1004 VDD pshort w=2 l=0.15 M=2
X39 a_10111_383 a_11033_943 a_10806_182 GND nshort w=3 l=0.15
X40 a_6149_943 a_6789_1004 VDD VDD pshort w=2 l=0.15 M=2
X41 a_9985_1004 a_10111_383 a_9880_73 GND nshort w=3 l=0.15
X42 VDD a_3473_1004 a_3599_383 VDD pshort w=2 l=0.15 M=2
X43 a_15044_181 a_3599_383 a_15430_73 GND nshort w=3 l=0.15
X44 VDD a_1265_943 a_3599_383 VDD pshort w=2 l=0.15 M=2
X45 a_14062_182 SN a_13781_75 GND nshort w=3 l=0.15
X46 a_1038_182 CLK a_757_75 GND nshort w=3 l=0.15
X47 VDD a_1265_943 a_343_383 VDD pshort w=2 l=0.15 M=2
X48 a_8483_383 a_8357_1004 VDD VDD pshort w=2 l=0.15 M=2
X49 VDD a_11033_943 a_13367_383 VDD pshort w=2 l=0.15 M=2
X50 VDD a_5101_1004 a_5227_383 VDD pshort w=2 l=0.15 M=2
X51 a_15533_1005 a_3599_383 a_14869_1005 VDD pshort w=2 l=0.15 M=2
X52 a_217_1004 D VDD VDD pshort w=2 l=0.15 M=2
X53 GND a_10111_383 a_13136_73 GND nshort w=3 l=0.15
X54 GND a_1905_1004 a_2702_73 GND nshort w=3 l=0.15
X55 VDD D a_9985_1004 VDD pshort w=2 l=0.15 M=2
X56 a_1905_1004 a_1265_943 VDD VDD pshort w=2 l=0.15 M=2
X57 GND a_13241_1004 a_13781_75 GND nshort w=3 l=0.15
X58 a_6789_1004 a_5101_1004 VDD VDD pshort w=2 l=0.15 M=2
X59 GND a_5227_383 a_8252_73 GND nshort w=3 l=0.15
X60 VDD a_9985_1004 a_11673_1004 VDD pshort w=2 l=0.15 M=2
X61 a_217_1004 a_343_383 a_112_73 GND nshort w=3 l=0.15
X62 a_3599_383 a_1265_943 a_4294_182 GND nshort w=3 l=0.15
X63 a_11673_1004 a_11033_943 a_11768_182 GND nshort w=3 l=0.15
X64 GND a_5101_1004 a_5641_75 GND nshort w=3 l=0.15
X65 a_15044_181 a_8483_383 a_15533_1005 VDD pshort w=2 l=0.15 M=2
X66 a_2000_182 SN a_1719_75 GND nshort w=3 l=0.15
X67 VDD SN a_3599_383 VDD pshort w=2 l=0.15 M=2
X68 VDD SN a_6789_1004 VDD pshort w=2 l=0.15 M=2
X69 GND a_13367_383 a_14764_73 GND nshort w=3 l=0.15
X70 a_3473_1004 a_3599_383 a_3368_73 GND nshort w=3 l=0.15
X71 a_1905_1004 SN VDD VDD pshort w=2 l=0.15 M=2
X72 a_15044_181 a_3599_383 a_15533_1005 VDD pshort w=2 l=0.15 M=2
X73 VDD a_8483_383 a_8357_1004 VDD pshort w=2 l=0.15 M=2
X74 GND a_5101_1004 a_6603_75 GND nshort w=3 l=0.15
X75 VDD a_6149_943 a_6789_1004 VDD pshort w=2 l=0.15 M=2
X76 GND a_3473_1004 a_4013_75 GND nshort w=3 l=0.15
X77 VDD a_10111_383 a_13241_1004 VDD pshort w=2 l=0.15 M=2
X78 a_15044_181 a_8483_383 a_14764_73 GND nshort w=3 l=0.15
X79 a_5922_182 CLK a_5641_75 GND nshort w=3 l=0.15
X80 a_11033_943 CLK VDD VDD pshort w=2 l=0.15 M=2
X81 a_5101_1004 D VDD VDD pshort w=2 l=0.15 M=2
X82 GND a_6789_1004 a_7586_73 GND nshort w=3 l=0.15
X83 GND a_3599_383 a_16096_73 GND nshort w=3 l=0.15
X84 GND a_9985_1004 a_10525_75 GND nshort w=3 l=0.15
X85 GND D a_4996_73 GND nshort w=3 l=0.15
X86 VDD CLK a_1265_943 VDD pshort w=2 l=0.15 M=2
X87 a_1265_943 CLK a_2702_73 GND nshort w=3 l=0.15
X88 a_8483_383 a_6149_943 a_9178_182 GND nshort w=3 l=0.15
X89 a_8357_1004 a_8483_383 a_8252_73 GND nshort w=3 l=0.15
X90 Q a_15044_181 GND GND nshort w=3 l=0.15
X91 a_6884_182 SN a_6603_75 GND nshort w=3 l=0.15
X92 a_13241_1004 a_13367_383 a_13136_73 GND nshort w=3 l=0.15
X93 a_4294_182 SN a_4013_75 GND nshort w=3 l=0.15
X94 GND a_9985_1004 a_11487_75 GND nshort w=3 l=0.15
X95 VDD CLK a_5227_383 VDD pshort w=2 l=0.15 M=2
X96 a_1905_1004 a_1265_943 a_2000_182 GND nshort w=3 l=0.15
X97 a_10806_182 CLK a_10525_75 GND nshort w=3 l=0.15
X98 GND a_11673_1004 a_12470_73 GND nshort w=3 l=0.15
X99 GND a_13367_383 a_15430_73 GND nshort w=3 l=0.15
X100 a_343_383 a_1265_943 a_1038_182 GND nshort w=3 l=0.15
X101 a_13367_383 a_11033_943 a_14062_182 GND nshort w=3 l=0.15
X102 a_11768_182 SN a_11487_75 GND nshort w=3 l=0.15
X103 a_6149_943 CLK a_7586_73 GND nshort w=3 l=0.15
C0 VDD a_343_383 3.07fF
C1 VDD CLK 5.43fF
C2 VDD a_11033_943 2.18fF
C3 VDD a_6789_1004 2.09fF
C4 a_11673_1004 VDD 2.09fF
C5 VDD a_5227_383 3.07fF
C6 VDD a_3599_383 3.32fF
C7 D a_3599_383 7.23fF
C8 SN a_3599_383 2.73fF
C9 a_343_383 a_1265_943 2.89fF
C10 a_5227_383 a_6149_943 2.89fF
C11 VDD a_1905_1004 2.09fF
C12 a_3599_383 a_6149_943 3.76fF
C13 CLK a_10111_383 3.20fF
C14 a_10111_383 a_11033_943 2.89fF
C15 a_13367_383 VDD 3.26fF
C16 a_3599_383 a_8483_383 6.79fF
C17 CLK a_343_383 2.96fF
C18 D SN 3.25fF
C19 VDD a_6149_943 2.17fF
C20 a_5227_383 CLK 3.80fF
C21 CLK a_3599_383 2.31fF
C22 a_3599_383 a_11033_943 3.76fF
C23 VDD a_8483_383 3.43fF
C24 VDD a_1265_943 2.17fF
C25 VDD a_10111_383 3.07fF
C26 SN a_8483_383 2.57fF
C27 SN GND 3.93fF
C28 VDD GND 40.56fF
C29 a_8483_383 GND 2.13fF **FLOATING
C30 a_3599_383 GND 3.57fF **FLOATING
.ends
