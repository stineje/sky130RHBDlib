// File: DFFSNRNX1.spi.pex
// Created: Tue Oct 15 15:47:46 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_DFFSNRNX1\%GND ( 1 51 55 58 63 73 81 91 99 109 117 127 135 145 160 \
 164 166 168 170 172 174 175 176 177 178 179 )
c308 ( 179 0 ) capacitor c=0.0226224f //x=24.935 //y=0.875
c309 ( 178 0 ) capacitor c=0.0226224f //x=20.125 //y=0.875
c310 ( 177 0 ) capacitor c=0.0226224f //x=15.315 //y=0.875
c311 ( 176 0 ) capacitor c=0.0226413f //x=10.505 //y=0.875
c312 ( 175 0 ) capacitor c=0.0226413f //x=5.695 //y=0.875
c313 ( 174 0 ) capacitor c=0.0226959f //x=0.885 //y=0.875
c314 ( 173 0 ) capacitor c=0.00440144f //x=25.125 //y=0
c315 ( 172 0 ) capacitor c=0.108597f //x=24.05 //y=0
c316 ( 171 0 ) capacitor c=0.00440144f //x=20.315 //y=0
c317 ( 170 0 ) capacitor c=0.108683f //x=19.24 //y=0
c318 ( 169 0 ) capacitor c=0.00440144f //x=15.505 //y=0
c319 ( 168 0 ) capacitor c=0.108636f //x=14.43 //y=0
c320 ( 167 0 ) capacitor c=0.00440144f //x=10.695 //y=0
c321 ( 166 0 ) capacitor c=0.107929f //x=9.62 //y=0
c322 ( 165 0 ) capacitor c=0.00440144f //x=5.885 //y=0
c323 ( 164 0 ) capacitor c=0.108262f //x=4.81 //y=0
c324 ( 163 0 ) capacitor c=0.00440144f //x=1.075 //y=0
c325 ( 160 0 ) capacitor c=0.321926f //x=28.12 //y=0
c326 ( 145 0 ) capacitor c=0.0339482f //x=25.04 //y=0
c327 ( 135 0 ) capacitor c=0.133515f //x=23.88 //y=0
c328 ( 127 0 ) capacitor c=0.0339482f //x=20.23 //y=0
c329 ( 117 0 ) capacitor c=0.133515f //x=19.07 //y=0
c330 ( 109 0 ) capacitor c=0.0339482f //x=15.42 //y=0
c331 ( 99 0 ) capacitor c=0.133551f //x=14.26 //y=0
c332 ( 91 0 ) capacitor c=0.0339619f //x=10.61 //y=0
c333 ( 81 0 ) capacitor c=0.13365f //x=9.45 //y=0
c334 ( 73 0 ) capacitor c=0.0339619f //x=5.8 //y=0
c335 ( 63 0 ) capacitor c=0.131658f //x=4.64 //y=0
c336 ( 58 0 ) capacitor c=0.178285f //x=0.74 //y=0
c337 ( 55 0 ) capacitor c=0.0367385f //x=0.99 //y=0
c338 ( 51 0 ) capacitor c=0.897892f //x=28.12 //y=0
r339 (  158 160 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=27.01 //y=0 //x2=28.12 //y2=0
r340 (  156 158 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=25.9 //y=0 //x2=27.01 //y2=0
r341 (  154 173 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.21 //y=0 //x2=25.125 //y2=0
r342 (  154 156 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=25.21 //y=0 //x2=25.9 //y2=0
r343 (  149 173 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.125 //y=0.17 //x2=25.125 //y2=0
r344 (  149 179 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=25.125 //y=0.17 //x2=25.125 //y2=0.965
r345 (  146 172 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.22 //y=0 //x2=24.05 //y2=0
r346 (  146 148 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.22 //y=0 //x2=24.79 //y2=0
r347 (  145 173 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.04 //y=0 //x2=25.125 //y2=0
r348 (  145 148 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=25.04 //y=0 //x2=24.79 //y2=0
r349 (  140 142 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=22.2 //y=0 //x2=23.31 //y2=0
r350 (  138 140 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=21.09 //y=0 //x2=22.2 //y2=0
r351 (  136 171 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.4 //y=0 //x2=20.315 //y2=0
r352 (  136 138 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=20.4 //y=0 //x2=21.09 //y2=0
r353 (  135 172 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.88 //y=0 //x2=24.05 //y2=0
r354 (  135 142 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=23.88 //y=0 //x2=23.31 //y2=0
r355 (  131 171 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.315 //y=0.17 //x2=20.315 //y2=0
r356 (  131 178 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=20.315 //y=0.17 //x2=20.315 //y2=0.965
r357 (  128 170 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.41 //y=0 //x2=19.24 //y2=0
r358 (  128 130 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.41 //y=0 //x2=19.98 //y2=0
r359 (  127 171 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.23 //y=0 //x2=20.315 //y2=0
r360 (  127 130 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=20.23 //y=0 //x2=19.98 //y2=0
r361 (  122 124 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=17.39 //y=0 //x2=18.5 //y2=0
r362 (  120 122 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=16.28 //y=0 //x2=17.39 //y2=0
r363 (  118 169 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.59 //y=0 //x2=15.505 //y2=0
r364 (  118 120 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=15.59 //y=0 //x2=16.28 //y2=0
r365 (  117 170 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.07 //y=0 //x2=19.24 //y2=0
r366 (  117 124 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.07 //y=0 //x2=18.5 //y2=0
r367 (  113 169 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.505 //y=0.17 //x2=15.505 //y2=0
r368 (  113 177 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=15.505 //y=0.17 //x2=15.505 //y2=0.965
r369 (  110 168 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.6 //y=0 //x2=14.43 //y2=0
r370 (  110 112 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.6 //y=0 //x2=15.17 //y2=0
r371 (  109 169 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.42 //y=0 //x2=15.505 //y2=0
r372 (  109 112 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=15.42 //y=0 //x2=15.17 //y2=0
r373 (  104 106 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=12.58 //y=0 //x2=13.69 //y2=0
r374 (  102 104 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=11.47 //y=0 //x2=12.58 //y2=0
r375 (  100 167 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.78 //y=0 //x2=10.695 //y2=0
r376 (  100 102 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=10.78 //y=0 //x2=11.47 //y2=0
r377 (  99 168 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.26 //y=0 //x2=14.43 //y2=0
r378 (  99 106 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.26 //y=0 //x2=13.69 //y2=0
r379 (  95 167 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.695 //y=0.17 //x2=10.695 //y2=0
r380 (  95 176 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=10.695 //y=0.17 //x2=10.695 //y2=0.965
r381 (  92 166 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.79 //y=0 //x2=9.62 //y2=0
r382 (  92 94 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.79 //y=0 //x2=10.36 //y2=0
r383 (  91 167 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.61 //y=0 //x2=10.695 //y2=0
r384 (  91 94 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=10.61 //y=0 //x2=10.36 //y2=0
r385 (  86 88 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=7.77 //y=0 //x2=8.88 //y2=0
r386 (  84 86 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r387 (  82 165 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.97 //y=0 //x2=5.885 //y2=0
r388 (  82 84 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=5.97 //y=0 //x2=6.66 //y2=0
r389 (  81 166 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.45 //y=0 //x2=9.62 //y2=0
r390 (  81 88 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.45 //y=0 //x2=8.88 //y2=0
r391 (  77 165 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.885 //y=0.17 //x2=5.885 //y2=0
r392 (  77 175 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=5.885 //y=0.17 //x2=5.885 //y2=0.965
r393 (  74 164 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=4.81 //y2=0
r394 (  74 76 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=5.55 //y2=0
r395 (  73 165 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.8 //y=0 //x2=5.885 //y2=0
r396 (  73 76 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=5.8 //y=0 //x2=5.55 //y2=0
r397 (  68 70 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=0 //x2=4.07 //y2=0
r398 (  66 68 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r399 (  64 163 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.075 //y2=0
r400 (  64 66 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.85 //y2=0
r401 (  63 164 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.81 //y2=0
r402 (  63 70 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.07 //y2=0
r403 (  59 163 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0
r404 (  59 174 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0.965
r405 (  55 163 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=1.075 //y2=0
r406 (  55 58 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=0.74 //y2=0
r407 (  51 160 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.12 //y=0 //x2=28.12 //y2=0
r408 (  49 158 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.01 //y=0 //x2=27.01 //y2=0
r409 (  49 51 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=27.01 //y=0 //x2=28.12 //y2=0
r410 (  47 156 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.9 //y=0 //x2=25.9 //y2=0
r411 (  47 49 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=25.9 //y=0 //x2=27.01 //y2=0
r412 (  45 148 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=0 //x2=24.79 //y2=0
r413 (  45 47 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=0 //x2=25.9 //y2=0
r414 (  43 142 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.31 //y=0 //x2=23.31 //y2=0
r415 (  43 45 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=23.31 //y=0 //x2=24.79 //y2=0
r416 (  41 140 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.2 //y=0 //x2=22.2 //y2=0
r417 (  41 43 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.2 //y=0 //x2=23.31 //y2=0
r418 (  39 138 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=0 //x2=21.09 //y2=0
r419 (  39 41 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=0 //x2=22.2 //y2=0
r420 (  37 130 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=0 //x2=19.98 //y2=0
r421 (  37 39 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=0 //x2=21.09 //y2=0
r422 (  35 124 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=0 //x2=18.5 //y2=0
r423 (  35 37 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=0 //x2=19.98 //y2=0
r424 (  33 122 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=0 //x2=17.39 //y2=0
r425 (  33 35 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=0 //x2=18.5 //y2=0
r426 (  31 120 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=0 //x2=16.28 //y2=0
r427 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=0 //x2=17.39 //y2=0
r428 (  29 112 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=0 //x2=15.17 //y2=0
r429 (  29 31 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=0 //x2=16.28 //y2=0
r430 (  26 106 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=0 //x2=13.69 //y2=0
r431 (  24 104 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=0 //x2=12.58 //y2=0
r432 (  24 26 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=0 //x2=13.69 //y2=0
r433 (  22 102 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=0 //x2=11.47 //y2=0
r434 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=0 //x2=12.58 //y2=0
r435 (  20 94 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r436 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=0 //x2=11.47 //y2=0
r437 (  18 88 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.88 //y=0 //x2=8.88 //y2=0
r438 (  18 20 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.88 //y=0 //x2=10.36 //y2=0
r439 (  16 86 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r440 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=8.88 //y2=0
r441 (  14 84 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r442 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r443 (  12 76 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r444 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r445 (  10 70 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r446 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=0 //x2=5.55 //y2=0
r447 (  8 68 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r448 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.07 //y2=0
r449 (  6 66 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r450 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r451 (  3 58 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r452 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r453 (  1 29 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=14.43 //y=0 //x2=15.17 //y2=0
r454 (  1 26 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=14.43 //y=0 //x2=13.69 //y2=0
ends PM_DFFSNRNX1\%GND

subckt PM_DFFSNRNX1\%VDD ( 1 51 58 65 75 83 93 99 109 119 127 137 143 153 163 \
 171 181 187 197 207 215 225 231 241 251 259 269 275 285 295 303 316 323 328 \
 333 338 343 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362 363 \
 364 365 366 367 368 369 370 371 )
c342 ( 371 0 ) capacitor c=0.0453711f //x=27.635 //y=5.02
c343 ( 370 0 ) capacitor c=0.02424f //x=26.755 //y=5.02
c344 ( 369 0 ) capacitor c=0.02424f //x=25.875 //y=5.02
c345 ( 368 0 ) capacitor c=0.0531793f //x=25.005 //y=5.02
c346 ( 367 0 ) capacitor c=0.0453059f //x=22.825 //y=5.02
c347 ( 366 0 ) capacitor c=0.02424f //x=21.945 //y=5.02
c348 ( 365 0 ) capacitor c=0.024152f //x=21.065 //y=5.02
c349 ( 364 0 ) capacitor c=0.053132f //x=20.195 //y=5.02
c350 ( 363 0 ) capacitor c=0.0452179f //x=18.015 //y=5.02
c351 ( 362 0 ) capacitor c=0.024152f //x=17.135 //y=5.02
c352 ( 361 0 ) capacitor c=0.024152f //x=16.255 //y=5.02
c353 ( 360 0 ) capacitor c=0.053132f //x=15.385 //y=5.02
c354 ( 359 0 ) capacitor c=0.0452179f //x=13.205 //y=5.02
c355 ( 358 0 ) capacitor c=0.024152f //x=12.325 //y=5.02
c356 ( 357 0 ) capacitor c=0.024152f //x=11.445 //y=5.02
c357 ( 356 0 ) capacitor c=0.053132f //x=10.575 //y=5.02
c358 ( 355 0 ) capacitor c=0.0452179f //x=8.395 //y=5.02
c359 ( 354 0 ) capacitor c=0.024152f //x=7.515 //y=5.02
c360 ( 353 0 ) capacitor c=0.024152f //x=6.635 //y=5.02
c361 ( 352 0 ) capacitor c=0.053132f //x=5.765 //y=5.02
c362 ( 351 0 ) capacitor c=0.0452179f //x=3.585 //y=5.02
c363 ( 350 0 ) capacitor c=0.024152f //x=2.705 //y=5.02
c364 ( 349 0 ) capacitor c=0.0244794f //x=1.825 //y=5.02
c365 ( 348 0 ) capacitor c=0.0533644f //x=0.955 //y=5.02
c366 ( 347 0 ) capacitor c=0.00591168f //x=27.78 //y=7.4
c367 ( 346 0 ) capacitor c=0.00591168f //x=26.9 //y=7.4
c368 ( 345 0 ) capacitor c=0.00591168f //x=26.02 //y=7.4
c369 ( 344 0 ) capacitor c=0.00591168f //x=25.14 //y=7.4
c370 ( 343 0 ) capacitor c=0.157232f //x=24.05 //y=7.4
c371 ( 342 0 ) capacitor c=0.00591168f //x=22.97 //y=7.4
c372 ( 341 0 ) capacitor c=0.00591168f //x=22.09 //y=7.4
c373 ( 340 0 ) capacitor c=0.00591168f //x=21.21 //y=7.4
c374 ( 339 0 ) capacitor c=0.00591168f //x=20.33 //y=7.4
c375 ( 338 0 ) capacitor c=0.154937f //x=19.24 //y=7.4
c376 ( 337 0 ) capacitor c=0.00591168f //x=18.16 //y=7.4
c377 ( 336 0 ) capacitor c=0.00591168f //x=17.28 //y=7.4
c378 ( 335 0 ) capacitor c=0.00591168f //x=16.4 //y=7.4
c379 ( 334 0 ) capacitor c=0.00591168f //x=15.52 //y=7.4
c380 ( 333 0 ) capacitor c=0.155149f //x=14.43 //y=7.4
c381 ( 332 0 ) capacitor c=0.00591168f //x=13.35 //y=7.4
c382 ( 331 0 ) capacitor c=0.00591168f //x=12.47 //y=7.4
c383 ( 330 0 ) capacitor c=0.00591168f //x=11.59 //y=7.4
c384 ( 329 0 ) capacitor c=0.00591168f //x=10.71 //y=7.4
c385 ( 328 0 ) capacitor c=0.15516f //x=9.62 //y=7.4
c386 ( 327 0 ) capacitor c=0.00591168f //x=8.54 //y=7.4
c387 ( 326 0 ) capacitor c=0.00591168f //x=7.66 //y=7.4
c388 ( 325 0 ) capacitor c=0.00591168f //x=6.78 //y=7.4
c389 ( 324 0 ) capacitor c=0.00591168f //x=5.9 //y=7.4
c390 ( 323 0 ) capacitor c=0.159704f //x=4.81 //y=7.4
c391 ( 322 0 ) capacitor c=0.00591168f //x=3.73 //y=7.4
c392 ( 321 0 ) capacitor c=0.00591168f //x=2.85 //y=7.4
c393 ( 320 0 ) capacitor c=0.00591168f //x=1.97 //y=7.4
c394 ( 319 0 ) capacitor c=0.00591168f //x=1.09 //y=7.4
c395 ( 316 0 ) capacitor c=0.272103f //x=28.12 //y=7.4
c396 ( 303 0 ) capacitor c=0.0288171f //x=27.695 //y=7.4
c397 ( 295 0 ) capacitor c=0.0287757f //x=26.815 //y=7.4
c398 ( 285 0 ) capacitor c=0.028511f //x=25.935 //y=7.4
c399 ( 275 0 ) capacitor c=0.0383672f //x=25.055 //y=7.4
c400 ( 269 0 ) capacitor c=0.0395236f //x=23.88 //y=7.4
c401 ( 259 0 ) capacitor c=0.0288769f //x=22.885 //y=7.4
c402 ( 251 0 ) capacitor c=0.0287624f //x=22.005 //y=7.4
c403 ( 241 0 ) capacitor c=0.0284966f //x=21.125 //y=7.4
c404 ( 231 0 ) capacitor c=0.0383672f //x=20.245 //y=7.4
c405 ( 225 0 ) capacitor c=0.0394667f //x=19.07 //y=7.4
c406 ( 215 0 ) capacitor c=0.028847f //x=18.075 //y=7.4
c407 ( 207 0 ) capacitor c=0.0287514f //x=17.195 //y=7.4
c408 ( 197 0 ) capacitor c=0.0284966f //x=16.315 //y=7.4
c409 ( 187 0 ) capacitor c=0.0383672f //x=15.435 //y=7.4
c410 ( 181 0 ) capacitor c=0.0394667f //x=14.26 //y=7.4
c411 ( 171 0 ) capacitor c=0.0288488f //x=13.265 //y=7.4
c412 ( 163 0 ) capacitor c=0.0287514f //x=12.385 //y=7.4
c413 ( 153 0 ) capacitor c=0.0284966f //x=11.505 //y=7.4
c414 ( 143 0 ) capacitor c=0.0383672f //x=10.625 //y=7.4
c415 ( 137 0 ) capacitor c=0.0394667f //x=9.45 //y=7.4
c416 ( 127 0 ) capacitor c=0.0288488f //x=8.455 //y=7.4
c417 ( 119 0 ) capacitor c=0.0287514f //x=7.575 //y=7.4
c418 ( 109 0 ) capacitor c=0.0284966f //x=6.695 //y=7.4
c419 ( 99 0 ) capacitor c=0.0383672f //x=5.815 //y=7.4
c420 ( 93 0 ) capacitor c=0.0394667f //x=4.64 //y=7.4
c421 ( 83 0 ) capacitor c=0.0288488f //x=3.645 //y=7.4
c422 ( 75 0 ) capacitor c=0.0287505f //x=2.765 //y=7.4
c423 ( 65 0 ) capacitor c=0.0292055f //x=1.885 //y=7.4
c424 ( 58 0 ) capacitor c=0.234703f //x=0.74 //y=7.4
c425 ( 55 0 ) capacitor c=0.0452081f //x=1.005 //y=7.4
c426 ( 51 0 ) capacitor c=1.00405f //x=28.12 //y=7.4
r427 (  314 347 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.865 //y=7.4 //x2=27.78 //y2=7.4
r428 (  314 316 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=27.865 //y=7.4 //x2=28.12 //y2=7.4
r429 (  307 347 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.78 //y=7.23 //x2=27.78 //y2=7.4
r430 (  307 371 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=27.78 //y=7.23 //x2=27.78 //y2=6.745
r431 (  304 346 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.985 //y=7.4 //x2=26.9 //y2=7.4
r432 (  304 306 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=26.985 //y=7.4 //x2=27.01 //y2=7.4
r433 (  303 347 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.695 //y=7.4 //x2=27.78 //y2=7.4
r434 (  303 306 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=27.695 //y=7.4 //x2=27.01 //y2=7.4
r435 (  297 346 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.9 //y=7.23 //x2=26.9 //y2=7.4
r436 (  297 370 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.9 //y=7.23 //x2=26.9 //y2=6.745
r437 (  296 345 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.105 //y=7.4 //x2=26.02 //y2=7.4
r438 (  295 346 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.815 //y=7.4 //x2=26.9 //y2=7.4
r439 (  295 296 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=26.815 //y=7.4 //x2=26.105 //y2=7.4
r440 (  289 345 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.02 //y=7.23 //x2=26.02 //y2=7.4
r441 (  289 369 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.02 //y=7.23 //x2=26.02 //y2=6.745
r442 (  286 344 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.225 //y=7.4 //x2=25.14 //y2=7.4
r443 (  286 288 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=25.225 //y=7.4 //x2=25.9 //y2=7.4
r444 (  285 345 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.935 //y=7.4 //x2=26.02 //y2=7.4
r445 (  285 288 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=25.935 //y=7.4 //x2=25.9 //y2=7.4
r446 (  279 344 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.14 //y=7.23 //x2=25.14 //y2=7.4
r447 (  279 368 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=25.14 //y=7.23 //x2=25.14 //y2=6.405
r448 (  276 343 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.22 //y=7.4 //x2=24.05 //y2=7.4
r449 (  276 278 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.22 //y=7.4 //x2=24.79 //y2=7.4
r450 (  275 344 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.055 //y=7.4 //x2=25.14 //y2=7.4
r451 (  275 278 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=25.055 //y=7.4 //x2=24.79 //y2=7.4
r452 (  270 342 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.055 //y=7.4 //x2=22.97 //y2=7.4
r453 (  270 272 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=23.055 //y=7.4 //x2=23.31 //y2=7.4
r454 (  269 343 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.88 //y=7.4 //x2=24.05 //y2=7.4
r455 (  269 272 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=23.88 //y=7.4 //x2=23.31 //y2=7.4
r456 (  263 342 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.97 //y=7.23 //x2=22.97 //y2=7.4
r457 (  263 367 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.97 //y=7.23 //x2=22.97 //y2=6.745
r458 (  260 341 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.175 //y=7.4 //x2=22.09 //y2=7.4
r459 (  260 262 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=22.175 //y=7.4 //x2=22.2 //y2=7.4
r460 (  259 342 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.885 //y=7.4 //x2=22.97 //y2=7.4
r461 (  259 262 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=22.885 //y=7.4 //x2=22.2 //y2=7.4
r462 (  253 341 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.09 //y=7.23 //x2=22.09 //y2=7.4
r463 (  253 366 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.09 //y=7.23 //x2=22.09 //y2=6.745
r464 (  252 340 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.295 //y=7.4 //x2=21.21 //y2=7.4
r465 (  251 341 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.005 //y=7.4 //x2=22.09 //y2=7.4
r466 (  251 252 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.005 //y=7.4 //x2=21.295 //y2=7.4
r467 (  245 340 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.21 //y=7.23 //x2=21.21 //y2=7.4
r468 (  245 365 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.21 //y=7.23 //x2=21.21 //y2=6.745
r469 (  242 339 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.415 //y=7.4 //x2=20.33 //y2=7.4
r470 (  242 244 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=20.415 //y=7.4 //x2=21.09 //y2=7.4
r471 (  241 340 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.125 //y=7.4 //x2=21.21 //y2=7.4
r472 (  241 244 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=21.125 //y=7.4 //x2=21.09 //y2=7.4
r473 (  235 339 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.33 //y=7.23 //x2=20.33 //y2=7.4
r474 (  235 364 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=20.33 //y=7.23 //x2=20.33 //y2=6.405
r475 (  232 338 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.41 //y=7.4 //x2=19.24 //y2=7.4
r476 (  232 234 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.41 //y=7.4 //x2=19.98 //y2=7.4
r477 (  231 339 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.245 //y=7.4 //x2=20.33 //y2=7.4
r478 (  231 234 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=20.245 //y=7.4 //x2=19.98 //y2=7.4
r479 (  226 337 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.245 //y=7.4 //x2=18.16 //y2=7.4
r480 (  226 228 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=18.245 //y=7.4 //x2=18.5 //y2=7.4
r481 (  225 338 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.07 //y=7.4 //x2=19.24 //y2=7.4
r482 (  225 228 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.07 //y=7.4 //x2=18.5 //y2=7.4
r483 (  219 337 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.16 //y=7.23 //x2=18.16 //y2=7.4
r484 (  219 363 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=18.16 //y=7.23 //x2=18.16 //y2=6.745
r485 (  216 336 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.365 //y=7.4 //x2=17.28 //y2=7.4
r486 (  216 218 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=17.365 //y=7.4 //x2=17.39 //y2=7.4
r487 (  215 337 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.075 //y=7.4 //x2=18.16 //y2=7.4
r488 (  215 218 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=18.075 //y=7.4 //x2=17.39 //y2=7.4
r489 (  209 336 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.28 //y=7.23 //x2=17.28 //y2=7.4
r490 (  209 362 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.28 //y=7.23 //x2=17.28 //y2=6.745
r491 (  208 335 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.485 //y=7.4 //x2=16.4 //y2=7.4
r492 (  207 336 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.195 //y=7.4 //x2=17.28 //y2=7.4
r493 (  207 208 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=17.195 //y=7.4 //x2=16.485 //y2=7.4
r494 (  201 335 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.4 //y=7.23 //x2=16.4 //y2=7.4
r495 (  201 361 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.4 //y=7.23 //x2=16.4 //y2=6.745
r496 (  198 334 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.605 //y=7.4 //x2=15.52 //y2=7.4
r497 (  198 200 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=15.605 //y=7.4 //x2=16.28 //y2=7.4
r498 (  197 335 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.315 //y=7.4 //x2=16.4 //y2=7.4
r499 (  197 200 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=16.315 //y=7.4 //x2=16.28 //y2=7.4
r500 (  191 334 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.52 //y=7.23 //x2=15.52 //y2=7.4
r501 (  191 360 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=15.52 //y=7.23 //x2=15.52 //y2=6.405
r502 (  188 333 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.6 //y=7.4 //x2=14.43 //y2=7.4
r503 (  188 190 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.6 //y=7.4 //x2=15.17 //y2=7.4
r504 (  187 334 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.435 //y=7.4 //x2=15.52 //y2=7.4
r505 (  187 190 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=15.435 //y=7.4 //x2=15.17 //y2=7.4
r506 (  182 332 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.435 //y=7.4 //x2=13.35 //y2=7.4
r507 (  182 184 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=13.435 //y=7.4 //x2=13.69 //y2=7.4
r508 (  181 333 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.26 //y=7.4 //x2=14.43 //y2=7.4
r509 (  181 184 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.26 //y=7.4 //x2=13.69 //y2=7.4
r510 (  175 332 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.35 //y=7.23 //x2=13.35 //y2=7.4
r511 (  175 359 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=13.35 //y=7.23 //x2=13.35 //y2=6.745
r512 (  172 331 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.555 //y=7.4 //x2=12.47 //y2=7.4
r513 (  172 174 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=12.555 //y=7.4 //x2=12.58 //y2=7.4
r514 (  171 332 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.265 //y=7.4 //x2=13.35 //y2=7.4
r515 (  171 174 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=13.265 //y=7.4 //x2=12.58 //y2=7.4
r516 (  165 331 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.47 //y=7.23 //x2=12.47 //y2=7.4
r517 (  165 358 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.47 //y=7.23 //x2=12.47 //y2=6.745
r518 (  164 330 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.675 //y=7.4 //x2=11.59 //y2=7.4
r519 (  163 331 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.385 //y=7.4 //x2=12.47 //y2=7.4
r520 (  163 164 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=12.385 //y=7.4 //x2=11.675 //y2=7.4
r521 (  157 330 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.59 //y=7.23 //x2=11.59 //y2=7.4
r522 (  157 357 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.59 //y=7.23 //x2=11.59 //y2=6.745
r523 (  154 329 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.795 //y=7.4 //x2=10.71 //y2=7.4
r524 (  154 156 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=10.795 //y=7.4 //x2=11.47 //y2=7.4
r525 (  153 330 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.505 //y=7.4 //x2=11.59 //y2=7.4
r526 (  153 156 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=11.505 //y=7.4 //x2=11.47 //y2=7.4
r527 (  147 329 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.71 //y=7.23 //x2=10.71 //y2=7.4
r528 (  147 356 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=10.71 //y=7.23 //x2=10.71 //y2=6.405
r529 (  144 328 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.79 //y=7.4 //x2=9.62 //y2=7.4
r530 (  144 146 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.79 //y=7.4 //x2=10.36 //y2=7.4
r531 (  143 329 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.625 //y=7.4 //x2=10.71 //y2=7.4
r532 (  143 146 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=10.625 //y=7.4 //x2=10.36 //y2=7.4
r533 (  138 327 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.625 //y=7.4 //x2=8.54 //y2=7.4
r534 (  138 140 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=8.625 //y=7.4 //x2=8.88 //y2=7.4
r535 (  137 328 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.45 //y=7.4 //x2=9.62 //y2=7.4
r536 (  137 140 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.45 //y=7.4 //x2=8.88 //y2=7.4
r537 (  131 327 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.54 //y=7.23 //x2=8.54 //y2=7.4
r538 (  131 355 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.54 //y=7.23 //x2=8.54 //y2=6.745
r539 (  128 326 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.745 //y=7.4 //x2=7.66 //y2=7.4
r540 (  128 130 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=7.745 //y=7.4 //x2=7.77 //y2=7.4
r541 (  127 327 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.455 //y=7.4 //x2=8.54 //y2=7.4
r542 (  127 130 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=8.455 //y=7.4 //x2=7.77 //y2=7.4
r543 (  121 326 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.66 //y=7.23 //x2=7.66 //y2=7.4
r544 (  121 354 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.66 //y=7.23 //x2=7.66 //y2=6.745
r545 (  120 325 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.865 //y=7.4 //x2=6.78 //y2=7.4
r546 (  119 326 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.575 //y=7.4 //x2=7.66 //y2=7.4
r547 (  119 120 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.575 //y=7.4 //x2=6.865 //y2=7.4
r548 (  113 325 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=7.4
r549 (  113 353 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=6.745
r550 (  110 324 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.985 //y=7.4 //x2=5.9 //y2=7.4
r551 (  110 112 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=5.985 //y=7.4 //x2=6.66 //y2=7.4
r552 (  109 325 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.78 //y2=7.4
r553 (  109 112 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.66 //y2=7.4
r554 (  103 324 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.9 //y=7.23 //x2=5.9 //y2=7.4
r555 (  103 352 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=5.9 //y=7.23 //x2=5.9 //y2=6.405
r556 (  100 323 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=4.81 //y2=7.4
r557 (  100 102 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=5.55 //y2=7.4
r558 (  99 324 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.815 //y=7.4 //x2=5.9 //y2=7.4
r559 (  99 102 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=5.815 //y=7.4 //x2=5.55 //y2=7.4
r560 (  94 322 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=3.73 //y2=7.4
r561 (  94 96 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=4.07 //y2=7.4
r562 (  93 323 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.81 //y2=7.4
r563 (  93 96 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.07 //y2=7.4
r564 (  87 322 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=7.4
r565 (  87 351 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=6.745
r566 (  84 321 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.85 //y2=7.4
r567 (  84 86 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.96 //y2=7.4
r568 (  83 322 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=3.73 //y2=7.4
r569 (  83 86 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=2.96 //y2=7.4
r570 (  77 321 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=7.4
r571 (  77 350 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=6.745
r572 (  76 320 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.055 //y=7.4 //x2=1.97 //y2=7.4
r573 (  75 321 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.85 //y2=7.4
r574 (  75 76 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.055 //y2=7.4
r575 (  69 320 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=7.4
r576 (  69 349 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=6.745
r577 (  66 319 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.09 //y2=7.4
r578 (  66 68 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.85 //y2=7.4
r579 (  65 320 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.97 //y2=7.4
r580 (  65 68 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.85 //y2=7.4
r581 (  59 319 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=7.4
r582 (  59 348 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=6.405
r583 (  55 319 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=1.09 //y2=7.4
r584 (  55 58 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=0.74 //y2=7.4
r585 (  51 316 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.12 //y=7.4 //x2=28.12 //y2=7.4
r586 (  49 306 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.01 //y=7.4 //x2=27.01 //y2=7.4
r587 (  49 51 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=27.01 //y=7.4 //x2=28.12 //y2=7.4
r588 (  47 288 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.9 //y=7.4 //x2=25.9 //y2=7.4
r589 (  47 49 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=25.9 //y=7.4 //x2=27.01 //y2=7.4
r590 (  45 278 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=7.4 //x2=24.79 //y2=7.4
r591 (  45 47 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=7.4 //x2=25.9 //y2=7.4
r592 (  43 272 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.31 //y=7.4 //x2=23.31 //y2=7.4
r593 (  43 45 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=23.31 //y=7.4 //x2=24.79 //y2=7.4
r594 (  41 262 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.2 //y=7.4 //x2=22.2 //y2=7.4
r595 (  41 43 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.2 //y=7.4 //x2=23.31 //y2=7.4
r596 (  39 244 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=7.4 //x2=21.09 //y2=7.4
r597 (  39 41 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=7.4 //x2=22.2 //y2=7.4
r598 (  37 234 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=7.4 //x2=19.98 //y2=7.4
r599 (  37 39 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=7.4 //x2=21.09 //y2=7.4
r600 (  35 228 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=7.4 //x2=18.5 //y2=7.4
r601 (  35 37 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=7.4 //x2=19.98 //y2=7.4
r602 (  33 218 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=7.4 //x2=17.39 //y2=7.4
r603 (  33 35 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=7.4 //x2=18.5 //y2=7.4
r604 (  31 200 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=7.4 //x2=16.28 //y2=7.4
r605 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=7.4 //x2=17.39 //y2=7.4
r606 (  29 190 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=7.4 //x2=15.17 //y2=7.4
r607 (  29 31 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=7.4 //x2=16.28 //y2=7.4
r608 (  26 184 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=7.4 //x2=13.69 //y2=7.4
r609 (  24 174 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=7.4 //x2=12.58 //y2=7.4
r610 (  24 26 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=7.4 //x2=13.69 //y2=7.4
r611 (  22 156 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=7.4 //x2=11.47 //y2=7.4
r612 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=7.4 //x2=12.58 //y2=7.4
r613 (  20 146 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r614 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=7.4 //x2=11.47 //y2=7.4
r615 (  18 140 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.88 //y=7.4 //x2=8.88 //y2=7.4
r616 (  18 20 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.88 //y=7.4 //x2=10.36 //y2=7.4
r617 (  16 130 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=7.4 //x2=7.77 //y2=7.4
r618 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=7.4 //x2=8.88 //y2=7.4
r619 (  14 112 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r620 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.4 //x2=7.77 //y2=7.4
r621 (  12 102 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r622 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.66 //y2=7.4
r623 (  10 96 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=7.4 //x2=4.07 //y2=7.4
r624 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=7.4 //x2=5.55 //y2=7.4
r625 (  8 86 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r626 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r627 (  6 68 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r628 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r629 (  3 58 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r630 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r631 (  1 29 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=14.43 //y=7.4 //x2=15.17 //y2=7.4
r632 (  1 26 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=14.43 //y=7.4 //x2=13.69 //y2=7.4
ends PM_DFFSNRNX1\%VDD

subckt PM_DFFSNRNX1\%noxref_3 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 63 64 \
 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 92 94 100 101 102 103 \
 123 125 126 127 )
c251 ( 127 0 ) capacitor c=0.023087f //x=3.145 //y=5.02
c252 ( 126 0 ) capacitor c=0.023519f //x=2.265 //y=5.02
c253 ( 125 0 ) capacitor c=0.0224735f //x=1.385 //y=5.02
c254 ( 123 0 ) capacitor c=0.00853354f //x=3.395 //y=0.915
c255 ( 103 0 ) capacitor c=0.0556143f //x=11.005 //y=4.79
c256 ( 102 0 ) capacitor c=0.0293157f //x=11.295 //y=4.79
c257 ( 101 0 ) capacitor c=0.0347816f //x=10.96 //y=1.22
c258 ( 100 0 ) capacitor c=0.0187487f //x=10.96 //y=0.875
c259 ( 94 0 ) capacitor c=0.0137055f //x=10.805 //y=1.375
c260 ( 92 0 ) capacitor c=0.0149861f //x=10.805 //y=0.72
c261 ( 91 0 ) capacitor c=0.0970408f //x=10.43 //y=1.915
c262 ( 90 0 ) capacitor c=0.0229444f //x=10.43 //y=1.53
c263 ( 89 0 ) capacitor c=0.0234352f //x=10.43 //y=1.22
c264 ( 88 0 ) capacitor c=0.0198724f //x=10.43 //y=0.875
c265 ( 84 0 ) capacitor c=0.0556143f //x=6.195 //y=4.79
c266 ( 83 0 ) capacitor c=0.0293157f //x=6.485 //y=4.79
c267 ( 82 0 ) capacitor c=0.0347816f //x=6.15 //y=1.22
c268 ( 81 0 ) capacitor c=0.0187487f //x=6.15 //y=0.875
c269 ( 75 0 ) capacitor c=0.0137055f //x=5.995 //y=1.375
c270 ( 73 0 ) capacitor c=0.0149861f //x=5.995 //y=0.72
c271 ( 72 0 ) capacitor c=0.0970408f //x=5.62 //y=1.915
c272 ( 71 0 ) capacitor c=0.0229444f //x=5.62 //y=1.53
c273 ( 70 0 ) capacitor c=0.0234352f //x=5.62 //y=1.22
c274 ( 69 0 ) capacitor c=0.0198724f //x=5.62 //y=0.875
c275 ( 68 0 ) capacitor c=0.110114f //x=11.37 //y=6.02
c276 ( 67 0 ) capacitor c=0.158956f //x=10.93 //y=6.02
c277 ( 66 0 ) capacitor c=0.110114f //x=6.56 //y=6.02
c278 ( 65 0 ) capacitor c=0.158956f //x=6.12 //y=6.02
c279 ( 62 0 ) capacitor c=0.00106608f //x=3.29 //y=5.155
c280 ( 61 0 ) capacitor c=0.00207162f //x=2.41 //y=5.155
c281 ( 54 0 ) capacitor c=0.0985621f //x=10.73 //y=2.08
c282 ( 46 0 ) capacitor c=0.104473f //x=5.92 //y=2.08
c283 ( 44 0 ) capacitor c=0.112493f //x=4.07 //y=2.965
c284 ( 40 0 ) capacitor c=0.0052078f //x=3.67 //y=1.665
c285 ( 39 0 ) capacitor c=0.0156949f //x=3.985 //y=1.665
c286 ( 33 0 ) capacitor c=0.0283082f //x=3.985 //y=5.155
c287 ( 25 0 ) capacitor c=0.0176454f //x=3.205 //y=5.155
c288 ( 18 0 ) capacitor c=0.00549987f //x=1.615 //y=5.155
c289 ( 17 0 ) capacitor c=0.020471f //x=2.325 //y=5.155
c290 ( 4 0 ) capacitor c=0.0060653f //x=6.035 //y=2.965
c291 ( 3 0 ) capacitor c=0.134092f //x=10.615 //y=2.965
c292 ( 2 0 ) capacitor c=0.0148225f //x=4.185 //y=2.965
c293 ( 1 0 ) capacitor c=0.0552687f //x=5.805 //y=2.965
r294 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=11.295 //y=4.79 //x2=11.37 //y2=4.865
r295 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=11.295 //y=4.79 //x2=11.005 //y2=4.79
r296 (  101 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.96 //y=1.22 //x2=10.92 //y2=1.375
r297 (  100 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.96 //y=0.875 //x2=10.92 //y2=0.72
r298 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.96 //y=0.875 //x2=10.96 //y2=1.22
r299 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.93 //y=4.865 //x2=11.005 //y2=4.79
r300 (  97 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=10.93 //y=4.865 //x2=10.73 //y2=4.7
r301 (  95 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.585 //y=1.375 //x2=10.47 //y2=1.375
r302 (  94 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.805 //y=1.375 //x2=10.92 //y2=1.375
r303 (  93 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.585 //y=0.72 //x2=10.47 //y2=0.72
r304 (  92 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.805 //y=0.72 //x2=10.92 //y2=0.72
r305 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.805 //y=0.72 //x2=10.585 //y2=0.72
r306 (  91 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.915 //x2=10.73 //y2=2.08
r307 (  90 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.53 //x2=10.47 //y2=1.375
r308 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.53 //x2=10.43 //y2=1.915
r309 (  89 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.22 //x2=10.47 //y2=1.375
r310 (  88 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.43 //y=0.875 //x2=10.47 //y2=0.72
r311 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.43 //y=0.875 //x2=10.43 //y2=1.22
r312 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.485 //y=4.79 //x2=6.56 //y2=4.865
r313 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=6.485 //y=4.79 //x2=6.195 //y2=4.79
r314 (  82 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.15 //y=1.22 //x2=6.11 //y2=1.375
r315 (  81 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.15 //y=0.875 //x2=6.11 //y2=0.72
r316 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.15 //y=0.875 //x2=6.15 //y2=1.22
r317 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.12 //y=4.865 //x2=6.195 //y2=4.79
r318 (  78 112 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=6.12 //y=4.865 //x2=5.92 //y2=4.7
r319 (  76 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.775 //y=1.375 //x2=5.66 //y2=1.375
r320 (  75 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.995 //y=1.375 //x2=6.11 //y2=1.375
r321 (  74 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.775 //y=0.72 //x2=5.66 //y2=0.72
r322 (  73 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.995 //y=0.72 //x2=6.11 //y2=0.72
r323 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=5.995 //y=0.72 //x2=5.775 //y2=0.72
r324 (  72 110 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.915 //x2=5.92 //y2=2.08
r325 (  71 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.53 //x2=5.66 //y2=1.375
r326 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.53 //x2=5.62 //y2=1.915
r327 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.22 //x2=5.66 //y2=1.375
r328 (  69 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=0.875 //x2=5.66 //y2=0.72
r329 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.62 //y=0.875 //x2=5.62 //y2=1.22
r330 (  68 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.37 //y=6.02 //x2=11.37 //y2=4.865
r331 (  67 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.93 //y=6.02 //x2=10.93 //y2=4.865
r332 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.56 //y=6.02 //x2=6.56 //y2=4.865
r333 (  65 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.12 //y=6.02 //x2=6.12 //y2=4.865
r334 (  64 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.695 //y=1.375 //x2=10.805 //y2=1.375
r335 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.695 //y=1.375 //x2=10.585 //y2=1.375
r336 (  63 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.375 //x2=5.995 //y2=1.375
r337 (  63 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.375 //x2=5.775 //y2=1.375
r338 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=4.7 //x2=10.73 //y2=4.7
r339 (  57 59 ) resistor r=118.759 //w=0.187 //l=1.735 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.965 //x2=10.73 //y2=4.7
r340 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=2.08 //x2=10.73 //y2=2.08
r341 (  54 57 ) resistor r=60.5775 //w=0.187 //l=0.885 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.08 //x2=10.73 //y2=2.965
r342 (  51 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=4.7 //x2=5.92 //y2=4.7
r343 (  49 51 ) resistor r=118.759 //w=0.187 //l=1.735 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.965 //x2=5.92 //y2=4.7
r344 (  46 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=2.08 //x2=5.92 //y2=2.08
r345 (  46 49 ) resistor r=60.5775 //w=0.187 //l=0.885 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.08 //x2=5.92 //y2=2.965
r346 (  42 44 ) resistor r=144.086 //w=0.187 //l=2.105 //layer=li \
 //thickness=0.1 //x=4.07 //y=5.07 //x2=4.07 //y2=2.965
r347 (  41 44 ) resistor r=83.1658 //w=0.187 //l=1.215 //layer=li \
 //thickness=0.1 //x=4.07 //y=1.75 //x2=4.07 //y2=2.965
r348 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=4.07 //y2=1.75
r349 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=3.67 //y2=1.665
r350 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.67 //y2=1.665
r351 (  35 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.585 //y2=1.01
r352 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.375 //y=5.155 //x2=3.29 //y2=5.155
r353 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=4.07 //y2=5.07
r354 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=3.375 //y2=5.155
r355 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.155
r356 (  27 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.725
r357 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.495 //y=5.155 //x2=2.41 //y2=5.155
r358 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=3.29 //y2=5.155
r359 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=2.495 //y2=5.155
r360 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.155
r361 (  19 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.725
r362 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=2.41 //y2=5.155
r363 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=1.615 //y2=5.155
r364 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.615 //y2=5.155
r365 (  11 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.53 //y2=5.725
r366 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.73 //y=2.965 //x2=10.73 //y2=2.965
r367 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.92 //y=2.965 //x2=5.92 //y2=2.965
r368 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=2.965 //x2=4.07 //y2=2.965
r369 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.035 //y=2.965 //x2=5.92 //y2=2.965
r370 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=2.965 //x2=10.73 //y2=2.965
r371 (  3 4 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=2.965 //x2=6.035 //y2=2.965
r372 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.185 //y=2.965 //x2=4.07 //y2=2.965
r373 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.805 //y=2.965 //x2=5.92 //y2=2.965
r374 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=5.805 //y=2.965 //x2=4.185 //y2=2.965
ends PM_DFFSNRNX1\%noxref_3

subckt PM_DFFSNRNX1\%noxref_4 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 54 \
 55 56 57 58 60 66 67 68 69 81 83 84 85 )
c160 ( 85 0 ) capacitor c=0.023087f //x=12.765 //y=5.02
c161 ( 84 0 ) capacitor c=0.023519f //x=11.885 //y=5.02
c162 ( 83 0 ) capacitor c=0.0224735f //x=11.005 //y=5.02
c163 ( 81 0 ) capacitor c=0.00853354f //x=13.015 //y=0.915
c164 ( 69 0 ) capacitor c=0.0556143f //x=15.815 //y=4.79
c165 ( 68 0 ) capacitor c=0.0293157f //x=16.105 //y=4.79
c166 ( 67 0 ) capacitor c=0.0347816f //x=15.77 //y=1.22
c167 ( 66 0 ) capacitor c=0.0187487f //x=15.77 //y=0.875
c168 ( 60 0 ) capacitor c=0.0137055f //x=15.615 //y=1.375
c169 ( 58 0 ) capacitor c=0.0149861f //x=15.615 //y=0.72
c170 ( 57 0 ) capacitor c=0.0965296f //x=15.24 //y=1.915
c171 ( 56 0 ) capacitor c=0.0229444f //x=15.24 //y=1.53
c172 ( 55 0 ) capacitor c=0.0234352f //x=15.24 //y=1.22
c173 ( 54 0 ) capacitor c=0.0198724f //x=15.24 //y=0.875
c174 ( 53 0 ) capacitor c=0.110114f //x=16.18 //y=6.02
c175 ( 52 0 ) capacitor c=0.158956f //x=15.74 //y=6.02
c176 ( 50 0 ) capacitor c=0.00106608f //x=12.91 //y=5.155
c177 ( 49 0 ) capacitor c=0.00207319f //x=12.03 //y=5.155
c178 ( 42 0 ) capacitor c=0.0961606f //x=15.54 //y=2.08
c179 ( 40 0 ) capacitor c=0.105233f //x=13.69 //y=2.96
c180 ( 36 0 ) capacitor c=0.00431225f //x=13.29 //y=1.665
c181 ( 35 0 ) capacitor c=0.0143009f //x=13.605 //y=1.665
c182 ( 29 0 ) capacitor c=0.0283082f //x=13.605 //y=5.155
c183 ( 21 0 ) capacitor c=0.0176454f //x=12.825 //y=5.155
c184 ( 14 0 ) capacitor c=0.00332903f //x=11.235 //y=5.155
c185 ( 13 0 ) capacitor c=0.0148427f //x=11.945 //y=5.155
c186 ( 2 0 ) capacitor c=0.00858068f //x=13.805 //y=2.96
c187 ( 1 0 ) capacitor c=0.0396798f //x=15.425 //y=2.96
r188 (  68 70 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=16.105 //y=4.79 //x2=16.18 //y2=4.865
r189 (  68 69 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=16.105 //y=4.79 //x2=15.815 //y2=4.79
r190 (  67 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.77 //y=1.22 //x2=15.73 //y2=1.375
r191 (  66 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.77 //y=0.875 //x2=15.73 //y2=0.72
r192 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.77 //y=0.875 //x2=15.77 //y2=1.22
r193 (  63 69 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.74 //y=4.865 //x2=15.815 //y2=4.79
r194 (  63 78 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=15.74 //y=4.865 //x2=15.54 //y2=4.7
r195 (  61 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.395 //y=1.375 //x2=15.28 //y2=1.375
r196 (  60 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.615 //y=1.375 //x2=15.73 //y2=1.375
r197 (  59 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.395 //y=0.72 //x2=15.28 //y2=0.72
r198 (  58 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.615 //y=0.72 //x2=15.73 //y2=0.72
r199 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=15.615 //y=0.72 //x2=15.395 //y2=0.72
r200 (  57 76 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.915 //x2=15.54 //y2=2.08
r201 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.53 //x2=15.28 //y2=1.375
r202 (  56 57 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.53 //x2=15.24 //y2=1.915
r203 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.22 //x2=15.28 //y2=1.375
r204 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.24 //y=0.875 //x2=15.28 //y2=0.72
r205 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.24 //y=0.875 //x2=15.24 //y2=1.22
r206 (  53 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.18 //y=6.02 //x2=16.18 //y2=4.865
r207 (  52 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.74 //y=6.02 //x2=15.74 //y2=4.865
r208 (  51 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.505 //y=1.375 //x2=15.615 //y2=1.375
r209 (  51 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.505 //y=1.375 //x2=15.395 //y2=1.375
r210 (  47 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.54 //y=4.7 //x2=15.54 //y2=4.7
r211 (  45 47 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=15.54 //y=2.96 //x2=15.54 //y2=4.7
r212 (  42 76 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.54 //y=2.08 //x2=15.54 //y2=2.08
r213 (  42 45 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=15.54 //y=2.08 //x2=15.54 //y2=2.96
r214 (  38 40 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=13.69 //y=5.07 //x2=13.69 //y2=2.96
r215 (  37 40 ) resistor r=82.8235 //w=0.187 //l=1.21 //layer=li \
 //thickness=0.1 //x=13.69 //y=1.75 //x2=13.69 //y2=2.96
r216 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.605 //y=1.665 //x2=13.69 //y2=1.75
r217 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=13.605 //y=1.665 //x2=13.29 //y2=1.665
r218 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.205 //y=1.58 //x2=13.29 //y2=1.665
r219 (  31 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=13.205 //y=1.58 //x2=13.205 //y2=1.01
r220 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.995 //y=5.155 //x2=12.91 //y2=5.155
r221 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.605 //y=5.155 //x2=13.69 //y2=5.07
r222 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=13.605 //y=5.155 //x2=12.995 //y2=5.155
r223 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.91 //y=5.24 //x2=12.91 //y2=5.155
r224 (  23 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.91 //y=5.24 //x2=12.91 //y2=5.725
r225 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.115 //y=5.155 //x2=12.03 //y2=5.155
r226 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.825 //y=5.155 //x2=12.91 //y2=5.155
r227 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=12.825 //y=5.155 //x2=12.115 //y2=5.155
r228 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.03 //y=5.24 //x2=12.03 //y2=5.155
r229 (  15 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.03 //y=5.24 //x2=12.03 //y2=5.725
r230 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.945 //y=5.155 //x2=12.03 //y2=5.155
r231 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.945 //y=5.155 //x2=11.235 //y2=5.155
r232 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.15 //y=5.24 //x2=11.235 //y2=5.155
r233 (  7 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.15 //y=5.24 //x2=11.15 //y2=5.725
r234 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.54 //y=2.96 //x2=15.54 //y2=2.96
r235 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=13.69 //y=2.96 //x2=13.69 //y2=2.96
r236 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.805 //y=2.96 //x2=13.69 //y2=2.96
r237 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.425 //y=2.96 //x2=15.54 //y2=2.96
r238 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=15.425 //y=2.96 //x2=13.805 //y2=2.96
ends PM_DFFSNRNX1\%noxref_4

subckt PM_DFFSNRNX1\%CLK ( 1 2 7 8 9 10 11 13 23 31 32 33 34 35 36 37 38 39 41 \
 47 48 49 50 51 56 57 58 60 66 67 68 69 70 78 89 )
c191 ( 89 0 ) capacitor c=0.0337106f //x=16.65 //y=4.7
c192 ( 78 0 ) capacitor c=0.0335551f //x=7.03 //y=4.7
c193 ( 70 0 ) capacitor c=0.0245352f //x=16.985 //y=4.79
c194 ( 69 0 ) capacitor c=0.0826403f //x=16.74 //y=1.915
c195 ( 68 0 ) capacitor c=0.0170266f //x=16.74 //y=1.45
c196 ( 67 0 ) capacitor c=0.018609f //x=16.74 //y=1.22
c197 ( 66 0 ) capacitor c=0.0187309f //x=16.74 //y=0.91
c198 ( 60 0 ) capacitor c=0.014725f //x=16.585 //y=1.375
c199 ( 58 0 ) capacitor c=0.0146567f //x=16.585 //y=0.755
c200 ( 57 0 ) capacitor c=0.0335408f //x=16.215 //y=1.22
c201 ( 56 0 ) capacitor c=0.0173761f //x=16.215 //y=0.91
c202 ( 51 0 ) capacitor c=0.0245352f //x=7.365 //y=4.79
c203 ( 50 0 ) capacitor c=0.0828223f //x=7.12 //y=1.915
c204 ( 49 0 ) capacitor c=0.0170266f //x=7.12 //y=1.45
c205 ( 48 0 ) capacitor c=0.018609f //x=7.12 //y=1.22
c206 ( 47 0 ) capacitor c=0.0187309f //x=7.12 //y=0.91
c207 ( 41 0 ) capacitor c=0.014725f //x=6.965 //y=1.375
c208 ( 39 0 ) capacitor c=0.0146567f //x=6.965 //y=0.755
c209 ( 38 0 ) capacitor c=0.0335408f //x=6.595 //y=1.22
c210 ( 37 0 ) capacitor c=0.0173761f //x=6.595 //y=0.91
c211 ( 36 0 ) capacitor c=0.110114f //x=17.06 //y=6.02
c212 ( 35 0 ) capacitor c=0.11012f //x=16.62 //y=6.02
c213 ( 34 0 ) capacitor c=0.110114f //x=7.44 //y=6.02
c214 ( 33 0 ) capacitor c=0.11012f //x=7 //y=6.02
c215 ( 23 0 ) capacitor c=0.0926339f //x=16.65 //y=2.08
c216 ( 13 0 ) capacitor c=0.0951886f //x=7.03 //y=2.08
c217 ( 2 0 ) capacitor c=0.0137564f //x=7.145 //y=3.33
c218 ( 1 0 ) capacitor c=0.169502f //x=16.535 //y=3.33
r219 (  91 92 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=16.65 //y=4.79 //x2=16.65 //y2=4.865
r220 (  89 91 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=16.65 //y=4.7 //x2=16.65 //y2=4.79
r221 (  80 81 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=7.03 //y=4.79 //x2=7.03 //y2=4.865
r222 (  78 80 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=7.03 //y=4.7 //x2=7.03 //y2=4.79
r223 (  71 91 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=16.785 //y=4.79 //x2=16.65 //y2=4.79
r224 (  70 72 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=16.985 //y=4.79 //x2=17.06 //y2=4.865
r225 (  70 71 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=16.985 //y=4.79 //x2=16.785 //y2=4.79
r226 (  69 96 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.915 //x2=16.665 //y2=2.08
r227 (  68 94 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.45 //x2=16.7 //y2=1.375
r228 (  68 69 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.45 //x2=16.74 //y2=1.915
r229 (  67 94 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.22 //x2=16.7 //y2=1.375
r230 (  66 93 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.74 //y=0.91 //x2=16.7 //y2=0.755
r231 (  66 67 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=16.74 //y=0.91 //x2=16.74 //y2=1.22
r232 (  61 87 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.37 //y=1.375 //x2=16.255 //y2=1.375
r233 (  60 94 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.585 //y=1.375 //x2=16.7 //y2=1.375
r234 (  59 86 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.37 //y=0.755 //x2=16.255 //y2=0.755
r235 (  58 93 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.585 //y=0.755 //x2=16.7 //y2=0.755
r236 (  58 59 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=16.585 //y=0.755 //x2=16.37 //y2=0.755
r237 (  57 87 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.215 //y=1.22 //x2=16.255 //y2=1.375
r238 (  56 86 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.215 //y=0.91 //x2=16.255 //y2=0.755
r239 (  56 57 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=16.215 //y=0.91 //x2=16.215 //y2=1.22
r240 (  52 80 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=7.165 //y=4.79 //x2=7.03 //y2=4.79
r241 (  51 53 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.365 //y=4.79 //x2=7.44 //y2=4.865
r242 (  51 52 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=7.365 //y=4.79 //x2=7.165 //y2=4.79
r243 (  50 85 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.915 //x2=7.045 //y2=2.08
r244 (  49 83 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.45 //x2=7.08 //y2=1.375
r245 (  49 50 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.45 //x2=7.12 //y2=1.915
r246 (  48 83 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.22 //x2=7.08 //y2=1.375
r247 (  47 82 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.12 //y=0.91 //x2=7.08 //y2=0.755
r248 (  47 48 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=7.12 //y=0.91 //x2=7.12 //y2=1.22
r249 (  42 76 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.75 //y=1.375 //x2=6.635 //y2=1.375
r250 (  41 83 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.965 //y=1.375 //x2=7.08 //y2=1.375
r251 (  40 75 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.75 //y=0.755 //x2=6.635 //y2=0.755
r252 (  39 82 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.965 //y=0.755 //x2=7.08 //y2=0.755
r253 (  39 40 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=6.965 //y=0.755 //x2=6.75 //y2=0.755
r254 (  38 76 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.595 //y=1.22 //x2=6.635 //y2=1.375
r255 (  37 75 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.595 //y=0.91 //x2=6.635 //y2=0.755
r256 (  37 38 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=6.595 //y=0.91 //x2=6.595 //y2=1.22
r257 (  36 72 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.06 //y=6.02 //x2=17.06 //y2=4.865
r258 (  35 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.62 //y=6.02 //x2=16.62 //y2=4.865
r259 (  34 53 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.44 //y=6.02 //x2=7.44 //y2=4.865
r260 (  33 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7 //y=6.02 //x2=7 //y2=4.865
r261 (  32 60 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=16.477 //y=1.375 //x2=16.585 //y2=1.375
r262 (  32 61 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=16.477 //y=1.375 //x2=16.37 //y2=1.375
r263 (  31 41 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=6.857 //y=1.375 //x2=6.965 //y2=1.375
r264 (  31 42 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=6.857 //y=1.375 //x2=6.75 //y2=1.375
r265 (  29 89 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.65 //y=4.7 //x2=16.65 //y2=4.7
r266 (  23 96 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.65 //y=2.08 //x2=16.65 //y2=2.08
r267 (  20 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.03 //y=4.7 //x2=7.03 //y2=4.7
r268 (  13 85 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.03 //y=2.08 //x2=7.03 //y2=2.08
r269 (  11 29 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=16.65 //y=3.33 //x2=16.65 //y2=4.7
r270 (  10 11 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=16.65 //y=2.96 //x2=16.65 //y2=3.33
r271 (  10 23 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=16.65 //y=2.96 //x2=16.65 //y2=2.08
r272 (  9 20 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li //thickness=0.1 \
 //x=7.03 //y=4.07 //x2=7.03 //y2=4.7
r273 (  8 9 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li //thickness=0.1 \
 //x=7.03 //y=3.33 //x2=7.03 //y2=4.07
r274 (  7 8 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li //thickness=0.1 \
 //x=7.03 //y=2.59 //x2=7.03 //y2=3.33
r275 (  7 13 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=7.03 //y=2.59 //x2=7.03 //y2=2.08
r276 (  6 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=16.65 //y=3.33 //x2=16.65 //y2=3.33
r277 (  4 8 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=7.03 \
 //y=3.33 //x2=7.03 //y2=3.33
r278 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.145 //y=3.33 //x2=7.03 //y2=3.33
r279 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.535 //y=3.33 //x2=16.65 //y2=3.33
r280 (  1 2 ) resistor r=8.95992 //w=0.131 //l=9.39 //layer=m1 \
 //thickness=0.36 //x=16.535 //y=3.33 //x2=7.145 //y2=3.33
ends PM_DFFSNRNX1\%CLK

subckt PM_DFFSNRNX1\%noxref_6 ( 1 2 3 4 12 25 26 33 41 47 48 52 54 61 62 63 64 \
 65 66 67 68 72 73 74 79 81 84 85 86 87 88 89 90 92 98 99 100 101 106 107 112 \
 123 125 126 127 )
c261 ( 127 0 ) capacitor c=0.023087f //x=7.955 //y=5.02
c262 ( 126 0 ) capacitor c=0.023519f //x=7.075 //y=5.02
c263 ( 125 0 ) capacitor c=0.0224735f //x=6.195 //y=5.02
c264 ( 123 0 ) capacitor c=0.00853354f //x=8.205 //y=0.915
c265 ( 112 0 ) capacitor c=0.058931f //x=3.33 //y=4.7
c266 ( 107 0 ) capacitor c=0.0273931f //x=3.33 //y=1.915
c267 ( 106 0 ) capacitor c=0.0471168f //x=3.33 //y=2.08
c268 ( 101 0 ) capacitor c=0.0556143f //x=20.625 //y=4.79
c269 ( 100 0 ) capacitor c=0.0293157f //x=20.915 //y=4.79
c270 ( 99 0 ) capacitor c=0.0347816f //x=20.58 //y=1.22
c271 ( 98 0 ) capacitor c=0.0187487f //x=20.58 //y=0.875
c272 ( 92 0 ) capacitor c=0.0137055f //x=20.425 //y=1.375
c273 ( 90 0 ) capacitor c=0.0149861f //x=20.425 //y=0.72
c274 ( 89 0 ) capacitor c=0.0965296f //x=20.05 //y=1.915
c275 ( 88 0 ) capacitor c=0.0229444f //x=20.05 //y=1.53
c276 ( 87 0 ) capacitor c=0.0234352f //x=20.05 //y=1.22
c277 ( 86 0 ) capacitor c=0.0198724f //x=20.05 //y=0.875
c278 ( 85 0 ) capacitor c=0.0432517f //x=3.85 //y=1.26
c279 ( 84 0 ) capacitor c=0.0200379f //x=3.85 //y=0.915
c280 ( 81 0 ) capacitor c=0.0158629f //x=3.695 //y=1.415
c281 ( 79 0 ) capacitor c=0.0157803f //x=3.695 //y=0.76
c282 ( 74 0 ) capacitor c=0.0218028f //x=3.32 //y=1.57
c283 ( 73 0 ) capacitor c=0.0207459f //x=3.32 //y=1.26
c284 ( 72 0 ) capacitor c=0.0194308f //x=3.32 //y=0.915
c285 ( 68 0 ) capacitor c=0.110114f //x=20.99 //y=6.02
c286 ( 67 0 ) capacitor c=0.158956f //x=20.55 //y=6.02
c287 ( 66 0 ) capacitor c=0.158794f //x=3.51 //y=6.02
c288 ( 65 0 ) capacitor c=0.110114f //x=3.07 //y=6.02
c289 ( 62 0 ) capacitor c=0.00104281f //x=8.1 //y=5.155
c290 ( 61 0 ) capacitor c=0.00207319f //x=7.22 //y=5.155
c291 ( 54 0 ) capacitor c=0.103455f //x=20.35 //y=2.08
c292 ( 52 0 ) capacitor c=0.10634f //x=8.88 //y=3.7
c293 ( 48 0 ) capacitor c=0.00463944f //x=8.48 //y=1.665
c294 ( 47 0 ) capacitor c=0.0148811f //x=8.795 //y=1.665
c295 ( 41 0 ) capacitor c=0.0283082f //x=8.795 //y=5.155
c296 ( 33 0 ) capacitor c=0.0176454f //x=8.015 //y=5.155
c297 ( 26 0 ) capacitor c=0.00332903f //x=6.425 //y=5.155
c298 ( 25 0 ) capacitor c=0.0148427f //x=7.135 //y=5.155
c299 ( 12 0 ) capacitor c=0.09073f //x=3.33 //y=2.08
c300 ( 4 0 ) capacitor c=0.0055354f //x=8.995 //y=3.7
c301 ( 3 0 ) capacitor c=0.195503f //x=20.235 //y=3.7
c302 ( 2 0 ) capacitor c=0.0166717f //x=3.445 //y=3.7
c303 ( 1 0 ) capacitor c=0.107088f //x=8.765 //y=3.7
r304 (  106 107 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.33 //y=2.08 //x2=3.33 //y2=1.915
r305 (  100 102 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.915 //y=4.79 //x2=20.99 //y2=4.865
r306 (  100 101 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=20.915 //y=4.79 //x2=20.625 //y2=4.79
r307 (  99 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.58 //y=1.22 //x2=20.54 //y2=1.375
r308 (  98 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.58 //y=0.875 //x2=20.54 //y2=0.72
r309 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.58 //y=0.875 //x2=20.58 //y2=1.22
r310 (  95 101 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.55 //y=4.865 //x2=20.625 //y2=4.79
r311 (  95 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=20.55 //y=4.865 //x2=20.35 //y2=4.7
r312 (  93 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.205 //y=1.375 //x2=20.09 //y2=1.375
r313 (  92 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.425 //y=1.375 //x2=20.54 //y2=1.375
r314 (  91 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.205 //y=0.72 //x2=20.09 //y2=0.72
r315 (  90 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.425 //y=0.72 //x2=20.54 //y2=0.72
r316 (  90 91 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=20.425 //y=0.72 //x2=20.205 //y2=0.72
r317 (  89 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.915 //x2=20.35 //y2=2.08
r318 (  88 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.53 //x2=20.09 //y2=1.375
r319 (  88 89 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.53 //x2=20.05 //y2=1.915
r320 (  87 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.22 //x2=20.09 //y2=1.375
r321 (  86 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.05 //y=0.875 //x2=20.09 //y2=0.72
r322 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.05 //y=0.875 //x2=20.05 //y2=1.22
r323 (  85 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=1.26 //x2=3.81 //y2=1.415
r324 (  84 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.81 //y2=0.76
r325 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.85 //y2=1.26
r326 (  82 110 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=1.415 //x2=3.36 //y2=1.415
r327 (  81 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=1.415 //x2=3.81 //y2=1.415
r328 (  80 109 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=0.76 //x2=3.36 //y2=0.76
r329 (  79 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.81 //y2=0.76
r330 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.475 //y2=0.76
r331 (  76 112 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=3.51 //y=4.865 //x2=3.33 //y2=4.7
r332 (  74 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.36 //y2=1.415
r333 (  74 107 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.32 //y2=1.915
r334 (  73 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.26 //x2=3.36 //y2=1.415
r335 (  72 109 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.36 //y2=0.76
r336 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.32 //y2=1.26
r337 (  69 112 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=3.07 //y=4.865 //x2=3.33 //y2=4.7
r338 (  68 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.99 //y=6.02 //x2=20.99 //y2=4.865
r339 (  67 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.55 //y=6.02 //x2=20.55 //y2=4.865
r340 (  66 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.51 //y=6.02 //x2=3.51 //y2=4.865
r341 (  65 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.07 //y=6.02 //x2=3.07 //y2=4.865
r342 (  64 92 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.315 //y=1.375 //x2=20.425 //y2=1.375
r343 (  64 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.315 //y=1.375 //x2=20.205 //y2=1.375
r344 (  63 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.695 //y2=1.415
r345 (  63 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.475 //y2=1.415
r346 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.35 //y=4.7 //x2=20.35 //y2=4.7
r347 (  57 59 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=20.35 //y=3.7 //x2=20.35 //y2=4.7
r348 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.35 //y=2.08 //x2=20.35 //y2=2.08
r349 (  54 57 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=20.35 //y=2.08 //x2=20.35 //y2=3.7
r350 (  50 52 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=8.88 //y=5.07 //x2=8.88 //y2=3.7
r351 (  49 52 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=8.88 //y=1.75 //x2=8.88 //y2=3.7
r352 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.795 //y=1.665 //x2=8.88 //y2=1.75
r353 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=8.795 //y=1.665 //x2=8.48 //y2=1.665
r354 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.395 //y=1.58 //x2=8.48 //y2=1.665
r355 (  43 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=8.395 //y=1.58 //x2=8.395 //y2=1.01
r356 (  42 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.185 //y=5.155 //x2=8.1 //y2=5.155
r357 (  41 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.795 //y=5.155 //x2=8.88 //y2=5.07
r358 (  41 42 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=8.795 //y=5.155 //x2=8.185 //y2=5.155
r359 (  35 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.1 //y=5.24 //x2=8.1 //y2=5.155
r360 (  35 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.1 //y=5.24 //x2=8.1 //y2=5.725
r361 (  34 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.305 //y=5.155 //x2=7.22 //y2=5.155
r362 (  33 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.015 //y=5.155 //x2=8.1 //y2=5.155
r363 (  33 34 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.015 //y=5.155 //x2=7.305 //y2=5.155
r364 (  27 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.24 //x2=7.22 //y2=5.155
r365 (  27 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.24 //x2=7.22 //y2=5.725
r366 (  25 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.155 //x2=7.22 //y2=5.155
r367 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.155 //x2=6.425 //y2=5.155
r368 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.24 //x2=6.425 //y2=5.155
r369 (  19 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.24 //x2=6.34 //y2=5.725
r370 (  17 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r371 (  15 17 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=3.33 //y=3.7 //x2=3.33 //y2=4.7
r372 (  12 106 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r373 (  12 15 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.08 //x2=3.33 //y2=3.7
r374 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=20.35 //y=3.7 //x2=20.35 //y2=3.7
r375 (  8 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.88 //y=3.7 //x2=8.88 //y2=3.7
r376 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=3.7 //x2=3.33 //y2=3.7
r377 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.995 //y=3.7 //x2=8.88 //y2=3.7
r378 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.235 //y=3.7 //x2=20.35 //y2=3.7
r379 (  3 4 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=20.235 //y=3.7 //x2=8.995 //y2=3.7
r380 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.445 //y=3.7 //x2=3.33 //y2=3.7
r381 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=3.7 //x2=8.88 //y2=3.7
r382 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=3.7 //x2=3.445 //y2=3.7
ends PM_DFFSNRNX1\%noxref_6

subckt PM_DFFSNRNX1\%RN ( 1 2 3 4 11 12 13 14 15 16 17 18 19 20 21 22 23 25 38 \
 48 58 59 60 61 62 63 64 65 66 67 68 69 71 77 78 79 80 81 89 90 91 96 98 101 \
 102 103 104 105 107 113 114 115 116 117 125 134 135 140 146 )
c309 ( 146 0 ) capacitor c=0.0334842f //x=21.46 //y=4.7
c310 ( 140 0 ) capacitor c=0.0587051f //x=17.76 //y=4.7
c311 ( 135 0 ) capacitor c=0.0273931f //x=17.76 //y=1.915
c312 ( 134 0 ) capacitor c=0.0457054f //x=17.76 //y=2.08
c313 ( 125 0 ) capacitor c=0.0334842f //x=2.22 //y=4.7
c314 ( 117 0 ) capacitor c=0.0249231f //x=21.795 //y=4.79
c315 ( 116 0 ) capacitor c=0.0826403f //x=21.55 //y=1.915
c316 ( 115 0 ) capacitor c=0.0170266f //x=21.55 //y=1.45
c317 ( 114 0 ) capacitor c=0.018609f //x=21.55 //y=1.22
c318 ( 113 0 ) capacitor c=0.0187309f //x=21.55 //y=0.91
c319 ( 107 0 ) capacitor c=0.014725f //x=21.395 //y=1.375
c320 ( 105 0 ) capacitor c=0.0146567f //x=21.395 //y=0.755
c321 ( 104 0 ) capacitor c=0.0335408f //x=21.025 //y=1.22
c322 ( 103 0 ) capacitor c=0.0173761f //x=21.025 //y=0.91
c323 ( 102 0 ) capacitor c=0.0432517f //x=18.28 //y=1.26
c324 ( 101 0 ) capacitor c=0.0200379f //x=18.28 //y=0.915
c325 ( 98 0 ) capacitor c=0.0158629f //x=18.125 //y=1.415
c326 ( 96 0 ) capacitor c=0.0157803f //x=18.125 //y=0.76
c327 ( 91 0 ) capacitor c=0.0218028f //x=17.75 //y=1.57
c328 ( 90 0 ) capacitor c=0.0207459f //x=17.75 //y=1.26
c329 ( 89 0 ) capacitor c=0.0194308f //x=17.75 //y=0.915
c330 ( 81 0 ) capacitor c=0.0245352f //x=2.555 //y=4.79
c331 ( 80 0 ) capacitor c=0.0850619f //x=2.31 //y=1.915
c332 ( 79 0 ) capacitor c=0.0170266f //x=2.31 //y=1.45
c333 ( 78 0 ) capacitor c=0.018609f //x=2.31 //y=1.22
c334 ( 77 0 ) capacitor c=0.0187309f //x=2.31 //y=0.91
c335 ( 71 0 ) capacitor c=0.014725f //x=2.155 //y=1.375
c336 ( 69 0 ) capacitor c=0.0146567f //x=2.155 //y=0.755
c337 ( 68 0 ) capacitor c=0.0335408f //x=1.785 //y=1.22
c338 ( 67 0 ) capacitor c=0.0173761f //x=1.785 //y=0.91
c339 ( 66 0 ) capacitor c=0.110114f //x=21.87 //y=6.02
c340 ( 65 0 ) capacitor c=0.11012f //x=21.43 //y=6.02
c341 ( 64 0 ) capacitor c=0.158794f //x=17.94 //y=6.02
c342 ( 63 0 ) capacitor c=0.110114f //x=17.5 //y=6.02
c343 ( 62 0 ) capacitor c=0.110114f //x=2.63 //y=6.02
c344 ( 61 0 ) capacitor c=0.11012f //x=2.19 //y=6.02
c345 ( 48 0 ) capacitor c=0.0968545f //x=21.46 //y=2.08
c346 ( 38 0 ) capacitor c=0.0856807f //x=17.76 //y=2.08
c347 ( 25 0 ) capacitor c=0.103016f //x=2.22 //y=2.08
c348 ( 4 0 ) capacitor c=0.00565359f //x=17.875 //y=4.44
c349 ( 3 0 ) capacitor c=0.0960334f //x=21.345 //y=4.44
c350 ( 2 0 ) capacitor c=0.0175929f //x=2.335 //y=4.44
c351 ( 1 0 ) capacitor c=0.377168f //x=17.645 //y=4.44
r352 (  148 149 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=21.46 //y=4.79 //x2=21.46 //y2=4.865
r353 (  146 148 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=21.46 //y=4.7 //x2=21.46 //y2=4.79
r354 (  134 135 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=17.76 //y=2.08 //x2=17.76 //y2=1.915
r355 (  127 128 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.79 //x2=2.22 //y2=4.865
r356 (  125 127 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.7 //x2=2.22 //y2=4.79
r357 (  118 148 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=21.595 //y=4.79 //x2=21.46 //y2=4.79
r358 (  117 119 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=21.795 //y=4.79 //x2=21.87 //y2=4.865
r359 (  117 118 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=21.795 //y=4.79 //x2=21.595 //y2=4.79
r360 (  116 153 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.915 //x2=21.475 //y2=2.08
r361 (  115 151 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.45 //x2=21.51 //y2=1.375
r362 (  115 116 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.45 //x2=21.55 //y2=1.915
r363 (  114 151 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.22 //x2=21.51 //y2=1.375
r364 (  113 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.55 //y=0.91 //x2=21.51 //y2=0.755
r365 (  113 114 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.55 //y=0.91 //x2=21.55 //y2=1.22
r366 (  108 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.18 //y=1.375 //x2=21.065 //y2=1.375
r367 (  107 151 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.395 //y=1.375 //x2=21.51 //y2=1.375
r368 (  106 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.18 //y=0.755 //x2=21.065 //y2=0.755
r369 (  105 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.755 //x2=21.51 //y2=0.755
r370 (  105 106 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.755 //x2=21.18 //y2=0.755
r371 (  104 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.025 //y=1.22 //x2=21.065 //y2=1.375
r372 (  103 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.025 //y=0.91 //x2=21.065 //y2=0.755
r373 (  103 104 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.025 //y=0.91 //x2=21.025 //y2=1.22
r374 (  102 142 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.28 //y=1.26 //x2=18.24 //y2=1.415
r375 (  101 141 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.28 //y=0.915 //x2=18.24 //y2=0.76
r376 (  101 102 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.28 //y=0.915 //x2=18.28 //y2=1.26
r377 (  99 138 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.905 //y=1.415 //x2=17.79 //y2=1.415
r378 (  98 142 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.125 //y=1.415 //x2=18.24 //y2=1.415
r379 (  97 137 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.905 //y=0.76 //x2=17.79 //y2=0.76
r380 (  96 141 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.125 //y=0.76 //x2=18.24 //y2=0.76
r381 (  96 97 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=18.125 //y=0.76 //x2=17.905 //y2=0.76
r382 (  93 140 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=17.94 //y=4.865 //x2=17.76 //y2=4.7
r383 (  91 138 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.75 //y=1.57 //x2=17.79 //y2=1.415
r384 (  91 135 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.75 //y=1.57 //x2=17.75 //y2=1.915
r385 (  90 138 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.75 //y=1.26 //x2=17.79 //y2=1.415
r386 (  89 137 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.75 //y=0.915 //x2=17.79 //y2=0.76
r387 (  89 90 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.75 //y=0.915 //x2=17.75 //y2=1.26
r388 (  86 140 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=17.5 //y=4.865 //x2=17.76 //y2=4.7
r389 (  82 127 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.355 //y=4.79 //x2=2.22 //y2=4.79
r390 (  81 83 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.63 //y2=4.865
r391 (  81 82 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.355 //y2=4.79
r392 (  80 132 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.915 //x2=2.235 //y2=2.08
r393 (  79 130 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.27 //y2=1.375
r394 (  79 80 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.31 //y2=1.915
r395 (  78 130 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.22 //x2=2.27 //y2=1.375
r396 (  77 129 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.27 //y2=0.755
r397 (  77 78 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.31 //y2=1.22
r398 (  72 123 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=1.375 //x2=1.825 //y2=1.375
r399 (  71 130 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=1.375 //x2=2.27 //y2=1.375
r400 (  70 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=0.755 //x2=1.825 //y2=0.755
r401 (  69 129 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=2.27 //y2=0.755
r402 (  69 70 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=1.94 //y2=0.755
r403 (  68 123 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=1.22 //x2=1.825 //y2=1.375
r404 (  67 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.825 //y2=0.755
r405 (  67 68 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.785 //y2=1.22
r406 (  66 119 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.87 //y=6.02 //x2=21.87 //y2=4.865
r407 (  65 149 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.43 //y=6.02 //x2=21.43 //y2=4.865
r408 (  64 93 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.94 //y=6.02 //x2=17.94 //y2=4.865
r409 (  63 86 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.5 //y=6.02 //x2=17.5 //y2=4.865
r410 (  62 83 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.63 //y=6.02 //x2=2.63 //y2=4.865
r411 (  61 128 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.19 //y=6.02 //x2=2.19 //y2=4.865
r412 (  60 107 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=21.287 //y=1.375 //x2=21.395 //y2=1.375
r413 (  60 108 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=21.287 //y=1.375 //x2=21.18 //y2=1.375
r414 (  59 98 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.015 //y=1.415 //x2=18.125 //y2=1.415
r415 (  59 99 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.015 //y=1.415 //x2=17.905 //y2=1.415
r416 (  58 71 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=2.155 //y2=1.375
r417 (  58 72 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=1.94 //y2=1.375
r418 (  56 146 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.46 //y=4.7 //x2=21.46 //y2=4.7
r419 (  48 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.46 //y=2.08 //x2=21.46 //y2=2.08
r420 (  45 140 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.76 //y=4.7 //x2=17.76 //y2=4.7
r421 (  38 134 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.76 //y=2.08 //x2=17.76 //y2=2.08
r422 (  35 125 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=4.7 //x2=2.22 //y2=4.7
r423 (  25 132 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=2.08
r424 (  23 56 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=21.46 //y=4.44 //x2=21.46 //y2=4.7
r425 (  22 23 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=21.46 //y=3.7 //x2=21.46 //y2=4.44
r426 (  21 22 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.46 //y=3.33 //x2=21.46 //y2=3.7
r427 (  20 21 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.96 //x2=21.46 //y2=3.33
r428 (  20 48 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.96 //x2=21.46 //y2=2.08
r429 (  19 45 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=17.76 //y=4.44 //x2=17.76 //y2=4.7
r430 (  18 19 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=17.76 //y=3.33 //x2=17.76 //y2=4.44
r431 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.96 //x2=17.76 //y2=3.33
r432 (  17 38 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.96 //x2=17.76 //y2=2.08
r433 (  16 35 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=2.22 //y=4.44 //x2=2.22 //y2=4.7
r434 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=4.07 //x2=2.22 //y2=4.44
r435 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.7 //x2=2.22 //y2=4.07
r436 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.33 //x2=2.22 //y2=3.7
r437 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.96 //x2=2.22 //y2=3.33
r438 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.59 //x2=2.22 //y2=2.96
r439 (  11 25 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.59 //x2=2.22 //y2=2.08
r440 (  10 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.46 //y=4.44 //x2=21.46 //y2=4.44
r441 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.76 //y=4.44 //x2=17.76 //y2=4.44
r442 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.22 //y=4.44 //x2=2.22 //y2=4.44
r443 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.875 //y=4.44 //x2=17.76 //y2=4.44
r444 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=4.44 //x2=21.46 //y2=4.44
r445 (  3 4 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=4.44 //x2=17.875 //y2=4.44
r446 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.335 //y=4.44 //x2=2.22 //y2=4.44
r447 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.645 //y=4.44 //x2=17.76 //y2=4.44
r448 (  1 2 ) resistor r=14.6088 //w=0.131 //l=15.31 //layer=m1 \
 //thickness=0.36 //x=17.645 //y=4.44 //x2=2.335 //y2=4.44
ends PM_DFFSNRNX1\%RN

subckt PM_DFFSNRNX1\%QN ( 1 2 7 8 9 10 11 12 13 14 21 22 29 37 43 44 53 63 64 \
 65 66 67 68 69 70 71 72 74 80 81 82 83 95 97 98 99 )
c157 ( 99 0 ) capacitor c=0.023087f //x=22.385 //y=5.02
c158 ( 98 0 ) capacitor c=0.023519f //x=21.505 //y=5.02
c159 ( 97 0 ) capacitor c=0.0224735f //x=20.625 //y=5.02
c160 ( 95 0 ) capacitor c=0.00853354f //x=22.635 //y=0.915
c161 ( 83 0 ) capacitor c=0.0558396f //x=25.435 //y=4.79
c162 ( 82 0 ) capacitor c=0.0298189f //x=25.725 //y=4.79
c163 ( 81 0 ) capacitor c=0.0347816f //x=25.39 //y=1.22
c164 ( 80 0 ) capacitor c=0.0187487f //x=25.39 //y=0.875
c165 ( 74 0 ) capacitor c=0.0137055f //x=25.235 //y=1.375
c166 ( 72 0 ) capacitor c=0.0149861f //x=25.235 //y=0.72
c167 ( 71 0 ) capacitor c=0.0965296f //x=24.86 //y=1.915
c168 ( 70 0 ) capacitor c=0.0229444f //x=24.86 //y=1.53
c169 ( 69 0 ) capacitor c=0.0234352f //x=24.86 //y=1.22
c170 ( 68 0 ) capacitor c=0.0198724f //x=24.86 //y=0.875
c171 ( 67 0 ) capacitor c=0.110114f //x=25.8 //y=6.02
c172 ( 66 0 ) capacitor c=0.158956f //x=25.36 //y=6.02
c173 ( 64 0 ) capacitor c=0.00116729f //x=22.53 //y=5.155
c174 ( 63 0 ) capacitor c=0.0021933f //x=21.65 //y=5.155
c175 ( 53 0 ) capacitor c=0.102092f //x=25.16 //y=2.08
c176 ( 44 0 ) capacitor c=0.00431225f //x=22.91 //y=1.665
c177 ( 43 0 ) capacitor c=0.0143009f //x=23.225 //y=1.665
c178 ( 37 0 ) capacitor c=0.0291119f //x=23.225 //y=5.155
c179 ( 29 0 ) capacitor c=0.0184197f //x=22.445 //y=5.155
c180 ( 22 0 ) capacitor c=0.00332903f //x=20.855 //y=5.155
c181 ( 21 0 ) capacitor c=0.014837f //x=21.565 //y=5.155
c182 ( 7 0 ) capacitor c=0.109457f //x=23.31 //y=2.22
c183 ( 2 0 ) capacitor c=0.0124102f //x=23.425 //y=3.33
c184 ( 1 0 ) capacitor c=0.0456899f //x=25.045 //y=3.33
r185 (  82 84 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=25.725 //y=4.79 //x2=25.8 //y2=4.865
r186 (  82 83 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=25.725 //y=4.79 //x2=25.435 //y2=4.79
r187 (  81 94 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.39 //y=1.22 //x2=25.35 //y2=1.375
r188 (  80 93 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.39 //y=0.875 //x2=25.35 //y2=0.72
r189 (  80 81 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=25.39 //y=0.875 //x2=25.39 //y2=1.22
r190 (  77 83 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=25.36 //y=4.865 //x2=25.435 //y2=4.79
r191 (  77 92 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=25.36 //y=4.865 //x2=25.16 //y2=4.7
r192 (  75 88 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.015 //y=1.375 //x2=24.9 //y2=1.375
r193 (  74 94 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.235 //y=1.375 //x2=25.35 //y2=1.375
r194 (  73 87 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.015 //y=0.72 //x2=24.9 //y2=0.72
r195 (  72 93 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.235 //y=0.72 //x2=25.35 //y2=0.72
r196 (  72 73 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=25.235 //y=0.72 //x2=25.015 //y2=0.72
r197 (  71 90 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.915 //x2=25.16 //y2=2.08
r198 (  70 88 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.53 //x2=24.9 //y2=1.375
r199 (  70 71 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.53 //x2=24.86 //y2=1.915
r200 (  69 88 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.22 //x2=24.9 //y2=1.375
r201 (  68 87 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.86 //y=0.875 //x2=24.9 //y2=0.72
r202 (  68 69 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.86 //y=0.875 //x2=24.86 //y2=1.22
r203 (  67 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=25.8 //y=6.02 //x2=25.8 //y2=4.865
r204 (  66 77 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=25.36 //y=6.02 //x2=25.36 //y2=4.865
r205 (  65 74 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.125 //y=1.375 //x2=25.235 //y2=1.375
r206 (  65 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.125 //y=1.375 //x2=25.015 //y2=1.375
r207 (  61 92 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=25.16 //y=4.7 //x2=25.16 //y2=4.7
r208 (  53 90 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=25.16 //y=2.08 //x2=25.16 //y2=2.08
r209 (  43 45 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.225 //y=1.665 //x2=23.31 //y2=1.75
r210 (  43 44 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=23.225 //y=1.665 //x2=22.91 //y2=1.665
r211 (  39 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=22.825 //y=1.58 //x2=22.91 //y2=1.665
r212 (  39 95 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=22.825 //y=1.58 //x2=22.825 //y2=1.01
r213 (  38 64 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.615 //y=5.155 //x2=22.53 //y2=5.155
r214 (  37 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.225 //y=5.155 //x2=23.31 //y2=5.07
r215 (  37 38 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=23.225 //y=5.155 //x2=22.615 //y2=5.155
r216 (  31 64 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.53 //y=5.24 //x2=22.53 //y2=5.155
r217 (  31 99 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.53 //y=5.24 //x2=22.53 //y2=5.725
r218 (  30 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.735 //y=5.155 //x2=21.65 //y2=5.155
r219 (  29 64 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.445 //y=5.155 //x2=22.53 //y2=5.155
r220 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.445 //y=5.155 //x2=21.735 //y2=5.155
r221 (  23 63 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.65 //y=5.24 //x2=21.65 //y2=5.155
r222 (  23 98 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.65 //y=5.24 //x2=21.65 //y2=5.725
r223 (  21 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.565 //y=5.155 //x2=21.65 //y2=5.155
r224 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=21.565 //y=5.155 //x2=20.855 //y2=5.155
r225 (  15 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.77 //y=5.24 //x2=20.855 //y2=5.155
r226 (  15 97 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.77 //y=5.24 //x2=20.77 //y2=5.725
r227 (  14 61 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=25.16 //y=4.44 //x2=25.16 //y2=4.7
r228 (  13 14 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=25.16 //y=3.33 //x2=25.16 //y2=4.44
r229 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=25.16 //y=2.96 //x2=25.16 //y2=3.33
r230 (  11 12 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=25.16 //y=2.22 //x2=25.16 //y2=2.96
r231 (  11 53 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=25.16 //y=2.22 //x2=25.16 //y2=2.08
r232 (  10 46 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=23.31 //y=4.44 //x2=23.31 //y2=5.07
r233 (  9 10 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=23.31 //y=3.33 //x2=23.31 //y2=4.44
r234 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=23.31 //y=2.96 //x2=23.31 //y2=3.33
r235 (  7 8 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li //thickness=0.1 \
 //x=23.31 //y=2.22 //x2=23.31 //y2=2.96
r236 (  7 45 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=23.31 //y=2.22 //x2=23.31 //y2=1.75
r237 (  6 13 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=25.16 //y=3.33 //x2=25.16 //y2=3.33
r238 (  4 9 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=23.31 //y=3.33 //x2=23.31 //y2=3.33
r239 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.425 //y=3.33 //x2=23.31 //y2=3.33
r240 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=25.045 //y=3.33 //x2=25.16 //y2=3.33
r241 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=25.045 //y=3.33 //x2=23.425 //y2=3.33
ends PM_DFFSNRNX1\%QN

subckt PM_DFFSNRNX1\%SN ( 1 2 7 8 9 10 11 12 14 23 33 34 35 36 37 38 39 40 41 \
 43 49 50 51 52 53 58 59 60 62 68 69 70 71 72 80 91 )
c229 ( 91 0 ) capacitor c=0.0336203f //x=26.27 //y=4.7
c230 ( 80 0 ) capacitor c=0.0335551f //x=11.84 //y=4.7
c231 ( 72 0 ) capacitor c=0.024933f //x=26.605 //y=4.79
c232 ( 71 0 ) capacitor c=0.0830584f //x=26.36 //y=1.915
c233 ( 70 0 ) capacitor c=0.0170266f //x=26.36 //y=1.45
c234 ( 69 0 ) capacitor c=0.018609f //x=26.36 //y=1.22
c235 ( 68 0 ) capacitor c=0.0187309f //x=26.36 //y=0.91
c236 ( 62 0 ) capacitor c=0.014725f //x=26.205 //y=1.375
c237 ( 60 0 ) capacitor c=0.0146567f //x=26.205 //y=0.755
c238 ( 59 0 ) capacitor c=0.0335408f //x=25.835 //y=1.22
c239 ( 58 0 ) capacitor c=0.0173761f //x=25.835 //y=0.91
c240 ( 53 0 ) capacitor c=0.0245352f //x=12.175 //y=4.79
c241 ( 52 0 ) capacitor c=0.0826363f //x=11.93 //y=1.915
c242 ( 51 0 ) capacitor c=0.0170266f //x=11.93 //y=1.45
c243 ( 50 0 ) capacitor c=0.018609f //x=11.93 //y=1.22
c244 ( 49 0 ) capacitor c=0.0187309f //x=11.93 //y=0.91
c245 ( 43 0 ) capacitor c=0.014725f //x=11.775 //y=1.375
c246 ( 41 0 ) capacitor c=0.0146567f //x=11.775 //y=0.755
c247 ( 40 0 ) capacitor c=0.0335408f //x=11.405 //y=1.22
c248 ( 39 0 ) capacitor c=0.0173761f //x=11.405 //y=0.91
c249 ( 38 0 ) capacitor c=0.110114f //x=26.68 //y=6.02
c250 ( 37 0 ) capacitor c=0.11012f //x=26.24 //y=6.02
c251 ( 36 0 ) capacitor c=0.110114f //x=12.25 //y=6.02
c252 ( 35 0 ) capacitor c=0.11012f //x=11.81 //y=6.02
c253 ( 23 0 ) capacitor c=0.0978636f //x=26.27 //y=2.08
c254 ( 14 0 ) capacitor c=0.0922012f //x=11.84 //y=2.08
c255 ( 2 0 ) capacitor c=0.0159757f //x=11.955 //y=2.59
c256 ( 1 0 ) capacitor c=0.395426f //x=26.155 //y=2.59
r257 (  93 94 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=26.27 //y=4.79 //x2=26.27 //y2=4.865
r258 (  91 93 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=26.27 //y=4.7 //x2=26.27 //y2=4.79
r259 (  82 83 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=11.84 //y=4.79 //x2=11.84 //y2=4.865
r260 (  80 82 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=11.84 //y=4.7 //x2=11.84 //y2=4.79
r261 (  73 93 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=26.405 //y=4.79 //x2=26.27 //y2=4.79
r262 (  72 74 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=26.605 //y=4.79 //x2=26.68 //y2=4.865
r263 (  72 73 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=26.605 //y=4.79 //x2=26.405 //y2=4.79
r264 (  71 98 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.915 //x2=26.285 //y2=2.08
r265 (  70 96 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.45 //x2=26.32 //y2=1.375
r266 (  70 71 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.45 //x2=26.36 //y2=1.915
r267 (  69 96 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.22 //x2=26.32 //y2=1.375
r268 (  68 95 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.36 //y=0.91 //x2=26.32 //y2=0.755
r269 (  68 69 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=26.36 //y=0.91 //x2=26.36 //y2=1.22
r270 (  63 89 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.99 //y=1.375 //x2=25.875 //y2=1.375
r271 (  62 96 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.205 //y=1.375 //x2=26.32 //y2=1.375
r272 (  61 88 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.99 //y=0.755 //x2=25.875 //y2=0.755
r273 (  60 95 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.205 //y=0.755 //x2=26.32 //y2=0.755
r274 (  60 61 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=26.205 //y=0.755 //x2=25.99 //y2=0.755
r275 (  59 89 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.835 //y=1.22 //x2=25.875 //y2=1.375
r276 (  58 88 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.835 //y=0.91 //x2=25.875 //y2=0.755
r277 (  58 59 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=25.835 //y=0.91 //x2=25.835 //y2=1.22
r278 (  54 82 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=11.975 //y=4.79 //x2=11.84 //y2=4.79
r279 (  53 55 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=12.175 //y=4.79 //x2=12.25 //y2=4.865
r280 (  53 54 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=12.175 //y=4.79 //x2=11.975 //y2=4.79
r281 (  52 87 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.915 //x2=11.855 //y2=2.08
r282 (  51 85 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.45 //x2=11.89 //y2=1.375
r283 (  51 52 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.45 //x2=11.93 //y2=1.915
r284 (  50 85 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.22 //x2=11.89 //y2=1.375
r285 (  49 84 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.93 //y=0.91 //x2=11.89 //y2=0.755
r286 (  49 50 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=11.93 //y=0.91 //x2=11.93 //y2=1.22
r287 (  44 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.56 //y=1.375 //x2=11.445 //y2=1.375
r288 (  43 85 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.775 //y=1.375 //x2=11.89 //y2=1.375
r289 (  42 77 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.56 //y=0.755 //x2=11.445 //y2=0.755
r290 (  41 84 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.775 //y=0.755 //x2=11.89 //y2=0.755
r291 (  41 42 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=11.775 //y=0.755 //x2=11.56 //y2=0.755
r292 (  40 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.405 //y=1.22 //x2=11.445 //y2=1.375
r293 (  39 77 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.405 //y=0.91 //x2=11.445 //y2=0.755
r294 (  39 40 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=11.405 //y=0.91 //x2=11.405 //y2=1.22
r295 (  38 74 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.68 //y=6.02 //x2=26.68 //y2=4.865
r296 (  37 94 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.24 //y=6.02 //x2=26.24 //y2=4.865
r297 (  36 55 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.25 //y=6.02 //x2=12.25 //y2=4.865
r298 (  35 83 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.81 //y=6.02 //x2=11.81 //y2=4.865
r299 (  34 62 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=26.097 //y=1.375 //x2=26.205 //y2=1.375
r300 (  34 63 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=26.097 //y=1.375 //x2=25.99 //y2=1.375
r301 (  33 43 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=11.667 //y=1.375 //x2=11.775 //y2=1.375
r302 (  33 44 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=11.667 //y=1.375 //x2=11.56 //y2=1.375
r303 (  31 91 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.27 //y=4.7 //x2=26.27 //y2=4.7
r304 (  23 98 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.27 //y=2.08 //x2=26.27 //y2=2.08
r305 (  20 80 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=4.7 //x2=11.84 //y2=4.7
r306 (  14 87 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=2.08 //x2=11.84 //y2=2.08
r307 (  12 31 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=26.27 //y=4.44 //x2=26.27 //y2=4.7
r308 (  11 12 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=26.27 //y=3.33 //x2=26.27 //y2=4.44
r309 (  10 11 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.96 //x2=26.27 //y2=3.33
r310 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.59 //x2=26.27 //y2=2.96
r311 (  9 23 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.59 //x2=26.27 //y2=2.08
r312 (  8 20 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.96 //x2=11.84 //y2=4.7
r313 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=11.84 //y=2.59 //x2=11.84 //y2=2.96
r314 (  7 14 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.59 //x2=11.84 //y2=2.08
r315 (  6 9 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=26.27 //y=2.59 //x2=26.27 //y2=2.59
r316 (  4 7 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.84 //y=2.59 //x2=11.84 //y2=2.59
r317 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.955 //y=2.59 //x2=11.84 //y2=2.59
r318 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=26.155 //y=2.59 //x2=26.27 //y2=2.59
r319 (  1 2 ) resistor r=13.5496 //w=0.131 //l=14.2 //layer=m1 \
 //thickness=0.36 //x=26.155 //y=2.59 //x2=11.955 //y2=2.59
ends PM_DFFSNRNX1\%SN

subckt PM_DFFSNRNX1\%noxref_10 ( 1 2 3 4 5 6 17 21 24 37 38 45 53 59 60 64 66 \
 74 77 78 79 80 81 82 83 84 85 86 87 91 92 93 98 100 103 104 108 109 110 115 \
 117 120 121 125 126 127 132 134 137 138 140 141 146 150 151 156 160 161 166 \
 169 171 172 173 )
c340 ( 173 0 ) capacitor c=0.023087f //x=17.575 //y=5.02
c341 ( 172 0 ) capacitor c=0.023519f //x=16.695 //y=5.02
c342 ( 171 0 ) capacitor c=0.0224735f //x=15.815 //y=5.02
c343 ( 169 0 ) capacitor c=0.00853354f //x=17.825 //y=0.915
c344 ( 166 0 ) capacitor c=0.0593979f //x=27.38 //y=4.7
c345 ( 161 0 ) capacitor c=0.0273931f //x=27.38 //y=1.915
c346 ( 160 0 ) capacitor c=0.0471168f //x=27.38 //y=2.08
c347 ( 156 0 ) capacitor c=0.0587755f //x=12.95 //y=4.7
c348 ( 151 0 ) capacitor c=0.0273931f //x=12.95 //y=1.915
c349 ( 150 0 ) capacitor c=0.0457054f //x=12.95 //y=2.08
c350 ( 146 0 ) capacitor c=0.0587602f //x=8.14 //y=4.7
c351 ( 141 0 ) capacitor c=0.0273931f //x=8.14 //y=1.915
c352 ( 140 0 ) capacitor c=0.0458344f //x=8.14 //y=2.08
c353 ( 138 0 ) capacitor c=0.0432517f //x=27.9 //y=1.26
c354 ( 137 0 ) capacitor c=0.0200379f //x=27.9 //y=0.915
c355 ( 134 0 ) capacitor c=0.0158629f //x=27.745 //y=1.415
c356 ( 132 0 ) capacitor c=0.0157803f //x=27.745 //y=0.76
c357 ( 127 0 ) capacitor c=0.0218028f //x=27.37 //y=1.57
c358 ( 126 0 ) capacitor c=0.0207459f //x=27.37 //y=1.26
c359 ( 125 0 ) capacitor c=0.0194308f //x=27.37 //y=0.915
c360 ( 121 0 ) capacitor c=0.0432517f //x=13.47 //y=1.26
c361 ( 120 0 ) capacitor c=0.0200379f //x=13.47 //y=0.915
c362 ( 117 0 ) capacitor c=0.0158629f //x=13.315 //y=1.415
c363 ( 115 0 ) capacitor c=0.0157803f //x=13.315 //y=0.76
c364 ( 110 0 ) capacitor c=0.0218028f //x=12.94 //y=1.57
c365 ( 109 0 ) capacitor c=0.0207459f //x=12.94 //y=1.26
c366 ( 108 0 ) capacitor c=0.0194308f //x=12.94 //y=0.915
c367 ( 104 0 ) capacitor c=0.0432517f //x=8.66 //y=1.26
c368 ( 103 0 ) capacitor c=0.0200379f //x=8.66 //y=0.915
c369 ( 100 0 ) capacitor c=0.0158629f //x=8.505 //y=1.415
c370 ( 98 0 ) capacitor c=0.0157803f //x=8.505 //y=0.76
c371 ( 93 0 ) capacitor c=0.0218028f //x=8.13 //y=1.57
c372 ( 92 0 ) capacitor c=0.0207459f //x=8.13 //y=1.26
c373 ( 91 0 ) capacitor c=0.0194308f //x=8.13 //y=0.915
c374 ( 87 0 ) capacitor c=0.158794f //x=27.56 //y=6.02
c375 ( 86 0 ) capacitor c=0.110114f //x=27.12 //y=6.02
c376 ( 85 0 ) capacitor c=0.158794f //x=13.13 //y=6.02
c377 ( 84 0 ) capacitor c=0.110114f //x=12.69 //y=6.02
c378 ( 83 0 ) capacitor c=0.158794f //x=8.32 //y=6.02
c379 ( 82 0 ) capacitor c=0.110114f //x=7.88 //y=6.02
c380 ( 78 0 ) capacitor c=0.00105927f //x=17.72 //y=5.155
c381 ( 77 0 ) capacitor c=0.00207319f //x=16.84 //y=5.155
c382 ( 74 0 ) capacitor c=0.0105673f //x=8.135 //y=4.07
c383 ( 66 0 ) capacitor c=0.090362f //x=27.38 //y=2.08
c384 ( 64 0 ) capacitor c=0.110121f //x=18.5 //y=4.07
c385 ( 60 0 ) capacitor c=0.00431225f //x=18.1 //y=1.665
c386 ( 59 0 ) capacitor c=0.0143009f //x=18.415 //y=1.665
c387 ( 53 0 ) capacitor c=0.0283032f //x=18.415 //y=5.155
c388 ( 45 0 ) capacitor c=0.0176454f //x=17.635 //y=5.155
c389 ( 38 0 ) capacitor c=0.00332903f //x=16.045 //y=5.155
c390 ( 37 0 ) capacitor c=0.0148427f //x=16.755 //y=5.155
c391 ( 24 0 ) capacitor c=0.0833947f //x=12.95 //y=2.08
c392 ( 21 0 ) capacitor c=0.0129218f //x=8.14 //y=4.7
c393 ( 17 0 ) capacitor c=0.0610714f //x=8.14 //y=2.08
c394 ( 6 0 ) capacitor c=0.00554824f //x=18.615 //y=4.07
c395 ( 5 0 ) capacitor c=0.218272f //x=27.265 //y=4.07
c396 ( 4 0 ) capacitor c=0.00562383f //x=13.065 //y=4.07
c397 ( 3 0 ) capacitor c=0.0724583f //x=18.385 //y=4.07
c398 ( 2 0 ) capacitor c=0.0138844f //x=8.25 //y=4.07
c399 ( 1 0 ) capacitor c=0.0638764f //x=12.835 //y=4.07
r400 (  160 161 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=27.38 //y=2.08 //x2=27.38 //y2=1.915
r401 (  150 151 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=12.95 //y=2.08 //x2=12.95 //y2=1.915
r402 (  140 141 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=8.14 //y=2.08 //x2=8.14 //y2=1.915
r403 (  138 168 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.9 //y=1.26 //x2=27.86 //y2=1.415
r404 (  137 167 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.9 //y=0.915 //x2=27.86 //y2=0.76
r405 (  137 138 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.9 //y=0.915 //x2=27.9 //y2=1.26
r406 (  135 164 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.525 //y=1.415 //x2=27.41 //y2=1.415
r407 (  134 168 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.745 //y=1.415 //x2=27.86 //y2=1.415
r408 (  133 163 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.525 //y=0.76 //x2=27.41 //y2=0.76
r409 (  132 167 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.745 //y=0.76 //x2=27.86 //y2=0.76
r410 (  132 133 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=27.745 //y=0.76 //x2=27.525 //y2=0.76
r411 (  129 166 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=27.56 //y=4.865 //x2=27.38 //y2=4.7
r412 (  127 164 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.37 //y=1.57 //x2=27.41 //y2=1.415
r413 (  127 161 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.37 //y=1.57 //x2=27.37 //y2=1.915
r414 (  126 164 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.37 //y=1.26 //x2=27.41 //y2=1.415
r415 (  125 163 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.37 //y=0.915 //x2=27.41 //y2=0.76
r416 (  125 126 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.37 //y=0.915 //x2=27.37 //y2=1.26
r417 (  122 166 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=27.12 //y=4.865 //x2=27.38 //y2=4.7
r418 (  121 158 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.47 //y=1.26 //x2=13.43 //y2=1.415
r419 (  120 157 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.47 //y=0.915 //x2=13.43 //y2=0.76
r420 (  120 121 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.47 //y=0.915 //x2=13.47 //y2=1.26
r421 (  118 154 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.095 //y=1.415 //x2=12.98 //y2=1.415
r422 (  117 158 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.315 //y=1.415 //x2=13.43 //y2=1.415
r423 (  116 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.095 //y=0.76 //x2=12.98 //y2=0.76
r424 (  115 157 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.315 //y=0.76 //x2=13.43 //y2=0.76
r425 (  115 116 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=13.315 //y=0.76 //x2=13.095 //y2=0.76
r426 (  112 156 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=13.13 //y=4.865 //x2=12.95 //y2=4.7
r427 (  110 154 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.94 //y=1.57 //x2=12.98 //y2=1.415
r428 (  110 151 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.94 //y=1.57 //x2=12.94 //y2=1.915
r429 (  109 154 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.94 //y=1.26 //x2=12.98 //y2=1.415
r430 (  108 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.94 //y=0.915 //x2=12.98 //y2=0.76
r431 (  108 109 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.94 //y=0.915 //x2=12.94 //y2=1.26
r432 (  105 156 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=12.69 //y=4.865 //x2=12.95 //y2=4.7
r433 (  104 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.66 //y=1.26 //x2=8.62 //y2=1.415
r434 (  103 147 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.66 //y=0.915 //x2=8.62 //y2=0.76
r435 (  103 104 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.66 //y=0.915 //x2=8.66 //y2=1.26
r436 (  101 144 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.285 //y=1.415 //x2=8.17 //y2=1.415
r437 (  100 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.505 //y=1.415 //x2=8.62 //y2=1.415
r438 (  99 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.285 //y=0.76 //x2=8.17 //y2=0.76
r439 (  98 147 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.505 //y=0.76 //x2=8.62 //y2=0.76
r440 (  98 99 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=8.505 //y=0.76 //x2=8.285 //y2=0.76
r441 (  95 146 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=8.32 //y=4.865 //x2=8.14 //y2=4.7
r442 (  93 144 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.57 //x2=8.17 //y2=1.415
r443 (  93 141 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.57 //x2=8.13 //y2=1.915
r444 (  92 144 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.26 //x2=8.17 //y2=1.415
r445 (  91 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=0.915 //x2=8.17 //y2=0.76
r446 (  91 92 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.13 //y=0.915 //x2=8.13 //y2=1.26
r447 (  88 146 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=7.88 //y=4.865 //x2=8.14 //y2=4.7
r448 (  87 129 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=27.56 //y=6.02 //x2=27.56 //y2=4.865
r449 (  86 122 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=27.12 //y=6.02 //x2=27.12 //y2=4.865
r450 (  85 112 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.13 //y=6.02 //x2=13.13 //y2=4.865
r451 (  84 105 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.69 //y=6.02 //x2=12.69 //y2=4.865
r452 (  83 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.32 //y=6.02 //x2=8.32 //y2=4.865
r453 (  82 88 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.88 //y=6.02 //x2=7.88 //y2=4.865
r454 (  81 134 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=27.635 //y=1.415 //x2=27.745 //y2=1.415
r455 (  81 135 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=27.635 //y=1.415 //x2=27.525 //y2=1.415
r456 (  80 117 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.205 //y=1.415 //x2=13.315 //y2=1.415
r457 (  80 118 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.205 //y=1.415 //x2=13.095 //y2=1.415
r458 (  79 100 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.395 //y=1.415 //x2=8.505 //y2=1.415
r459 (  79 101 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.395 //y=1.415 //x2=8.285 //y2=1.415
r460 (  74 76 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=8.137 //y=4.07 //x2=8.137 //y2=4.235
r461 (  74 75 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=8.137 //y=4.07 //x2=8.137 //y2=3.905
r462 (  71 166 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=27.38 //y=4.7 //x2=27.38 //y2=4.7
r463 (  69 71 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=27.38 //y=4.07 //x2=27.38 //y2=4.7
r464 (  66 160 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=27.38 //y=2.08 //x2=27.38 //y2=2.08
r465 (  66 69 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=27.38 //y=2.08 //x2=27.38 //y2=4.07
r466 (  62 64 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=18.5 //y=5.07 //x2=18.5 //y2=4.07
r467 (  61 64 ) resistor r=158.802 //w=0.187 //l=2.32 //layer=li \
 //thickness=0.1 //x=18.5 //y=1.75 //x2=18.5 //y2=4.07
r468 (  59 61 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.415 //y=1.665 //x2=18.5 //y2=1.75
r469 (  59 60 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=18.415 //y=1.665 //x2=18.1 //y2=1.665
r470 (  55 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.015 //y=1.58 //x2=18.1 //y2=1.665
r471 (  55 169 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=18.015 //y=1.58 //x2=18.015 //y2=1.01
r472 (  54 78 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.805 //y=5.155 //x2=17.72 //y2=5.155
r473 (  53 62 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.415 //y=5.155 //x2=18.5 //y2=5.07
r474 (  53 54 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=18.415 //y=5.155 //x2=17.805 //y2=5.155
r475 (  47 78 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.72 //y=5.24 //x2=17.72 //y2=5.155
r476 (  47 173 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.72 //y=5.24 //x2=17.72 //y2=5.725
r477 (  46 77 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.925 //y=5.155 //x2=16.84 //y2=5.155
r478 (  45 78 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.635 //y=5.155 //x2=17.72 //y2=5.155
r479 (  45 46 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=17.635 //y=5.155 //x2=16.925 //y2=5.155
r480 (  39 77 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.84 //y=5.24 //x2=16.84 //y2=5.155
r481 (  39 172 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.84 //y=5.24 //x2=16.84 //y2=5.725
r482 (  37 77 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.755 //y=5.155 //x2=16.84 //y2=5.155
r483 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=16.755 //y=5.155 //x2=16.045 //y2=5.155
r484 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.96 //y=5.24 //x2=16.045 //y2=5.155
r485 (  31 171 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.96 //y=5.24 //x2=15.96 //y2=5.725
r486 (  29 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.95 //y=4.7 //x2=12.95 //y2=4.7
r487 (  27 29 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=12.95 //y=4.07 //x2=12.95 //y2=4.7
r488 (  24 150 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.95 //y=2.08 //x2=12.95 //y2=2.08
r489 (  24 27 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=12.95 //y=2.08 //x2=12.95 //y2=4.07
r490 (  21 146 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.14 //y=4.7 //x2=8.14 //y2=4.7
r491 (  21 76 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=8.14 //y=4.7 //x2=8.14 //y2=4.235
r492 (  17 140 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.14 //y=2.08 //x2=8.14 //y2=2.08
r493 (  17 75 ) resistor r=124.92 //w=0.187 //l=1.825 //layer=li \
 //thickness=0.1 //x=8.14 //y=2.08 //x2=8.14 //y2=3.905
r494 (  14 69 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=27.38 //y=4.07 //x2=27.38 //y2=4.07
r495 (  12 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.5 //y=4.07 //x2=18.5 //y2=4.07
r496 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.95 //y=4.07 //x2=12.95 //y2=4.07
r497 (  8 74 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.135 //y=4.07 //x2=8.135 //y2=4.07
r498 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.615 //y=4.07 //x2=18.5 //y2=4.07
r499 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=27.265 //y=4.07 //x2=27.38 //y2=4.07
r500 (  5 6 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=27.265 //y=4.07 //x2=18.615 //y2=4.07
r501 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.065 //y=4.07 //x2=12.95 //y2=4.07
r502 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.385 //y=4.07 //x2=18.5 //y2=4.07
r503 (  3 4 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=18.385 //y=4.07 //x2=13.065 //y2=4.07
r504 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.25 //y=4.07 //x2=8.135 //y2=4.07
r505 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.835 //y=4.07 //x2=12.95 //y2=4.07
r506 (  1 2 ) resistor r=4.375 //w=0.131 //l=4.585 //layer=m1 //thickness=0.36 \
 //x=12.835 //y=4.07 //x2=8.25 //y2=4.07
ends PM_DFFSNRNX1\%noxref_10

subckt PM_DFFSNRNX1\%Q ( 1 2 7 8 9 10 11 12 13 14 15 16 17 18 19 21 38 39 46 \
 54 60 61 73 74 75 76 77 81 82 83 88 90 93 94 96 97 102 105 107 108 109 )
c157 ( 109 0 ) capacitor c=0.023087f //x=27.195 //y=5.02
c158 ( 108 0 ) capacitor c=0.023519f //x=26.315 //y=5.02
c159 ( 107 0 ) capacitor c=0.0224735f //x=25.435 //y=5.02
c160 ( 105 0 ) capacitor c=0.00853354f //x=27.445 //y=0.915
c161 ( 102 0 ) capacitor c=0.0593675f //x=22.57 //y=4.7
c162 ( 97 0 ) capacitor c=0.0273931f //x=22.57 //y=1.915
c163 ( 96 0 ) capacitor c=0.0457054f //x=22.57 //y=2.08
c164 ( 94 0 ) capacitor c=0.0432517f //x=23.09 //y=1.26
c165 ( 93 0 ) capacitor c=0.0200379f //x=23.09 //y=0.915
c166 ( 90 0 ) capacitor c=0.0158629f //x=22.935 //y=1.415
c167 ( 88 0 ) capacitor c=0.0157803f //x=22.935 //y=0.76
c168 ( 83 0 ) capacitor c=0.0218028f //x=22.56 //y=1.57
c169 ( 82 0 ) capacitor c=0.0207459f //x=22.56 //y=1.26
c170 ( 81 0 ) capacitor c=0.0194308f //x=22.56 //y=0.915
c171 ( 77 0 ) capacitor c=0.158794f //x=22.75 //y=6.02
c172 ( 76 0 ) capacitor c=0.110114f //x=22.31 //y=6.02
c173 ( 74 0 ) capacitor c=0.00116099f //x=27.34 //y=5.155
c174 ( 73 0 ) capacitor c=0.00226015f //x=26.46 //y=5.155
c175 ( 61 0 ) capacitor c=0.0052078f //x=27.72 //y=1.665
c176 ( 60 0 ) capacitor c=0.0158856f //x=28.035 //y=1.665
c177 ( 54 0 ) capacitor c=0.0297779f //x=28.035 //y=5.155
c178 ( 46 0 ) capacitor c=0.0184197f //x=27.255 //y=5.155
c179 ( 39 0 ) capacitor c=0.00351598f //x=25.665 //y=5.155
c180 ( 38 0 ) capacitor c=0.0155255f //x=26.375 //y=5.155
c181 ( 21 0 ) capacitor c=0.088301f //x=22.57 //y=2.08
c182 ( 12 0 ) capacitor c=0.129879f //x=28.12 //y=2.22
c183 ( 2 0 ) capacitor c=0.00997231f //x=22.685 //y=3.7
c184 ( 1 0 ) capacitor c=0.132281f //x=28.005 //y=3.7
r185 (  96 97 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=22.57 //y=2.08 //x2=22.57 //y2=1.915
r186 (  94 104 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.09 //y=1.26 //x2=23.05 //y2=1.415
r187 (  93 103 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.09 //y=0.915 //x2=23.05 //y2=0.76
r188 (  93 94 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=23.09 //y=0.915 //x2=23.09 //y2=1.26
r189 (  91 100 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.715 //y=1.415 //x2=22.6 //y2=1.415
r190 (  90 104 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.935 //y=1.415 //x2=23.05 //y2=1.415
r191 (  89 99 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.715 //y=0.76 //x2=22.6 //y2=0.76
r192 (  88 103 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.935 //y=0.76 //x2=23.05 //y2=0.76
r193 (  88 89 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=22.935 //y=0.76 //x2=22.715 //y2=0.76
r194 (  85 102 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=22.75 //y=4.865 //x2=22.57 //y2=4.7
r195 (  83 100 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.56 //y=1.57 //x2=22.6 //y2=1.415
r196 (  83 97 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.56 //y=1.57 //x2=22.56 //y2=1.915
r197 (  82 100 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.56 //y=1.26 //x2=22.6 //y2=1.415
r198 (  81 99 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.56 //y=0.915 //x2=22.6 //y2=0.76
r199 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.56 //y=0.915 //x2=22.56 //y2=1.26
r200 (  78 102 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=22.31 //y=4.865 //x2=22.57 //y2=4.7
r201 (  77 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.75 //y=6.02 //x2=22.75 //y2=4.865
r202 (  76 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.31 //y=6.02 //x2=22.31 //y2=4.865
r203 (  75 90 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=22.825 //y=1.415 //x2=22.935 //y2=1.415
r204 (  75 91 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=22.825 //y=1.415 //x2=22.715 //y2=1.415
r205 (  60 62 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=28.035 //y=1.665 //x2=28.12 //y2=1.75
r206 (  60 61 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=28.035 //y=1.665 //x2=27.72 //y2=1.665
r207 (  56 61 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=27.635 //y=1.58 //x2=27.72 //y2=1.665
r208 (  56 105 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=27.635 //y=1.58 //x2=27.635 //y2=1.01
r209 (  55 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.425 //y=5.155 //x2=27.34 //y2=5.155
r210 (  54 63 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=28.035 //y=5.155 //x2=28.12 //y2=5.07
r211 (  54 55 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=28.035 //y=5.155 //x2=27.425 //y2=5.155
r212 (  48 74 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.34 //y=5.24 //x2=27.34 //y2=5.155
r213 (  48 109 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=27.34 //y=5.24 //x2=27.34 //y2=5.725
r214 (  47 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.545 //y=5.155 //x2=26.46 //y2=5.155
r215 (  46 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.255 //y=5.155 //x2=27.34 //y2=5.155
r216 (  46 47 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=27.255 //y=5.155 //x2=26.545 //y2=5.155
r217 (  40 73 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.46 //y=5.24 //x2=26.46 //y2=5.155
r218 (  40 108 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.46 //y=5.24 //x2=26.46 //y2=5.725
r219 (  38 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.375 //y=5.155 //x2=26.46 //y2=5.155
r220 (  38 39 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=26.375 //y=5.155 //x2=25.665 //y2=5.155
r221 (  32 39 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.58 //y=5.24 //x2=25.665 //y2=5.155
r222 (  32 107 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=25.58 //y=5.24 //x2=25.58 //y2=5.725
r223 (  30 102 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.57 //y=4.7 //x2=22.57 //y2=4.7
r224 (  21 96 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.57 //y=2.08 //x2=22.57 //y2=2.08
r225 (  19 63 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=28.12 //y=4.81 //x2=28.12 //y2=5.07
r226 (  18 19 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=28.12 //y=4.44 //x2=28.12 //y2=4.81
r227 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=28.12 //y=4.07 //x2=28.12 //y2=4.44
r228 (  16 17 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=28.12 //y=3.7 //x2=28.12 //y2=4.07
r229 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=28.12 //y=3.33 //x2=28.12 //y2=3.7
r230 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=28.12 //y=2.96 //x2=28.12 //y2=3.33
r231 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=28.12 //y=2.59 //x2=28.12 //y2=2.96
r232 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=28.12 //y=2.22 //x2=28.12 //y2=2.59
r233 (  12 62 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=28.12 //y=2.22 //x2=28.12 //y2=1.75
r234 (  11 30 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=22.57 //y=4.44 //x2=22.57 //y2=4.7
r235 (  10 11 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=22.57 //y=3.7 //x2=22.57 //y2=4.44
r236 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=22.57 //y=3.33 //x2=22.57 //y2=3.7
r237 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=22.57 //y=2.96 //x2=22.57 //y2=3.33
r238 (  7 8 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li //thickness=0.1 \
 //x=22.57 //y=2.22 //x2=22.57 //y2=2.96
r239 (  7 21 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=22.57 //y=2.22 //x2=22.57 //y2=2.08
r240 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=28.12 //y=3.7 //x2=28.12 //y2=3.7
r241 (  4 10 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=22.57 //y=3.7 //x2=22.57 //y2=3.7
r242 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=22.685 //y=3.7 //x2=22.57 //y2=3.7
r243 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=28.005 //y=3.7 //x2=28.12 //y2=3.7
r244 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=28.005 //y=3.7 //x2=22.685 //y2=3.7
ends PM_DFFSNRNX1\%Q

subckt PM_DFFSNRNX1\%D ( 1 2 3 4 5 6 8 19 20 21 22 23 24 25 26 28 34 35 36 37 )
c56 ( 37 0 ) capacitor c=0.06002f //x=1.385 //y=4.79
c57 ( 36 0 ) capacitor c=0.0375015f //x=1.675 //y=4.79
c58 ( 35 0 ) capacitor c=0.0347816f //x=1.34 //y=1.22
c59 ( 34 0 ) capacitor c=0.0187487f //x=1.34 //y=0.875
c60 ( 28 0 ) capacitor c=0.0137055f //x=1.185 //y=1.375
c61 ( 26 0 ) capacitor c=0.0149861f //x=1.185 //y=0.72
c62 ( 25 0 ) capacitor c=0.102158f //x=0.81 //y=1.915
c63 ( 24 0 ) capacitor c=0.0229444f //x=0.81 //y=1.53
c64 ( 23 0 ) capacitor c=0.0234352f //x=0.81 //y=1.22
c65 ( 22 0 ) capacitor c=0.0198724f //x=0.81 //y=0.875
c66 ( 21 0 ) capacitor c=0.110114f //x=1.75 //y=6.02
c67 ( 20 0 ) capacitor c=0.158956f //x=1.31 //y=6.02
c68 ( 8 0 ) capacitor c=0.127598f //x=1.11 //y=2.08
r69 (  36 38 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.75 //y2=4.865
r70 (  36 37 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.385 //y2=4.79
r71 (  35 48 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=1.22 //x2=1.3 //y2=1.375
r72 (  34 47 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.3 //y2=0.72
r73 (  34 35 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.34 //y2=1.22
r74 (  31 37 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.385 //y2=4.79
r75 (  31 46 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.11 //y2=4.7
r76 (  29 42 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=1.375 //x2=0.85 //y2=1.375
r77 (  28 48 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=1.375 //x2=1.3 //y2=1.375
r78 (  27 41 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=0.72 //x2=0.85 //y2=0.72
r79 (  26 47 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=1.3 //y2=0.72
r80 (  26 27 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=0.965 //y2=0.72
r81 (  25 44 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.915 //x2=1.11 //y2=2.08
r82 (  24 42 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.85 //y2=1.375
r83 (  24 25 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.81 //y2=1.915
r84 (  23 42 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.22 //x2=0.85 //y2=1.375
r85 (  22 41 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.85 //y2=0.72
r86 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.81 //y2=1.22
r87 (  21 38 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.75 //y=6.02 //x2=1.75 //y2=4.865
r88 (  20 31 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.31 //y=6.02 //x2=1.31 //y2=4.865
r89 (  19 28 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=1.185 //y2=1.375
r90 (  19 29 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=0.965 //y2=1.375
r91 (  17 46 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r92 (  8 44 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r93 (  6 17 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.44 //x2=1.11 //y2=4.7
r94 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.44
r95 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=3.7 //x2=1.11 //y2=4.07
r96 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=3.33 //x2=1.11 //y2=3.7
r97 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.96 //x2=1.11 //y2=3.33
r98 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.59 //x2=1.11 //y2=2.96
r99 (  1 8 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.59 //x2=1.11 //y2=2.08
ends PM_DFFSNRNX1\%D

subckt PM_DFFSNRNX1\%noxref_13 ( 1 5 9 13 17 35 )
c46 ( 35 0 ) capacitor c=0.0731773f //x=0.455 //y=0.375
c47 ( 17 0 ) capacitor c=0.0259594f //x=2.445 //y=1.59
c48 ( 13 0 ) capacitor c=0.0156939f //x=2.445 //y=0.54
c49 ( 9 0 ) capacitor c=0.00678203f //x=1.56 //y=0.625
c50 ( 5 0 ) capacitor c=0.0236189f //x=1.475 //y=1.59
c51 ( 1 0 ) capacitor c=0.0109947f //x=0.59 //y=1.505
r52 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=1.59 //x2=1.56 //y2=1.63
r53 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=1.59 //x2=2.045 //y2=1.59
r54 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=1.59 //x2=2.53 //y2=1.59
r55 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=1.59 //x2=2.045 //y2=1.59
r56 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=0.54 //x2=1.56 //y2=0.5
r57 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=0.54 //x2=2.045 //y2=0.54
r58 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=0.54 //x2=2.53 //y2=0.54
r59 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=0.54 //x2=2.045 //y2=0.54
r60 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=1.63
r61 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=0.89
r62 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.5
r63 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.89
r64 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.675 //y=1.59 //x2=0.59 //y2=1.63
r65 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.675 //y=1.59 //x2=1.075 //y2=1.59
r66 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.475 //y=1.59 //x2=1.56 //y2=1.63
r67 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.475 //y=1.59 //x2=1.075 //y2=1.59
r68 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.59 //y=1.505 //x2=0.59 //y2=1.63
r69 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.59 //y=1.505 //x2=0.59 //y2=0.89
ends PM_DFFSNRNX1\%noxref_13

subckt PM_DFFSNRNX1\%noxref_14 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0432447f //x=2.965 //y=0.375
c54 ( 28 0 ) capacitor c=0.00466591f //x=1.86 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=3.1 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=4.07 //y=0.625
c57 ( 11 0 ) capacitor c=0.0152133f //x=3.985 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=3.1 //y=0.625
c59 ( 1 0 ) capacitor c=0.0255948f //x=3.015 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.185 //y=0.54 //x2=3.1 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.185 //y=0.54 //x2=3.585 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.985 //y=0.54 //x2=4.07 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.985 //y=0.54 //x2=3.585 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.135 //y=0.995 //x2=2.05 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=3.1 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=2.135 //y2=0.995
ends PM_DFFSNRNX1\%noxref_14

subckt PM_DFFSNRNX1\%noxref_15 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0686862f //x=5.265 //y=0.375
c53 ( 17 0 ) capacitor c=0.019765f //x=7.255 //y=1.59
c54 ( 13 0 ) capacitor c=0.0155888f //x=7.255 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=6.37 //y=0.625
c56 ( 5 0 ) capacitor c=0.0177541f //x=6.285 //y=1.59
c57 ( 1 0 ) capacitor c=0.00762097f //x=5.4 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.455 //y=1.59 //x2=6.37 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.455 //y=1.59 //x2=6.855 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.255 //y=1.59 //x2=7.34 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.255 //y=1.59 //x2=6.855 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.455 //y=0.54 //x2=6.37 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.455 //y=0.54 //x2=6.855 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.255 //y=0.54 //x2=7.34 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.255 //y=0.54 //x2=6.855 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=6.37 //y=1.505 //x2=6.37 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.37 //y=1.505 //x2=6.37 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.37 //y=0.625 //x2=6.37 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.37 //y=0.625 //x2=6.37 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.485 //y=1.59 //x2=5.4 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.485 //y=1.59 //x2=5.885 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.285 //y=1.59 //x2=6.37 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.285 //y=1.59 //x2=5.885 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=5.4 //y=1.505 //x2=5.4 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=5.4 //y=1.505 //x2=5.4 //y2=0.89
ends PM_DFFSNRNX1\%noxref_15

subckt PM_DFFSNRNX1\%noxref_16 ( 1 3 11 15 25 28 29 )
c54 ( 29 0 ) capacitor c=0.0422014f //x=7.775 //y=0.375
c55 ( 28 0 ) capacitor c=0.00461992f //x=6.67 //y=0.91
c56 ( 25 0 ) capacitor c=0.00156479f //x=7.91 //y=0.995
c57 ( 15 0 ) capacitor c=0.00737666f //x=8.88 //y=0.625
c58 ( 11 0 ) capacitor c=0.0147502f //x=8.795 //y=0.54
c59 ( 3 0 ) capacitor c=0.00718386f //x=7.91 //y=0.625
c60 ( 1 0 ) capacitor c=0.0234542f //x=7.825 //y=0.995
r61 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=8.88 //y=0.625 //x2=8.88 //y2=0.5
r62 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=8.88 //y=0.625 //x2=8.88 //y2=0.89
r63 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.995 //y=0.54 //x2=7.91 //y2=0.5
r64 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.995 //y=0.54 //x2=8.395 //y2=0.54
r65 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.795 //y=0.54 //x2=8.88 //y2=0.5
r66 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.795 //y=0.54 //x2=8.395 //y2=0.54
r67 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.91 //y=1.08 //x2=7.91 //y2=0.995
r68 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=7.91 //y=1.08 //x2=7.91 //y2=1.23
r69 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.91 //x2=7.91 //y2=0.995
r70 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.91 //x2=7.91 //y2=0.89
r71 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.625 //x2=7.91 //y2=0.5
r72 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.625 //x2=7.91 //y2=0.89
r73 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.945 //y=0.995 //x2=6.86 //y2=0.995
r74 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.825 //y=0.995 //x2=7.91 //y2=0.995
r75 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=7.825 //y=0.995 //x2=6.945 //y2=0.995
ends PM_DFFSNRNX1\%noxref_16

subckt PM_DFFSNRNX1\%noxref_17 ( 1 5 9 13 17 35 )
c54 ( 35 0 ) capacitor c=0.0686255f //x=10.075 //y=0.375
c55 ( 17 0 ) capacitor c=0.020294f //x=12.065 //y=1.59
c56 ( 13 0 ) capacitor c=0.0155578f //x=12.065 //y=0.54
c57 ( 9 0 ) capacitor c=0.00678203f //x=11.18 //y=0.625
c58 ( 5 0 ) capacitor c=0.0181206f //x=11.095 //y=1.59
c59 ( 1 0 ) capacitor c=0.00762097f //x=10.21 //y=1.505
r60 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.265 //y=1.59 //x2=11.18 //y2=1.63
r61 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.265 //y=1.59 //x2=11.665 //y2=1.59
r62 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.065 //y=1.59 //x2=12.15 //y2=1.59
r63 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.065 //y=1.59 //x2=11.665 //y2=1.59
r64 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.265 //y=0.54 //x2=11.18 //y2=0.5
r65 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.265 //y=0.54 //x2=11.665 //y2=0.54
r66 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.065 //y=0.54 //x2=12.15 //y2=0.54
r67 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.065 //y=0.54 //x2=11.665 //y2=0.54
r68 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=11.18 //y=1.505 //x2=11.18 //y2=1.63
r69 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=11.18 //y=1.505 //x2=11.18 //y2=0.89
r70 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=11.18 //y=0.625 //x2=11.18 //y2=0.5
r71 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=11.18 //y=0.625 //x2=11.18 //y2=0.89
r72 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.295 //y=1.59 //x2=10.21 //y2=1.63
r73 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.295 //y=1.59 //x2=10.695 //y2=1.59
r74 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.095 //y=1.59 //x2=11.18 //y2=1.63
r75 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.095 //y=1.59 //x2=10.695 //y2=1.59
r76 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=10.21 //y=1.505 //x2=10.21 //y2=1.63
r77 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=10.21 //y=1.505 //x2=10.21 //y2=0.89
ends PM_DFFSNRNX1\%noxref_17

subckt PM_DFFSNRNX1\%noxref_18 ( 1 3 11 15 25 28 29 )
c54 ( 29 0 ) capacitor c=0.0418028f //x=12.585 //y=0.375
c55 ( 28 0 ) capacitor c=0.00462171f //x=11.48 //y=0.91
c56 ( 25 0 ) capacitor c=0.00156479f //x=12.72 //y=0.995
c57 ( 15 0 ) capacitor c=0.00737666f //x=13.69 //y=0.625
c58 ( 11 0 ) capacitor c=0.0145763f //x=13.605 //y=0.54
c59 ( 3 0 ) capacitor c=0.00718386f //x=12.72 //y=0.625
c60 ( 1 0 ) capacitor c=0.0227139f //x=12.635 //y=0.995
r61 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=13.69 //y=0.625 //x2=13.69 //y2=0.5
r62 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=13.69 //y=0.625 //x2=13.69 //y2=0.89
r63 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.805 //y=0.54 //x2=12.72 //y2=0.5
r64 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.805 //y=0.54 //x2=13.205 //y2=0.54
r65 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.605 //y=0.54 //x2=13.69 //y2=0.5
r66 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.605 //y=0.54 //x2=13.205 //y2=0.54
r67 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=12.72 //y=1.08 //x2=12.72 //y2=0.995
r68 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=12.72 //y=1.08 //x2=12.72 //y2=1.23
r69 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.91 //x2=12.72 //y2=0.995
r70 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.91 //x2=12.72 //y2=0.89
r71 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.625 //x2=12.72 //y2=0.5
r72 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.625 //x2=12.72 //y2=0.89
r73 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.755 //y=0.995 //x2=11.67 //y2=0.995
r74 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=12.635 //y=0.995 //x2=12.72 //y2=0.995
r75 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=12.635 //y=0.995 //x2=11.755 //y2=0.995
ends PM_DFFSNRNX1\%noxref_18

subckt PM_DFFSNRNX1\%noxref_19 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0679963f //x=14.885 //y=0.375
c51 ( 17 0 ) capacitor c=0.018806f //x=16.875 //y=1.59
c52 ( 13 0 ) capacitor c=0.0155484f //x=16.875 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=15.99 //y=0.625
c54 ( 5 0 ) capacitor c=0.0170872f //x=15.905 //y=1.59
c55 ( 1 0 ) capacitor c=0.00729042f //x=15.02 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.075 //y=1.59 //x2=15.99 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.075 //y=1.59 //x2=16.475 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.875 //y=1.59 //x2=16.96 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.875 //y=1.59 //x2=16.475 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.075 //y=0.54 //x2=15.99 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.075 //y=0.54 //x2=16.475 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.875 //y=0.54 //x2=16.96 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.875 //y=0.54 //x2=16.475 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=15.99 //y=1.505 //x2=15.99 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=15.99 //y=1.505 //x2=15.99 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=15.99 //y=0.625 //x2=15.99 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=15.99 //y=0.625 //x2=15.99 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.105 //y=1.59 //x2=15.02 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.105 //y=1.59 //x2=15.505 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.905 //y=1.59 //x2=15.99 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.905 //y=1.59 //x2=15.505 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=15.02 //y=1.505 //x2=15.02 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=15.02 //y=1.505 //x2=15.02 //y2=0.89
ends PM_DFFSNRNX1\%noxref_19

subckt PM_DFFSNRNX1\%noxref_20 ( 1 3 11 15 25 28 29 )
c54 ( 29 0 ) capacitor c=0.0418028f //x=17.395 //y=0.375
c55 ( 28 0 ) capacitor c=0.00460056f //x=16.29 //y=0.91
c56 ( 25 0 ) capacitor c=0.00156479f //x=17.53 //y=0.995
c57 ( 15 0 ) capacitor c=0.00737666f //x=18.5 //y=0.625
c58 ( 11 0 ) capacitor c=0.0145763f //x=18.415 //y=0.54
c59 ( 3 0 ) capacitor c=0.00718386f //x=17.53 //y=0.625
c60 ( 1 0 ) capacitor c=0.022715f //x=17.445 //y=0.995
r61 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=18.5 //y=0.625 //x2=18.5 //y2=0.5
r62 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=18.5 //y=0.625 //x2=18.5 //y2=0.89
r63 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.615 //y=0.54 //x2=17.53 //y2=0.5
r64 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.615 //y=0.54 //x2=18.015 //y2=0.54
r65 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.415 //y=0.54 //x2=18.5 //y2=0.5
r66 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.415 //y=0.54 //x2=18.015 //y2=0.54
r67 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.53 //y=1.08 //x2=17.53 //y2=0.995
r68 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=17.53 //y=1.08 //x2=17.53 //y2=1.23
r69 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.91 //x2=17.53 //y2=0.995
r70 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.91 //x2=17.53 //y2=0.89
r71 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.625 //x2=17.53 //y2=0.5
r72 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.625 //x2=17.53 //y2=0.89
r73 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.565 //y=0.995 //x2=16.48 //y2=0.995
r74 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.445 //y=0.995 //x2=17.53 //y2=0.995
r75 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=17.445 //y=0.995 //x2=16.565 //y2=0.995
ends PM_DFFSNRNX1\%noxref_20

subckt PM_DFFSNRNX1\%noxref_21 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0679963f //x=19.695 //y=0.375
c51 ( 17 0 ) capacitor c=0.018806f //x=21.685 //y=1.59
c52 ( 13 0 ) capacitor c=0.0155484f //x=21.685 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=20.8 //y=0.625
c54 ( 5 0 ) capacitor c=0.0170872f //x=20.715 //y=1.59
c55 ( 1 0 ) capacitor c=0.00729042f //x=19.83 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.885 //y=1.59 //x2=20.8 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.885 //y=1.59 //x2=21.285 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.685 //y=1.59 //x2=21.77 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.685 //y=1.59 //x2=21.285 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.885 //y=0.54 //x2=20.8 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.885 //y=0.54 //x2=21.285 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.685 //y=0.54 //x2=21.77 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.685 //y=0.54 //x2=21.285 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=20.8 //y=1.505 //x2=20.8 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=20.8 //y=1.505 //x2=20.8 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=20.8 //y=0.625 //x2=20.8 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=20.8 //y=0.625 //x2=20.8 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.915 //y=1.59 //x2=19.83 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.915 //y=1.59 //x2=20.315 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.715 //y=1.59 //x2=20.8 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.715 //y=1.59 //x2=20.315 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=19.83 //y=1.505 //x2=19.83 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=19.83 //y=1.505 //x2=19.83 //y2=0.89
ends PM_DFFSNRNX1\%noxref_21

subckt PM_DFFSNRNX1\%noxref_22 ( 1 3 11 15 25 28 29 )
c54 ( 29 0 ) capacitor c=0.0418028f //x=22.205 //y=0.375
c55 ( 28 0 ) capacitor c=0.00460056f //x=21.1 //y=0.91
c56 ( 25 0 ) capacitor c=0.00156479f //x=22.34 //y=0.995
c57 ( 15 0 ) capacitor c=0.00737666f //x=23.31 //y=0.625
c58 ( 11 0 ) capacitor c=0.0145763f //x=23.225 //y=0.54
c59 ( 3 0 ) capacitor c=0.00718386f //x=22.34 //y=0.625
c60 ( 1 0 ) capacitor c=0.022715f //x=22.255 //y=0.995
r61 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=23.31 //y=0.625 //x2=23.31 //y2=0.5
r62 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=23.31 //y=0.625 //x2=23.31 //y2=0.89
r63 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=22.425 //y=0.54 //x2=22.34 //y2=0.5
r64 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.425 //y=0.54 //x2=22.825 //y2=0.54
r65 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.225 //y=0.54 //x2=23.31 //y2=0.5
r66 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.225 //y=0.54 //x2=22.825 //y2=0.54
r67 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.34 //y=1.08 //x2=22.34 //y2=0.995
r68 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=22.34 //y=1.08 //x2=22.34 //y2=1.23
r69 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.91 //x2=22.34 //y2=0.995
r70 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.91 //x2=22.34 //y2=0.89
r71 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.625 //x2=22.34 //y2=0.5
r72 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.625 //x2=22.34 //y2=0.89
r73 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.375 //y=0.995 //x2=21.29 //y2=0.995
r74 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.255 //y=0.995 //x2=22.34 //y2=0.995
r75 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=22.255 //y=0.995 //x2=21.375 //y2=0.995
ends PM_DFFSNRNX1\%noxref_22

subckt PM_DFFSNRNX1\%noxref_23 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0689605f //x=24.505 //y=0.375
c51 ( 17 0 ) capacitor c=0.0190974f //x=26.495 //y=1.59
c52 ( 13 0 ) capacitor c=0.0155819f //x=26.495 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=25.61 //y=0.625
c54 ( 5 0 ) capacitor c=0.0170872f //x=25.525 //y=1.59
c55 ( 1 0 ) capacitor c=0.00729042f //x=24.64 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.695 //y=1.59 //x2=25.61 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.695 //y=1.59 //x2=26.095 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.495 //y=1.59 //x2=26.58 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.495 //y=1.59 //x2=26.095 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.695 //y=0.54 //x2=25.61 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.695 //y=0.54 //x2=26.095 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.495 //y=0.54 //x2=26.58 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.495 //y=0.54 //x2=26.095 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=25.61 //y=1.505 //x2=25.61 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=25.61 //y=1.505 //x2=25.61 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=25.61 //y=0.625 //x2=25.61 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=25.61 //y=0.625 //x2=25.61 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=24.725 //y=1.59 //x2=24.64 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=24.725 //y=1.59 //x2=25.125 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.525 //y=1.59 //x2=25.61 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.525 //y=1.59 //x2=25.125 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=24.64 //y=1.505 //x2=24.64 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=24.64 //y=1.505 //x2=24.64 //y2=0.89
ends PM_DFFSNRNX1\%noxref_23

subckt PM_DFFSNRNX1\%noxref_24 ( 1 3 11 15 25 28 29 )
c50 ( 29 0 ) capacitor c=0.0428586f //x=27.015 //y=0.375
c51 ( 28 0 ) capacitor c=0.00460023f //x=25.91 //y=0.91
c52 ( 25 0 ) capacitor c=0.00156479f //x=27.15 //y=0.995
c53 ( 15 0 ) capacitor c=0.00737666f //x=28.12 //y=0.625
c54 ( 11 0 ) capacitor c=0.0148675f //x=28.035 //y=0.54
c55 ( 3 0 ) capacitor c=0.00718386f //x=27.15 //y=0.625
c56 ( 1 0 ) capacitor c=0.024626f //x=27.065 //y=0.995
r57 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=28.12 //y=0.625 //x2=28.12 //y2=0.5
r58 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=28.12 //y=0.625 //x2=28.12 //y2=0.89
r59 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=27.235 //y=0.54 //x2=27.15 //y2=0.5
r60 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=27.235 //y=0.54 //x2=27.635 //y2=0.54
r61 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=28.035 //y=0.54 //x2=28.12 //y2=0.5
r62 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=28.035 //y=0.54 //x2=27.635 //y2=0.54
r63 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.15 //y=1.08 //x2=27.15 //y2=0.995
r64 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=27.15 //y=1.08 //x2=27.15 //y2=1.23
r65 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.91 //x2=27.15 //y2=0.995
r66 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.91 //x2=27.15 //y2=0.89
r67 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.625 //x2=27.15 //y2=0.5
r68 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.625 //x2=27.15 //y2=0.89
r69 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.185 //y=0.995 //x2=26.1 //y2=0.995
r70 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.065 //y=0.995 //x2=27.15 //y2=0.995
r71 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=27.065 //y=0.995 //x2=26.185 //y2=0.995
ends PM_DFFSNRNX1\%noxref_24

