* SPICE3 file created from TIELO.ext - technology: sky130A

.subckt TIELO YN VPB VNB
M1000 a_121_383.t3 a_121_383.t2 VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VPB.t0 a_121_383.t0 a_121_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
R0 a_121_383.n0 a_121_383.t0 512.525
R1 a_121_383.n0 a_121_383.t2 371.139
R2 a_121_383.n1 a_121_383.t4 312.699
R3 a_121_383.n2 a_121_383.n1 75.63
R4 a_121_383.n1 a_121_383.n0 58.377
R5 a_121_383.n2 a_121_383.t1 14.282
R6 a_121_383.t3 a_121_383.n2 14.282
R7 VPB VPB.n62 126.832
R8 VPB.n52 VPB.n51 76
R9 VPB.n44 VPB.n15 76
R10 VPB.n55 VPB.n54 76
R11 VPB.n42 VPB.n41 66.753
R12 VPB.n46 VPB.n45 66.753
R13 VPB.n14 VPB.t1 55.106
R14 VPB.n40 VPB.t0 55.106
R15 VPB.n59 VPB.n55 20.452
R16 VPB.n39 VPB.n36 20.452
R17 VPB.n39 VPB.n38 13.653
R18 VPB.n38 VPB.n37 13.653
R19 VPB.n44 VPB.n43 13.653
R20 VPB.n43 VPB.n42 13.653
R21 VPB.n51 VPB.n50 13.653
R22 VPB.n50 VPB.n49 13.653
R23 VPB.n48 VPB.n47 13.653
R24 VPB.n47 VPB.n46 13.653
R25 VPB.n55 VPB.n0 13.653
R26 VPB VPB.n0 13.653
R27 VPB.n59 VPB.n58 13.276
R28 VPB.n58 VPB.n56 13.276
R29 VPB.n51 VPB.n44 13.276
R30 VPB.n51 VPB.n48 13.276
R31 VPB.n36 VPB.n18 13.276
R32 VPB.n18 VPB.n16 13.276
R33 VPB.n23 VPB.n21 12.796
R34 VPB.n23 VPB.n22 12.564
R35 VPB.n31 VPB.n30 12.198
R36 VPB.n27 VPB.n26 12.198
R37 VPB.n31 VPB.n28 12.198
R38 VPB.n40 VPB.n39 10.764
R39 VPB.n55 VPB.n14 10.764
R40 VPB.n36 VPB.n35 7.5
R41 VPB.n21 VPB.n20 7.5
R42 VPB.n26 VPB.n25 7.5
R43 VPB.n30 VPB.n29 7.5
R44 VPB.n18 VPB.n17 7.5
R45 VPB.n33 VPB.n19 7.5
R46 VPB.n58 VPB.n57 7.5
R47 VPB.n12 VPB.n11 7.5
R48 VPB.n6 VPB.n5 7.5
R49 VPB.n8 VPB.n7 7.5
R50 VPB.n2 VPB.n1 7.5
R51 VPB.n60 VPB.n59 7.5
R52 VPB.n13 VPB.n10 6.729
R53 VPB.n9 VPB.n6 6.729
R54 VPB.n4 VPB.n2 6.729
R55 VPB.n4 VPB.n3 6.728
R56 VPB.n9 VPB.n8 6.728
R57 VPB.n13 VPB.n12 6.728
R58 VPB.n61 VPB.n60 6.728
R59 VPB.n35 VPB.n34 6.398
R60 VPB.n44 VPB.n40 2.511
R61 VPB.n48 VPB.n14 2.511
R62 VPB.n33 VPB.n24 1.402
R63 VPB.n33 VPB.n27 1.402
R64 VPB.n33 VPB.n31 1.402
R65 VPB.n33 VPB.n32 1.402
R66 VPB.n34 VPB.n33 0.735
R67 VPB.n33 VPB.n23 0.735
R68 VPB.n62 VPB.n13 0.387
R69 VPB.n62 VPB.n9 0.387
R70 VPB.n62 VPB.n4 0.387
R71 VPB.n62 VPB.n61 0.387
R72 VPB.n54 VPB 0.198
R73 VPB.n52 VPB.n15 0.136
R74 VPB.n53 VPB.n52 0.136
R75 VPB.n54 VPB.n53 0.136
R76 VNB VNB.n58 1525
R77 VNB.n58 VNB 1525
R78 VNB.n33 VNB.n6 76
R79 VNB.n38 VNB.n37 76
R80 VNB.n56 VNB.n40 76
R81 VNB.n3 VNB.t0 39.412
R82 VNB.n13 VNB.n12 35.01
R83 VNB.n30 VNB.n28 20.452
R84 VNB.n56 VNB.n55 20.452
R85 VNB.n37 VNB.n9 19.735
R86 VNB.n31 VNB.n13 19.735
R87 VNB.n5 VNB.n4 19.735
R88 VNB.n13 VNB.n11 19.017
R89 VNB.n17 VNB.n14 18.356
R90 VNB.n44 VNB.n41 18.356
R91 VNB.n3 VNB.n2 17.185
R92 VNB.n20 VNB.n17 13.919
R93 VNB.n47 VNB.n44 13.919
R94 VNB.n36 VNB.n35 13.653
R95 VNB.n37 VNB.n34 13.653
R96 VNB.n33 VNB.n32 13.653
R97 VNB.n30 VNB.n29 13.653
R98 VNB.n57 VNB.n56 13.653
R99 VNB.n58 VNB.n57 13.653
R100 VNB.n23 VNB.n20 13.276
R101 VNB.n26 VNB.n23 13.276
R102 VNB.n28 VNB.n26 13.276
R103 VNB.n50 VNB.n47 13.276
R104 VNB.n53 VNB.n50 13.276
R105 VNB.n55 VNB.n53 13.276
R106 VNB.n37 VNB.n33 13.276
R107 VNB.n37 VNB.n36 13.276
R108 VNB.n56 VNB.n5 9.329
R109 VNB.n31 VNB.n30 8.97
R110 VNB.n11 VNB.n10 7.5
R111 VNB.n9 VNB.n8 7.5
R112 VNB.n28 VNB.n27 7.5
R113 VNB.n16 VNB.n15 7.5
R114 VNB.n20 VNB.n19 7.5
R115 VNB.n19 VNB.n18 7.5
R116 VNB.n23 VNB.n22 7.5
R117 VNB.n22 VNB.n21 7.5
R118 VNB.n26 VNB.n25 7.5
R119 VNB.n43 VNB.n42 7.5
R120 VNB.n55 VNB.n54 7.5
R121 VNB.n53 VNB.n52 7.5
R122 VNB.n50 VNB.n49 7.5
R123 VNB.n49 VNB.n48 7.5
R124 VNB.n47 VNB.n46 7.5
R125 VNB.n46 VNB.n45 7.5
R126 VNB.n17 VNB.n16 6.627
R127 VNB.n44 VNB.n43 6.627
R128 VNB.n4 VNB.n3 6.139
R129 VNB.n1 VNB.n0 4.551
R130 VNB.n33 VNB.n31 4.305
R131 VNB.n36 VNB.n5 3.947
R132 VNB.t0 VNB.n1 2.238
R133 VNB.n8 VNB.n7 1.935
R134 VNB.n25 VNB.n24 0.454
R135 VNB.n52 VNB.n51 0.454
R136 VNB.n40 VNB 0.198
R137 VNB.n38 VNB.n6 0.136
R138 VNB.n39 VNB.n38 0.136
R139 VNB.n40 VNB.n39 0.136
R140 a_185_181.n1 a_185_181.n0 27.232
C0 VPB VNB 2.90fF
C1 a_185_181.n0 VNB 0.37fF
C2 a_185_181.n1 VNB 0.39fF
C3 VPB.n0 VNB 0.03fF
C4 VPB.n1 VNB 0.03fF
C5 VPB.n2 VNB 0.02fF
C6 VPB.n3 VNB 0.09fF
C7 VPB.n5 VNB 0.02fF
C8 VPB.n6 VNB 0.02fF
C9 VPB.n7 VNB 0.02fF
C10 VPB.n8 VNB 0.02fF
C11 VPB.n10 VNB 0.02fF
C12 VPB.n11 VNB 0.02fF
C13 VPB.n12 VNB 0.02fF
C14 VPB.n14 VNB 0.05fF
C15 VPB.n15 VNB 0.06fF
C16 VPB.n16 VNB 0.02fF
C17 VPB.n17 VNB 0.02fF
C18 VPB.n18 VNB 0.02fF
C19 VPB.n19 VNB 0.09fF
C20 VPB.n20 VNB 0.02fF
C21 VPB.n21 VNB 0.02fF
C22 VPB.n22 VNB 0.04fF
C23 VPB.n23 VNB 0.01fF
C24 VPB.n25 VNB 0.02fF
C25 VPB.n26 VNB 0.02fF
C26 VPB.n28 VNB 0.02fF
C27 VPB.n29 VNB 0.02fF
C28 VPB.n30 VNB 0.02fF
C29 VPB.n33 VNB 0.39fF
C30 VPB.n35 VNB 0.03fF
C31 VPB.n36 VNB 0.03fF
C32 VPB.n37 VNB 0.23fF
C33 VPB.n38 VNB 0.03fF
C34 VPB.n39 VNB 0.03fF
C35 VPB.n40 VNB 0.05fF
C36 VPB.n41 VNB 0.12fF
C37 VPB.n42 VNB 0.16fF
C38 VPB.n43 VNB 0.02fF
C39 VPB.n44 VNB 0.01fF
C40 VPB.n45 VNB 0.12fF
C41 VPB.n46 VNB 0.16fF
C42 VPB.n47 VNB 0.02fF
C43 VPB.n48 VNB 0.01fF
C44 VPB.n49 VNB 0.14fF
C45 VPB.n50 VNB 0.02fF
C46 VPB.n51 VNB 0.02fF
C47 VPB.n52 VNB 0.02fF
C48 VPB.n53 VNB 0.02fF
C49 VPB.n54 VNB 0.03fF
C50 VPB.n55 VNB 0.03fF
C51 VPB.n56 VNB 0.02fF
C52 VPB.n57 VNB 0.02fF
C53 VPB.n58 VNB 0.02fF
C54 VPB.n59 VNB 0.03fF
C55 VPB.n60 VNB 0.03fF
C56 VPB.n62 VNB 0.36fF
C57 a_121_383.t4 VNB 0.40fF
C58 a_121_383.n0 VNB 0.15fF
C59 a_121_383.n1 VNB 0.33fF
C60 a_121_383.n2 VNB 0.40fF
.ends
