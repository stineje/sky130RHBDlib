// File: dffsnrnx1_pcell.spi.pex
// Created: Tue Oct 15 15:56:04 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_DFFSNRNX1_PCELL\%noxref_1 ( 49 53 56 61 71 79 89 97 107 115 125 133 \
 143 158 162 164 166 168 170 172 173 174 175 176 177 )
c312 ( 177 0 ) capacitor c=0.0226424f //x=24.935 //y=0.875
c313 ( 176 0 ) capacitor c=0.0225954f //x=20.125 //y=0.875
c314 ( 175 0 ) capacitor c=0.0225954f //x=15.315 //y=0.875
c315 ( 174 0 ) capacitor c=0.0225954f //x=10.505 //y=0.875
c316 ( 173 0 ) capacitor c=0.0225954f //x=5.695 //y=0.875
c317 ( 172 0 ) capacitor c=0.0226959f //x=0.885 //y=0.875
c318 ( 171 0 ) capacitor c=0.00440144f //x=25.125 //y=0
c319 ( 170 0 ) capacitor c=0.108076f //x=24.05 //y=0
c320 ( 169 0 ) capacitor c=0.00440144f //x=20.315 //y=0
c321 ( 168 0 ) capacitor c=0.106903f //x=19.24 //y=0
c322 ( 167 0 ) capacitor c=0.00440144f //x=15.505 //y=0
c323 ( 166 0 ) capacitor c=0.107052f //x=14.43 //y=0
c324 ( 165 0 ) capacitor c=0.00440144f //x=10.695 //y=0
c325 ( 164 0 ) capacitor c=0.107294f //x=9.62 //y=0
c326 ( 163 0 ) capacitor c=0.00440144f //x=5.885 //y=0
c327 ( 162 0 ) capacitor c=0.10703f //x=4.81 //y=0
c328 ( 161 0 ) capacitor c=0.00440144f //x=1.075 //y=0
c329 ( 158 0 ) capacitor c=0.322126f //x=28.12 //y=0
c330 ( 143 0 ) capacitor c=0.0339617f //x=25.04 //y=0
c331 ( 133 0 ) capacitor c=0.133607f //x=23.88 //y=0
c332 ( 125 0 ) capacitor c=0.0339325f //x=20.23 //y=0
c333 ( 115 0 ) capacitor c=0.133561f //x=19.07 //y=0
c334 ( 107 0 ) capacitor c=0.0339325f //x=15.42 //y=0
c335 ( 97 0 ) capacitor c=0.133362f //x=14.26 //y=0
c336 ( 89 0 ) capacitor c=0.0339325f //x=10.61 //y=0
c337 ( 79 0 ) capacitor c=0.133362f //x=9.45 //y=0
c338 ( 71 0 ) capacitor c=0.0339325f //x=5.8 //y=0
c339 ( 61 0 ) capacitor c=0.133402f //x=4.64 //y=0
c340 ( 56 0 ) capacitor c=0.178058f //x=0.74 //y=0
c341 ( 53 0 ) capacitor c=0.0367385f //x=0.99 //y=0
c342 ( 49 0 ) capacitor c=0.892258f //x=28.12 //y=0
r343 (  156 158 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=27.01 //y=0 //x2=28.12 //y2=0
r344 (  154 156 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=25.9 //y=0 //x2=27.01 //y2=0
r345 (  152 171 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.21 //y=0 //x2=25.125 //y2=0
r346 (  152 154 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=25.21 //y=0 //x2=25.9 //y2=0
r347 (  147 171 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.125 //y=0.17 //x2=25.125 //y2=0
r348 (  147 177 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=25.125 //y=0.17 //x2=25.125 //y2=0.965
r349 (  144 170 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.22 //y=0 //x2=24.05 //y2=0
r350 (  144 146 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.22 //y=0 //x2=24.79 //y2=0
r351 (  143 171 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.04 //y=0 //x2=25.125 //y2=0
r352 (  143 146 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=25.04 //y=0 //x2=24.79 //y2=0
r353 (  138 140 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=22.2 //y=0 //x2=23.31 //y2=0
r354 (  136 138 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=21.09 //y=0 //x2=22.2 //y2=0
r355 (  134 169 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.4 //y=0 //x2=20.315 //y2=0
r356 (  134 136 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=20.4 //y=0 //x2=21.09 //y2=0
r357 (  133 170 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.88 //y=0 //x2=24.05 //y2=0
r358 (  133 140 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=23.88 //y=0 //x2=23.31 //y2=0
r359 (  129 169 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.315 //y=0.17 //x2=20.315 //y2=0
r360 (  129 176 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=20.315 //y=0.17 //x2=20.315 //y2=0.965
r361 (  126 168 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.41 //y=0 //x2=19.24 //y2=0
r362 (  126 128 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.41 //y=0 //x2=19.98 //y2=0
r363 (  125 169 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.23 //y=0 //x2=20.315 //y2=0
r364 (  125 128 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=20.23 //y=0 //x2=19.98 //y2=0
r365 (  120 122 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=17.39 //y=0 //x2=18.5 //y2=0
r366 (  118 120 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=16.28 //y=0 //x2=17.39 //y2=0
r367 (  116 167 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.59 //y=0 //x2=15.505 //y2=0
r368 (  116 118 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=15.59 //y=0 //x2=16.28 //y2=0
r369 (  115 168 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.07 //y=0 //x2=19.24 //y2=0
r370 (  115 122 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.07 //y=0 //x2=18.5 //y2=0
r371 (  111 167 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.505 //y=0.17 //x2=15.505 //y2=0
r372 (  111 175 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=15.505 //y=0.17 //x2=15.505 //y2=0.965
r373 (  108 166 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.6 //y=0 //x2=14.43 //y2=0
r374 (  108 110 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.6 //y=0 //x2=15.17 //y2=0
r375 (  107 167 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.42 //y=0 //x2=15.505 //y2=0
r376 (  107 110 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=15.42 //y=0 //x2=15.17 //y2=0
r377 (  102 104 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=12.58 //y=0 //x2=13.69 //y2=0
r378 (  100 102 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=11.47 //y=0 //x2=12.58 //y2=0
r379 (  98 165 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.78 //y=0 //x2=10.695 //y2=0
r380 (  98 100 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=10.78 //y=0 //x2=11.47 //y2=0
r381 (  97 166 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.26 //y=0 //x2=14.43 //y2=0
r382 (  97 104 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.26 //y=0 //x2=13.69 //y2=0
r383 (  93 165 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.695 //y=0.17 //x2=10.695 //y2=0
r384 (  93 174 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=10.695 //y=0.17 //x2=10.695 //y2=0.965
r385 (  90 164 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.79 //y=0 //x2=9.62 //y2=0
r386 (  90 92 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.79 //y=0 //x2=10.36 //y2=0
r387 (  89 165 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.61 //y=0 //x2=10.695 //y2=0
r388 (  89 92 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=10.61 //y=0 //x2=10.36 //y2=0
r389 (  84 86 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=7.77 //y=0 //x2=8.88 //y2=0
r390 (  82 84 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r391 (  80 163 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.97 //y=0 //x2=5.885 //y2=0
r392 (  80 82 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=5.97 //y=0 //x2=6.66 //y2=0
r393 (  79 164 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.45 //y=0 //x2=9.62 //y2=0
r394 (  79 86 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.45 //y=0 //x2=8.88 //y2=0
r395 (  75 163 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.885 //y=0.17 //x2=5.885 //y2=0
r396 (  75 173 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=5.885 //y=0.17 //x2=5.885 //y2=0.965
r397 (  72 162 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=4.81 //y2=0
r398 (  72 74 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=5.55 //y2=0
r399 (  71 163 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.8 //y=0 //x2=5.885 //y2=0
r400 (  71 74 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=5.8 //y=0 //x2=5.55 //y2=0
r401 (  66 68 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=0 //x2=4.07 //y2=0
r402 (  64 66 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r403 (  62 161 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.075 //y2=0
r404 (  62 64 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.85 //y2=0
r405 (  61 162 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.81 //y2=0
r406 (  61 68 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.07 //y2=0
r407 (  57 161 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0
r408 (  57 172 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0.965
r409 (  53 161 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=1.075 //y2=0
r410 (  53 56 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=0.74 //y2=0
r411 (  49 158 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.12 //y=0 //x2=28.12 //y2=0
r412 (  47 156 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.01 //y=0 //x2=27.01 //y2=0
r413 (  47 49 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=27.01 //y=0 //x2=28.12 //y2=0
r414 (  45 154 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.9 //y=0 //x2=25.9 //y2=0
r415 (  45 47 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=25.9 //y=0 //x2=27.01 //y2=0
r416 (  43 146 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=0 //x2=24.79 //y2=0
r417 (  43 45 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=0 //x2=25.9 //y2=0
r418 (  41 140 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.31 //y=0 //x2=23.31 //y2=0
r419 (  41 43 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=23.31 //y=0 //x2=24.79 //y2=0
r420 (  39 138 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.2 //y=0 //x2=22.2 //y2=0
r421 (  39 41 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.2 //y=0 //x2=23.31 //y2=0
r422 (  37 136 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=0 //x2=21.09 //y2=0
r423 (  37 39 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=0 //x2=22.2 //y2=0
r424 (  35 128 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=0 //x2=19.98 //y2=0
r425 (  35 37 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=0 //x2=21.09 //y2=0
r426 (  33 122 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=0 //x2=18.5 //y2=0
r427 (  33 35 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=0 //x2=19.98 //y2=0
r428 (  31 120 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=0 //x2=17.39 //y2=0
r429 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=0 //x2=18.5 //y2=0
r430 (  29 118 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=0 //x2=16.28 //y2=0
r431 (  29 31 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=0 //x2=17.39 //y2=0
r432 (  27 110 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=0 //x2=15.17 //y2=0
r433 (  27 29 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=0 //x2=16.28 //y2=0
r434 (  25 104 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=0 //x2=13.69 //y2=0
r435 (  25 27 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=13.69 //y=0 //x2=15.17 //y2=0
r436 (  23 102 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=0 //x2=12.58 //y2=0
r437 (  23 25 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=0 //x2=13.69 //y2=0
r438 (  21 100 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=0 //x2=11.47 //y2=0
r439 (  21 23 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=0 //x2=12.58 //y2=0
r440 (  19 92 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r441 (  19 21 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=0 //x2=11.47 //y2=0
r442 (  17 86 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.88 //y=0 //x2=8.88 //y2=0
r443 (  17 19 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.88 //y=0 //x2=10.36 //y2=0
r444 (  15 84 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r445 (  15 17 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=8.88 //y2=0
r446 (  13 82 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r447 (  13 15 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r448 (  11 74 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r449 (  11 13 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r450 (  9 68 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r451 (  9 11 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=0 //x2=5.55 //y2=0
r452 (  7 66 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r453 (  7 9 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.07 //y2=0
r454 (  5 64 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r455 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r456 (  2 56 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r457 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
ends PM_DFFSNRNX1_PCELL\%noxref_1

subckt PM_DFFSNRNX1_PCELL\%noxref_2 ( 49 56 63 73 81 91 107 117 125 135 141 \
 151 161 169 179 185 195 205 213 223 239 249 257 267 283 293 301 314 321 326 \
 331 336 341 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 \
 362 363 364 365 366 367 368 369 )
c331 ( 369 0 ) capacitor c=0.0455453f //x=27.635 //y=5.02
c332 ( 368 0 ) capacitor c=0.0243052f //x=26.755 //y=5.02
c333 ( 367 0 ) capacitor c=0.0243052f //x=25.875 //y=5.02
c334 ( 366 0 ) capacitor c=0.0532177f //x=25.005 //y=5.02
c335 ( 365 0 ) capacitor c=0.0453711f //x=22.825 //y=5.02
c336 ( 364 0 ) capacitor c=0.0243052f //x=21.945 //y=5.02
c337 ( 363 0 ) capacitor c=0.0243052f //x=21.065 //y=5.02
c338 ( 362 0 ) capacitor c=0.0532177f //x=20.195 //y=5.02
c339 ( 361 0 ) capacitor c=0.0453711f //x=18.015 //y=5.02
c340 ( 360 0 ) capacitor c=0.0243052f //x=17.135 //y=5.02
c341 ( 359 0 ) capacitor c=0.024152f //x=16.255 //y=5.02
c342 ( 358 0 ) capacitor c=0.053132f //x=15.385 //y=5.02
c343 ( 357 0 ) capacitor c=0.0452179f //x=13.205 //y=5.02
c344 ( 356 0 ) capacitor c=0.024152f //x=12.325 //y=5.02
c345 ( 355 0 ) capacitor c=0.024152f //x=11.445 //y=5.02
c346 ( 354 0 ) capacitor c=0.053132f //x=10.575 //y=5.02
c347 ( 353 0 ) capacitor c=0.0452179f //x=8.395 //y=5.02
c348 ( 352 0 ) capacitor c=0.024152f //x=7.515 //y=5.02
c349 ( 351 0 ) capacitor c=0.0243529f //x=6.635 //y=5.02
c350 ( 350 0 ) capacitor c=0.0532483f //x=5.765 //y=5.02
c351 ( 349 0 ) capacitor c=0.0454188f //x=3.585 //y=5.02
c352 ( 348 0 ) capacitor c=0.0244314f //x=2.705 //y=5.02
c353 ( 347 0 ) capacitor c=0.0244794f //x=1.825 //y=5.02
c354 ( 346 0 ) capacitor c=0.0533644f //x=0.955 //y=5.02
c355 ( 345 0 ) capacitor c=0.00591168f //x=27.78 //y=7.4
c356 ( 344 0 ) capacitor c=0.00591168f //x=26.9 //y=7.4
c357 ( 343 0 ) capacitor c=0.00591168f //x=26.02 //y=7.4
c358 ( 342 0 ) capacitor c=0.00591168f //x=25.14 //y=7.4
c359 ( 341 0 ) capacitor c=0.159571f //x=24.05 //y=7.4
c360 ( 340 0 ) capacitor c=0.00591168f //x=22.97 //y=7.4
c361 ( 339 0 ) capacitor c=0.00591168f //x=22.09 //y=7.4
c362 ( 338 0 ) capacitor c=0.00591168f //x=21.21 //y=7.4
c363 ( 337 0 ) capacitor c=0.00591168f //x=20.33 //y=7.4
c364 ( 336 0 ) capacitor c=0.15939f //x=19.24 //y=7.4
c365 ( 335 0 ) capacitor c=0.00591168f //x=18.16 //y=7.4
c366 ( 334 0 ) capacitor c=0.00591168f //x=17.28 //y=7.4
c367 ( 333 0 ) capacitor c=0.00591168f //x=16.4 //y=7.4
c368 ( 332 0 ) capacitor c=0.00591168f //x=15.52 //y=7.4
c369 ( 331 0 ) capacitor c=0.159721f //x=14.43 //y=7.4
c370 ( 330 0 ) capacitor c=0.00591168f //x=13.35 //y=7.4
c371 ( 329 0 ) capacitor c=0.00591168f //x=12.47 //y=7.4
c372 ( 328 0 ) capacitor c=0.00591168f //x=11.59 //y=7.4
c373 ( 327 0 ) capacitor c=0.00591168f //x=10.71 //y=7.4
c374 ( 326 0 ) capacitor c=0.159745f //x=9.62 //y=7.4
c375 ( 325 0 ) capacitor c=0.00591168f //x=8.54 //y=7.4
c376 ( 324 0 ) capacitor c=0.00591168f //x=7.66 //y=7.4
c377 ( 323 0 ) capacitor c=0.00591168f //x=6.78 //y=7.4
c378 ( 322 0 ) capacitor c=0.00591168f //x=5.9 //y=7.4
c379 ( 321 0 ) capacitor c=0.159817f //x=4.81 //y=7.4
c380 ( 320 0 ) capacitor c=0.00591168f //x=3.73 //y=7.4
c381 ( 319 0 ) capacitor c=0.00591168f //x=2.85 //y=7.4
c382 ( 318 0 ) capacitor c=0.00591168f //x=1.97 //y=7.4
c383 ( 317 0 ) capacitor c=0.00591168f //x=1.09 //y=7.4
c384 ( 314 0 ) capacitor c=0.272255f //x=28.12 //y=7.4
c385 ( 301 0 ) capacitor c=0.028513f //x=27.695 //y=7.4
c386 ( 293 0 ) capacitor c=0.0287069f //x=26.815 //y=7.4
c387 ( 283 0 ) capacitor c=0.0292055f //x=25.935 //y=7.4
c388 ( 273 0 ) capacitor c=0.0452081f //x=25.055 //y=7.4
c389 ( 267 0 ) capacitor c=0.0418861f //x=23.88 //y=7.4
c390 ( 257 0 ) capacitor c=0.028513f //x=22.885 //y=7.4
c391 ( 249 0 ) capacitor c=0.0287069f //x=22.005 //y=7.4
c392 ( 239 0 ) capacitor c=0.0292055f //x=21.125 //y=7.4
c393 ( 229 0 ) capacitor c=0.0452081f //x=20.245 //y=7.4
c394 ( 223 0 ) capacitor c=0.0418861f //x=19.07 //y=7.4
c395 ( 213 0 ) capacitor c=0.028513f //x=18.075 //y=7.4
c396 ( 205 0 ) capacitor c=0.0288775f //x=17.195 //y=7.4
c397 ( 195 0 ) capacitor c=0.0284966f //x=16.315 //y=7.4
c398 ( 185 0 ) capacitor c=0.0383672f //x=15.435 //y=7.4
c399 ( 179 0 ) capacitor c=0.0394667f //x=14.26 //y=7.4
c400 ( 169 0 ) capacitor c=0.0288488f //x=13.265 //y=7.4
c401 ( 161 0 ) capacitor c=0.0287514f //x=12.385 //y=7.4
c402 ( 151 0 ) capacitor c=0.0284966f //x=11.505 //y=7.4
c403 ( 141 0 ) capacitor c=0.0383672f //x=10.625 //y=7.4
c404 ( 135 0 ) capacitor c=0.0394667f //x=9.45 //y=7.4
c405 ( 125 0 ) capacitor c=0.0288488f //x=8.455 //y=7.4
c406 ( 117 0 ) capacitor c=0.0287505f //x=7.575 //y=7.4
c407 ( 107 0 ) capacitor c=0.0292055f //x=6.695 //y=7.4
c408 ( 97 0 ) capacitor c=0.0452081f //x=5.815 //y=7.4
c409 ( 91 0 ) capacitor c=0.0418861f //x=4.64 //y=7.4
c410 ( 81 0 ) capacitor c=0.028513f //x=3.645 //y=7.4
c411 ( 73 0 ) capacitor c=0.0287069f //x=2.765 //y=7.4
c412 ( 63 0 ) capacitor c=0.0292055f //x=1.885 //y=7.4
c413 ( 56 0 ) capacitor c=0.235022f //x=0.74 //y=7.4
c414 ( 53 0 ) capacitor c=0.0452081f //x=1.005 //y=7.4
c415 ( 49 0 ) capacitor c=1.0243f //x=28.12 //y=7.4
r416 (  312 345 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.865 //y=7.4 //x2=27.78 //y2=7.4
r417 (  312 314 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=27.865 //y=7.4 //x2=28.12 //y2=7.4
r418 (  305 345 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.78 //y=7.23 //x2=27.78 //y2=7.4
r419 (  305 369 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=27.78 //y=7.23 //x2=27.78 //y2=6.745
r420 (  302 344 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.985 //y=7.4 //x2=26.9 //y2=7.4
r421 (  302 304 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=26.985 //y=7.4 //x2=27.01 //y2=7.4
r422 (  301 345 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.695 //y=7.4 //x2=27.78 //y2=7.4
r423 (  301 304 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=27.695 //y=7.4 //x2=27.01 //y2=7.4
r424 (  295 344 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.9 //y=7.23 //x2=26.9 //y2=7.4
r425 (  295 368 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.9 //y=7.23 //x2=26.9 //y2=6.745
r426 (  294 343 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.105 //y=7.4 //x2=26.02 //y2=7.4
r427 (  293 344 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.815 //y=7.4 //x2=26.9 //y2=7.4
r428 (  293 294 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=26.815 //y=7.4 //x2=26.105 //y2=7.4
r429 (  287 343 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.02 //y=7.23 //x2=26.02 //y2=7.4
r430 (  287 367 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.02 //y=7.23 //x2=26.02 //y2=6.745
r431 (  284 342 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.225 //y=7.4 //x2=25.14 //y2=7.4
r432 (  284 286 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=25.225 //y=7.4 //x2=25.9 //y2=7.4
r433 (  283 343 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.935 //y=7.4 //x2=26.02 //y2=7.4
r434 (  283 286 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=25.935 //y=7.4 //x2=25.9 //y2=7.4
r435 (  277 342 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.14 //y=7.23 //x2=25.14 //y2=7.4
r436 (  277 366 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=25.14 //y=7.23 //x2=25.14 //y2=6.405
r437 (  274 341 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.22 //y=7.4 //x2=24.05 //y2=7.4
r438 (  274 276 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.22 //y=7.4 //x2=24.79 //y2=7.4
r439 (  273 342 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.055 //y=7.4 //x2=25.14 //y2=7.4
r440 (  273 276 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=25.055 //y=7.4 //x2=24.79 //y2=7.4
r441 (  268 340 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.055 //y=7.4 //x2=22.97 //y2=7.4
r442 (  268 270 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=23.055 //y=7.4 //x2=23.31 //y2=7.4
r443 (  267 341 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.88 //y=7.4 //x2=24.05 //y2=7.4
r444 (  267 270 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=23.88 //y=7.4 //x2=23.31 //y2=7.4
r445 (  261 340 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.97 //y=7.23 //x2=22.97 //y2=7.4
r446 (  261 365 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.97 //y=7.23 //x2=22.97 //y2=6.745
r447 (  258 339 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.175 //y=7.4 //x2=22.09 //y2=7.4
r448 (  258 260 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=22.175 //y=7.4 //x2=22.2 //y2=7.4
r449 (  257 340 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.885 //y=7.4 //x2=22.97 //y2=7.4
r450 (  257 260 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=22.885 //y=7.4 //x2=22.2 //y2=7.4
r451 (  251 339 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.09 //y=7.23 //x2=22.09 //y2=7.4
r452 (  251 364 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.09 //y=7.23 //x2=22.09 //y2=6.745
r453 (  250 338 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.295 //y=7.4 //x2=21.21 //y2=7.4
r454 (  249 339 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.005 //y=7.4 //x2=22.09 //y2=7.4
r455 (  249 250 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.005 //y=7.4 //x2=21.295 //y2=7.4
r456 (  243 338 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.21 //y=7.23 //x2=21.21 //y2=7.4
r457 (  243 363 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.21 //y=7.23 //x2=21.21 //y2=6.745
r458 (  240 337 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.415 //y=7.4 //x2=20.33 //y2=7.4
r459 (  240 242 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=20.415 //y=7.4 //x2=21.09 //y2=7.4
r460 (  239 338 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.125 //y=7.4 //x2=21.21 //y2=7.4
r461 (  239 242 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=21.125 //y=7.4 //x2=21.09 //y2=7.4
r462 (  233 337 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.33 //y=7.23 //x2=20.33 //y2=7.4
r463 (  233 362 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=20.33 //y=7.23 //x2=20.33 //y2=6.405
r464 (  230 336 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.41 //y=7.4 //x2=19.24 //y2=7.4
r465 (  230 232 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.41 //y=7.4 //x2=19.98 //y2=7.4
r466 (  229 337 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.245 //y=7.4 //x2=20.33 //y2=7.4
r467 (  229 232 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=20.245 //y=7.4 //x2=19.98 //y2=7.4
r468 (  224 335 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.245 //y=7.4 //x2=18.16 //y2=7.4
r469 (  224 226 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=18.245 //y=7.4 //x2=18.5 //y2=7.4
r470 (  223 336 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.07 //y=7.4 //x2=19.24 //y2=7.4
r471 (  223 226 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.07 //y=7.4 //x2=18.5 //y2=7.4
r472 (  217 335 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.16 //y=7.23 //x2=18.16 //y2=7.4
r473 (  217 361 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=18.16 //y=7.23 //x2=18.16 //y2=6.745
r474 (  214 334 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.365 //y=7.4 //x2=17.28 //y2=7.4
r475 (  214 216 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=17.365 //y=7.4 //x2=17.39 //y2=7.4
r476 (  213 335 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.075 //y=7.4 //x2=18.16 //y2=7.4
r477 (  213 216 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=18.075 //y=7.4 //x2=17.39 //y2=7.4
r478 (  207 334 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.28 //y=7.23 //x2=17.28 //y2=7.4
r479 (  207 360 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.28 //y=7.23 //x2=17.28 //y2=6.745
r480 (  206 333 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.485 //y=7.4 //x2=16.4 //y2=7.4
r481 (  205 334 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.195 //y=7.4 //x2=17.28 //y2=7.4
r482 (  205 206 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=17.195 //y=7.4 //x2=16.485 //y2=7.4
r483 (  199 333 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.4 //y=7.23 //x2=16.4 //y2=7.4
r484 (  199 359 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.4 //y=7.23 //x2=16.4 //y2=6.745
r485 (  196 332 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.605 //y=7.4 //x2=15.52 //y2=7.4
r486 (  196 198 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=15.605 //y=7.4 //x2=16.28 //y2=7.4
r487 (  195 333 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.315 //y=7.4 //x2=16.4 //y2=7.4
r488 (  195 198 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=16.315 //y=7.4 //x2=16.28 //y2=7.4
r489 (  189 332 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.52 //y=7.23 //x2=15.52 //y2=7.4
r490 (  189 358 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=15.52 //y=7.23 //x2=15.52 //y2=6.405
r491 (  186 331 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.6 //y=7.4 //x2=14.43 //y2=7.4
r492 (  186 188 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.6 //y=7.4 //x2=15.17 //y2=7.4
r493 (  185 332 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.435 //y=7.4 //x2=15.52 //y2=7.4
r494 (  185 188 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=15.435 //y=7.4 //x2=15.17 //y2=7.4
r495 (  180 330 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.435 //y=7.4 //x2=13.35 //y2=7.4
r496 (  180 182 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=13.435 //y=7.4 //x2=13.69 //y2=7.4
r497 (  179 331 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.26 //y=7.4 //x2=14.43 //y2=7.4
r498 (  179 182 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=14.26 //y=7.4 //x2=13.69 //y2=7.4
r499 (  173 330 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.35 //y=7.23 //x2=13.35 //y2=7.4
r500 (  173 357 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=13.35 //y=7.23 //x2=13.35 //y2=6.745
r501 (  170 329 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.555 //y=7.4 //x2=12.47 //y2=7.4
r502 (  170 172 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=12.555 //y=7.4 //x2=12.58 //y2=7.4
r503 (  169 330 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.265 //y=7.4 //x2=13.35 //y2=7.4
r504 (  169 172 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=13.265 //y=7.4 //x2=12.58 //y2=7.4
r505 (  163 329 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.47 //y=7.23 //x2=12.47 //y2=7.4
r506 (  163 356 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.47 //y=7.23 //x2=12.47 //y2=6.745
r507 (  162 328 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.675 //y=7.4 //x2=11.59 //y2=7.4
r508 (  161 329 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.385 //y=7.4 //x2=12.47 //y2=7.4
r509 (  161 162 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=12.385 //y=7.4 //x2=11.675 //y2=7.4
r510 (  155 328 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.59 //y=7.23 //x2=11.59 //y2=7.4
r511 (  155 355 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.59 //y=7.23 //x2=11.59 //y2=6.745
r512 (  152 327 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.795 //y=7.4 //x2=10.71 //y2=7.4
r513 (  152 154 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=10.795 //y=7.4 //x2=11.47 //y2=7.4
r514 (  151 328 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.505 //y=7.4 //x2=11.59 //y2=7.4
r515 (  151 154 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=11.505 //y=7.4 //x2=11.47 //y2=7.4
r516 (  145 327 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.71 //y=7.23 //x2=10.71 //y2=7.4
r517 (  145 354 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=10.71 //y=7.23 //x2=10.71 //y2=6.405
r518 (  142 326 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.79 //y=7.4 //x2=9.62 //y2=7.4
r519 (  142 144 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.79 //y=7.4 //x2=10.36 //y2=7.4
r520 (  141 327 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.625 //y=7.4 //x2=10.71 //y2=7.4
r521 (  141 144 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=10.625 //y=7.4 //x2=10.36 //y2=7.4
r522 (  136 325 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.625 //y=7.4 //x2=8.54 //y2=7.4
r523 (  136 138 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=8.625 //y=7.4 //x2=8.88 //y2=7.4
r524 (  135 326 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.45 //y=7.4 //x2=9.62 //y2=7.4
r525 (  135 138 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.45 //y=7.4 //x2=8.88 //y2=7.4
r526 (  129 325 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.54 //y=7.23 //x2=8.54 //y2=7.4
r527 (  129 353 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.54 //y=7.23 //x2=8.54 //y2=6.745
r528 (  126 324 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.745 //y=7.4 //x2=7.66 //y2=7.4
r529 (  126 128 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=7.745 //y=7.4 //x2=7.77 //y2=7.4
r530 (  125 325 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.455 //y=7.4 //x2=8.54 //y2=7.4
r531 (  125 128 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=8.455 //y=7.4 //x2=7.77 //y2=7.4
r532 (  119 324 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.66 //y=7.23 //x2=7.66 //y2=7.4
r533 (  119 352 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.66 //y=7.23 //x2=7.66 //y2=6.745
r534 (  118 323 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.865 //y=7.4 //x2=6.78 //y2=7.4
r535 (  117 324 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.575 //y=7.4 //x2=7.66 //y2=7.4
r536 (  117 118 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.575 //y=7.4 //x2=6.865 //y2=7.4
r537 (  111 323 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=7.4
r538 (  111 351 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=6.745
r539 (  108 322 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.985 //y=7.4 //x2=5.9 //y2=7.4
r540 (  108 110 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=5.985 //y=7.4 //x2=6.66 //y2=7.4
r541 (  107 323 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.78 //y2=7.4
r542 (  107 110 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.66 //y2=7.4
r543 (  101 322 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.9 //y=7.23 //x2=5.9 //y2=7.4
r544 (  101 350 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=5.9 //y=7.23 //x2=5.9 //y2=6.405
r545 (  98 321 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=4.81 //y2=7.4
r546 (  98 100 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=5.55 //y2=7.4
r547 (  97 322 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.815 //y=7.4 //x2=5.9 //y2=7.4
r548 (  97 100 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=5.815 //y=7.4 //x2=5.55 //y2=7.4
r549 (  92 320 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=3.73 //y2=7.4
r550 (  92 94 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=4.07 //y2=7.4
r551 (  91 321 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.81 //y2=7.4
r552 (  91 94 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.07 //y2=7.4
r553 (  85 320 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=7.4
r554 (  85 349 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=6.745
r555 (  82 319 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.85 //y2=7.4
r556 (  82 84 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.96 //y2=7.4
r557 (  81 320 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=3.73 //y2=7.4
r558 (  81 84 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=2.96 //y2=7.4
r559 (  75 319 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=7.4
r560 (  75 348 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=6.745
r561 (  74 318 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.055 //y=7.4 //x2=1.97 //y2=7.4
r562 (  73 319 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.85 //y2=7.4
r563 (  73 74 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.055 //y2=7.4
r564 (  67 318 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=7.4
r565 (  67 347 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=6.745
r566 (  64 317 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.09 //y2=7.4
r567 (  64 66 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.85 //y2=7.4
r568 (  63 318 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.97 //y2=7.4
r569 (  63 66 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.85 //y2=7.4
r570 (  57 317 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=7.4
r571 (  57 346 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=6.405
r572 (  53 317 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=1.09 //y2=7.4
r573 (  53 56 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=0.74 //y2=7.4
r574 (  49 314 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.12 //y=7.4 //x2=28.12 //y2=7.4
r575 (  47 304 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.01 //y=7.4 //x2=27.01 //y2=7.4
r576 (  47 49 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=27.01 //y=7.4 //x2=28.12 //y2=7.4
r577 (  45 286 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.9 //y=7.4 //x2=25.9 //y2=7.4
r578 (  45 47 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=25.9 //y=7.4 //x2=27.01 //y2=7.4
r579 (  43 276 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=7.4 //x2=24.79 //y2=7.4
r580 (  43 45 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=7.4 //x2=25.9 //y2=7.4
r581 (  41 270 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.31 //y=7.4 //x2=23.31 //y2=7.4
r582 (  41 43 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=23.31 //y=7.4 //x2=24.79 //y2=7.4
r583 (  39 260 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.2 //y=7.4 //x2=22.2 //y2=7.4
r584 (  39 41 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.2 //y=7.4 //x2=23.31 //y2=7.4
r585 (  37 242 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=7.4 //x2=21.09 //y2=7.4
r586 (  37 39 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=7.4 //x2=22.2 //y2=7.4
r587 (  35 232 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=7.4 //x2=19.98 //y2=7.4
r588 (  35 37 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=7.4 //x2=21.09 //y2=7.4
r589 (  33 226 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.5 //y=7.4 //x2=18.5 //y2=7.4
r590 (  33 35 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.5 //y=7.4 //x2=19.98 //y2=7.4
r591 (  31 216 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=7.4 //x2=17.39 //y2=7.4
r592 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=7.4 //x2=18.5 //y2=7.4
r593 (  29 198 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=7.4 //x2=16.28 //y2=7.4
r594 (  29 31 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=7.4 //x2=17.39 //y2=7.4
r595 (  27 188 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=7.4 //x2=15.17 //y2=7.4
r596 (  27 29 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=7.4 //x2=16.28 //y2=7.4
r597 (  25 182 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=13.69 //y=7.4 //x2=13.69 //y2=7.4
r598 (  25 27 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=13.69 //y=7.4 //x2=15.17 //y2=7.4
r599 (  23 172 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=7.4 //x2=12.58 //y2=7.4
r600 (  23 25 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=7.4 //x2=13.69 //y2=7.4
r601 (  21 154 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=7.4 //x2=11.47 //y2=7.4
r602 (  21 23 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=7.4 //x2=12.58 //y2=7.4
r603 (  19 144 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r604 (  19 21 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=7.4 //x2=11.47 //y2=7.4
r605 (  17 138 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.88 //y=7.4 //x2=8.88 //y2=7.4
r606 (  17 19 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.88 //y=7.4 //x2=10.36 //y2=7.4
r607 (  15 128 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=7.4 //x2=7.77 //y2=7.4
r608 (  15 17 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=7.4 //x2=8.88 //y2=7.4
r609 (  13 110 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r610 (  13 15 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.4 //x2=7.77 //y2=7.4
r611 (  11 100 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r612 (  11 13 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.66 //y2=7.4
r613 (  9 94 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=7.4 //x2=4.07 //y2=7.4
r614 (  9 11 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=7.4 //x2=5.55 //y2=7.4
r615 (  7 84 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r616 (  7 9 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r617 (  5 66 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r618 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r619 (  2 56 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r620 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_DFFSNRNX1_PCELL\%noxref_2

subckt PM_DFFSNRNX1_PCELL\%noxref_3 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 \
 63 64 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 92 94 100 101 102 \
 103 123 125 126 127 )
c237 ( 127 0 ) capacitor c=0.023087f //x=3.145 //y=5.02
c238 ( 126 0 ) capacitor c=0.023519f //x=2.265 //y=5.02
c239 ( 125 0 ) capacitor c=0.0224735f //x=1.385 //y=5.02
c240 ( 123 0 ) capacitor c=0.00853354f //x=3.395 //y=0.915
c241 ( 103 0 ) capacitor c=0.0556143f //x=11.005 //y=4.79
c242 ( 102 0 ) capacitor c=0.0293157f //x=11.295 //y=4.79
c243 ( 101 0 ) capacitor c=0.0347816f //x=10.96 //y=1.22
c244 ( 100 0 ) capacitor c=0.0187487f //x=10.96 //y=0.875
c245 ( 94 0 ) capacitor c=0.0137055f //x=10.805 //y=1.375
c246 ( 92 0 ) capacitor c=0.0149861f //x=10.805 //y=0.72
c247 ( 91 0 ) capacitor c=0.096037f //x=10.43 //y=1.915
c248 ( 90 0 ) capacitor c=0.0228993f //x=10.43 //y=1.53
c249 ( 89 0 ) capacitor c=0.0234352f //x=10.43 //y=1.22
c250 ( 88 0 ) capacitor c=0.0198724f //x=10.43 //y=0.875
c251 ( 84 0 ) capacitor c=0.06002f //x=6.195 //y=4.79
c252 ( 83 0 ) capacitor c=0.0375015f //x=6.485 //y=4.79
c253 ( 82 0 ) capacitor c=0.0347816f //x=6.15 //y=1.22
c254 ( 81 0 ) capacitor c=0.0187487f //x=6.15 //y=0.875
c255 ( 75 0 ) capacitor c=0.0137055f //x=5.995 //y=1.375
c256 ( 73 0 ) capacitor c=0.0149861f //x=5.995 //y=0.72
c257 ( 72 0 ) capacitor c=0.096037f //x=5.62 //y=1.915
c258 ( 71 0 ) capacitor c=0.0228993f //x=5.62 //y=1.53
c259 ( 70 0 ) capacitor c=0.0234352f //x=5.62 //y=1.22
c260 ( 69 0 ) capacitor c=0.0198724f //x=5.62 //y=0.875
c261 ( 68 0 ) capacitor c=0.110114f //x=11.37 //y=6.02
c262 ( 67 0 ) capacitor c=0.158956f //x=10.93 //y=6.02
c263 ( 66 0 ) capacitor c=0.110114f //x=6.56 //y=6.02
c264 ( 65 0 ) capacitor c=0.158956f //x=6.12 //y=6.02
c265 ( 62 0 ) capacitor c=0.0013314f //x=3.29 //y=5.155
c266 ( 61 0 ) capacitor c=0.00300453f //x=2.41 //y=5.155
c267 ( 54 0 ) capacitor c=0.100268f //x=10.73 //y=2.08
c268 ( 46 0 ) capacitor c=0.105472f //x=5.92 //y=2.08
c269 ( 44 0 ) capacitor c=0.114369f //x=4.07 //y=2.59
c270 ( 40 0 ) capacitor c=0.00398962f //x=3.67 //y=1.665
c271 ( 39 0 ) capacitor c=0.0137288f //x=3.985 //y=1.665
c272 ( 33 0 ) capacitor c=0.0305699f //x=3.985 //y=5.155
c273 ( 25 0 ) capacitor c=0.0214251f //x=3.205 //y=5.155
c274 ( 18 0 ) capacitor c=0.00549987f //x=1.615 //y=5.155
c275 ( 17 0 ) capacitor c=0.0209329f //x=2.325 //y=5.155
c276 ( 4 0 ) capacitor c=0.00440131f //x=6.035 //y=2.59
c277 ( 3 0 ) capacitor c=0.0870935f //x=10.615 //y=2.59
c278 ( 2 0 ) capacitor c=0.0124623f //x=4.185 //y=2.59
c279 ( 1 0 ) capacitor c=0.0300768f //x=5.805 //y=2.59
r280 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=11.295 //y=4.79 //x2=11.37 //y2=4.865
r281 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=11.295 //y=4.79 //x2=11.005 //y2=4.79
r282 (  101 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.96 //y=1.22 //x2=10.92 //y2=1.375
r283 (  100 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.96 //y=0.875 //x2=10.92 //y2=0.72
r284 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.96 //y=0.875 //x2=10.96 //y2=1.22
r285 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.93 //y=4.865 //x2=11.005 //y2=4.79
r286 (  97 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=10.93 //y=4.865 //x2=10.73 //y2=4.7
r287 (  95 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.585 //y=1.375 //x2=10.47 //y2=1.375
r288 (  94 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.805 //y=1.375 //x2=10.92 //y2=1.375
r289 (  93 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.585 //y=0.72 //x2=10.47 //y2=0.72
r290 (  92 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.805 //y=0.72 //x2=10.92 //y2=0.72
r291 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.805 //y=0.72 //x2=10.585 //y2=0.72
r292 (  91 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.915 //x2=10.73 //y2=2.08
r293 (  90 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.53 //x2=10.47 //y2=1.375
r294 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.53 //x2=10.43 //y2=1.915
r295 (  89 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.43 //y=1.22 //x2=10.47 //y2=1.375
r296 (  88 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.43 //y=0.875 //x2=10.47 //y2=0.72
r297 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.43 //y=0.875 //x2=10.43 //y2=1.22
r298 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.485 //y=4.79 //x2=6.56 //y2=4.865
r299 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=6.485 //y=4.79 //x2=6.195 //y2=4.79
r300 (  82 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.15 //y=1.22 //x2=6.11 //y2=1.375
r301 (  81 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.15 //y=0.875 //x2=6.11 //y2=0.72
r302 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.15 //y=0.875 //x2=6.15 //y2=1.22
r303 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.12 //y=4.865 //x2=6.195 //y2=4.79
r304 (  78 112 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=6.12 //y=4.865 //x2=5.92 //y2=4.7
r305 (  76 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.775 //y=1.375 //x2=5.66 //y2=1.375
r306 (  75 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.995 //y=1.375 //x2=6.11 //y2=1.375
r307 (  74 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.775 //y=0.72 //x2=5.66 //y2=0.72
r308 (  73 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.995 //y=0.72 //x2=6.11 //y2=0.72
r309 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=5.995 //y=0.72 //x2=5.775 //y2=0.72
r310 (  72 110 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.915 //x2=5.92 //y2=2.08
r311 (  71 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.53 //x2=5.66 //y2=1.375
r312 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.53 //x2=5.62 //y2=1.915
r313 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.22 //x2=5.66 //y2=1.375
r314 (  69 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=0.875 //x2=5.66 //y2=0.72
r315 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.62 //y=0.875 //x2=5.62 //y2=1.22
r316 (  68 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.37 //y=6.02 //x2=11.37 //y2=4.865
r317 (  67 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.93 //y=6.02 //x2=10.93 //y2=4.865
r318 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.56 //y=6.02 //x2=6.56 //y2=4.865
r319 (  65 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.12 //y=6.02 //x2=6.12 //y2=4.865
r320 (  64 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.695 //y=1.375 //x2=10.805 //y2=1.375
r321 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.695 //y=1.375 //x2=10.585 //y2=1.375
r322 (  63 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.375 //x2=5.995 //y2=1.375
r323 (  63 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.375 //x2=5.775 //y2=1.375
r324 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=4.7 //x2=10.73 //y2=4.7
r325 (  57 59 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.59 //x2=10.73 //y2=4.7
r326 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=2.08 //x2=10.73 //y2=2.08
r327 (  54 57 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.08 //x2=10.73 //y2=2.59
r328 (  51 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=4.7 //x2=5.92 //y2=4.7
r329 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.59 //x2=5.92 //y2=4.7
r330 (  46 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=2.08 //x2=5.92 //y2=2.08
r331 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.08 //x2=5.92 //y2=2.59
r332 (  42 44 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=4.07 //y=5.07 //x2=4.07 //y2=2.59
r333 (  41 44 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=4.07 //y=1.75 //x2=4.07 //y2=2.59
r334 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=4.07 //y2=1.75
r335 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=3.67 //y2=1.665
r336 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.67 //y2=1.665
r337 (  35 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.585 //y2=1.01
r338 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.375 //y=5.155 //x2=3.29 //y2=5.155
r339 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=4.07 //y2=5.07
r340 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=3.375 //y2=5.155
r341 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.155
r342 (  27 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.725
r343 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.495 //y=5.155 //x2=2.41 //y2=5.155
r344 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=3.29 //y2=5.155
r345 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=2.495 //y2=5.155
r346 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.155
r347 (  19 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.725
r348 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=2.41 //y2=5.155
r349 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=1.615 //y2=5.155
r350 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.615 //y2=5.155
r351 (  11 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.53 //y2=5.725
r352 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.73 //y=2.59 //x2=10.73 //y2=2.59
r353 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.92 //y=2.59 //x2=5.92 //y2=2.59
r354 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=2.59 //x2=4.07 //y2=2.59
r355 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.035 //y=2.59 //x2=5.92 //y2=2.59
r356 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=2.59 //x2=10.73 //y2=2.59
r357 (  3 4 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=2.59 //x2=6.035 //y2=2.59
r358 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.185 //y=2.59 //x2=4.07 //y2=2.59
r359 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.805 //y=2.59 //x2=5.92 //y2=2.59
r360 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=5.805 //y=2.59 //x2=4.185 //y2=2.59
ends PM_DFFSNRNX1_PCELL\%noxref_3

subckt PM_DFFSNRNX1_PCELL\%noxref_4 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 \
 53 54 55 56 57 58 60 66 67 68 69 81 83 84 85 )
c162 ( 85 0 ) capacitor c=0.023087f //x=12.765 //y=5.02
c163 ( 84 0 ) capacitor c=0.023519f //x=11.885 //y=5.02
c164 ( 83 0 ) capacitor c=0.0224735f //x=11.005 //y=5.02
c165 ( 81 0 ) capacitor c=0.00853354f //x=13.015 //y=0.915
c166 ( 69 0 ) capacitor c=0.0556143f //x=15.815 //y=4.79
c167 ( 68 0 ) capacitor c=0.0293157f //x=16.105 //y=4.79
c168 ( 67 0 ) capacitor c=0.0347816f //x=15.77 //y=1.22
c169 ( 66 0 ) capacitor c=0.0187487f //x=15.77 //y=0.875
c170 ( 60 0 ) capacitor c=0.0137055f //x=15.615 //y=1.375
c171 ( 58 0 ) capacitor c=0.0149861f //x=15.615 //y=0.72
c172 ( 57 0 ) capacitor c=0.096037f //x=15.24 //y=1.915
c173 ( 56 0 ) capacitor c=0.0228993f //x=15.24 //y=1.53
c174 ( 55 0 ) capacitor c=0.0234352f //x=15.24 //y=1.22
c175 ( 54 0 ) capacitor c=0.0198724f //x=15.24 //y=0.875
c176 ( 53 0 ) capacitor c=0.110114f //x=16.18 //y=6.02
c177 ( 52 0 ) capacitor c=0.158956f //x=15.74 //y=6.02
c178 ( 50 0 ) capacitor c=0.00106608f //x=12.91 //y=5.155
c179 ( 49 0 ) capacitor c=0.00207319f //x=12.03 //y=5.155
c180 ( 42 0 ) capacitor c=0.0970641f //x=15.54 //y=2.08
c181 ( 40 0 ) capacitor c=0.106809f //x=13.69 //y=2.59
c182 ( 36 0 ) capacitor c=0.00398962f //x=13.29 //y=1.665
c183 ( 35 0 ) capacitor c=0.0137288f //x=13.605 //y=1.665
c184 ( 29 0 ) capacitor c=0.0283082f //x=13.605 //y=5.155
c185 ( 21 0 ) capacitor c=0.0176454f //x=12.825 //y=5.155
c186 ( 14 0 ) capacitor c=0.00332903f //x=11.235 //y=5.155
c187 ( 13 0 ) capacitor c=0.0148427f //x=11.945 //y=5.155
c188 ( 2 0 ) capacitor c=0.00808366f //x=13.805 //y=2.59
c189 ( 1 0 ) capacitor c=0.0352679f //x=15.425 //y=2.59
r190 (  68 70 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=16.105 //y=4.79 //x2=16.18 //y2=4.865
r191 (  68 69 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=16.105 //y=4.79 //x2=15.815 //y2=4.79
r192 (  67 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.77 //y=1.22 //x2=15.73 //y2=1.375
r193 (  66 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.77 //y=0.875 //x2=15.73 //y2=0.72
r194 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.77 //y=0.875 //x2=15.77 //y2=1.22
r195 (  63 69 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.74 //y=4.865 //x2=15.815 //y2=4.79
r196 (  63 78 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=15.74 //y=4.865 //x2=15.54 //y2=4.7
r197 (  61 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.395 //y=1.375 //x2=15.28 //y2=1.375
r198 (  60 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.615 //y=1.375 //x2=15.73 //y2=1.375
r199 (  59 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.395 //y=0.72 //x2=15.28 //y2=0.72
r200 (  58 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.615 //y=0.72 //x2=15.73 //y2=0.72
r201 (  58 59 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=15.615 //y=0.72 //x2=15.395 //y2=0.72
r202 (  57 76 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.915 //x2=15.54 //y2=2.08
r203 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.53 //x2=15.28 //y2=1.375
r204 (  56 57 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.53 //x2=15.24 //y2=1.915
r205 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.24 //y=1.22 //x2=15.28 //y2=1.375
r206 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.24 //y=0.875 //x2=15.28 //y2=0.72
r207 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.24 //y=0.875 //x2=15.24 //y2=1.22
r208 (  53 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.18 //y=6.02 //x2=16.18 //y2=4.865
r209 (  52 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.74 //y=6.02 //x2=15.74 //y2=4.865
r210 (  51 60 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.505 //y=1.375 //x2=15.615 //y2=1.375
r211 (  51 61 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.505 //y=1.375 //x2=15.395 //y2=1.375
r212 (  47 78 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.54 //y=4.7 //x2=15.54 //y2=4.7
r213 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=15.54 //y=2.59 //x2=15.54 //y2=4.7
r214 (  42 76 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.54 //y=2.08 //x2=15.54 //y2=2.08
r215 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=15.54 //y=2.08 //x2=15.54 //y2=2.59
r216 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=13.69 //y=5.07 //x2=13.69 //y2=2.59
r217 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=13.69 //y=1.75 //x2=13.69 //y2=2.59
r218 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.605 //y=1.665 //x2=13.69 //y2=1.75
r219 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=13.605 //y=1.665 //x2=13.29 //y2=1.665
r220 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.205 //y=1.58 //x2=13.29 //y2=1.665
r221 (  31 81 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=13.205 //y=1.58 //x2=13.205 //y2=1.01
r222 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.995 //y=5.155 //x2=12.91 //y2=5.155
r223 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=13.605 //y=5.155 //x2=13.69 //y2=5.07
r224 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=13.605 //y=5.155 //x2=12.995 //y2=5.155
r225 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.91 //y=5.24 //x2=12.91 //y2=5.155
r226 (  23 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.91 //y=5.24 //x2=12.91 //y2=5.725
r227 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.115 //y=5.155 //x2=12.03 //y2=5.155
r228 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.825 //y=5.155 //x2=12.91 //y2=5.155
r229 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=12.825 //y=5.155 //x2=12.115 //y2=5.155
r230 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.03 //y=5.24 //x2=12.03 //y2=5.155
r231 (  15 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.03 //y=5.24 //x2=12.03 //y2=5.725
r232 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.945 //y=5.155 //x2=12.03 //y2=5.155
r233 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.945 //y=5.155 //x2=11.235 //y2=5.155
r234 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.15 //y=5.24 //x2=11.235 //y2=5.155
r235 (  7 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.15 //y=5.24 //x2=11.15 //y2=5.725
r236 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.54 //y=2.59 //x2=15.54 //y2=2.59
r237 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=13.69 //y=2.59 //x2=13.69 //y2=2.59
r238 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.805 //y=2.59 //x2=13.69 //y2=2.59
r239 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.425 //y=2.59 //x2=15.54 //y2=2.59
r240 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=15.425 //y=2.59 //x2=13.805 //y2=2.59
ends PM_DFFSNRNX1_PCELL\%noxref_4

subckt PM_DFFSNRNX1_PCELL\%noxref_5 ( 1 2 8 16 23 24 25 26 27 28 29 30 31 33 \
 39 40 41 42 43 48 49 50 52 58 59 60 61 62 70 81 )
c204 ( 81 0 ) capacitor c=0.0334842f //x=16.65 //y=4.7
c205 ( 70 0 ) capacitor c=0.0334842f //x=7.03 //y=4.7
c206 ( 62 0 ) capacitor c=0.0255071f //x=16.985 //y=4.79
c207 ( 61 0 ) capacitor c=0.0825763f //x=16.74 //y=1.915
c208 ( 60 0 ) capacitor c=0.0170266f //x=16.74 //y=1.45
c209 ( 59 0 ) capacitor c=0.018609f //x=16.74 //y=1.22
c210 ( 58 0 ) capacitor c=0.0187309f //x=16.74 //y=0.91
c211 ( 52 0 ) capacitor c=0.014725f //x=16.585 //y=1.375
c212 ( 50 0 ) capacitor c=0.0146567f //x=16.585 //y=0.755
c213 ( 49 0 ) capacitor c=0.0335408f //x=16.215 //y=1.22
c214 ( 48 0 ) capacitor c=0.0173761f //x=16.215 //y=0.91
c215 ( 43 0 ) capacitor c=0.0245352f //x=7.365 //y=4.79
c216 ( 42 0 ) capacitor c=0.0825763f //x=7.12 //y=1.915
c217 ( 41 0 ) capacitor c=0.0170266f //x=7.12 //y=1.45
c218 ( 40 0 ) capacitor c=0.018609f //x=7.12 //y=1.22
c219 ( 39 0 ) capacitor c=0.0187309f //x=7.12 //y=0.91
c220 ( 33 0 ) capacitor c=0.014725f //x=6.965 //y=1.375
c221 ( 31 0 ) capacitor c=0.0146567f //x=6.965 //y=0.755
c222 ( 30 0 ) capacitor c=0.0335408f //x=6.595 //y=1.22
c223 ( 29 0 ) capacitor c=0.0173761f //x=6.595 //y=0.91
c224 ( 28 0 ) capacitor c=0.110114f //x=17.06 //y=6.02
c225 ( 27 0 ) capacitor c=0.11012f //x=16.62 //y=6.02
c226 ( 26 0 ) capacitor c=0.110114f //x=7.44 //y=6.02
c227 ( 25 0 ) capacitor c=0.11012f //x=7 //y=6.02
c228 ( 16 0 ) capacitor c=0.0926307f //x=16.65 //y=2.08
c229 ( 8 0 ) capacitor c=0.0951701f //x=7.03 //y=2.08
c230 ( 2 0 ) capacitor c=0.0161259f //x=7.145 //y=4.44
c231 ( 1 0 ) capacitor c=0.263506f //x=16.535 //y=4.44
r232 (  83 84 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=16.65 //y=4.79 //x2=16.65 //y2=4.865
r233 (  81 83 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=16.65 //y=4.7 //x2=16.65 //y2=4.79
r234 (  72 73 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=7.03 //y=4.79 //x2=7.03 //y2=4.865
r235 (  70 72 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=7.03 //y=4.7 //x2=7.03 //y2=4.79
r236 (  63 83 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=16.785 //y=4.79 //x2=16.65 //y2=4.79
r237 (  62 64 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=16.985 //y=4.79 //x2=17.06 //y2=4.865
r238 (  62 63 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=16.985 //y=4.79 //x2=16.785 //y2=4.79
r239 (  61 88 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.915 //x2=16.665 //y2=2.08
r240 (  60 86 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.45 //x2=16.7 //y2=1.375
r241 (  60 61 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.45 //x2=16.74 //y2=1.915
r242 (  59 86 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.74 //y=1.22 //x2=16.7 //y2=1.375
r243 (  58 85 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.74 //y=0.91 //x2=16.7 //y2=0.755
r244 (  58 59 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=16.74 //y=0.91 //x2=16.74 //y2=1.22
r245 (  53 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.37 //y=1.375 //x2=16.255 //y2=1.375
r246 (  52 86 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.585 //y=1.375 //x2=16.7 //y2=1.375
r247 (  51 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.37 //y=0.755 //x2=16.255 //y2=0.755
r248 (  50 85 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.585 //y=0.755 //x2=16.7 //y2=0.755
r249 (  50 51 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=16.585 //y=0.755 //x2=16.37 //y2=0.755
r250 (  49 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.215 //y=1.22 //x2=16.255 //y2=1.375
r251 (  48 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.215 //y=0.91 //x2=16.255 //y2=0.755
r252 (  48 49 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=16.215 //y=0.91 //x2=16.215 //y2=1.22
r253 (  44 72 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=7.165 //y=4.79 //x2=7.03 //y2=4.79
r254 (  43 45 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.365 //y=4.79 //x2=7.44 //y2=4.865
r255 (  43 44 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=7.365 //y=4.79 //x2=7.165 //y2=4.79
r256 (  42 77 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.915 //x2=7.045 //y2=2.08
r257 (  41 75 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.45 //x2=7.08 //y2=1.375
r258 (  41 42 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.45 //x2=7.12 //y2=1.915
r259 (  40 75 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.22 //x2=7.08 //y2=1.375
r260 (  39 74 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.12 //y=0.91 //x2=7.08 //y2=0.755
r261 (  39 40 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=7.12 //y=0.91 //x2=7.12 //y2=1.22
r262 (  34 68 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.75 //y=1.375 //x2=6.635 //y2=1.375
r263 (  33 75 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.965 //y=1.375 //x2=7.08 //y2=1.375
r264 (  32 67 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.75 //y=0.755 //x2=6.635 //y2=0.755
r265 (  31 74 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.965 //y=0.755 //x2=7.08 //y2=0.755
r266 (  31 32 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=6.965 //y=0.755 //x2=6.75 //y2=0.755
r267 (  30 68 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.595 //y=1.22 //x2=6.635 //y2=1.375
r268 (  29 67 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.595 //y=0.91 //x2=6.635 //y2=0.755
r269 (  29 30 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=6.595 //y=0.91 //x2=6.595 //y2=1.22
r270 (  28 64 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.06 //y=6.02 //x2=17.06 //y2=4.865
r271 (  27 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.62 //y=6.02 //x2=16.62 //y2=4.865
r272 (  26 45 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.44 //y=6.02 //x2=7.44 //y2=4.865
r273 (  25 73 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7 //y=6.02 //x2=7 //y2=4.865
r274 (  24 52 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=16.477 //y=1.375 //x2=16.585 //y2=1.375
r275 (  24 53 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=16.477 //y=1.375 //x2=16.37 //y2=1.375
r276 (  23 33 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=6.857 //y=1.375 //x2=6.965 //y2=1.375
r277 (  23 34 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=6.857 //y=1.375 //x2=6.75 //y2=1.375
r278 (  21 81 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.65 //y=4.7 //x2=16.65 //y2=4.7
r279 (  19 21 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=16.65 //y=4.44 //x2=16.65 //y2=4.7
r280 (  16 88 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.65 //y=2.08 //x2=16.65 //y2=2.08
r281 (  16 19 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=16.65 //y=2.08 //x2=16.65 //y2=4.44
r282 (  13 70 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.03 //y=4.7 //x2=7.03 //y2=4.7
r283 (  11 13 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=7.03 //y=4.44 //x2=7.03 //y2=4.7
r284 (  8 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.03 //y=2.08 //x2=7.03 //y2=2.08
r285 (  8 11 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li //thickness=0.1 \
 //x=7.03 //y=2.08 //x2=7.03 //y2=4.44
r286 (  6 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=16.65 //y=4.44 //x2=16.65 //y2=4.44
r287 (  4 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.03 //y=4.44 //x2=7.03 //y2=4.44
r288 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.145 //y=4.44 //x2=7.03 //y2=4.44
r289 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.535 //y=4.44 //x2=16.65 //y2=4.44
r290 (  1 2 ) resistor r=8.95992 //w=0.131 //l=9.39 //layer=m1 \
 //thickness=0.36 //x=16.535 //y=4.44 //x2=7.145 //y2=4.44
ends PM_DFFSNRNX1_PCELL\%noxref_5

subckt PM_DFFSNRNX1_PCELL\%noxref_6 ( 1 2 3 4 12 25 26 33 41 47 48 52 54 61 62 \
 63 64 65 66 67 68 72 73 74 79 81 84 85 86 87 88 89 90 92 98 99 100 101 106 \
 107 112 123 125 126 127 )
c264 ( 127 0 ) capacitor c=0.023087f //x=7.955 //y=5.02
c265 ( 126 0 ) capacitor c=0.023519f //x=7.075 //y=5.02
c266 ( 125 0 ) capacitor c=0.0224735f //x=6.195 //y=5.02
c267 ( 123 0 ) capacitor c=0.00853354f //x=8.205 //y=0.915
c268 ( 112 0 ) capacitor c=0.0672371f //x=3.33 //y=4.7
c269 ( 107 0 ) capacitor c=0.0273931f //x=3.33 //y=1.915
c270 ( 106 0 ) capacitor c=0.045877f //x=3.33 //y=2.08
c271 ( 101 0 ) capacitor c=0.0562318f //x=20.625 //y=4.79
c272 ( 100 0 ) capacitor c=0.0305765f //x=20.915 //y=4.79
c273 ( 99 0 ) capacitor c=0.0347816f //x=20.58 //y=1.22
c274 ( 98 0 ) capacitor c=0.0187487f //x=20.58 //y=0.875
c275 ( 92 0 ) capacitor c=0.0137055f //x=20.425 //y=1.375
c276 ( 90 0 ) capacitor c=0.0149861f //x=20.425 //y=0.72
c277 ( 89 0 ) capacitor c=0.096037f //x=20.05 //y=1.915
c278 ( 88 0 ) capacitor c=0.0228993f //x=20.05 //y=1.53
c279 ( 87 0 ) capacitor c=0.0234352f //x=20.05 //y=1.22
c280 ( 86 0 ) capacitor c=0.0198724f //x=20.05 //y=0.875
c281 ( 85 0 ) capacitor c=0.0432517f //x=3.85 //y=1.26
c282 ( 84 0 ) capacitor c=0.0200379f //x=3.85 //y=0.915
c283 ( 81 0 ) capacitor c=0.0148873f //x=3.695 //y=1.415
c284 ( 79 0 ) capacitor c=0.0157803f //x=3.695 //y=0.76
c285 ( 74 0 ) capacitor c=0.0218028f //x=3.32 //y=1.57
c286 ( 73 0 ) capacitor c=0.0207459f //x=3.32 //y=1.26
c287 ( 72 0 ) capacitor c=0.0194308f //x=3.32 //y=0.915
c288 ( 68 0 ) capacitor c=0.110114f //x=20.99 //y=6.02
c289 ( 67 0 ) capacitor c=0.158956f //x=20.55 //y=6.02
c290 ( 66 0 ) capacitor c=0.158794f //x=3.51 //y=6.02
c291 ( 65 0 ) capacitor c=0.110114f //x=3.07 //y=6.02
c292 ( 62 0 ) capacitor c=0.00106608f //x=8.1 //y=5.155
c293 ( 61 0 ) capacitor c=0.00207162f //x=7.22 //y=5.155
c294 ( 54 0 ) capacitor c=0.101888f //x=20.35 //y=2.08
c295 ( 52 0 ) capacitor c=0.109321f //x=8.88 //y=3.33
c296 ( 48 0 ) capacitor c=0.00398962f //x=8.48 //y=1.665
c297 ( 47 0 ) capacitor c=0.0137288f //x=8.795 //y=1.665
c298 ( 41 0 ) capacitor c=0.0283082f //x=8.795 //y=5.155
c299 ( 33 0 ) capacitor c=0.0176454f //x=8.015 //y=5.155
c300 ( 26 0 ) capacitor c=0.00385842f //x=6.425 //y=5.155
c301 ( 25 0 ) capacitor c=0.016487f //x=7.135 //y=5.155
c302 ( 12 0 ) capacitor c=0.0907612f //x=3.33 //y=2.08
c303 ( 4 0 ) capacitor c=0.00578611f //x=8.995 //y=3.33
c304 ( 3 0 ) capacitor c=0.189113f //x=20.235 //y=3.33
c305 ( 2 0 ) capacitor c=0.0166611f //x=3.445 //y=3.33
c306 ( 1 0 ) capacitor c=0.156035f //x=8.765 //y=3.33
r307 (  106 107 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.33 //y=2.08 //x2=3.33 //y2=1.915
r308 (  100 102 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.915 //y=4.79 //x2=20.99 //y2=4.865
r309 (  100 101 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=20.915 //y=4.79 //x2=20.625 //y2=4.79
r310 (  99 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.58 //y=1.22 //x2=20.54 //y2=1.375
r311 (  98 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.58 //y=0.875 //x2=20.54 //y2=0.72
r312 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.58 //y=0.875 //x2=20.58 //y2=1.22
r313 (  95 101 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.55 //y=4.865 //x2=20.625 //y2=4.79
r314 (  95 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=20.55 //y=4.865 //x2=20.35 //y2=4.7
r315 (  93 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.205 //y=1.375 //x2=20.09 //y2=1.375
r316 (  92 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.425 //y=1.375 //x2=20.54 //y2=1.375
r317 (  91 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.205 //y=0.72 //x2=20.09 //y2=0.72
r318 (  90 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.425 //y=0.72 //x2=20.54 //y2=0.72
r319 (  90 91 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=20.425 //y=0.72 //x2=20.205 //y2=0.72
r320 (  89 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.915 //x2=20.35 //y2=2.08
r321 (  88 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.53 //x2=20.09 //y2=1.375
r322 (  88 89 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.53 //x2=20.05 //y2=1.915
r323 (  87 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.05 //y=1.22 //x2=20.09 //y2=1.375
r324 (  86 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.05 //y=0.875 //x2=20.09 //y2=0.72
r325 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.05 //y=0.875 //x2=20.05 //y2=1.22
r326 (  85 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=1.26 //x2=3.81 //y2=1.415
r327 (  84 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.81 //y2=0.76
r328 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.85 //y2=1.26
r329 (  82 110 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=1.415 //x2=3.36 //y2=1.415
r330 (  81 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=1.415 //x2=3.81 //y2=1.415
r331 (  80 109 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=0.76 //x2=3.36 //y2=0.76
r332 (  79 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.81 //y2=0.76
r333 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.475 //y2=0.76
r334 (  76 112 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=3.51 //y=4.865 //x2=3.33 //y2=4.7
r335 (  74 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.36 //y2=1.415
r336 (  74 107 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.32 //y2=1.915
r337 (  73 110 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.26 //x2=3.36 //y2=1.415
r338 (  72 109 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.36 //y2=0.76
r339 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.32 //y2=1.26
r340 (  69 112 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=3.07 //y=4.865 //x2=3.33 //y2=4.7
r341 (  68 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.99 //y=6.02 //x2=20.99 //y2=4.865
r342 (  67 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.55 //y=6.02 //x2=20.55 //y2=4.865
r343 (  66 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.51 //y=6.02 //x2=3.51 //y2=4.865
r344 (  65 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.07 //y=6.02 //x2=3.07 //y2=4.865
r345 (  64 92 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.315 //y=1.375 //x2=20.425 //y2=1.375
r346 (  64 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.315 //y=1.375 //x2=20.205 //y2=1.375
r347 (  63 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.695 //y2=1.415
r348 (  63 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.475 //y2=1.415
r349 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.35 //y=4.7 //x2=20.35 //y2=4.7
r350 (  57 59 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=20.35 //y=3.33 //x2=20.35 //y2=4.7
r351 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.35 //y=2.08 //x2=20.35 //y2=2.08
r352 (  54 57 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=20.35 //y=2.08 //x2=20.35 //y2=3.33
r353 (  50 52 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=8.88 //y=5.07 //x2=8.88 //y2=3.33
r354 (  49 52 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=8.88 //y=1.75 //x2=8.88 //y2=3.33
r355 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.795 //y=1.665 //x2=8.88 //y2=1.75
r356 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=8.795 //y=1.665 //x2=8.48 //y2=1.665
r357 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.395 //y=1.58 //x2=8.48 //y2=1.665
r358 (  43 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=8.395 //y=1.58 //x2=8.395 //y2=1.01
r359 (  42 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.185 //y=5.155 //x2=8.1 //y2=5.155
r360 (  41 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.795 //y=5.155 //x2=8.88 //y2=5.07
r361 (  41 42 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=8.795 //y=5.155 //x2=8.185 //y2=5.155
r362 (  35 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.1 //y=5.24 //x2=8.1 //y2=5.155
r363 (  35 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.1 //y=5.24 //x2=8.1 //y2=5.725
r364 (  34 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.305 //y=5.155 //x2=7.22 //y2=5.155
r365 (  33 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.015 //y=5.155 //x2=8.1 //y2=5.155
r366 (  33 34 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.015 //y=5.155 //x2=7.305 //y2=5.155
r367 (  27 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.24 //x2=7.22 //y2=5.155
r368 (  27 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.24 //x2=7.22 //y2=5.725
r369 (  25 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.155 //x2=7.22 //y2=5.155
r370 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.155 //x2=6.425 //y2=5.155
r371 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.24 //x2=6.425 //y2=5.155
r372 (  19 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.24 //x2=6.34 //y2=5.725
r373 (  17 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r374 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=3.33 //x2=3.33 //y2=4.7
r375 (  12 106 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r376 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.08 //x2=3.33 //y2=3.33
r377 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=20.35 //y=3.33 //x2=20.35 //y2=3.33
r378 (  8 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.88 //y=3.33 //x2=8.88 //y2=3.33
r379 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=3.33 //x2=3.33 //y2=3.33
r380 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.995 //y=3.33 //x2=8.88 //y2=3.33
r381 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.235 //y=3.33 //x2=20.35 //y2=3.33
r382 (  3 4 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=20.235 //y=3.33 //x2=8.995 //y2=3.33
r383 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.445 //y=3.33 //x2=3.33 //y2=3.33
r384 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=3.33 //x2=8.88 //y2=3.33
r385 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=3.33 //x2=3.445 //y2=3.33
ends PM_DFFSNRNX1_PCELL\%noxref_6

subckt PM_DFFSNRNX1_PCELL\%noxref_7 ( 1 2 3 4 12 20 28 35 36 37 38 39 40 41 42 \
 43 44 45 46 48 54 55 56 57 58 66 67 68 73 75 78 79 80 81 82 84 90 91 92 93 94 \
 102 111 112 117 123 )
c316 ( 123 0 ) capacitor c=0.0337728f //x=21.46 //y=4.7
c317 ( 117 0 ) capacitor c=0.0600797f //x=17.76 //y=4.7
c318 ( 112 0 ) capacitor c=0.0273931f //x=17.76 //y=1.915
c319 ( 111 0 ) capacitor c=0.0455604f //x=17.76 //y=2.08
c320 ( 102 0 ) capacitor c=0.0354872f //x=2.22 //y=4.7
c321 ( 94 0 ) capacitor c=0.025532f //x=21.795 //y=4.79
c322 ( 93 0 ) capacitor c=0.0827272f //x=21.55 //y=1.915
c323 ( 92 0 ) capacitor c=0.0170266f //x=21.55 //y=1.45
c324 ( 91 0 ) capacitor c=0.018609f //x=21.55 //y=1.22
c325 ( 90 0 ) capacitor c=0.0187309f //x=21.55 //y=0.91
c326 ( 84 0 ) capacitor c=0.014725f //x=21.395 //y=1.375
c327 ( 82 0 ) capacitor c=0.0146567f //x=21.395 //y=0.755
c328 ( 81 0 ) capacitor c=0.0335408f //x=21.025 //y=1.22
c329 ( 80 0 ) capacitor c=0.0173761f //x=21.025 //y=0.91
c330 ( 79 0 ) capacitor c=0.0432517f //x=18.28 //y=1.26
c331 ( 78 0 ) capacitor c=0.0200379f //x=18.28 //y=0.915
c332 ( 75 0 ) capacitor c=0.0148873f //x=18.125 //y=1.415
c333 ( 73 0 ) capacitor c=0.0157803f //x=18.125 //y=0.76
c334 ( 68 0 ) capacitor c=0.0218028f //x=17.75 //y=1.57
c335 ( 67 0 ) capacitor c=0.0207459f //x=17.75 //y=1.26
c336 ( 66 0 ) capacitor c=0.0194308f //x=17.75 //y=0.915
c337 ( 58 0 ) capacitor c=0.0307682f //x=2.555 //y=4.79
c338 ( 57 0 ) capacitor c=0.0826756f //x=2.31 //y=1.915
c339 ( 56 0 ) capacitor c=0.0170266f //x=2.31 //y=1.45
c340 ( 55 0 ) capacitor c=0.018609f //x=2.31 //y=1.22
c341 ( 54 0 ) capacitor c=0.0187309f //x=2.31 //y=0.91
c342 ( 48 0 ) capacitor c=0.014725f //x=2.155 //y=1.375
c343 ( 46 0 ) capacitor c=0.0146567f //x=2.155 //y=0.755
c344 ( 45 0 ) capacitor c=0.0335408f //x=1.785 //y=1.22
c345 ( 44 0 ) capacitor c=0.0173761f //x=1.785 //y=0.91
c346 ( 43 0 ) capacitor c=0.110114f //x=21.87 //y=6.02
c347 ( 42 0 ) capacitor c=0.11012f //x=21.43 //y=6.02
c348 ( 41 0 ) capacitor c=0.158794f //x=17.94 //y=6.02
c349 ( 40 0 ) capacitor c=0.110114f //x=17.5 //y=6.02
c350 ( 39 0 ) capacitor c=0.110114f //x=2.63 //y=6.02
c351 ( 38 0 ) capacitor c=0.11012f //x=2.19 //y=6.02
c352 ( 28 0 ) capacitor c=0.0980911f //x=21.46 //y=2.08
c353 ( 20 0 ) capacitor c=0.0858438f //x=17.76 //y=2.08
c354 ( 12 0 ) capacitor c=0.10298f //x=2.22 //y=2.08
c355 ( 4 0 ) capacitor c=0.00626813f //x=17.875 //y=2.22
c356 ( 3 0 ) capacitor c=0.0949894f //x=21.345 //y=2.22
c357 ( 2 0 ) capacitor c=0.0179508f //x=2.335 //y=2.22
c358 ( 1 0 ) capacitor c=0.340196f //x=17.645 //y=2.22
r359 (  125 126 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=21.46 //y=4.79 //x2=21.46 //y2=4.865
r360 (  123 125 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=21.46 //y=4.7 //x2=21.46 //y2=4.79
r361 (  111 112 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=17.76 //y=2.08 //x2=17.76 //y2=1.915
r362 (  104 105 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.79 //x2=2.22 //y2=4.865
r363 (  102 104 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.7 //x2=2.22 //y2=4.79
r364 (  95 125 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=21.595 //y=4.79 //x2=21.46 //y2=4.79
r365 (  94 96 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=21.795 //y=4.79 //x2=21.87 //y2=4.865
r366 (  94 95 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=21.795 //y=4.79 //x2=21.595 //y2=4.79
r367 (  93 130 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.915 //x2=21.475 //y2=2.08
r368 (  92 128 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.45 //x2=21.51 //y2=1.375
r369 (  92 93 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.45 //x2=21.55 //y2=1.915
r370 (  91 128 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.22 //x2=21.51 //y2=1.375
r371 (  90 127 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.55 //y=0.91 //x2=21.51 //y2=0.755
r372 (  90 91 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.55 //y=0.91 //x2=21.55 //y2=1.22
r373 (  85 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.18 //y=1.375 //x2=21.065 //y2=1.375
r374 (  84 128 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.395 //y=1.375 //x2=21.51 //y2=1.375
r375 (  83 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.18 //y=0.755 //x2=21.065 //y2=0.755
r376 (  82 127 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.755 //x2=21.51 //y2=0.755
r377 (  82 83 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.755 //x2=21.18 //y2=0.755
r378 (  81 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.025 //y=1.22 //x2=21.065 //y2=1.375
r379 (  80 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.025 //y=0.91 //x2=21.065 //y2=0.755
r380 (  80 81 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.025 //y=0.91 //x2=21.025 //y2=1.22
r381 (  79 119 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.28 //y=1.26 //x2=18.24 //y2=1.415
r382 (  78 118 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.28 //y=0.915 //x2=18.24 //y2=0.76
r383 (  78 79 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.28 //y=0.915 //x2=18.28 //y2=1.26
r384 (  76 115 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.905 //y=1.415 //x2=17.79 //y2=1.415
r385 (  75 119 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.125 //y=1.415 //x2=18.24 //y2=1.415
r386 (  74 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.905 //y=0.76 //x2=17.79 //y2=0.76
r387 (  73 118 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.125 //y=0.76 //x2=18.24 //y2=0.76
r388 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=18.125 //y=0.76 //x2=17.905 //y2=0.76
r389 (  70 117 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=17.94 //y=4.865 //x2=17.76 //y2=4.7
r390 (  68 115 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.75 //y=1.57 //x2=17.79 //y2=1.415
r391 (  68 112 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.75 //y=1.57 //x2=17.75 //y2=1.915
r392 (  67 115 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.75 //y=1.26 //x2=17.79 //y2=1.415
r393 (  66 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.75 //y=0.915 //x2=17.79 //y2=0.76
r394 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.75 //y=0.915 //x2=17.75 //y2=1.26
r395 (  63 117 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=17.5 //y=4.865 //x2=17.76 //y2=4.7
r396 (  59 104 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.355 //y=4.79 //x2=2.22 //y2=4.79
r397 (  58 60 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.63 //y2=4.865
r398 (  58 59 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.355 //y2=4.79
r399 (  57 109 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.915 //x2=2.235 //y2=2.08
r400 (  56 107 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.27 //y2=1.375
r401 (  56 57 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.31 //y2=1.915
r402 (  55 107 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.22 //x2=2.27 //y2=1.375
r403 (  54 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.27 //y2=0.755
r404 (  54 55 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.31 //y2=1.22
r405 (  49 100 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=1.375 //x2=1.825 //y2=1.375
r406 (  48 107 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=1.375 //x2=2.27 //y2=1.375
r407 (  47 99 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=0.755 //x2=1.825 //y2=0.755
r408 (  46 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=2.27 //y2=0.755
r409 (  46 47 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=1.94 //y2=0.755
r410 (  45 100 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=1.22 //x2=1.825 //y2=1.375
r411 (  44 99 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.825 //y2=0.755
r412 (  44 45 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.785 //y2=1.22
r413 (  43 96 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.87 //y=6.02 //x2=21.87 //y2=4.865
r414 (  42 126 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.43 //y=6.02 //x2=21.43 //y2=4.865
r415 (  41 70 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.94 //y=6.02 //x2=17.94 //y2=4.865
r416 (  40 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.5 //y=6.02 //x2=17.5 //y2=4.865
r417 (  39 60 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.63 //y=6.02 //x2=2.63 //y2=4.865
r418 (  38 105 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.19 //y=6.02 //x2=2.19 //y2=4.865
r419 (  37 84 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=21.287 //y=1.375 //x2=21.395 //y2=1.375
r420 (  37 85 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=21.287 //y=1.375 //x2=21.18 //y2=1.375
r421 (  36 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.015 //y=1.415 //x2=18.125 //y2=1.415
r422 (  36 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.015 //y=1.415 //x2=17.905 //y2=1.415
r423 (  35 48 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=2.155 //y2=1.375
r424 (  35 49 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=1.94 //y2=1.375
r425 (  33 123 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.46 //y=4.7 //x2=21.46 //y2=4.7
r426 (  31 33 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.22 //x2=21.46 //y2=4.7
r427 (  28 130 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.46 //y=2.08 //x2=21.46 //y2=2.08
r428 (  28 31 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=21.46 //y=2.08 //x2=21.46 //y2=2.22
r429 (  25 117 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.76 //y=4.7 //x2=17.76 //y2=4.7
r430 (  23 25 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.22 //x2=17.76 //y2=4.7
r431 (  20 111 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.76 //y=2.08 //x2=17.76 //y2=2.08
r432 (  20 23 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=17.76 //y=2.08 //x2=17.76 //y2=2.22
r433 (  17 102 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=4.7 //x2=2.22 //y2=4.7
r434 (  15 17 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.22 //x2=2.22 //y2=4.7
r435 (  12 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=2.08
r436 (  12 15 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.08 //x2=2.22 //y2=2.22
r437 (  10 31 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.46 //y=2.22 //x2=21.46 //y2=2.22
r438 (  8 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.76 //y=2.22 //x2=17.76 //y2=2.22
r439 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.22 //y=2.22 //x2=2.22 //y2=2.22
r440 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.875 //y=2.22 //x2=17.76 //y2=2.22
r441 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=2.22 //x2=21.46 //y2=2.22
r442 (  3 4 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=21.345 //y=2.22 //x2=17.875 //y2=2.22
r443 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.335 //y=2.22 //x2=2.22 //y2=2.22
r444 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.645 //y=2.22 //x2=17.76 //y2=2.22
r445 (  1 2 ) resistor r=14.6088 //w=0.131 //l=15.31 //layer=m1 \
 //thickness=0.36 //x=17.645 //y=2.22 //x2=2.335 //y2=2.22
ends PM_DFFSNRNX1_PCELL\%noxref_7

subckt PM_DFFSNRNX1_PCELL\%noxref_8 ( 1 2 8 16 23 24 25 26 27 28 29 30 31 33 \
 39 40 41 42 43 48 49 50 52 58 59 60 61 62 70 81 )
c201 ( 81 0 ) capacitor c=0.0337728f //x=26.27 //y=4.7
c202 ( 70 0 ) capacitor c=0.0335551f //x=11.84 //y=4.7
c203 ( 62 0 ) capacitor c=0.025532f //x=26.605 //y=4.79
c204 ( 61 0 ) capacitor c=0.0832009f //x=26.36 //y=1.915
c205 ( 60 0 ) capacitor c=0.0170266f //x=26.36 //y=1.45
c206 ( 59 0 ) capacitor c=0.018609f //x=26.36 //y=1.22
c207 ( 58 0 ) capacitor c=0.0187309f //x=26.36 //y=0.91
c208 ( 52 0 ) capacitor c=0.014725f //x=26.205 //y=1.375
c209 ( 50 0 ) capacitor c=0.0146567f //x=26.205 //y=0.755
c210 ( 49 0 ) capacitor c=0.0335408f //x=25.835 //y=1.22
c211 ( 48 0 ) capacitor c=0.0173761f //x=25.835 //y=0.91
c212 ( 43 0 ) capacitor c=0.0245352f //x=12.175 //y=4.79
c213 ( 42 0 ) capacitor c=0.0825763f //x=11.93 //y=1.915
c214 ( 41 0 ) capacitor c=0.0170266f //x=11.93 //y=1.45
c215 ( 40 0 ) capacitor c=0.018609f //x=11.93 //y=1.22
c216 ( 39 0 ) capacitor c=0.0187309f //x=11.93 //y=0.91
c217 ( 33 0 ) capacitor c=0.014725f //x=11.775 //y=1.375
c218 ( 31 0 ) capacitor c=0.0146567f //x=11.775 //y=0.755
c219 ( 30 0 ) capacitor c=0.0335408f //x=11.405 //y=1.22
c220 ( 29 0 ) capacitor c=0.0173761f //x=11.405 //y=0.91
c221 ( 28 0 ) capacitor c=0.110114f //x=26.68 //y=6.02
c222 ( 27 0 ) capacitor c=0.11012f //x=26.24 //y=6.02
c223 ( 26 0 ) capacitor c=0.110114f //x=12.25 //y=6.02
c224 ( 25 0 ) capacitor c=0.11012f //x=11.81 //y=6.02
c225 ( 16 0 ) capacitor c=0.10144f //x=26.27 //y=2.08
c226 ( 8 0 ) capacitor c=0.0921574f //x=11.84 //y=2.08
c227 ( 2 0 ) capacitor c=0.0141295f //x=11.955 //y=2.96
c228 ( 1 0 ) capacitor c=0.307352f //x=26.155 //y=2.96
r229 (  83 84 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=26.27 //y=4.79 //x2=26.27 //y2=4.865
r230 (  81 83 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=26.27 //y=4.7 //x2=26.27 //y2=4.79
r231 (  72 73 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=11.84 //y=4.79 //x2=11.84 //y2=4.865
r232 (  70 72 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=11.84 //y=4.7 //x2=11.84 //y2=4.79
r233 (  63 83 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=26.405 //y=4.79 //x2=26.27 //y2=4.79
r234 (  62 64 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=26.605 //y=4.79 //x2=26.68 //y2=4.865
r235 (  62 63 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=26.605 //y=4.79 //x2=26.405 //y2=4.79
r236 (  61 88 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.915 //x2=26.285 //y2=2.08
r237 (  60 86 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.45 //x2=26.32 //y2=1.375
r238 (  60 61 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.45 //x2=26.36 //y2=1.915
r239 (  59 86 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.36 //y=1.22 //x2=26.32 //y2=1.375
r240 (  58 85 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.36 //y=0.91 //x2=26.32 //y2=0.755
r241 (  58 59 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=26.36 //y=0.91 //x2=26.36 //y2=1.22
r242 (  53 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.99 //y=1.375 //x2=25.875 //y2=1.375
r243 (  52 86 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.205 //y=1.375 //x2=26.32 //y2=1.375
r244 (  51 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.99 //y=0.755 //x2=25.875 //y2=0.755
r245 (  50 85 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.205 //y=0.755 //x2=26.32 //y2=0.755
r246 (  50 51 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=26.205 //y=0.755 //x2=25.99 //y2=0.755
r247 (  49 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.835 //y=1.22 //x2=25.875 //y2=1.375
r248 (  48 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.835 //y=0.91 //x2=25.875 //y2=0.755
r249 (  48 49 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=25.835 //y=0.91 //x2=25.835 //y2=1.22
r250 (  44 72 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=11.975 //y=4.79 //x2=11.84 //y2=4.79
r251 (  43 45 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=12.175 //y=4.79 //x2=12.25 //y2=4.865
r252 (  43 44 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=12.175 //y=4.79 //x2=11.975 //y2=4.79
r253 (  42 77 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.915 //x2=11.855 //y2=2.08
r254 (  41 75 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.45 //x2=11.89 //y2=1.375
r255 (  41 42 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.45 //x2=11.93 //y2=1.915
r256 (  40 75 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.93 //y=1.22 //x2=11.89 //y2=1.375
r257 (  39 74 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.93 //y=0.91 //x2=11.89 //y2=0.755
r258 (  39 40 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=11.93 //y=0.91 //x2=11.93 //y2=1.22
r259 (  34 68 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.56 //y=1.375 //x2=11.445 //y2=1.375
r260 (  33 75 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.775 //y=1.375 //x2=11.89 //y2=1.375
r261 (  32 67 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.56 //y=0.755 //x2=11.445 //y2=0.755
r262 (  31 74 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.775 //y=0.755 //x2=11.89 //y2=0.755
r263 (  31 32 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=11.775 //y=0.755 //x2=11.56 //y2=0.755
r264 (  30 68 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.405 //y=1.22 //x2=11.445 //y2=1.375
r265 (  29 67 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.405 //y=0.91 //x2=11.445 //y2=0.755
r266 (  29 30 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=11.405 //y=0.91 //x2=11.405 //y2=1.22
r267 (  28 64 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.68 //y=6.02 //x2=26.68 //y2=4.865
r268 (  27 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.24 //y=6.02 //x2=26.24 //y2=4.865
r269 (  26 45 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.25 //y=6.02 //x2=12.25 //y2=4.865
r270 (  25 73 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.81 //y=6.02 //x2=11.81 //y2=4.865
r271 (  24 52 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=26.097 //y=1.375 //x2=26.205 //y2=1.375
r272 (  24 53 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=26.097 //y=1.375 //x2=25.99 //y2=1.375
r273 (  23 33 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=11.667 //y=1.375 //x2=11.775 //y2=1.375
r274 (  23 34 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=11.667 //y=1.375 //x2=11.56 //y2=1.375
r275 (  21 81 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.27 //y=4.7 //x2=26.27 //y2=4.7
r276 (  19 21 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.96 //x2=26.27 //y2=4.7
r277 (  16 88 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.27 //y=2.08 //x2=26.27 //y2=2.08
r278 (  16 19 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.08 //x2=26.27 //y2=2.96
r279 (  13 70 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=4.7 //x2=11.84 //y2=4.7
r280 (  11 13 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.96 //x2=11.84 //y2=4.7
r281 (  8 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.84 //y=2.08 //x2=11.84 //y2=2.08
r282 (  8 11 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=11.84 //y=2.08 //x2=11.84 //y2=2.96
r283 (  6 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=26.27 //y=2.96 //x2=26.27 //y2=2.96
r284 (  4 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.84 //y=2.96 //x2=11.84 //y2=2.96
r285 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.955 //y=2.96 //x2=11.84 //y2=2.96
r286 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=26.155 //y=2.96 //x2=26.27 //y2=2.96
r287 (  1 2 ) resistor r=13.5496 //w=0.131 //l=14.2 //layer=m1 \
 //thickness=0.36 //x=26.155 //y=2.96 //x2=11.955 //y2=2.96
ends PM_DFFSNRNX1_PCELL\%noxref_8

subckt PM_DFFSNRNX1_PCELL\%noxref_9 ( 1 2 3 4 5 6 16 24 37 38 45 53 59 60 64 \
 66 73 74 75 76 77 78 79 80 81 82 83 87 88 89 94 96 99 100 104 105 106 111 113 \
 116 117 121 122 123 128 130 133 134 136 137 142 146 147 152 156 157 162 165 \
 167 168 169 )
c336 ( 169 0 ) capacitor c=0.023087f //x=17.575 //y=5.02
c337 ( 168 0 ) capacitor c=0.023519f //x=16.695 //y=5.02
c338 ( 167 0 ) capacitor c=0.0224735f //x=15.815 //y=5.02
c339 ( 165 0 ) capacitor c=0.00853354f //x=17.825 //y=0.915
c340 ( 162 0 ) capacitor c=0.0617593f //x=27.38 //y=4.7
c341 ( 157 0 ) capacitor c=0.0273931f //x=27.38 //y=1.915
c342 ( 156 0 ) capacitor c=0.0471168f //x=27.38 //y=2.08
c343 ( 152 0 ) capacitor c=0.0587755f //x=12.95 //y=4.7
c344 ( 147 0 ) capacitor c=0.0273931f //x=12.95 //y=1.915
c345 ( 146 0 ) capacitor c=0.0456313f //x=12.95 //y=2.08
c346 ( 142 0 ) capacitor c=0.058931f //x=8.14 //y=4.7
c347 ( 137 0 ) capacitor c=0.0273931f //x=8.14 //y=1.915
c348 ( 136 0 ) capacitor c=0.0456313f //x=8.14 //y=2.08
c349 ( 134 0 ) capacitor c=0.0432517f //x=27.9 //y=1.26
c350 ( 133 0 ) capacitor c=0.0200379f //x=27.9 //y=0.915
c351 ( 130 0 ) capacitor c=0.0158629f //x=27.745 //y=1.415
c352 ( 128 0 ) capacitor c=0.0157803f //x=27.745 //y=0.76
c353 ( 123 0 ) capacitor c=0.0218028f //x=27.37 //y=1.57
c354 ( 122 0 ) capacitor c=0.0207459f //x=27.37 //y=1.26
c355 ( 121 0 ) capacitor c=0.0194308f //x=27.37 //y=0.915
c356 ( 117 0 ) capacitor c=0.0432517f //x=13.47 //y=1.26
c357 ( 116 0 ) capacitor c=0.0200379f //x=13.47 //y=0.915
c358 ( 113 0 ) capacitor c=0.0148873f //x=13.315 //y=1.415
c359 ( 111 0 ) capacitor c=0.0157803f //x=13.315 //y=0.76
c360 ( 106 0 ) capacitor c=0.0218028f //x=12.94 //y=1.57
c361 ( 105 0 ) capacitor c=0.0207459f //x=12.94 //y=1.26
c362 ( 104 0 ) capacitor c=0.0194308f //x=12.94 //y=0.915
c363 ( 100 0 ) capacitor c=0.0432517f //x=8.66 //y=1.26
c364 ( 99 0 ) capacitor c=0.0200379f //x=8.66 //y=0.915
c365 ( 96 0 ) capacitor c=0.0148873f //x=8.505 //y=1.415
c366 ( 94 0 ) capacitor c=0.0157803f //x=8.505 //y=0.76
c367 ( 89 0 ) capacitor c=0.0218028f //x=8.13 //y=1.57
c368 ( 88 0 ) capacitor c=0.0207459f //x=8.13 //y=1.26
c369 ( 87 0 ) capacitor c=0.0194308f //x=8.13 //y=0.915
c370 ( 83 0 ) capacitor c=0.158794f //x=27.56 //y=6.02
c371 ( 82 0 ) capacitor c=0.110114f //x=27.12 //y=6.02
c372 ( 81 0 ) capacitor c=0.158794f //x=13.13 //y=6.02
c373 ( 80 0 ) capacitor c=0.110114f //x=12.69 //y=6.02
c374 ( 79 0 ) capacitor c=0.158794f //x=8.32 //y=6.02
c375 ( 78 0 ) capacitor c=0.110114f //x=7.88 //y=6.02
c376 ( 74 0 ) capacitor c=0.00125776f //x=17.72 //y=5.155
c377 ( 73 0 ) capacitor c=0.0023095f //x=16.84 //y=5.155
c378 ( 66 0 ) capacitor c=0.0932167f //x=27.38 //y=2.08
c379 ( 64 0 ) capacitor c=0.109929f //x=18.5 //y=3.7
c380 ( 60 0 ) capacitor c=0.00398962f //x=18.1 //y=1.665
c381 ( 59 0 ) capacitor c=0.0137288f //x=18.415 //y=1.665
c382 ( 53 0 ) capacitor c=0.0298716f //x=18.415 //y=5.155
c383 ( 45 0 ) capacitor c=0.0191592f //x=17.635 //y=5.155
c384 ( 38 0 ) capacitor c=0.00332903f //x=16.045 //y=5.155
c385 ( 37 0 ) capacitor c=0.014837f //x=16.755 //y=5.155
c386 ( 24 0 ) capacitor c=0.0833868f //x=12.95 //y=2.08
c387 ( 16 0 ) capacitor c=0.0842881f //x=8.14 //y=2.08
c388 ( 6 0 ) capacitor c=0.00717893f //x=18.615 //y=3.7
c389 ( 5 0 ) capacitor c=0.301821f //x=27.265 //y=3.7
c390 ( 4 0 ) capacitor c=0.00584265f //x=13.065 //y=3.7
c391 ( 3 0 ) capacitor c=0.107948f //x=18.385 //y=3.7
c392 ( 2 0 ) capacitor c=0.0142286f //x=8.255 //y=3.7
c393 ( 1 0 ) capacitor c=0.080604f //x=12.835 //y=3.7
r394 (  156 157 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=27.38 //y=2.08 //x2=27.38 //y2=1.915
r395 (  146 147 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=12.95 //y=2.08 //x2=12.95 //y2=1.915
r396 (  136 137 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=8.14 //y=2.08 //x2=8.14 //y2=1.915
r397 (  134 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.9 //y=1.26 //x2=27.86 //y2=1.415
r398 (  133 163 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.9 //y=0.915 //x2=27.86 //y2=0.76
r399 (  133 134 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.9 //y=0.915 //x2=27.9 //y2=1.26
r400 (  131 160 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.525 //y=1.415 //x2=27.41 //y2=1.415
r401 (  130 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.745 //y=1.415 //x2=27.86 //y2=1.415
r402 (  129 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.525 //y=0.76 //x2=27.41 //y2=0.76
r403 (  128 163 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.745 //y=0.76 //x2=27.86 //y2=0.76
r404 (  128 129 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=27.745 //y=0.76 //x2=27.525 //y2=0.76
r405 (  125 162 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=27.56 //y=4.865 //x2=27.38 //y2=4.7
r406 (  123 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.37 //y=1.57 //x2=27.41 //y2=1.415
r407 (  123 157 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.37 //y=1.57 //x2=27.37 //y2=1.915
r408 (  122 160 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.37 //y=1.26 //x2=27.41 //y2=1.415
r409 (  121 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.37 //y=0.915 //x2=27.41 //y2=0.76
r410 (  121 122 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.37 //y=0.915 //x2=27.37 //y2=1.26
r411 (  118 162 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=27.12 //y=4.865 //x2=27.38 //y2=4.7
r412 (  117 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.47 //y=1.26 //x2=13.43 //y2=1.415
r413 (  116 153 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.47 //y=0.915 //x2=13.43 //y2=0.76
r414 (  116 117 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.47 //y=0.915 //x2=13.47 //y2=1.26
r415 (  114 150 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.095 //y=1.415 //x2=12.98 //y2=1.415
r416 (  113 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.315 //y=1.415 //x2=13.43 //y2=1.415
r417 (  112 149 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.095 //y=0.76 //x2=12.98 //y2=0.76
r418 (  111 153 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.315 //y=0.76 //x2=13.43 //y2=0.76
r419 (  111 112 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=13.315 //y=0.76 //x2=13.095 //y2=0.76
r420 (  108 152 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=13.13 //y=4.865 //x2=12.95 //y2=4.7
r421 (  106 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.94 //y=1.57 //x2=12.98 //y2=1.415
r422 (  106 147 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.94 //y=1.57 //x2=12.94 //y2=1.915
r423 (  105 150 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.94 //y=1.26 //x2=12.98 //y2=1.415
r424 (  104 149 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.94 //y=0.915 //x2=12.98 //y2=0.76
r425 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.94 //y=0.915 //x2=12.94 //y2=1.26
r426 (  101 152 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=12.69 //y=4.865 //x2=12.95 //y2=4.7
r427 (  100 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.66 //y=1.26 //x2=8.62 //y2=1.415
r428 (  99 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.66 //y=0.915 //x2=8.62 //y2=0.76
r429 (  99 100 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.66 //y=0.915 //x2=8.66 //y2=1.26
r430 (  97 140 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.285 //y=1.415 //x2=8.17 //y2=1.415
r431 (  96 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.505 //y=1.415 //x2=8.62 //y2=1.415
r432 (  95 139 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.285 //y=0.76 //x2=8.17 //y2=0.76
r433 (  94 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.505 //y=0.76 //x2=8.62 //y2=0.76
r434 (  94 95 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=8.505 //y=0.76 //x2=8.285 //y2=0.76
r435 (  91 142 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=8.32 //y=4.865 //x2=8.14 //y2=4.7
r436 (  89 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.57 //x2=8.17 //y2=1.415
r437 (  89 137 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.57 //x2=8.13 //y2=1.915
r438 (  88 140 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.26 //x2=8.17 //y2=1.415
r439 (  87 139 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=0.915 //x2=8.17 //y2=0.76
r440 (  87 88 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.13 //y=0.915 //x2=8.13 //y2=1.26
r441 (  84 142 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=7.88 //y=4.865 //x2=8.14 //y2=4.7
r442 (  83 125 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=27.56 //y=6.02 //x2=27.56 //y2=4.865
r443 (  82 118 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=27.12 //y=6.02 //x2=27.12 //y2=4.865
r444 (  81 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.13 //y=6.02 //x2=13.13 //y2=4.865
r445 (  80 101 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=12.69 //y=6.02 //x2=12.69 //y2=4.865
r446 (  79 91 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.32 //y=6.02 //x2=8.32 //y2=4.865
r447 (  78 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.88 //y=6.02 //x2=7.88 //y2=4.865
r448 (  77 130 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=27.635 //y=1.415 //x2=27.745 //y2=1.415
r449 (  77 131 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=27.635 //y=1.415 //x2=27.525 //y2=1.415
r450 (  76 113 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.205 //y=1.415 //x2=13.315 //y2=1.415
r451 (  76 114 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=13.205 //y=1.415 //x2=13.095 //y2=1.415
r452 (  75 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.395 //y=1.415 //x2=8.505 //y2=1.415
r453 (  75 97 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.395 //y=1.415 //x2=8.285 //y2=1.415
r454 (  71 162 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=27.38 //y=4.7 //x2=27.38 //y2=4.7
r455 (  69 71 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=27.38 //y=3.7 //x2=27.38 //y2=4.7
r456 (  66 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=27.38 //y=2.08 //x2=27.38 //y2=2.08
r457 (  66 69 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=27.38 //y=2.08 //x2=27.38 //y2=3.7
r458 (  62 64 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=18.5 //y=5.07 //x2=18.5 //y2=3.7
r459 (  61 64 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=18.5 //y=1.75 //x2=18.5 //y2=3.7
r460 (  59 61 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.415 //y=1.665 //x2=18.5 //y2=1.75
r461 (  59 60 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=18.415 //y=1.665 //x2=18.1 //y2=1.665
r462 (  55 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.015 //y=1.58 //x2=18.1 //y2=1.665
r463 (  55 165 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=18.015 //y=1.58 //x2=18.015 //y2=1.01
r464 (  54 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.805 //y=5.155 //x2=17.72 //y2=5.155
r465 (  53 62 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.415 //y=5.155 //x2=18.5 //y2=5.07
r466 (  53 54 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=18.415 //y=5.155 //x2=17.805 //y2=5.155
r467 (  47 74 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.72 //y=5.24 //x2=17.72 //y2=5.155
r468 (  47 169 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.72 //y=5.24 //x2=17.72 //y2=5.725
r469 (  46 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.925 //y=5.155 //x2=16.84 //y2=5.155
r470 (  45 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.635 //y=5.155 //x2=17.72 //y2=5.155
r471 (  45 46 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=17.635 //y=5.155 //x2=16.925 //y2=5.155
r472 (  39 73 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.84 //y=5.24 //x2=16.84 //y2=5.155
r473 (  39 168 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.84 //y=5.24 //x2=16.84 //y2=5.725
r474 (  37 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.755 //y=5.155 //x2=16.84 //y2=5.155
r475 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=16.755 //y=5.155 //x2=16.045 //y2=5.155
r476 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.96 //y=5.24 //x2=16.045 //y2=5.155
r477 (  31 167 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.96 //y=5.24 //x2=15.96 //y2=5.725
r478 (  29 152 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.95 //y=4.7 //x2=12.95 //y2=4.7
r479 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=12.95 //y=3.7 //x2=12.95 //y2=4.7
r480 (  24 146 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=12.95 //y=2.08 //x2=12.95 //y2=2.08
r481 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=12.95 //y=2.08 //x2=12.95 //y2=3.7
r482 (  21 142 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.14 //y=4.7 //x2=8.14 //y2=4.7
r483 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=8.14 //y=3.7 //x2=8.14 //y2=4.7
r484 (  16 136 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.14 //y=2.08 //x2=8.14 //y2=2.08
r485 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=8.14 //y=2.08 //x2=8.14 //y2=3.7
r486 (  14 69 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=27.38 //y=3.7 //x2=27.38 //y2=3.7
r487 (  12 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.5 //y=3.7 //x2=18.5 //y2=3.7
r488 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.95 //y=3.7 //x2=12.95 //y2=3.7
r489 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.14 //y=3.7 //x2=8.14 //y2=3.7
r490 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.615 //y=3.7 //x2=18.5 //y2=3.7
r491 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=27.265 //y=3.7 //x2=27.38 //y2=3.7
r492 (  5 6 ) resistor r=8.25382 //w=0.131 //l=8.65 //layer=m1 \
 //thickness=0.36 //x=27.265 //y=3.7 //x2=18.615 //y2=3.7
r493 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.065 //y=3.7 //x2=12.95 //y2=3.7
r494 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.385 //y=3.7 //x2=18.5 //y2=3.7
r495 (  3 4 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=18.385 //y=3.7 //x2=13.065 //y2=3.7
r496 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.255 //y=3.7 //x2=8.14 //y2=3.7
r497 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.835 //y=3.7 //x2=12.95 //y2=3.7
r498 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=12.835 //y=3.7 //x2=8.255 //y2=3.7
ends PM_DFFSNRNX1_PCELL\%noxref_9

subckt PM_DFFSNRNX1_PCELL\%noxref_10 ( 2 7 8 9 10 11 12 13 14 16 22 23 24 25 )
c57 ( 25 0 ) capacitor c=0.0598646f //x=1.385 //y=4.79
c58 ( 24 0 ) capacitor c=0.0375015f //x=1.675 //y=4.79
c59 ( 23 0 ) capacitor c=0.0347816f //x=1.34 //y=1.22
c60 ( 22 0 ) capacitor c=0.0187487f //x=1.34 //y=0.875
c61 ( 16 0 ) capacitor c=0.0137055f //x=1.185 //y=1.375
c62 ( 14 0 ) capacitor c=0.0149861f //x=1.185 //y=0.72
c63 ( 13 0 ) capacitor c=0.102158f //x=0.81 //y=1.915
c64 ( 12 0 ) capacitor c=0.0229444f //x=0.81 //y=1.53
c65 ( 11 0 ) capacitor c=0.0234352f //x=0.81 //y=1.22
c66 ( 10 0 ) capacitor c=0.0198724f //x=0.81 //y=0.875
c67 ( 9 0 ) capacitor c=0.110114f //x=1.75 //y=6.02
c68 ( 8 0 ) capacitor c=0.158956f //x=1.31 //y=6.02
c69 ( 2 0 ) capacitor c=0.128033f //x=1.11 //y=2.08
r70 (  24 26 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.75 //y2=4.865
r71 (  24 25 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.385 //y2=4.79
r72 (  23 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=1.22 //x2=1.3 //y2=1.375
r73 (  22 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.3 //y2=0.72
r74 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.34 //y2=1.22
r75 (  19 25 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.385 //y2=4.79
r76 (  19 34 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.11 //y2=4.7
r77 (  17 30 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=1.375 //x2=0.85 //y2=1.375
r78 (  16 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=1.375 //x2=1.3 //y2=1.375
r79 (  15 29 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=0.72 //x2=0.85 //y2=0.72
r80 (  14 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=1.3 //y2=0.72
r81 (  14 15 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=0.965 //y2=0.72
r82 (  13 32 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.915 //x2=1.11 //y2=2.08
r83 (  12 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.85 //y2=1.375
r84 (  12 13 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.81 //y2=1.915
r85 (  11 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.22 //x2=0.85 //y2=1.375
r86 (  10 29 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.85 //y2=0.72
r87 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.81 //y2=1.22
r88 (  9 26 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.75 //y=6.02 //x2=1.75 //y2=4.865
r89 (  8 19 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.31 //y=6.02 //x2=1.31 //y2=4.865
r90 (  7 16 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=1.185 //y2=1.375
r91 (  7 17 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=0.965 //y2=1.375
r92 (  5 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r93 (  2 32 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r94 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=4.7
ends PM_DFFSNRNX1_PCELL\%noxref_10

subckt PM_DFFSNRNX1_PCELL\%noxref_11 ( 1 5 9 13 17 35 )
c46 ( 35 0 ) capacitor c=0.0713324f //x=0.455 //y=0.375
c47 ( 17 0 ) capacitor c=0.0250784f //x=2.445 //y=1.59
c48 ( 13 0 ) capacitor c=0.015523f //x=2.445 //y=0.54
c49 ( 9 0 ) capacitor c=0.00678203f //x=1.56 //y=0.625
c50 ( 5 0 ) capacitor c=0.0236189f //x=1.475 //y=1.59
c51 ( 1 0 ) capacitor c=0.0109947f //x=0.59 //y=1.505
r52 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=1.59 //x2=1.56 //y2=1.63
r53 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=1.59 //x2=2.045 //y2=1.59
r54 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=1.59 //x2=2.53 //y2=1.59
r55 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=1.59 //x2=2.045 //y2=1.59
r56 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=0.54 //x2=1.56 //y2=0.5
r57 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=0.54 //x2=2.045 //y2=0.54
r58 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=0.54 //x2=2.53 //y2=0.54
r59 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=0.54 //x2=2.045 //y2=0.54
r60 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=1.63
r61 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=0.89
r62 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.5
r63 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.89
r64 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.675 //y=1.59 //x2=0.59 //y2=1.63
r65 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.675 //y=1.59 //x2=1.075 //y2=1.59
r66 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.475 //y=1.59 //x2=1.56 //y2=1.63
r67 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.475 //y=1.59 //x2=1.075 //y2=1.59
r68 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.59 //y=1.505 //x2=0.59 //y2=1.63
r69 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.59 //y=1.505 //x2=0.59 //y2=0.89
ends PM_DFFSNRNX1_PCELL\%noxref_11

subckt PM_DFFSNRNX1_PCELL\%noxref_12 ( 1 3 11 15 25 28 29 )
c54 ( 29 0 ) capacitor c=0.0414744f //x=2.965 //y=0.375
c55 ( 28 0 ) capacitor c=0.0046366f //x=1.86 //y=0.91
c56 ( 25 0 ) capacitor c=0.00156479f //x=3.1 //y=0.995
c57 ( 15 0 ) capacitor c=0.00737666f //x=4.07 //y=0.625
c58 ( 11 0 ) capacitor c=0.0144274f //x=3.985 //y=0.54
c59 ( 3 0 ) capacitor c=0.00718386f //x=3.1 //y=0.625
c60 ( 1 0 ) capacitor c=0.0218873f //x=3.015 //y=0.995
r61 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.5
r62 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.89
r63 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.185 //y=0.54 //x2=3.1 //y2=0.5
r64 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.185 //y=0.54 //x2=3.585 //y2=0.54
r65 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.985 //y=0.54 //x2=4.07 //y2=0.5
r66 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.985 //y=0.54 //x2=3.585 //y2=0.54
r67 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=0.995
r68 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=1.23
r69 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.995
r70 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.89
r71 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.5
r72 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.89
r73 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.135 //y=0.995 //x2=2.05 //y2=0.995
r74 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=3.1 //y2=0.995
r75 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=2.135 //y2=0.995
ends PM_DFFSNRNX1_PCELL\%noxref_12

subckt PM_DFFSNRNX1_PCELL\%noxref_13 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0673029f //x=5.265 //y=0.375
c51 ( 17 0 ) capacitor c=0.0178317f //x=7.255 //y=1.59
c52 ( 13 0 ) capacitor c=0.0154936f //x=7.255 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=6.37 //y=0.625
c54 ( 5 0 ) capacitor c=0.0164013f //x=6.285 //y=1.59
c55 ( 1 0 ) capacitor c=0.00696517f //x=5.4 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.455 //y=1.59 //x2=6.37 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.455 //y=1.59 //x2=6.855 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.255 //y=1.59 //x2=7.34 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.255 //y=1.59 //x2=6.855 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.455 //y=0.54 //x2=6.37 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.455 //y=0.54 //x2=6.855 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.255 //y=0.54 //x2=7.34 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.255 //y=0.54 //x2=6.855 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=6.37 //y=1.505 //x2=6.37 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.37 //y=1.505 //x2=6.37 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.37 //y=0.625 //x2=6.37 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.37 //y=0.625 //x2=6.37 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.485 //y=1.59 //x2=5.4 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.485 //y=1.59 //x2=5.885 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.285 //y=1.59 //x2=6.37 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.285 //y=1.59 //x2=5.885 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=5.4 //y=1.505 //x2=5.4 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=5.4 //y=1.505 //x2=5.4 //y2=0.89
ends PM_DFFSNRNX1_PCELL\%noxref_13

subckt PM_DFFSNRNX1_PCELL\%noxref_14 ( 1 3 11 15 25 28 29 )
c54 ( 29 0 ) capacitor c=0.0413887f //x=7.775 //y=0.375
c55 ( 28 0 ) capacitor c=0.0045748f //x=6.67 //y=0.91
c56 ( 25 0 ) capacitor c=0.00156479f //x=7.91 //y=0.995
c57 ( 15 0 ) capacitor c=0.00737666f //x=8.88 //y=0.625
c58 ( 11 0 ) capacitor c=0.0144274f //x=8.795 //y=0.54
c59 ( 3 0 ) capacitor c=0.00718386f //x=7.91 //y=0.625
c60 ( 1 0 ) capacitor c=0.0218888f //x=7.825 //y=0.995
r61 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=8.88 //y=0.625 //x2=8.88 //y2=0.5
r62 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=8.88 //y=0.625 //x2=8.88 //y2=0.89
r63 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.995 //y=0.54 //x2=7.91 //y2=0.5
r64 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.995 //y=0.54 //x2=8.395 //y2=0.54
r65 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.795 //y=0.54 //x2=8.88 //y2=0.5
r66 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.795 //y=0.54 //x2=8.395 //y2=0.54
r67 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.91 //y=1.08 //x2=7.91 //y2=0.995
r68 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=7.91 //y=1.08 //x2=7.91 //y2=1.23
r69 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.91 //x2=7.91 //y2=0.995
r70 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.91 //x2=7.91 //y2=0.89
r71 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.625 //x2=7.91 //y2=0.5
r72 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.625 //x2=7.91 //y2=0.89
r73 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.945 //y=0.995 //x2=6.86 //y2=0.995
r74 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.825 //y=0.995 //x2=7.91 //y2=0.995
r75 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=7.825 //y=0.995 //x2=6.945 //y2=0.995
ends PM_DFFSNRNX1_PCELL\%noxref_14

subckt PM_DFFSNRNX1_PCELL\%noxref_15 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0673029f //x=10.075 //y=0.375
c51 ( 17 0 ) capacitor c=0.0178317f //x=12.065 //y=1.59
c52 ( 13 0 ) capacitor c=0.0154936f //x=12.065 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=11.18 //y=0.625
c54 ( 5 0 ) capacitor c=0.0164013f //x=11.095 //y=1.59
c55 ( 1 0 ) capacitor c=0.00696517f //x=10.21 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.265 //y=1.59 //x2=11.18 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.265 //y=1.59 //x2=11.665 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.065 //y=1.59 //x2=12.15 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.065 //y=1.59 //x2=11.665 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.265 //y=0.54 //x2=11.18 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.265 //y=0.54 //x2=11.665 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.065 //y=0.54 //x2=12.15 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.065 //y=0.54 //x2=11.665 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=11.18 //y=1.505 //x2=11.18 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=11.18 //y=1.505 //x2=11.18 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=11.18 //y=0.625 //x2=11.18 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=11.18 //y=0.625 //x2=11.18 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.295 //y=1.59 //x2=10.21 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.295 //y=1.59 //x2=10.695 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.095 //y=1.59 //x2=11.18 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.095 //y=1.59 //x2=10.695 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=10.21 //y=1.505 //x2=10.21 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=10.21 //y=1.505 //x2=10.21 //y2=0.89
ends PM_DFFSNRNX1_PCELL\%noxref_15

subckt PM_DFFSNRNX1_PCELL\%noxref_16 ( 1 3 11 15 25 28 29 )
c54 ( 29 0 ) capacitor c=0.0414744f //x=12.585 //y=0.375
c55 ( 28 0 ) capacitor c=0.0045748f //x=11.48 //y=0.91
c56 ( 25 0 ) capacitor c=0.00156479f //x=12.72 //y=0.995
c57 ( 15 0 ) capacitor c=0.00737666f //x=13.69 //y=0.625
c58 ( 11 0 ) capacitor c=0.0144274f //x=13.605 //y=0.54
c59 ( 3 0 ) capacitor c=0.00718386f //x=12.72 //y=0.625
c60 ( 1 0 ) capacitor c=0.0218888f //x=12.635 //y=0.995
r61 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=13.69 //y=0.625 //x2=13.69 //y2=0.5
r62 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=13.69 //y=0.625 //x2=13.69 //y2=0.89
r63 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.805 //y=0.54 //x2=12.72 //y2=0.5
r64 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.805 //y=0.54 //x2=13.205 //y2=0.54
r65 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.605 //y=0.54 //x2=13.69 //y2=0.5
r66 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.605 //y=0.54 //x2=13.205 //y2=0.54
r67 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=12.72 //y=1.08 //x2=12.72 //y2=0.995
r68 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=12.72 //y=1.08 //x2=12.72 //y2=1.23
r69 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.91 //x2=12.72 //y2=0.995
r70 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.91 //x2=12.72 //y2=0.89
r71 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.625 //x2=12.72 //y2=0.5
r72 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=12.72 //y=0.625 //x2=12.72 //y2=0.89
r73 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.755 //y=0.995 //x2=11.67 //y2=0.995
r74 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=12.635 //y=0.995 //x2=12.72 //y2=0.995
r75 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=12.635 //y=0.995 //x2=11.755 //y2=0.995
ends PM_DFFSNRNX1_PCELL\%noxref_16

subckt PM_DFFSNRNX1_PCELL\%noxref_17 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0673029f //x=14.885 //y=0.375
c51 ( 17 0 ) capacitor c=0.0178317f //x=16.875 //y=1.59
c52 ( 13 0 ) capacitor c=0.0154936f //x=16.875 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=15.99 //y=0.625
c54 ( 5 0 ) capacitor c=0.0164013f //x=15.905 //y=1.59
c55 ( 1 0 ) capacitor c=0.00696517f //x=15.02 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.075 //y=1.59 //x2=15.99 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.075 //y=1.59 //x2=16.475 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.875 //y=1.59 //x2=16.96 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.875 //y=1.59 //x2=16.475 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.075 //y=0.54 //x2=15.99 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.075 //y=0.54 //x2=16.475 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.875 //y=0.54 //x2=16.96 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.875 //y=0.54 //x2=16.475 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=15.99 //y=1.505 //x2=15.99 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=15.99 //y=1.505 //x2=15.99 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=15.99 //y=0.625 //x2=15.99 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=15.99 //y=0.625 //x2=15.99 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.105 //y=1.59 //x2=15.02 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.105 //y=1.59 //x2=15.505 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.905 //y=1.59 //x2=15.99 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.905 //y=1.59 //x2=15.505 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=15.02 //y=1.505 //x2=15.02 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=15.02 //y=1.505 //x2=15.02 //y2=0.89
ends PM_DFFSNRNX1_PCELL\%noxref_17

subckt PM_DFFSNRNX1_PCELL\%noxref_18 ( 1 3 11 15 25 28 29 )
c55 ( 29 0 ) capacitor c=0.0413887f //x=17.395 //y=0.375
c56 ( 28 0 ) capacitor c=0.0045748f //x=16.29 //y=0.91
c57 ( 25 0 ) capacitor c=0.00156479f //x=17.53 //y=0.995
c58 ( 15 0 ) capacitor c=0.00737666f //x=18.5 //y=0.625
c59 ( 11 0 ) capacitor c=0.0144218f //x=18.415 //y=0.54
c60 ( 3 0 ) capacitor c=0.00718386f //x=17.53 //y=0.625
c61 ( 1 0 ) capacitor c=0.0218888f //x=17.445 //y=0.995
r62 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=18.5 //y=0.625 //x2=18.5 //y2=0.5
r63 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=18.5 //y=0.625 //x2=18.5 //y2=0.89
r64 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.615 //y=0.54 //x2=17.53 //y2=0.5
r65 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.615 //y=0.54 //x2=18.015 //y2=0.54
r66 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.415 //y=0.54 //x2=18.5 //y2=0.5
r67 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.415 //y=0.54 //x2=18.015 //y2=0.54
r68 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.53 //y=1.08 //x2=17.53 //y2=0.995
r69 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=17.53 //y=1.08 //x2=17.53 //y2=1.23
r70 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.91 //x2=17.53 //y2=0.995
r71 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.91 //x2=17.53 //y2=0.89
r72 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.625 //x2=17.53 //y2=0.5
r73 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=17.53 //y=0.625 //x2=17.53 //y2=0.89
r74 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.565 //y=0.995 //x2=16.48 //y2=0.995
r75 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=17.445 //y=0.995 //x2=17.53 //y2=0.995
r76 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=17.445 //y=0.995 //x2=16.565 //y2=0.995
ends PM_DFFSNRNX1_PCELL\%noxref_18

subckt PM_DFFSNRNX1_PCELL\%noxref_19 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0680259f //x=19.695 //y=0.375
c53 ( 17 0 ) capacitor c=0.0180446f //x=21.685 //y=1.59
c54 ( 13 0 ) capacitor c=0.0155283f //x=21.685 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=20.8 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=20.715 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=19.83 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.885 //y=1.59 //x2=20.8 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.885 //y=1.59 //x2=21.285 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.685 //y=1.59 //x2=21.77 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.685 //y=1.59 //x2=21.285 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.885 //y=0.54 //x2=20.8 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.885 //y=0.54 //x2=21.285 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.685 //y=0.54 //x2=21.77 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.685 //y=0.54 //x2=21.285 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=20.8 //y=1.505 //x2=20.8 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=20.8 //y=1.505 //x2=20.8 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=20.8 //y=0.625 //x2=20.8 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=20.8 //y=0.625 //x2=20.8 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.915 //y=1.59 //x2=19.83 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.915 //y=1.59 //x2=20.315 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.715 //y=1.59 //x2=20.8 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.715 //y=1.59 //x2=20.315 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=19.83 //y=1.505 //x2=19.83 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=19.83 //y=1.505 //x2=19.83 //y2=0.89
ends PM_DFFSNRNX1_PCELL\%noxref_19

subckt PM_DFFSNRNX1_PCELL\%noxref_20 ( 2 7 8 9 13 14 15 20 22 25 26 28 29 34 )
c59 ( 34 0 ) capacitor c=0.0599242f //x=22.57 //y=4.7
c60 ( 29 0 ) capacitor c=0.0273931f //x=22.57 //y=1.915
c61 ( 28 0 ) capacitor c=0.0458323f //x=22.57 //y=2.08
c62 ( 26 0 ) capacitor c=0.0432517f //x=23.09 //y=1.26
c63 ( 25 0 ) capacitor c=0.0200379f //x=23.09 //y=0.915
c64 ( 22 0 ) capacitor c=0.0158629f //x=22.935 //y=1.415
c65 ( 20 0 ) capacitor c=0.0157803f //x=22.935 //y=0.76
c66 ( 15 0 ) capacitor c=0.0218028f //x=22.56 //y=1.57
c67 ( 14 0 ) capacitor c=0.0207459f //x=22.56 //y=1.26
c68 ( 13 0 ) capacitor c=0.0194308f //x=22.56 //y=0.915
c69 ( 9 0 ) capacitor c=0.158794f //x=22.75 //y=6.02
c70 ( 8 0 ) capacitor c=0.110114f //x=22.31 //y=6.02
c71 ( 2 0 ) capacitor c=0.0914217f //x=22.57 //y=2.08
r72 (  28 29 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=22.57 //y=2.08 //x2=22.57 //y2=1.915
r73 (  26 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.09 //y=1.26 //x2=23.05 //y2=1.415
r74 (  25 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.09 //y=0.915 //x2=23.05 //y2=0.76
r75 (  25 26 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=23.09 //y=0.915 //x2=23.09 //y2=1.26
r76 (  23 32 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.715 //y=1.415 //x2=22.6 //y2=1.415
r77 (  22 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.935 //y=1.415 //x2=23.05 //y2=1.415
r78 (  21 31 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.715 //y=0.76 //x2=22.6 //y2=0.76
r79 (  20 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=22.935 //y=0.76 //x2=23.05 //y2=0.76
r80 (  20 21 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=22.935 //y=0.76 //x2=22.715 //y2=0.76
r81 (  17 34 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=22.75 //y=4.865 //x2=22.57 //y2=4.7
r82 (  15 32 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.56 //y=1.57 //x2=22.6 //y2=1.415
r83 (  15 29 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.56 //y=1.57 //x2=22.56 //y2=1.915
r84 (  14 32 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.56 //y=1.26 //x2=22.6 //y2=1.415
r85 (  13 31 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.56 //y=0.915 //x2=22.6 //y2=0.76
r86 (  13 14 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.56 //y=0.915 //x2=22.56 //y2=1.26
r87 (  10 34 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=22.31 //y=4.865 //x2=22.57 //y2=4.7
r88 (  9 17 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.75 //y=6.02 //x2=22.75 //y2=4.865
r89 (  8 10 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.31 //y=6.02 //x2=22.31 //y2=4.865
r90 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=22.825 //y=1.415 //x2=22.935 //y2=1.415
r91 (  7 23 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=22.825 //y=1.415 //x2=22.715 //y2=1.415
r92 (  5 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.57 //y=4.7 //x2=22.57 //y2=4.7
r93 (  2 28 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.57 //y=2.08 //x2=22.57 //y2=2.08
r94 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=22.57 //y=2.08 //x2=22.57 //y2=4.7
ends PM_DFFSNRNX1_PCELL\%noxref_20

subckt PM_DFFSNRNX1_PCELL\%noxref_21 ( 7 8 15 23 29 30 32 33 34 35 37 38 39 )
c84 ( 39 0 ) capacitor c=0.023087f //x=22.385 //y=5.02
c85 ( 38 0 ) capacitor c=0.023519f //x=21.505 //y=5.02
c86 ( 37 0 ) capacitor c=0.0224735f //x=20.625 //y=5.02
c87 ( 35 0 ) capacitor c=0.00853354f //x=22.635 //y=0.915
c88 ( 34 0 ) capacitor c=0.00125776f //x=22.53 //y=5.155
c89 ( 33 0 ) capacitor c=0.00243871f //x=21.65 //y=5.155
c90 ( 32 0 ) capacitor c=0.114994f //x=23.31 //y=5.07
c91 ( 30 0 ) capacitor c=0.00463522f //x=22.91 //y=1.665
c92 ( 29 0 ) capacitor c=0.0148737f //x=23.225 //y=1.665
c93 ( 23 0 ) capacitor c=0.0298756f //x=23.225 //y=5.155
c94 ( 15 0 ) capacitor c=0.0191592f //x=22.445 //y=5.155
c95 ( 8 0 ) capacitor c=0.00369455f //x=20.855 //y=5.155
c96 ( 7 0 ) capacitor c=0.0161734f //x=21.565 //y=5.155
r97 (  31 32 ) resistor r=227.251 //w=0.187 //l=3.32 //layer=li \
 //thickness=0.1 //x=23.31 //y=1.75 //x2=23.31 //y2=5.07
r98 (  29 31 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.225 //y=1.665 //x2=23.31 //y2=1.75
r99 (  29 30 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=23.225 //y=1.665 //x2=22.91 //y2=1.665
r100 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=22.825 //y=1.58 //x2=22.91 //y2=1.665
r101 (  25 35 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=22.825 //y=1.58 //x2=22.825 //y2=1.01
r102 (  24 34 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.615 //y=5.155 //x2=22.53 //y2=5.155
r103 (  23 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.225 //y=5.155 //x2=23.31 //y2=5.07
r104 (  23 24 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=23.225 //y=5.155 //x2=22.615 //y2=5.155
r105 (  17 34 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.53 //y=5.24 //x2=22.53 //y2=5.155
r106 (  17 39 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.53 //y=5.24 //x2=22.53 //y2=5.725
r107 (  16 33 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.735 //y=5.155 //x2=21.65 //y2=5.155
r108 (  15 34 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.445 //y=5.155 //x2=22.53 //y2=5.155
r109 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.445 //y=5.155 //x2=21.735 //y2=5.155
r110 (  9 33 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.65 //y=5.24 //x2=21.65 //y2=5.155
r111 (  9 38 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.65 //y=5.24 //x2=21.65 //y2=5.725
r112 (  7 33 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=21.565 //y=5.155 //x2=21.65 //y2=5.155
r113 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=21.565 //y=5.155 //x2=20.855 //y2=5.155
r114 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=20.77 //y=5.24 //x2=20.855 //y2=5.155
r115 (  1 37 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.77 //y=5.24 //x2=20.77 //y2=5.725
ends PM_DFFSNRNX1_PCELL\%noxref_21

subckt PM_DFFSNRNX1_PCELL\%noxref_22 ( 1 3 11 15 25 28 29 )
c54 ( 29 0 ) capacitor c=0.0421963f //x=22.205 //y=0.375
c55 ( 28 0 ) capacitor c=0.00457437f //x=21.1 //y=0.91
c56 ( 25 0 ) capacitor c=0.00156479f //x=22.34 //y=0.995
c57 ( 15 0 ) capacitor c=0.00737666f //x=23.31 //y=0.625
c58 ( 11 0 ) capacitor c=0.014695f //x=23.225 //y=0.54
c59 ( 3 0 ) capacitor c=0.00718386f //x=22.34 //y=0.625
c60 ( 1 0 ) capacitor c=0.0234159f //x=22.255 //y=0.995
r61 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=23.31 //y=0.625 //x2=23.31 //y2=0.5
r62 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=23.31 //y=0.625 //x2=23.31 //y2=0.89
r63 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=22.425 //y=0.54 //x2=22.34 //y2=0.5
r64 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.425 //y=0.54 //x2=22.825 //y2=0.54
r65 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.225 //y=0.54 //x2=23.31 //y2=0.5
r66 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.225 //y=0.54 //x2=22.825 //y2=0.54
r67 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.34 //y=1.08 //x2=22.34 //y2=0.995
r68 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=22.34 //y=1.08 //x2=22.34 //y2=1.23
r69 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.91 //x2=22.34 //y2=0.995
r70 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.91 //x2=22.34 //y2=0.89
r71 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.625 //x2=22.34 //y2=0.5
r72 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=22.34 //y=0.625 //x2=22.34 //y2=0.89
r73 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.375 //y=0.995 //x2=21.29 //y2=0.995
r74 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.255 //y=0.995 //x2=22.34 //y2=0.995
r75 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=22.255 //y=0.995 //x2=21.375 //y2=0.995
ends PM_DFFSNRNX1_PCELL\%noxref_22

subckt PM_DFFSNRNX1_PCELL\%noxref_23 ( 2 7 8 9 10 11 12 13 14 16 22 23 24 25 )
c61 ( 25 0 ) capacitor c=0.0562318f //x=25.435 //y=4.79
c62 ( 24 0 ) capacitor c=0.0305765f //x=25.725 //y=4.79
c63 ( 23 0 ) capacitor c=0.0347816f //x=25.39 //y=1.22
c64 ( 22 0 ) capacitor c=0.0187487f //x=25.39 //y=0.875
c65 ( 16 0 ) capacitor c=0.0137055f //x=25.235 //y=1.375
c66 ( 14 0 ) capacitor c=0.0149861f //x=25.235 //y=0.72
c67 ( 13 0 ) capacitor c=0.0970405f //x=24.86 //y=1.915
c68 ( 12 0 ) capacitor c=0.0229444f //x=24.86 //y=1.53
c69 ( 11 0 ) capacitor c=0.0234352f //x=24.86 //y=1.22
c70 ( 10 0 ) capacitor c=0.0198724f //x=24.86 //y=0.875
c71 ( 9 0 ) capacitor c=0.110114f //x=25.8 //y=6.02
c72 ( 8 0 ) capacitor c=0.158956f //x=25.36 //y=6.02
c73 ( 2 0 ) capacitor c=0.108162f //x=25.16 //y=2.08
r74 (  24 26 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=25.725 //y=4.79 //x2=25.8 //y2=4.865
r75 (  24 25 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=25.725 //y=4.79 //x2=25.435 //y2=4.79
r76 (  23 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.39 //y=1.22 //x2=25.35 //y2=1.375
r77 (  22 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.39 //y=0.875 //x2=25.35 //y2=0.72
r78 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=25.39 //y=0.875 //x2=25.39 //y2=1.22
r79 (  19 25 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=25.36 //y=4.865 //x2=25.435 //y2=4.79
r80 (  19 34 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=25.36 //y=4.865 //x2=25.16 //y2=4.7
r81 (  17 30 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.015 //y=1.375 //x2=24.9 //y2=1.375
r82 (  16 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.235 //y=1.375 //x2=25.35 //y2=1.375
r83 (  15 29 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.015 //y=0.72 //x2=24.9 //y2=0.72
r84 (  14 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.235 //y=0.72 //x2=25.35 //y2=0.72
r85 (  14 15 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=25.235 //y=0.72 //x2=25.015 //y2=0.72
r86 (  13 32 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.915 //x2=25.16 //y2=2.08
r87 (  12 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.53 //x2=24.9 //y2=1.375
r88 (  12 13 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.53 //x2=24.86 //y2=1.915
r89 (  11 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.86 //y=1.22 //x2=24.9 //y2=1.375
r90 (  10 29 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.86 //y=0.875 //x2=24.9 //y2=0.72
r91 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.86 //y=0.875 //x2=24.86 //y2=1.22
r92 (  9 26 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=25.8 //y=6.02 //x2=25.8 //y2=4.865
r93 (  8 19 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=25.36 //y=6.02 //x2=25.36 //y2=4.865
r94 (  7 16 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.125 //y=1.375 //x2=25.235 //y2=1.375
r95 (  7 17 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.125 //y=1.375 //x2=25.015 //y2=1.375
r96 (  5 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=25.16 //y=4.7 //x2=25.16 //y2=4.7
r97 (  2 32 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=25.16 //y=2.08 //x2=25.16 //y2=2.08
r98 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=25.16 //y=2.08 //x2=25.16 //y2=4.7
ends PM_DFFSNRNX1_PCELL\%noxref_23

subckt PM_DFFSNRNX1_PCELL\%noxref_24 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0692867f //x=24.505 //y=0.375
c51 ( 17 0 ) capacitor c=0.0199379f //x=26.495 //y=1.59
c52 ( 13 0 ) capacitor c=0.0156068f //x=26.495 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=25.61 //y=0.625
c54 ( 5 0 ) capacitor c=0.0177503f //x=25.525 //y=1.59
c55 ( 1 0 ) capacitor c=0.0076167f //x=24.64 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.695 //y=1.59 //x2=25.61 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.695 //y=1.59 //x2=26.095 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.495 //y=1.59 //x2=26.58 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.495 //y=1.59 //x2=26.095 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.695 //y=0.54 //x2=25.61 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.695 //y=0.54 //x2=26.095 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.495 //y=0.54 //x2=26.58 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.495 //y=0.54 //x2=26.095 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=25.61 //y=1.505 //x2=25.61 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=25.61 //y=1.505 //x2=25.61 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=25.61 //y=0.625 //x2=25.61 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=25.61 //y=0.625 //x2=25.61 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=24.725 //y=1.59 //x2=24.64 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=24.725 //y=1.59 //x2=25.125 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.525 //y=1.59 //x2=25.61 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.525 //y=1.59 //x2=25.125 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=24.64 //y=1.505 //x2=24.64 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=24.64 //y=1.505 //x2=24.64 //y2=0.89
ends PM_DFFSNRNX1_PCELL\%noxref_24

subckt PM_DFFSNRNX1_PCELL\%noxref_25 ( 7 8 15 23 29 30 32 33 34 35 37 38 39 )
c77 ( 39 0 ) capacitor c=0.023087f //x=27.195 //y=5.02
c78 ( 38 0 ) capacitor c=0.023519f //x=26.315 //y=5.02
c79 ( 37 0 ) capacitor c=0.0224735f //x=25.435 //y=5.02
c80 ( 35 0 ) capacitor c=0.00853354f //x=27.445 //y=0.915
c81 ( 34 0 ) capacitor c=0.00125237f //x=27.34 //y=5.155
c82 ( 33 0 ) capacitor c=0.00243871f //x=26.46 //y=5.155
c83 ( 32 0 ) capacitor c=0.133928f //x=28.12 //y=5.07
c84 ( 30 0 ) capacitor c=0.00777616f //x=27.72 //y=1.665
c85 ( 29 0 ) capacitor c=0.0191287f //x=28.035 //y=1.665
c86 ( 23 0 ) capacitor c=0.0349602f //x=28.035 //y=5.155
c87 ( 15 0 ) capacitor c=0.0191592f //x=27.255 //y=5.155
c88 ( 8 0 ) capacitor c=0.00369455f //x=25.665 //y=5.155
c89 ( 7 0 ) capacitor c=0.0161734f //x=26.375 //y=5.155
r90 (  31 32 ) resistor r=227.251 //w=0.187 //l=3.32 //layer=li \
 //thickness=0.1 //x=28.12 //y=1.75 //x2=28.12 //y2=5.07
r91 (  29 31 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=28.035 //y=1.665 //x2=28.12 //y2=1.75
r92 (  29 30 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=28.035 //y=1.665 //x2=27.72 //y2=1.665
r93 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=27.635 //y=1.58 //x2=27.72 //y2=1.665
r94 (  25 35 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=27.635 //y=1.58 //x2=27.635 //y2=1.01
r95 (  24 34 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.425 //y=5.155 //x2=27.34 //y2=5.155
r96 (  23 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=28.035 //y=5.155 //x2=28.12 //y2=5.07
r97 (  23 24 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li //thickness=0.1 \
 //x=28.035 //y=5.155 //x2=27.425 //y2=5.155
r98 (  17 34 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.34 //y=5.24 //x2=27.34 //y2=5.155
r99 (  17 39 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=27.34 //y=5.24 //x2=27.34 //y2=5.725
r100 (  16 33 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.545 //y=5.155 //x2=26.46 //y2=5.155
r101 (  15 34 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.255 //y=5.155 //x2=27.34 //y2=5.155
r102 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=27.255 //y=5.155 //x2=26.545 //y2=5.155
r103 (  9 33 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.46 //y=5.24 //x2=26.46 //y2=5.155
r104 (  9 38 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.46 //y=5.24 //x2=26.46 //y2=5.725
r105 (  7 33 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=26.375 //y=5.155 //x2=26.46 //y2=5.155
r106 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=26.375 //y=5.155 //x2=25.665 //y2=5.155
r107 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.58 //y=5.24 //x2=25.665 //y2=5.155
r108 (  1 37 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=25.58 //y=5.24 //x2=25.58 //y2=5.725
ends PM_DFFSNRNX1_PCELL\%noxref_25

subckt PM_DFFSNRNX1_PCELL\%noxref_26 ( 1 3 11 15 25 28 29 )
c50 ( 29 0 ) capacitor c=0.0429573f //x=27.015 //y=0.375
c51 ( 28 0 ) capacitor c=0.00461946f //x=25.91 //y=0.91
c52 ( 25 0 ) capacitor c=0.00156479f //x=27.15 //y=0.995
c53 ( 15 0 ) capacitor c=0.00737666f //x=28.12 //y=0.625
c54 ( 11 0 ) capacitor c=0.0150034f //x=28.035 //y=0.54
c55 ( 3 0 ) capacitor c=0.00718386f //x=27.15 //y=0.625
c56 ( 1 0 ) capacitor c=0.024638f //x=27.065 //y=0.995
r57 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=28.12 //y=0.625 //x2=28.12 //y2=0.5
r58 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=28.12 //y=0.625 //x2=28.12 //y2=0.89
r59 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=27.235 //y=0.54 //x2=27.15 //y2=0.5
r60 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=27.235 //y=0.54 //x2=27.635 //y2=0.54
r61 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=28.035 //y=0.54 //x2=28.12 //y2=0.5
r62 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=28.035 //y=0.54 //x2=27.635 //y2=0.54
r63 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.15 //y=1.08 //x2=27.15 //y2=0.995
r64 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=27.15 //y=1.08 //x2=27.15 //y2=1.23
r65 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.91 //x2=27.15 //y2=0.995
r66 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.91 //x2=27.15 //y2=0.89
r67 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.625 //x2=27.15 //y2=0.5
r68 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=27.15 //y=0.625 //x2=27.15 //y2=0.89
r69 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.185 //y=0.995 //x2=26.1 //y2=0.995
r70 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=27.065 //y=0.995 //x2=27.15 //y2=0.995
r71 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=27.065 //y=0.995 //x2=26.185 //y2=0.995
ends PM_DFFSNRNX1_PCELL\%noxref_26

