* SPICE3 file created from XOR2X1.ext - technology: sky130A

.subckt XOR2X1 Y A B VDD GND
X0 GND A xor2X1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X1 GND xor2X1_pcell_0/m1_939_797# xor2X1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X2 VDD A xor2X1_pcell_0/a_761_1330# VDD pshort w=2 l=0.15
X3 Y xor2X1_pcell_0/m1_315_501# xor2X1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X4 Y B xor2X1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X5 Y xor2X1_pcell_0/m1_939_797# xor2X1_pcell_0/a_761_1330# VDD pshort w=2 l=0.15
X6 VDD B xor2X1_pcell_0/a_1427_1330# VDD pshort w=2 l=0.15
X7 Y xor2X1_pcell_0/m1_315_501# xor2X1_pcell_0/a_1427_1330# VDD pshort w=2 l=0.15
X8 xor2X1_pcell_0/m1_315_501# A GND GND nshort w=3 l=0.15
X9 VDD A xor2X1_pcell_0/m1_315_501# VDD pshort w=2 l=0.15
X10 xor2X1_pcell_0/m1_939_797# B xor2X1_pcell_0/li1_M1_contact_2/VSUBS xor2X1_pcell_0/li1_M1_contact_2/VSUBS nshort w=3 l=0.15
X11 VDD B xor2X1_pcell_0/m1_939_797# VDD pshort w=2 l=0.15
C0 xor2X1_pcell_0/m1_939_797# B 2.08fF
C1 VDD xor2X1_pcell_0/li1_M1_contact_2/VSUBS 14.15fF
.ends
