magic
tech sky130A
magscale 1 2
timestamp 1652387157
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 205 871 239 905
rect 353 871 387 905
rect 1019 871 1053 905
rect 1685 871 1719 905
rect 2277 871 2311 905
rect 205 797 239 831
rect 353 797 387 831
rect 1019 797 1053 831
rect 1685 797 1719 831
rect 2277 797 2311 831
rect 205 723 239 757
rect 353 723 387 757
rect 1019 723 1053 757
rect 1685 723 1719 757
rect 2277 723 2311 757
rect 205 649 239 683
rect 353 649 387 683
rect 1019 649 1053 683
rect 1685 649 1719 683
rect 2277 649 2311 683
rect 205 575 239 609
rect 353 575 387 609
rect 1019 575 1053 609
rect 1685 575 1719 609
rect 2277 575 2311 609
rect 205 501 239 535
rect 353 501 387 535
rect 1019 501 1053 535
rect 1685 501 1719 535
rect 2277 501 2311 535
rect 205 427 239 461
rect 353 427 387 461
rect 1019 427 1053 461
rect 1685 427 1719 461
rect 2277 427 2311 461
<< metal1 >>
rect -34 1446 2476 1514
rect -34 -34 2476 34
use aoa4x1_pcell  aoa4x1_pcell_0 pcells
timestamp 1652367678
transform 1 0 0 0 1 0
box -87 -34 2529 1550
<< labels >>
rlabel locali 2277 575 2311 609 1 Y
port 1 nsew signal output
rlabel locali 2277 501 2311 535 1 Y
port 1 nsew signal output
rlabel locali 2277 427 2311 461 1 Y
port 1 nsew signal output
rlabel locali 2277 649 2311 683 1 Y
port 1 nsew signal output
rlabel locali 2277 723 2311 757 1 Y
port 1 nsew signal output
rlabel locali 2277 797 2311 831 1 Y
port 1 nsew signal output
rlabel locali 2277 871 2311 905 1 Y
port 1 nsew signal output
rlabel locali 205 575 239 609 1 A
port 2 nsew signal input
rlabel locali 205 501 239 535 1 A
port 2 nsew signal input
rlabel locali 205 427 239 461 1 A
port 2 nsew signal input
rlabel locali 205 649 239 683 1 A
port 2 nsew signal input
rlabel locali 205 723 239 757 1 A
port 2 nsew signal input
rlabel locali 205 797 239 831 1 A
port 2 nsew signal input
rlabel locali 205 871 239 905 1 A
port 2 nsew signal input
rlabel locali 353 649 387 683 1 B
port 3 nsew signal input
rlabel locali 353 723 387 757 1 B
port 3 nsew signal input
rlabel locali 353 871 387 905 1 B
port 3 nsew signal input
rlabel locali 353 797 387 831 1 B
port 3 nsew signal input
rlabel locali 353 575 387 609 1 B
port 3 nsew signal input
rlabel locali 353 501 387 535 1 B
port 3 nsew signal input
rlabel locali 353 427 387 461 1 B
port 3 nsew signal input
rlabel locali 1019 723 1053 757 1 C
port 4 nsew signal input
rlabel locali 1019 797 1053 831 1 C
port 4 nsew signal input
rlabel locali 1019 871 1053 905 1 C
port 4 nsew signal input
rlabel locali 1019 649 1053 683 1 C
port 4 nsew signal input
rlabel locali 1019 575 1053 609 1 C
port 4 nsew signal input
rlabel locali 1019 501 1053 535 1 C
port 4 nsew signal input
rlabel locali 1019 427 1053 461 1 C
port 4 nsew signal input
rlabel locali 1685 797 1719 831 1 D
port 5 nsew signal input
rlabel locali 1685 723 1719 757 1 D
port 5 nsew signal input
rlabel locali 1685 649 1719 683 1 D
port 5 nsew signal input
rlabel locali 1685 575 1719 609 1 D
port 5 nsew signal input
rlabel locali 1685 501 1719 535 1 D
port 5 nsew signal input
rlabel locali 1685 427 1719 461 1 D
port 5 nsew signal input
rlabel locali 1685 871 1719 905 1 D
port 5 nsew signal input
rlabel metal1 -34 1446 2476 1514 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 -34 -34 2476 34 1 VGND
port 7 nsew ground bidirectional abutment
rlabel nwell 57 1463 91 1497 1 VPB
port 8 nsew power bidirectional 
rlabel pwell 57 -17 91 17 1 VNB
port 9 nsew ground bidirectional 
<< properties >>
string LEFclass CORE
string LEFsite unithd
string FIXED_BBOX 0 0 2442 1480
string LEFsymmetry X Y R90
<< end >>
