magic
tech sky130A
magscale 1 2
timestamp 1670281621
<< nwell >>
rect -87 786 1197 1550
<< pwell >>
rect -34 -34 1144 544
<< nmos >>
rect 168 288 198 349
tri 198 288 214 304 sw
rect 362 296 392 349
tri 392 296 408 312 sw
rect 168 258 274 288
tri 274 258 304 288 sw
rect 362 266 468 296
tri 468 266 498 296 sw
rect 168 157 198 258
tri 198 242 214 258 nw
tri 258 242 274 258 ne
tri 198 157 214 173 sw
tri 258 157 274 173 se
rect 274 157 304 258
rect 362 165 392 266
tri 392 250 408 266 nw
tri 452 250 468 266 ne
tri 392 165 408 181 sw
tri 452 165 468 181 se
rect 468 165 498 266
tri 168 127 198 157 ne
rect 198 127 274 157
tri 274 127 304 157 nw
tri 362 135 392 165 ne
rect 392 135 468 165
tri 468 135 498 165 nw
rect 821 297 851 350
tri 851 297 867 313 sw
rect 821 267 927 297
tri 927 267 957 297 sw
rect 821 166 851 267
tri 851 251 867 267 nw
tri 911 251 927 267 ne
tri 851 166 867 182 sw
tri 911 166 927 182 se
rect 927 166 957 267
tri 821 136 851 166 ne
rect 851 136 927 166
tri 927 136 957 166 nw
<< pmos >>
rect 187 1004 217 1404
rect 275 1004 305 1404
rect 363 1004 393 1404
rect 451 1004 481 1404
rect 830 1004 860 1404
rect 918 1004 948 1404
<< ndiff >>
rect 112 333 168 349
rect 112 299 122 333
rect 156 299 168 333
rect 112 261 168 299
rect 198 333 362 349
rect 198 304 219 333
tri 198 288 214 304 ne
rect 214 299 219 304
rect 253 299 316 333
rect 350 299 362 333
rect 214 288 362 299
rect 392 312 554 349
tri 392 296 408 312 ne
rect 408 296 554 312
rect 112 227 122 261
rect 156 227 168 261
tri 274 258 304 288 ne
rect 304 261 362 288
tri 468 266 498 296 ne
rect 112 193 168 227
rect 112 159 122 193
rect 156 159 168 193
rect 112 127 168 159
tri 198 242 214 258 se
rect 214 242 258 258
tri 258 242 274 258 sw
rect 198 208 274 242
rect 198 174 219 208
rect 253 174 274 208
rect 198 173 274 174
tri 198 157 214 173 ne
rect 214 157 258 173
tri 258 157 274 173 nw
rect 304 227 316 261
rect 350 227 362 261
rect 304 193 362 227
rect 304 159 316 193
rect 350 159 362 193
tri 392 250 408 266 se
rect 408 250 452 266
tri 452 250 468 266 sw
rect 392 217 468 250
rect 392 183 413 217
rect 447 183 468 217
rect 392 181 468 183
tri 392 165 408 181 ne
rect 408 165 452 181
tri 452 165 468 181 nw
rect 498 261 554 296
rect 498 227 510 261
rect 544 227 554 261
rect 498 193 554 227
tri 168 127 198 157 sw
tri 274 127 304 157 se
rect 304 135 362 159
tri 362 135 392 165 sw
tri 468 135 498 165 se
rect 498 159 510 193
rect 544 159 554 193
rect 498 135 554 159
rect 304 127 554 135
rect 112 123 554 127
rect 112 89 122 123
rect 156 89 316 123
rect 350 89 413 123
rect 447 89 510 123
rect 544 89 554 123
rect 112 73 554 89
rect 765 334 821 350
rect 765 300 775 334
rect 809 300 821 334
rect 765 262 821 300
rect 851 334 1011 350
rect 851 313 969 334
tri 851 297 867 313 ne
rect 867 300 969 313
rect 1003 300 1011 334
rect 867 297 1011 300
tri 927 267 957 297 ne
rect 765 228 775 262
rect 809 228 821 262
rect 765 194 821 228
rect 765 160 775 194
rect 809 160 821 194
tri 851 251 867 267 se
rect 867 251 911 267
tri 911 251 927 267 sw
rect 851 218 927 251
rect 851 184 871 218
rect 905 184 927 218
rect 851 182 927 184
tri 851 166 867 182 ne
rect 867 166 911 182
tri 911 166 927 182 nw
rect 957 262 1011 297
rect 957 228 969 262
rect 1003 228 1011 262
rect 957 194 1011 228
rect 765 136 821 160
tri 821 136 851 166 sw
tri 927 136 957 166 se
rect 957 160 969 194
rect 1003 160 1011 194
rect 957 136 1011 160
rect 765 124 1011 136
rect 765 90 775 124
rect 809 90 871 124
rect 905 90 969 124
rect 1003 90 1011 124
rect 765 74 1011 90
<< pdiff >>
rect 131 1366 187 1404
rect 131 1332 141 1366
rect 175 1332 187 1366
rect 131 1298 187 1332
rect 131 1264 141 1298
rect 175 1264 187 1298
rect 131 1230 187 1264
rect 131 1196 141 1230
rect 175 1196 187 1230
rect 131 1162 187 1196
rect 131 1128 141 1162
rect 175 1128 187 1162
rect 131 1093 187 1128
rect 131 1059 141 1093
rect 175 1059 187 1093
rect 131 1004 187 1059
rect 217 1366 275 1404
rect 217 1332 229 1366
rect 263 1332 275 1366
rect 217 1298 275 1332
rect 217 1264 229 1298
rect 263 1264 275 1298
rect 217 1230 275 1264
rect 217 1196 229 1230
rect 263 1196 275 1230
rect 217 1162 275 1196
rect 217 1128 229 1162
rect 263 1128 275 1162
rect 217 1093 275 1128
rect 217 1059 229 1093
rect 263 1059 275 1093
rect 217 1004 275 1059
rect 305 1366 363 1404
rect 305 1332 317 1366
rect 351 1332 363 1366
rect 305 1298 363 1332
rect 305 1264 317 1298
rect 351 1264 363 1298
rect 305 1230 363 1264
rect 305 1196 317 1230
rect 351 1196 363 1230
rect 305 1162 363 1196
rect 305 1128 317 1162
rect 351 1128 363 1162
rect 305 1004 363 1128
rect 393 1366 451 1404
rect 393 1332 405 1366
rect 439 1332 451 1366
rect 393 1298 451 1332
rect 393 1264 405 1298
rect 439 1264 451 1298
rect 393 1230 451 1264
rect 393 1196 405 1230
rect 439 1196 451 1230
rect 393 1162 451 1196
rect 393 1128 405 1162
rect 439 1128 451 1162
rect 393 1093 451 1128
rect 393 1059 405 1093
rect 439 1059 451 1093
rect 393 1004 451 1059
rect 481 1366 535 1404
rect 481 1332 493 1366
rect 527 1332 535 1366
rect 481 1298 535 1332
rect 481 1264 493 1298
rect 527 1264 535 1298
rect 481 1230 535 1264
rect 481 1196 493 1230
rect 527 1196 535 1230
rect 481 1162 535 1196
rect 481 1128 493 1162
rect 527 1128 535 1162
rect 481 1004 535 1128
rect 774 1366 830 1404
rect 774 1332 784 1366
rect 818 1332 830 1366
rect 774 1298 830 1332
rect 774 1264 784 1298
rect 818 1264 830 1298
rect 774 1230 830 1264
rect 774 1196 784 1230
rect 818 1196 830 1230
rect 774 1162 830 1196
rect 774 1128 784 1162
rect 818 1128 830 1162
rect 774 1093 830 1128
rect 774 1059 784 1093
rect 818 1059 830 1093
rect 774 1004 830 1059
rect 860 1366 918 1404
rect 860 1332 872 1366
rect 906 1332 918 1366
rect 860 1298 918 1332
rect 860 1264 872 1298
rect 906 1264 918 1298
rect 860 1230 918 1264
rect 860 1196 872 1230
rect 906 1196 918 1230
rect 860 1162 918 1196
rect 860 1128 872 1162
rect 906 1128 918 1162
rect 860 1093 918 1128
rect 860 1059 872 1093
rect 906 1059 918 1093
rect 860 1004 918 1059
rect 948 1366 1002 1404
rect 948 1332 960 1366
rect 994 1332 1002 1366
rect 948 1298 1002 1332
rect 948 1264 960 1298
rect 994 1264 1002 1298
rect 948 1230 1002 1264
rect 948 1196 960 1230
rect 994 1196 1002 1230
rect 948 1162 1002 1196
rect 948 1128 960 1162
rect 994 1128 1002 1162
rect 948 1093 1002 1128
rect 948 1059 960 1093
rect 994 1059 1002 1093
rect 948 1004 1002 1059
<< ndiffc >>
rect 122 299 156 333
rect 219 299 253 333
rect 316 299 350 333
rect 122 227 156 261
rect 122 159 156 193
rect 219 174 253 208
rect 316 227 350 261
rect 316 159 350 193
rect 413 183 447 217
rect 510 227 544 261
rect 510 159 544 193
rect 122 89 156 123
rect 316 89 350 123
rect 413 89 447 123
rect 510 89 544 123
rect 775 300 809 334
rect 969 300 1003 334
rect 775 228 809 262
rect 775 160 809 194
rect 871 184 905 218
rect 969 228 1003 262
rect 969 160 1003 194
rect 775 90 809 124
rect 871 90 905 124
rect 969 90 1003 124
<< pdiffc >>
rect 141 1332 175 1366
rect 141 1264 175 1298
rect 141 1196 175 1230
rect 141 1128 175 1162
rect 141 1059 175 1093
rect 229 1332 263 1366
rect 229 1264 263 1298
rect 229 1196 263 1230
rect 229 1128 263 1162
rect 229 1059 263 1093
rect 317 1332 351 1366
rect 317 1264 351 1298
rect 317 1196 351 1230
rect 317 1128 351 1162
rect 405 1332 439 1366
rect 405 1264 439 1298
rect 405 1196 439 1230
rect 405 1128 439 1162
rect 405 1059 439 1093
rect 493 1332 527 1366
rect 493 1264 527 1298
rect 493 1196 527 1230
rect 493 1128 527 1162
rect 784 1332 818 1366
rect 784 1264 818 1298
rect 784 1196 818 1230
rect 784 1128 818 1162
rect 784 1059 818 1093
rect 872 1332 906 1366
rect 872 1264 906 1298
rect 872 1196 906 1230
rect 872 1128 906 1162
rect 872 1059 906 1093
rect 960 1332 994 1366
rect 960 1264 994 1298
rect 960 1196 994 1230
rect 960 1128 994 1162
rect 960 1059 994 1093
<< psubdiff >>
rect -34 482 1144 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 632 461 700 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 632 427 649 461
rect 683 427 700 461
rect 1076 461 1144 482
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect 1076 427 1093 461
rect 1127 427 1144 461
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 632 313 700 353
rect 1076 387 1144 427
rect 1076 353 1093 387
rect 1127 353 1144 387
rect 632 279 649 313
rect 683 279 700 313
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect -34 17 34 57
rect 632 57 649 91
rect 683 57 700 91
rect 1076 313 1144 353
rect 1076 279 1093 313
rect 1127 279 1144 313
rect 1076 239 1144 279
rect 1076 205 1093 239
rect 1127 205 1144 239
rect 1076 165 1144 205
rect 1076 131 1093 165
rect 1127 131 1144 165
rect 1076 91 1144 131
rect 632 17 700 57
rect 1076 57 1093 91
rect 1127 57 1144 91
rect 1076 17 1144 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1144 17
rect -34 -34 1144 -17
<< nsubdiff >>
rect -34 1497 1144 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1144 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 632 1423 700 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 1076 1423 1144 1463
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 632 979 700 1019
rect 1076 1389 1093 1423
rect 1127 1389 1144 1423
rect 1076 1349 1144 1389
rect 1076 1315 1093 1349
rect 1127 1315 1144 1349
rect 1076 1275 1144 1315
rect 1076 1241 1093 1275
rect 1127 1241 1144 1275
rect 1076 1201 1144 1241
rect 1076 1167 1093 1201
rect 1127 1167 1144 1201
rect 1076 1127 1144 1167
rect 1076 1093 1093 1127
rect 1127 1093 1144 1127
rect 1076 1053 1144 1093
rect 1076 1019 1093 1053
rect 1127 1019 1144 1053
rect 632 945 649 979
rect 683 945 700 979
rect -34 871 -17 905
rect 17 884 34 905
rect 632 905 700 945
rect 1076 979 1144 1019
rect 1076 945 1093 979
rect 1127 945 1144 979
rect 632 884 649 905
rect 17 871 649 884
rect 683 884 700 905
rect 1076 905 1144 945
rect 1076 884 1093 905
rect 683 871 1093 884
rect 1127 871 1144 905
rect -34 822 1144 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 649 427 683 461
rect 649 353 683 387
rect 1093 427 1127 461
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1093 353 1127 387
rect 649 279 683 313
rect 649 205 683 239
rect 649 131 683 165
rect 649 57 683 91
rect 1093 279 1127 313
rect 1093 205 1127 239
rect 1093 131 1127 165
rect 1093 57 1127 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 649 1389 683 1423
rect 649 1315 683 1349
rect 649 1241 683 1275
rect 649 1167 683 1201
rect 649 1093 683 1127
rect 649 1019 683 1053
rect -17 945 17 979
rect 1093 1389 1127 1423
rect 1093 1315 1127 1349
rect 1093 1241 1127 1275
rect 1093 1167 1127 1201
rect 1093 1093 1127 1127
rect 1093 1019 1127 1053
rect 649 945 683 979
rect -17 871 17 905
rect 1093 945 1127 979
rect 649 871 683 905
rect 1093 871 1127 905
<< poly >>
rect 187 1404 217 1430
rect 275 1404 305 1430
rect 363 1404 393 1430
rect 451 1404 481 1430
rect 830 1404 860 1430
rect 918 1404 948 1430
rect 187 973 217 1004
rect 275 973 305 1004
rect 363 973 393 1004
rect 451 973 481 1004
rect 187 957 305 973
rect 187 943 205 957
rect 195 923 205 943
rect 239 943 305 957
rect 349 957 481 973
rect 239 923 249 943
rect 195 907 249 923
rect 349 923 359 957
rect 393 943 481 957
rect 830 973 860 1004
rect 918 973 948 1004
rect 393 923 403 943
rect 349 907 403 923
rect 787 957 948 973
rect 787 923 797 957
rect 831 943 948 957
rect 831 923 841 943
rect 787 907 841 923
rect 195 433 249 449
rect 195 413 205 433
rect 168 399 205 413
rect 239 399 249 433
rect 168 383 249 399
rect 343 433 397 449
rect 343 399 353 433
rect 387 399 397 433
rect 343 383 397 399
rect 168 349 198 383
rect 362 349 392 383
rect 787 434 841 450
rect 787 400 797 434
rect 831 413 841 434
rect 831 400 851 413
rect 787 384 851 400
rect 821 350 851 384
<< polycont >>
rect 205 923 239 957
rect 359 923 393 957
rect 797 923 831 957
rect 205 399 239 433
rect 353 399 387 433
rect 797 400 831 434
<< locali >>
rect -34 1497 1144 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1144 1497
rect -34 1446 1144 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 141 1366 175 1446
rect 141 1298 175 1332
rect 141 1230 175 1264
rect 141 1162 175 1196
rect 141 1093 175 1128
rect 141 1027 175 1059
rect 229 1366 263 1404
rect 229 1298 263 1332
rect 229 1230 263 1264
rect 229 1162 263 1196
rect 229 1093 263 1128
rect 317 1366 351 1446
rect 317 1298 351 1332
rect 317 1230 351 1264
rect 317 1162 351 1196
rect 317 1111 351 1128
rect 405 1366 439 1404
rect 405 1298 439 1332
rect 405 1230 439 1264
rect 405 1162 439 1196
rect 229 1057 263 1059
rect 405 1093 439 1128
rect 493 1366 527 1446
rect 493 1298 527 1332
rect 493 1230 527 1264
rect 493 1162 527 1196
rect 493 1111 527 1128
rect 632 1423 700 1446
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 405 1057 439 1059
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 229 1023 535 1057
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect 359 957 393 973
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 923
rect 205 383 239 399
rect 353 923 359 942
rect 353 907 393 923
rect 353 433 387 907
rect 353 383 387 399
rect 501 683 535 1023
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect 784 1366 818 1446
rect 784 1298 818 1332
rect 784 1230 818 1264
rect 784 1162 818 1196
rect 784 1093 818 1128
rect 784 1037 818 1059
rect 872 1366 906 1404
rect 872 1298 906 1332
rect 872 1230 906 1264
rect 872 1162 906 1196
rect 872 1093 906 1128
rect 632 979 700 1019
rect 632 945 649 979
rect 683 945 700 979
rect 632 905 700 945
rect 632 871 649 905
rect 683 871 700 905
rect 632 822 700 871
rect 797 957 831 973
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 122 333 156 349
rect 316 333 350 349
rect 501 348 535 649
rect 797 683 831 923
rect 872 933 906 1059
rect 960 1366 994 1446
rect 960 1298 994 1332
rect 960 1230 994 1264
rect 960 1162 994 1196
rect 960 1093 994 1128
rect 960 1037 994 1059
rect 1076 1423 1144 1446
rect 1076 1389 1093 1423
rect 1127 1389 1144 1423
rect 1076 1349 1144 1389
rect 1076 1315 1093 1349
rect 1127 1315 1144 1349
rect 1076 1275 1144 1315
rect 1076 1241 1093 1275
rect 1127 1241 1144 1275
rect 1076 1201 1144 1241
rect 1076 1167 1093 1201
rect 1127 1167 1144 1201
rect 1076 1127 1144 1167
rect 1076 1093 1093 1127
rect 1127 1093 1144 1127
rect 1076 1053 1144 1093
rect 1076 1019 1093 1053
rect 1127 1019 1144 1053
rect 1076 979 1144 1019
rect 1076 945 1093 979
rect 1127 945 1144 979
rect 872 899 979 933
rect 156 299 219 333
rect 253 299 316 333
rect 122 261 156 299
rect 122 193 156 227
rect 316 261 350 299
rect 122 123 156 159
rect 122 73 156 89
rect 219 208 253 224
rect -34 34 34 57
rect 219 34 253 174
rect 316 193 350 227
rect 413 314 535 348
rect 632 461 700 544
rect 632 427 649 461
rect 683 427 700 461
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect 797 434 831 649
rect 945 433 979 899
rect 1076 905 1144 945
rect 1076 871 1093 905
rect 1127 871 1144 905
rect 1076 822 1144 871
rect 797 384 831 400
rect 871 399 979 433
rect 1076 461 1144 544
rect 1076 427 1093 461
rect 1127 427 1144 461
rect 413 217 447 314
rect 632 313 700 353
rect 632 279 649 313
rect 683 279 700 313
rect 413 167 447 183
rect 510 261 544 277
rect 510 193 544 227
rect 316 123 350 159
rect 510 123 544 159
rect 350 89 413 123
rect 447 89 510 123
rect 316 73 350 89
rect 510 73 544 89
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect 632 57 649 91
rect 683 57 700 91
rect 632 34 700 57
rect 775 334 809 350
rect 775 262 809 300
rect 775 194 809 228
rect 871 218 905 399
rect 1076 387 1144 427
rect 1076 353 1093 387
rect 1127 353 1144 387
rect 871 168 905 184
rect 969 334 1003 350
rect 969 262 1003 300
rect 969 194 1003 228
rect 775 124 809 160
rect 969 124 1003 160
rect 809 90 871 124
rect 905 90 969 124
rect 775 34 809 90
rect 872 34 906 90
rect 969 34 1003 90
rect 1076 313 1144 353
rect 1076 279 1093 313
rect 1127 279 1144 313
rect 1076 239 1144 279
rect 1076 205 1093 239
rect 1127 205 1144 239
rect 1076 165 1144 205
rect 1076 131 1093 165
rect 1127 131 1144 165
rect 1076 91 1144 131
rect 1076 57 1093 91
rect 1127 57 1144 91
rect 1076 34 1144 57
rect -34 17 1144 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1144 17
rect -34 -34 1144 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 501 649 535 683
rect 797 649 831 683
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
<< metal1 >>
rect -34 1497 1144 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1144 1497
rect -34 1446 1144 1463
rect 495 683 541 689
rect 791 683 837 689
rect 489 649 501 683
rect 535 649 797 683
rect 831 649 843 683
rect 495 643 541 649
rect 791 643 837 649
rect -34 17 1144 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1144 17
rect -34 -34 1144 -17
<< labels >>
rlabel locali 945 575 979 609 1 Y
port 1 nsew signal output
rlabel locali 945 501 979 535 1 Y
port 1 nsew signal output
rlabel locali 945 427 979 461 1 Y
port 1 nsew signal output
rlabel locali 945 649 979 683 1 Y
port 1 nsew signal output
rlabel locali 945 723 979 757 1 Y
port 1 nsew signal output
rlabel locali 945 797 979 831 1 Y
port 1 nsew signal output
rlabel locali 945 871 979 905 1 Y
port 1 nsew signal output
rlabel locali 205 427 239 461 1 A
port 2 nsew signal input
rlabel locali 205 501 239 535 1 A
port 2 nsew signal input
rlabel locali 205 575 239 609 1 A
port 2 nsew signal input
rlabel locali 205 649 239 683 1 A
port 2 nsew signal input
rlabel locali 205 723 239 757 1 A
port 2 nsew signal input
rlabel locali 205 797 239 831 1 A
port 2 nsew signal input
rlabel locali 205 871 239 905 1 A
port 2 nsew signal input
rlabel locali 353 871 387 905 1 B
port 3 nsew signal input
rlabel locali 353 797 387 831 1 B
port 3 nsew signal input
rlabel locali 353 723 387 757 1 B
port 3 nsew signal input
rlabel locali 353 649 387 683 1 B
port 3 nsew signal input
rlabel locali 353 575 387 609 1 B
port 3 nsew signal input
rlabel locali 353 501 387 535 1 B
port 3 nsew signal input
rlabel locali 353 427 387 461 1 B
port 3 nsew signal input
rlabel metal1 -34 1446 1144 1514 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 -34 -34 1144 34 1 GND
port 5 nsew ground bidirectional abutment
<< end >>
