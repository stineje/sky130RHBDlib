// File: TMRDFFRNQNX1.spi.pex
// Created: Tue Oct 15 15:52:03 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_TMRDFFRNQNX1\%GND ( 1 147 151 154 159 169 177 187 195 203 209 219 \
 225 235 241 247 255 265 273 283 291 299 307 317 325 335 343 351 357 367 373 \
 383 389 395 403 413 421 431 439 447 455 463 469 475 488 492 494 496 499 502 \
 505 507 509 511 513 515 517 520 523 526 528 530 532 534 537 539 540 541 542 \
 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 )
c991 ( 559 0 ) capacitor c=0.0215012f //x=85.35 //y=0.865
c992 ( 558 0 ) capacitor c=0.0215012f //x=82.02 //y=0.865
c993 ( 557 0 ) capacitor c=0.0207524f //x=78.69 //y=0.865
c994 ( 556 0 ) capacitor c=0.0207873f //x=75.36 //y=0.865
c995 ( 555 0 ) capacitor c=0.0225954f //x=70.445 //y=0.875
c996 ( 554 0 ) capacitor c=0.0226075f //x=65.635 //y=0.875
c997 ( 553 0 ) capacitor c=0.0207407f //x=62.41 //y=0.865
c998 ( 552 0 ) capacitor c=0.0225954f //x=57.495 //y=0.875
c999 ( 551 0 ) capacitor c=0.0226075f //x=52.685 //y=0.875
c1000 ( 550 0 ) capacitor c=0.0207407f //x=49.46 //y=0.865
c1001 ( 549 0 ) capacitor c=0.0225954f //x=44.545 //y=0.875
c1002 ( 548 0 ) capacitor c=0.0226075f //x=39.735 //y=0.875
c1003 ( 547 0 ) capacitor c=0.0207407f //x=36.51 //y=0.865
c1004 ( 546 0 ) capacitor c=0.0225954f //x=31.595 //y=0.875
c1005 ( 545 0 ) capacitor c=0.0226075f //x=26.785 //y=0.875
c1006 ( 544 0 ) capacitor c=0.0207407f //x=23.56 //y=0.865
c1007 ( 543 0 ) capacitor c=0.0225954f //x=18.645 //y=0.875
c1008 ( 542 0 ) capacitor c=0.0226075f //x=13.835 //y=0.875
c1009 ( 541 0 ) capacitor c=0.0207407f //x=10.61 //y=0.865
c1010 ( 540 0 ) capacitor c=0.0226571f //x=5.695 //y=0.875
c1011 ( 539 0 ) capacitor c=0.022675f //x=0.885 //y=0.875
c1012 ( 538 0 ) capacitor c=0.00440095f //x=85.54 //y=0
c1013 ( 537 0 ) capacitor c=0.101477f //x=84.36 //y=0
c1014 ( 536 0 ) capacitor c=0.00440095f //x=82.14 //y=0
c1015 ( 534 0 ) capacitor c=0.116475f //x=81.03 //y=0
c1016 ( 533 0 ) capacitor c=0.00440095f //x=78.88 //y=0
c1017 ( 532 0 ) capacitor c=0.104074f //x=77.7 //y=0
c1018 ( 531 0 ) capacitor c=0.00440095f //x=75.55 //y=0
c1019 ( 530 0 ) capacitor c=0.109295f //x=74.37 //y=0
c1020 ( 529 0 ) capacitor c=0.00440144f //x=70.635 //y=0
c1021 ( 528 0 ) capacitor c=0.106903f //x=69.56 //y=0
c1022 ( 527 0 ) capacitor c=0.00440144f //x=65.825 //y=0
c1023 ( 526 0 ) capacitor c=0.10413f //x=64.75 //y=0
c1024 ( 525 0 ) capacitor c=0.00440095f //x=62.53 //y=0
c1025 ( 523 0 ) capacitor c=0.10799f //x=61.42 //y=0
c1026 ( 522 0 ) capacitor c=0.00440144f //x=57.72 //y=0
c1027 ( 520 0 ) capacitor c=0.107403f //x=56.61 //y=0
c1028 ( 519 0 ) capacitor c=0.00440144f //x=52.91 //y=0
c1029 ( 517 0 ) capacitor c=0.104579f //x=51.8 //y=0
c1030 ( 516 0 ) capacitor c=0.00440095f //x=49.65 //y=0
c1031 ( 515 0 ) capacitor c=0.108685f //x=48.47 //y=0
c1032 ( 514 0 ) capacitor c=0.00440144f //x=44.735 //y=0
c1033 ( 513 0 ) capacitor c=0.107329f //x=43.66 //y=0
c1034 ( 512 0 ) capacitor c=0.00440144f //x=39.925 //y=0
c1035 ( 511 0 ) capacitor c=0.104555f //x=38.85 //y=0
c1036 ( 510 0 ) capacitor c=0.00440095f //x=36.7 //y=0
c1037 ( 509 0 ) capacitor c=0.108565f //x=35.52 //y=0
c1038 ( 508 0 ) capacitor c=0.00440144f //x=31.785 //y=0
c1039 ( 507 0 ) capacitor c=0.107403f //x=30.71 //y=0
c1040 ( 506 0 ) capacitor c=0.00440144f //x=26.975 //y=0
c1041 ( 505 0 ) capacitor c=0.104579f //x=25.9 //y=0
c1042 ( 504 0 ) capacitor c=0.00440095f //x=23.68 //y=0
c1043 ( 502 0 ) capacitor c=0.108685f //x=22.57 //y=0
c1044 ( 501 0 ) capacitor c=0.00440144f //x=18.87 //y=0
c1045 ( 499 0 ) capacitor c=0.107329f //x=17.76 //y=0
c1046 ( 498 0 ) capacitor c=0.00440144f //x=14.06 //y=0
c1047 ( 496 0 ) capacitor c=0.104555f //x=12.95 //y=0
c1048 ( 495 0 ) capacitor c=0.00440095f //x=10.8 //y=0
c1049 ( 494 0 ) capacitor c=0.108565f //x=9.62 //y=0
c1050 ( 493 0 ) capacitor c=0.00440144f //x=5.885 //y=0
c1051 ( 492 0 ) capacitor c=0.108357f //x=4.81 //y=0
c1052 ( 491 0 ) capacitor c=0.00440144f //x=1.075 //y=0
c1053 ( 488 0 ) capacitor c=0.258637f //x=86.95 //y=0
c1054 ( 475 0 ) capacitor c=0.0389876f //x=85.455 //y=0
c1055 ( 469 0 ) capacitor c=0.0716428f //x=84.19 //y=0
c1056 ( 463 0 ) capacitor c=0.0388276f //x=82.125 //y=0
c1057 ( 455 0 ) capacitor c=0.0717666f //x=80.86 //y=0
c1058 ( 447 0 ) capacitor c=0.0391432f //x=78.795 //y=0
c1059 ( 439 0 ) capacitor c=0.0718766f //x=77.53 //y=0
c1060 ( 431 0 ) capacitor c=0.0389171f //x=75.465 //y=0
c1061 ( 421 0 ) capacitor c=0.133607f //x=74.2 //y=0
c1062 ( 413 0 ) capacitor c=0.0339325f //x=70.55 //y=0
c1063 ( 403 0 ) capacitor c=0.133561f //x=69.39 //y=0
c1064 ( 395 0 ) capacitor c=0.0339325f //x=65.74 //y=0
c1065 ( 389 0 ) capacitor c=0.0718026f //x=64.58 //y=0
c1066 ( 383 0 ) capacitor c=0.0388888f //x=62.515 //y=0
c1067 ( 373 0 ) capacitor c=0.133561f //x=61.25 //y=0
c1068 ( 367 0 ) capacitor c=0.0339325f //x=57.6 //y=0
c1069 ( 357 0 ) capacitor c=0.133362f //x=56.44 //y=0
c1070 ( 351 0 ) capacitor c=0.0339325f //x=52.79 //y=0
c1071 ( 343 0 ) capacitor c=0.0718026f //x=51.63 //y=0
c1072 ( 335 0 ) capacitor c=0.0388888f //x=49.565 //y=0
c1073 ( 325 0 ) capacitor c=0.133362f //x=48.3 //y=0
c1074 ( 317 0 ) capacitor c=0.0339325f //x=44.65 //y=0
c1075 ( 307 0 ) capacitor c=0.133561f //x=43.49 //y=0
c1076 ( 299 0 ) capacitor c=0.0339325f //x=39.84 //y=0
c1077 ( 291 0 ) capacitor c=0.0718026f //x=38.68 //y=0
c1078 ( 283 0 ) capacitor c=0.0388888f //x=36.615 //y=0
c1079 ( 273 0 ) capacitor c=0.133561f //x=35.35 //y=0
c1080 ( 265 0 ) capacitor c=0.0339325f //x=31.7 //y=0
c1081 ( 255 0 ) capacitor c=0.133362f //x=30.54 //y=0
c1082 ( 247 0 ) capacitor c=0.0339325f //x=26.89 //y=0
c1083 ( 241 0 ) capacitor c=0.0718026f //x=25.73 //y=0
c1084 ( 235 0 ) capacitor c=0.0388888f //x=23.665 //y=0
c1085 ( 225 0 ) capacitor c=0.133362f //x=22.4 //y=0
c1086 ( 219 0 ) capacitor c=0.0339325f //x=18.75 //y=0
c1087 ( 209 0 ) capacitor c=0.133561f //x=17.59 //y=0
c1088 ( 203 0 ) capacitor c=0.0339325f //x=13.94 //y=0
c1089 ( 195 0 ) capacitor c=0.0718026f //x=12.78 //y=0
c1090 ( 187 0 ) capacitor c=0.0388888f //x=10.715 //y=0
c1091 ( 177 0 ) capacitor c=0.133526f //x=9.45 //y=0
c1092 ( 169 0 ) capacitor c=0.0339738f //x=5.8 //y=0
c1093 ( 159 0 ) capacitor c=0.131745f //x=4.64 //y=0
c1094 ( 154 0 ) capacitor c=0.178285f //x=0.74 //y=0
c1095 ( 151 0 ) capacitor c=0.0367385f //x=0.99 //y=0
c1096 ( 147 0 ) capacitor c=2.63764f //x=86.95 //y=0
r1097 (  486 488 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=85.84 //y=0 //x2=86.95 //y2=0
r1098 (  484 538 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=85.625 //y=0 //x2=85.54 //y2=0
r1099 (  484 486 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=85.625 //y=0 //x2=85.84 //y2=0
r1100 (  479 538 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=85.54 //y=0.17 //x2=85.54 //y2=0
r1101 (  479 559 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=85.54 //y=0.17 //x2=85.54 //y2=0.955
r1102 (  476 537 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=84.53 //y=0 //x2=84.36 //y2=0
r1103 (  476 478 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=84.53 //y=0 //x2=84.73 //y2=0
r1104 (  475 538 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=85.455 //y=0 //x2=85.54 //y2=0
r1105 (  475 478 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=85.455 //y=0 //x2=84.73 //y2=0
r1106 (  470 536 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.295 //y=0 //x2=82.21 //y2=0
r1107 (  470 472 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=82.295 //y=0 //x2=83.25 //y2=0
r1108 (  469 537 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=84.19 //y=0 //x2=84.36 //y2=0
r1109 (  469 472 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=84.19 //y=0 //x2=83.25 //y2=0
r1110 (  465 536 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=82.21 //y=0.17 //x2=82.21 //y2=0
r1111 (  465 558 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=82.21 //y=0.17 //x2=82.21 //y2=0.955
r1112 (  464 534 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=81.2 //y=0 //x2=81.03 //y2=0
r1113 (  463 536 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.125 //y=0 //x2=82.21 //y2=0
r1114 (  463 464 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=82.125 //y=0 //x2=81.2 //y2=0
r1115 (  458 460 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=79.55 //y=0 //x2=80.66 //y2=0
r1116 (  456 533 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.965 //y=0 //x2=78.88 //y2=0
r1117 (  456 458 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=78.965 //y=0 //x2=79.55 //y2=0
r1118 (  455 534 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=80.86 //y=0 //x2=81.03 //y2=0
r1119 (  455 460 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=80.86 //y=0 //x2=80.66 //y2=0
r1120 (  451 533 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=78.88 //y=0.17 //x2=78.88 //y2=0
r1121 (  451 557 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=78.88 //y=0.17 //x2=78.88 //y2=0.955
r1122 (  448 532 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=77.87 //y=0 //x2=77.7 //y2=0
r1123 (  448 450 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=77.87 //y=0 //x2=78.44 //y2=0
r1124 (  447 533 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.795 //y=0 //x2=78.88 //y2=0
r1125 (  447 450 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=78.795 //y=0 //x2=78.44 //y2=0
r1126 (  442 444 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=75.85 //y=0 //x2=76.96 //y2=0
r1127 (  440 531 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.635 //y=0 //x2=75.55 //y2=0
r1128 (  440 442 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=75.635 //y=0 //x2=75.85 //y2=0
r1129 (  439 532 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=77.53 //y=0 //x2=77.7 //y2=0
r1130 (  439 444 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=77.53 //y=0 //x2=76.96 //y2=0
r1131 (  435 531 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=75.55 //y=0.17 //x2=75.55 //y2=0
r1132 (  435 556 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=75.55 //y=0.17 //x2=75.55 //y2=0.955
r1133 (  432 530 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=74.54 //y=0 //x2=74.37 //y2=0
r1134 (  432 434 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=74.54 //y=0 //x2=74.74 //y2=0
r1135 (  431 531 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.465 //y=0 //x2=75.55 //y2=0
r1136 (  431 434 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=75.465 //y=0 //x2=74.74 //y2=0
r1137 (  426 428 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=72.15 //y=0 //x2=73.26 //y2=0
r1138 (  424 426 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=71.04 //y=0 //x2=72.15 //y2=0
r1139 (  422 529 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.72 //y=0 //x2=70.635 //y2=0
r1140 (  422 424 ) resistor r=11.4734 //w=0.357 //l=0.32 //layer=li \
 //thickness=0.1 //x=70.72 //y=0 //x2=71.04 //y2=0
r1141 (  421 530 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=74.2 //y=0 //x2=74.37 //y2=0
r1142 (  421 428 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=74.2 //y=0 //x2=73.26 //y2=0
r1143 (  417 529 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=70.635 //y=0.17 //x2=70.635 //y2=0
r1144 (  417 555 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=70.635 //y=0.17 //x2=70.635 //y2=0.965
r1145 (  414 528 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=69.73 //y=0 //x2=69.56 //y2=0
r1146 (  414 416 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=69.73 //y=0 //x2=69.93 //y2=0
r1147 (  413 529 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.55 //y=0 //x2=70.635 //y2=0
r1148 (  413 416 ) resistor r=22.2297 //w=0.357 //l=0.62 //layer=li \
 //thickness=0.1 //x=70.55 //y=0 //x2=69.93 //y2=0
r1149 (  408 410 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=67.34 //y=0 //x2=68.45 //y2=0
r1150 (  406 408 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=66.23 //y=0 //x2=67.34 //y2=0
r1151 (  404 527 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.91 //y=0 //x2=65.825 //y2=0
r1152 (  404 406 ) resistor r=11.4734 //w=0.357 //l=0.32 //layer=li \
 //thickness=0.1 //x=65.91 //y=0 //x2=66.23 //y2=0
r1153 (  403 528 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=69.39 //y=0 //x2=69.56 //y2=0
r1154 (  403 410 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=69.39 //y=0 //x2=68.45 //y2=0
r1155 (  399 527 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=65.825 //y=0.17 //x2=65.825 //y2=0
r1156 (  399 554 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=65.825 //y=0.17 //x2=65.825 //y2=0.965
r1157 (  396 526 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.92 //y=0 //x2=64.75 //y2=0
r1158 (  396 398 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=64.92 //y=0 //x2=65.12 //y2=0
r1159 (  395 527 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.74 //y=0 //x2=65.825 //y2=0
r1160 (  395 398 ) resistor r=22.2297 //w=0.357 //l=0.62 //layer=li \
 //thickness=0.1 //x=65.74 //y=0 //x2=65.12 //y2=0
r1161 (  390 525 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.685 //y=0 //x2=62.6 //y2=0
r1162 (  390 392 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=62.685 //y=0 //x2=63.64 //y2=0
r1163 (  389 526 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.58 //y=0 //x2=64.75 //y2=0
r1164 (  389 392 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=64.58 //y=0 //x2=63.64 //y2=0
r1165 (  385 525 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.6 //y=0.17 //x2=62.6 //y2=0
r1166 (  385 553 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=62.6 //y=0.17 //x2=62.6 //y2=0.955
r1167 (  384 523 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.59 //y=0 //x2=61.42 //y2=0
r1168 (  383 525 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.515 //y=0 //x2=62.6 //y2=0
r1169 (  383 384 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=62.515 //y=0 //x2=61.59 //y2=0
r1170 (  378 380 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=59.94 //y=0 //x2=61.05 //y2=0
r1171 (  376 378 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=58.83 //y=0 //x2=59.94 //y2=0
r1172 (  374 522 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=57.77 //y=0 //x2=57.685 //y2=0
r1173 (  374 376 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=57.77 //y=0 //x2=58.83 //y2=0
r1174 (  373 523 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.25 //y=0 //x2=61.42 //y2=0
r1175 (  373 380 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=61.25 //y=0 //x2=61.05 //y2=0
r1176 (  369 522 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.685 //y=0.17 //x2=57.685 //y2=0
r1177 (  369 552 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=57.685 //y=0.17 //x2=57.685 //y2=0.965
r1178 (  368 520 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=56.78 //y=0 //x2=56.61 //y2=0
r1179 (  367 522 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=57.6 //y=0 //x2=57.685 //y2=0
r1180 (  367 368 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=57.6 //y=0 //x2=56.78 //y2=0
r1181 (  362 364 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=55.13 //y=0 //x2=56.24 //y2=0
r1182 (  360 362 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=54.02 //y=0 //x2=55.13 //y2=0
r1183 (  358 519 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=52.96 //y=0 //x2=52.875 //y2=0
r1184 (  358 360 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=52.96 //y=0 //x2=54.02 //y2=0
r1185 (  357 520 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=56.44 //y=0 //x2=56.61 //y2=0
r1186 (  357 364 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=56.44 //y=0 //x2=56.24 //y2=0
r1187 (  353 519 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=52.875 //y=0.17 //x2=52.875 //y2=0
r1188 (  353 551 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=52.875 //y=0.17 //x2=52.875 //y2=0.965
r1189 (  352 517 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=51.97 //y=0 //x2=51.8 //y2=0
r1190 (  351 519 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=52.79 //y=0 //x2=52.875 //y2=0
r1191 (  351 352 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=52.79 //y=0 //x2=51.97 //y2=0
r1192 (  346 348 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=50.32 //y=0 //x2=51.43 //y2=0
r1193 (  344 516 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.735 //y=0 //x2=49.65 //y2=0
r1194 (  344 346 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=49.735 //y=0 //x2=50.32 //y2=0
r1195 (  343 517 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=51.63 //y=0 //x2=51.8 //y2=0
r1196 (  343 348 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=51.63 //y=0 //x2=51.43 //y2=0
r1197 (  339 516 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.65 //y=0.17 //x2=49.65 //y2=0
r1198 (  339 550 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=49.65 //y=0.17 //x2=49.65 //y2=0.955
r1199 (  336 515 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.64 //y=0 //x2=48.47 //y2=0
r1200 (  336 338 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=48.64 //y=0 //x2=49.21 //y2=0
r1201 (  335 516 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.565 //y=0 //x2=49.65 //y2=0
r1202 (  335 338 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=49.565 //y=0 //x2=49.21 //y2=0
r1203 (  330 332 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=46.62 //y=0 //x2=47.73 //y2=0
r1204 (  328 330 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=45.51 //y=0 //x2=46.62 //y2=0
r1205 (  326 514 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.82 //y=0 //x2=44.735 //y2=0
r1206 (  326 328 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=44.82 //y=0 //x2=45.51 //y2=0
r1207 (  325 515 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.3 //y=0 //x2=48.47 //y2=0
r1208 (  325 332 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=48.3 //y=0 //x2=47.73 //y2=0
r1209 (  321 514 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=44.735 //y=0.17 //x2=44.735 //y2=0
r1210 (  321 549 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=44.735 //y=0.17 //x2=44.735 //y2=0.965
r1211 (  318 513 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.83 //y=0 //x2=43.66 //y2=0
r1212 (  318 320 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.83 //y=0 //x2=44.4 //y2=0
r1213 (  317 514 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.65 //y=0 //x2=44.735 //y2=0
r1214 (  317 320 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=44.65 //y=0 //x2=44.4 //y2=0
r1215 (  312 314 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=41.81 //y=0 //x2=42.92 //y2=0
r1216 (  310 312 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=40.7 //y=0 //x2=41.81 //y2=0
r1217 (  308 512 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.01 //y=0 //x2=39.925 //y2=0
r1218 (  308 310 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=40.01 //y=0 //x2=40.7 //y2=0
r1219 (  307 513 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.49 //y=0 //x2=43.66 //y2=0
r1220 (  307 314 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.49 //y=0 //x2=42.92 //y2=0
r1221 (  303 512 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.925 //y=0.17 //x2=39.925 //y2=0
r1222 (  303 548 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=39.925 //y=0.17 //x2=39.925 //y2=0.965
r1223 (  300 511 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.02 //y=0 //x2=38.85 //y2=0
r1224 (  300 302 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=39.02 //y=0 //x2=39.59 //y2=0
r1225 (  299 512 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.84 //y=0 //x2=39.925 //y2=0
r1226 (  299 302 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=39.84 //y=0 //x2=39.59 //y2=0
r1227 (  294 296 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=37 //y=0 //x2=38.11 //y2=0
r1228 (  292 510 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.785 //y=0 //x2=36.7 //y2=0
r1229 (  292 294 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=36.785 //y=0 //x2=37 //y2=0
r1230 (  291 511 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.68 //y=0 //x2=38.85 //y2=0
r1231 (  291 296 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=38.68 //y=0 //x2=38.11 //y2=0
r1232 (  287 510 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.7 //y=0.17 //x2=36.7 //y2=0
r1233 (  287 547 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=36.7 //y=0.17 //x2=36.7 //y2=0.955
r1234 (  284 509 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=35.69 //y=0 //x2=35.52 //y2=0
r1235 (  284 286 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=35.69 //y=0 //x2=35.89 //y2=0
r1236 (  283 510 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.615 //y=0 //x2=36.7 //y2=0
r1237 (  283 286 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=36.615 //y=0 //x2=35.89 //y2=0
r1238 (  278 280 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=33.3 //y=0 //x2=34.41 //y2=0
r1239 (  276 278 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=32.19 //y=0 //x2=33.3 //y2=0
r1240 (  274 508 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.87 //y=0 //x2=31.785 //y2=0
r1241 (  274 276 ) resistor r=11.4734 //w=0.357 //l=0.32 //layer=li \
 //thickness=0.1 //x=31.87 //y=0 //x2=32.19 //y2=0
r1242 (  273 509 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=35.35 //y=0 //x2=35.52 //y2=0
r1243 (  273 280 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=35.35 //y=0 //x2=34.41 //y2=0
r1244 (  269 508 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=31.785 //y=0.17 //x2=31.785 //y2=0
r1245 (  269 546 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=31.785 //y=0.17 //x2=31.785 //y2=0.965
r1246 (  266 507 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.88 //y=0 //x2=30.71 //y2=0
r1247 (  266 268 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=30.88 //y=0 //x2=31.08 //y2=0
r1248 (  265 508 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.7 //y=0 //x2=31.785 //y2=0
r1249 (  265 268 ) resistor r=22.2297 //w=0.357 //l=0.62 //layer=li \
 //thickness=0.1 //x=31.7 //y=0 //x2=31.08 //y2=0
r1250 (  260 262 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=28.49 //y=0 //x2=29.6 //y2=0
r1251 (  258 260 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=27.38 //y=0 //x2=28.49 //y2=0
r1252 (  256 506 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.06 //y=0 //x2=26.975 //y2=0
r1253 (  256 258 ) resistor r=11.4734 //w=0.357 //l=0.32 //layer=li \
 //thickness=0.1 //x=27.06 //y=0 //x2=27.38 //y2=0
r1254 (  255 507 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.54 //y=0 //x2=30.71 //y2=0
r1255 (  255 262 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=30.54 //y=0 //x2=29.6 //y2=0
r1256 (  251 506 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.975 //y=0.17 //x2=26.975 //y2=0
r1257 (  251 545 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=26.975 //y=0.17 //x2=26.975 //y2=0.965
r1258 (  248 505 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.07 //y=0 //x2=25.9 //y2=0
r1259 (  248 250 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=26.07 //y=0 //x2=26.27 //y2=0
r1260 (  247 506 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.89 //y=0 //x2=26.975 //y2=0
r1261 (  247 250 ) resistor r=22.2297 //w=0.357 //l=0.62 //layer=li \
 //thickness=0.1 //x=26.89 //y=0 //x2=26.27 //y2=0
r1262 (  242 504 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.835 //y=0 //x2=23.75 //y2=0
r1263 (  242 244 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=23.835 //y=0 //x2=24.79 //y2=0
r1264 (  241 505 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.73 //y=0 //x2=25.9 //y2=0
r1265 (  241 244 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=25.73 //y=0 //x2=24.79 //y2=0
r1266 (  237 504 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.75 //y=0.17 //x2=23.75 //y2=0
r1267 (  237 544 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=23.75 //y=0.17 //x2=23.75 //y2=0.955
r1268 (  236 502 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.74 //y=0 //x2=22.57 //y2=0
r1269 (  235 504 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.665 //y=0 //x2=23.75 //y2=0
r1270 (  235 236 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=23.665 //y=0 //x2=22.74 //y2=0
r1271 (  230 232 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=21.09 //y=0 //x2=22.2 //y2=0
r1272 (  228 230 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=19.98 //y=0 //x2=21.09 //y2=0
r1273 (  226 501 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.92 //y=0 //x2=18.835 //y2=0
r1274 (  226 228 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=18.92 //y=0 //x2=19.98 //y2=0
r1275 (  225 502 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.4 //y=0 //x2=22.57 //y2=0
r1276 (  225 232 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=22.4 //y=0 //x2=22.2 //y2=0
r1277 (  221 501 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.835 //y=0.17 //x2=18.835 //y2=0
r1278 (  221 543 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=18.835 //y=0.17 //x2=18.835 //y2=0.965
r1279 (  220 499 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.93 //y=0 //x2=17.76 //y2=0
r1280 (  219 501 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.75 //y=0 //x2=18.835 //y2=0
r1281 (  219 220 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=18.75 //y=0 //x2=17.93 //y2=0
r1282 (  214 216 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=16.28 //y=0 //x2=17.39 //y2=0
r1283 (  212 214 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=15.17 //y=0 //x2=16.28 //y2=0
r1284 (  210 498 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.11 //y=0 //x2=14.025 //y2=0
r1285 (  210 212 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=14.11 //y=0 //x2=15.17 //y2=0
r1286 (  209 499 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.59 //y=0 //x2=17.76 //y2=0
r1287 (  209 216 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=17.59 //y=0 //x2=17.39 //y2=0
r1288 (  205 498 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.025 //y=0.17 //x2=14.025 //y2=0
r1289 (  205 542 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=14.025 //y=0.17 //x2=14.025 //y2=0.965
r1290 (  204 496 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.12 //y=0 //x2=12.95 //y2=0
r1291 (  203 498 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.94 //y=0 //x2=14.025 //y2=0
r1292 (  203 204 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=13.94 //y=0 //x2=13.12 //y2=0
r1293 (  198 200 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=11.47 //y=0 //x2=12.58 //y2=0
r1294 (  196 495 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.885 //y=0 //x2=10.8 //y2=0
r1295 (  196 198 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=10.885 //y=0 //x2=11.47 //y2=0
r1296 (  195 496 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.78 //y=0 //x2=12.95 //y2=0
r1297 (  195 200 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.78 //y=0 //x2=12.58 //y2=0
r1298 (  191 495 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.8 //y=0.17 //x2=10.8 //y2=0
r1299 (  191 541 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=10.8 //y=0.17 //x2=10.8 //y2=0.955
r1300 (  188 494 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.79 //y=0 //x2=9.62 //y2=0
r1301 (  188 190 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.79 //y=0 //x2=10.36 //y2=0
r1302 (  187 495 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.715 //y=0 //x2=10.8 //y2=0
r1303 (  187 190 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=10.715 //y=0 //x2=10.36 //y2=0
r1304 (  182 184 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=7.77 //y=0 //x2=8.88 //y2=0
r1305 (  180 182 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r1306 (  178 493 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.97 //y=0 //x2=5.885 //y2=0
r1307 (  178 180 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=5.97 //y=0 //x2=6.66 //y2=0
r1308 (  177 494 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.45 //y=0 //x2=9.62 //y2=0
r1309 (  177 184 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.45 //y=0 //x2=8.88 //y2=0
r1310 (  173 493 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.885 //y=0.17 //x2=5.885 //y2=0
r1311 (  173 540 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=5.885 //y=0.17 //x2=5.885 //y2=0.965
r1312 (  170 492 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=4.81 //y2=0
r1313 (  170 172 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=5.55 //y2=0
r1314 (  169 493 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.8 //y=0 //x2=5.885 //y2=0
r1315 (  169 172 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=5.8 //y=0 //x2=5.55 //y2=0
r1316 (  164 166 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=0 //x2=4.07 //y2=0
r1317 (  162 164 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r1318 (  160 491 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.075 //y2=0
r1319 (  160 162 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.85 //y2=0
r1320 (  159 492 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.81 //y2=0
r1321 (  159 166 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.07 //y2=0
r1322 (  155 491 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0
r1323 (  155 539 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0.965
r1324 (  151 491 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=1.075 //y2=0
r1325 (  151 154 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=0.74 //y2=0
r1326 (  147 488 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=86.95 //y=0 //x2=86.95 //y2=0
r1327 (  145 486 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=85.84 //y=0 //x2=85.84 //y2=0
r1328 (  145 147 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=85.84 //y=0 //x2=86.95 //y2=0
r1329 (  143 478 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=84.73 //y=0 //x2=84.73 //y2=0
r1330 (  143 145 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=84.73 //y=0 //x2=85.84 //y2=0
r1331 (  141 472 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=83.25 //y=0 //x2=83.25 //y2=0
r1332 (  141 143 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=83.25 //y=0 //x2=84.73 //y2=0
r1333 (  139 536 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=82.14 //y=0 //x2=82.14 //y2=0
r1334 (  139 141 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=82.14 //y=0 //x2=83.25 //y2=0
r1335 (  137 460 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=80.66 //y=0 //x2=80.66 //y2=0
r1336 (  137 139 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=80.66 //y=0 //x2=82.14 //y2=0
r1337 (  135 458 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=79.55 //y=0 //x2=79.55 //y2=0
r1338 (  135 137 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=79.55 //y=0 //x2=80.66 //y2=0
r1339 (  133 450 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=78.44 //y=0 //x2=78.44 //y2=0
r1340 (  133 135 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=78.44 //y=0 //x2=79.55 //y2=0
r1341 (  131 444 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=76.96 //y=0 //x2=76.96 //y2=0
r1342 (  131 133 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=76.96 //y=0 //x2=78.44 //y2=0
r1343 (  129 442 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=75.85 //y=0 //x2=75.85 //y2=0
r1344 (  129 131 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=75.85 //y=0 //x2=76.96 //y2=0
r1345 (  127 434 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=74.74 //y=0 //x2=74.74 //y2=0
r1346 (  127 129 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=74.74 //y=0 //x2=75.85 //y2=0
r1347 (  125 428 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=73.26 //y=0 //x2=73.26 //y2=0
r1348 (  125 127 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=73.26 //y=0 //x2=74.74 //y2=0
r1349 (  123 426 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=72.15 //y=0 //x2=72.15 //y2=0
r1350 (  123 125 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=72.15 //y=0 //x2=73.26 //y2=0
r1351 (  121 424 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=71.04 //y=0 //x2=71.04 //y2=0
r1352 (  121 123 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=71.04 //y=0 //x2=72.15 //y2=0
r1353 (  119 416 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=69.93 //y=0 //x2=69.93 //y2=0
r1354 (  119 121 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=69.93 //y=0 //x2=71.04 //y2=0
r1355 (  117 410 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=68.45 //y=0 //x2=68.45 //y2=0
r1356 (  117 119 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=68.45 //y=0 //x2=69.93 //y2=0
r1357 (  115 408 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=67.34 //y=0 //x2=67.34 //y2=0
r1358 (  115 117 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=67.34 //y=0 //x2=68.45 //y2=0
r1359 (  113 406 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=66.23 //y=0 //x2=66.23 //y2=0
r1360 (  113 115 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=66.23 //y=0 //x2=67.34 //y2=0
r1361 (  111 398 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=65.12 //y=0 //x2=65.12 //y2=0
r1362 (  111 113 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=65.12 //y=0 //x2=66.23 //y2=0
r1363 (  109 392 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=63.64 //y=0 //x2=63.64 //y2=0
r1364 (  109 111 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=63.64 //y=0 //x2=65.12 //y2=0
r1365 (  107 525 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=62.53 //y=0 //x2=62.53 //y2=0
r1366 (  107 109 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=62.53 //y=0 //x2=63.64 //y2=0
r1367 (  105 380 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=61.05 //y=0 //x2=61.05 //y2=0
r1368 (  105 107 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=61.05 //y=0 //x2=62.53 //y2=0
r1369 (  103 378 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=59.94 //y=0 //x2=59.94 //y2=0
r1370 (  103 105 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=59.94 //y=0 //x2=61.05 //y2=0
r1371 (  101 376 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=58.83 //y=0 //x2=58.83 //y2=0
r1372 (  101 103 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=58.83 //y=0 //x2=59.94 //y2=0
r1373 (  99 522 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=57.72 //y=0 //x2=57.72 //y2=0
r1374 (  99 101 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=57.72 //y=0 //x2=58.83 //y2=0
r1375 (  97 364 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=56.24 //y=0 //x2=56.24 //y2=0
r1376 (  97 99 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=56.24 //y=0 //x2=57.72 //y2=0
r1377 (  95 362 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=55.13 //y=0 //x2=55.13 //y2=0
r1378 (  95 97 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=55.13 //y=0 //x2=56.24 //y2=0
r1379 (  93 360 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=54.02 //y=0 //x2=54.02 //y2=0
r1380 (  93 95 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=54.02 //y=0 //x2=55.13 //y2=0
r1381 (  91 519 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=52.91 //y=0 //x2=52.91 //y2=0
r1382 (  91 93 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=52.91 //y=0 //x2=54.02 //y2=0
r1383 (  89 348 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=51.43 //y=0 //x2=51.43 //y2=0
r1384 (  89 91 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=51.43 //y=0 //x2=52.91 //y2=0
r1385 (  87 346 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=50.32 //y=0 //x2=50.32 //y2=0
r1386 (  87 89 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=50.32 //y=0 //x2=51.43 //y2=0
r1387 (  85 338 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=49.21 //y=0 //x2=49.21 //y2=0
r1388 (  85 87 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=49.21 //y=0 //x2=50.32 //y2=0
r1389 (  83 332 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=47.73 //y=0 //x2=47.73 //y2=0
r1390 (  83 85 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=47.73 //y=0 //x2=49.21 //y2=0
r1391 (  81 330 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=46.62 //y=0 //x2=46.62 //y2=0
r1392 (  81 83 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=46.62 //y=0 //x2=47.73 //y2=0
r1393 (  79 328 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=45.51 //y=0 //x2=45.51 //y2=0
r1394 (  79 81 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=45.51 //y=0 //x2=46.62 //y2=0
r1395 (  77 320 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=44.4 //y=0 //x2=44.4 //y2=0
r1396 (  77 79 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=44.4 //y=0 //x2=45.51 //y2=0
r1397 (  74 314 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=42.92 //y=0 //x2=42.92 //y2=0
r1398 (  72 312 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=41.81 //y=0 //x2=41.81 //y2=0
r1399 (  72 74 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=41.81 //y=0 //x2=42.92 //y2=0
r1400 (  70 310 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=40.7 //y=0 //x2=40.7 //y2=0
r1401 (  70 72 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=40.7 //y=0 //x2=41.81 //y2=0
r1402 (  68 302 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=39.59 //y=0 //x2=39.59 //y2=0
r1403 (  68 70 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=39.59 //y=0 //x2=40.7 //y2=0
r1404 (  66 296 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=38.11 //y=0 //x2=38.11 //y2=0
r1405 (  66 68 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=38.11 //y=0 //x2=39.59 //y2=0
r1406 (  64 294 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37 //y=0 //x2=37 //y2=0
r1407 (  64 66 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=37 //y=0 //x2=38.11 //y2=0
r1408 (  62 286 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.89 //y=0 //x2=35.89 //y2=0
r1409 (  62 64 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=35.89 //y=0 //x2=37 //y2=0
r1410 (  60 280 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.41 //y=0 //x2=34.41 //y2=0
r1411 (  60 62 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=34.41 //y=0 //x2=35.89 //y2=0
r1412 (  58 278 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=33.3 //y=0 //x2=33.3 //y2=0
r1413 (  58 60 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=33.3 //y=0 //x2=34.41 //y2=0
r1414 (  56 276 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.19 //y=0 //x2=32.19 //y2=0
r1415 (  56 58 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=32.19 //y=0 //x2=33.3 //y2=0
r1416 (  54 268 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.08 //y=0 //x2=31.08 //y2=0
r1417 (  54 56 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.08 //y=0 //x2=32.19 //y2=0
r1418 (  52 262 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=29.6 //y=0 //x2=29.6 //y2=0
r1419 (  52 54 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=29.6 //y=0 //x2=31.08 //y2=0
r1420 (  50 260 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.49 //y=0 //x2=28.49 //y2=0
r1421 (  50 52 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=28.49 //y=0 //x2=29.6 //y2=0
r1422 (  48 258 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.38 //y=0 //x2=27.38 //y2=0
r1423 (  48 50 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=27.38 //y=0 //x2=28.49 //y2=0
r1424 (  46 250 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=26.27 //y=0 //x2=26.27 //y2=0
r1425 (  46 48 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=26.27 //y=0 //x2=27.38 //y2=0
r1426 (  44 244 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=0 //x2=24.79 //y2=0
r1427 (  44 46 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=0 //x2=26.27 //y2=0
r1428 (  42 504 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=0 //x2=23.68 //y2=0
r1429 (  42 44 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=23.68 //y=0 //x2=24.79 //y2=0
r1430 (  40 232 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.2 //y=0 //x2=22.2 //y2=0
r1431 (  40 42 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=22.2 //y=0 //x2=23.68 //y2=0
r1432 (  38 230 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=0 //x2=21.09 //y2=0
r1433 (  38 40 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=0 //x2=22.2 //y2=0
r1434 (  36 228 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=0 //x2=19.98 //y2=0
r1435 (  36 38 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=0 //x2=21.09 //y2=0
r1436 (  34 501 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.87 //y=0 //x2=18.87 //y2=0
r1437 (  34 36 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=18.87 //y=0 //x2=19.98 //y2=0
r1438 (  32 216 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=0 //x2=17.39 //y2=0
r1439 (  32 34 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=0 //x2=18.87 //y2=0
r1440 (  30 214 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=0 //x2=16.28 //y2=0
r1441 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=0 //x2=17.39 //y2=0
r1442 (  28 212 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=0 //x2=15.17 //y2=0
r1443 (  28 30 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=0 //x2=16.28 //y2=0
r1444 (  26 498 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=0 //x2=14.06 //y2=0
r1445 (  26 28 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=0 //x2=15.17 //y2=0
r1446 (  24 200 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=0 //x2=12.58 //y2=0
r1447 (  24 26 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=0 //x2=14.06 //y2=0
r1448 (  22 198 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=0 //x2=11.47 //y2=0
r1449 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=0 //x2=12.58 //y2=0
r1450 (  20 190 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r1451 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=0 //x2=11.47 //y2=0
r1452 (  18 184 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.88 //y=0 //x2=8.88 //y2=0
r1453 (  18 20 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.88 //y=0 //x2=10.36 //y2=0
r1454 (  16 182 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r1455 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=8.88 //y2=0
r1456 (  14 180 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r1457 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r1458 (  12 172 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r1459 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r1460 (  10 166 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r1461 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=0 //x2=5.55 //y2=0
r1462 (  8 164 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r1463 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.07 //y2=0
r1464 (  6 162 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r1465 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r1466 (  3 154 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r1467 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r1468 (  1 77 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=43.845 //y=0 //x2=44.4 //y2=0
r1469 (  1 74 ) resistor r=0.384136 //w=0.301 //l=0.925 //layer=m1 \
 //thickness=0.36 //x=43.845 //y=0 //x2=42.92 //y2=0
ends PM_TMRDFFRNQNX1\%GND

subckt PM_TMRDFFRNQNX1\%VDD ( 1 147 154 161 171 179 189 195 205 215 223 233 \
 239 247 255 265 271 279 287 297 307 313 321 329 339 349 355 363 373 383 387 \
 397 407 417 425 429 439 449 459 467 471 481 491 499 503 513 523 531 541 547 \
 557 567 575 585 591 599 607 617 623 631 639 649 659 665 673 681 691 701 707 \
 715 725 735 739 749 759 769 777 781 791 801 811 819 823 833 843 855 863 871 \
 881 887 902 909 914 919 925 931 935 941 947 952 957 962 967 973 979 983 989 \
 995 1000 1005 1006 1007 1008 1009 1010 1011 1012 1013 1014 1015 1016 1017 \
 1018 1019 1020 1021 1022 1023 1024 1025 1026 1027 1028 1029 1030 1031 1032 \
 1033 1034 1035 1036 1037 1038 1039 1040 1041 1042 1043 1044 1045 1046 1047 \
 1048 1049 1050 1051 1052 1053 1054 1055 1056 1057 1058 1059 1060 1061 1062 \
 1063 1064 1065 1066 1067 1068 1069 1070 1071 1072 1073 1074 1075 )
c1101 ( 1075 0 ) capacitor c=0.0476806f //x=80.105 //y=5.025
c1102 ( 1074 0 ) capacitor c=0.0241714f //x=79.225 //y=5.025
c1103 ( 1073 0 ) capacitor c=0.0467094f //x=78.355 //y=5.025
c1104 ( 1072 0 ) capacitor c=0.0382077f //x=76.775 //y=5.02
c1105 ( 1071 0 ) capacitor c=0.0240874f //x=75.895 //y=5.02
c1106 ( 1070 0 ) capacitor c=0.0495444f //x=75.025 //y=5.02
c1107 ( 1069 0 ) capacitor c=0.0453059f //x=73.145 //y=5.02
c1108 ( 1068 0 ) capacitor c=0.02424f //x=72.265 //y=5.02
c1109 ( 1067 0 ) capacitor c=0.02424f //x=71.385 //y=5.02
c1110 ( 1066 0 ) capacitor c=0.0531793f //x=70.515 //y=5.02
c1111 ( 1065 0 ) capacitor c=0.0453059f //x=68.335 //y=5.02
c1112 ( 1064 0 ) capacitor c=0.02424f //x=67.455 //y=5.02
c1113 ( 1063 0 ) capacitor c=0.024152f //x=66.575 //y=5.02
c1114 ( 1062 0 ) capacitor c=0.0531894f //x=65.705 //y=5.02
c1115 ( 1061 0 ) capacitor c=0.0380679f //x=63.825 //y=5.02
c1116 ( 1060 0 ) capacitor c=0.024008f //x=62.945 //y=5.02
c1117 ( 1059 0 ) capacitor c=0.049209f //x=62.075 //y=5.02
c1118 ( 1058 0 ) capacitor c=0.0452179f //x=60.195 //y=5.02
c1119 ( 1057 0 ) capacitor c=0.024152f //x=59.315 //y=5.02
c1120 ( 1056 0 ) capacitor c=0.024152f //x=58.435 //y=5.02
c1121 ( 1055 0 ) capacitor c=0.053132f //x=57.565 //y=5.02
c1122 ( 1054 0 ) capacitor c=0.0452179f //x=55.385 //y=5.02
c1123 ( 1053 0 ) capacitor c=0.024152f //x=54.505 //y=5.02
c1124 ( 1052 0 ) capacitor c=0.024152f //x=53.625 //y=5.02
c1125 ( 1051 0 ) capacitor c=0.0531894f //x=52.755 //y=5.02
c1126 ( 1050 0 ) capacitor c=0.0380679f //x=50.875 //y=5.02
c1127 ( 1049 0 ) capacitor c=0.024008f //x=49.995 //y=5.02
c1128 ( 1048 0 ) capacitor c=0.049209f //x=49.125 //y=5.02
c1129 ( 1047 0 ) capacitor c=0.0452179f //x=47.245 //y=5.02
c1130 ( 1046 0 ) capacitor c=0.024152f //x=46.365 //y=5.02
c1131 ( 1045 0 ) capacitor c=0.024152f //x=45.485 //y=5.02
c1132 ( 1044 0 ) capacitor c=0.053132f //x=44.615 //y=5.02
c1133 ( 1043 0 ) capacitor c=0.0452179f //x=42.435 //y=5.02
c1134 ( 1042 0 ) capacitor c=0.024152f //x=41.555 //y=5.02
c1135 ( 1041 0 ) capacitor c=0.024152f //x=40.675 //y=5.02
c1136 ( 1040 0 ) capacitor c=0.0531894f //x=39.805 //y=5.02
c1137 ( 1039 0 ) capacitor c=0.0380679f //x=37.925 //y=5.02
c1138 ( 1038 0 ) capacitor c=0.024008f //x=37.045 //y=5.02
c1139 ( 1037 0 ) capacitor c=0.049209f //x=36.175 //y=5.02
c1140 ( 1036 0 ) capacitor c=0.0452179f //x=34.295 //y=5.02
c1141 ( 1035 0 ) capacitor c=0.024152f //x=33.415 //y=5.02
c1142 ( 1034 0 ) capacitor c=0.024152f //x=32.535 //y=5.02
c1143 ( 1033 0 ) capacitor c=0.053132f //x=31.665 //y=5.02
c1144 ( 1032 0 ) capacitor c=0.0452179f //x=29.485 //y=5.02
c1145 ( 1031 0 ) capacitor c=0.024152f //x=28.605 //y=5.02
c1146 ( 1030 0 ) capacitor c=0.024152f //x=27.725 //y=5.02
c1147 ( 1029 0 ) capacitor c=0.0531894f //x=26.855 //y=5.02
c1148 ( 1028 0 ) capacitor c=0.0380679f //x=24.975 //y=5.02
c1149 ( 1027 0 ) capacitor c=0.024008f //x=24.095 //y=5.02
c1150 ( 1026 0 ) capacitor c=0.049209f //x=23.225 //y=5.02
c1151 ( 1025 0 ) capacitor c=0.0452179f //x=21.345 //y=5.02
c1152 ( 1024 0 ) capacitor c=0.024152f //x=20.465 //y=5.02
c1153 ( 1023 0 ) capacitor c=0.024152f //x=19.585 //y=5.02
c1154 ( 1022 0 ) capacitor c=0.053132f //x=18.715 //y=5.02
c1155 ( 1021 0 ) capacitor c=0.0452179f //x=16.535 //y=5.02
c1156 ( 1020 0 ) capacitor c=0.024152f //x=15.655 //y=5.02
c1157 ( 1019 0 ) capacitor c=0.024152f //x=14.775 //y=5.02
c1158 ( 1018 0 ) capacitor c=0.0531894f //x=13.905 //y=5.02
c1159 ( 1017 0 ) capacitor c=0.0380679f //x=12.025 //y=5.02
c1160 ( 1016 0 ) capacitor c=0.024008f //x=11.145 //y=5.02
c1161 ( 1015 0 ) capacitor c=0.049209f //x=10.275 //y=5.02
c1162 ( 1014 0 ) capacitor c=0.0452179f //x=8.395 //y=5.02
c1163 ( 1013 0 ) capacitor c=0.024152f //x=7.515 //y=5.02
c1164 ( 1012 0 ) capacitor c=0.024152f //x=6.635 //y=5.02
c1165 ( 1011 0 ) capacitor c=0.053132f //x=5.765 //y=5.02
c1166 ( 1010 0 ) capacitor c=0.0452179f //x=3.585 //y=5.02
c1167 ( 1009 0 ) capacitor c=0.024152f //x=2.705 //y=5.02
c1168 ( 1008 0 ) capacitor c=0.02424f //x=1.825 //y=5.02
c1169 ( 1007 0 ) capacitor c=0.0531407f //x=0.955 //y=5.02
c1170 ( 1006 0 ) capacitor c=0.113329f //x=84.36 //y=7.4
c1171 ( 1005 0 ) capacitor c=0.121198f //x=81.03 //y=7.4
c1172 ( 1004 0 ) capacitor c=0.00591168f //x=80.25 //y=7.4
c1173 ( 1003 0 ) capacitor c=0.00591168f //x=79.37 //y=7.4
c1174 ( 1002 0 ) capacitor c=0.00591168f //x=78.44 //y=7.4
c1175 ( 1000 0 ) capacitor c=0.115506f //x=77.7 //y=7.4
c1176 ( 999 0 ) capacitor c=0.00591168f //x=76.96 //y=7.4
c1177 ( 997 0 ) capacitor c=0.00591168f //x=76.04 //y=7.4
c1178 ( 996 0 ) capacitor c=0.00591168f //x=75.16 //y=7.4
c1179 ( 995 0 ) capacitor c=0.136591f //x=74.37 //y=7.4
c1180 ( 994 0 ) capacitor c=0.00591168f //x=73.26 //y=7.4
c1181 ( 992 0 ) capacitor c=0.00591168f //x=72.41 //y=7.4
c1182 ( 991 0 ) capacitor c=0.00591168f //x=71.53 //y=7.4
c1183 ( 990 0 ) capacitor c=0.00591168f //x=70.65 //y=7.4
c1184 ( 989 0 ) capacitor c=0.15714f //x=69.56 //y=7.4
c1185 ( 988 0 ) capacitor c=0.00591168f //x=68.45 //y=7.4
c1186 ( 986 0 ) capacitor c=0.00591168f //x=67.6 //y=7.4
c1187 ( 985 0 ) capacitor c=0.00591168f //x=66.72 //y=7.4
c1188 ( 984 0 ) capacitor c=0.00591168f //x=65.84 //y=7.4
c1189 ( 983 0 ) capacitor c=0.135038f //x=64.75 //y=7.4
c1190 ( 982 0 ) capacitor c=0.00591168f //x=63.97 //y=7.4
c1191 ( 981 0 ) capacitor c=0.00591168f //x=63.09 //y=7.4
c1192 ( 980 0 ) capacitor c=0.00591168f //x=62.21 //y=7.4
c1193 ( 979 0 ) capacitor c=0.134558f //x=61.42 //y=7.4
c1194 ( 978 0 ) capacitor c=0.00591168f //x=60.34 //y=7.4
c1195 ( 977 0 ) capacitor c=0.00591168f //x=59.46 //y=7.4
c1196 ( 976 0 ) capacitor c=0.00591168f //x=58.58 //y=7.4
c1197 ( 975 0 ) capacitor c=0.00591168f //x=57.72 //y=7.4
c1198 ( 973 0 ) capacitor c=0.15519f //x=56.61 //y=7.4
c1199 ( 972 0 ) capacitor c=0.00591168f //x=55.53 //y=7.4
c1200 ( 971 0 ) capacitor c=0.00591168f //x=54.65 //y=7.4
c1201 ( 970 0 ) capacitor c=0.00591168f //x=53.77 //y=7.4
c1202 ( 969 0 ) capacitor c=0.00591168f //x=52.91 //y=7.4
c1203 ( 967 0 ) capacitor c=0.139223f //x=51.8 //y=7.4
c1204 ( 966 0 ) capacitor c=0.00591168f //x=51.02 //y=7.4
c1205 ( 965 0 ) capacitor c=0.00591168f //x=50.14 //y=7.4
c1206 ( 964 0 ) capacitor c=0.00591168f //x=49.21 //y=7.4
c1207 ( 962 0 ) capacitor c=0.134558f //x=48.47 //y=7.4
c1208 ( 961 0 ) capacitor c=0.00591168f //x=47.39 //y=7.4
c1209 ( 960 0 ) capacitor c=0.00591168f //x=46.51 //y=7.4
c1210 ( 959 0 ) capacitor c=0.00591168f //x=45.63 //y=7.4
c1211 ( 958 0 ) capacitor c=0.00591168f //x=44.75 //y=7.4
c1212 ( 957 0 ) capacitor c=0.155081f //x=43.66 //y=7.4
c1213 ( 956 0 ) capacitor c=0.00591168f //x=42.58 //y=7.4
c1214 ( 955 0 ) capacitor c=0.00591168f //x=41.7 //y=7.4
c1215 ( 954 0 ) capacitor c=0.00591168f //x=40.82 //y=7.4
c1216 ( 953 0 ) capacitor c=0.00591168f //x=39.94 //y=7.4
c1217 ( 952 0 ) capacitor c=0.135038f //x=38.85 //y=7.4
c1218 ( 951 0 ) capacitor c=0.00591168f //x=38.11 //y=7.4
c1219 ( 949 0 ) capacitor c=0.00591168f //x=37.19 //y=7.4
c1220 ( 948 0 ) capacitor c=0.00591168f //x=36.31 //y=7.4
c1221 ( 947 0 ) capacitor c=0.134558f //x=35.52 //y=7.4
c1222 ( 946 0 ) capacitor c=0.00591168f //x=34.41 //y=7.4
c1223 ( 944 0 ) capacitor c=0.00591168f //x=33.56 //y=7.4
c1224 ( 943 0 ) capacitor c=0.00591168f //x=32.68 //y=7.4
c1225 ( 942 0 ) capacitor c=0.00591168f //x=31.8 //y=7.4
c1226 ( 941 0 ) capacitor c=0.15519f //x=30.71 //y=7.4
c1227 ( 940 0 ) capacitor c=0.00591168f //x=29.6 //y=7.4
c1228 ( 938 0 ) capacitor c=0.00591168f //x=28.75 //y=7.4
c1229 ( 937 0 ) capacitor c=0.00591168f //x=27.87 //y=7.4
c1230 ( 936 0 ) capacitor c=0.00591168f //x=26.99 //y=7.4
c1231 ( 935 0 ) capacitor c=0.139223f //x=25.9 //y=7.4
c1232 ( 934 0 ) capacitor c=0.00591168f //x=25.12 //y=7.4
c1233 ( 933 0 ) capacitor c=0.00591168f //x=24.24 //y=7.4
c1234 ( 932 0 ) capacitor c=0.00591168f //x=23.36 //y=7.4
c1235 ( 931 0 ) capacitor c=0.134712f //x=22.57 //y=7.4
c1236 ( 930 0 ) capacitor c=0.00591168f //x=21.49 //y=7.4
c1237 ( 929 0 ) capacitor c=0.00591168f //x=20.61 //y=7.4
c1238 ( 928 0 ) capacitor c=0.00591168f //x=19.73 //y=7.4
c1239 ( 927 0 ) capacitor c=0.00591168f //x=18.87 //y=7.4
c1240 ( 925 0 ) capacitor c=0.155081f //x=17.76 //y=7.4
c1241 ( 924 0 ) capacitor c=0.00591168f //x=16.68 //y=7.4
c1242 ( 923 0 ) capacitor c=0.00591168f //x=15.8 //y=7.4
c1243 ( 922 0 ) capacitor c=0.00591168f //x=14.92 //y=7.4
c1244 ( 921 0 ) capacitor c=0.00591168f //x=14.06 //y=7.4
c1245 ( 919 0 ) capacitor c=0.135038f //x=12.95 //y=7.4
c1246 ( 918 0 ) capacitor c=0.00591168f //x=12.17 //y=7.4
c1247 ( 917 0 ) capacitor c=0.00591168f //x=11.29 //y=7.4
c1248 ( 916 0 ) capacitor c=0.00591168f //x=10.36 //y=7.4
c1249 ( 914 0 ) capacitor c=0.134558f //x=9.62 //y=7.4
c1250 ( 913 0 ) capacitor c=0.00591168f //x=8.54 //y=7.4
c1251 ( 912 0 ) capacitor c=0.00591168f //x=7.66 //y=7.4
c1252 ( 911 0 ) capacitor c=0.00591168f //x=6.78 //y=7.4
c1253 ( 910 0 ) capacitor c=0.00591168f //x=5.9 //y=7.4
c1254 ( 909 0 ) capacitor c=0.15519f //x=4.81 //y=7.4
c1255 ( 908 0 ) capacitor c=0.00591168f //x=3.73 //y=7.4
c1256 ( 907 0 ) capacitor c=0.00591168f //x=2.85 //y=7.4
c1257 ( 906 0 ) capacitor c=0.00591168f //x=1.97 //y=7.4
c1258 ( 905 0 ) capacitor c=0.00591168f //x=1.09 //y=7.4
c1259 ( 902 0 ) capacitor c=0.334471f //x=86.95 //y=7.4
c1260 ( 887 0 ) capacitor c=0.120978f //x=84.19 //y=7.4
c1261 ( 881 0 ) capacitor c=0.0236224f //x=80.86 //y=7.4
c1262 ( 871 0 ) capacitor c=0.028539f //x=80.165 //y=7.4
c1263 ( 863 0 ) capacitor c=0.0285075f //x=79.285 //y=7.4
c1264 ( 855 0 ) capacitor c=0.0275884f //x=78.405 //y=7.4
c1265 ( 851 0 ) capacitor c=0.0275781f //x=77.53 //y=7.4
c1266 ( 843 0 ) capacitor c=0.0284327f //x=76.835 //y=7.4
c1267 ( 833 0 ) capacitor c=0.028862f //x=75.955 //y=7.4
c1268 ( 823 0 ) capacitor c=0.0240981f //x=75.075 //y=7.4
c1269 ( 819 0 ) capacitor c=0.0395206f //x=74.2 //y=7.4
c1270 ( 811 0 ) capacitor c=0.0288769f //x=73.205 //y=7.4
c1271 ( 801 0 ) capacitor c=0.0287757f //x=72.325 //y=7.4
c1272 ( 791 0 ) capacitor c=0.028511f //x=71.445 //y=7.4
c1273 ( 781 0 ) capacitor c=0.0383672f //x=70.565 //y=7.4
c1274 ( 777 0 ) capacitor c=0.0395206f //x=69.39 //y=7.4
c1275 ( 769 0 ) capacitor c=0.0288769f //x=68.395 //y=7.4
c1276 ( 759 0 ) capacitor c=0.0287624f //x=67.515 //y=7.4
c1277 ( 749 0 ) capacitor c=0.0284966f //x=66.635 //y=7.4
c1278 ( 739 0 ) capacitor c=0.0383672f //x=65.755 //y=7.4
c1279 ( 735 0 ) capacitor c=0.0236224f //x=64.58 //y=7.4
c1280 ( 725 0 ) capacitor c=0.0288359f //x=63.885 //y=7.4
c1281 ( 715 0 ) capacitor c=0.0288369f //x=63.005 //y=7.4
c1282 ( 707 0 ) capacitor c=0.0240981f //x=62.125 //y=7.4
c1283 ( 701 0 ) capacitor c=0.0394667f //x=61.25 //y=7.4
c1284 ( 691 0 ) capacitor c=0.0288488f //x=60.255 //y=7.4
c1285 ( 681 0 ) capacitor c=0.0287514f //x=59.375 //y=7.4
c1286 ( 673 0 ) capacitor c=0.0284966f //x=58.495 //y=7.4
c1287 ( 665 0 ) capacitor c=0.0383672f //x=57.615 //y=7.4
c1288 ( 659 0 ) capacitor c=0.0394667f //x=56.44 //y=7.4
c1289 ( 649 0 ) capacitor c=0.0288488f //x=55.445 //y=7.4
c1290 ( 639 0 ) capacitor c=0.0287505f //x=54.565 //y=7.4
c1291 ( 631 0 ) capacitor c=0.0284966f //x=53.685 //y=7.4
c1292 ( 623 0 ) capacitor c=0.0383672f //x=52.805 //y=7.4
c1293 ( 617 0 ) capacitor c=0.0236224f //x=51.63 //y=7.4
c1294 ( 607 0 ) capacitor c=0.0288359f //x=50.935 //y=7.4
c1295 ( 599 0 ) capacitor c=0.0288369f //x=50.055 //y=7.4
c1296 ( 591 0 ) capacitor c=0.0240981f //x=49.175 //y=7.4
c1297 ( 585 0 ) capacitor c=0.0394667f //x=48.3 //y=7.4
c1298 ( 575 0 ) capacitor c=0.0288488f //x=47.305 //y=7.4
c1299 ( 567 0 ) capacitor c=0.0287514f //x=46.425 //y=7.4
c1300 ( 557 0 ) capacitor c=0.0284966f //x=45.545 //y=7.4
c1301 ( 547 0 ) capacitor c=0.0383672f //x=44.665 //y=7.4
c1302 ( 541 0 ) capacitor c=0.0394667f //x=43.49 //y=7.4
c1303 ( 531 0 ) capacitor c=0.0288488f //x=42.495 //y=7.4
c1304 ( 523 0 ) capacitor c=0.0287505f //x=41.615 //y=7.4
c1305 ( 513 0 ) capacitor c=0.0284966f //x=40.735 //y=7.4
c1306 ( 503 0 ) capacitor c=0.0383672f //x=39.855 //y=7.4
c1307 ( 499 0 ) capacitor c=0.0236224f //x=38.68 //y=7.4
c1308 ( 491 0 ) capacitor c=0.0288359f //x=37.985 //y=7.4
c1309 ( 481 0 ) capacitor c=0.0288369f //x=37.105 //y=7.4
c1310 ( 471 0 ) capacitor c=0.0240981f //x=36.225 //y=7.4
c1311 ( 467 0 ) capacitor c=0.0394667f //x=35.35 //y=7.4
c1312 ( 459 0 ) capacitor c=0.0288488f //x=34.355 //y=7.4
c1313 ( 449 0 ) capacitor c=0.0287514f //x=33.475 //y=7.4
c1314 ( 439 0 ) capacitor c=0.0284966f //x=32.595 //y=7.4
c1315 ( 429 0 ) capacitor c=0.0383672f //x=31.715 //y=7.4
c1316 ( 425 0 ) capacitor c=0.0394667f //x=30.54 //y=7.4
c1317 ( 417 0 ) capacitor c=0.0288488f //x=29.545 //y=7.4
c1318 ( 407 0 ) capacitor c=0.0287505f //x=28.665 //y=7.4
c1319 ( 397 0 ) capacitor c=0.0284966f //x=27.785 //y=7.4
c1320 ( 387 0 ) capacitor c=0.0383672f //x=26.905 //y=7.4
c1321 ( 383 0 ) capacitor c=0.0236224f //x=25.73 //y=7.4
c1322 ( 373 0 ) capacitor c=0.0288359f //x=25.035 //y=7.4
c1323 ( 363 0 ) capacitor c=0.0288369f //x=24.155 //y=7.4
c1324 ( 355 0 ) capacitor c=0.0240981f //x=23.275 //y=7.4
c1325 ( 349 0 ) capacitor c=0.0394667f //x=22.4 //y=7.4
c1326 ( 339 0 ) capacitor c=0.0288488f //x=21.405 //y=7.4
c1327 ( 329 0 ) capacitor c=0.0287514f //x=20.525 //y=7.4
c1328 ( 321 0 ) capacitor c=0.0284966f //x=19.645 //y=7.4
c1329 ( 313 0 ) capacitor c=0.0383672f //x=18.765 //y=7.4
c1330 ( 307 0 ) capacitor c=0.0394667f //x=17.59 //y=7.4
c1331 ( 297 0 ) capacitor c=0.0288488f //x=16.595 //y=7.4
c1332 ( 287 0 ) capacitor c=0.0287505f //x=15.715 //y=7.4
c1333 ( 279 0 ) capacitor c=0.0284966f //x=14.835 //y=7.4
c1334 ( 271 0 ) capacitor c=0.0383672f //x=13.955 //y=7.4
c1335 ( 265 0 ) capacitor c=0.0236224f //x=12.78 //y=7.4
c1336 ( 255 0 ) capacitor c=0.0288359f //x=12.085 //y=7.4
c1337 ( 247 0 ) capacitor c=0.0288369f //x=11.205 //y=7.4
c1338 ( 239 0 ) capacitor c=0.0240981f //x=10.325 //y=7.4
c1339 ( 233 0 ) capacitor c=0.0394667f //x=9.45 //y=7.4
c1340 ( 223 0 ) capacitor c=0.0288488f //x=8.455 //y=7.4
c1341 ( 215 0 ) capacitor c=0.0287514f //x=7.575 //y=7.4
c1342 ( 205 0 ) capacitor c=0.0284966f //x=6.695 //y=7.4
c1343 ( 195 0 ) capacitor c=0.0383672f //x=5.815 //y=7.4
c1344 ( 189 0 ) capacitor c=0.0394667f //x=4.64 //y=7.4
c1345 ( 179 0 ) capacitor c=0.0288488f //x=3.645 //y=7.4
c1346 ( 171 0 ) capacitor c=0.0287505f //x=2.765 //y=7.4
c1347 ( 161 0 ) capacitor c=0.028511f //x=1.885 //y=7.4
c1348 ( 154 0 ) capacitor c=0.234426f //x=0.74 //y=7.4
c1349 ( 151 0 ) capacitor c=0.0452081f //x=1.005 //y=7.4
c1350 ( 147 0 ) capacitor c=2.90576f //x=86.95 //y=7.4
r1351 (  900 902 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=85.84 //y=7.4 //x2=86.95 //y2=7.4
r1352 (  898 900 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=84.73 //y=7.4 //x2=85.84 //y2=7.4
r1353 (  896 1006 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=84.53 //y=7.4 //x2=84.36 //y2=7.4
r1354 (  896 898 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=84.53 //y=7.4 //x2=84.73 //y2=7.4
r1355 (  890 892 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=82.14 //y=7.4 //x2=83.25 //y2=7.4
r1356 (  888 1005 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=81.2 //y=7.4 //x2=81.03 //y2=7.4
r1357 (  888 890 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=81.2 //y=7.4 //x2=82.14 //y2=7.4
r1358 (  887 1006 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=84.19 //y=7.4 //x2=84.36 //y2=7.4
r1359 (  887 892 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=84.19 //y=7.4 //x2=83.25 //y2=7.4
r1360 (  882 1004 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.335 //y=7.4 //x2=80.25 //y2=7.4
r1361 (  882 884 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=80.335 //y=7.4 //x2=80.66 //y2=7.4
r1362 (  881 1005 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=80.86 //y=7.4 //x2=81.03 //y2=7.4
r1363 (  881 884 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=80.86 //y=7.4 //x2=80.66 //y2=7.4
r1364 (  875 1004 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=80.25 //y=7.23 //x2=80.25 //y2=7.4
r1365 (  875 1075 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=80.25 //y=7.23 //x2=80.25 //y2=6.4
r1366 (  872 1003 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.455 //y=7.4 //x2=79.37 //y2=7.4
r1367 (  872 874 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=79.455 //y=7.4 //x2=79.55 //y2=7.4
r1368 (  871 1004 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.165 //y=7.4 //x2=80.25 //y2=7.4
r1369 (  871 874 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=80.165 //y=7.4 //x2=79.55 //y2=7.4
r1370 (  865 1003 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=79.37 //y=7.23 //x2=79.37 //y2=7.4
r1371 (  865 1074 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=79.37 //y=7.23 //x2=79.37 //y2=6.74
r1372 (  864 1002 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.575 //y=7.4 //x2=78.49 //y2=7.4
r1373 (  863 1003 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.285 //y=7.4 //x2=79.37 //y2=7.4
r1374 (  863 864 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=79.285 //y=7.4 //x2=78.575 //y2=7.4
r1375 (  857 1002 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=78.49 //y=7.23 //x2=78.49 //y2=7.4
r1376 (  857 1073 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=78.49 //y=7.23 //x2=78.49 //y2=6.4
r1377 (  856 1000 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=77.87 //y=7.4 //x2=77.7 //y2=7.4
r1378 (  855 1002 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.405 //y=7.4 //x2=78.49 //y2=7.4
r1379 (  855 856 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=78.405 //y=7.4 //x2=77.87 //y2=7.4
r1380 (  852 999 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=77.005 //y=7.4 //x2=76.92 //y2=7.4
r1381 (  851 1000 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=77.53 //y=7.4 //x2=77.7 //y2=7.4
r1382 (  851 852 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=77.53 //y=7.4 //x2=77.005 //y2=7.4
r1383 (  845 999 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.92 //y=7.23 //x2=76.92 //y2=7.4
r1384 (  845 1072 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=76.92 //y=7.23 //x2=76.92 //y2=6.745
r1385 (  844 997 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=76.125 //y=7.4 //x2=76.04 //y2=7.4
r1386 (  843 999 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=76.835 //y=7.4 //x2=76.92 //y2=7.4
r1387 (  843 844 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=76.835 //y=7.4 //x2=76.125 //y2=7.4
r1388 (  837 997 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.04 //y=7.23 //x2=76.04 //y2=7.4
r1389 (  837 1071 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=76.04 //y=7.23 //x2=76.04 //y2=6.745
r1390 (  834 996 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.245 //y=7.4 //x2=75.16 //y2=7.4
r1391 (  834 836 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=75.245 //y=7.4 //x2=75.85 //y2=7.4
r1392 (  833 997 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.955 //y=7.4 //x2=76.04 //y2=7.4
r1393 (  833 836 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=75.955 //y=7.4 //x2=75.85 //y2=7.4
r1394 (  827 996 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=75.16 //y=7.23 //x2=75.16 //y2=7.4
r1395 (  827 1070 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=75.16 //y=7.23 //x2=75.16 //y2=6.405
r1396 (  824 995 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=74.54 //y=7.4 //x2=74.37 //y2=7.4
r1397 (  824 826 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=74.54 //y=7.4 //x2=74.74 //y2=7.4
r1398 (  823 996 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.075 //y=7.4 //x2=75.16 //y2=7.4
r1399 (  823 826 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=75.075 //y=7.4 //x2=74.74 //y2=7.4
r1400 (  820 994 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.375 //y=7.4 //x2=73.29 //y2=7.4
r1401 (  819 995 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=74.2 //y=7.4 //x2=74.37 //y2=7.4
r1402 (  819 820 ) resistor r=29.5798 //w=0.357 //l=0.825 //layer=li \
 //thickness=0.1 //x=74.2 //y=7.4 //x2=73.375 //y2=7.4
r1403 (  813 994 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.29 //y=7.23 //x2=73.29 //y2=7.4
r1404 (  813 1069 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=73.29 //y=7.23 //x2=73.29 //y2=6.745
r1405 (  812 992 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.495 //y=7.4 //x2=72.41 //y2=7.4
r1406 (  811 994 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.205 //y=7.4 //x2=73.29 //y2=7.4
r1407 (  811 812 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=73.205 //y=7.4 //x2=72.495 //y2=7.4
r1408 (  805 992 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=72.41 //y=7.23 //x2=72.41 //y2=7.4
r1409 (  805 1068 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=72.41 //y=7.23 //x2=72.41 //y2=6.745
r1410 (  802 991 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.615 //y=7.4 //x2=71.53 //y2=7.4
r1411 (  802 804 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=71.615 //y=7.4 //x2=72.15 //y2=7.4
r1412 (  801 992 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.325 //y=7.4 //x2=72.41 //y2=7.4
r1413 (  801 804 ) resistor r=6.27451 //w=0.357 //l=0.175 //layer=li \
 //thickness=0.1 //x=72.325 //y=7.4 //x2=72.15 //y2=7.4
r1414 (  795 991 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=71.53 //y=7.23 //x2=71.53 //y2=7.4
r1415 (  795 1067 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=71.53 //y=7.23 //x2=71.53 //y2=6.745
r1416 (  792 990 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.735 //y=7.4 //x2=70.65 //y2=7.4
r1417 (  792 794 ) resistor r=10.9356 //w=0.357 //l=0.305 //layer=li \
 //thickness=0.1 //x=70.735 //y=7.4 //x2=71.04 //y2=7.4
r1418 (  791 991 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.445 //y=7.4 //x2=71.53 //y2=7.4
r1419 (  791 794 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=71.445 //y=7.4 //x2=71.04 //y2=7.4
r1420 (  785 990 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=70.65 //y=7.23 //x2=70.65 //y2=7.4
r1421 (  785 1066 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=70.65 //y=7.23 //x2=70.65 //y2=6.405
r1422 (  782 989 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=69.73 //y=7.4 //x2=69.56 //y2=7.4
r1423 (  782 784 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=69.73 //y=7.4 //x2=69.93 //y2=7.4
r1424 (  781 990 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.565 //y=7.4 //x2=70.65 //y2=7.4
r1425 (  781 784 ) resistor r=22.7675 //w=0.357 //l=0.635 //layer=li \
 //thickness=0.1 //x=70.565 //y=7.4 //x2=69.93 //y2=7.4
r1426 (  778 988 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.565 //y=7.4 //x2=68.48 //y2=7.4
r1427 (  777 989 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=69.39 //y=7.4 //x2=69.56 //y2=7.4
r1428 (  777 778 ) resistor r=29.5798 //w=0.357 //l=0.825 //layer=li \
 //thickness=0.1 //x=69.39 //y=7.4 //x2=68.565 //y2=7.4
r1429 (  771 988 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.48 //y=7.23 //x2=68.48 //y2=7.4
r1430 (  771 1065 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=68.48 //y=7.23 //x2=68.48 //y2=6.745
r1431 (  770 986 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.685 //y=7.4 //x2=67.6 //y2=7.4
r1432 (  769 988 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.395 //y=7.4 //x2=68.48 //y2=7.4
r1433 (  769 770 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=68.395 //y=7.4 //x2=67.685 //y2=7.4
r1434 (  763 986 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.6 //y=7.23 //x2=67.6 //y2=7.4
r1435 (  763 1064 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=67.6 //y=7.23 //x2=67.6 //y2=6.745
r1436 (  760 985 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.805 //y=7.4 //x2=66.72 //y2=7.4
r1437 (  760 762 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=66.805 //y=7.4 //x2=67.34 //y2=7.4
r1438 (  759 986 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.515 //y=7.4 //x2=67.6 //y2=7.4
r1439 (  759 762 ) resistor r=6.27451 //w=0.357 //l=0.175 //layer=li \
 //thickness=0.1 //x=67.515 //y=7.4 //x2=67.34 //y2=7.4
r1440 (  753 985 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=66.72 //y=7.23 //x2=66.72 //y2=7.4
r1441 (  753 1063 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=66.72 //y=7.23 //x2=66.72 //y2=6.745
r1442 (  750 984 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.925 //y=7.4 //x2=65.84 //y2=7.4
r1443 (  750 752 ) resistor r=10.9356 //w=0.357 //l=0.305 //layer=li \
 //thickness=0.1 //x=65.925 //y=7.4 //x2=66.23 //y2=7.4
r1444 (  749 985 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.635 //y=7.4 //x2=66.72 //y2=7.4
r1445 (  749 752 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=66.635 //y=7.4 //x2=66.23 //y2=7.4
r1446 (  743 984 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=65.84 //y=7.23 //x2=65.84 //y2=7.4
r1447 (  743 1062 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=65.84 //y=7.23 //x2=65.84 //y2=6.405
r1448 (  740 983 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.92 //y=7.4 //x2=64.75 //y2=7.4
r1449 (  740 742 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=64.92 //y=7.4 //x2=65.12 //y2=7.4
r1450 (  739 984 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.755 //y=7.4 //x2=65.84 //y2=7.4
r1451 (  739 742 ) resistor r=22.7675 //w=0.357 //l=0.635 //layer=li \
 //thickness=0.1 //x=65.755 //y=7.4 //x2=65.12 //y2=7.4
r1452 (  736 982 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.055 //y=7.4 //x2=63.97 //y2=7.4
r1453 (  735 983 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.58 //y=7.4 //x2=64.75 //y2=7.4
r1454 (  735 736 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=64.58 //y=7.4 //x2=64.055 //y2=7.4
r1455 (  729 982 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=63.97 //y=7.23 //x2=63.97 //y2=7.4
r1456 (  729 1061 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=63.97 //y=7.23 //x2=63.97 //y2=6.745
r1457 (  726 981 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.175 //y=7.4 //x2=63.09 //y2=7.4
r1458 (  726 728 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=63.175 //y=7.4 //x2=63.64 //y2=7.4
r1459 (  725 982 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.885 //y=7.4 //x2=63.97 //y2=7.4
r1460 (  725 728 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=63.885 //y=7.4 //x2=63.64 //y2=7.4
r1461 (  719 981 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=63.09 //y=7.23 //x2=63.09 //y2=7.4
r1462 (  719 1060 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=63.09 //y=7.23 //x2=63.09 //y2=6.745
r1463 (  716 980 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.295 //y=7.4 //x2=62.21 //y2=7.4
r1464 (  716 718 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=62.295 //y=7.4 //x2=62.53 //y2=7.4
r1465 (  715 981 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.005 //y=7.4 //x2=63.09 //y2=7.4
r1466 (  715 718 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=63.005 //y=7.4 //x2=62.53 //y2=7.4
r1467 (  709 980 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.21 //y=7.23 //x2=62.21 //y2=7.4
r1468 (  709 1059 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=62.21 //y=7.23 //x2=62.21 //y2=6.405
r1469 (  708 979 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.59 //y=7.4 //x2=61.42 //y2=7.4
r1470 (  707 980 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.125 //y=7.4 //x2=62.21 //y2=7.4
r1471 (  707 708 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=62.125 //y=7.4 //x2=61.59 //y2=7.4
r1472 (  702 978 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.425 //y=7.4 //x2=60.34 //y2=7.4
r1473 (  702 704 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=60.425 //y=7.4 //x2=61.05 //y2=7.4
r1474 (  701 979 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.25 //y=7.4 //x2=61.42 //y2=7.4
r1475 (  701 704 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=61.25 //y=7.4 //x2=61.05 //y2=7.4
r1476 (  695 978 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=60.34 //y=7.23 //x2=60.34 //y2=7.4
r1477 (  695 1058 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=60.34 //y=7.23 //x2=60.34 //y2=6.745
r1478 (  692 977 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.545 //y=7.4 //x2=59.46 //y2=7.4
r1479 (  692 694 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=59.545 //y=7.4 //x2=59.94 //y2=7.4
r1480 (  691 978 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.255 //y=7.4 //x2=60.34 //y2=7.4
r1481 (  691 694 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=60.255 //y=7.4 //x2=59.94 //y2=7.4
r1482 (  685 977 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=59.46 //y=7.23 //x2=59.46 //y2=7.4
r1483 (  685 1057 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=59.46 //y=7.23 //x2=59.46 //y2=6.745
r1484 (  682 976 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.665 //y=7.4 //x2=58.58 //y2=7.4
r1485 (  682 684 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=58.665 //y=7.4 //x2=58.83 //y2=7.4
r1486 (  681 977 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.375 //y=7.4 //x2=59.46 //y2=7.4
r1487 (  681 684 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=59.375 //y=7.4 //x2=58.83 //y2=7.4
r1488 (  675 976 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.58 //y=7.23 //x2=58.58 //y2=7.4
r1489 (  675 1056 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=58.58 //y=7.23 //x2=58.58 //y2=6.745
r1490 (  674 975 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=57.785 //y=7.4 //x2=57.7 //y2=7.4
r1491 (  673 976 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.495 //y=7.4 //x2=58.58 //y2=7.4
r1492 (  673 674 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=58.495 //y=7.4 //x2=57.785 //y2=7.4
r1493 (  667 975 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.7 //y=7.23 //x2=57.7 //y2=7.4
r1494 (  667 1055 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=57.7 //y=7.23 //x2=57.7 //y2=6.405
r1495 (  666 973 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=56.78 //y=7.4 //x2=56.61 //y2=7.4
r1496 (  665 975 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=57.615 //y=7.4 //x2=57.7 //y2=7.4
r1497 (  665 666 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=57.615 //y=7.4 //x2=56.78 //y2=7.4
r1498 (  660 972 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.615 //y=7.4 //x2=55.53 //y2=7.4
r1499 (  660 662 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=55.615 //y=7.4 //x2=56.24 //y2=7.4
r1500 (  659 973 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=56.44 //y=7.4 //x2=56.61 //y2=7.4
r1501 (  659 662 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=56.44 //y=7.4 //x2=56.24 //y2=7.4
r1502 (  653 972 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=55.53 //y=7.23 //x2=55.53 //y2=7.4
r1503 (  653 1054 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=55.53 //y=7.23 //x2=55.53 //y2=6.745
r1504 (  650 971 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.735 //y=7.4 //x2=54.65 //y2=7.4
r1505 (  650 652 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=54.735 //y=7.4 //x2=55.13 //y2=7.4
r1506 (  649 972 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.445 //y=7.4 //x2=55.53 //y2=7.4
r1507 (  649 652 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=55.445 //y=7.4 //x2=55.13 //y2=7.4
r1508 (  643 971 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=54.65 //y=7.23 //x2=54.65 //y2=7.4
r1509 (  643 1053 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=54.65 //y=7.23 //x2=54.65 //y2=6.745
r1510 (  640 970 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.855 //y=7.4 //x2=53.77 //y2=7.4
r1511 (  640 642 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=53.855 //y=7.4 //x2=54.02 //y2=7.4
r1512 (  639 971 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.565 //y=7.4 //x2=54.65 //y2=7.4
r1513 (  639 642 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=54.565 //y=7.4 //x2=54.02 //y2=7.4
r1514 (  633 970 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=53.77 //y=7.23 //x2=53.77 //y2=7.4
r1515 (  633 1052 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=53.77 //y=7.23 //x2=53.77 //y2=6.745
r1516 (  632 969 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=52.975 //y=7.4 //x2=52.89 //y2=7.4
r1517 (  631 970 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.685 //y=7.4 //x2=53.77 //y2=7.4
r1518 (  631 632 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=53.685 //y=7.4 //x2=52.975 //y2=7.4
r1519 (  625 969 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=52.89 //y=7.23 //x2=52.89 //y2=7.4
r1520 (  625 1051 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=52.89 //y=7.23 //x2=52.89 //y2=6.405
r1521 (  624 967 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=51.97 //y=7.4 //x2=51.8 //y2=7.4
r1522 (  623 969 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=52.805 //y=7.4 //x2=52.89 //y2=7.4
r1523 (  623 624 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=52.805 //y=7.4 //x2=51.97 //y2=7.4
r1524 (  618 966 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.105 //y=7.4 //x2=51.02 //y2=7.4
r1525 (  618 620 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=51.105 //y=7.4 //x2=51.43 //y2=7.4
r1526 (  617 967 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=51.63 //y=7.4 //x2=51.8 //y2=7.4
r1527 (  617 620 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=51.63 //y=7.4 //x2=51.43 //y2=7.4
r1528 (  611 966 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=51.02 //y=7.23 //x2=51.02 //y2=7.4
r1529 (  611 1050 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=51.02 //y=7.23 //x2=51.02 //y2=6.745
r1530 (  608 965 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.225 //y=7.4 //x2=50.14 //y2=7.4
r1531 (  608 610 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=50.225 //y=7.4 //x2=50.32 //y2=7.4
r1532 (  607 966 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.935 //y=7.4 //x2=51.02 //y2=7.4
r1533 (  607 610 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=50.935 //y=7.4 //x2=50.32 //y2=7.4
r1534 (  601 965 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=50.14 //y=7.23 //x2=50.14 //y2=7.4
r1535 (  601 1049 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=50.14 //y=7.23 //x2=50.14 //y2=6.745
r1536 (  600 964 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.345 //y=7.4 //x2=49.26 //y2=7.4
r1537 (  599 965 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.055 //y=7.4 //x2=50.14 //y2=7.4
r1538 (  599 600 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=50.055 //y=7.4 //x2=49.345 //y2=7.4
r1539 (  593 964 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.26 //y=7.23 //x2=49.26 //y2=7.4
r1540 (  593 1048 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=49.26 //y=7.23 //x2=49.26 //y2=6.405
r1541 (  592 962 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.64 //y=7.4 //x2=48.47 //y2=7.4
r1542 (  591 964 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.175 //y=7.4 //x2=49.26 //y2=7.4
r1543 (  591 592 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=49.175 //y=7.4 //x2=48.64 //y2=7.4
r1544 (  586 961 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.475 //y=7.4 //x2=47.39 //y2=7.4
r1545 (  586 588 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=47.475 //y=7.4 //x2=47.73 //y2=7.4
r1546 (  585 962 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.3 //y=7.4 //x2=48.47 //y2=7.4
r1547 (  585 588 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=48.3 //y=7.4 //x2=47.73 //y2=7.4
r1548 (  579 961 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.39 //y=7.23 //x2=47.39 //y2=7.4
r1549 (  579 1047 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=47.39 //y=7.23 //x2=47.39 //y2=6.745
r1550 (  576 960 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.595 //y=7.4 //x2=46.51 //y2=7.4
r1551 (  576 578 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=46.595 //y=7.4 //x2=46.62 //y2=7.4
r1552 (  575 961 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.305 //y=7.4 //x2=47.39 //y2=7.4
r1553 (  575 578 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=47.305 //y=7.4 //x2=46.62 //y2=7.4
r1554 (  569 960 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=46.51 //y=7.23 //x2=46.51 //y2=7.4
r1555 (  569 1046 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.51 //y=7.23 //x2=46.51 //y2=6.745
r1556 (  568 959 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.715 //y=7.4 //x2=45.63 //y2=7.4
r1557 (  567 960 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.425 //y=7.4 //x2=46.51 //y2=7.4
r1558 (  567 568 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=46.425 //y=7.4 //x2=45.715 //y2=7.4
r1559 (  561 959 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=45.63 //y=7.23 //x2=45.63 //y2=7.4
r1560 (  561 1045 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=45.63 //y=7.23 //x2=45.63 //y2=6.745
r1561 (  558 958 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.835 //y=7.4 //x2=44.75 //y2=7.4
r1562 (  558 560 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=44.835 //y=7.4 //x2=45.51 //y2=7.4
r1563 (  557 959 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.545 //y=7.4 //x2=45.63 //y2=7.4
r1564 (  557 560 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=45.545 //y=7.4 //x2=45.51 //y2=7.4
r1565 (  551 958 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=44.75 //y=7.23 //x2=44.75 //y2=7.4
r1566 (  551 1044 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=44.75 //y=7.23 //x2=44.75 //y2=6.405
r1567 (  548 957 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.83 //y=7.4 //x2=43.66 //y2=7.4
r1568 (  548 550 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.83 //y=7.4 //x2=44.4 //y2=7.4
r1569 (  547 958 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=44.665 //y=7.4 //x2=44.75 //y2=7.4
r1570 (  547 550 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=44.665 //y=7.4 //x2=44.4 //y2=7.4
r1571 (  542 956 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.665 //y=7.4 //x2=42.58 //y2=7.4
r1572 (  542 544 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=42.665 //y=7.4 //x2=42.92 //y2=7.4
r1573 (  541 957 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.49 //y=7.4 //x2=43.66 //y2=7.4
r1574 (  541 544 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.49 //y=7.4 //x2=42.92 //y2=7.4
r1575 (  535 956 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=42.58 //y=7.23 //x2=42.58 //y2=7.4
r1576 (  535 1043 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=42.58 //y=7.23 //x2=42.58 //y2=6.745
r1577 (  532 955 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.785 //y=7.4 //x2=41.7 //y2=7.4
r1578 (  532 534 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=41.785 //y=7.4 //x2=41.81 //y2=7.4
r1579 (  531 956 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.495 //y=7.4 //x2=42.58 //y2=7.4
r1580 (  531 534 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=42.495 //y=7.4 //x2=41.81 //y2=7.4
r1581 (  525 955 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=41.7 //y=7.23 //x2=41.7 //y2=7.4
r1582 (  525 1042 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=41.7 //y=7.23 //x2=41.7 //y2=6.745
r1583 (  524 954 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.905 //y=7.4 //x2=40.82 //y2=7.4
r1584 (  523 955 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.615 //y=7.4 //x2=41.7 //y2=7.4
r1585 (  523 524 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=41.615 //y=7.4 //x2=40.905 //y2=7.4
r1586 (  517 954 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.82 //y=7.23 //x2=40.82 //y2=7.4
r1587 (  517 1041 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=40.82 //y=7.23 //x2=40.82 //y2=6.745
r1588 (  514 953 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.025 //y=7.4 //x2=39.94 //y2=7.4
r1589 (  514 516 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=40.025 //y=7.4 //x2=40.7 //y2=7.4
r1590 (  513 954 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.735 //y=7.4 //x2=40.82 //y2=7.4
r1591 (  513 516 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=40.735 //y=7.4 //x2=40.7 //y2=7.4
r1592 (  507 953 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.94 //y=7.23 //x2=39.94 //y2=7.4
r1593 (  507 1040 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=39.94 //y=7.23 //x2=39.94 //y2=6.405
r1594 (  504 952 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.02 //y=7.4 //x2=38.85 //y2=7.4
r1595 (  504 506 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=39.02 //y=7.4 //x2=39.59 //y2=7.4
r1596 (  503 953 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.855 //y=7.4 //x2=39.94 //y2=7.4
r1597 (  503 506 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=39.855 //y=7.4 //x2=39.59 //y2=7.4
r1598 (  500 951 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.155 //y=7.4 //x2=38.07 //y2=7.4
r1599 (  499 952 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.68 //y=7.4 //x2=38.85 //y2=7.4
r1600 (  499 500 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=38.68 //y=7.4 //x2=38.155 //y2=7.4
r1601 (  493 951 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.07 //y=7.23 //x2=38.07 //y2=7.4
r1602 (  493 1039 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=38.07 //y=7.23 //x2=38.07 //y2=6.745
r1603 (  492 949 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.275 //y=7.4 //x2=37.19 //y2=7.4
r1604 (  491 951 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.985 //y=7.4 //x2=38.07 //y2=7.4
r1605 (  491 492 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=37.985 //y=7.4 //x2=37.275 //y2=7.4
r1606 (  485 949 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.19 //y=7.23 //x2=37.19 //y2=7.4
r1607 (  485 1038 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=37.19 //y=7.23 //x2=37.19 //y2=6.745
r1608 (  482 948 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.395 //y=7.4 //x2=36.31 //y2=7.4
r1609 (  482 484 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=36.395 //y=7.4 //x2=37 //y2=7.4
r1610 (  481 949 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.105 //y=7.4 //x2=37.19 //y2=7.4
r1611 (  481 484 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=37.105 //y=7.4 //x2=37 //y2=7.4
r1612 (  475 948 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.31 //y=7.23 //x2=36.31 //y2=7.4
r1613 (  475 1037 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=36.31 //y=7.23 //x2=36.31 //y2=6.405
r1614 (  472 947 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=35.69 //y=7.4 //x2=35.52 //y2=7.4
r1615 (  472 474 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=35.69 //y=7.4 //x2=35.89 //y2=7.4
r1616 (  471 948 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.225 //y=7.4 //x2=36.31 //y2=7.4
r1617 (  471 474 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=36.225 //y=7.4 //x2=35.89 //y2=7.4
r1618 (  468 946 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.525 //y=7.4 //x2=34.44 //y2=7.4
r1619 (  467 947 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=35.35 //y=7.4 //x2=35.52 //y2=7.4
r1620 (  467 468 ) resistor r=29.5798 //w=0.357 //l=0.825 //layer=li \
 //thickness=0.1 //x=35.35 //y=7.4 //x2=34.525 //y2=7.4
r1621 (  461 946 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=34.44 //y=7.23 //x2=34.44 //y2=7.4
r1622 (  461 1036 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=34.44 //y=7.23 //x2=34.44 //y2=6.745
r1623 (  460 944 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.645 //y=7.4 //x2=33.56 //y2=7.4
r1624 (  459 946 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.355 //y=7.4 //x2=34.44 //y2=7.4
r1625 (  459 460 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=34.355 //y=7.4 //x2=33.645 //y2=7.4
r1626 (  453 944 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.56 //y=7.23 //x2=33.56 //y2=7.4
r1627 (  453 1035 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=33.56 //y=7.23 //x2=33.56 //y2=6.745
r1628 (  450 943 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.765 //y=7.4 //x2=32.68 //y2=7.4
r1629 (  450 452 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=32.765 //y=7.4 //x2=33.3 //y2=7.4
r1630 (  449 944 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.475 //y=7.4 //x2=33.56 //y2=7.4
r1631 (  449 452 ) resistor r=6.27451 //w=0.357 //l=0.175 //layer=li \
 //thickness=0.1 //x=33.475 //y=7.4 //x2=33.3 //y2=7.4
r1632 (  443 943 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.68 //y=7.23 //x2=32.68 //y2=7.4
r1633 (  443 1034 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=32.68 //y=7.23 //x2=32.68 //y2=6.745
r1634 (  440 942 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.885 //y=7.4 //x2=31.8 //y2=7.4
r1635 (  440 442 ) resistor r=10.9356 //w=0.357 //l=0.305 //layer=li \
 //thickness=0.1 //x=31.885 //y=7.4 //x2=32.19 //y2=7.4
r1636 (  439 943 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.595 //y=7.4 //x2=32.68 //y2=7.4
r1637 (  439 442 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=32.595 //y=7.4 //x2=32.19 //y2=7.4
r1638 (  433 942 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=31.8 //y=7.23 //x2=31.8 //y2=7.4
r1639 (  433 1033 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=31.8 //y=7.23 //x2=31.8 //y2=6.405
r1640 (  430 941 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.88 //y=7.4 //x2=30.71 //y2=7.4
r1641 (  430 432 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=30.88 //y=7.4 //x2=31.08 //y2=7.4
r1642 (  429 942 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.715 //y=7.4 //x2=31.8 //y2=7.4
r1643 (  429 432 ) resistor r=22.7675 //w=0.357 //l=0.635 //layer=li \
 //thickness=0.1 //x=31.715 //y=7.4 //x2=31.08 //y2=7.4
r1644 (  426 940 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.715 //y=7.4 //x2=29.63 //y2=7.4
r1645 (  425 941 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.54 //y=7.4 //x2=30.71 //y2=7.4
r1646 (  425 426 ) resistor r=29.5798 //w=0.357 //l=0.825 //layer=li \
 //thickness=0.1 //x=30.54 //y=7.4 //x2=29.715 //y2=7.4
r1647 (  419 940 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.63 //y=7.23 //x2=29.63 //y2=7.4
r1648 (  419 1032 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=29.63 //y=7.23 //x2=29.63 //y2=6.745
r1649 (  418 938 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.835 //y=7.4 //x2=28.75 //y2=7.4
r1650 (  417 940 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.545 //y=7.4 //x2=29.63 //y2=7.4
r1651 (  417 418 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=29.545 //y=7.4 //x2=28.835 //y2=7.4
r1652 (  411 938 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=28.75 //y=7.23 //x2=28.75 //y2=7.4
r1653 (  411 1031 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=28.75 //y=7.23 //x2=28.75 //y2=6.745
r1654 (  408 937 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.955 //y=7.4 //x2=27.87 //y2=7.4
r1655 (  408 410 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=27.955 //y=7.4 //x2=28.49 //y2=7.4
r1656 (  407 938 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.665 //y=7.4 //x2=28.75 //y2=7.4
r1657 (  407 410 ) resistor r=6.27451 //w=0.357 //l=0.175 //layer=li \
 //thickness=0.1 //x=28.665 //y=7.4 //x2=28.49 //y2=7.4
r1658 (  401 937 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.87 //y=7.23 //x2=27.87 //y2=7.4
r1659 (  401 1030 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=27.87 //y=7.23 //x2=27.87 //y2=6.745
r1660 (  398 936 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.075 //y=7.4 //x2=26.99 //y2=7.4
r1661 (  398 400 ) resistor r=10.9356 //w=0.357 //l=0.305 //layer=li \
 //thickness=0.1 //x=27.075 //y=7.4 //x2=27.38 //y2=7.4
r1662 (  397 937 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.785 //y=7.4 //x2=27.87 //y2=7.4
r1663 (  397 400 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=27.785 //y=7.4 //x2=27.38 //y2=7.4
r1664 (  391 936 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.99 //y=7.23 //x2=26.99 //y2=7.4
r1665 (  391 1029 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=26.99 //y=7.23 //x2=26.99 //y2=6.405
r1666 (  388 935 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.07 //y=7.4 //x2=25.9 //y2=7.4
r1667 (  388 390 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=26.07 //y=7.4 //x2=26.27 //y2=7.4
r1668 (  387 936 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.905 //y=7.4 //x2=26.99 //y2=7.4
r1669 (  387 390 ) resistor r=22.7675 //w=0.357 //l=0.635 //layer=li \
 //thickness=0.1 //x=26.905 //y=7.4 //x2=26.27 //y2=7.4
r1670 (  384 934 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.205 //y=7.4 //x2=25.12 //y2=7.4
r1671 (  383 935 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.73 //y=7.4 //x2=25.9 //y2=7.4
r1672 (  383 384 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=25.73 //y=7.4 //x2=25.205 //y2=7.4
r1673 (  377 934 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.12 //y=7.23 //x2=25.12 //y2=7.4
r1674 (  377 1028 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=25.12 //y=7.23 //x2=25.12 //y2=6.745
r1675 (  374 933 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.325 //y=7.4 //x2=24.24 //y2=7.4
r1676 (  374 376 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=24.325 //y=7.4 //x2=24.79 //y2=7.4
r1677 (  373 934 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.035 //y=7.4 //x2=25.12 //y2=7.4
r1678 (  373 376 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=25.035 //y=7.4 //x2=24.79 //y2=7.4
r1679 (  367 933 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.24 //y=7.23 //x2=24.24 //y2=7.4
r1680 (  367 1027 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=24.24 //y=7.23 //x2=24.24 //y2=6.745
r1681 (  364 932 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.445 //y=7.4 //x2=23.36 //y2=7.4
r1682 (  364 366 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=23.445 //y=7.4 //x2=23.68 //y2=7.4
r1683 (  363 933 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.155 //y=7.4 //x2=24.24 //y2=7.4
r1684 (  363 366 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=24.155 //y=7.4 //x2=23.68 //y2=7.4
r1685 (  357 932 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.36 //y=7.23 //x2=23.36 //y2=7.4
r1686 (  357 1026 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=23.36 //y=7.23 //x2=23.36 //y2=6.405
r1687 (  356 931 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.74 //y=7.4 //x2=22.57 //y2=7.4
r1688 (  355 932 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.275 //y=7.4 //x2=23.36 //y2=7.4
r1689 (  355 356 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=23.275 //y=7.4 //x2=22.74 //y2=7.4
r1690 (  350 930 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.575 //y=7.4 //x2=21.49 //y2=7.4
r1691 (  350 352 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=21.575 //y=7.4 //x2=22.2 //y2=7.4
r1692 (  349 931 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.4 //y=7.4 //x2=22.57 //y2=7.4
r1693 (  349 352 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=22.4 //y=7.4 //x2=22.2 //y2=7.4
r1694 (  343 930 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.49 //y=7.23 //x2=21.49 //y2=7.4
r1695 (  343 1025 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.49 //y=7.23 //x2=21.49 //y2=6.745
r1696 (  340 929 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.695 //y=7.4 //x2=20.61 //y2=7.4
r1697 (  340 342 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=20.695 //y=7.4 //x2=21.09 //y2=7.4
r1698 (  339 930 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.405 //y=7.4 //x2=21.49 //y2=7.4
r1699 (  339 342 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=21.405 //y=7.4 //x2=21.09 //y2=7.4
r1700 (  333 929 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.61 //y=7.23 //x2=20.61 //y2=7.4
r1701 (  333 1024 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.61 //y=7.23 //x2=20.61 //y2=6.745
r1702 (  330 928 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.815 //y=7.4 //x2=19.73 //y2=7.4
r1703 (  330 332 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=19.815 //y=7.4 //x2=19.98 //y2=7.4
r1704 (  329 929 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.525 //y=7.4 //x2=20.61 //y2=7.4
r1705 (  329 332 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=20.525 //y=7.4 //x2=19.98 //y2=7.4
r1706 (  323 928 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.73 //y=7.23 //x2=19.73 //y2=7.4
r1707 (  323 1023 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=19.73 //y=7.23 //x2=19.73 //y2=6.745
r1708 (  322 927 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.935 //y=7.4 //x2=18.85 //y2=7.4
r1709 (  321 928 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.645 //y=7.4 //x2=19.73 //y2=7.4
r1710 (  321 322 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=19.645 //y=7.4 //x2=18.935 //y2=7.4
r1711 (  315 927 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.85 //y=7.23 //x2=18.85 //y2=7.4
r1712 (  315 1022 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=18.85 //y=7.23 //x2=18.85 //y2=6.405
r1713 (  314 925 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.93 //y=7.4 //x2=17.76 //y2=7.4
r1714 (  313 927 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.765 //y=7.4 //x2=18.85 //y2=7.4
r1715 (  313 314 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=18.765 //y=7.4 //x2=17.93 //y2=7.4
r1716 (  308 924 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.765 //y=7.4 //x2=16.68 //y2=7.4
r1717 (  308 310 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=16.765 //y=7.4 //x2=17.39 //y2=7.4
r1718 (  307 925 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.59 //y=7.4 //x2=17.76 //y2=7.4
r1719 (  307 310 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=17.59 //y=7.4 //x2=17.39 //y2=7.4
r1720 (  301 924 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.68 //y=7.23 //x2=16.68 //y2=7.4
r1721 (  301 1021 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.68 //y=7.23 //x2=16.68 //y2=6.745
r1722 (  298 923 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.885 //y=7.4 //x2=15.8 //y2=7.4
r1723 (  298 300 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=15.885 //y=7.4 //x2=16.28 //y2=7.4
r1724 (  297 924 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.595 //y=7.4 //x2=16.68 //y2=7.4
r1725 (  297 300 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=16.595 //y=7.4 //x2=16.28 //y2=7.4
r1726 (  291 923 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.8 //y=7.23 //x2=15.8 //y2=7.4
r1727 (  291 1020 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.8 //y=7.23 //x2=15.8 //y2=6.745
r1728 (  288 922 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.005 //y=7.4 //x2=14.92 //y2=7.4
r1729 (  288 290 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=15.005 //y=7.4 //x2=15.17 //y2=7.4
r1730 (  287 923 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.715 //y=7.4 //x2=15.8 //y2=7.4
r1731 (  287 290 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=15.715 //y=7.4 //x2=15.17 //y2=7.4
r1732 (  281 922 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.92 //y=7.23 //x2=14.92 //y2=7.4
r1733 (  281 1019 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.92 //y=7.23 //x2=14.92 //y2=6.745
r1734 (  280 921 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.125 //y=7.4 //x2=14.04 //y2=7.4
r1735 (  279 922 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.835 //y=7.4 //x2=14.92 //y2=7.4
r1736 (  279 280 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=14.835 //y=7.4 //x2=14.125 //y2=7.4
r1737 (  273 921 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.04 //y=7.23 //x2=14.04 //y2=7.4
r1738 (  273 1018 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=14.04 //y=7.23 //x2=14.04 //y2=6.405
r1739 (  272 919 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.12 //y=7.4 //x2=12.95 //y2=7.4
r1740 (  271 921 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.955 //y=7.4 //x2=14.04 //y2=7.4
r1741 (  271 272 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=13.955 //y=7.4 //x2=13.12 //y2=7.4
r1742 (  266 918 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.255 //y=7.4 //x2=12.17 //y2=7.4
r1743 (  266 268 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=12.255 //y=7.4 //x2=12.58 //y2=7.4
r1744 (  265 919 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.78 //y=7.4 //x2=12.95 //y2=7.4
r1745 (  265 268 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.78 //y=7.4 //x2=12.58 //y2=7.4
r1746 (  259 918 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.17 //y=7.23 //x2=12.17 //y2=7.4
r1747 (  259 1017 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.17 //y=7.23 //x2=12.17 //y2=6.745
r1748 (  256 917 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.375 //y=7.4 //x2=11.29 //y2=7.4
r1749 (  256 258 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=11.375 //y=7.4 //x2=11.47 //y2=7.4
r1750 (  255 918 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.085 //y=7.4 //x2=12.17 //y2=7.4
r1751 (  255 258 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=12.085 //y=7.4 //x2=11.47 //y2=7.4
r1752 (  249 917 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.29 //y=7.23 //x2=11.29 //y2=7.4
r1753 (  249 1016 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.29 //y=7.23 //x2=11.29 //y2=6.745
r1754 (  248 916 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.495 //y=7.4 //x2=10.41 //y2=7.4
r1755 (  247 917 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.205 //y=7.4 //x2=11.29 //y2=7.4
r1756 (  247 248 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.205 //y=7.4 //x2=10.495 //y2=7.4
r1757 (  241 916 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.41 //y=7.23 //x2=10.41 //y2=7.4
r1758 (  241 1015 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=10.41 //y=7.23 //x2=10.41 //y2=6.405
r1759 (  240 914 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.79 //y=7.4 //x2=9.62 //y2=7.4
r1760 (  239 916 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.325 //y=7.4 //x2=10.41 //y2=7.4
r1761 (  239 240 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=10.325 //y=7.4 //x2=9.79 //y2=7.4
r1762 (  234 913 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.625 //y=7.4 //x2=8.54 //y2=7.4
r1763 (  234 236 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=8.625 //y=7.4 //x2=8.88 //y2=7.4
r1764 (  233 914 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.45 //y=7.4 //x2=9.62 //y2=7.4
r1765 (  233 236 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.45 //y=7.4 //x2=8.88 //y2=7.4
r1766 (  227 913 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.54 //y=7.23 //x2=8.54 //y2=7.4
r1767 (  227 1014 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.54 //y=7.23 //x2=8.54 //y2=6.745
r1768 (  224 912 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.745 //y=7.4 //x2=7.66 //y2=7.4
r1769 (  224 226 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=7.745 //y=7.4 //x2=7.77 //y2=7.4
r1770 (  223 913 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.455 //y=7.4 //x2=8.54 //y2=7.4
r1771 (  223 226 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=8.455 //y=7.4 //x2=7.77 //y2=7.4
r1772 (  217 912 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.66 //y=7.23 //x2=7.66 //y2=7.4
r1773 (  217 1013 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.66 //y=7.23 //x2=7.66 //y2=6.745
r1774 (  216 911 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.865 //y=7.4 //x2=6.78 //y2=7.4
r1775 (  215 912 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.575 //y=7.4 //x2=7.66 //y2=7.4
r1776 (  215 216 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.575 //y=7.4 //x2=6.865 //y2=7.4
r1777 (  209 911 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=7.4
r1778 (  209 1012 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=6.745
r1779 (  206 910 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.985 //y=7.4 //x2=5.9 //y2=7.4
r1780 (  206 208 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=5.985 //y=7.4 //x2=6.66 //y2=7.4
r1781 (  205 911 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.78 //y2=7.4
r1782 (  205 208 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.66 //y2=7.4
r1783 (  199 910 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.9 //y=7.23 //x2=5.9 //y2=7.4
r1784 (  199 1011 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=5.9 //y=7.23 //x2=5.9 //y2=6.405
r1785 (  196 909 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=4.81 //y2=7.4
r1786 (  196 198 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=5.55 //y2=7.4
r1787 (  195 910 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.815 //y=7.4 //x2=5.9 //y2=7.4
r1788 (  195 198 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=5.815 //y=7.4 //x2=5.55 //y2=7.4
r1789 (  190 908 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=3.73 //y2=7.4
r1790 (  190 192 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=4.07 //y2=7.4
r1791 (  189 909 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.81 //y2=7.4
r1792 (  189 192 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.07 //y2=7.4
r1793 (  183 908 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=7.4
r1794 (  183 1010 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=6.745
r1795 (  180 907 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.85 //y2=7.4
r1796 (  180 182 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.96 //y2=7.4
r1797 (  179 908 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=3.73 //y2=7.4
r1798 (  179 182 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=2.96 //y2=7.4
r1799 (  173 907 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=7.4
r1800 (  173 1009 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=6.745
r1801 (  172 906 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.055 //y=7.4 //x2=1.97 //y2=7.4
r1802 (  171 907 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.85 //y2=7.4
r1803 (  171 172 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.055 //y2=7.4
r1804 (  165 906 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=7.4
r1805 (  165 1008 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=6.745
r1806 (  162 905 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.09 //y2=7.4
r1807 (  162 164 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.85 //y2=7.4
r1808 (  161 906 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.97 //y2=7.4
r1809 (  161 164 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.85 //y2=7.4
r1810 (  155 905 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=7.4
r1811 (  155 1007 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=6.405
r1812 (  151 905 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=1.09 //y2=7.4
r1813 (  151 154 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=0.74 //y2=7.4
r1814 (  147 902 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=86.95 //y=7.4 //x2=86.95 //y2=7.4
r1815 (  145 900 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=85.84 //y=7.4 //x2=85.84 //y2=7.4
r1816 (  145 147 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=85.84 //y=7.4 //x2=86.95 //y2=7.4
r1817 (  143 898 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=84.73 //y=7.4 //x2=84.73 //y2=7.4
r1818 (  143 145 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=84.73 //y=7.4 //x2=85.84 //y2=7.4
r1819 (  141 892 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=83.25 //y=7.4 //x2=83.25 //y2=7.4
r1820 (  141 143 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=83.25 //y=7.4 //x2=84.73 //y2=7.4
r1821 (  139 890 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=82.14 //y=7.4 //x2=82.14 //y2=7.4
r1822 (  139 141 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=82.14 //y=7.4 //x2=83.25 //y2=7.4
r1823 (  137 884 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=80.66 //y=7.4 //x2=80.66 //y2=7.4
r1824 (  137 139 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=80.66 //y=7.4 //x2=82.14 //y2=7.4
r1825 (  135 874 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=79.55 //y=7.4 //x2=79.55 //y2=7.4
r1826 (  135 137 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=79.55 //y=7.4 //x2=80.66 //y2=7.4
r1827 (  133 1002 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=78.44 //y=7.4 //x2=78.44 //y2=7.4
r1828 (  133 135 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=78.44 //y=7.4 //x2=79.55 //y2=7.4
r1829 (  131 999 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=76.96 //y=7.4 //x2=76.96 //y2=7.4
r1830 (  131 133 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=76.96 //y=7.4 //x2=78.44 //y2=7.4
r1831 (  129 836 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=75.85 //y=7.4 //x2=75.85 //y2=7.4
r1832 (  129 131 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=75.85 //y=7.4 //x2=76.96 //y2=7.4
r1833 (  127 826 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=74.74 //y=7.4 //x2=74.74 //y2=7.4
r1834 (  127 129 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=74.74 //y=7.4 //x2=75.85 //y2=7.4
r1835 (  125 994 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=73.26 //y=7.4 //x2=73.26 //y2=7.4
r1836 (  125 127 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=73.26 //y=7.4 //x2=74.74 //y2=7.4
r1837 (  123 804 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=72.15 //y=7.4 //x2=72.15 //y2=7.4
r1838 (  123 125 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=72.15 //y=7.4 //x2=73.26 //y2=7.4
r1839 (  121 794 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=71.04 //y=7.4 //x2=71.04 //y2=7.4
r1840 (  121 123 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=71.04 //y=7.4 //x2=72.15 //y2=7.4
r1841 (  119 784 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=69.93 //y=7.4 //x2=69.93 //y2=7.4
r1842 (  119 121 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=69.93 //y=7.4 //x2=71.04 //y2=7.4
r1843 (  117 988 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=68.45 //y=7.4 //x2=68.45 //y2=7.4
r1844 (  117 119 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=68.45 //y=7.4 //x2=69.93 //y2=7.4
r1845 (  115 762 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=67.34 //y=7.4 //x2=67.34 //y2=7.4
r1846 (  115 117 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=67.34 //y=7.4 //x2=68.45 //y2=7.4
r1847 (  113 752 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=66.23 //y=7.4 //x2=66.23 //y2=7.4
r1848 (  113 115 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=66.23 //y=7.4 //x2=67.34 //y2=7.4
r1849 (  111 742 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=65.12 //y=7.4 //x2=65.12 //y2=7.4
r1850 (  111 113 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=65.12 //y=7.4 //x2=66.23 //y2=7.4
r1851 (  109 728 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=63.64 //y=7.4 //x2=63.64 //y2=7.4
r1852 (  109 111 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=63.64 //y=7.4 //x2=65.12 //y2=7.4
r1853 (  107 718 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=62.53 //y=7.4 //x2=62.53 //y2=7.4
r1854 (  107 109 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=62.53 //y=7.4 //x2=63.64 //y2=7.4
r1855 (  105 704 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=61.05 //y=7.4 //x2=61.05 //y2=7.4
r1856 (  105 107 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=61.05 //y=7.4 //x2=62.53 //y2=7.4
r1857 (  103 694 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=59.94 //y=7.4 //x2=59.94 //y2=7.4
r1858 (  103 105 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=59.94 //y=7.4 //x2=61.05 //y2=7.4
r1859 (  101 684 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=58.83 //y=7.4 //x2=58.83 //y2=7.4
r1860 (  101 103 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=58.83 //y=7.4 //x2=59.94 //y2=7.4
r1861 (  99 975 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=57.72 //y=7.4 //x2=57.72 //y2=7.4
r1862 (  99 101 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=57.72 //y=7.4 //x2=58.83 //y2=7.4
r1863 (  97 662 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=56.24 //y=7.4 //x2=56.24 //y2=7.4
r1864 (  97 99 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=56.24 //y=7.4 //x2=57.72 //y2=7.4
r1865 (  95 652 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=55.13 //y=7.4 //x2=55.13 //y2=7.4
r1866 (  95 97 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=55.13 //y=7.4 //x2=56.24 //y2=7.4
r1867 (  93 642 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=54.02 //y=7.4 //x2=54.02 //y2=7.4
r1868 (  93 95 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=54.02 //y=7.4 //x2=55.13 //y2=7.4
r1869 (  91 969 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=52.91 //y=7.4 //x2=52.91 //y2=7.4
r1870 (  91 93 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=52.91 //y=7.4 //x2=54.02 //y2=7.4
r1871 (  89 620 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=51.43 //y=7.4 //x2=51.43 //y2=7.4
r1872 (  89 91 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=51.43 //y=7.4 //x2=52.91 //y2=7.4
r1873 (  87 610 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=50.32 //y=7.4 //x2=50.32 //y2=7.4
r1874 (  87 89 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=50.32 //y=7.4 //x2=51.43 //y2=7.4
r1875 (  85 964 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=49.21 //y=7.4 //x2=49.21 //y2=7.4
r1876 (  85 87 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=49.21 //y=7.4 //x2=50.32 //y2=7.4
r1877 (  83 588 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=47.73 //y=7.4 //x2=47.73 //y2=7.4
r1878 (  83 85 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=47.73 //y=7.4 //x2=49.21 //y2=7.4
r1879 (  81 578 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=46.62 //y=7.4 //x2=46.62 //y2=7.4
r1880 (  81 83 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=46.62 //y=7.4 //x2=47.73 //y2=7.4
r1881 (  79 560 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=45.51 //y=7.4 //x2=45.51 //y2=7.4
r1882 (  79 81 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=45.51 //y=7.4 //x2=46.62 //y2=7.4
r1883 (  77 550 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=44.4 //y=7.4 //x2=44.4 //y2=7.4
r1884 (  77 79 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=44.4 //y=7.4 //x2=45.51 //y2=7.4
r1885 (  74 544 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=42.92 //y=7.4 //x2=42.92 //y2=7.4
r1886 (  72 534 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=41.81 //y=7.4 //x2=41.81 //y2=7.4
r1887 (  72 74 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=41.81 //y=7.4 //x2=42.92 //y2=7.4
r1888 (  70 516 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=40.7 //y=7.4 //x2=40.7 //y2=7.4
r1889 (  70 72 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=40.7 //y=7.4 //x2=41.81 //y2=7.4
r1890 (  68 506 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=39.59 //y=7.4 //x2=39.59 //y2=7.4
r1891 (  68 70 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=39.59 //y=7.4 //x2=40.7 //y2=7.4
r1892 (  66 951 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=38.11 //y=7.4 //x2=38.11 //y2=7.4
r1893 (  66 68 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=38.11 //y=7.4 //x2=39.59 //y2=7.4
r1894 (  64 484 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37 //y=7.4 //x2=37 //y2=7.4
r1895 (  64 66 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=37 //y=7.4 //x2=38.11 //y2=7.4
r1896 (  62 474 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.89 //y=7.4 //x2=35.89 //y2=7.4
r1897 (  62 64 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=35.89 //y=7.4 //x2=37 //y2=7.4
r1898 (  60 946 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.41 //y=7.4 //x2=34.41 //y2=7.4
r1899 (  60 62 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=34.41 //y=7.4 //x2=35.89 //y2=7.4
r1900 (  58 452 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=33.3 //y=7.4 //x2=33.3 //y2=7.4
r1901 (  58 60 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=33.3 //y=7.4 //x2=34.41 //y2=7.4
r1902 (  56 442 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.19 //y=7.4 //x2=32.19 //y2=7.4
r1903 (  56 58 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=32.19 //y=7.4 //x2=33.3 //y2=7.4
r1904 (  54 432 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.08 //y=7.4 //x2=31.08 //y2=7.4
r1905 (  54 56 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.08 //y=7.4 //x2=32.19 //y2=7.4
r1906 (  52 940 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=29.6 //y=7.4 //x2=29.6 //y2=7.4
r1907 (  52 54 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=29.6 //y=7.4 //x2=31.08 //y2=7.4
r1908 (  50 410 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.49 //y=7.4 //x2=28.49 //y2=7.4
r1909 (  50 52 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=28.49 //y=7.4 //x2=29.6 //y2=7.4
r1910 (  48 400 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.38 //y=7.4 //x2=27.38 //y2=7.4
r1911 (  48 50 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=27.38 //y=7.4 //x2=28.49 //y2=7.4
r1912 (  46 390 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=26.27 //y=7.4 //x2=26.27 //y2=7.4
r1913 (  46 48 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=26.27 //y=7.4 //x2=27.38 //y2=7.4
r1914 (  44 376 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=7.4 //x2=24.79 //y2=7.4
r1915 (  44 46 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=7.4 //x2=26.27 //y2=7.4
r1916 (  42 366 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=7.4 //x2=23.68 //y2=7.4
r1917 (  42 44 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=23.68 //y=7.4 //x2=24.79 //y2=7.4
r1918 (  40 352 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.2 //y=7.4 //x2=22.2 //y2=7.4
r1919 (  40 42 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=22.2 //y=7.4 //x2=23.68 //y2=7.4
r1920 (  38 342 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=7.4 //x2=21.09 //y2=7.4
r1921 (  38 40 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=7.4 //x2=22.2 //y2=7.4
r1922 (  36 332 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=7.4 //x2=19.98 //y2=7.4
r1923 (  36 38 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=7.4 //x2=21.09 //y2=7.4
r1924 (  34 927 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.87 //y=7.4 //x2=18.87 //y2=7.4
r1925 (  34 36 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=18.87 //y=7.4 //x2=19.98 //y2=7.4
r1926 (  32 310 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=7.4 //x2=17.39 //y2=7.4
r1927 (  32 34 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=7.4 //x2=18.87 //y2=7.4
r1928 (  30 300 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=7.4 //x2=16.28 //y2=7.4
r1929 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=7.4 //x2=17.39 //y2=7.4
r1930 (  28 290 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=7.4 //x2=15.17 //y2=7.4
r1931 (  28 30 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=7.4 //x2=16.28 //y2=7.4
r1932 (  26 921 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=7.4 //x2=14.06 //y2=7.4
r1933 (  26 28 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=7.4 //x2=15.17 //y2=7.4
r1934 (  24 268 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=7.4 //x2=12.58 //y2=7.4
r1935 (  24 26 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=7.4 //x2=14.06 //y2=7.4
r1936 (  22 258 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=7.4 //x2=11.47 //y2=7.4
r1937 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=7.4 //x2=12.58 //y2=7.4
r1938 (  20 916 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r1939 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=7.4 //x2=11.47 //y2=7.4
r1940 (  18 236 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.88 //y=7.4 //x2=8.88 //y2=7.4
r1941 (  18 20 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.88 //y=7.4 //x2=10.36 //y2=7.4
r1942 (  16 226 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=7.4 //x2=7.77 //y2=7.4
r1943 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=7.4 //x2=8.88 //y2=7.4
r1944 (  14 208 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r1945 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.4 //x2=7.77 //y2=7.4
r1946 (  12 198 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r1947 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.66 //y2=7.4
r1948 (  10 192 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=7.4 //x2=4.07 //y2=7.4
r1949 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=7.4 //x2=5.55 //y2=7.4
r1950 (  8 182 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r1951 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r1952 (  6 164 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r1953 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r1954 (  3 154 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r1955 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r1956 (  1 77 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=43.845 //y=7.4 //x2=44.4 //y2=7.4
r1957 (  1 74 ) resistor r=0.384136 //w=0.301 //l=0.925 //layer=m1 \
 //thickness=0.36 //x=43.845 //y=7.4 //x2=42.92 //y2=7.4
ends PM_TMRDFFRNQNX1\%VDD

subckt PM_TMRDFFRNQNX1\%noxref_3 ( 1 2 3 4 12 25 26 33 41 47 48 52 54 61 62 63 \
 64 65 66 67 68 72 73 74 79 81 84 85 86 87 88 89 93 95 98 99 104 105 110 119 \
 122 124 125 126 )
c250 ( 126 0 ) capacitor c=0.023087f //x=7.955 //y=5.02
c251 ( 125 0 ) capacitor c=0.023519f //x=7.075 //y=5.02
c252 ( 124 0 ) capacitor c=0.0224735f //x=6.195 //y=5.02
c253 ( 122 0 ) capacitor c=0.00872971f //x=8.205 //y=0.915
c254 ( 119 0 ) capacitor c=0.0588816f //x=10.73 //y=4.7
c255 ( 110 0 ) capacitor c=0.058931f //x=3.33 //y=4.7
c256 ( 105 0 ) capacitor c=0.0273931f //x=3.33 //y=1.915
c257 ( 104 0 ) capacitor c=0.0464411f //x=3.33 //y=2.08
c258 ( 99 0 ) capacitor c=0.0318948f //x=11.065 //y=1.21
c259 ( 98 0 ) capacitor c=0.0187384f //x=11.065 //y=0.865
c260 ( 95 0 ) capacitor c=0.0141798f //x=10.91 //y=1.365
c261 ( 93 0 ) capacitor c=0.0149844f //x=10.91 //y=0.71
c262 ( 89 0 ) capacitor c=0.0813322f //x=10.535 //y=1.915
c263 ( 88 0 ) capacitor c=0.0229267f //x=10.535 //y=1.52
c264 ( 87 0 ) capacitor c=0.0234352f //x=10.535 //y=1.21
c265 ( 86 0 ) capacitor c=0.0199343f //x=10.535 //y=0.865
c266 ( 85 0 ) capacitor c=0.0432517f //x=3.85 //y=1.26
c267 ( 84 0 ) capacitor c=0.0200379f //x=3.85 //y=0.915
c268 ( 81 0 ) capacitor c=0.0158629f //x=3.695 //y=1.415
c269 ( 79 0 ) capacitor c=0.0157803f //x=3.695 //y=0.76
c270 ( 74 0 ) capacitor c=0.0218028f //x=3.32 //y=1.57
c271 ( 73 0 ) capacitor c=0.0207459f //x=3.32 //y=1.26
c272 ( 72 0 ) capacitor c=0.0194308f //x=3.32 //y=0.915
c273 ( 68 0 ) capacitor c=0.110275f //x=11.07 //y=6.02
c274 ( 67 0 ) capacitor c=0.154305f //x=10.63 //y=6.02
c275 ( 66 0 ) capacitor c=0.158794f //x=3.51 //y=6.02
c276 ( 65 0 ) capacitor c=0.110114f //x=3.07 //y=6.02
c277 ( 62 0 ) capacitor c=0.00106608f //x=8.1 //y=5.155
c278 ( 61 0 ) capacitor c=0.00207319f //x=7.22 //y=5.155
c279 ( 54 0 ) capacitor c=0.0872487f //x=10.73 //y=2.08
c280 ( 52 0 ) capacitor c=0.10679f //x=8.88 //y=3.33
c281 ( 48 0 ) capacitor c=0.00398962f //x=8.48 //y=1.665
c282 ( 47 0 ) capacitor c=0.0137288f //x=8.795 //y=1.665
c283 ( 41 0 ) capacitor c=0.0284988f //x=8.795 //y=5.155
c284 ( 33 0 ) capacitor c=0.0176454f //x=8.015 //y=5.155
c285 ( 26 0 ) capacitor c=0.00332903f //x=6.425 //y=5.155
c286 ( 25 0 ) capacitor c=0.0148427f //x=7.135 //y=5.155
c287 ( 12 0 ) capacitor c=0.0883349f //x=3.33 //y=2.08
c288 ( 4 0 ) capacitor c=0.00455264f //x=8.995 //y=3.33
c289 ( 3 0 ) capacitor c=0.0402401f //x=10.615 //y=3.33
c290 ( 2 0 ) capacitor c=0.0164246f //x=3.445 //y=3.33
c291 ( 1 0 ) capacitor c=0.130412f //x=8.765 //y=3.33
r292 (  117 119 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=10.63 //y=4.7 //x2=10.73 //y2=4.7
r293 (  104 105 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.33 //y=2.08 //x2=3.33 //y2=1.915
r294 (  100 119 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=11.07 //y=4.865 //x2=10.73 //y2=4.7
r295 (  99 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.065 //y=1.21 //x2=11.025 //y2=1.365
r296 (  98 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.065 //y=0.865 //x2=11.025 //y2=0.71
r297 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.065 //y=0.865 //x2=11.065 //y2=1.21
r298 (  96 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.69 //y=1.365 //x2=10.575 //y2=1.365
r299 (  95 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.91 //y=1.365 //x2=11.025 //y2=1.365
r300 (  94 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.69 //y=0.71 //x2=10.575 //y2=0.71
r301 (  93 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.91 //y=0.71 //x2=11.025 //y2=0.71
r302 (  93 94 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.91 //y=0.71 //x2=10.69 //y2=0.71
r303 (  90 117 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=10.63 //y=4.865 //x2=10.63 //y2=4.7
r304 (  89 114 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=10.535 //y=1.915 //x2=10.73 //y2=2.08
r305 (  88 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.535 //y=1.52 //x2=10.575 //y2=1.365
r306 (  88 89 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=10.535 //y=1.52 //x2=10.535 //y2=1.915
r307 (  87 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.535 //y=1.21 //x2=10.575 //y2=1.365
r308 (  86 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.535 //y=0.865 //x2=10.575 //y2=0.71
r309 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.535 //y=0.865 //x2=10.535 //y2=1.21
r310 (  85 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=1.26 //x2=3.81 //y2=1.415
r311 (  84 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.81 //y2=0.76
r312 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.85 //y2=1.26
r313 (  82 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=1.415 //x2=3.36 //y2=1.415
r314 (  81 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=1.415 //x2=3.81 //y2=1.415
r315 (  80 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=0.76 //x2=3.36 //y2=0.76
r316 (  79 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.81 //y2=0.76
r317 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.475 //y2=0.76
r318 (  76 110 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=3.51 //y=4.865 //x2=3.33 //y2=4.7
r319 (  74 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.36 //y2=1.415
r320 (  74 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.32 //y2=1.915
r321 (  73 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.26 //x2=3.36 //y2=1.415
r322 (  72 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.36 //y2=0.76
r323 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.32 //y2=1.26
r324 (  69 110 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=3.07 //y=4.865 //x2=3.33 //y2=4.7
r325 (  68 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.07 //y=6.02 //x2=11.07 //y2=4.865
r326 (  67 90 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.63 //y=6.02 //x2=10.63 //y2=4.865
r327 (  66 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.51 //y=6.02 //x2=3.51 //y2=4.865
r328 (  65 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.07 //y=6.02 //x2=3.07 //y2=4.865
r329 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.8 //y=1.365 //x2=10.91 //y2=1.365
r330 (  64 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.8 //y=1.365 //x2=10.69 //y2=1.365
r331 (  63 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.695 //y2=1.415
r332 (  63 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.475 //y2=1.415
r333 (  59 119 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=4.7 //x2=10.73 //y2=4.7
r334 (  57 59 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=10.73 //y=3.33 //x2=10.73 //y2=4.7
r335 (  54 114 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=2.08 //x2=10.73 //y2=2.08
r336 (  54 57 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.08 //x2=10.73 //y2=3.33
r337 (  50 52 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=8.88 //y=5.07 //x2=8.88 //y2=3.33
r338 (  49 52 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=8.88 //y=1.75 //x2=8.88 //y2=3.33
r339 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.795 //y=1.665 //x2=8.88 //y2=1.75
r340 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=8.795 //y=1.665 //x2=8.48 //y2=1.665
r341 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.395 //y=1.58 //x2=8.48 //y2=1.665
r342 (  43 122 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=8.395 //y=1.58 //x2=8.395 //y2=1.01
r343 (  42 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.185 //y=5.155 //x2=8.1 //y2=5.155
r344 (  41 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.795 //y=5.155 //x2=8.88 //y2=5.07
r345 (  41 42 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=8.795 //y=5.155 //x2=8.185 //y2=5.155
r346 (  35 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.1 //y=5.24 //x2=8.1 //y2=5.155
r347 (  35 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.1 //y=5.24 //x2=8.1 //y2=5.725
r348 (  34 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.305 //y=5.155 //x2=7.22 //y2=5.155
r349 (  33 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.015 //y=5.155 //x2=8.1 //y2=5.155
r350 (  33 34 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.015 //y=5.155 //x2=7.305 //y2=5.155
r351 (  27 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.24 //x2=7.22 //y2=5.155
r352 (  27 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.24 //x2=7.22 //y2=5.725
r353 (  25 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.155 //x2=7.22 //y2=5.155
r354 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.155 //x2=6.425 //y2=5.155
r355 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.24 //x2=6.425 //y2=5.155
r356 (  19 124 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.24 //x2=6.34 //y2=5.725
r357 (  17 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r358 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=3.33 //x2=3.33 //y2=4.7
r359 (  12 104 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r360 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.08 //x2=3.33 //y2=3.33
r361 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.73 //y=3.33 //x2=10.73 //y2=3.33
r362 (  8 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.88 //y=3.33 //x2=8.88 //y2=3.33
r363 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=3.33 //x2=3.33 //y2=3.33
r364 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.995 //y=3.33 //x2=8.88 //y2=3.33
r365 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=3.33 //x2=10.73 //y2=3.33
r366 (  3 4 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=10.615 //y=3.33 //x2=8.995 //y2=3.33
r367 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.445 //y=3.33 //x2=3.33 //y2=3.33
r368 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=3.33 //x2=8.88 //y2=3.33
r369 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=3.33 //x2=3.445 //y2=3.33
ends PM_TMRDFFRNQNX1\%noxref_3

subckt PM_TMRDFFRNQNX1\%noxref_4 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 \
 47 48 49 51 57 58 59 60 72 74 75 )
c152 ( 75 0 ) capacitor c=0.0220291f //x=11.585 //y=5.02
c153 ( 74 0 ) capacitor c=0.0217503f //x=10.705 //y=5.02
c154 ( 72 0 ) capacitor c=0.0084702f //x=11.58 //y=0.905
c155 ( 60 0 ) capacitor c=0.0557698f //x=14.335 //y=4.79
c156 ( 59 0 ) capacitor c=0.0293157f //x=14.625 //y=4.79
c157 ( 58 0 ) capacitor c=0.0347816f //x=14.29 //y=1.22
c158 ( 57 0 ) capacitor c=0.0187487f //x=14.29 //y=0.875
c159 ( 51 0 ) capacitor c=0.0137055f //x=14.135 //y=1.375
c160 ( 49 0 ) capacitor c=0.0149861f //x=14.135 //y=0.72
c161 ( 48 0 ) capacitor c=0.096037f //x=13.76 //y=1.915
c162 ( 47 0 ) capacitor c=0.0228993f //x=13.76 //y=1.53
c163 ( 46 0 ) capacitor c=0.0234352f //x=13.76 //y=1.22
c164 ( 45 0 ) capacitor c=0.0198724f //x=13.76 //y=0.875
c165 ( 44 0 ) capacitor c=0.110114f //x=14.7 //y=6.02
c166 ( 43 0 ) capacitor c=0.158956f //x=14.26 //y=6.02
c167 ( 41 0 ) capacitor c=0.00211606f //x=11.73 //y=5.2
c168 ( 34 0 ) capacitor c=0.0970289f //x=14.06 //y=2.08
c169 ( 32 0 ) capacitor c=0.105815f //x=12.21 //y=3.33
c170 ( 28 0 ) capacitor c=0.00404073f //x=11.855 //y=1.655
c171 ( 27 0 ) capacitor c=0.0122201f //x=12.125 //y=1.655
c172 ( 25 0 ) capacitor c=0.0137995f //x=12.125 //y=5.2
c173 ( 14 0 ) capacitor c=0.00251635f //x=10.935 //y=5.2
c174 ( 13 0 ) capacitor c=0.0143649f //x=11.645 //y=5.2
c175 ( 2 0 ) capacitor c=0.00703116f //x=12.325 //y=3.33
c176 ( 1 0 ) capacitor c=0.0456992f //x=13.945 //y=3.33
r177 (  59 61 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=14.625 //y=4.79 //x2=14.7 //y2=4.865
r178 (  59 60 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=14.625 //y=4.79 //x2=14.335 //y2=4.79
r179 (  58 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.29 //y=1.22 //x2=14.25 //y2=1.375
r180 (  57 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.29 //y=0.875 //x2=14.25 //y2=0.72
r181 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.29 //y=0.875 //x2=14.29 //y2=1.22
r182 (  54 60 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=14.26 //y=4.865 //x2=14.335 //y2=4.79
r183 (  54 69 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=14.26 //y=4.865 //x2=14.06 //y2=4.7
r184 (  52 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.915 //y=1.375 //x2=13.8 //y2=1.375
r185 (  51 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.135 //y=1.375 //x2=14.25 //y2=1.375
r186 (  50 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.915 //y=0.72 //x2=13.8 //y2=0.72
r187 (  49 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.135 //y=0.72 //x2=14.25 //y2=0.72
r188 (  49 50 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=14.135 //y=0.72 //x2=13.915 //y2=0.72
r189 (  48 67 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=13.76 //y=1.915 //x2=14.06 //y2=2.08
r190 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.76 //y=1.53 //x2=13.8 //y2=1.375
r191 (  47 48 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=13.76 //y=1.53 //x2=13.76 //y2=1.915
r192 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.76 //y=1.22 //x2=13.8 //y2=1.375
r193 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.76 //y=0.875 //x2=13.8 //y2=0.72
r194 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.76 //y=0.875 //x2=13.76 //y2=1.22
r195 (  44 61 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.7 //y=6.02 //x2=14.7 //y2=4.865
r196 (  43 54 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.26 //y=6.02 //x2=14.26 //y2=4.865
r197 (  42 51 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.025 //y=1.375 //x2=14.135 //y2=1.375
r198 (  42 52 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.025 //y=1.375 //x2=13.915 //y2=1.375
r199 (  39 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=4.7 //x2=14.06 //y2=4.7
r200 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=14.06 //y=3.33 //x2=14.06 //y2=4.7
r201 (  34 67 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=2.08 //x2=14.06 //y2=2.08
r202 (  34 37 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=14.06 //y=2.08 //x2=14.06 //y2=3.33
r203 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=12.21 //y=5.115 //x2=12.21 //y2=3.33
r204 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=12.21 //y=1.74 //x2=12.21 //y2=3.33
r205 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.125 //y=1.655 //x2=12.21 //y2=1.74
r206 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=12.125 //y=1.655 //x2=11.855 //y2=1.655
r207 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.815 //y=5.2 //x2=11.73 //y2=5.2
r208 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.125 //y=5.2 //x2=12.21 //y2=5.115
r209 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=12.125 //y=5.2 //x2=11.815 //y2=5.2
r210 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.77 //y=1.57 //x2=11.855 //y2=1.655
r211 (  21 72 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=11.77 //y=1.57 //x2=11.77 //y2=1
r212 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.73 //y=5.285 //x2=11.73 //y2=5.2
r213 (  15 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=11.73 //y=5.285 //x2=11.73 //y2=5.725
r214 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.645 //y=5.2 //x2=11.73 //y2=5.2
r215 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.645 //y=5.2 //x2=10.935 //y2=5.2
r216 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.85 //y=5.285 //x2=10.935 //y2=5.2
r217 (  7 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=10.85 //y=5.285 //x2=10.85 //y2=5.725
r218 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.06 //y=3.33 //x2=14.06 //y2=3.33
r219 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.21 //y=3.33 //x2=12.21 //y2=3.33
r220 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.325 //y=3.33 //x2=12.21 //y2=3.33
r221 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=3.33 //x2=14.06 //y2=3.33
r222 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=13.945 //y=3.33 //x2=12.325 //y2=3.33
ends PM_TMRDFFRNQNX1\%noxref_4

subckt PM_TMRDFFRNQNX1\%noxref_5 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 63 \
 64 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 92 94 100 101 102 \
 103 123 125 126 127 )
c253 ( 127 0 ) capacitor c=0.023087f //x=3.145 //y=5.02
c254 ( 126 0 ) capacitor c=0.023519f //x=2.265 //y=5.02
c255 ( 125 0 ) capacitor c=0.0224735f //x=1.385 //y=5.02
c256 ( 123 0 ) capacitor c=0.00853354f //x=3.395 //y=0.915
c257 ( 103 0 ) capacitor c=0.0556143f //x=19.145 //y=4.79
c258 ( 102 0 ) capacitor c=0.0293157f //x=19.435 //y=4.79
c259 ( 101 0 ) capacitor c=0.0347816f //x=19.1 //y=1.22
c260 ( 100 0 ) capacitor c=0.0187487f //x=19.1 //y=0.875
c261 ( 94 0 ) capacitor c=0.0137055f //x=18.945 //y=1.375
c262 ( 92 0 ) capacitor c=0.0149861f //x=18.945 //y=0.72
c263 ( 91 0 ) capacitor c=0.096037f //x=18.57 //y=1.915
c264 ( 90 0 ) capacitor c=0.0228993f //x=18.57 //y=1.53
c265 ( 89 0 ) capacitor c=0.0234352f //x=18.57 //y=1.22
c266 ( 88 0 ) capacitor c=0.0198724f //x=18.57 //y=0.875
c267 ( 84 0 ) capacitor c=0.0556143f //x=6.195 //y=4.79
c268 ( 83 0 ) capacitor c=0.0293157f //x=6.485 //y=4.79
c269 ( 82 0 ) capacitor c=0.0347816f //x=6.15 //y=1.22
c270 ( 81 0 ) capacitor c=0.0187487f //x=6.15 //y=0.875
c271 ( 75 0 ) capacitor c=0.0137055f //x=5.995 //y=1.375
c272 ( 73 0 ) capacitor c=0.0149861f //x=5.995 //y=0.72
c273 ( 72 0 ) capacitor c=0.102158f //x=5.62 //y=1.915
c274 ( 71 0 ) capacitor c=0.0229444f //x=5.62 //y=1.53
c275 ( 70 0 ) capacitor c=0.0234352f //x=5.62 //y=1.22
c276 ( 69 0 ) capacitor c=0.0198724f //x=5.62 //y=0.875
c277 ( 68 0 ) capacitor c=0.110114f //x=19.51 //y=6.02
c278 ( 67 0 ) capacitor c=0.158956f //x=19.07 //y=6.02
c279 ( 66 0 ) capacitor c=0.110114f //x=6.56 //y=6.02
c280 ( 65 0 ) capacitor c=0.158956f //x=6.12 //y=6.02
c281 ( 62 0 ) capacitor c=0.00106608f //x=3.29 //y=5.155
c282 ( 61 0 ) capacitor c=0.00207162f //x=2.41 //y=5.155
c283 ( 54 0 ) capacitor c=0.100095f //x=18.87 //y=2.08
c284 ( 46 0 ) capacitor c=0.101432f //x=5.92 //y=2.08
c285 ( 44 0 ) capacitor c=0.109588f //x=4.07 //y=3.7
c286 ( 40 0 ) capacitor c=0.00493499f //x=3.67 //y=1.665
c287 ( 39 0 ) capacitor c=0.0154052f //x=3.985 //y=1.665
c288 ( 33 0 ) capacitor c=0.0283082f //x=3.985 //y=5.155
c289 ( 25 0 ) capacitor c=0.0176454f //x=3.205 //y=5.155
c290 ( 18 0 ) capacitor c=0.00351598f //x=1.615 //y=5.155
c291 ( 17 0 ) capacitor c=0.0154196f //x=2.325 //y=5.155
c292 ( 4 0 ) capacitor c=0.00424246f //x=6.035 //y=3.7
c293 ( 3 0 ) capacitor c=0.229463f //x=18.755 //y=3.7
c294 ( 2 0 ) capacitor c=0.0125346f //x=4.185 //y=3.7
c295 ( 1 0 ) capacitor c=0.0288301f //x=5.805 //y=3.7
r296 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=19.435 //y=4.79 //x2=19.51 //y2=4.865
r297 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=19.435 //y=4.79 //x2=19.145 //y2=4.79
r298 (  101 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.1 //y=1.22 //x2=19.06 //y2=1.375
r299 (  100 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.1 //y=0.875 //x2=19.06 //y2=0.72
r300 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=19.1 //y=0.875 //x2=19.1 //y2=1.22
r301 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=19.07 //y=4.865 //x2=19.145 //y2=4.79
r302 (  97 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=19.07 //y=4.865 //x2=18.87 //y2=4.7
r303 (  95 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.725 //y=1.375 //x2=18.61 //y2=1.375
r304 (  94 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.945 //y=1.375 //x2=19.06 //y2=1.375
r305 (  93 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.725 //y=0.72 //x2=18.61 //y2=0.72
r306 (  92 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.945 //y=0.72 //x2=19.06 //y2=0.72
r307 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=18.945 //y=0.72 //x2=18.725 //y2=0.72
r308 (  91 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=18.57 //y=1.915 //x2=18.87 //y2=2.08
r309 (  90 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.57 //y=1.53 //x2=18.61 //y2=1.375
r310 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=18.57 //y=1.53 //x2=18.57 //y2=1.915
r311 (  89 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.57 //y=1.22 //x2=18.61 //y2=1.375
r312 (  88 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.57 //y=0.875 //x2=18.61 //y2=0.72
r313 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.57 //y=0.875 //x2=18.57 //y2=1.22
r314 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.485 //y=4.79 //x2=6.56 //y2=4.865
r315 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=6.485 //y=4.79 //x2=6.195 //y2=4.79
r316 (  82 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.15 //y=1.22 //x2=6.11 //y2=1.375
r317 (  81 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.15 //y=0.875 //x2=6.11 //y2=0.72
r318 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.15 //y=0.875 //x2=6.15 //y2=1.22
r319 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.12 //y=4.865 //x2=6.195 //y2=4.79
r320 (  78 112 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=6.12 //y=4.865 //x2=5.92 //y2=4.7
r321 (  76 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.775 //y=1.375 //x2=5.66 //y2=1.375
r322 (  75 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.995 //y=1.375 //x2=6.11 //y2=1.375
r323 (  74 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.775 //y=0.72 //x2=5.66 //y2=0.72
r324 (  73 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.995 //y=0.72 //x2=6.11 //y2=0.72
r325 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=5.995 //y=0.72 //x2=5.775 //y2=0.72
r326 (  72 110 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.915 //x2=5.92 //y2=2.08
r327 (  71 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.53 //x2=5.66 //y2=1.375
r328 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.53 //x2=5.62 //y2=1.915
r329 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.22 //x2=5.66 //y2=1.375
r330 (  69 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=0.875 //x2=5.66 //y2=0.72
r331 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.62 //y=0.875 //x2=5.62 //y2=1.22
r332 (  68 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.51 //y=6.02 //x2=19.51 //y2=4.865
r333 (  67 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.07 //y=6.02 //x2=19.07 //y2=4.865
r334 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.56 //y=6.02 //x2=6.56 //y2=4.865
r335 (  65 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.12 //y=6.02 //x2=6.12 //y2=4.865
r336 (  64 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.835 //y=1.375 //x2=18.945 //y2=1.375
r337 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.835 //y=1.375 //x2=18.725 //y2=1.375
r338 (  63 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.375 //x2=5.995 //y2=1.375
r339 (  63 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.375 //x2=5.775 //y2=1.375
r340 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.87 //y=4.7 //x2=18.87 //y2=4.7
r341 (  57 59 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=18.87 //y=3.7 //x2=18.87 //y2=4.7
r342 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.87 //y=2.08 //x2=18.87 //y2=2.08
r343 (  54 57 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=18.87 //y=2.08 //x2=18.87 //y2=3.7
r344 (  51 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=4.7 //x2=5.92 //y2=4.7
r345 (  49 51 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=5.92 //y=3.7 //x2=5.92 //y2=4.7
r346 (  46 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=2.08 //x2=5.92 //y2=2.08
r347 (  46 49 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.08 //x2=5.92 //y2=3.7
r348 (  42 44 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=4.07 //y=5.07 //x2=4.07 //y2=3.7
r349 (  41 44 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=4.07 //y=1.75 //x2=4.07 //y2=3.7
r350 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=4.07 //y2=1.75
r351 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=3.67 //y2=1.665
r352 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.67 //y2=1.665
r353 (  35 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.585 //y2=1.01
r354 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.375 //y=5.155 //x2=3.29 //y2=5.155
r355 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=4.07 //y2=5.07
r356 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=3.375 //y2=5.155
r357 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.155
r358 (  27 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.725
r359 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.495 //y=5.155 //x2=2.41 //y2=5.155
r360 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=3.29 //y2=5.155
r361 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=2.495 //y2=5.155
r362 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.155
r363 (  19 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.725
r364 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=2.41 //y2=5.155
r365 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=1.615 //y2=5.155
r366 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.615 //y2=5.155
r367 (  11 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.53 //y2=5.725
r368 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.87 //y=3.7 //x2=18.87 //y2=3.7
r369 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.92 //y=3.7 //x2=5.92 //y2=3.7
r370 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=3.7 //x2=4.07 //y2=3.7
r371 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.035 //y=3.7 //x2=5.92 //y2=3.7
r372 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.755 //y=3.7 //x2=18.87 //y2=3.7
r373 (  3 4 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=18.755 //y=3.7 //x2=6.035 //y2=3.7
r374 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.185 //y=3.7 //x2=4.07 //y2=3.7
r375 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.805 //y=3.7 //x2=5.92 //y2=3.7
r376 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=5.805 //y=3.7 //x2=4.185 //y2=3.7
ends PM_TMRDFFRNQNX1\%noxref_5

subckt PM_TMRDFFRNQNX1\%noxref_6 ( 1 2 3 4 5 6 7 8 9 10 24 31 33 43 44 51 59 \
 65 66 70 77 78 85 93 99 100 104 106 113 115 121 122 123 124 127 128 129 130 \
 131 132 133 134 135 136 137 138 139 140 141 142 143 145 151 152 153 154 158 \
 159 160 165 167 169 175 176 177 178 179 180 184 186 189 190 194 195 196 201 \
 203 205 211 212 222 223 226 240 244 245 248 256 257 260 261 262 263 264 265 )
c485 ( 265 0 ) capacitor c=0.023087f //x=20.905 //y=5.02
c486 ( 264 0 ) capacitor c=0.023519f //x=20.025 //y=5.02
c487 ( 263 0 ) capacitor c=0.0224735f //x=19.145 //y=5.02
c488 ( 262 0 ) capacitor c=0.023087f //x=16.095 //y=5.02
c489 ( 261 0 ) capacitor c=0.023519f //x=15.215 //y=5.02
c490 ( 260 0 ) capacitor c=0.0224735f //x=14.335 //y=5.02
c491 ( 257 0 ) capacitor c=0.00872971f //x=21.155 //y=0.915
c492 ( 256 0 ) capacitor c=0.00853354f //x=16.345 //y=0.915
c493 ( 248 0 ) capacitor c=0.0339723f //x=24.45 //y=4.7
c494 ( 245 0 ) capacitor c=0.0292616f //x=24.42 //y=1.915
c495 ( 244 0 ) capacitor c=0.0430486f //x=24.42 //y=2.08
c496 ( 240 0 ) capacitor c=0.0598414f //x=23.68 //y=4.7
c497 ( 226 0 ) capacitor c=0.0331095f //x=11.5 //y=4.7
c498 ( 223 0 ) capacitor c=0.0279499f //x=11.47 //y=1.915
c499 ( 222 0 ) capacitor c=0.0421676f //x=11.47 //y=2.08
c500 ( 212 0 ) capacitor c=0.0431781f //x=24.985 //y=1.25
c501 ( 211 0 ) capacitor c=0.0197948f //x=24.985 //y=0.905
c502 ( 205 0 ) capacitor c=0.0148884f //x=24.83 //y=1.405
c503 ( 203 0 ) capacitor c=0.0157803f //x=24.83 //y=0.75
c504 ( 201 0 ) capacitor c=0.0295235f //x=24.825 //y=4.79
c505 ( 196 0 ) capacitor c=0.02098f //x=24.455 //y=1.56
c506 ( 195 0 ) capacitor c=0.0179879f //x=24.455 //y=1.25
c507 ( 194 0 ) capacitor c=0.0177928f //x=24.455 //y=0.905
c508 ( 190 0 ) capacitor c=0.0338875f //x=24.015 //y=1.21
c509 ( 189 0 ) capacitor c=0.0189263f //x=24.015 //y=0.865
c510 ( 186 0 ) capacitor c=0.0141798f //x=23.86 //y=1.365
c511 ( 184 0 ) capacitor c=0.0149844f //x=23.86 //y=0.71
c512 ( 180 0 ) capacitor c=0.0828193f //x=23.485 //y=1.915
c513 ( 179 0 ) capacitor c=0.0230657f //x=23.485 //y=1.52
c514 ( 178 0 ) capacitor c=0.0234352f //x=23.485 //y=1.21
c515 ( 177 0 ) capacitor c=0.0201338f //x=23.485 //y=0.865
c516 ( 176 0 ) capacitor c=0.0429696f //x=12.035 //y=1.25
c517 ( 175 0 ) capacitor c=0.0192208f //x=12.035 //y=0.905
c518 ( 169 0 ) capacitor c=0.0148884f //x=11.88 //y=1.405
c519 ( 167 0 ) capacitor c=0.0157803f //x=11.88 //y=0.75
c520 ( 165 0 ) capacitor c=0.0295235f //x=11.875 //y=4.79
c521 ( 160 0 ) capacitor c=0.0204188f //x=11.505 //y=1.56
c522 ( 159 0 ) capacitor c=0.0168481f //x=11.505 //y=1.25
c523 ( 158 0 ) capacitor c=0.0174783f //x=11.505 //y=0.905
c524 ( 154 0 ) capacitor c=0.0559896f //x=1.385 //y=4.79
c525 ( 153 0 ) capacitor c=0.0298189f //x=1.675 //y=4.79
c526 ( 152 0 ) capacitor c=0.0347816f //x=1.34 //y=1.22
c527 ( 151 0 ) capacitor c=0.0187487f //x=1.34 //y=0.875
c528 ( 145 0 ) capacitor c=0.0137055f //x=1.185 //y=1.375
c529 ( 143 0 ) capacitor c=0.0149861f //x=1.185 //y=0.72
c530 ( 142 0 ) capacitor c=0.102158f //x=0.81 //y=1.915
c531 ( 141 0 ) capacitor c=0.0229444f //x=0.81 //y=1.53
c532 ( 140 0 ) capacitor c=0.0234352f //x=0.81 //y=1.22
c533 ( 139 0 ) capacitor c=0.0198724f //x=0.81 //y=0.875
c534 ( 138 0 ) capacitor c=0.15358f //x=24.9 //y=6.02
c535 ( 137 0 ) capacitor c=0.116098f //x=24.46 //y=6.02
c536 ( 136 0 ) capacitor c=0.116091f //x=24.02 //y=6.02
c537 ( 135 0 ) capacitor c=0.154305f //x=23.58 //y=6.02
c538 ( 134 0 ) capacitor c=0.15358f //x=11.95 //y=6.02
c539 ( 133 0 ) capacitor c=0.110281f //x=11.51 //y=6.02
c540 ( 132 0 ) capacitor c=0.110114f //x=1.75 //y=6.02
c541 ( 131 0 ) capacitor c=0.158956f //x=1.31 //y=6.02
c542 ( 124 0 ) capacitor c=0.00106608f //x=21.05 //y=5.155
c543 ( 123 0 ) capacitor c=0.00207319f //x=20.17 //y=5.155
c544 ( 122 0 ) capacitor c=0.00106608f //x=16.24 //y=5.155
c545 ( 121 0 ) capacitor c=0.00207162f //x=15.36 //y=5.155
c546 ( 115 0 ) capacitor c=0.0695278f //x=24.42 //y=2.08
c547 ( 113 0 ) capacitor c=0.00453889f //x=24.42 //y=4.535
c548 ( 106 0 ) capacitor c=0.0878398f //x=23.68 //y=2.08
c549 ( 104 0 ) capacitor c=0.109391f //x=21.83 //y=4.07
c550 ( 100 0 ) capacitor c=0.00398962f //x=21.43 //y=1.665
c551 ( 99 0 ) capacitor c=0.0137288f //x=21.745 //y=1.665
c552 ( 93 0 ) capacitor c=0.0284988f //x=21.745 //y=5.155
c553 ( 85 0 ) capacitor c=0.0176454f //x=20.965 //y=5.155
c554 ( 78 0 ) capacitor c=0.00332903f //x=19.375 //y=5.155
c555 ( 77 0 ) capacitor c=0.0148427f //x=20.085 //y=5.155
c556 ( 70 0 ) capacitor c=0.109457f //x=17.02 //y=4.07
c557 ( 66 0 ) capacitor c=0.00398962f //x=16.62 //y=1.665
c558 ( 65 0 ) capacitor c=0.0137288f //x=16.935 //y=1.665
c559 ( 59 0 ) capacitor c=0.0283082f //x=16.935 //y=5.155
c560 ( 51 0 ) capacitor c=0.0176454f //x=16.155 //y=5.155
c561 ( 44 0 ) capacitor c=0.00332903f //x=14.565 //y=5.155
c562 ( 43 0 ) capacitor c=0.014837f //x=15.275 //y=5.155
c563 ( 33 0 ) capacitor c=0.0700114f //x=11.47 //y=2.08
c564 ( 31 0 ) capacitor c=0.00453889f //x=11.47 //y=4.535
c565 ( 24 0 ) capacitor c=0.124161f //x=1.11 //y=2.08
c566 ( 10 0 ) capacitor c=0.00274864f //x=23.795 //y=4.07
c567 ( 9 0 ) capacitor c=0.0190681f //x=24.305 //y=4.07
c568 ( 8 0 ) capacitor c=0.00457352f //x=21.945 //y=4.07
c569 ( 7 0 ) capacitor c=0.0387588f //x=23.565 //y=4.07
c570 ( 6 0 ) capacitor c=0.00554824f //x=17.135 //y=4.07
c571 ( 5 0 ) capacitor c=0.0842645f //x=21.715 //y=4.07
c572 ( 4 0 ) capacitor c=0.00557292f //x=11.585 //y=4.07
c573 ( 3 0 ) capacitor c=0.0725278f //x=16.905 //y=4.07
c574 ( 2 0 ) capacitor c=0.0160831f //x=1.225 //y=4.07
c575 ( 1 0 ) capacitor c=0.183938f //x=11.355 //y=4.07
r576 (  250 251 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=24.45 //y=4.79 //x2=24.45 //y2=4.865
r577 (  248 250 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=24.45 //y=4.7 //x2=24.45 //y2=4.79
r578 (  244 245 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=24.42 //y=2.08 //x2=24.42 //y2=1.915
r579 (  238 240 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=23.58 //y=4.7 //x2=23.68 //y2=4.7
r580 (  228 229 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=11.5 //y=4.79 //x2=11.5 //y2=4.865
r581 (  226 228 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=11.5 //y=4.7 //x2=11.5 //y2=4.79
r582 (  222 223 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=11.47 //y=2.08 //x2=11.47 //y2=1.915
r583 (  212 255 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.985 //y=1.25 //x2=24.945 //y2=1.405
r584 (  211 254 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.985 //y=0.905 //x2=24.945 //y2=0.75
r585 (  211 212 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.985 //y=0.905 //x2=24.985 //y2=1.25
r586 (  206 253 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.61 //y=1.405 //x2=24.495 //y2=1.405
r587 (  205 255 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.83 //y=1.405 //x2=24.945 //y2=1.405
r588 (  204 252 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.61 //y=0.75 //x2=24.495 //y2=0.75
r589 (  203 254 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.83 //y=0.75 //x2=24.945 //y2=0.75
r590 (  203 204 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=24.83 //y=0.75 //x2=24.61 //y2=0.75
r591 (  202 250 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=24.585 //y=4.79 //x2=24.45 //y2=4.79
r592 (  201 208 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=24.825 //y=4.79 //x2=24.9 //y2=4.865
r593 (  201 202 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=24.825 //y=4.79 //x2=24.585 //y2=4.79
r594 (  196 253 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.455 //y=1.56 //x2=24.495 //y2=1.405
r595 (  196 245 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=24.455 //y=1.56 //x2=24.455 //y2=1.915
r596 (  195 253 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.455 //y=1.25 //x2=24.495 //y2=1.405
r597 (  194 252 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.455 //y=0.905 //x2=24.495 //y2=0.75
r598 (  194 195 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.455 //y=0.905 //x2=24.455 //y2=1.25
r599 (  191 240 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=24.02 //y=4.865 //x2=23.68 //y2=4.7
r600 (  190 242 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.015 //y=1.21 //x2=23.975 //y2=1.365
r601 (  189 241 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.015 //y=0.865 //x2=23.975 //y2=0.71
r602 (  189 190 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.015 //y=0.865 //x2=24.015 //y2=1.21
r603 (  187 237 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.64 //y=1.365 //x2=23.525 //y2=1.365
r604 (  186 242 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.86 //y=1.365 //x2=23.975 //y2=1.365
r605 (  185 236 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.64 //y=0.71 //x2=23.525 //y2=0.71
r606 (  184 241 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.86 //y=0.71 //x2=23.975 //y2=0.71
r607 (  184 185 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=23.86 //y=0.71 //x2=23.64 //y2=0.71
r608 (  181 238 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=23.58 //y=4.865 //x2=23.58 //y2=4.7
r609 (  180 235 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=23.485 //y=1.915 //x2=23.68 //y2=2.08
r610 (  179 237 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.485 //y=1.52 //x2=23.525 //y2=1.365
r611 (  179 180 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=23.485 //y=1.52 //x2=23.485 //y2=1.915
r612 (  178 237 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.485 //y=1.21 //x2=23.525 //y2=1.365
r613 (  177 236 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.485 //y=0.865 //x2=23.525 //y2=0.71
r614 (  177 178 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=23.485 //y=0.865 //x2=23.485 //y2=1.21
r615 (  176 233 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.035 //y=1.25 //x2=11.995 //y2=1.405
r616 (  175 232 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.035 //y=0.905 //x2=11.995 //y2=0.75
r617 (  175 176 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.035 //y=0.905 //x2=12.035 //y2=1.25
r618 (  170 231 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.66 //y=1.405 //x2=11.545 //y2=1.405
r619 (  169 233 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.88 //y=1.405 //x2=11.995 //y2=1.405
r620 (  168 230 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.66 //y=0.75 //x2=11.545 //y2=0.75
r621 (  167 232 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.88 //y=0.75 //x2=11.995 //y2=0.75
r622 (  167 168 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=11.88 //y=0.75 //x2=11.66 //y2=0.75
r623 (  166 228 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=11.635 //y=4.79 //x2=11.5 //y2=4.79
r624 (  165 172 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=11.875 //y=4.79 //x2=11.95 //y2=4.865
r625 (  165 166 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=11.875 //y=4.79 //x2=11.635 //y2=4.79
r626 (  160 231 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.505 //y=1.56 //x2=11.545 //y2=1.405
r627 (  160 223 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=11.505 //y=1.56 //x2=11.505 //y2=1.915
r628 (  159 231 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.505 //y=1.25 //x2=11.545 //y2=1.405
r629 (  158 230 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.505 //y=0.905 //x2=11.545 //y2=0.75
r630 (  158 159 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.505 //y=0.905 //x2=11.505 //y2=1.25
r631 (  153 155 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.75 //y2=4.865
r632 (  153 154 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.385 //y2=4.79
r633 (  152 220 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=1.22 //x2=1.3 //y2=1.375
r634 (  151 219 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.3 //y2=0.72
r635 (  151 152 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.34 //y2=1.22
r636 (  148 154 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.385 //y2=4.79
r637 (  148 218 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.11 //y2=4.7
r638 (  146 214 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=1.375 //x2=0.85 //y2=1.375
r639 (  145 220 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=1.375 //x2=1.3 //y2=1.375
r640 (  144 213 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=0.72 //x2=0.85 //y2=0.72
r641 (  143 219 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=1.3 //y2=0.72
r642 (  143 144 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=0.965 //y2=0.72
r643 (  142 216 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.915 //x2=1.11 //y2=2.08
r644 (  141 214 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.85 //y2=1.375
r645 (  141 142 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.81 //y2=1.915
r646 (  140 214 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.22 //x2=0.85 //y2=1.375
r647 (  139 213 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.85 //y2=0.72
r648 (  139 140 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.81 //y2=1.22
r649 (  138 208 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=24.9 //y=6.02 //x2=24.9 //y2=4.865
r650 (  137 251 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=24.46 //y=6.02 //x2=24.46 //y2=4.865
r651 (  136 191 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=24.02 //y=6.02 //x2=24.02 //y2=4.865
r652 (  135 181 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=23.58 //y=6.02 //x2=23.58 //y2=4.865
r653 (  134 172 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.95 //y=6.02 //x2=11.95 //y2=4.865
r654 (  133 229 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.51 //y=6.02 //x2=11.51 //y2=4.865
r655 (  132 155 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.75 //y=6.02 //x2=1.75 //y2=4.865
r656 (  131 148 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.31 //y=6.02 //x2=1.31 //y2=4.865
r657 (  130 205 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=24.72 //y=1.405 //x2=24.83 //y2=1.405
r658 (  130 206 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=24.72 //y=1.405 //x2=24.61 //y2=1.405
r659 (  129 186 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.75 //y=1.365 //x2=23.86 //y2=1.365
r660 (  129 187 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.75 //y=1.365 //x2=23.64 //y2=1.365
r661 (  128 169 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.77 //y=1.405 //x2=11.88 //y2=1.405
r662 (  128 170 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.77 //y=1.405 //x2=11.66 //y2=1.405
r663 (  127 145 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=1.185 //y2=1.375
r664 (  127 146 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=0.965 //y2=1.375
r665 (  126 248 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=24.45 //y=4.7 //x2=24.45 //y2=4.7
r666 (  120 226 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.5 //y=4.7 //x2=11.5 //y2=4.7
r667 (  115 244 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=24.42 //y=2.08 //x2=24.42 //y2=2.08
r668 (  115 118 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=24.42 //y=2.08 //x2=24.42 //y2=4.07
r669 (  113 126 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=24.42 //y=4.535 //x2=24.435 //y2=4.7
r670 (  113 118 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=24.42 //y=4.535 //x2=24.42 //y2=4.07
r671 (  111 240 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=23.68 //y=4.7 //x2=23.68 //y2=4.7
r672 (  109 111 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=23.68 //y=4.07 //x2=23.68 //y2=4.7
r673 (  106 235 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=23.68 //y=2.08 //x2=23.68 //y2=2.08
r674 (  106 109 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=23.68 //y=2.08 //x2=23.68 //y2=4.07
r675 (  102 104 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li \
 //thickness=0.1 //x=21.83 //y=5.07 //x2=21.83 //y2=4.07
r676 (  101 104 ) resistor r=158.802 //w=0.187 //l=2.32 //layer=li \
 //thickness=0.1 //x=21.83 //y=1.75 //x2=21.83 //y2=4.07
r677 (  99 101 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.745 //y=1.665 //x2=21.83 //y2=1.75
r678 (  99 100 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=21.745 //y=1.665 //x2=21.43 //y2=1.665
r679 (  95 100 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.345 //y=1.58 //x2=21.43 //y2=1.665
r680 (  95 257 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=21.345 //y=1.58 //x2=21.345 //y2=1.01
r681 (  94 124 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.135 //y=5.155 //x2=21.05 //y2=5.155
r682 (  93 102 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.745 //y=5.155 //x2=21.83 //y2=5.07
r683 (  93 94 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=21.745 //y=5.155 //x2=21.135 //y2=5.155
r684 (  87 124 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.05 //y=5.24 //x2=21.05 //y2=5.155
r685 (  87 265 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.05 //y=5.24 //x2=21.05 //y2=5.725
r686 (  86 123 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.255 //y=5.155 //x2=20.17 //y2=5.155
r687 (  85 124 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.965 //y=5.155 //x2=21.05 //y2=5.155
r688 (  85 86 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=20.965 //y=5.155 //x2=20.255 //y2=5.155
r689 (  79 123 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.17 //y=5.24 //x2=20.17 //y2=5.155
r690 (  79 264 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.17 //y=5.24 //x2=20.17 //y2=5.725
r691 (  77 123 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.085 //y=5.155 //x2=20.17 //y2=5.155
r692 (  77 78 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=20.085 //y=5.155 //x2=19.375 //y2=5.155
r693 (  71 78 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=19.29 //y=5.24 //x2=19.375 //y2=5.155
r694 (  71 263 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=19.29 //y=5.24 //x2=19.29 //y2=5.725
r695 (  68 70 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=17.02 //y=5.07 //x2=17.02 //y2=4.07
r696 (  67 70 ) resistor r=158.802 //w=0.187 //l=2.32 //layer=li \
 //thickness=0.1 //x=17.02 //y=1.75 //x2=17.02 //y2=4.07
r697 (  65 67 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.935 //y=1.665 //x2=17.02 //y2=1.75
r698 (  65 66 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=16.935 //y=1.665 //x2=16.62 //y2=1.665
r699 (  61 66 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.535 //y=1.58 //x2=16.62 //y2=1.665
r700 (  61 256 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=16.535 //y=1.58 //x2=16.535 //y2=1.01
r701 (  60 122 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.325 //y=5.155 //x2=16.24 //y2=5.155
r702 (  59 68 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.935 //y=5.155 //x2=17.02 //y2=5.07
r703 (  59 60 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=16.935 //y=5.155 //x2=16.325 //y2=5.155
r704 (  53 122 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.24 //y=5.24 //x2=16.24 //y2=5.155
r705 (  53 262 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.24 //y=5.24 //x2=16.24 //y2=5.725
r706 (  52 121 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.445 //y=5.155 //x2=15.36 //y2=5.155
r707 (  51 122 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.155 //y=5.155 //x2=16.24 //y2=5.155
r708 (  51 52 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=16.155 //y=5.155 //x2=15.445 //y2=5.155
r709 (  45 121 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.36 //y=5.24 //x2=15.36 //y2=5.155
r710 (  45 261 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.36 //y=5.24 //x2=15.36 //y2=5.725
r711 (  43 121 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.275 //y=5.155 //x2=15.36 //y2=5.155
r712 (  43 44 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=15.275 //y=5.155 //x2=14.565 //y2=5.155
r713 (  37 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.48 //y=5.24 //x2=14.565 //y2=5.155
r714 (  37 260 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.48 //y=5.24 //x2=14.48 //y2=5.725
r715 (  33 222 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.47 //y=2.08 //x2=11.47 //y2=2.08
r716 (  33 36 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=11.47 //y=2.08 //x2=11.47 //y2=4.07
r717 (  31 120 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=11.47 //y=4.535 //x2=11.485 //y2=4.7
r718 (  31 36 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=11.47 //y=4.535 //x2=11.47 //y2=4.07
r719 (  29 218 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r720 (  27 29 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.07 //x2=1.11 //y2=4.7
r721 (  24 216 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r722 (  24 27 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.08 //x2=1.11 //y2=4.07
r723 (  22 118 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=24.42 //y=4.07 //x2=24.42 //y2=4.07
r724 (  20 109 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=23.68 //y=4.07 //x2=23.68 //y2=4.07
r725 (  18 104 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.83 //y=4.07 //x2=21.83 //y2=4.07
r726 (  16 70 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.02 //y=4.07 //x2=17.02 //y2=4.07
r727 (  14 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.47 //y=4.07 //x2=11.47 //y2=4.07
r728 (  12 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.07
r729 (  10 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.795 //y=4.07 //x2=23.68 //y2=4.07
r730 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=24.305 //y=4.07 //x2=24.42 //y2=4.07
r731 (  9 10 ) resistor r=0.486641 //w=0.131 //l=0.51 //layer=m1 \
 //thickness=0.36 //x=24.305 //y=4.07 //x2=23.795 //y2=4.07
r732 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.945 //y=4.07 //x2=21.83 //y2=4.07
r733 (  7 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.565 //y=4.07 //x2=23.68 //y2=4.07
r734 (  7 8 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=23.565 //y=4.07 //x2=21.945 //y2=4.07
r735 (  6 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.135 //y=4.07 //x2=17.02 //y2=4.07
r736 (  5 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.715 //y=4.07 //x2=21.83 //y2=4.07
r737 (  5 6 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=21.715 //y=4.07 //x2=17.135 //y2=4.07
r738 (  4 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.585 //y=4.07 //x2=11.47 //y2=4.07
r739 (  3 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.905 //y=4.07 //x2=17.02 //y2=4.07
r740 (  3 4 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=16.905 //y=4.07 //x2=11.585 //y2=4.07
r741 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.225 //y=4.07 //x2=1.11 //y2=4.07
r742 (  1 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.355 //y=4.07 //x2=11.47 //y2=4.07
r743 (  1 2 ) resistor r=9.66603 //w=0.131 //l=10.13 //layer=m1 \
 //thickness=0.36 //x=11.355 //y=4.07 //x2=1.225 //y2=4.07
ends PM_TMRDFFRNQNX1\%noxref_6

subckt PM_TMRDFFRNQNX1\%noxref_7 ( 1 2 3 4 12 25 26 33 41 47 48 52 54 61 62 63 \
 64 65 66 67 68 72 73 74 79 81 84 85 86 87 88 89 93 95 98 99 104 105 110 119 \
 122 124 125 126 )
c247 ( 126 0 ) capacitor c=0.023087f //x=33.855 //y=5.02
c248 ( 125 0 ) capacitor c=0.023519f //x=32.975 //y=5.02
c249 ( 124 0 ) capacitor c=0.0224735f //x=32.095 //y=5.02
c250 ( 122 0 ) capacitor c=0.00872971f //x=34.105 //y=0.915
c251 ( 119 0 ) capacitor c=0.0588816f //x=36.63 //y=4.7
c252 ( 110 0 ) capacitor c=0.058931f //x=29.23 //y=4.7
c253 ( 105 0 ) capacitor c=0.0273931f //x=29.23 //y=1.915
c254 ( 104 0 ) capacitor c=0.0456313f //x=29.23 //y=2.08
c255 ( 99 0 ) capacitor c=0.0318948f //x=36.965 //y=1.21
c256 ( 98 0 ) capacitor c=0.0187384f //x=36.965 //y=0.865
c257 ( 95 0 ) capacitor c=0.0141798f //x=36.81 //y=1.365
c258 ( 93 0 ) capacitor c=0.0149844f //x=36.81 //y=0.71
c259 ( 89 0 ) capacitor c=0.0813322f //x=36.435 //y=1.915
c260 ( 88 0 ) capacitor c=0.0229267f //x=36.435 //y=1.52
c261 ( 87 0 ) capacitor c=0.0234352f //x=36.435 //y=1.21
c262 ( 86 0 ) capacitor c=0.0199343f //x=36.435 //y=0.865
c263 ( 85 0 ) capacitor c=0.0432517f //x=29.75 //y=1.26
c264 ( 84 0 ) capacitor c=0.0200379f //x=29.75 //y=0.915
c265 ( 81 0 ) capacitor c=0.0148873f //x=29.595 //y=1.415
c266 ( 79 0 ) capacitor c=0.0157803f //x=29.595 //y=0.76
c267 ( 74 0 ) capacitor c=0.0218028f //x=29.22 //y=1.57
c268 ( 73 0 ) capacitor c=0.0207459f //x=29.22 //y=1.26
c269 ( 72 0 ) capacitor c=0.0194308f //x=29.22 //y=0.915
c270 ( 68 0 ) capacitor c=0.110275f //x=36.97 //y=6.02
c271 ( 67 0 ) capacitor c=0.154305f //x=36.53 //y=6.02
c272 ( 66 0 ) capacitor c=0.158794f //x=29.41 //y=6.02
c273 ( 65 0 ) capacitor c=0.110114f //x=28.97 //y=6.02
c274 ( 62 0 ) capacitor c=0.00106608f //x=34 //y=5.155
c275 ( 61 0 ) capacitor c=0.00207319f //x=33.12 //y=5.155
c276 ( 54 0 ) capacitor c=0.084205f //x=36.63 //y=2.08
c277 ( 52 0 ) capacitor c=0.103747f //x=34.78 //y=3.33
c278 ( 48 0 ) capacitor c=0.00398962f //x=34.38 //y=1.665
c279 ( 47 0 ) capacitor c=0.0137288f //x=34.695 //y=1.665
c280 ( 41 0 ) capacitor c=0.0284988f //x=34.695 //y=5.155
c281 ( 33 0 ) capacitor c=0.0176454f //x=33.915 //y=5.155
c282 ( 26 0 ) capacitor c=0.00332903f //x=32.325 //y=5.155
c283 ( 25 0 ) capacitor c=0.0148427f //x=33.035 //y=5.155
c284 ( 12 0 ) capacitor c=0.081384f //x=29.23 //y=2.08
c285 ( 4 0 ) capacitor c=0.00427986f //x=34.895 //y=3.33
c286 ( 3 0 ) capacitor c=0.0347042f //x=36.515 //y=3.33
c287 ( 2 0 ) capacitor c=0.0141678f //x=29.345 //y=3.33
c288 ( 1 0 ) capacitor c=0.077708f //x=34.665 //y=3.33
r289 (  117 119 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=36.53 //y=4.7 //x2=36.63 //y2=4.7
r290 (  104 105 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=29.23 //y=2.08 //x2=29.23 //y2=1.915
r291 (  100 119 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=36.97 //y=4.865 //x2=36.63 //y2=4.7
r292 (  99 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.965 //y=1.21 //x2=36.925 //y2=1.365
r293 (  98 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.965 //y=0.865 //x2=36.925 //y2=0.71
r294 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=36.965 //y=0.865 //x2=36.965 //y2=1.21
r295 (  96 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=36.59 //y=1.365 //x2=36.475 //y2=1.365
r296 (  95 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=36.81 //y=1.365 //x2=36.925 //y2=1.365
r297 (  94 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=36.59 //y=0.71 //x2=36.475 //y2=0.71
r298 (  93 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=36.81 //y=0.71 //x2=36.925 //y2=0.71
r299 (  93 94 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=36.81 //y=0.71 //x2=36.59 //y2=0.71
r300 (  90 117 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=36.53 //y=4.865 //x2=36.53 //y2=4.7
r301 (  89 114 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=36.435 //y=1.915 //x2=36.63 //y2=2.08
r302 (  88 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.435 //y=1.52 //x2=36.475 //y2=1.365
r303 (  88 89 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=36.435 //y=1.52 //x2=36.435 //y2=1.915
r304 (  87 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.435 //y=1.21 //x2=36.475 //y2=1.365
r305 (  86 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.435 //y=0.865 //x2=36.475 //y2=0.71
r306 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=36.435 //y=0.865 //x2=36.435 //y2=1.21
r307 (  85 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.75 //y=1.26 //x2=29.71 //y2=1.415
r308 (  84 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.75 //y=0.915 //x2=29.71 //y2=0.76
r309 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=29.75 //y=0.915 //x2=29.75 //y2=1.26
r310 (  82 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.375 //y=1.415 //x2=29.26 //y2=1.415
r311 (  81 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.595 //y=1.415 //x2=29.71 //y2=1.415
r312 (  80 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.375 //y=0.76 //x2=29.26 //y2=0.76
r313 (  79 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.595 //y=0.76 //x2=29.71 //y2=0.76
r314 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=29.595 //y=0.76 //x2=29.375 //y2=0.76
r315 (  76 110 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=29.41 //y=4.865 //x2=29.23 //y2=4.7
r316 (  74 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.22 //y=1.57 //x2=29.26 //y2=1.415
r317 (  74 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=29.22 //y=1.57 //x2=29.22 //y2=1.915
r318 (  73 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.22 //y=1.26 //x2=29.26 //y2=1.415
r319 (  72 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.22 //y=0.915 //x2=29.26 //y2=0.76
r320 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=29.22 //y=0.915 //x2=29.22 //y2=1.26
r321 (  69 110 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=28.97 //y=4.865 //x2=29.23 //y2=4.7
r322 (  68 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=36.97 //y=6.02 //x2=36.97 //y2=4.865
r323 (  67 90 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=36.53 //y=6.02 //x2=36.53 //y2=4.865
r324 (  66 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=29.41 //y=6.02 //x2=29.41 //y2=4.865
r325 (  65 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=28.97 //y=6.02 //x2=28.97 //y2=4.865
r326 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=36.7 //y=1.365 //x2=36.81 //y2=1.365
r327 (  64 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=36.7 //y=1.365 //x2=36.59 //y2=1.365
r328 (  63 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=29.485 //y=1.415 //x2=29.595 //y2=1.415
r329 (  63 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=29.485 //y=1.415 //x2=29.375 //y2=1.415
r330 (  59 119 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=36.63 //y=4.7 //x2=36.63 //y2=4.7
r331 (  57 59 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=36.63 //y=3.33 //x2=36.63 //y2=4.7
r332 (  54 114 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=36.63 //y=2.08 //x2=36.63 //y2=2.08
r333 (  54 57 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=36.63 //y=2.08 //x2=36.63 //y2=3.33
r334 (  50 52 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=34.78 //y=5.07 //x2=34.78 //y2=3.33
r335 (  49 52 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=34.78 //y=1.75 //x2=34.78 //y2=3.33
r336 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=34.695 //y=1.665 //x2=34.78 //y2=1.75
r337 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=34.695 //y=1.665 //x2=34.38 //y2=1.665
r338 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=34.295 //y=1.58 //x2=34.38 //y2=1.665
r339 (  43 122 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=34.295 //y=1.58 //x2=34.295 //y2=1.01
r340 (  42 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.085 //y=5.155 //x2=34 //y2=5.155
r341 (  41 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=34.695 //y=5.155 //x2=34.78 //y2=5.07
r342 (  41 42 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=34.695 //y=5.155 //x2=34.085 //y2=5.155
r343 (  35 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34 //y=5.24 //x2=34 //y2=5.155
r344 (  35 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=34 //y=5.24 //x2=34 //y2=5.725
r345 (  34 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.205 //y=5.155 //x2=33.12 //y2=5.155
r346 (  33 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.915 //y=5.155 //x2=34 //y2=5.155
r347 (  33 34 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=33.915 //y=5.155 //x2=33.205 //y2=5.155
r348 (  27 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.12 //y=5.24 //x2=33.12 //y2=5.155
r349 (  27 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=33.12 //y=5.24 //x2=33.12 //y2=5.725
r350 (  25 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.035 //y=5.155 //x2=33.12 //y2=5.155
r351 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=33.035 //y=5.155 //x2=32.325 //y2=5.155
r352 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=32.24 //y=5.24 //x2=32.325 //y2=5.155
r353 (  19 124 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=32.24 //y=5.24 //x2=32.24 //y2=5.725
r354 (  17 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=29.23 //y=4.7 //x2=29.23 //y2=4.7
r355 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=29.23 //y=3.33 //x2=29.23 //y2=4.7
r356 (  12 104 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=29.23 //y=2.08 //x2=29.23 //y2=2.08
r357 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=29.23 //y=2.08 //x2=29.23 //y2=3.33
r358 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=36.63 //y=3.33 //x2=36.63 //y2=3.33
r359 (  8 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=34.78 //y=3.33 //x2=34.78 //y2=3.33
r360 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=29.23 //y=3.33 //x2=29.23 //y2=3.33
r361 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.895 //y=3.33 //x2=34.78 //y2=3.33
r362 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=36.515 //y=3.33 //x2=36.63 //y2=3.33
r363 (  3 4 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=36.515 //y=3.33 //x2=34.895 //y2=3.33
r364 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=29.345 //y=3.33 //x2=29.23 //y2=3.33
r365 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.665 //y=3.33 //x2=34.78 //y2=3.33
r366 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=34.665 //y=3.33 //x2=29.345 //y2=3.33
ends PM_TMRDFFRNQNX1\%noxref_7

subckt PM_TMRDFFRNQNX1\%noxref_8 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 \
 47 48 49 51 57 58 59 60 72 74 75 )
c153 ( 75 0 ) capacitor c=0.0220291f //x=37.485 //y=5.02
c154 ( 74 0 ) capacitor c=0.0217503f //x=36.605 //y=5.02
c155 ( 72 0 ) capacitor c=0.0084702f //x=37.48 //y=0.905
c156 ( 60 0 ) capacitor c=0.0557698f //x=40.235 //y=4.79
c157 ( 59 0 ) capacitor c=0.0293157f //x=40.525 //y=4.79
c158 ( 58 0 ) capacitor c=0.0347816f //x=40.19 //y=1.22
c159 ( 57 0 ) capacitor c=0.0187487f //x=40.19 //y=0.875
c160 ( 51 0 ) capacitor c=0.0137055f //x=40.035 //y=1.375
c161 ( 49 0 ) capacitor c=0.0149861f //x=40.035 //y=0.72
c162 ( 48 0 ) capacitor c=0.096037f //x=39.66 //y=1.915
c163 ( 47 0 ) capacitor c=0.0228993f //x=39.66 //y=1.53
c164 ( 46 0 ) capacitor c=0.0234352f //x=39.66 //y=1.22
c165 ( 45 0 ) capacitor c=0.0198724f //x=39.66 //y=0.875
c166 ( 44 0 ) capacitor c=0.110114f //x=40.6 //y=6.02
c167 ( 43 0 ) capacitor c=0.158956f //x=40.16 //y=6.02
c168 ( 41 0 ) capacitor c=0.00211606f //x=37.63 //y=5.2
c169 ( 34 0 ) capacitor c=0.0936549f //x=39.96 //y=2.08
c170 ( 32 0 ) capacitor c=0.102772f //x=38.11 //y=3.33
c171 ( 28 0 ) capacitor c=0.00404073f //x=37.755 //y=1.655
c172 ( 27 0 ) capacitor c=0.0122201f //x=38.025 //y=1.655
c173 ( 25 0 ) capacitor c=0.0137995f //x=38.025 //y=5.2
c174 ( 14 0 ) capacitor c=0.00251635f //x=36.835 //y=5.2
c175 ( 13 0 ) capacitor c=0.0143649f //x=37.545 //y=5.2
c176 ( 2 0 ) capacitor c=0.00668619f //x=38.225 //y=3.33
c177 ( 1 0 ) capacitor c=0.0402621f //x=39.845 //y=3.33
r178 (  59 61 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=40.525 //y=4.79 //x2=40.6 //y2=4.865
r179 (  59 60 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=40.525 //y=4.79 //x2=40.235 //y2=4.79
r180 (  58 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.19 //y=1.22 //x2=40.15 //y2=1.375
r181 (  57 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.19 //y=0.875 //x2=40.15 //y2=0.72
r182 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=40.19 //y=0.875 //x2=40.19 //y2=1.22
r183 (  54 60 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=40.16 //y=4.865 //x2=40.235 //y2=4.79
r184 (  54 69 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=40.16 //y=4.865 //x2=39.96 //y2=4.7
r185 (  52 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.815 //y=1.375 //x2=39.7 //y2=1.375
r186 (  51 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.035 //y=1.375 //x2=40.15 //y2=1.375
r187 (  50 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.815 //y=0.72 //x2=39.7 //y2=0.72
r188 (  49 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.035 //y=0.72 //x2=40.15 //y2=0.72
r189 (  49 50 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=40.035 //y=0.72 //x2=39.815 //y2=0.72
r190 (  48 67 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=39.66 //y=1.915 //x2=39.96 //y2=2.08
r191 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.66 //y=1.53 //x2=39.7 //y2=1.375
r192 (  47 48 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=39.66 //y=1.53 //x2=39.66 //y2=1.915
r193 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.66 //y=1.22 //x2=39.7 //y2=1.375
r194 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.66 //y=0.875 //x2=39.7 //y2=0.72
r195 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=39.66 //y=0.875 //x2=39.66 //y2=1.22
r196 (  44 61 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=40.6 //y=6.02 //x2=40.6 //y2=4.865
r197 (  43 54 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=40.16 //y=6.02 //x2=40.16 //y2=4.865
r198 (  42 51 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=39.925 //y=1.375 //x2=40.035 //y2=1.375
r199 (  42 52 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=39.925 //y=1.375 //x2=39.815 //y2=1.375
r200 (  39 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=39.96 //y=4.7 //x2=39.96 //y2=4.7
r201 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=39.96 //y=3.33 //x2=39.96 //y2=4.7
r202 (  34 67 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=39.96 //y=2.08 //x2=39.96 //y2=2.08
r203 (  34 37 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=39.96 //y=2.08 //x2=39.96 //y2=3.33
r204 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=38.11 //y=5.115 //x2=38.11 //y2=3.33
r205 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=38.11 //y=1.74 //x2=38.11 //y2=3.33
r206 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=38.025 //y=1.655 //x2=38.11 //y2=1.74
r207 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=38.025 //y=1.655 //x2=37.755 //y2=1.655
r208 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.715 //y=5.2 //x2=37.63 //y2=5.2
r209 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=38.025 //y=5.2 //x2=38.11 //y2=5.115
r210 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=38.025 //y=5.2 //x2=37.715 //y2=5.2
r211 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=37.67 //y=1.57 //x2=37.755 //y2=1.655
r212 (  21 72 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=37.67 //y=1.57 //x2=37.67 //y2=1
r213 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.63 //y=5.285 //x2=37.63 //y2=5.2
r214 (  15 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=37.63 //y=5.285 //x2=37.63 //y2=5.725
r215 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=37.545 //y=5.2 //x2=37.63 //y2=5.2
r216 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=37.545 //y=5.2 //x2=36.835 //y2=5.2
r217 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=36.75 //y=5.285 //x2=36.835 //y2=5.2
r218 (  7 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=36.75 //y=5.285 //x2=36.75 //y2=5.725
r219 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=39.96 //y=3.33 //x2=39.96 //y2=3.33
r220 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=38.11 //y=3.33 //x2=38.11 //y2=3.33
r221 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=38.225 //y=3.33 //x2=38.11 //y2=3.33
r222 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=39.845 //y=3.33 //x2=39.96 //y2=3.33
r223 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=39.845 //y=3.33 //x2=38.225 //y2=3.33
ends PM_TMRDFFRNQNX1\%noxref_8

subckt PM_TMRDFFRNQNX1\%noxref_9 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 63 \
 64 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 92 94 100 101 102 \
 103 123 125 126 127 )
c262 ( 127 0 ) capacitor c=0.023087f //x=29.045 //y=5.02
c263 ( 126 0 ) capacitor c=0.023519f //x=28.165 //y=5.02
c264 ( 125 0 ) capacitor c=0.0224735f //x=27.285 //y=5.02
c265 ( 123 0 ) capacitor c=0.00853354f //x=29.295 //y=0.915
c266 ( 103 0 ) capacitor c=0.0556143f //x=45.045 //y=4.79
c267 ( 102 0 ) capacitor c=0.0293157f //x=45.335 //y=4.79
c268 ( 101 0 ) capacitor c=0.0347816f //x=45 //y=1.22
c269 ( 100 0 ) capacitor c=0.0187487f //x=45 //y=0.875
c270 ( 94 0 ) capacitor c=0.0137055f //x=44.845 //y=1.375
c271 ( 92 0 ) capacitor c=0.0149861f //x=44.845 //y=0.72
c272 ( 91 0 ) capacitor c=0.096037f //x=44.47 //y=1.915
c273 ( 90 0 ) capacitor c=0.0228993f //x=44.47 //y=1.53
c274 ( 89 0 ) capacitor c=0.0234352f //x=44.47 //y=1.22
c275 ( 88 0 ) capacitor c=0.0198724f //x=44.47 //y=0.875
c276 ( 84 0 ) capacitor c=0.0556143f //x=32.095 //y=4.79
c277 ( 83 0 ) capacitor c=0.0293157f //x=32.385 //y=4.79
c278 ( 82 0 ) capacitor c=0.0347816f //x=32.05 //y=1.22
c279 ( 81 0 ) capacitor c=0.0187487f //x=32.05 //y=0.875
c280 ( 75 0 ) capacitor c=0.0137055f //x=31.895 //y=1.375
c281 ( 73 0 ) capacitor c=0.0149861f //x=31.895 //y=0.72
c282 ( 72 0 ) capacitor c=0.096037f //x=31.52 //y=1.915
c283 ( 71 0 ) capacitor c=0.0228993f //x=31.52 //y=1.53
c284 ( 70 0 ) capacitor c=0.0234352f //x=31.52 //y=1.22
c285 ( 69 0 ) capacitor c=0.0198724f //x=31.52 //y=0.875
c286 ( 68 0 ) capacitor c=0.110114f //x=45.41 //y=6.02
c287 ( 67 0 ) capacitor c=0.158956f //x=44.97 //y=6.02
c288 ( 66 0 ) capacitor c=0.110114f //x=32.46 //y=6.02
c289 ( 65 0 ) capacitor c=0.158956f //x=32.02 //y=6.02
c290 ( 62 0 ) capacitor c=0.00106608f //x=29.19 //y=5.155
c291 ( 61 0 ) capacitor c=0.00207162f //x=28.31 //y=5.155
c292 ( 54 0 ) capacitor c=0.0974046f //x=44.77 //y=2.08
c293 ( 46 0 ) capacitor c=0.0936123f //x=31.82 //y=2.08
c294 ( 44 0 ) capacitor c=0.103742f //x=29.97 //y=3.7
c295 ( 40 0 ) capacitor c=0.00398962f //x=29.57 //y=1.665
c296 ( 39 0 ) capacitor c=0.0137288f //x=29.885 //y=1.665
c297 ( 33 0 ) capacitor c=0.0283082f //x=29.885 //y=5.155
c298 ( 25 0 ) capacitor c=0.0176454f //x=29.105 //y=5.155
c299 ( 18 0 ) capacitor c=0.00332903f //x=27.515 //y=5.155
c300 ( 17 0 ) capacitor c=0.014837f //x=28.225 //y=5.155
c301 ( 4 0 ) capacitor c=0.00424246f //x=31.935 //y=3.7
c302 ( 3 0 ) capacitor c=0.210233f //x=44.655 //y=3.7
c303 ( 2 0 ) capacitor c=0.0125346f //x=30.085 //y=3.7
c304 ( 1 0 ) capacitor c=0.0288301f //x=31.705 //y=3.7
r305 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=45.335 //y=4.79 //x2=45.41 //y2=4.865
r306 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=45.335 //y=4.79 //x2=45.045 //y2=4.79
r307 (  101 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45 //y=1.22 //x2=44.96 //y2=1.375
r308 (  100 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45 //y=0.875 //x2=44.96 //y2=0.72
r309 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=45 //y=0.875 //x2=45 //y2=1.22
r310 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=44.97 //y=4.865 //x2=45.045 //y2=4.79
r311 (  97 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=44.97 //y=4.865 //x2=44.77 //y2=4.7
r312 (  95 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.625 //y=1.375 //x2=44.51 //y2=1.375
r313 (  94 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.845 //y=1.375 //x2=44.96 //y2=1.375
r314 (  93 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.625 //y=0.72 //x2=44.51 //y2=0.72
r315 (  92 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.845 //y=0.72 //x2=44.96 //y2=0.72
r316 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=44.845 //y=0.72 //x2=44.625 //y2=0.72
r317 (  91 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=44.47 //y=1.915 //x2=44.77 //y2=2.08
r318 (  90 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.47 //y=1.53 //x2=44.51 //y2=1.375
r319 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=44.47 //y=1.53 //x2=44.47 //y2=1.915
r320 (  89 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.47 //y=1.22 //x2=44.51 //y2=1.375
r321 (  88 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.47 //y=0.875 //x2=44.51 //y2=0.72
r322 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=44.47 //y=0.875 //x2=44.47 //y2=1.22
r323 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=32.385 //y=4.79 //x2=32.46 //y2=4.865
r324 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=32.385 //y=4.79 //x2=32.095 //y2=4.79
r325 (  82 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.05 //y=1.22 //x2=32.01 //y2=1.375
r326 (  81 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.05 //y=0.875 //x2=32.01 //y2=0.72
r327 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=32.05 //y=0.875 //x2=32.05 //y2=1.22
r328 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=32.02 //y=4.865 //x2=32.095 //y2=4.79
r329 (  78 112 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=32.02 //y=4.865 //x2=31.82 //y2=4.7
r330 (  76 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.675 //y=1.375 //x2=31.56 //y2=1.375
r331 (  75 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.895 //y=1.375 //x2=32.01 //y2=1.375
r332 (  74 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.675 //y=0.72 //x2=31.56 //y2=0.72
r333 (  73 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.895 //y=0.72 //x2=32.01 //y2=0.72
r334 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=31.895 //y=0.72 //x2=31.675 //y2=0.72
r335 (  72 110 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=31.52 //y=1.915 //x2=31.82 //y2=2.08
r336 (  71 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.52 //y=1.53 //x2=31.56 //y2=1.375
r337 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=31.52 //y=1.53 //x2=31.52 //y2=1.915
r338 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.52 //y=1.22 //x2=31.56 //y2=1.375
r339 (  69 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.52 //y=0.875 //x2=31.56 //y2=0.72
r340 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=31.52 //y=0.875 //x2=31.52 //y2=1.22
r341 (  68 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.41 //y=6.02 //x2=45.41 //y2=4.865
r342 (  67 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=44.97 //y=6.02 //x2=44.97 //y2=4.865
r343 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=32.46 //y=6.02 //x2=32.46 //y2=4.865
r344 (  65 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=32.02 //y=6.02 //x2=32.02 //y2=4.865
r345 (  64 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=44.735 //y=1.375 //x2=44.845 //y2=1.375
r346 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=44.735 //y=1.375 //x2=44.625 //y2=1.375
r347 (  63 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=31.785 //y=1.375 //x2=31.895 //y2=1.375
r348 (  63 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=31.785 //y=1.375 //x2=31.675 //y2=1.375
r349 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=44.77 //y=4.7 //x2=44.77 //y2=4.7
r350 (  57 59 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=44.77 //y=3.7 //x2=44.77 //y2=4.7
r351 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=44.77 //y=2.08 //x2=44.77 //y2=2.08
r352 (  54 57 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=44.77 //y=2.08 //x2=44.77 //y2=3.7
r353 (  51 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.82 //y=4.7 //x2=31.82 //y2=4.7
r354 (  49 51 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=31.82 //y=3.7 //x2=31.82 //y2=4.7
r355 (  46 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.82 //y=2.08 //x2=31.82 //y2=2.08
r356 (  46 49 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=31.82 //y=2.08 //x2=31.82 //y2=3.7
r357 (  42 44 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=29.97 //y=5.07 //x2=29.97 //y2=3.7
r358 (  41 44 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=29.97 //y=1.75 //x2=29.97 //y2=3.7
r359 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=29.885 //y=1.665 //x2=29.97 //y2=1.75
r360 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=29.885 //y=1.665 //x2=29.57 //y2=1.665
r361 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=29.485 //y=1.58 //x2=29.57 //y2=1.665
r362 (  35 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=29.485 //y=1.58 //x2=29.485 //y2=1.01
r363 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.275 //y=5.155 //x2=29.19 //y2=5.155
r364 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=29.885 //y=5.155 //x2=29.97 //y2=5.07
r365 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=29.885 //y=5.155 //x2=29.275 //y2=5.155
r366 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.19 //y=5.24 //x2=29.19 //y2=5.155
r367 (  27 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=29.19 //y=5.24 //x2=29.19 //y2=5.725
r368 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.395 //y=5.155 //x2=28.31 //y2=5.155
r369 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.105 //y=5.155 //x2=29.19 //y2=5.155
r370 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=29.105 //y=5.155 //x2=28.395 //y2=5.155
r371 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.31 //y=5.24 //x2=28.31 //y2=5.155
r372 (  19 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=28.31 //y=5.24 //x2=28.31 //y2=5.725
r373 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.225 //y=5.155 //x2=28.31 //y2=5.155
r374 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=28.225 //y=5.155 //x2=27.515 //y2=5.155
r375 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=27.43 //y=5.24 //x2=27.515 //y2=5.155
r376 (  11 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=27.43 //y=5.24 //x2=27.43 //y2=5.725
r377 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=44.77 //y=3.7 //x2=44.77 //y2=3.7
r378 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=31.82 //y=3.7 //x2=31.82 //y2=3.7
r379 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=29.97 //y=3.7 //x2=29.97 //y2=3.7
r380 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.935 //y=3.7 //x2=31.82 //y2=3.7
r381 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=44.655 //y=3.7 //x2=44.77 //y2=3.7
r382 (  3 4 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=44.655 //y=3.7 //x2=31.935 //y2=3.7
r383 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=30.085 //y=3.7 //x2=29.97 //y2=3.7
r384 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.705 //y=3.7 //x2=31.82 //y2=3.7
r385 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=31.705 //y=3.7 //x2=30.085 //y2=3.7
ends PM_TMRDFFRNQNX1\%noxref_9

subckt PM_TMRDFFRNQNX1\%noxref_10 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 \
 54 55 56 57 61 63 66 67 77 80 82 83 84 )
c163 ( 84 0 ) capacitor c=0.023087f //x=46.805 //y=5.02
c164 ( 83 0 ) capacitor c=0.023519f //x=45.925 //y=5.02
c165 ( 82 0 ) capacitor c=0.0224735f //x=45.045 //y=5.02
c166 ( 80 0 ) capacitor c=0.00872971f //x=47.055 //y=0.915
c167 ( 77 0 ) capacitor c=0.0588816f //x=49.58 //y=4.7
c168 ( 67 0 ) capacitor c=0.0318948f //x=49.915 //y=1.21
c169 ( 66 0 ) capacitor c=0.0187384f //x=49.915 //y=0.865
c170 ( 63 0 ) capacitor c=0.0141798f //x=49.76 //y=1.365
c171 ( 61 0 ) capacitor c=0.0149844f //x=49.76 //y=0.71
c172 ( 57 0 ) capacitor c=0.0813322f //x=49.385 //y=1.915
c173 ( 56 0 ) capacitor c=0.0229267f //x=49.385 //y=1.52
c174 ( 55 0 ) capacitor c=0.0234352f //x=49.385 //y=1.21
c175 ( 54 0 ) capacitor c=0.0199343f //x=49.385 //y=0.865
c176 ( 53 0 ) capacitor c=0.110275f //x=49.92 //y=6.02
c177 ( 52 0 ) capacitor c=0.154305f //x=49.48 //y=6.02
c178 ( 50 0 ) capacitor c=0.00106608f //x=46.95 //y=5.155
c179 ( 49 0 ) capacitor c=0.00207319f //x=46.07 //y=5.155
c180 ( 42 0 ) capacitor c=0.0836545f //x=49.58 //y=2.08
c181 ( 40 0 ) capacitor c=0.104238f //x=47.73 //y=3.7
c182 ( 36 0 ) capacitor c=0.00398962f //x=47.33 //y=1.665
c183 ( 35 0 ) capacitor c=0.0137288f //x=47.645 //y=1.665
c184 ( 29 0 ) capacitor c=0.0284988f //x=47.645 //y=5.155
c185 ( 21 0 ) capacitor c=0.0176454f //x=46.865 //y=5.155
c186 ( 14 0 ) capacitor c=0.00332903f //x=45.275 //y=5.155
c187 ( 13 0 ) capacitor c=0.0148427f //x=45.985 //y=5.155
c188 ( 2 0 ) capacitor c=0.00854301f //x=47.845 //y=3.7
c189 ( 1 0 ) capacitor c=0.0405342f //x=49.465 //y=3.7
r190 (  75 77 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=49.48 //y=4.7 //x2=49.58 //y2=4.7
r191 (  68 77 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=49.92 //y=4.865 //x2=49.58 //y2=4.7
r192 (  67 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.915 //y=1.21 //x2=49.875 //y2=1.365
r193 (  66 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.915 //y=0.865 //x2=49.875 //y2=0.71
r194 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=49.915 //y=0.865 //x2=49.915 //y2=1.21
r195 (  64 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.54 //y=1.365 //x2=49.425 //y2=1.365
r196 (  63 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.76 //y=1.365 //x2=49.875 //y2=1.365
r197 (  62 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.54 //y=0.71 //x2=49.425 //y2=0.71
r198 (  61 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.76 //y=0.71 //x2=49.875 //y2=0.71
r199 (  61 62 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=49.76 //y=0.71 //x2=49.54 //y2=0.71
r200 (  58 75 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=49.48 //y=4.865 //x2=49.48 //y2=4.7
r201 (  57 72 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=49.385 //y=1.915 //x2=49.58 //y2=2.08
r202 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.385 //y=1.52 //x2=49.425 //y2=1.365
r203 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=49.385 //y=1.52 //x2=49.385 //y2=1.915
r204 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.385 //y=1.21 //x2=49.425 //y2=1.365
r205 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.385 //y=0.865 //x2=49.425 //y2=0.71
r206 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=49.385 //y=0.865 //x2=49.385 //y2=1.21
r207 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=49.92 //y=6.02 //x2=49.92 //y2=4.865
r208 (  52 58 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=49.48 //y=6.02 //x2=49.48 //y2=4.865
r209 (  51 63 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=49.65 //y=1.365 //x2=49.76 //y2=1.365
r210 (  51 64 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=49.65 //y=1.365 //x2=49.54 //y2=1.365
r211 (  47 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=49.58 //y=4.7 //x2=49.58 //y2=4.7
r212 (  45 47 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=49.58 //y=3.7 //x2=49.58 //y2=4.7
r213 (  42 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=49.58 //y=2.08 //x2=49.58 //y2=2.08
r214 (  42 45 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=49.58 //y=2.08 //x2=49.58 //y2=3.7
r215 (  38 40 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=47.73 //y=5.07 //x2=47.73 //y2=3.7
r216 (  37 40 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=47.73 //y=1.75 //x2=47.73 //y2=3.7
r217 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=47.645 //y=1.665 //x2=47.73 //y2=1.75
r218 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=47.645 //y=1.665 //x2=47.33 //y2=1.665
r219 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=47.245 //y=1.58 //x2=47.33 //y2=1.665
r220 (  31 80 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=47.245 //y=1.58 //x2=47.245 //y2=1.01
r221 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.035 //y=5.155 //x2=46.95 //y2=5.155
r222 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=47.645 //y=5.155 //x2=47.73 //y2=5.07
r223 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=47.645 //y=5.155 //x2=47.035 //y2=5.155
r224 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.95 //y=5.24 //x2=46.95 //y2=5.155
r225 (  23 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.95 //y=5.24 //x2=46.95 //y2=5.725
r226 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.155 //y=5.155 //x2=46.07 //y2=5.155
r227 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.865 //y=5.155 //x2=46.95 //y2=5.155
r228 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=46.865 //y=5.155 //x2=46.155 //y2=5.155
r229 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.07 //y=5.24 //x2=46.07 //y2=5.155
r230 (  15 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.07 //y=5.24 //x2=46.07 //y2=5.725
r231 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.985 //y=5.155 //x2=46.07 //y2=5.155
r232 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=45.985 //y=5.155 //x2=45.275 //y2=5.155
r233 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=45.19 //y=5.24 //x2=45.275 //y2=5.155
r234 (  7 82 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=45.19 //y=5.24 //x2=45.19 //y2=5.725
r235 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=49.58 //y=3.7 //x2=49.58 //y2=3.7
r236 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=47.73 //y=3.7 //x2=47.73 //y2=3.7
r237 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=47.845 //y=3.7 //x2=47.73 //y2=3.7
r238 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=49.465 //y=3.7 //x2=49.58 //y2=3.7
r239 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=49.465 //y=3.7 //x2=47.845 //y2=3.7
ends PM_TMRDFFRNQNX1\%noxref_10

subckt PM_TMRDFFRNQNX1\%noxref_11 ( 1 2 3 4 5 6 16 23 25 35 36 43 51 57 58 62 \
 63 65 71 72 75 76 77 78 79 80 81 82 83 84 85 86 87 88 90 96 97 98 99 103 104 \
 105 110 112 114 120 121 122 123 124 129 131 133 139 140 150 151 154 163 164 \
 167 175 177 178 179 )
c376 ( 179 0 ) capacitor c=0.023087f //x=41.995 //y=5.02
c377 ( 178 0 ) capacitor c=0.023519f //x=41.115 //y=5.02
c378 ( 177 0 ) capacitor c=0.0224735f //x=40.235 //y=5.02
c379 ( 175 0 ) capacitor c=0.00853354f //x=42.245 //y=0.915
c380 ( 167 0 ) capacitor c=0.0331095f //x=50.35 //y=4.7
c381 ( 164 0 ) capacitor c=0.0279499f //x=50.32 //y=1.915
c382 ( 163 0 ) capacitor c=0.0421676f //x=50.32 //y=2.08
c383 ( 154 0 ) capacitor c=0.0331095f //x=37.4 //y=4.7
c384 ( 151 0 ) capacitor c=0.0279499f //x=37.37 //y=1.915
c385 ( 150 0 ) capacitor c=0.0421676f //x=37.37 //y=2.08
c386 ( 140 0 ) capacitor c=0.0429696f //x=50.885 //y=1.25
c387 ( 139 0 ) capacitor c=0.0192208f //x=50.885 //y=0.905
c388 ( 133 0 ) capacitor c=0.0148884f //x=50.73 //y=1.405
c389 ( 131 0 ) capacitor c=0.0157803f //x=50.73 //y=0.75
c390 ( 129 0 ) capacitor c=0.0295235f //x=50.725 //y=4.79
c391 ( 124 0 ) capacitor c=0.0204188f //x=50.355 //y=1.56
c392 ( 123 0 ) capacitor c=0.0168481f //x=50.355 //y=1.25
c393 ( 122 0 ) capacitor c=0.0174783f //x=50.355 //y=0.905
c394 ( 121 0 ) capacitor c=0.0429696f //x=37.935 //y=1.25
c395 ( 120 0 ) capacitor c=0.0192208f //x=37.935 //y=0.905
c396 ( 114 0 ) capacitor c=0.0148884f //x=37.78 //y=1.405
c397 ( 112 0 ) capacitor c=0.0157803f //x=37.78 //y=0.75
c398 ( 110 0 ) capacitor c=0.0295235f //x=37.775 //y=4.79
c399 ( 105 0 ) capacitor c=0.0204188f //x=37.405 //y=1.56
c400 ( 104 0 ) capacitor c=0.0168481f //x=37.405 //y=1.25
c401 ( 103 0 ) capacitor c=0.0174783f //x=37.405 //y=0.905
c402 ( 99 0 ) capacitor c=0.0557698f //x=27.285 //y=4.79
c403 ( 98 0 ) capacitor c=0.0293157f //x=27.575 //y=4.79
c404 ( 97 0 ) capacitor c=0.0347816f //x=27.24 //y=1.22
c405 ( 96 0 ) capacitor c=0.0187487f //x=27.24 //y=0.875
c406 ( 90 0 ) capacitor c=0.0137055f //x=27.085 //y=1.375
c407 ( 88 0 ) capacitor c=0.0149861f //x=27.085 //y=0.72
c408 ( 87 0 ) capacitor c=0.096037f //x=26.71 //y=1.915
c409 ( 86 0 ) capacitor c=0.0228993f //x=26.71 //y=1.53
c410 ( 85 0 ) capacitor c=0.0234352f //x=26.71 //y=1.22
c411 ( 84 0 ) capacitor c=0.0198724f //x=26.71 //y=0.875
c412 ( 83 0 ) capacitor c=0.15358f //x=50.8 //y=6.02
c413 ( 82 0 ) capacitor c=0.110281f //x=50.36 //y=6.02
c414 ( 81 0 ) capacitor c=0.15358f //x=37.85 //y=6.02
c415 ( 80 0 ) capacitor c=0.110281f //x=37.41 //y=6.02
c416 ( 79 0 ) capacitor c=0.110114f //x=27.65 //y=6.02
c417 ( 78 0 ) capacitor c=0.158956f //x=27.21 //y=6.02
c418 ( 72 0 ) capacitor c=0.00106608f //x=42.14 //y=5.155
c419 ( 71 0 ) capacitor c=0.00207162f //x=41.26 //y=5.155
c420 ( 65 0 ) capacitor c=0.0690311f //x=50.32 //y=2.08
c421 ( 63 0 ) capacitor c=0.00453889f //x=50.32 //y=4.535
c422 ( 62 0 ) capacitor c=0.106357f //x=42.92 //y=4.07
c423 ( 58 0 ) capacitor c=0.00398962f //x=42.52 //y=1.665
c424 ( 57 0 ) capacitor c=0.0137288f //x=42.835 //y=1.665
c425 ( 51 0 ) capacitor c=0.0283082f //x=42.835 //y=5.155
c426 ( 43 0 ) capacitor c=0.0176454f //x=42.055 //y=5.155
c427 ( 36 0 ) capacitor c=0.00332903f //x=40.465 //y=5.155
c428 ( 35 0 ) capacitor c=0.014837f //x=41.175 //y=5.155
c429 ( 25 0 ) capacitor c=0.0680284f //x=37.37 //y=2.08
c430 ( 23 0 ) capacitor c=0.00453889f //x=37.37 //y=4.535
c431 ( 16 0 ) capacitor c=0.100832f //x=27.01 //y=2.08
c432 ( 6 0 ) capacitor c=0.00554824f //x=43.035 //y=4.07
c433 ( 5 0 ) capacitor c=0.124977f //x=50.205 //y=4.07
c434 ( 4 0 ) capacitor c=0.00557292f //x=37.485 //y=4.07
c435 ( 3 0 ) capacitor c=0.0725278f //x=42.805 //y=4.07
c436 ( 2 0 ) capacitor c=0.0102374f //x=27.125 //y=4.07
c437 ( 1 0 ) capacitor c=0.151078f //x=37.255 //y=4.07
r438 (  169 170 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=50.35 //y=4.79 //x2=50.35 //y2=4.865
r439 (  167 169 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=50.35 //y=4.7 //x2=50.35 //y2=4.79
r440 (  163 164 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=50.32 //y=2.08 //x2=50.32 //y2=1.915
r441 (  156 157 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=37.4 //y=4.79 //x2=37.4 //y2=4.865
r442 (  154 156 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=37.4 //y=4.7 //x2=37.4 //y2=4.79
r443 (  150 151 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=37.37 //y=2.08 //x2=37.37 //y2=1.915
r444 (  140 174 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.885 //y=1.25 //x2=50.845 //y2=1.405
r445 (  139 173 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.885 //y=0.905 //x2=50.845 //y2=0.75
r446 (  139 140 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=50.885 //y=0.905 //x2=50.885 //y2=1.25
r447 (  134 172 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.51 //y=1.405 //x2=50.395 //y2=1.405
r448 (  133 174 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.73 //y=1.405 //x2=50.845 //y2=1.405
r449 (  132 171 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.51 //y=0.75 //x2=50.395 //y2=0.75
r450 (  131 173 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.73 //y=0.75 //x2=50.845 //y2=0.75
r451 (  131 132 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=50.73 //y=0.75 //x2=50.51 //y2=0.75
r452 (  130 169 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=50.485 //y=4.79 //x2=50.35 //y2=4.79
r453 (  129 136 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=50.725 //y=4.79 //x2=50.8 //y2=4.865
r454 (  129 130 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=50.725 //y=4.79 //x2=50.485 //y2=4.79
r455 (  124 172 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.355 //y=1.56 //x2=50.395 //y2=1.405
r456 (  124 164 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=50.355 //y=1.56 //x2=50.355 //y2=1.915
r457 (  123 172 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.355 //y=1.25 //x2=50.395 //y2=1.405
r458 (  122 171 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.355 //y=0.905 //x2=50.395 //y2=0.75
r459 (  122 123 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=50.355 //y=0.905 //x2=50.355 //y2=1.25
r460 (  121 161 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.935 //y=1.25 //x2=37.895 //y2=1.405
r461 (  120 160 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.935 //y=0.905 //x2=37.895 //y2=0.75
r462 (  120 121 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=37.935 //y=0.905 //x2=37.935 //y2=1.25
r463 (  115 159 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.56 //y=1.405 //x2=37.445 //y2=1.405
r464 (  114 161 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.78 //y=1.405 //x2=37.895 //y2=1.405
r465 (  113 158 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.56 //y=0.75 //x2=37.445 //y2=0.75
r466 (  112 160 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=37.78 //y=0.75 //x2=37.895 //y2=0.75
r467 (  112 113 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=37.78 //y=0.75 //x2=37.56 //y2=0.75
r468 (  111 156 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=37.535 //y=4.79 //x2=37.4 //y2=4.79
r469 (  110 117 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=37.775 //y=4.79 //x2=37.85 //y2=4.865
r470 (  110 111 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=37.775 //y=4.79 //x2=37.535 //y2=4.79
r471 (  105 159 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.405 //y=1.56 //x2=37.445 //y2=1.405
r472 (  105 151 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=37.405 //y=1.56 //x2=37.405 //y2=1.915
r473 (  104 159 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.405 //y=1.25 //x2=37.445 //y2=1.405
r474 (  103 158 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=37.405 //y=0.905 //x2=37.445 //y2=0.75
r475 (  103 104 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=37.405 //y=0.905 //x2=37.405 //y2=1.25
r476 (  98 100 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=27.575 //y=4.79 //x2=27.65 //y2=4.865
r477 (  98 99 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=27.575 //y=4.79 //x2=27.285 //y2=4.79
r478 (  97 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.24 //y=1.22 //x2=27.2 //y2=1.375
r479 (  96 147 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.24 //y=0.875 //x2=27.2 //y2=0.72
r480 (  96 97 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=27.24 //y=0.875 //x2=27.24 //y2=1.22
r481 (  93 99 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=27.21 //y=4.865 //x2=27.285 //y2=4.79
r482 (  93 146 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=27.21 //y=4.865 //x2=27.01 //y2=4.7
r483 (  91 142 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.865 //y=1.375 //x2=26.75 //y2=1.375
r484 (  90 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.085 //y=1.375 //x2=27.2 //y2=1.375
r485 (  89 141 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.865 //y=0.72 //x2=26.75 //y2=0.72
r486 (  88 147 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.085 //y=0.72 //x2=27.2 //y2=0.72
r487 (  88 89 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=27.085 //y=0.72 //x2=26.865 //y2=0.72
r488 (  87 144 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=26.71 //y=1.915 //x2=27.01 //y2=2.08
r489 (  86 142 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.71 //y=1.53 //x2=26.75 //y2=1.375
r490 (  86 87 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=26.71 //y=1.53 //x2=26.71 //y2=1.915
r491 (  85 142 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.71 //y=1.22 //x2=26.75 //y2=1.375
r492 (  84 141 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.71 //y=0.875 //x2=26.75 //y2=0.72
r493 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=26.71 //y=0.875 //x2=26.71 //y2=1.22
r494 (  83 136 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=50.8 //y=6.02 //x2=50.8 //y2=4.865
r495 (  82 170 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=50.36 //y=6.02 //x2=50.36 //y2=4.865
r496 (  81 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=37.85 //y=6.02 //x2=37.85 //y2=4.865
r497 (  80 157 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=37.41 //y=6.02 //x2=37.41 //y2=4.865
r498 (  79 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=27.65 //y=6.02 //x2=27.65 //y2=4.865
r499 (  78 93 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=27.21 //y=6.02 //x2=27.21 //y2=4.865
r500 (  77 133 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=50.62 //y=1.405 //x2=50.73 //y2=1.405
r501 (  77 134 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=50.62 //y=1.405 //x2=50.51 //y2=1.405
r502 (  76 114 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=37.67 //y=1.405 //x2=37.78 //y2=1.405
r503 (  76 115 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=37.67 //y=1.405 //x2=37.56 //y2=1.405
r504 (  75 90 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=26.975 //y=1.375 //x2=27.085 //y2=1.375
r505 (  75 91 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=26.975 //y=1.375 //x2=26.865 //y2=1.375
r506 (  74 167 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=50.35 //y=4.7 //x2=50.35 //y2=4.7
r507 (  70 154 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=37.4 //y=4.7 //x2=37.4 //y2=4.7
r508 (  65 163 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=50.32 //y=2.08 //x2=50.32 //y2=2.08
r509 (  65 68 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=50.32 //y=2.08 //x2=50.32 //y2=4.07
r510 (  63 74 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=50.32 //y=4.535 //x2=50.335 //y2=4.7
r511 (  63 68 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=50.32 //y=4.535 //x2=50.32 //y2=4.07
r512 (  60 62 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=42.92 //y=5.07 //x2=42.92 //y2=4.07
r513 (  59 62 ) resistor r=158.802 //w=0.187 //l=2.32 //layer=li \
 //thickness=0.1 //x=42.92 //y=1.75 //x2=42.92 //y2=4.07
r514 (  57 59 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.835 //y=1.665 //x2=42.92 //y2=1.75
r515 (  57 58 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=42.835 //y=1.665 //x2=42.52 //y2=1.665
r516 (  53 58 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.435 //y=1.58 //x2=42.52 //y2=1.665
r517 (  53 175 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=42.435 //y=1.58 //x2=42.435 //y2=1.01
r518 (  52 72 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.225 //y=5.155 //x2=42.14 //y2=5.155
r519 (  51 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.835 //y=5.155 //x2=42.92 //y2=5.07
r520 (  51 52 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=42.835 //y=5.155 //x2=42.225 //y2=5.155
r521 (  45 72 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.14 //y=5.24 //x2=42.14 //y2=5.155
r522 (  45 179 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=42.14 //y=5.24 //x2=42.14 //y2=5.725
r523 (  44 71 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.345 //y=5.155 //x2=41.26 //y2=5.155
r524 (  43 72 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.055 //y=5.155 //x2=42.14 //y2=5.155
r525 (  43 44 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=42.055 //y=5.155 //x2=41.345 //y2=5.155
r526 (  37 71 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.26 //y=5.24 //x2=41.26 //y2=5.155
r527 (  37 178 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=41.26 //y=5.24 //x2=41.26 //y2=5.725
r528 (  35 71 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.175 //y=5.155 //x2=41.26 //y2=5.155
r529 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=41.175 //y=5.155 //x2=40.465 //y2=5.155
r530 (  29 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=40.38 //y=5.24 //x2=40.465 //y2=5.155
r531 (  29 177 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=40.38 //y=5.24 //x2=40.38 //y2=5.725
r532 (  25 150 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=37.37 //y=2.08 //x2=37.37 //y2=2.08
r533 (  25 28 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=37.37 //y=2.08 //x2=37.37 //y2=4.07
r534 (  23 70 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=37.37 //y=4.535 //x2=37.385 //y2=4.7
r535 (  23 28 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=37.37 //y=4.535 //x2=37.37 //y2=4.07
r536 (  21 146 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=27.01 //y=4.7 //x2=27.01 //y2=4.7
r537 (  19 21 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=27.01 //y=4.07 //x2=27.01 //y2=4.7
r538 (  16 144 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=27.01 //y=2.08 //x2=27.01 //y2=2.08
r539 (  16 19 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=27.01 //y=2.08 //x2=27.01 //y2=4.07
r540 (  14 68 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=50.32 //y=4.07 //x2=50.32 //y2=4.07
r541 (  12 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=42.92 //y=4.07 //x2=42.92 //y2=4.07
r542 (  10 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=37.37 //y=4.07 //x2=37.37 //y2=4.07
r543 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=27.01 //y=4.07 //x2=27.01 //y2=4.07
r544 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=43.035 //y=4.07 //x2=42.92 //y2=4.07
r545 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=50.205 //y=4.07 //x2=50.32 //y2=4.07
r546 (  5 6 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=50.205 //y=4.07 //x2=43.035 //y2=4.07
r547 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=37.485 //y=4.07 //x2=37.37 //y2=4.07
r548 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=42.805 //y=4.07 //x2=42.92 //y2=4.07
r549 (  3 4 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=42.805 //y=4.07 //x2=37.485 //y2=4.07
r550 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=27.125 //y=4.07 //x2=27.01 //y2=4.07
r551 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=37.255 //y=4.07 //x2=37.37 //y2=4.07
r552 (  1 2 ) resistor r=9.66603 //w=0.131 //l=10.13 //layer=m1 \
 //thickness=0.36 //x=37.255 //y=4.07 //x2=27.125 //y2=4.07
ends PM_TMRDFFRNQNX1\%noxref_11

subckt PM_TMRDFFRNQNX1\%D ( 1 2 3 4 11 12 14 23 31 38 39 40 41 42 43 44 45 46 \
 47 48 49 51 57 58 59 60 61 66 67 68 70 76 77 78 79 80 85 86 87 89 95 96 97 98 \
 99 107 118 129 )
c368 ( 129 0 ) capacitor c=0.0335551f //x=58.83 //y=4.7
c369 ( 118 0 ) capacitor c=0.0335551f //x=32.93 //y=4.7
c370 ( 107 0 ) capacitor c=0.0335551f //x=7.03 //y=4.7
c371 ( 99 0 ) capacitor c=0.0245352f //x=59.165 //y=4.79
c372 ( 98 0 ) capacitor c=0.0825763f //x=58.92 //y=1.915
c373 ( 97 0 ) capacitor c=0.0170266f //x=58.92 //y=1.45
c374 ( 96 0 ) capacitor c=0.018609f //x=58.92 //y=1.22
c375 ( 95 0 ) capacitor c=0.0187309f //x=58.92 //y=0.91
c376 ( 89 0 ) capacitor c=0.014725f //x=58.765 //y=1.375
c377 ( 87 0 ) capacitor c=0.0146567f //x=58.765 //y=0.755
c378 ( 86 0 ) capacitor c=0.0335408f //x=58.395 //y=1.22
c379 ( 85 0 ) capacitor c=0.0173761f //x=58.395 //y=0.91
c380 ( 80 0 ) capacitor c=0.0245352f //x=33.265 //y=4.79
c381 ( 79 0 ) capacitor c=0.0825763f //x=33.02 //y=1.915
c382 ( 78 0 ) capacitor c=0.0170266f //x=33.02 //y=1.45
c383 ( 77 0 ) capacitor c=0.018609f //x=33.02 //y=1.22
c384 ( 76 0 ) capacitor c=0.0187309f //x=33.02 //y=0.91
c385 ( 70 0 ) capacitor c=0.014725f //x=32.865 //y=1.375
c386 ( 68 0 ) capacitor c=0.0146567f //x=32.865 //y=0.755
c387 ( 67 0 ) capacitor c=0.0335408f //x=32.495 //y=1.22
c388 ( 66 0 ) capacitor c=0.0173761f //x=32.495 //y=0.91
c389 ( 61 0 ) capacitor c=0.0245352f //x=7.365 //y=4.79
c390 ( 60 0 ) capacitor c=0.0826363f //x=7.12 //y=1.915
c391 ( 59 0 ) capacitor c=0.0170266f //x=7.12 //y=1.45
c392 ( 58 0 ) capacitor c=0.018609f //x=7.12 //y=1.22
c393 ( 57 0 ) capacitor c=0.0187309f //x=7.12 //y=0.91
c394 ( 51 0 ) capacitor c=0.014725f //x=6.965 //y=1.375
c395 ( 49 0 ) capacitor c=0.0146567f //x=6.965 //y=0.755
c396 ( 48 0 ) capacitor c=0.0335408f //x=6.595 //y=1.22
c397 ( 47 0 ) capacitor c=0.0173761f //x=6.595 //y=0.91
c398 ( 46 0 ) capacitor c=0.110114f //x=59.24 //y=6.02
c399 ( 45 0 ) capacitor c=0.11012f //x=58.8 //y=6.02
c400 ( 44 0 ) capacitor c=0.110114f //x=33.34 //y=6.02
c401 ( 43 0 ) capacitor c=0.11012f //x=32.9 //y=6.02
c402 ( 42 0 ) capacitor c=0.110114f //x=7.44 //y=6.02
c403 ( 41 0 ) capacitor c=0.11012f //x=7 //y=6.02
c404 ( 31 0 ) capacitor c=0.0879663f //x=58.83 //y=2.08
c405 ( 23 0 ) capacitor c=0.0879663f //x=32.93 //y=2.08
c406 ( 14 0 ) capacitor c=0.0930795f //x=7.03 //y=2.08
c407 ( 4 0 ) capacitor c=0.00558494f //x=33.045 //y=2.59
c408 ( 3 0 ) capacitor c=0.34213f //x=58.715 //y=2.59
c409 ( 2 0 ) capacitor c=0.0159757f //x=7.145 //y=2.59
c410 ( 1 0 ) capacitor c=0.411825f //x=32.815 //y=2.59
r411 (  131 132 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=58.83 //y=4.79 //x2=58.83 //y2=4.865
r412 (  129 131 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=58.83 //y=4.7 //x2=58.83 //y2=4.79
r413 (  120 121 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=32.93 //y=4.79 //x2=32.93 //y2=4.865
r414 (  118 120 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=32.93 //y=4.7 //x2=32.93 //y2=4.79
r415 (  109 110 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=7.03 //y=4.79 //x2=7.03 //y2=4.865
r416 (  107 109 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=7.03 //y=4.7 //x2=7.03 //y2=4.79
r417 (  100 131 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=58.965 //y=4.79 //x2=58.83 //y2=4.79
r418 (  99 101 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=59.165 //y=4.79 //x2=59.24 //y2=4.865
r419 (  99 100 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=59.165 //y=4.79 //x2=58.965 //y2=4.79
r420 (  98 136 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=58.92 //y=1.915 //x2=58.845 //y2=2.08
r421 (  97 134 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=58.92 //y=1.45 //x2=58.88 //y2=1.375
r422 (  97 98 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=58.92 //y=1.45 //x2=58.92 //y2=1.915
r423 (  96 134 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.92 //y=1.22 //x2=58.88 //y2=1.375
r424 (  95 133 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.92 //y=0.91 //x2=58.88 //y2=0.755
r425 (  95 96 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=58.92 //y=0.91 //x2=58.92 //y2=1.22
r426 (  90 127 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.55 //y=1.375 //x2=58.435 //y2=1.375
r427 (  89 134 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.765 //y=1.375 //x2=58.88 //y2=1.375
r428 (  88 126 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.55 //y=0.755 //x2=58.435 //y2=0.755
r429 (  87 133 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.765 //y=0.755 //x2=58.88 //y2=0.755
r430 (  87 88 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=58.765 //y=0.755 //x2=58.55 //y2=0.755
r431 (  86 127 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.395 //y=1.22 //x2=58.435 //y2=1.375
r432 (  85 126 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.395 //y=0.91 //x2=58.435 //y2=0.755
r433 (  85 86 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=58.395 //y=0.91 //x2=58.395 //y2=1.22
r434 (  81 120 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=33.065 //y=4.79 //x2=32.93 //y2=4.79
r435 (  80 82 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=33.265 //y=4.79 //x2=33.34 //y2=4.865
r436 (  80 81 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=33.265 //y=4.79 //x2=33.065 //y2=4.79
r437 (  79 125 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=33.02 //y=1.915 //x2=32.945 //y2=2.08
r438 (  78 123 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=33.02 //y=1.45 //x2=32.98 //y2=1.375
r439 (  78 79 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=33.02 //y=1.45 //x2=33.02 //y2=1.915
r440 (  77 123 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.02 //y=1.22 //x2=32.98 //y2=1.375
r441 (  76 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.02 //y=0.91 //x2=32.98 //y2=0.755
r442 (  76 77 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=33.02 //y=0.91 //x2=33.02 //y2=1.22
r443 (  71 116 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.65 //y=1.375 //x2=32.535 //y2=1.375
r444 (  70 123 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.865 //y=1.375 //x2=32.98 //y2=1.375
r445 (  69 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.65 //y=0.755 //x2=32.535 //y2=0.755
r446 (  68 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=32.865 //y=0.755 //x2=32.98 //y2=0.755
r447 (  68 69 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=32.865 //y=0.755 //x2=32.65 //y2=0.755
r448 (  67 116 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.495 //y=1.22 //x2=32.535 //y2=1.375
r449 (  66 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=32.495 //y=0.91 //x2=32.535 //y2=0.755
r450 (  66 67 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=32.495 //y=0.91 //x2=32.495 //y2=1.22
r451 (  62 109 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=7.165 //y=4.79 //x2=7.03 //y2=4.79
r452 (  61 63 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.365 //y=4.79 //x2=7.44 //y2=4.865
r453 (  61 62 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=7.365 //y=4.79 //x2=7.165 //y2=4.79
r454 (  60 114 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.915 //x2=7.045 //y2=2.08
r455 (  59 112 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.45 //x2=7.08 //y2=1.375
r456 (  59 60 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.45 //x2=7.12 //y2=1.915
r457 (  58 112 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.22 //x2=7.08 //y2=1.375
r458 (  57 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.12 //y=0.91 //x2=7.08 //y2=0.755
r459 (  57 58 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=7.12 //y=0.91 //x2=7.12 //y2=1.22
r460 (  52 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.75 //y=1.375 //x2=6.635 //y2=1.375
r461 (  51 112 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.965 //y=1.375 //x2=7.08 //y2=1.375
r462 (  50 104 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.75 //y=0.755 //x2=6.635 //y2=0.755
r463 (  49 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.965 //y=0.755 //x2=7.08 //y2=0.755
r464 (  49 50 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=6.965 //y=0.755 //x2=6.75 //y2=0.755
r465 (  48 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.595 //y=1.22 //x2=6.635 //y2=1.375
r466 (  47 104 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.595 //y=0.91 //x2=6.635 //y2=0.755
r467 (  47 48 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=6.595 //y=0.91 //x2=6.595 //y2=1.22
r468 (  46 101 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.24 //y=6.02 //x2=59.24 //y2=4.865
r469 (  45 132 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=58.8 //y=6.02 //x2=58.8 //y2=4.865
r470 (  44 82 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=33.34 //y=6.02 //x2=33.34 //y2=4.865
r471 (  43 121 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=32.9 //y=6.02 //x2=32.9 //y2=4.865
r472 (  42 63 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.44 //y=6.02 //x2=7.44 //y2=4.865
r473 (  41 110 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7 //y=6.02 //x2=7 //y2=4.865
r474 (  40 89 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=58.657 //y=1.375 //x2=58.765 //y2=1.375
r475 (  40 90 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=58.657 //y=1.375 //x2=58.55 //y2=1.375
r476 (  39 70 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=32.757 //y=1.375 //x2=32.865 //y2=1.375
r477 (  39 71 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=32.757 //y=1.375 //x2=32.65 //y2=1.375
r478 (  38 51 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=6.857 //y=1.375 //x2=6.965 //y2=1.375
r479 (  38 52 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=6.857 //y=1.375 //x2=6.75 //y2=1.375
r480 (  36 129 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=58.83 //y=4.7 //x2=58.83 //y2=4.7
r481 (  34 36 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=58.83 //y=2.59 //x2=58.83 //y2=4.7
r482 (  31 136 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=58.83 //y=2.08 //x2=58.83 //y2=2.08
r483 (  31 34 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=58.83 //y=2.08 //x2=58.83 //y2=2.59
r484 (  28 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=32.93 //y=4.7 //x2=32.93 //y2=4.7
r485 (  26 28 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=32.93 //y=2.59 //x2=32.93 //y2=4.7
r486 (  23 125 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=32.93 //y=2.08 //x2=32.93 //y2=2.08
r487 (  23 26 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=32.93 //y=2.08 //x2=32.93 //y2=2.59
r488 (  20 107 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.03 //y=4.7 //x2=7.03 //y2=4.7
r489 (  14 114 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.03 //y=2.08 //x2=7.03 //y2=2.08
r490 (  12 20 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=7.03 //y=2.96 //x2=7.03 //y2=4.7
r491 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=7.03 //y=2.59 //x2=7.03 //y2=2.96
r492 (  11 14 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=7.03 //y=2.59 //x2=7.03 //y2=2.08
r493 (  10 34 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=58.83 //y=2.59 //x2=58.83 //y2=2.59
r494 (  8 26 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=32.93 //y=2.59 //x2=32.93 //y2=2.59
r495 (  6 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.03 //y=2.59 //x2=7.03 //y2=2.59
r496 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=33.045 //y=2.59 //x2=32.93 //y2=2.59
r497 (  3 10 ) resistor r=0.0738079 //w=0.207 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=58.715 //y=2.59 //x2=58.83 //y2=2.59
r498 (  3 4 ) resistor r=24.4943 //w=0.131 //l=25.67 //layer=m1 \
 //thickness=0.36 //x=58.715 //y=2.59 //x2=33.045 //y2=2.59
r499 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.145 //y=2.59 //x2=7.03 //y2=2.59
r500 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=32.815 //y=2.59 //x2=32.93 //y2=2.59
r501 (  1 2 ) resistor r=24.4943 //w=0.131 //l=25.67 //layer=m1 \
 //thickness=0.36 //x=32.815 //y=2.59 //x2=7.145 //y2=2.59
ends PM_TMRDFFRNQNX1\%D

subckt PM_TMRDFFRNQNX1\%CLK ( 1 2 3 4 5 6 7 8 9 10 23 24 25 26 27 28 29 30 31 \
 32 33 34 35 36 37 38 40 52 62 72 81 90 97 98 99 100 101 102 103 104 105 106 \
 107 108 109 110 111 112 113 114 115 116 117 119 125 126 127 128 129 134 135 \
 136 138 144 145 146 147 148 153 154 155 157 163 164 165 166 167 172 173 174 \
 176 182 183 184 185 186 191 192 193 195 201 202 203 204 205 210 211 212 214 \
 220 221 222 223 224 232 243 254 265 276 287 )
c785 ( 287 0 ) capacitor c=0.0334842f //x=66.97 //y=4.7
c786 ( 276 0 ) capacitor c=0.0334842f //x=54.02 //y=4.7
c787 ( 265 0 ) capacitor c=0.0334842f //x=41.07 //y=4.7
c788 ( 254 0 ) capacitor c=0.0334842f //x=28.12 //y=4.7
c789 ( 243 0 ) capacitor c=0.0334842f //x=15.17 //y=4.7
c790 ( 232 0 ) capacitor c=0.0334842f //x=2.22 //y=4.7
c791 ( 224 0 ) capacitor c=0.0249231f //x=67.305 //y=4.79
c792 ( 223 0 ) capacitor c=0.0825763f //x=67.06 //y=1.915
c793 ( 222 0 ) capacitor c=0.0170266f //x=67.06 //y=1.45
c794 ( 221 0 ) capacitor c=0.018609f //x=67.06 //y=1.22
c795 ( 220 0 ) capacitor c=0.0187309f //x=67.06 //y=0.91
c796 ( 214 0 ) capacitor c=0.014725f //x=66.905 //y=1.375
c797 ( 212 0 ) capacitor c=0.0146567f //x=66.905 //y=0.755
c798 ( 211 0 ) capacitor c=0.0335408f //x=66.535 //y=1.22
c799 ( 210 0 ) capacitor c=0.0173761f //x=66.535 //y=0.91
c800 ( 205 0 ) capacitor c=0.0245352f //x=54.355 //y=4.79
c801 ( 204 0 ) capacitor c=0.0825763f //x=54.11 //y=1.915
c802 ( 203 0 ) capacitor c=0.0170266f //x=54.11 //y=1.45
c803 ( 202 0 ) capacitor c=0.018609f //x=54.11 //y=1.22
c804 ( 201 0 ) capacitor c=0.0187309f //x=54.11 //y=0.91
c805 ( 195 0 ) capacitor c=0.014725f //x=53.955 //y=1.375
c806 ( 193 0 ) capacitor c=0.0146567f //x=53.955 //y=0.755
c807 ( 192 0 ) capacitor c=0.0335408f //x=53.585 //y=1.22
c808 ( 191 0 ) capacitor c=0.0173761f //x=53.585 //y=0.91
c809 ( 186 0 ) capacitor c=0.0245352f //x=41.405 //y=4.79
c810 ( 185 0 ) capacitor c=0.0825763f //x=41.16 //y=1.915
c811 ( 184 0 ) capacitor c=0.0170266f //x=41.16 //y=1.45
c812 ( 183 0 ) capacitor c=0.018609f //x=41.16 //y=1.22
c813 ( 182 0 ) capacitor c=0.0187309f //x=41.16 //y=0.91
c814 ( 176 0 ) capacitor c=0.014725f //x=41.005 //y=1.375
c815 ( 174 0 ) capacitor c=0.0146567f //x=41.005 //y=0.755
c816 ( 173 0 ) capacitor c=0.0335408f //x=40.635 //y=1.22
c817 ( 172 0 ) capacitor c=0.0173761f //x=40.635 //y=0.91
c818 ( 167 0 ) capacitor c=0.0245352f //x=28.455 //y=4.79
c819 ( 166 0 ) capacitor c=0.0825763f //x=28.21 //y=1.915
c820 ( 165 0 ) capacitor c=0.0170266f //x=28.21 //y=1.45
c821 ( 164 0 ) capacitor c=0.018609f //x=28.21 //y=1.22
c822 ( 163 0 ) capacitor c=0.0187309f //x=28.21 //y=0.91
c823 ( 157 0 ) capacitor c=0.014725f //x=28.055 //y=1.375
c824 ( 155 0 ) capacitor c=0.0146567f //x=28.055 //y=0.755
c825 ( 154 0 ) capacitor c=0.0335408f //x=27.685 //y=1.22
c826 ( 153 0 ) capacitor c=0.0173761f //x=27.685 //y=0.91
c827 ( 148 0 ) capacitor c=0.0245352f //x=15.505 //y=4.79
c828 ( 147 0 ) capacitor c=0.0825763f //x=15.26 //y=1.915
c829 ( 146 0 ) capacitor c=0.0170266f //x=15.26 //y=1.45
c830 ( 145 0 ) capacitor c=0.018609f //x=15.26 //y=1.22
c831 ( 144 0 ) capacitor c=0.0187309f //x=15.26 //y=0.91
c832 ( 138 0 ) capacitor c=0.014725f //x=15.105 //y=1.375
c833 ( 136 0 ) capacitor c=0.0146567f //x=15.105 //y=0.755
c834 ( 135 0 ) capacitor c=0.0335408f //x=14.735 //y=1.22
c835 ( 134 0 ) capacitor c=0.0173761f //x=14.735 //y=0.91
c836 ( 129 0 ) capacitor c=0.0245352f //x=2.555 //y=4.79
c837 ( 128 0 ) capacitor c=0.0850619f //x=2.31 //y=1.915
c838 ( 127 0 ) capacitor c=0.0170266f //x=2.31 //y=1.45
c839 ( 126 0 ) capacitor c=0.018609f //x=2.31 //y=1.22
c840 ( 125 0 ) capacitor c=0.0187309f //x=2.31 //y=0.91
c841 ( 119 0 ) capacitor c=0.014725f //x=2.155 //y=1.375
c842 ( 117 0 ) capacitor c=0.0146567f //x=2.155 //y=0.755
c843 ( 116 0 ) capacitor c=0.0335408f //x=1.785 //y=1.22
c844 ( 115 0 ) capacitor c=0.0173761f //x=1.785 //y=0.91
c845 ( 114 0 ) capacitor c=0.110114f //x=67.38 //y=6.02
c846 ( 113 0 ) capacitor c=0.11012f //x=66.94 //y=6.02
c847 ( 112 0 ) capacitor c=0.110114f //x=54.43 //y=6.02
c848 ( 111 0 ) capacitor c=0.11012f //x=53.99 //y=6.02
c849 ( 110 0 ) capacitor c=0.110114f //x=41.48 //y=6.02
c850 ( 109 0 ) capacitor c=0.11012f //x=41.04 //y=6.02
c851 ( 108 0 ) capacitor c=0.110114f //x=28.53 //y=6.02
c852 ( 107 0 ) capacitor c=0.11012f //x=28.09 //y=6.02
c853 ( 106 0 ) capacitor c=0.110114f //x=15.58 //y=6.02
c854 ( 105 0 ) capacitor c=0.11012f //x=15.14 //y=6.02
c855 ( 104 0 ) capacitor c=0.110114f //x=2.63 //y=6.02
c856 ( 103 0 ) capacitor c=0.11012f //x=2.19 //y=6.02
c857 ( 90 0 ) capacitor c=0.0906039f //x=66.97 //y=2.08
c858 ( 81 0 ) capacitor c=0.0901246f //x=54.02 //y=2.08
c859 ( 72 0 ) capacitor c=0.0899873f //x=41.07 //y=2.08
c860 ( 62 0 ) capacitor c=0.0921514f //x=28.12 //y=2.08
c861 ( 52 0 ) capacitor c=0.0926307f //x=15.17 //y=2.08
c862 ( 40 0 ) capacitor c=0.100158f //x=2.22 //y=2.08
c863 ( 10 0 ) capacitor c=0.00697397f //x=54.135 //y=4.44
c864 ( 9 0 ) capacitor c=0.301662f //x=66.855 //y=4.44
c865 ( 8 0 ) capacitor c=0.00697397f //x=41.185 //y=4.44
c866 ( 7 0 ) capacitor c=0.301789f //x=53.905 //y=4.44
c867 ( 6 0 ) capacitor c=0.00697397f //x=28.235 //y=4.44
c868 ( 5 0 ) capacitor c=0.286372f //x=40.955 //y=4.44
c869 ( 4 0 ) capacitor c=0.00697397f //x=15.285 //y=4.44
c870 ( 3 0 ) capacitor c=0.307121f //x=28.005 //y=4.44
c871 ( 2 0 ) capacitor c=0.0154455f //x=2.335 //y=4.44
c872 ( 1 0 ) capacitor c=0.286372f //x=15.055 //y=4.44
r873 (  289 290 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=66.97 //y=4.79 //x2=66.97 //y2=4.865
r874 (  287 289 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=66.97 //y=4.7 //x2=66.97 //y2=4.79
r875 (  278 279 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=54.02 //y=4.79 //x2=54.02 //y2=4.865
r876 (  276 278 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=54.02 //y=4.7 //x2=54.02 //y2=4.79
r877 (  267 268 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=41.07 //y=4.79 //x2=41.07 //y2=4.865
r878 (  265 267 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=41.07 //y=4.7 //x2=41.07 //y2=4.79
r879 (  256 257 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=28.12 //y=4.79 //x2=28.12 //y2=4.865
r880 (  254 256 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=28.12 //y=4.7 //x2=28.12 //y2=4.79
r881 (  245 246 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=15.17 //y=4.79 //x2=15.17 //y2=4.865
r882 (  243 245 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=15.17 //y=4.7 //x2=15.17 //y2=4.79
r883 (  234 235 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.79 //x2=2.22 //y2=4.865
r884 (  232 234 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.7 //x2=2.22 //y2=4.79
r885 (  225 289 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=67.105 //y=4.79 //x2=66.97 //y2=4.79
r886 (  224 226 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=67.305 //y=4.79 //x2=67.38 //y2=4.865
r887 (  224 225 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=67.305 //y=4.79 //x2=67.105 //y2=4.79
r888 (  223 294 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=67.06 //y=1.915 //x2=66.985 //y2=2.08
r889 (  222 292 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=67.06 //y=1.45 //x2=67.02 //y2=1.375
r890 (  222 223 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=67.06 //y=1.45 //x2=67.06 //y2=1.915
r891 (  221 292 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=67.06 //y=1.22 //x2=67.02 //y2=1.375
r892 (  220 291 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=67.06 //y=0.91 //x2=67.02 //y2=0.755
r893 (  220 221 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=67.06 //y=0.91 //x2=67.06 //y2=1.22
r894 (  215 285 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.69 //y=1.375 //x2=66.575 //y2=1.375
r895 (  214 292 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.905 //y=1.375 //x2=67.02 //y2=1.375
r896 (  213 284 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.69 //y=0.755 //x2=66.575 //y2=0.755
r897 (  212 291 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.905 //y=0.755 //x2=67.02 //y2=0.755
r898 (  212 213 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=66.905 //y=0.755 //x2=66.69 //y2=0.755
r899 (  211 285 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.535 //y=1.22 //x2=66.575 //y2=1.375
r900 (  210 284 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.535 //y=0.91 //x2=66.575 //y2=0.755
r901 (  210 211 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=66.535 //y=0.91 //x2=66.535 //y2=1.22
r902 (  206 278 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=54.155 //y=4.79 //x2=54.02 //y2=4.79
r903 (  205 207 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=54.355 //y=4.79 //x2=54.43 //y2=4.865
r904 (  205 206 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=54.355 //y=4.79 //x2=54.155 //y2=4.79
r905 (  204 283 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=54.11 //y=1.915 //x2=54.035 //y2=2.08
r906 (  203 281 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=54.11 //y=1.45 //x2=54.07 //y2=1.375
r907 (  203 204 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=54.11 //y=1.45 //x2=54.11 //y2=1.915
r908 (  202 281 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.11 //y=1.22 //x2=54.07 //y2=1.375
r909 (  201 280 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.11 //y=0.91 //x2=54.07 //y2=0.755
r910 (  201 202 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=54.11 //y=0.91 //x2=54.11 //y2=1.22
r911 (  196 274 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.74 //y=1.375 //x2=53.625 //y2=1.375
r912 (  195 281 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.955 //y=1.375 //x2=54.07 //y2=1.375
r913 (  194 273 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.74 //y=0.755 //x2=53.625 //y2=0.755
r914 (  193 280 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.955 //y=0.755 //x2=54.07 //y2=0.755
r915 (  193 194 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=53.955 //y=0.755 //x2=53.74 //y2=0.755
r916 (  192 274 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.585 //y=1.22 //x2=53.625 //y2=1.375
r917 (  191 273 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.585 //y=0.91 //x2=53.625 //y2=0.755
r918 (  191 192 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=53.585 //y=0.91 //x2=53.585 //y2=1.22
r919 (  187 267 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=41.205 //y=4.79 //x2=41.07 //y2=4.79
r920 (  186 188 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=41.405 //y=4.79 //x2=41.48 //y2=4.865
r921 (  186 187 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=41.405 //y=4.79 //x2=41.205 //y2=4.79
r922 (  185 272 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=41.16 //y=1.915 //x2=41.085 //y2=2.08
r923 (  184 270 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=41.16 //y=1.45 //x2=41.12 //y2=1.375
r924 (  184 185 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=41.16 //y=1.45 //x2=41.16 //y2=1.915
r925 (  183 270 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.16 //y=1.22 //x2=41.12 //y2=1.375
r926 (  182 269 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.16 //y=0.91 //x2=41.12 //y2=0.755
r927 (  182 183 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=41.16 //y=0.91 //x2=41.16 //y2=1.22
r928 (  177 263 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.79 //y=1.375 //x2=40.675 //y2=1.375
r929 (  176 270 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.005 //y=1.375 //x2=41.12 //y2=1.375
r930 (  175 262 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=40.79 //y=0.755 //x2=40.675 //y2=0.755
r931 (  174 269 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.005 //y=0.755 //x2=41.12 //y2=0.755
r932 (  174 175 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=41.005 //y=0.755 //x2=40.79 //y2=0.755
r933 (  173 263 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.635 //y=1.22 //x2=40.675 //y2=1.375
r934 (  172 262 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=40.635 //y=0.91 //x2=40.675 //y2=0.755
r935 (  172 173 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=40.635 //y=0.91 //x2=40.635 //y2=1.22
r936 (  168 256 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=28.255 //y=4.79 //x2=28.12 //y2=4.79
r937 (  167 169 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=28.455 //y=4.79 //x2=28.53 //y2=4.865
r938 (  167 168 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=28.455 //y=4.79 //x2=28.255 //y2=4.79
r939 (  166 261 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=28.21 //y=1.915 //x2=28.135 //y2=2.08
r940 (  165 259 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=28.21 //y=1.45 //x2=28.17 //y2=1.375
r941 (  165 166 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=28.21 //y=1.45 //x2=28.21 //y2=1.915
r942 (  164 259 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.21 //y=1.22 //x2=28.17 //y2=1.375
r943 (  163 258 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.21 //y=0.91 //x2=28.17 //y2=0.755
r944 (  163 164 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=28.21 //y=0.91 //x2=28.21 //y2=1.22
r945 (  158 252 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.84 //y=1.375 //x2=27.725 //y2=1.375
r946 (  157 259 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.055 //y=1.375 //x2=28.17 //y2=1.375
r947 (  156 251 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=27.84 //y=0.755 //x2=27.725 //y2=0.755
r948 (  155 258 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.055 //y=0.755 //x2=28.17 //y2=0.755
r949 (  155 156 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=28.055 //y=0.755 //x2=27.84 //y2=0.755
r950 (  154 252 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.685 //y=1.22 //x2=27.725 //y2=1.375
r951 (  153 251 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=27.685 //y=0.91 //x2=27.725 //y2=0.755
r952 (  153 154 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=27.685 //y=0.91 //x2=27.685 //y2=1.22
r953 (  149 245 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=15.305 //y=4.79 //x2=15.17 //y2=4.79
r954 (  148 150 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.505 //y=4.79 //x2=15.58 //y2=4.865
r955 (  148 149 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=15.505 //y=4.79 //x2=15.305 //y2=4.79
r956 (  147 250 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=15.26 //y=1.915 //x2=15.185 //y2=2.08
r957 (  146 248 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=15.26 //y=1.45 //x2=15.22 //y2=1.375
r958 (  146 147 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=15.26 //y=1.45 //x2=15.26 //y2=1.915
r959 (  145 248 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.26 //y=1.22 //x2=15.22 //y2=1.375
r960 (  144 247 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.26 //y=0.91 //x2=15.22 //y2=0.755
r961 (  144 145 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=15.26 //y=0.91 //x2=15.26 //y2=1.22
r962 (  139 241 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.89 //y=1.375 //x2=14.775 //y2=1.375
r963 (  138 248 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.105 //y=1.375 //x2=15.22 //y2=1.375
r964 (  137 240 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.89 //y=0.755 //x2=14.775 //y2=0.755
r965 (  136 247 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.105 //y=0.755 //x2=15.22 //y2=0.755
r966 (  136 137 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=15.105 //y=0.755 //x2=14.89 //y2=0.755
r967 (  135 241 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.735 //y=1.22 //x2=14.775 //y2=1.375
r968 (  134 240 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.735 //y=0.91 //x2=14.775 //y2=0.755
r969 (  134 135 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=14.735 //y=0.91 //x2=14.735 //y2=1.22
r970 (  130 234 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.355 //y=4.79 //x2=2.22 //y2=4.79
r971 (  129 131 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.63 //y2=4.865
r972 (  129 130 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.355 //y2=4.79
r973 (  128 239 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.915 //x2=2.235 //y2=2.08
r974 (  127 237 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.27 //y2=1.375
r975 (  127 128 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.31 //y2=1.915
r976 (  126 237 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.22 //x2=2.27 //y2=1.375
r977 (  125 236 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.27 //y2=0.755
r978 (  125 126 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.31 //y2=1.22
r979 (  120 230 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=1.375 //x2=1.825 //y2=1.375
r980 (  119 237 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=1.375 //x2=2.27 //y2=1.375
r981 (  118 229 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=0.755 //x2=1.825 //y2=0.755
r982 (  117 236 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=2.27 //y2=0.755
r983 (  117 118 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=1.94 //y2=0.755
r984 (  116 230 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=1.22 //x2=1.825 //y2=1.375
r985 (  115 229 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.825 //y2=0.755
r986 (  115 116 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.785 //y2=1.22
r987 (  114 226 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=67.38 //y=6.02 //x2=67.38 //y2=4.865
r988 (  113 290 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=66.94 //y=6.02 //x2=66.94 //y2=4.865
r989 (  112 207 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=54.43 //y=6.02 //x2=54.43 //y2=4.865
r990 (  111 279 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=53.99 //y=6.02 //x2=53.99 //y2=4.865
r991 (  110 188 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.48 //y=6.02 //x2=41.48 //y2=4.865
r992 (  109 268 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.04 //y=6.02 //x2=41.04 //y2=4.865
r993 (  108 169 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=28.53 //y=6.02 //x2=28.53 //y2=4.865
r994 (  107 257 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=28.09 //y=6.02 //x2=28.09 //y2=4.865
r995 (  106 150 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.58 //y=6.02 //x2=15.58 //y2=4.865
r996 (  105 246 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.14 //y=6.02 //x2=15.14 //y2=4.865
r997 (  104 131 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.63 //y=6.02 //x2=2.63 //y2=4.865
r998 (  103 235 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.19 //y=6.02 //x2=2.19 //y2=4.865
r999 (  102 214 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=66.797 //y=1.375 //x2=66.905 //y2=1.375
r1000 (  102 215 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=66.797 //y=1.375 //x2=66.69 //y2=1.375
r1001 (  101 195 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=53.847 //y=1.375 //x2=53.955 //y2=1.375
r1002 (  101 196 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=53.847 //y=1.375 //x2=53.74 //y2=1.375
r1003 (  100 176 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=40.897 //y=1.375 //x2=41.005 //y2=1.375
r1004 (  100 177 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=40.897 //y=1.375 //x2=40.79 //y2=1.375
r1005 (  99 157 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=27.947 //y=1.375 //x2=28.055 //y2=1.375
r1006 (  99 158 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=27.947 //y=1.375 //x2=27.84 //y2=1.375
r1007 (  98 138 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=14.997 //y=1.375 //x2=15.105 //y2=1.375
r1008 (  98 139 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=14.997 //y=1.375 //x2=14.89 //y2=1.375
r1009 (  97 119 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=2.155 //y2=1.375
r1010 (  97 120 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=1.94 //y2=1.375
r1011 (  95 287 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=66.97 //y=4.7 //x2=66.97 //y2=4.7
r1012 (  90 294 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=66.97 //y=2.08 //x2=66.97 //y2=2.08
r1013 (  87 276 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=54.02 //y=4.7 //x2=54.02 //y2=4.7
r1014 (  81 283 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=54.02 //y=2.08 //x2=54.02 //y2=2.08
r1015 (  78 265 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=41.07 //y=4.7 //x2=41.07 //y2=4.7
r1016 (  72 272 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=41.07 //y=2.08 //x2=41.07 //y2=2.08
r1017 (  69 254 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=28.12 //y=4.7 //x2=28.12 //y2=4.7
r1018 (  62 261 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=28.12 //y=2.08 //x2=28.12 //y2=2.08
r1019 (  59 243 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.17 //y=4.7 //x2=15.17 //y2=4.7
r1020 (  52 250 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.17 //y=2.08 //x2=15.17 //y2=2.08
r1021 (  49 232 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=4.7 //x2=2.22 //y2=4.7
r1022 (  40 239 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=2.08
r1023 (  38 95 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=66.97 //y=4.44 //x2=66.97 //y2=4.7
r1024 (  38 90 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=66.97 //y=4.44 //x2=66.97 //y2=2.08
r1025 (  37 87 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=54.02 //y=4.44 //x2=54.02 //y2=4.7
r1026 (  36 37 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=54.02 //y=3.7 //x2=54.02 //y2=4.44
r1027 (  36 81 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=54.02 //y=3.7 //x2=54.02 //y2=2.08
r1028 (  35 78 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=41.07 //y=4.44 //x2=41.07 //y2=4.7
r1029 (  34 35 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=41.07 //y=3.33 //x2=41.07 //y2=4.44
r1030 (  34 72 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=41.07 //y=3.33 //x2=41.07 //y2=2.08
r1031 (  33 69 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=28.12 //y=4.44 //x2=28.12 //y2=4.7
r1032 (  32 33 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=28.12 //y=3.7 //x2=28.12 //y2=4.44
r1033 (  31 32 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=28.12 //y=3.33 //x2=28.12 //y2=3.7
r1034 (  31 62 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=28.12 //y=3.33 //x2=28.12 //y2=2.08
r1035 (  30 59 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=15.17 //y=4.44 //x2=15.17 //y2=4.7
r1036 (  29 30 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=15.17 //y=3.33 //x2=15.17 //y2=4.44
r1037 (  28 29 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=15.17 //y=2.96 //x2=15.17 //y2=3.33
r1038 (  28 52 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=15.17 //y=2.96 //x2=15.17 //y2=2.08
r1039 (  27 49 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=2.22 //y=4.44 //x2=2.22 //y2=4.7
r1040 (  26 27 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.7 //x2=2.22 //y2=4.44
r1041 (  25 26 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.33 //x2=2.22 //y2=3.7
r1042 (  24 25 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.96 //x2=2.22 //y2=3.33
r1043 (  23 24 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.59 //x2=2.22 //y2=2.96
r1044 (  23 40 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.59 //x2=2.22 //y2=2.08
r1045 (  22 38 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=66.97 //y=4.44 //x2=66.97 //y2=4.44
r1046 (  20 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=54.02 //y=4.44 //x2=54.02 //y2=4.44
r1047 (  18 35 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=41.07 //y=4.44 //x2=41.07 //y2=4.44
r1048 (  16 33 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=28.12 //y=4.44 //x2=28.12 //y2=4.44
r1049 (  14 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.17 //y=4.44 //x2=15.17 //y2=4.44
r1050 (  12 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.22 //y=4.44 //x2=2.22 //y2=4.44
r1051 (  10 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=54.135 //y=4.44 //x2=54.02 //y2=4.44
r1052 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=66.855 //y=4.44 //x2=66.97 //y2=4.44
r1053 (  9 10 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=66.855 //y=4.44 //x2=54.135 //y2=4.44
r1054 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=41.185 //y=4.44 //x2=41.07 //y2=4.44
r1055 (  7 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=53.905 //y=4.44 //x2=54.02 //y2=4.44
r1056 (  7 8 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=53.905 //y=4.44 //x2=41.185 //y2=4.44
r1057 (  6 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=28.235 //y=4.44 //x2=28.12 //y2=4.44
r1058 (  5 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=40.955 //y=4.44 //x2=41.07 //y2=4.44
r1059 (  5 6 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=40.955 //y=4.44 //x2=28.235 //y2=4.44
r1060 (  4 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.285 //y=4.44 //x2=15.17 //y2=4.44
r1061 (  3 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=28.005 //y=4.44 //x2=28.12 //y2=4.44
r1062 (  3 4 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=28.005 //y=4.44 //x2=15.285 //y2=4.44
r1063 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.335 //y=4.44 //x2=2.22 //y2=4.44
r1064 (  1 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.055 //y=4.44 //x2=15.17 //y2=4.44
r1065 (  1 2 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=15.055 //y=4.44 //x2=2.335 //y2=4.44
ends PM_TMRDFFRNQNX1\%CLK

subckt PM_TMRDFFRNQNX1\%noxref_14 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 \
 63 64 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 92 94 100 101 102 \
 103 123 125 126 127 )
c259 ( 127 0 ) capacitor c=0.023087f //x=54.945 //y=5.02
c260 ( 126 0 ) capacitor c=0.023519f //x=54.065 //y=5.02
c261 ( 125 0 ) capacitor c=0.0224735f //x=53.185 //y=5.02
c262 ( 123 0 ) capacitor c=0.00853354f //x=55.195 //y=0.915
c263 ( 103 0 ) capacitor c=0.0558396f //x=70.945 //y=4.79
c264 ( 102 0 ) capacitor c=0.0298189f //x=71.235 //y=4.79
c265 ( 101 0 ) capacitor c=0.0347816f //x=70.9 //y=1.22
c266 ( 100 0 ) capacitor c=0.0187487f //x=70.9 //y=0.875
c267 ( 94 0 ) capacitor c=0.0137055f //x=70.745 //y=1.375
c268 ( 92 0 ) capacitor c=0.0149861f //x=70.745 //y=0.72
c269 ( 91 0 ) capacitor c=0.096037f //x=70.37 //y=1.915
c270 ( 90 0 ) capacitor c=0.0228993f //x=70.37 //y=1.53
c271 ( 89 0 ) capacitor c=0.0234352f //x=70.37 //y=1.22
c272 ( 88 0 ) capacitor c=0.0198724f //x=70.37 //y=0.875
c273 ( 84 0 ) capacitor c=0.0556143f //x=57.995 //y=4.79
c274 ( 83 0 ) capacitor c=0.0293157f //x=58.285 //y=4.79
c275 ( 82 0 ) capacitor c=0.0347816f //x=57.95 //y=1.22
c276 ( 81 0 ) capacitor c=0.0187487f //x=57.95 //y=0.875
c277 ( 75 0 ) capacitor c=0.0137055f //x=57.795 //y=1.375
c278 ( 73 0 ) capacitor c=0.0149861f //x=57.795 //y=0.72
c279 ( 72 0 ) capacitor c=0.096037f //x=57.42 //y=1.915
c280 ( 71 0 ) capacitor c=0.0228993f //x=57.42 //y=1.53
c281 ( 70 0 ) capacitor c=0.0234352f //x=57.42 //y=1.22
c282 ( 69 0 ) capacitor c=0.0198724f //x=57.42 //y=0.875
c283 ( 68 0 ) capacitor c=0.110114f //x=71.31 //y=6.02
c284 ( 67 0 ) capacitor c=0.158956f //x=70.87 //y=6.02
c285 ( 66 0 ) capacitor c=0.110114f //x=58.36 //y=6.02
c286 ( 65 0 ) capacitor c=0.158956f //x=57.92 //y=6.02
c287 ( 62 0 ) capacitor c=0.00106608f //x=55.09 //y=5.155
c288 ( 61 0 ) capacitor c=0.00207162f //x=54.21 //y=5.155
c289 ( 54 0 ) capacitor c=0.0992856f //x=70.67 //y=2.08
c290 ( 46 0 ) capacitor c=0.0936123f //x=57.72 //y=2.08
c291 ( 44 0 ) capacitor c=0.103742f //x=55.87 //y=3.7
c292 ( 40 0 ) capacitor c=0.00398962f //x=55.47 //y=1.665
c293 ( 39 0 ) capacitor c=0.0137288f //x=55.785 //y=1.665
c294 ( 33 0 ) capacitor c=0.0283082f //x=55.785 //y=5.155
c295 ( 25 0 ) capacitor c=0.0176454f //x=55.005 //y=5.155
c296 ( 18 0 ) capacitor c=0.00332903f //x=53.415 //y=5.155
c297 ( 17 0 ) capacitor c=0.014837f //x=54.125 //y=5.155
c298 ( 4 0 ) capacitor c=0.00424246f //x=57.835 //y=3.7
c299 ( 3 0 ) capacitor c=0.191185f //x=70.555 //y=3.7
c300 ( 2 0 ) capacitor c=0.0125346f //x=55.985 //y=3.7
c301 ( 1 0 ) capacitor c=0.0288301f //x=57.605 //y=3.7
r302 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=71.235 //y=4.79 //x2=71.31 //y2=4.865
r303 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=71.235 //y=4.79 //x2=70.945 //y2=4.79
r304 (  101 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.9 //y=1.22 //x2=70.86 //y2=1.375
r305 (  100 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.9 //y=0.875 //x2=70.86 //y2=0.72
r306 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=70.9 //y=0.875 //x2=70.9 //y2=1.22
r307 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=70.87 //y=4.865 //x2=70.945 //y2=4.79
r308 (  97 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=70.87 //y=4.865 //x2=70.67 //y2=4.7
r309 (  95 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.525 //y=1.375 //x2=70.41 //y2=1.375
r310 (  94 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.745 //y=1.375 //x2=70.86 //y2=1.375
r311 (  93 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.525 //y=0.72 //x2=70.41 //y2=0.72
r312 (  92 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.745 //y=0.72 //x2=70.86 //y2=0.72
r313 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=70.745 //y=0.72 //x2=70.525 //y2=0.72
r314 (  91 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=70.37 //y=1.915 //x2=70.67 //y2=2.08
r315 (  90 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.37 //y=1.53 //x2=70.41 //y2=1.375
r316 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=70.37 //y=1.53 //x2=70.37 //y2=1.915
r317 (  89 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.37 //y=1.22 //x2=70.41 //y2=1.375
r318 (  88 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.37 //y=0.875 //x2=70.41 //y2=0.72
r319 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=70.37 //y=0.875 //x2=70.37 //y2=1.22
r320 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=58.285 //y=4.79 //x2=58.36 //y2=4.865
r321 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=58.285 //y=4.79 //x2=57.995 //y2=4.79
r322 (  82 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=57.95 //y=1.22 //x2=57.91 //y2=1.375
r323 (  81 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=57.95 //y=0.875 //x2=57.91 //y2=0.72
r324 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=57.95 //y=0.875 //x2=57.95 //y2=1.22
r325 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=57.92 //y=4.865 //x2=57.995 //y2=4.79
r326 (  78 112 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=57.92 //y=4.865 //x2=57.72 //y2=4.7
r327 (  76 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=57.575 //y=1.375 //x2=57.46 //y2=1.375
r328 (  75 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=57.795 //y=1.375 //x2=57.91 //y2=1.375
r329 (  74 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=57.575 //y=0.72 //x2=57.46 //y2=0.72
r330 (  73 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=57.795 //y=0.72 //x2=57.91 //y2=0.72
r331 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=57.795 //y=0.72 //x2=57.575 //y2=0.72
r332 (  72 110 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=57.42 //y=1.915 //x2=57.72 //y2=2.08
r333 (  71 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=57.42 //y=1.53 //x2=57.46 //y2=1.375
r334 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=57.42 //y=1.53 //x2=57.42 //y2=1.915
r335 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=57.42 //y=1.22 //x2=57.46 //y2=1.375
r336 (  69 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=57.42 //y=0.875 //x2=57.46 //y2=0.72
r337 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=57.42 //y=0.875 //x2=57.42 //y2=1.22
r338 (  68 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=71.31 //y=6.02 //x2=71.31 //y2=4.865
r339 (  67 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=70.87 //y=6.02 //x2=70.87 //y2=4.865
r340 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=58.36 //y=6.02 //x2=58.36 //y2=4.865
r341 (  65 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=57.92 //y=6.02 //x2=57.92 //y2=4.865
r342 (  64 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=70.635 //y=1.375 //x2=70.745 //y2=1.375
r343 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=70.635 //y=1.375 //x2=70.525 //y2=1.375
r344 (  63 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=57.685 //y=1.375 //x2=57.795 //y2=1.375
r345 (  63 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=57.685 //y=1.375 //x2=57.575 //y2=1.375
r346 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=70.67 //y=4.7 //x2=70.67 //y2=4.7
r347 (  57 59 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=70.67 //y=3.7 //x2=70.67 //y2=4.7
r348 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=70.67 //y=2.08 //x2=70.67 //y2=2.08
r349 (  54 57 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=70.67 //y=2.08 //x2=70.67 //y2=3.7
r350 (  51 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=57.72 //y=4.7 //x2=57.72 //y2=4.7
r351 (  49 51 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=57.72 //y=3.7 //x2=57.72 //y2=4.7
r352 (  46 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=57.72 //y=2.08 //x2=57.72 //y2=2.08
r353 (  46 49 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=57.72 //y=2.08 //x2=57.72 //y2=3.7
r354 (  42 44 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=55.87 //y=5.07 //x2=55.87 //y2=3.7
r355 (  41 44 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=55.87 //y=1.75 //x2=55.87 //y2=3.7
r356 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=55.785 //y=1.665 //x2=55.87 //y2=1.75
r357 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=55.785 //y=1.665 //x2=55.47 //y2=1.665
r358 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=55.385 //y=1.58 //x2=55.47 //y2=1.665
r359 (  35 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=55.385 //y=1.58 //x2=55.385 //y2=1.01
r360 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.175 //y=5.155 //x2=55.09 //y2=5.155
r361 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=55.785 //y=5.155 //x2=55.87 //y2=5.07
r362 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=55.785 //y=5.155 //x2=55.175 //y2=5.155
r363 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.09 //y=5.24 //x2=55.09 //y2=5.155
r364 (  27 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=55.09 //y=5.24 //x2=55.09 //y2=5.725
r365 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.295 //y=5.155 //x2=54.21 //y2=5.155
r366 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.005 //y=5.155 //x2=55.09 //y2=5.155
r367 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=55.005 //y=5.155 //x2=54.295 //y2=5.155
r368 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.21 //y=5.24 //x2=54.21 //y2=5.155
r369 (  19 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=54.21 //y=5.24 //x2=54.21 //y2=5.725
r370 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.125 //y=5.155 //x2=54.21 //y2=5.155
r371 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=54.125 //y=5.155 //x2=53.415 //y2=5.155
r372 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=53.33 //y=5.24 //x2=53.415 //y2=5.155
r373 (  11 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=53.33 //y=5.24 //x2=53.33 //y2=5.725
r374 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=70.67 //y=3.7 //x2=70.67 //y2=3.7
r375 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=57.72 //y=3.7 //x2=57.72 //y2=3.7
r376 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=55.87 //y=3.7 //x2=55.87 //y2=3.7
r377 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=57.835 //y=3.7 //x2=57.72 //y2=3.7
r378 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=70.555 //y=3.7 //x2=70.67 //y2=3.7
r379 (  3 4 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=70.555 //y=3.7 //x2=57.835 //y2=3.7
r380 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=55.985 //y=3.7 //x2=55.87 //y2=3.7
r381 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=57.605 //y=3.7 //x2=57.72 //y2=3.7
r382 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=57.605 //y=3.7 //x2=55.985 //y2=3.7
ends PM_TMRDFFRNQNX1\%noxref_14

subckt PM_TMRDFFRNQNX1\%RN ( 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 35 36 37 \
 38 39 40 41 42 43 44 46 55 65 75 83 92 102 110 118 126 127 128 129 130 131 \
 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149 150 \
 151 152 156 157 158 163 165 168 169 173 174 175 180 182 185 186 187 188 189 \
 191 197 198 199 200 201 209 210 211 216 218 221 222 226 227 228 233 235 238 \
 239 240 241 242 244 250 251 252 253 254 262 263 264 269 271 274 275 279 280 \
 281 286 288 291 292 293 294 295 297 303 304 305 306 307 313 314 319 323 324 \
 329 335 344 345 350 354 355 360 366 375 376 381 385 386 391 397 )
c955 ( 397 0 ) capacitor c=0.0336203f //x=71.78 //y=4.7
c956 ( 391 0 ) capacitor c=0.0593675f //x=68.08 //y=4.7
c957 ( 386 0 ) capacitor c=0.0273931f //x=68.08 //y=1.915
c958 ( 385 0 ) capacitor c=0.0455604f //x=68.08 //y=2.08
c959 ( 381 0 ) capacitor c=0.0587755f //x=59.94 //y=4.7
c960 ( 376 0 ) capacitor c=0.0273931f //x=59.94 //y=1.915
c961 ( 375 0 ) capacitor c=0.0455604f //x=59.94 //y=2.08
c962 ( 366 0 ) capacitor c=0.0335551f //x=45.88 //y=4.7
c963 ( 360 0 ) capacitor c=0.058931f //x=42.18 //y=4.7
c964 ( 355 0 ) capacitor c=0.0273931f //x=42.18 //y=1.915
c965 ( 354 0 ) capacitor c=0.0455604f //x=42.18 //y=2.08
c966 ( 350 0 ) capacitor c=0.0587755f //x=34.04 //y=4.7
c967 ( 345 0 ) capacitor c=0.0273931f //x=34.04 //y=1.915
c968 ( 344 0 ) capacitor c=0.0455604f //x=34.04 //y=2.08
c969 ( 335 0 ) capacitor c=0.0335551f //x=19.98 //y=4.7
c970 ( 329 0 ) capacitor c=0.058931f //x=16.28 //y=4.7
c971 ( 324 0 ) capacitor c=0.0273931f //x=16.28 //y=1.915
c972 ( 323 0 ) capacitor c=0.0455604f //x=16.28 //y=2.08
c973 ( 319 0 ) capacitor c=0.0587755f //x=8.14 //y=4.7
c974 ( 314 0 ) capacitor c=0.0273931f //x=8.14 //y=1.915
c975 ( 313 0 ) capacitor c=0.0457326f //x=8.14 //y=2.08
c976 ( 307 0 ) capacitor c=0.024933f //x=72.115 //y=4.79
c977 ( 306 0 ) capacitor c=0.0827272f //x=71.87 //y=1.915
c978 ( 305 0 ) capacitor c=0.0170266f //x=71.87 //y=1.45
c979 ( 304 0 ) capacitor c=0.018609f //x=71.87 //y=1.22
c980 ( 303 0 ) capacitor c=0.0187309f //x=71.87 //y=0.91
c981 ( 297 0 ) capacitor c=0.014725f //x=71.715 //y=1.375
c982 ( 295 0 ) capacitor c=0.0146567f //x=71.715 //y=0.755
c983 ( 294 0 ) capacitor c=0.0335408f //x=71.345 //y=1.22
c984 ( 293 0 ) capacitor c=0.0173761f //x=71.345 //y=0.91
c985 ( 292 0 ) capacitor c=0.0432517f //x=68.6 //y=1.26
c986 ( 291 0 ) capacitor c=0.0200379f //x=68.6 //y=0.915
c987 ( 288 0 ) capacitor c=0.0148873f //x=68.445 //y=1.415
c988 ( 286 0 ) capacitor c=0.0157803f //x=68.445 //y=0.76
c989 ( 281 0 ) capacitor c=0.0218028f //x=68.07 //y=1.57
c990 ( 280 0 ) capacitor c=0.0207459f //x=68.07 //y=1.26
c991 ( 279 0 ) capacitor c=0.0194308f //x=68.07 //y=0.915
c992 ( 275 0 ) capacitor c=0.0432517f //x=60.46 //y=1.26
c993 ( 274 0 ) capacitor c=0.0200379f //x=60.46 //y=0.915
c994 ( 271 0 ) capacitor c=0.0148873f //x=60.305 //y=1.415
c995 ( 269 0 ) capacitor c=0.0157803f //x=60.305 //y=0.76
c996 ( 264 0 ) capacitor c=0.0218028f //x=59.93 //y=1.57
c997 ( 263 0 ) capacitor c=0.0207459f //x=59.93 //y=1.26
c998 ( 262 0 ) capacitor c=0.0194308f //x=59.93 //y=0.915
c999 ( 254 0 ) capacitor c=0.0245352f //x=46.215 //y=4.79
c1000 ( 253 0 ) capacitor c=0.0825033f //x=45.97 //y=1.915
c1001 ( 252 0 ) capacitor c=0.0170266f //x=45.97 //y=1.45
c1002 ( 251 0 ) capacitor c=0.018609f //x=45.97 //y=1.22
c1003 ( 250 0 ) capacitor c=0.0187309f //x=45.97 //y=0.91
c1004 ( 244 0 ) capacitor c=0.014725f //x=45.815 //y=1.375
c1005 ( 242 0 ) capacitor c=0.0146567f //x=45.815 //y=0.755
c1006 ( 241 0 ) capacitor c=0.0335408f //x=45.445 //y=1.22
c1007 ( 240 0 ) capacitor c=0.0173761f //x=45.445 //y=0.91
c1008 ( 239 0 ) capacitor c=0.0432517f //x=42.7 //y=1.26
c1009 ( 238 0 ) capacitor c=0.0200379f //x=42.7 //y=0.915
c1010 ( 235 0 ) capacitor c=0.0148873f //x=42.545 //y=1.415
c1011 ( 233 0 ) capacitor c=0.0157803f //x=42.545 //y=0.76
c1012 ( 228 0 ) capacitor c=0.0218028f //x=42.17 //y=1.57
c1013 ( 227 0 ) capacitor c=0.0207459f //x=42.17 //y=1.26
c1014 ( 226 0 ) capacitor c=0.0194308f //x=42.17 //y=0.915
c1015 ( 222 0 ) capacitor c=0.0432517f //x=34.56 //y=1.26
c1016 ( 221 0 ) capacitor c=0.0200379f //x=34.56 //y=0.915
c1017 ( 218 0 ) capacitor c=0.0148873f //x=34.405 //y=1.415
c1018 ( 216 0 ) capacitor c=0.0157803f //x=34.405 //y=0.76
c1019 ( 211 0 ) capacitor c=0.0218028f //x=34.03 //y=1.57
c1020 ( 210 0 ) capacitor c=0.0207459f //x=34.03 //y=1.26
c1021 ( 209 0 ) capacitor c=0.0194308f //x=34.03 //y=0.915
c1022 ( 201 0 ) capacitor c=0.0245352f //x=20.315 //y=4.79
c1023 ( 200 0 ) capacitor c=0.0825033f //x=20.07 //y=1.915
c1024 ( 199 0 ) capacitor c=0.0170266f //x=20.07 //y=1.45
c1025 ( 198 0 ) capacitor c=0.018609f //x=20.07 //y=1.22
c1026 ( 197 0 ) capacitor c=0.0187309f //x=20.07 //y=0.91
c1027 ( 191 0 ) capacitor c=0.014725f //x=19.915 //y=1.375
c1028 ( 189 0 ) capacitor c=0.0146567f //x=19.915 //y=0.755
c1029 ( 188 0 ) capacitor c=0.0335408f //x=19.545 //y=1.22
c1030 ( 187 0 ) capacitor c=0.0173761f //x=19.545 //y=0.91
c1031 ( 186 0 ) capacitor c=0.0432517f //x=16.8 //y=1.26
c1032 ( 185 0 ) capacitor c=0.0200379f //x=16.8 //y=0.915
c1033 ( 182 0 ) capacitor c=0.0148873f //x=16.645 //y=1.415
c1034 ( 180 0 ) capacitor c=0.0157803f //x=16.645 //y=0.76
c1035 ( 175 0 ) capacitor c=0.0218028f //x=16.27 //y=1.57
c1036 ( 174 0 ) capacitor c=0.0207459f //x=16.27 //y=1.26
c1037 ( 173 0 ) capacitor c=0.0194308f //x=16.27 //y=0.915
c1038 ( 169 0 ) capacitor c=0.0432517f //x=8.66 //y=1.26
c1039 ( 168 0 ) capacitor c=0.0200379f //x=8.66 //y=0.915
c1040 ( 165 0 ) capacitor c=0.0148873f //x=8.505 //y=1.415
c1041 ( 163 0 ) capacitor c=0.0157803f //x=8.505 //y=0.76
c1042 ( 158 0 ) capacitor c=0.0218028f //x=8.13 //y=1.57
c1043 ( 157 0 ) capacitor c=0.0207459f //x=8.13 //y=1.26
c1044 ( 156 0 ) capacitor c=0.0194308f //x=8.13 //y=0.915
c1045 ( 152 0 ) capacitor c=0.110114f //x=72.19 //y=6.02
c1046 ( 151 0 ) capacitor c=0.11012f //x=71.75 //y=6.02
c1047 ( 150 0 ) capacitor c=0.158794f //x=68.26 //y=6.02
c1048 ( 149 0 ) capacitor c=0.110114f //x=67.82 //y=6.02
c1049 ( 148 0 ) capacitor c=0.158794f //x=60.12 //y=6.02
c1050 ( 147 0 ) capacitor c=0.110114f //x=59.68 //y=6.02
c1051 ( 146 0 ) capacitor c=0.110114f //x=46.29 //y=6.02
c1052 ( 145 0 ) capacitor c=0.11012f //x=45.85 //y=6.02
c1053 ( 144 0 ) capacitor c=0.158794f //x=42.36 //y=6.02
c1054 ( 143 0 ) capacitor c=0.110114f //x=41.92 //y=6.02
c1055 ( 142 0 ) capacitor c=0.158794f //x=34.22 //y=6.02
c1056 ( 141 0 ) capacitor c=0.110114f //x=33.78 //y=6.02
c1057 ( 140 0 ) capacitor c=0.110114f //x=20.39 //y=6.02
c1058 ( 139 0 ) capacitor c=0.11012f //x=19.95 //y=6.02
c1059 ( 138 0 ) capacitor c=0.158794f //x=16.46 //y=6.02
c1060 ( 137 0 ) capacitor c=0.110114f //x=16.02 //y=6.02
c1061 ( 136 0 ) capacitor c=0.158794f //x=8.32 //y=6.02
c1062 ( 135 0 ) capacitor c=0.110114f //x=7.88 //y=6.02
c1063 ( 118 0 ) capacitor c=0.0945052f //x=71.78 //y=2.08
c1064 ( 110 0 ) capacitor c=0.0837702f //x=68.08 //y=2.08
c1065 ( 102 0 ) capacitor c=0.0813451f //x=59.94 //y=2.08
c1066 ( 92 0 ) capacitor c=0.0915318f //x=45.88 //y=2.08
c1067 ( 83 0 ) capacitor c=0.081834f //x=42.18 //y=2.08
c1068 ( 75 0 ) capacitor c=0.0797116f //x=34.04 //y=2.08
c1069 ( 65 0 ) capacitor c=0.0945052f //x=19.98 //y=2.08
c1070 ( 55 0 ) capacitor c=0.0841472f //x=16.28 //y=2.08
c1071 ( 46 0 ) capacitor c=0.0820248f //x=8.14 //y=2.08
c1072 ( 16 0 ) capacitor c=0.00626813f //x=68.195 //y=2.22
c1073 ( 15 0 ) capacitor c=0.0949894f //x=71.665 //y=2.22
c1074 ( 14 0 ) capacitor c=0.00730636f //x=60.055 //y=2.22
c1075 ( 13 0 ) capacitor c=0.180678f //x=67.965 //y=2.22
c1076 ( 12 0 ) capacitor c=0.00575878f //x=45.995 //y=2.22
c1077 ( 11 0 ) capacitor c=0.271811f //x=59.825 //y=2.22
c1078 ( 10 0 ) capacitor c=0.00601486f //x=42.295 //y=2.22
c1079 ( 9 0 ) capacitor c=0.0680922f //x=45.765 //y=2.22
c1080 ( 8 0 ) capacitor c=0.00705309f //x=34.155 //y=2.22
c1081 ( 7 0 ) capacitor c=0.153868f //x=42.065 //y=2.22
c1082 ( 6 0 ) capacitor c=0.00575878f //x=20.095 //y=2.22
c1083 ( 5 0 ) capacitor c=0.269152f //x=33.925 //y=2.22
c1084 ( 4 0 ) capacitor c=0.00601486f //x=16.395 //y=2.22
c1085 ( 3 0 ) capacitor c=0.0680922f //x=19.865 //y=2.22
c1086 ( 2 0 ) capacitor c=0.0153965f //x=8.255 //y=2.22
c1087 ( 1 0 ) capacitor c=0.153868f //x=16.165 //y=2.22
r1088 (  399 400 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=71.78 //y=4.79 //x2=71.78 //y2=4.865
r1089 (  397 399 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=71.78 //y=4.7 //x2=71.78 //y2=4.79
r1090 (  385 386 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=68.08 //y=2.08 //x2=68.08 //y2=1.915
r1091 (  375 376 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=59.94 //y=2.08 //x2=59.94 //y2=1.915
r1092 (  368 369 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=45.88 //y=4.79 //x2=45.88 //y2=4.865
r1093 (  366 368 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=45.88 //y=4.7 //x2=45.88 //y2=4.79
r1094 (  354 355 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=42.18 //y=2.08 //x2=42.18 //y2=1.915
r1095 (  344 345 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=34.04 //y=2.08 //x2=34.04 //y2=1.915
r1096 (  337 338 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=19.98 //y=4.79 //x2=19.98 //y2=4.865
r1097 (  335 337 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=19.98 //y=4.7 //x2=19.98 //y2=4.79
r1098 (  323 324 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=16.28 //y=2.08 //x2=16.28 //y2=1.915
r1099 (  313 314 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=8.14 //y=2.08 //x2=8.14 //y2=1.915
r1100 (  308 399 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=71.915 //y=4.79 //x2=71.78 //y2=4.79
r1101 (  307 309 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=72.115 //y=4.79 //x2=72.19 //y2=4.865
r1102 (  307 308 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=72.115 //y=4.79 //x2=71.915 //y2=4.79
r1103 (  306 404 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=71.87 //y=1.915 //x2=71.795 //y2=2.08
r1104 (  305 402 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=71.87 //y=1.45 //x2=71.83 //y2=1.375
r1105 (  305 306 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=71.87 //y=1.45 //x2=71.87 //y2=1.915
r1106 (  304 402 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.87 //y=1.22 //x2=71.83 //y2=1.375
r1107 (  303 401 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.87 //y=0.91 //x2=71.83 //y2=0.755
r1108 (  303 304 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=71.87 //y=0.91 //x2=71.87 //y2=1.22
r1109 (  298 395 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=71.5 //y=1.375 //x2=71.385 //y2=1.375
r1110 (  297 402 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=71.715 //y=1.375 //x2=71.83 //y2=1.375
r1111 (  296 394 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=71.5 //y=0.755 //x2=71.385 //y2=0.755
r1112 (  295 401 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=71.715 //y=0.755 //x2=71.83 //y2=0.755
r1113 (  295 296 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=71.715 //y=0.755 //x2=71.5 //y2=0.755
r1114 (  294 395 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.345 //y=1.22 //x2=71.385 //y2=1.375
r1115 (  293 394 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.345 //y=0.91 //x2=71.385 //y2=0.755
r1116 (  293 294 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=71.345 //y=0.91 //x2=71.345 //y2=1.22
r1117 (  292 393 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.6 //y=1.26 //x2=68.56 //y2=1.415
r1118 (  291 392 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.6 //y=0.915 //x2=68.56 //y2=0.76
r1119 (  291 292 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=68.6 //y=0.915 //x2=68.6 //y2=1.26
r1120 (  289 389 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.225 //y=1.415 //x2=68.11 //y2=1.415
r1121 (  288 393 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.445 //y=1.415 //x2=68.56 //y2=1.415
r1122 (  287 388 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.225 //y=0.76 //x2=68.11 //y2=0.76
r1123 (  286 392 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=68.445 //y=0.76 //x2=68.56 //y2=0.76
r1124 (  286 287 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=68.445 //y=0.76 //x2=68.225 //y2=0.76
r1125 (  283 391 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=68.26 //y=4.865 //x2=68.08 //y2=4.7
r1126 (  281 389 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.07 //y=1.57 //x2=68.11 //y2=1.415
r1127 (  281 386 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=68.07 //y=1.57 //x2=68.07 //y2=1.915
r1128 (  280 389 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.07 //y=1.26 //x2=68.11 //y2=1.415
r1129 (  279 388 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=68.07 //y=0.915 //x2=68.11 //y2=0.76
r1130 (  279 280 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=68.07 //y=0.915 //x2=68.07 //y2=1.26
r1131 (  276 391 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=67.82 //y=4.865 //x2=68.08 //y2=4.7
r1132 (  275 383 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.46 //y=1.26 //x2=60.42 //y2=1.415
r1133 (  274 382 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.46 //y=0.915 //x2=60.42 //y2=0.76
r1134 (  274 275 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=60.46 //y=0.915 //x2=60.46 //y2=1.26
r1135 (  272 379 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=60.085 //y=1.415 //x2=59.97 //y2=1.415
r1136 (  271 383 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=60.305 //y=1.415 //x2=60.42 //y2=1.415
r1137 (  270 378 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=60.085 //y=0.76 //x2=59.97 //y2=0.76
r1138 (  269 382 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=60.305 //y=0.76 //x2=60.42 //y2=0.76
r1139 (  269 270 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=60.305 //y=0.76 //x2=60.085 //y2=0.76
r1140 (  266 381 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=60.12 //y=4.865 //x2=59.94 //y2=4.7
r1141 (  264 379 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.93 //y=1.57 //x2=59.97 //y2=1.415
r1142 (  264 376 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=59.93 //y=1.57 //x2=59.93 //y2=1.915
r1143 (  263 379 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.93 //y=1.26 //x2=59.97 //y2=1.415
r1144 (  262 378 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.93 //y=0.915 //x2=59.97 //y2=0.76
r1145 (  262 263 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=59.93 //y=0.915 //x2=59.93 //y2=1.26
r1146 (  259 381 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=59.68 //y=4.865 //x2=59.94 //y2=4.7
r1147 (  255 368 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=46.015 //y=4.79 //x2=45.88 //y2=4.79
r1148 (  254 256 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=46.215 //y=4.79 //x2=46.29 //y2=4.865
r1149 (  254 255 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=46.215 //y=4.79 //x2=46.015 //y2=4.79
r1150 (  253 373 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=45.97 //y=1.915 //x2=45.895 //y2=2.08
r1151 (  252 371 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=45.97 //y=1.45 //x2=45.93 //y2=1.375
r1152 (  252 253 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=45.97 //y=1.45 //x2=45.97 //y2=1.915
r1153 (  251 371 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.97 //y=1.22 //x2=45.93 //y2=1.375
r1154 (  250 370 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.97 //y=0.91 //x2=45.93 //y2=0.755
r1155 (  250 251 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=45.97 //y=0.91 //x2=45.97 //y2=1.22
r1156 (  245 364 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.6 //y=1.375 //x2=45.485 //y2=1.375
r1157 (  244 371 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.815 //y=1.375 //x2=45.93 //y2=1.375
r1158 (  243 363 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.6 //y=0.755 //x2=45.485 //y2=0.755
r1159 (  242 370 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.815 //y=0.755 //x2=45.93 //y2=0.755
r1160 (  242 243 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=45.815 //y=0.755 //x2=45.6 //y2=0.755
r1161 (  241 364 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.445 //y=1.22 //x2=45.485 //y2=1.375
r1162 (  240 363 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.445 //y=0.91 //x2=45.485 //y2=0.755
r1163 (  240 241 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=45.445 //y=0.91 //x2=45.445 //y2=1.22
r1164 (  239 362 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.7 //y=1.26 //x2=42.66 //y2=1.415
r1165 (  238 361 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.7 //y=0.915 //x2=42.66 //y2=0.76
r1166 (  238 239 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=42.7 //y=0.915 //x2=42.7 //y2=1.26
r1167 (  236 358 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.325 //y=1.415 //x2=42.21 //y2=1.415
r1168 (  235 362 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.545 //y=1.415 //x2=42.66 //y2=1.415
r1169 (  234 357 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.325 //y=0.76 //x2=42.21 //y2=0.76
r1170 (  233 361 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.545 //y=0.76 //x2=42.66 //y2=0.76
r1171 (  233 234 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=42.545 //y=0.76 //x2=42.325 //y2=0.76
r1172 (  230 360 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=42.36 //y=4.865 //x2=42.18 //y2=4.7
r1173 (  228 358 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.17 //y=1.57 //x2=42.21 //y2=1.415
r1174 (  228 355 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=42.17 //y=1.57 //x2=42.17 //y2=1.915
r1175 (  227 358 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.17 //y=1.26 //x2=42.21 //y2=1.415
r1176 (  226 357 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.17 //y=0.915 //x2=42.21 //y2=0.76
r1177 (  226 227 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=42.17 //y=0.915 //x2=42.17 //y2=1.26
r1178 (  223 360 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=41.92 //y=4.865 //x2=42.18 //y2=4.7
r1179 (  222 352 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.56 //y=1.26 //x2=34.52 //y2=1.415
r1180 (  221 351 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.56 //y=0.915 //x2=34.52 //y2=0.76
r1181 (  221 222 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=34.56 //y=0.915 //x2=34.56 //y2=1.26
r1182 (  219 348 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.185 //y=1.415 //x2=34.07 //y2=1.415
r1183 (  218 352 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.405 //y=1.415 //x2=34.52 //y2=1.415
r1184 (  217 347 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.185 //y=0.76 //x2=34.07 //y2=0.76
r1185 (  216 351 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.405 //y=0.76 //x2=34.52 //y2=0.76
r1186 (  216 217 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=34.405 //y=0.76 //x2=34.185 //y2=0.76
r1187 (  213 350 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=34.22 //y=4.865 //x2=34.04 //y2=4.7
r1188 (  211 348 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.03 //y=1.57 //x2=34.07 //y2=1.415
r1189 (  211 345 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=34.03 //y=1.57 //x2=34.03 //y2=1.915
r1190 (  210 348 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.03 //y=1.26 //x2=34.07 //y2=1.415
r1191 (  209 347 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.03 //y=0.915 //x2=34.07 //y2=0.76
r1192 (  209 210 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=34.03 //y=0.915 //x2=34.03 //y2=1.26
r1193 (  206 350 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=33.78 //y=4.865 //x2=34.04 //y2=4.7
r1194 (  202 337 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=20.115 //y=4.79 //x2=19.98 //y2=4.79
r1195 (  201 203 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.315 //y=4.79 //x2=20.39 //y2=4.865
r1196 (  201 202 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=20.315 //y=4.79 //x2=20.115 //y2=4.79
r1197 (  200 342 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=20.07 //y=1.915 //x2=19.995 //y2=2.08
r1198 (  199 340 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=20.07 //y=1.45 //x2=20.03 //y2=1.375
r1199 (  199 200 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=20.07 //y=1.45 //x2=20.07 //y2=1.915
r1200 (  198 340 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.07 //y=1.22 //x2=20.03 //y2=1.375
r1201 (  197 339 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.07 //y=0.91 //x2=20.03 //y2=0.755
r1202 (  197 198 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=20.07 //y=0.91 //x2=20.07 //y2=1.22
r1203 (  192 333 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.7 //y=1.375 //x2=19.585 //y2=1.375
r1204 (  191 340 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.915 //y=1.375 //x2=20.03 //y2=1.375
r1205 (  190 332 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.7 //y=0.755 //x2=19.585 //y2=0.755
r1206 (  189 339 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.915 //y=0.755 //x2=20.03 //y2=0.755
r1207 (  189 190 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=19.915 //y=0.755 //x2=19.7 //y2=0.755
r1208 (  188 333 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.545 //y=1.22 //x2=19.585 //y2=1.375
r1209 (  187 332 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.545 //y=0.91 //x2=19.585 //y2=0.755
r1210 (  187 188 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=19.545 //y=0.91 //x2=19.545 //y2=1.22
r1211 (  186 331 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.8 //y=1.26 //x2=16.76 //y2=1.415
r1212 (  185 330 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.8 //y=0.915 //x2=16.76 //y2=0.76
r1213 (  185 186 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.8 //y=0.915 //x2=16.8 //y2=1.26
r1214 (  183 327 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.425 //y=1.415 //x2=16.31 //y2=1.415
r1215 (  182 331 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.645 //y=1.415 //x2=16.76 //y2=1.415
r1216 (  181 326 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.425 //y=0.76 //x2=16.31 //y2=0.76
r1217 (  180 330 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.645 //y=0.76 //x2=16.76 //y2=0.76
r1218 (  180 181 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=16.645 //y=0.76 //x2=16.425 //y2=0.76
r1219 (  177 329 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=16.46 //y=4.865 //x2=16.28 //y2=4.7
r1220 (  175 327 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.27 //y=1.57 //x2=16.31 //y2=1.415
r1221 (  175 324 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.27 //y=1.57 //x2=16.27 //y2=1.915
r1222 (  174 327 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.27 //y=1.26 //x2=16.31 //y2=1.415
r1223 (  173 326 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.27 //y=0.915 //x2=16.31 //y2=0.76
r1224 (  173 174 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.27 //y=0.915 //x2=16.27 //y2=1.26
r1225 (  170 329 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=16.02 //y=4.865 //x2=16.28 //y2=4.7
r1226 (  169 321 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.66 //y=1.26 //x2=8.62 //y2=1.415
r1227 (  168 320 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.66 //y=0.915 //x2=8.62 //y2=0.76
r1228 (  168 169 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.66 //y=0.915 //x2=8.66 //y2=1.26
r1229 (  166 317 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.285 //y=1.415 //x2=8.17 //y2=1.415
r1230 (  165 321 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.505 //y=1.415 //x2=8.62 //y2=1.415
r1231 (  164 316 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.285 //y=0.76 //x2=8.17 //y2=0.76
r1232 (  163 320 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.505 //y=0.76 //x2=8.62 //y2=0.76
r1233 (  163 164 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=8.505 //y=0.76 //x2=8.285 //y2=0.76
r1234 (  160 319 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=8.32 //y=4.865 //x2=8.14 //y2=4.7
r1235 (  158 317 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.57 //x2=8.17 //y2=1.415
r1236 (  158 314 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.57 //x2=8.13 //y2=1.915
r1237 (  157 317 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.26 //x2=8.17 //y2=1.415
r1238 (  156 316 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=0.915 //x2=8.17 //y2=0.76
r1239 (  156 157 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.13 //y=0.915 //x2=8.13 //y2=1.26
r1240 (  153 319 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=7.88 //y=4.865 //x2=8.14 //y2=4.7
r1241 (  152 309 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=72.19 //y=6.02 //x2=72.19 //y2=4.865
r1242 (  151 400 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=71.75 //y=6.02 //x2=71.75 //y2=4.865
r1243 (  150 283 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=68.26 //y=6.02 //x2=68.26 //y2=4.865
r1244 (  149 276 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=67.82 //y=6.02 //x2=67.82 //y2=4.865
r1245 (  148 266 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=60.12 //y=6.02 //x2=60.12 //y2=4.865
r1246 (  147 259 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.68 //y=6.02 //x2=59.68 //y2=4.865
r1247 (  146 256 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=46.29 //y=6.02 //x2=46.29 //y2=4.865
r1248 (  145 369 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.85 //y=6.02 //x2=45.85 //y2=4.865
r1249 (  144 230 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=42.36 //y=6.02 //x2=42.36 //y2=4.865
r1250 (  143 223 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.92 //y=6.02 //x2=41.92 //y2=4.865
r1251 (  142 213 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=34.22 //y=6.02 //x2=34.22 //y2=4.865
r1252 (  141 206 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=33.78 //y=6.02 //x2=33.78 //y2=4.865
r1253 (  140 203 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.39 //y=6.02 //x2=20.39 //y2=4.865
r1254 (  139 338 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.95 //y=6.02 //x2=19.95 //y2=4.865
r1255 (  138 177 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.46 //y=6.02 //x2=16.46 //y2=4.865
r1256 (  137 170 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.02 //y=6.02 //x2=16.02 //y2=4.865
r1257 (  136 160 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.32 //y=6.02 //x2=8.32 //y2=4.865
r1258 (  135 153 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.88 //y=6.02 //x2=7.88 //y2=4.865
r1259 (  134 297 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=71.607 //y=1.375 //x2=71.715 //y2=1.375
r1260 (  134 298 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=71.607 //y=1.375 //x2=71.5 //y2=1.375
r1261 (  133 288 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=68.335 //y=1.415 //x2=68.445 //y2=1.415
r1262 (  133 289 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=68.335 //y=1.415 //x2=68.225 //y2=1.415
r1263 (  132 271 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=60.195 //y=1.415 //x2=60.305 //y2=1.415
r1264 (  132 272 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=60.195 //y=1.415 //x2=60.085 //y2=1.415
r1265 (  131 244 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=45.707 //y=1.375 //x2=45.815 //y2=1.375
r1266 (  131 245 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=45.707 //y=1.375 //x2=45.6 //y2=1.375
r1267 (  130 235 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=42.435 //y=1.415 //x2=42.545 //y2=1.415
r1268 (  130 236 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=42.435 //y=1.415 //x2=42.325 //y2=1.415
r1269 (  129 218 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=34.295 //y=1.415 //x2=34.405 //y2=1.415
r1270 (  129 219 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=34.295 //y=1.415 //x2=34.185 //y2=1.415
r1271 (  128 191 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=19.807 //y=1.375 //x2=19.915 //y2=1.375
r1272 (  128 192 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=19.807 //y=1.375 //x2=19.7 //y2=1.375
r1273 (  127 182 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=16.535 //y=1.415 //x2=16.645 //y2=1.415
r1274 (  127 183 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=16.535 //y=1.415 //x2=16.425 //y2=1.415
r1275 (  126 165 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.395 //y=1.415 //x2=8.505 //y2=1.415
r1276 (  126 166 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.395 //y=1.415 //x2=8.285 //y2=1.415
r1277 (  124 397 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=71.78 //y=4.7 //x2=71.78 //y2=4.7
r1278 (  118 404 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=71.78 //y=2.08 //x2=71.78 //y2=2.08
r1279 (  118 121 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=71.78 //y=2.08 //x2=71.78 //y2=2.22
r1280 (  115 391 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=68.08 //y=4.7 //x2=68.08 //y2=4.7
r1281 (  113 115 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=68.08 //y=2.22 //x2=68.08 //y2=4.7
r1282 (  110 385 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=68.08 //y=2.08 //x2=68.08 //y2=2.08
r1283 (  110 113 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=68.08 //y=2.08 //x2=68.08 //y2=2.22
r1284 (  107 381 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=59.94 //y=4.7 //x2=59.94 //y2=4.7
r1285 (  105 107 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=59.94 //y=2.22 //x2=59.94 //y2=4.7
r1286 (  102 375 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=59.94 //y=2.08 //x2=59.94 //y2=2.08
r1287 (  102 105 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=59.94 //y=2.08 //x2=59.94 //y2=2.22
r1288 (  99 366 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=45.88 //y=4.7 //x2=45.88 //y2=4.7
r1289 (  92 373 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=45.88 //y=2.08 //x2=45.88 //y2=2.08
r1290 (  92 95 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=45.88 //y=2.08 //x2=45.88 //y2=2.22
r1291 (  89 360 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=42.18 //y=4.7 //x2=42.18 //y2=4.7
r1292 (  83 354 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=42.18 //y=2.08 //x2=42.18 //y2=2.08
r1293 (  83 86 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=42.18 //y=2.08 //x2=42.18 //y2=2.22
r1294 (  80 350 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.04 //y=4.7 //x2=34.04 //y2=4.7
r1295 (  78 80 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=34.04 //y=2.22 //x2=34.04 //y2=4.7
r1296 (  75 344 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.04 //y=2.08 //x2=34.04 //y2=2.08
r1297 (  75 78 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=34.04 //y=2.08 //x2=34.04 //y2=2.22
r1298 (  72 335 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.98 //y=4.7 //x2=19.98 //y2=4.7
r1299 (  65 342 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.98 //y=2.08 //x2=19.98 //y2=2.08
r1300 (  65 68 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.08 //x2=19.98 //y2=2.22
r1301 (  62 329 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.28 //y=4.7 //x2=16.28 //y2=4.7
r1302 (  55 323 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.28 //y=2.08 //x2=16.28 //y2=2.08
r1303 (  55 58 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=16.28 //y=2.08 //x2=16.28 //y2=2.22
r1304 (  52 319 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.14 //y=4.7 //x2=8.14 //y2=4.7
r1305 (  46 313 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.14 //y=2.08 //x2=8.14 //y2=2.08
r1306 (  44 124 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li \
 //thickness=0.1 //x=71.78 //y=3.7 //x2=71.78 //y2=4.7
r1307 (  44 121 ) resistor r=101.305 //w=0.187 //l=1.48 //layer=li \
 //thickness=0.1 //x=71.78 //y=3.7 //x2=71.78 //y2=2.22
r1308 (  43 99 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=45.88 //y=3.7 //x2=45.88 //y2=4.7
r1309 (  42 43 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=45.88 //y=3.33 //x2=45.88 //y2=3.7
r1310 (  42 95 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=45.88 //y=3.33 //x2=45.88 //y2=2.22
r1311 (  41 89 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=42.18 //y=3.33 //x2=42.18 //y2=4.7
r1312 (  41 86 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=42.18 //y=3.33 //x2=42.18 //y2=2.22
r1313 (  40 72 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=19.98 //y=3.33 //x2=19.98 //y2=4.7
r1314 (  39 40 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.96 //x2=19.98 //y2=3.33
r1315 (  39 68 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.96 //x2=19.98 //y2=2.22
r1316 (  38 62 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=16.28 //y=3.33 //x2=16.28 //y2=4.7
r1317 (  37 38 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=16.28 //y=2.96 //x2=16.28 //y2=3.33
r1318 (  37 58 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=16.28 //y=2.96 //x2=16.28 //y2=2.22
r1319 (  36 52 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=8.14 //y=2.96 //x2=8.14 //y2=4.7
r1320 (  35 36 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=8.14 //y=2.22 //x2=8.14 //y2=2.96
r1321 (  35 46 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=8.14 //y=2.22 //x2=8.14 //y2=2.08
r1322 (  34 121 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=71.78 //y=2.22 //x2=71.78 //y2=2.22
r1323 (  32 113 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=68.08 //y=2.22 //x2=68.08 //y2=2.22
r1324 (  30 105 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=59.94 //y=2.22 //x2=59.94 //y2=2.22
r1325 (  28 95 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=45.88 //y=2.22 //x2=45.88 //y2=2.22
r1326 (  26 86 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=42.18 //y=2.22 //x2=42.18 //y2=2.22
r1327 (  24 78 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=34.04 //y=2.22 //x2=34.04 //y2=2.22
r1328 (  22 68 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=19.98 //y=2.22 //x2=19.98 //y2=2.22
r1329 (  20 58 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=16.28 //y=2.22 //x2=16.28 //y2=2.22
r1330 (  18 35 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.14 //y=2.22 //x2=8.14 //y2=2.22
r1331 (  16 32 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=68.195 //y=2.22 //x2=68.08 //y2=2.22
r1332 (  15 34 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=71.665 //y=2.22 //x2=71.78 //y2=2.22
r1333 (  15 16 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=71.665 //y=2.22 //x2=68.195 //y2=2.22
r1334 (  14 30 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=60.055 //y=2.22 //x2=59.94 //y2=2.22
r1335 (  13 32 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=67.965 //y=2.22 //x2=68.08 //y2=2.22
r1336 (  13 14 ) resistor r=7.54771 //w=0.131 //l=7.91 //layer=m1 \
 //thickness=0.36 //x=67.965 //y=2.22 //x2=60.055 //y2=2.22
r1337 (  12 28 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=45.995 //y=2.22 //x2=45.88 //y2=2.22
r1338 (  11 30 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=59.825 //y=2.22 //x2=59.94 //y2=2.22
r1339 (  11 12 ) resistor r=13.1966 //w=0.131 //l=13.83 //layer=m1 \
 //thickness=0.36 //x=59.825 //y=2.22 //x2=45.995 //y2=2.22
r1340 (  10 26 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=42.295 //y=2.22 //x2=42.18 //y2=2.22
r1341 (  9 28 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=45.765 //y=2.22 //x2=45.88 //y2=2.22
r1342 (  9 10 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=45.765 //y=2.22 //x2=42.295 //y2=2.22
r1343 (  8 24 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.155 //y=2.22 //x2=34.04 //y2=2.22
r1344 (  7 26 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=42.065 //y=2.22 //x2=42.18 //y2=2.22
r1345 (  7 8 ) resistor r=7.54771 //w=0.131 //l=7.91 //layer=m1 \
 //thickness=0.36 //x=42.065 //y=2.22 //x2=34.155 //y2=2.22
r1346 (  6 22 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.095 //y=2.22 //x2=19.98 //y2=2.22
r1347 (  5 24 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=33.925 //y=2.22 //x2=34.04 //y2=2.22
r1348 (  5 6 ) resistor r=13.1966 //w=0.131 //l=13.83 //layer=m1 \
 //thickness=0.36 //x=33.925 //y=2.22 //x2=20.095 //y2=2.22
r1349 (  4 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.395 //y=2.22 //x2=16.28 //y2=2.22
r1350 (  3 22 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=19.865 //y=2.22 //x2=19.98 //y2=2.22
r1351 (  3 4 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=19.865 //y=2.22 //x2=16.395 //y2=2.22
r1352 (  2 18 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.255 //y=2.22 //x2=8.14 //y2=2.22
r1353 (  1 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.165 //y=2.22 //x2=16.28 //y2=2.22
r1354 (  1 2 ) resistor r=7.54771 //w=0.131 //l=7.91 //layer=m1 \
 //thickness=0.36 //x=16.165 //y=2.22 //x2=8.255 //y2=2.22
ends PM_TMRDFFRNQNX1\%RN

subckt PM_TMRDFFRNQNX1\%noxref_16 ( 1 2 3 4 5 6 7 8 9 10 24 31 33 43 44 51 59 \
 65 66 70 77 78 85 93 99 100 104 106 113 115 121 122 123 124 127 128 129 130 \
 131 132 133 134 135 136 137 138 139 140 141 142 143 145 151 152 153 154 158 \
 159 160 165 167 169 175 176 177 178 179 180 184 186 189 190 194 195 196 201 \
 203 205 211 212 222 223 226 240 244 245 248 256 257 260 261 262 263 264 265 )
c500 ( 265 0 ) capacitor c=0.023087f //x=72.705 //y=5.02
c501 ( 264 0 ) capacitor c=0.023519f //x=71.825 //y=5.02
c502 ( 263 0 ) capacitor c=0.0224735f //x=70.945 //y=5.02
c503 ( 262 0 ) capacitor c=0.023087f //x=67.895 //y=5.02
c504 ( 261 0 ) capacitor c=0.023519f //x=67.015 //y=5.02
c505 ( 260 0 ) capacitor c=0.0224735f //x=66.135 //y=5.02
c506 ( 257 0 ) capacitor c=0.00872971f //x=72.955 //y=0.915
c507 ( 256 0 ) capacitor c=0.00853354f //x=68.145 //y=0.915
c508 ( 248 0 ) capacitor c=0.0340473f //x=76.25 //y=4.7
c509 ( 245 0 ) capacitor c=0.0292616f //x=76.22 //y=1.915
c510 ( 244 0 ) capacitor c=0.0436018f //x=76.22 //y=2.08
c511 ( 240 0 ) capacitor c=0.0602694f //x=75.48 //y=4.7
c512 ( 226 0 ) capacitor c=0.0331095f //x=63.3 //y=4.7
c513 ( 223 0 ) capacitor c=0.0279499f //x=63.27 //y=1.915
c514 ( 222 0 ) capacitor c=0.0421676f //x=63.27 //y=2.08
c515 ( 212 0 ) capacitor c=0.0431781f //x=76.785 //y=1.25
c516 ( 211 0 ) capacitor c=0.0197948f //x=76.785 //y=0.905
c517 ( 205 0 ) capacitor c=0.0158629f //x=76.63 //y=1.405
c518 ( 203 0 ) capacitor c=0.0157803f //x=76.63 //y=0.75
c519 ( 201 0 ) capacitor c=0.0307199f //x=76.625 //y=4.79
c520 ( 196 0 ) capacitor c=0.0210775f //x=76.255 //y=1.56
c521 ( 195 0 ) capacitor c=0.0179879f //x=76.255 //y=1.25
c522 ( 194 0 ) capacitor c=0.0177928f //x=76.255 //y=0.905
c523 ( 190 0 ) capacitor c=0.0338875f //x=75.815 //y=1.21
c524 ( 189 0 ) capacitor c=0.0189263f //x=75.815 //y=0.865
c525 ( 186 0 ) capacitor c=0.0141798f //x=75.66 //y=1.365
c526 ( 184 0 ) capacitor c=0.0149844f //x=75.66 //y=0.71
c527 ( 180 0 ) capacitor c=0.083929f //x=75.285 //y=1.915
c528 ( 179 0 ) capacitor c=0.0231111f //x=75.285 //y=1.52
c529 ( 178 0 ) capacitor c=0.0234352f //x=75.285 //y=1.21
c530 ( 177 0 ) capacitor c=0.0201338f //x=75.285 //y=0.865
c531 ( 176 0 ) capacitor c=0.0429696f //x=63.835 //y=1.25
c532 ( 175 0 ) capacitor c=0.0192208f //x=63.835 //y=0.905
c533 ( 169 0 ) capacitor c=0.0148884f //x=63.68 //y=1.405
c534 ( 167 0 ) capacitor c=0.0157803f //x=63.68 //y=0.75
c535 ( 165 0 ) capacitor c=0.0295235f //x=63.675 //y=4.79
c536 ( 160 0 ) capacitor c=0.0205163f //x=63.305 //y=1.56
c537 ( 159 0 ) capacitor c=0.0168481f //x=63.305 //y=1.25
c538 ( 158 0 ) capacitor c=0.0174783f //x=63.305 //y=0.905
c539 ( 154 0 ) capacitor c=0.0557698f //x=53.185 //y=4.79
c540 ( 153 0 ) capacitor c=0.0293157f //x=53.475 //y=4.79
c541 ( 152 0 ) capacitor c=0.0347816f //x=53.14 //y=1.22
c542 ( 151 0 ) capacitor c=0.0187487f //x=53.14 //y=0.875
c543 ( 145 0 ) capacitor c=0.0137055f //x=52.985 //y=1.375
c544 ( 143 0 ) capacitor c=0.0149861f //x=52.985 //y=0.72
c545 ( 142 0 ) capacitor c=0.096037f //x=52.61 //y=1.915
c546 ( 141 0 ) capacitor c=0.0228993f //x=52.61 //y=1.53
c547 ( 140 0 ) capacitor c=0.0234352f //x=52.61 //y=1.22
c548 ( 139 0 ) capacitor c=0.0198724f //x=52.61 //y=0.875
c549 ( 138 0 ) capacitor c=0.15358f //x=76.7 //y=6.02
c550 ( 137 0 ) capacitor c=0.116098f //x=76.26 //y=6.02
c551 ( 136 0 ) capacitor c=0.116091f //x=75.82 //y=6.02
c552 ( 135 0 ) capacitor c=0.154305f //x=75.38 //y=6.02
c553 ( 134 0 ) capacitor c=0.15358f //x=63.75 //y=6.02
c554 ( 133 0 ) capacitor c=0.110281f //x=63.31 //y=6.02
c555 ( 132 0 ) capacitor c=0.110114f //x=53.55 //y=6.02
c556 ( 131 0 ) capacitor c=0.158956f //x=53.11 //y=6.02
c557 ( 124 0 ) capacitor c=0.00116729f //x=72.85 //y=5.155
c558 ( 123 0 ) capacitor c=0.00226015f //x=71.97 //y=5.155
c559 ( 122 0 ) capacitor c=0.00116729f //x=68.04 //y=5.155
c560 ( 121 0 ) capacitor c=0.0021933f //x=67.16 //y=5.155
c561 ( 115 0 ) capacitor c=0.0711582f //x=76.22 //y=2.08
c562 ( 113 0 ) capacitor c=0.00453889f //x=76.22 //y=4.535
c563 ( 106 0 ) capacitor c=0.0883483f //x=75.48 //y=2.08
c564 ( 104 0 ) capacitor c=0.108107f //x=73.63 //y=4.07
c565 ( 100 0 ) capacitor c=0.00463522f //x=73.23 //y=1.665
c566 ( 99 0 ) capacitor c=0.0148737f //x=73.545 //y=1.665
c567 ( 93 0 ) capacitor c=0.0292981f //x=73.545 //y=5.155
c568 ( 85 0 ) capacitor c=0.0184197f //x=72.765 //y=5.155
c569 ( 78 0 ) capacitor c=0.00351598f //x=71.175 //y=5.155
c570 ( 77 0 ) capacitor c=0.0155255f //x=71.885 //y=5.155
c571 ( 70 0 ) capacitor c=0.106966f //x=68.82 //y=4.07
c572 ( 66 0 ) capacitor c=0.00398962f //x=68.42 //y=1.665
c573 ( 65 0 ) capacitor c=0.0137288f //x=68.735 //y=1.665
c574 ( 59 0 ) capacitor c=0.0291076f //x=68.735 //y=5.155
c575 ( 51 0 ) capacitor c=0.0184197f //x=67.955 //y=5.155
c576 ( 44 0 ) capacitor c=0.00332903f //x=66.365 //y=5.155
c577 ( 43 0 ) capacitor c=0.014837f //x=67.075 //y=5.155
c578 ( 33 0 ) capacitor c=0.0693025f //x=63.27 //y=2.08
c579 ( 31 0 ) capacitor c=0.00453889f //x=63.27 //y=4.535
c580 ( 24 0 ) capacitor c=0.0974753f //x=52.91 //y=2.08
c581 ( 10 0 ) capacitor c=0.00400147f //x=75.595 //y=4.07
c582 ( 9 0 ) capacitor c=0.0236326f //x=76.105 //y=4.07
c583 ( 8 0 ) capacitor c=0.00570859f //x=73.745 //y=4.07
c584 ( 7 0 ) capacitor c=0.0482058f //x=75.365 //y=4.07
c585 ( 6 0 ) capacitor c=0.00720076f //x=68.935 //y=4.07
c586 ( 5 0 ) capacitor c=0.124606f //x=73.515 //y=4.07
c587 ( 4 0 ) capacitor c=0.00557292f //x=63.385 //y=4.07
c588 ( 3 0 ) capacitor c=0.0897132f //x=68.705 //y=4.07
c589 ( 2 0 ) capacitor c=0.00985259f //x=53.025 //y=4.07
c590 ( 1 0 ) capacitor c=0.145635f //x=63.155 //y=4.07
r591 (  250 251 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=76.25 //y=4.79 //x2=76.25 //y2=4.865
r592 (  248 250 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=76.25 //y=4.7 //x2=76.25 //y2=4.79
r593 (  244 245 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=76.22 //y=2.08 //x2=76.22 //y2=1.915
r594 (  238 240 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=75.38 //y=4.7 //x2=75.48 //y2=4.7
r595 (  228 229 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=63.3 //y=4.79 //x2=63.3 //y2=4.865
r596 (  226 228 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=63.3 //y=4.7 //x2=63.3 //y2=4.79
r597 (  222 223 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=63.27 //y=2.08 //x2=63.27 //y2=1.915
r598 (  212 255 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=76.785 //y=1.25 //x2=76.745 //y2=1.405
r599 (  211 254 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=76.785 //y=0.905 //x2=76.745 //y2=0.75
r600 (  211 212 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=76.785 //y=0.905 //x2=76.785 //y2=1.25
r601 (  206 253 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=76.41 //y=1.405 //x2=76.295 //y2=1.405
r602 (  205 255 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=76.63 //y=1.405 //x2=76.745 //y2=1.405
r603 (  204 252 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=76.41 //y=0.75 //x2=76.295 //y2=0.75
r604 (  203 254 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=76.63 //y=0.75 //x2=76.745 //y2=0.75
r605 (  203 204 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=76.63 //y=0.75 //x2=76.41 //y2=0.75
r606 (  202 250 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=76.385 //y=4.79 //x2=76.25 //y2=4.79
r607 (  201 208 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=76.625 //y=4.79 //x2=76.7 //y2=4.865
r608 (  201 202 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=76.625 //y=4.79 //x2=76.385 //y2=4.79
r609 (  196 253 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=76.255 //y=1.56 //x2=76.295 //y2=1.405
r610 (  196 245 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=76.255 //y=1.56 //x2=76.255 //y2=1.915
r611 (  195 253 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=76.255 //y=1.25 //x2=76.295 //y2=1.405
r612 (  194 252 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=76.255 //y=0.905 //x2=76.295 //y2=0.75
r613 (  194 195 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=76.255 //y=0.905 //x2=76.255 //y2=1.25
r614 (  191 240 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=75.82 //y=4.865 //x2=75.48 //y2=4.7
r615 (  190 242 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.815 //y=1.21 //x2=75.775 //y2=1.365
r616 (  189 241 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.815 //y=0.865 //x2=75.775 //y2=0.71
r617 (  189 190 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=75.815 //y=0.865 //x2=75.815 //y2=1.21
r618 (  187 237 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.44 //y=1.365 //x2=75.325 //y2=1.365
r619 (  186 242 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.66 //y=1.365 //x2=75.775 //y2=1.365
r620 (  185 236 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.44 //y=0.71 //x2=75.325 //y2=0.71
r621 (  184 241 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.66 //y=0.71 //x2=75.775 //y2=0.71
r622 (  184 185 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=75.66 //y=0.71 //x2=75.44 //y2=0.71
r623 (  181 238 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=75.38 //y=4.865 //x2=75.38 //y2=4.7
r624 (  180 235 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=75.285 //y=1.915 //x2=75.48 //y2=2.08
r625 (  179 237 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.285 //y=1.52 //x2=75.325 //y2=1.365
r626 (  179 180 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=75.285 //y=1.52 //x2=75.285 //y2=1.915
r627 (  178 237 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.285 //y=1.21 //x2=75.325 //y2=1.365
r628 (  177 236 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.285 //y=0.865 //x2=75.325 //y2=0.71
r629 (  177 178 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=75.285 //y=0.865 //x2=75.285 //y2=1.21
r630 (  176 233 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.835 //y=1.25 //x2=63.795 //y2=1.405
r631 (  175 232 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.835 //y=0.905 //x2=63.795 //y2=0.75
r632 (  175 176 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=63.835 //y=0.905 //x2=63.835 //y2=1.25
r633 (  170 231 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.46 //y=1.405 //x2=63.345 //y2=1.405
r634 (  169 233 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.68 //y=1.405 //x2=63.795 //y2=1.405
r635 (  168 230 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.46 //y=0.75 //x2=63.345 //y2=0.75
r636 (  167 232 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.68 //y=0.75 //x2=63.795 //y2=0.75
r637 (  167 168 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=63.68 //y=0.75 //x2=63.46 //y2=0.75
r638 (  166 228 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=63.435 //y=4.79 //x2=63.3 //y2=4.79
r639 (  165 172 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=63.675 //y=4.79 //x2=63.75 //y2=4.865
r640 (  165 166 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=63.675 //y=4.79 //x2=63.435 //y2=4.79
r641 (  160 231 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.305 //y=1.56 //x2=63.345 //y2=1.405
r642 (  160 223 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=63.305 //y=1.56 //x2=63.305 //y2=1.915
r643 (  159 231 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.305 //y=1.25 //x2=63.345 //y2=1.405
r644 (  158 230 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.305 //y=0.905 //x2=63.345 //y2=0.75
r645 (  158 159 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=63.305 //y=0.905 //x2=63.305 //y2=1.25
r646 (  153 155 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=53.475 //y=4.79 //x2=53.55 //y2=4.865
r647 (  153 154 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=53.475 //y=4.79 //x2=53.185 //y2=4.79
r648 (  152 220 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.14 //y=1.22 //x2=53.1 //y2=1.375
r649 (  151 219 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.14 //y=0.875 //x2=53.1 //y2=0.72
r650 (  151 152 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=53.14 //y=0.875 //x2=53.14 //y2=1.22
r651 (  148 154 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=53.11 //y=4.865 //x2=53.185 //y2=4.79
r652 (  148 218 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=53.11 //y=4.865 //x2=52.91 //y2=4.7
r653 (  146 214 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=52.765 //y=1.375 //x2=52.65 //y2=1.375
r654 (  145 220 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=52.985 //y=1.375 //x2=53.1 //y2=1.375
r655 (  144 213 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=52.765 //y=0.72 //x2=52.65 //y2=0.72
r656 (  143 219 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=52.985 //y=0.72 //x2=53.1 //y2=0.72
r657 (  143 144 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=52.985 //y=0.72 //x2=52.765 //y2=0.72
r658 (  142 216 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=52.61 //y=1.915 //x2=52.91 //y2=2.08
r659 (  141 214 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.61 //y=1.53 //x2=52.65 //y2=1.375
r660 (  141 142 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=52.61 //y=1.53 //x2=52.61 //y2=1.915
r661 (  140 214 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.61 //y=1.22 //x2=52.65 //y2=1.375
r662 (  139 213 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.61 //y=0.875 //x2=52.65 //y2=0.72
r663 (  139 140 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=52.61 //y=0.875 //x2=52.61 //y2=1.22
r664 (  138 208 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=76.7 //y=6.02 //x2=76.7 //y2=4.865
r665 (  137 251 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=76.26 //y=6.02 //x2=76.26 //y2=4.865
r666 (  136 191 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=75.82 //y=6.02 //x2=75.82 //y2=4.865
r667 (  135 181 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=75.38 //y=6.02 //x2=75.38 //y2=4.865
r668 (  134 172 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=63.75 //y=6.02 //x2=63.75 //y2=4.865
r669 (  133 229 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=63.31 //y=6.02 //x2=63.31 //y2=4.865
r670 (  132 155 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=53.55 //y=6.02 //x2=53.55 //y2=4.865
r671 (  131 148 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=53.11 //y=6.02 //x2=53.11 //y2=4.865
r672 (  130 205 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=76.52 //y=1.405 //x2=76.63 //y2=1.405
r673 (  130 206 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=76.52 //y=1.405 //x2=76.41 //y2=1.405
r674 (  129 186 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=75.55 //y=1.365 //x2=75.66 //y2=1.365
r675 (  129 187 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=75.55 //y=1.365 //x2=75.44 //y2=1.365
r676 (  128 169 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=63.57 //y=1.405 //x2=63.68 //y2=1.405
r677 (  128 170 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=63.57 //y=1.405 //x2=63.46 //y2=1.405
r678 (  127 145 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=52.875 //y=1.375 //x2=52.985 //y2=1.375
r679 (  127 146 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=52.875 //y=1.375 //x2=52.765 //y2=1.375
r680 (  126 248 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=76.25 //y=4.7 //x2=76.25 //y2=4.7
r681 (  120 226 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=63.3 //y=4.7 //x2=63.3 //y2=4.7
r682 (  115 244 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=76.22 //y=2.08 //x2=76.22 //y2=2.08
r683 (  115 118 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=76.22 //y=2.08 //x2=76.22 //y2=4.07
r684 (  113 126 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=76.22 //y=4.535 //x2=76.235 //y2=4.7
r685 (  113 118 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=76.22 //y=4.535 //x2=76.22 //y2=4.07
r686 (  111 240 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=75.48 //y=4.7 //x2=75.48 //y2=4.7
r687 (  109 111 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=75.48 //y=4.07 //x2=75.48 //y2=4.7
r688 (  106 235 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=75.48 //y=2.08 //x2=75.48 //y2=2.08
r689 (  106 109 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=75.48 //y=2.08 //x2=75.48 //y2=4.07
r690 (  102 104 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li \
 //thickness=0.1 //x=73.63 //y=5.07 //x2=73.63 //y2=4.07
r691 (  101 104 ) resistor r=158.802 //w=0.187 //l=2.32 //layer=li \
 //thickness=0.1 //x=73.63 //y=1.75 //x2=73.63 //y2=4.07
r692 (  99 101 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=73.545 //y=1.665 //x2=73.63 //y2=1.75
r693 (  99 100 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=73.545 //y=1.665 //x2=73.23 //y2=1.665
r694 (  95 100 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=73.145 //y=1.58 //x2=73.23 //y2=1.665
r695 (  95 257 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=73.145 //y=1.58 //x2=73.145 //y2=1.01
r696 (  94 124 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.935 //y=5.155 //x2=72.85 //y2=5.155
r697 (  93 102 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=73.545 //y=5.155 //x2=73.63 //y2=5.07
r698 (  93 94 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=73.545 //y=5.155 //x2=72.935 //y2=5.155
r699 (  87 124 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.85 //y=5.24 //x2=72.85 //y2=5.155
r700 (  87 265 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=72.85 //y=5.24 //x2=72.85 //y2=5.725
r701 (  86 123 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.055 //y=5.155 //x2=71.97 //y2=5.155
r702 (  85 124 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.765 //y=5.155 //x2=72.85 //y2=5.155
r703 (  85 86 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=72.765 //y=5.155 //x2=72.055 //y2=5.155
r704 (  79 123 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.97 //y=5.24 //x2=71.97 //y2=5.155
r705 (  79 264 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=71.97 //y=5.24 //x2=71.97 //y2=5.725
r706 (  77 123 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.885 //y=5.155 //x2=71.97 //y2=5.155
r707 (  77 78 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=71.885 //y=5.155 //x2=71.175 //y2=5.155
r708 (  71 78 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=71.09 //y=5.24 //x2=71.175 //y2=5.155
r709 (  71 263 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=71.09 //y=5.24 //x2=71.09 //y2=5.725
r710 (  68 70 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=68.82 //y=5.07 //x2=68.82 //y2=4.07
r711 (  67 70 ) resistor r=158.802 //w=0.187 //l=2.32 //layer=li \
 //thickness=0.1 //x=68.82 //y=1.75 //x2=68.82 //y2=4.07
r712 (  65 67 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=68.735 //y=1.665 //x2=68.82 //y2=1.75
r713 (  65 66 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=68.735 //y=1.665 //x2=68.42 //y2=1.665
r714 (  61 66 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=68.335 //y=1.58 //x2=68.42 //y2=1.665
r715 (  61 256 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=68.335 //y=1.58 //x2=68.335 //y2=1.01
r716 (  60 122 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.125 //y=5.155 //x2=68.04 //y2=5.155
r717 (  59 68 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=68.735 //y=5.155 //x2=68.82 //y2=5.07
r718 (  59 60 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=68.735 //y=5.155 //x2=68.125 //y2=5.155
r719 (  53 122 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=68.04 //y=5.24 //x2=68.04 //y2=5.155
r720 (  53 262 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=68.04 //y=5.24 //x2=68.04 //y2=5.725
r721 (  52 121 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.245 //y=5.155 //x2=67.16 //y2=5.155
r722 (  51 122 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.955 //y=5.155 //x2=68.04 //y2=5.155
r723 (  51 52 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=67.955 //y=5.155 //x2=67.245 //y2=5.155
r724 (  45 121 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.16 //y=5.24 //x2=67.16 //y2=5.155
r725 (  45 261 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=67.16 //y=5.24 //x2=67.16 //y2=5.725
r726 (  43 121 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.075 //y=5.155 //x2=67.16 //y2=5.155
r727 (  43 44 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=67.075 //y=5.155 //x2=66.365 //y2=5.155
r728 (  37 44 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=66.28 //y=5.24 //x2=66.365 //y2=5.155
r729 (  37 260 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=66.28 //y=5.24 //x2=66.28 //y2=5.725
r730 (  33 222 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=63.27 //y=2.08 //x2=63.27 //y2=2.08
r731 (  33 36 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=63.27 //y=2.08 //x2=63.27 //y2=4.07
r732 (  31 120 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=63.27 //y=4.535 //x2=63.285 //y2=4.7
r733 (  31 36 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=63.27 //y=4.535 //x2=63.27 //y2=4.07
r734 (  29 218 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=52.91 //y=4.7 //x2=52.91 //y2=4.7
r735 (  27 29 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=52.91 //y=4.07 //x2=52.91 //y2=4.7
r736 (  24 216 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=52.91 //y=2.08 //x2=52.91 //y2=2.08
r737 (  24 27 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=52.91 //y=2.08 //x2=52.91 //y2=4.07
r738 (  22 118 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=76.22 //y=4.07 //x2=76.22 //y2=4.07
r739 (  20 109 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=75.48 //y=4.07 //x2=75.48 //y2=4.07
r740 (  18 104 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=73.63 //y=4.07 //x2=73.63 //y2=4.07
r741 (  16 70 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=68.82 //y=4.07 //x2=68.82 //y2=4.07
r742 (  14 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=63.27 //y=4.07 //x2=63.27 //y2=4.07
r743 (  12 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=52.91 //y=4.07 //x2=52.91 //y2=4.07
r744 (  10 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=75.595 //y=4.07 //x2=75.48 //y2=4.07
r745 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=76.105 //y=4.07 //x2=76.22 //y2=4.07
r746 (  9 10 ) resistor r=0.486641 //w=0.131 //l=0.51 //layer=m1 \
 //thickness=0.36 //x=76.105 //y=4.07 //x2=75.595 //y2=4.07
r747 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=73.745 //y=4.07 //x2=73.63 //y2=4.07
r748 (  7 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=75.365 //y=4.07 //x2=75.48 //y2=4.07
r749 (  7 8 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=75.365 //y=4.07 //x2=73.745 //y2=4.07
r750 (  6 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=68.935 //y=4.07 //x2=68.82 //y2=4.07
r751 (  5 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=73.515 //y=4.07 //x2=73.63 //y2=4.07
r752 (  5 6 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=73.515 //y=4.07 //x2=68.935 //y2=4.07
r753 (  4 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=63.385 //y=4.07 //x2=63.27 //y2=4.07
r754 (  3 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=68.705 //y=4.07 //x2=68.82 //y2=4.07
r755 (  3 4 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=68.705 //y=4.07 //x2=63.385 //y2=4.07
r756 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=53.025 //y=4.07 //x2=52.91 //y2=4.07
r757 (  1 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=63.155 //y=4.07 //x2=63.27 //y2=4.07
r758 (  1 2 ) resistor r=9.66603 //w=0.131 //l=10.13 //layer=m1 \
 //thickness=0.36 //x=63.155 //y=4.07 //x2=53.025 //y2=4.07
ends PM_TMRDFFRNQNX1\%noxref_16

subckt PM_TMRDFFRNQNX1\%noxref_17 ( 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 38 \
 51 52 63 65 66 70 72 85 86 93 101 107 108 112 114 127 128 139 141 142 146 148 \
 156 166 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 189 \
 190 191 192 193 194 198 199 200 205 207 210 211 215 216 217 222 224 227 228 \
 229 230 231 232 236 238 241 242 246 247 248 249 250 252 258 259 260 261 265 \
 266 267 268 272 274 277 278 279 280 284 285 286 287 291 293 299 300 302 303 \
 308 312 313 318 327 339 352 355 356 357 361 362 363 364 365 366 367 )
c763 ( 367 0 ) capacitor c=0.0220291f //x=63.385 //y=5.02
c764 ( 366 0 ) capacitor c=0.0217503f //x=62.505 //y=5.02
c765 ( 365 0 ) capacitor c=0.023087f //x=59.755 //y=5.02
c766 ( 364 0 ) capacitor c=0.023519f //x=58.875 //y=5.02
c767 ( 363 0 ) capacitor c=0.0224735f //x=57.995 //y=5.02
c768 ( 362 0 ) capacitor c=0.0220291f //x=50.435 //y=5.02
c769 ( 361 0 ) capacitor c=0.0217503f //x=49.555 //y=5.02
c770 ( 357 0 ) capacitor c=0.0084702f //x=63.38 //y=0.905
c771 ( 356 0 ) capacitor c=0.00872971f //x=60.005 //y=0.915
c772 ( 355 0 ) capacitor c=0.0084702f //x=50.43 //y=0.905
c773 ( 352 0 ) capacitor c=0.0655948f //x=82.14 //y=4.705
c774 ( 339 0 ) capacitor c=0.0545009f //x=78.44 //y=2.08
c775 ( 327 0 ) capacitor c=0.0588816f //x=62.53 //y=4.7
c776 ( 318 0 ) capacitor c=0.058931f //x=55.13 //y=4.7
c777 ( 313 0 ) capacitor c=0.0273931f //x=55.13 //y=1.915
c778 ( 312 0 ) capacitor c=0.0456313f //x=55.13 //y=2.08
c779 ( 308 0 ) capacitor c=0.0587755f //x=46.99 //y=4.7
c780 ( 303 0 ) capacitor c=0.0273931f //x=46.99 //y=1.915
c781 ( 302 0 ) capacitor c=0.0456313f //x=46.99 //y=2.08
c782 ( 300 0 ) capacitor c=0.0342409f //x=82.475 //y=1.21
c783 ( 299 0 ) capacitor c=0.0187384f //x=82.475 //y=0.865
c784 ( 293 0 ) capacitor c=0.0141797f //x=82.32 //y=1.365
c785 ( 291 0 ) capacitor c=0.0149844f //x=82.32 //y=0.71
c786 ( 287 0 ) capacitor c=0.0979048f //x=81.945 //y=1.915
c787 ( 286 0 ) capacitor c=0.0225105f //x=81.945 //y=1.52
c788 ( 285 0 ) capacitor c=0.0234376f //x=81.945 //y=1.21
c789 ( 284 0 ) capacitor c=0.0199343f //x=81.945 //y=0.865
c790 ( 280 0 ) capacitor c=0.0318948f //x=79.145 //y=1.21
c791 ( 279 0 ) capacitor c=0.0187384f //x=79.145 //y=0.865
c792 ( 278 0 ) capacitor c=0.0606536f //x=78.785 //y=4.795
c793 ( 277 0 ) capacitor c=0.0292043f //x=79.075 //y=4.795
c794 ( 274 0 ) capacitor c=0.0157913f //x=78.99 //y=1.365
c795 ( 272 0 ) capacitor c=0.0149844f //x=78.99 //y=0.71
c796 ( 268 0 ) capacitor c=0.0302441f //x=78.615 //y=1.915
c797 ( 267 0 ) capacitor c=0.0238107f //x=78.615 //y=1.52
c798 ( 266 0 ) capacitor c=0.0234352f //x=78.615 //y=1.21
c799 ( 265 0 ) capacitor c=0.0199931f //x=78.615 //y=0.865
c800 ( 261 0 ) capacitor c=0.0556143f //x=66.135 //y=4.79
c801 ( 260 0 ) capacitor c=0.0293157f //x=66.425 //y=4.79
c802 ( 259 0 ) capacitor c=0.0347816f //x=66.09 //y=1.22
c803 ( 258 0 ) capacitor c=0.0187487f //x=66.09 //y=0.875
c804 ( 252 0 ) capacitor c=0.0137055f //x=65.935 //y=1.375
c805 ( 250 0 ) capacitor c=0.0149861f //x=65.935 //y=0.72
c806 ( 249 0 ) capacitor c=0.096037f //x=65.56 //y=1.915
c807 ( 248 0 ) capacitor c=0.0228993f //x=65.56 //y=1.53
c808 ( 247 0 ) capacitor c=0.0234352f //x=65.56 //y=1.22
c809 ( 246 0 ) capacitor c=0.0198724f //x=65.56 //y=0.875
c810 ( 242 0 ) capacitor c=0.0318948f //x=62.865 //y=1.21
c811 ( 241 0 ) capacitor c=0.0187384f //x=62.865 //y=0.865
c812 ( 238 0 ) capacitor c=0.0141798f //x=62.71 //y=1.365
c813 ( 236 0 ) capacitor c=0.0149844f //x=62.71 //y=0.71
c814 ( 232 0 ) capacitor c=0.0813322f //x=62.335 //y=1.915
c815 ( 231 0 ) capacitor c=0.0229267f //x=62.335 //y=1.52
c816 ( 230 0 ) capacitor c=0.0234352f //x=62.335 //y=1.21
c817 ( 229 0 ) capacitor c=0.0199343f //x=62.335 //y=0.865
c818 ( 228 0 ) capacitor c=0.0432517f //x=55.65 //y=1.26
c819 ( 227 0 ) capacitor c=0.0200379f //x=55.65 //y=0.915
c820 ( 224 0 ) capacitor c=0.0148873f //x=55.495 //y=1.415
c821 ( 222 0 ) capacitor c=0.0157803f //x=55.495 //y=0.76
c822 ( 217 0 ) capacitor c=0.0218028f //x=55.12 //y=1.57
c823 ( 216 0 ) capacitor c=0.0207459f //x=55.12 //y=1.26
c824 ( 215 0 ) capacitor c=0.0194308f //x=55.12 //y=0.915
c825 ( 211 0 ) capacitor c=0.0432517f //x=47.51 //y=1.26
c826 ( 210 0 ) capacitor c=0.0200379f //x=47.51 //y=0.915
c827 ( 207 0 ) capacitor c=0.0148873f //x=47.355 //y=1.415
c828 ( 205 0 ) capacitor c=0.0157803f //x=47.355 //y=0.76
c829 ( 200 0 ) capacitor c=0.0218028f //x=46.98 //y=1.57
c830 ( 199 0 ) capacitor c=0.0207459f //x=46.98 //y=1.26
c831 ( 198 0 ) capacitor c=0.0194308f //x=46.98 //y=0.915
c832 ( 194 0 ) capacitor c=0.110336f //x=82.47 //y=6.025
c833 ( 193 0 ) capacitor c=0.154049f //x=82.03 //y=6.025
c834 ( 192 0 ) capacitor c=0.110003f //x=79.15 //y=6.025
c835 ( 191 0 ) capacitor c=0.15424f //x=78.71 //y=6.025
c836 ( 190 0 ) capacitor c=0.110114f //x=66.5 //y=6.02
c837 ( 189 0 ) capacitor c=0.158956f //x=66.06 //y=6.02
c838 ( 188 0 ) capacitor c=0.110275f //x=62.87 //y=6.02
c839 ( 187 0 ) capacitor c=0.154305f //x=62.43 //y=6.02
c840 ( 186 0 ) capacitor c=0.158794f //x=55.31 //y=6.02
c841 ( 185 0 ) capacitor c=0.110114f //x=54.87 //y=6.02
c842 ( 184 0 ) capacitor c=0.158794f //x=47.17 //y=6.02
c843 ( 183 0 ) capacitor c=0.110114f //x=46.73 //y=6.02
c844 ( 176 0 ) capacitor c=0.00211606f //x=63.53 //y=5.2
c845 ( 175 0 ) capacitor c=0.00106608f //x=59.9 //y=5.155
c846 ( 174 0 ) capacitor c=0.00207319f //x=59.02 //y=5.155
c847 ( 173 0 ) capacitor c=0.00211606f //x=50.58 //y=5.2
c848 ( 166 0 ) capacitor c=0.117496f //x=82.14 //y=2.08
c849 ( 156 0 ) capacitor c=0.0945553f //x=78.44 //y=2.08
c850 ( 148 0 ) capacitor c=0.096212f //x=65.86 //y=2.08
c851 ( 146 0 ) capacitor c=0.104337f //x=64.01 //y=3.33
c852 ( 142 0 ) capacitor c=0.00404073f //x=63.655 //y=1.655
c853 ( 141 0 ) capacitor c=0.0122201f //x=63.925 //y=1.655
c854 ( 139 0 ) capacitor c=0.0137995f //x=63.925 //y=5.2
c855 ( 128 0 ) capacitor c=0.00249378f //x=62.735 //y=5.2
c856 ( 127 0 ) capacitor c=0.0143649f //x=63.445 //y=5.2
c857 ( 114 0 ) capacitor c=0.0860657f //x=62.53 //y=2.08
c858 ( 112 0 ) capacitor c=0.105397f //x=60.68 //y=3.33
c859 ( 108 0 ) capacitor c=0.00398962f //x=60.28 //y=1.665
c860 ( 107 0 ) capacitor c=0.0137288f //x=60.595 //y=1.665
c861 ( 101 0 ) capacitor c=0.0284518f //x=60.595 //y=5.155
c862 ( 93 0 ) capacitor c=0.0176454f //x=59.815 //y=5.155
c863 ( 86 0 ) capacitor c=0.00332903f //x=58.225 //y=5.155
c864 ( 85 0 ) capacitor c=0.0148427f //x=58.935 //y=5.155
c865 ( 72 0 ) capacitor c=0.081384f //x=55.13 //y=2.08
c866 ( 70 0 ) capacitor c=0.106559f //x=51.06 //y=3.33
c867 ( 66 0 ) capacitor c=0.00404073f //x=50.705 //y=1.655
c868 ( 65 0 ) capacitor c=0.0122201f //x=50.975 //y=1.655
c869 ( 63 0 ) capacitor c=0.0137995f //x=50.975 //y=5.2
c870 ( 52 0 ) capacitor c=0.00251635f //x=49.785 //y=5.2
c871 ( 51 0 ) capacitor c=0.0143649f //x=50.495 //y=5.2
c872 ( 38 0 ) capacitor c=0.0811555f //x=46.99 //y=2.08
c873 ( 16 0 ) capacitor c=0.0152968f //x=78.555 //y=4.44
c874 ( 15 0 ) capacitor c=0.0828557f //x=82.025 //y=4.44
c875 ( 14 0 ) capacitor c=0.004304f //x=65.975 //y=3.33
c876 ( 13 0 ) capacitor c=0.195727f //x=78.325 //y=3.33
c877 ( 12 0 ) capacitor c=0.00246264f //x=64.125 //y=3.33
c878 ( 11 0 ) capacitor c=0.0280612f //x=65.745 //y=3.33
c879 ( 10 0 ) capacitor c=0.00253051f //x=62.645 //y=3.33
c880 ( 9 0 ) capacitor c=0.0166351f //x=63.895 //y=3.33
c881 ( 8 0 ) capacitor c=0.00424937f //x=60.795 //y=3.33
c882 ( 7 0 ) capacitor c=0.0279453f //x=62.415 //y=3.33
c883 ( 6 0 ) capacitor c=0.00458481f //x=55.245 //y=3.33
c884 ( 5 0 ) capacitor c=0.077708f //x=60.565 //y=3.33
c885 ( 4 0 ) capacitor c=0.00376077f //x=51.175 //y=3.33
c886 ( 3 0 ) capacitor c=0.0767635f //x=55.015 //y=3.33
c887 ( 2 0 ) capacitor c=0.0127233f //x=47.105 //y=3.33
c888 ( 1 0 ) capacitor c=0.060553f //x=50.945 //y=3.33
r889 (  350 352 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=82.03 //y=4.705 //x2=82.14 //y2=4.705
r890 (  325 327 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=62.43 //y=4.7 //x2=62.53 //y2=4.7
r891 (  312 313 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=55.13 //y=2.08 //x2=55.13 //y2=1.915
r892 (  302 303 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=46.99 //y=2.08 //x2=46.99 //y2=1.915
r893 (  300 354 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=82.475 //y=1.21 //x2=82.435 //y2=1.365
r894 (  299 353 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=82.475 //y=0.865 //x2=82.435 //y2=0.71
r895 (  299 300 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=82.475 //y=0.865 //x2=82.475 //y2=1.21
r896 (  296 352 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=82.47 //y=4.87 //x2=82.14 //y2=4.705
r897 (  294 349 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.1 //y=1.365 //x2=81.985 //y2=1.365
r898 (  293 354 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.32 //y=1.365 //x2=82.435 //y2=1.365
r899 (  292 348 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.1 //y=0.71 //x2=81.985 //y2=0.71
r900 (  291 353 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.32 //y=0.71 //x2=82.435 //y2=0.71
r901 (  291 292 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=82.32 //y=0.71 //x2=82.1 //y2=0.71
r902 (  288 350 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=82.03 //y=4.87 //x2=82.03 //y2=4.705
r903 (  287 347 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=81.945 //y=1.915 //x2=82.14 //y2=2.08
r904 (  286 349 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=81.945 //y=1.52 //x2=81.985 //y2=1.365
r905 (  286 287 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=81.945 //y=1.52 //x2=81.945 //y2=1.915
r906 (  285 349 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=81.945 //y=1.21 //x2=81.985 //y2=1.365
r907 (  284 348 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=81.945 //y=0.865 //x2=81.985 //y2=0.71
r908 (  284 285 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=81.945 //y=0.865 //x2=81.945 //y2=1.21
r909 (  280 345 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.145 //y=1.21 //x2=79.105 //y2=1.365
r910 (  279 344 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.145 //y=0.865 //x2=79.105 //y2=0.71
r911 (  279 280 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=79.145 //y=0.865 //x2=79.145 //y2=1.21
r912 (  277 281 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=79.075 //y=4.795 //x2=79.15 //y2=4.87
r913 (  277 278 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=79.075 //y=4.795 //x2=78.785 //y2=4.795
r914 (  275 343 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.77 //y=1.365 //x2=78.655 //y2=1.365
r915 (  274 345 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.99 //y=1.365 //x2=79.105 //y2=1.365
r916 (  273 342 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.77 //y=0.71 //x2=78.655 //y2=0.71
r917 (  272 344 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.99 //y=0.71 //x2=79.105 //y2=0.71
r918 (  272 273 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=78.99 //y=0.71 //x2=78.77 //y2=0.71
r919 (  269 278 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=78.71 //y=4.87 //x2=78.785 //y2=4.795
r920 (  269 341 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=78.71 //y=4.87 //x2=78.44 //y2=4.705
r921 (  268 339 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=78.615 //y=1.915 //x2=78.44 //y2=2.08
r922 (  267 343 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.615 //y=1.52 //x2=78.655 //y2=1.365
r923 (  267 268 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=78.615 //y=1.52 //x2=78.615 //y2=1.915
r924 (  266 343 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.615 //y=1.21 //x2=78.655 //y2=1.365
r925 (  265 342 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.615 //y=0.865 //x2=78.655 //y2=0.71
r926 (  265 266 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=78.615 //y=0.865 //x2=78.615 //y2=1.21
r927 (  260 262 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=66.425 //y=4.79 //x2=66.5 //y2=4.865
r928 (  260 261 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=66.425 //y=4.79 //x2=66.135 //y2=4.79
r929 (  259 337 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.09 //y=1.22 //x2=66.05 //y2=1.375
r930 (  258 336 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.09 //y=0.875 //x2=66.05 //y2=0.72
r931 (  258 259 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=66.09 //y=0.875 //x2=66.09 //y2=1.22
r932 (  255 261 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=66.06 //y=4.865 //x2=66.135 //y2=4.79
r933 (  255 335 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=66.06 //y=4.865 //x2=65.86 //y2=4.7
r934 (  253 331 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=65.715 //y=1.375 //x2=65.6 //y2=1.375
r935 (  252 337 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=65.935 //y=1.375 //x2=66.05 //y2=1.375
r936 (  251 330 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=65.715 //y=0.72 //x2=65.6 //y2=0.72
r937 (  250 336 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=65.935 //y=0.72 //x2=66.05 //y2=0.72
r938 (  250 251 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=65.935 //y=0.72 //x2=65.715 //y2=0.72
r939 (  249 333 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=65.56 //y=1.915 //x2=65.86 //y2=2.08
r940 (  248 331 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.56 //y=1.53 //x2=65.6 //y2=1.375
r941 (  248 249 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=65.56 //y=1.53 //x2=65.56 //y2=1.915
r942 (  247 331 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.56 //y=1.22 //x2=65.6 //y2=1.375
r943 (  246 330 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=65.56 //y=0.875 //x2=65.6 //y2=0.72
r944 (  246 247 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=65.56 //y=0.875 //x2=65.56 //y2=1.22
r945 (  243 327 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=62.87 //y=4.865 //x2=62.53 //y2=4.7
r946 (  242 329 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.865 //y=1.21 //x2=62.825 //y2=1.365
r947 (  241 328 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.865 //y=0.865 //x2=62.825 //y2=0.71
r948 (  241 242 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=62.865 //y=0.865 //x2=62.865 //y2=1.21
r949 (  239 324 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=62.49 //y=1.365 //x2=62.375 //y2=1.365
r950 (  238 329 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=62.71 //y=1.365 //x2=62.825 //y2=1.365
r951 (  237 323 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=62.49 //y=0.71 //x2=62.375 //y2=0.71
r952 (  236 328 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=62.71 //y=0.71 //x2=62.825 //y2=0.71
r953 (  236 237 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=62.71 //y=0.71 //x2=62.49 //y2=0.71
r954 (  233 325 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=62.43 //y=4.865 //x2=62.43 //y2=4.7
r955 (  232 322 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=62.335 //y=1.915 //x2=62.53 //y2=2.08
r956 (  231 324 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.335 //y=1.52 //x2=62.375 //y2=1.365
r957 (  231 232 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=62.335 //y=1.52 //x2=62.335 //y2=1.915
r958 (  230 324 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.335 //y=1.21 //x2=62.375 //y2=1.365
r959 (  229 323 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.335 //y=0.865 //x2=62.375 //y2=0.71
r960 (  229 230 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=62.335 //y=0.865 //x2=62.335 //y2=1.21
r961 (  228 320 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.65 //y=1.26 //x2=55.61 //y2=1.415
r962 (  227 319 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.65 //y=0.915 //x2=55.61 //y2=0.76
r963 (  227 228 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=55.65 //y=0.915 //x2=55.65 //y2=1.26
r964 (  225 316 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.275 //y=1.415 //x2=55.16 //y2=1.415
r965 (  224 320 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.495 //y=1.415 //x2=55.61 //y2=1.415
r966 (  223 315 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.275 //y=0.76 //x2=55.16 //y2=0.76
r967 (  222 319 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.495 //y=0.76 //x2=55.61 //y2=0.76
r968 (  222 223 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=55.495 //y=0.76 //x2=55.275 //y2=0.76
r969 (  219 318 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=55.31 //y=4.865 //x2=55.13 //y2=4.7
r970 (  217 316 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.12 //y=1.57 //x2=55.16 //y2=1.415
r971 (  217 313 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=55.12 //y=1.57 //x2=55.12 //y2=1.915
r972 (  216 316 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.12 //y=1.26 //x2=55.16 //y2=1.415
r973 (  215 315 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.12 //y=0.915 //x2=55.16 //y2=0.76
r974 (  215 216 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=55.12 //y=0.915 //x2=55.12 //y2=1.26
r975 (  212 318 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=54.87 //y=4.865 //x2=55.13 //y2=4.7
r976 (  211 310 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.51 //y=1.26 //x2=47.47 //y2=1.415
r977 (  210 309 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.51 //y=0.915 //x2=47.47 //y2=0.76
r978 (  210 211 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=47.51 //y=0.915 //x2=47.51 //y2=1.26
r979 (  208 306 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=47.135 //y=1.415 //x2=47.02 //y2=1.415
r980 (  207 310 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=47.355 //y=1.415 //x2=47.47 //y2=1.415
r981 (  206 305 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=47.135 //y=0.76 //x2=47.02 //y2=0.76
r982 (  205 309 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=47.355 //y=0.76 //x2=47.47 //y2=0.76
r983 (  205 206 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=47.355 //y=0.76 //x2=47.135 //y2=0.76
r984 (  202 308 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=47.17 //y=4.865 //x2=46.99 //y2=4.7
r985 (  200 306 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.98 //y=1.57 //x2=47.02 //y2=1.415
r986 (  200 303 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=46.98 //y=1.57 //x2=46.98 //y2=1.915
r987 (  199 306 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.98 //y=1.26 //x2=47.02 //y2=1.415
r988 (  198 305 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.98 //y=0.915 //x2=47.02 //y2=0.76
r989 (  198 199 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=46.98 //y=0.915 //x2=46.98 //y2=1.26
r990 (  195 308 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=46.73 //y=4.865 //x2=46.99 //y2=4.7
r991 (  194 296 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=82.47 //y=6.025 //x2=82.47 //y2=4.87
r992 (  193 288 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=82.03 //y=6.025 //x2=82.03 //y2=4.87
r993 (  192 281 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=79.15 //y=6.025 //x2=79.15 //y2=4.87
r994 (  191 269 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=78.71 //y=6.025 //x2=78.71 //y2=4.87
r995 (  190 262 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=66.5 //y=6.02 //x2=66.5 //y2=4.865
r996 (  189 255 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=66.06 //y=6.02 //x2=66.06 //y2=4.865
r997 (  188 243 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=62.87 //y=6.02 //x2=62.87 //y2=4.865
r998 (  187 233 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=62.43 //y=6.02 //x2=62.43 //y2=4.865
r999 (  186 219 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.31 //y=6.02 //x2=55.31 //y2=4.865
r1000 (  185 212 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=54.87 //y=6.02 //x2=54.87 //y2=4.865
r1001 (  184 202 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=47.17 //y=6.02 //x2=47.17 //y2=4.865
r1002 (  183 195 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=46.73 //y=6.02 //x2=46.73 //y2=4.865
r1003 (  182 293 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=82.21 //y=1.365 //x2=82.32 //y2=1.365
r1004 (  182 294 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=82.21 //y=1.365 //x2=82.1 //y2=1.365
r1005 (  181 274 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=78.88 //y=1.365 //x2=78.99 //y2=1.365
r1006 (  181 275 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=78.88 //y=1.365 //x2=78.77 //y2=1.365
r1007 (  180 252 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=65.825 //y=1.375 //x2=65.935 //y2=1.375
r1008 (  180 253 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=65.825 //y=1.375 //x2=65.715 //y2=1.375
r1009 (  179 238 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=62.6 //y=1.365 //x2=62.71 //y2=1.365
r1010 (  179 239 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=62.6 //y=1.365 //x2=62.49 //y2=1.365
r1011 (  178 224 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=55.385 //y=1.415 //x2=55.495 //y2=1.415
r1012 (  178 225 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=55.385 //y=1.415 //x2=55.275 //y2=1.415
r1013 (  177 207 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=47.245 //y=1.415 //x2=47.355 //y2=1.415
r1014 (  177 208 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=47.245 //y=1.415 //x2=47.135 //y2=1.415
r1015 (  171 352 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=82.14 //y=4.705 //x2=82.14 //y2=4.705
r1016 (  169 171 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=82.14 //y=4.44 //x2=82.14 //y2=4.705
r1017 (  166 347 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=82.14 //y=2.08 //x2=82.14 //y2=2.08
r1018 (  166 169 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=82.14 //y=2.08 //x2=82.14 //y2=4.44
r1019 (  163 341 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=78.44 //y=4.705 //x2=78.44 //y2=4.705
r1020 (  161 163 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=78.44 //y=4.44 //x2=78.44 //y2=4.705
r1021 (  159 161 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=78.44 //y=3.33 //x2=78.44 //y2=4.44
r1022 (  156 339 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=78.44 //y=2.08 //x2=78.44 //y2=2.08
r1023 (  156 159 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=78.44 //y=2.08 //x2=78.44 //y2=3.33
r1024 (  153 335 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=65.86 //y=4.7 //x2=65.86 //y2=4.7
r1025 (  151 153 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=65.86 //y=3.33 //x2=65.86 //y2=4.7
r1026 (  148 333 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=65.86 //y=2.08 //x2=65.86 //y2=2.08
r1027 (  148 151 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=65.86 //y=2.08 //x2=65.86 //y2=3.33
r1028 (  144 146 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=64.01 //y=5.115 //x2=64.01 //y2=3.33
r1029 (  143 146 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=64.01 //y=1.74 //x2=64.01 //y2=3.33
r1030 (  141 143 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=63.925 //y=1.655 //x2=64.01 //y2=1.74
r1031 (  141 142 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=63.925 //y=1.655 //x2=63.655 //y2=1.655
r1032 (  140 176 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.615 //y=5.2 //x2=63.53 //y2=5.2
r1033 (  139 144 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=63.925 //y=5.2 //x2=64.01 //y2=5.115
r1034 (  139 140 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=63.925 //y=5.2 //x2=63.615 //y2=5.2
r1035 (  135 142 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=63.57 //y=1.57 //x2=63.655 //y2=1.655
r1036 (  135 357 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=63.57 //y=1.57 //x2=63.57 //y2=1
r1037 (  129 176 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.53 //y=5.285 //x2=63.53 //y2=5.2
r1038 (  129 367 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=63.53 //y=5.285 //x2=63.53 //y2=5.725
r1039 (  127 176 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.445 //y=5.2 //x2=63.53 //y2=5.2
r1040 (  127 128 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=63.445 //y=5.2 //x2=62.735 //y2=5.2
r1041 (  121 128 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=62.65 //y=5.285 //x2=62.735 //y2=5.2
r1042 (  121 366 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=62.65 //y=5.285 //x2=62.65 //y2=5.725
r1043 (  119 327 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=62.53 //y=4.7 //x2=62.53 //y2=4.7
r1044 (  117 119 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=62.53 //y=3.33 //x2=62.53 //y2=4.7
r1045 (  114 322 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=62.53 //y=2.08 //x2=62.53 //y2=2.08
r1046 (  114 117 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=62.53 //y=2.08 //x2=62.53 //y2=3.33
r1047 (  110 112 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=60.68 //y=5.07 //x2=60.68 //y2=3.33
r1048 (  109 112 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=60.68 //y=1.75 //x2=60.68 //y2=3.33
r1049 (  107 109 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=60.595 //y=1.665 //x2=60.68 //y2=1.75
r1050 (  107 108 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=60.595 //y=1.665 //x2=60.28 //y2=1.665
r1051 (  103 108 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=60.195 //y=1.58 //x2=60.28 //y2=1.665
r1052 (  103 356 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=60.195 //y=1.58 //x2=60.195 //y2=1.01
r1053 (  102 175 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.985 //y=5.155 //x2=59.9 //y2=5.155
r1054 (  101 110 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=60.595 //y=5.155 //x2=60.68 //y2=5.07
r1055 (  101 102 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=60.595 //y=5.155 //x2=59.985 //y2=5.155
r1056 (  95 175 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.9 //y=5.24 //x2=59.9 //y2=5.155
r1057 (  95 365 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=59.9 //y=5.24 //x2=59.9 //y2=5.725
r1058 (  94 174 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.105 //y=5.155 //x2=59.02 //y2=5.155
r1059 (  93 175 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.815 //y=5.155 //x2=59.9 //y2=5.155
r1060 (  93 94 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=59.815 //y=5.155 //x2=59.105 //y2=5.155
r1061 (  87 174 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.02 //y=5.24 //x2=59.02 //y2=5.155
r1062 (  87 364 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=59.02 //y=5.24 //x2=59.02 //y2=5.725
r1063 (  85 174 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.935 //y=5.155 //x2=59.02 //y2=5.155
r1064 (  85 86 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=58.935 //y=5.155 //x2=58.225 //y2=5.155
r1065 (  79 86 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=58.14 //y=5.24 //x2=58.225 //y2=5.155
r1066 (  79 363 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=58.14 //y=5.24 //x2=58.14 //y2=5.725
r1067 (  77 318 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=55.13 //y=4.7 //x2=55.13 //y2=4.7
r1068 (  75 77 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=55.13 //y=3.33 //x2=55.13 //y2=4.7
r1069 (  72 312 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=55.13 //y=2.08 //x2=55.13 //y2=2.08
r1070 (  72 75 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=55.13 //y=2.08 //x2=55.13 //y2=3.33
r1071 (  68 70 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=51.06 //y=5.115 //x2=51.06 //y2=3.33
r1072 (  67 70 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=51.06 //y=1.74 //x2=51.06 //y2=3.33
r1073 (  65 67 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=50.975 //y=1.655 //x2=51.06 //y2=1.74
r1074 (  65 66 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=50.975 //y=1.655 //x2=50.705 //y2=1.655
r1075 (  64 173 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.665 //y=5.2 //x2=50.58 //y2=5.2
r1076 (  63 68 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=50.975 //y=5.2 //x2=51.06 //y2=5.115
r1077 (  63 64 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=50.975 //y=5.2 //x2=50.665 //y2=5.2
r1078 (  59 66 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=50.62 //y=1.57 //x2=50.705 //y2=1.655
r1079 (  59 355 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=50.62 //y=1.57 //x2=50.62 //y2=1
r1080 (  53 173 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.58 //y=5.285 //x2=50.58 //y2=5.2
r1081 (  53 362 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=50.58 //y=5.285 //x2=50.58 //y2=5.725
r1082 (  51 173 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.495 //y=5.2 //x2=50.58 //y2=5.2
r1083 (  51 52 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=50.495 //y=5.2 //x2=49.785 //y2=5.2
r1084 (  45 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=49.7 //y=5.285 //x2=49.785 //y2=5.2
r1085 (  45 361 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=49.7 //y=5.285 //x2=49.7 //y2=5.725
r1086 (  43 308 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=46.99 //y=4.7 //x2=46.99 //y2=4.7
r1087 (  41 43 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=46.99 //y=3.33 //x2=46.99 //y2=4.7
r1088 (  38 302 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=46.99 //y=2.08 //x2=46.99 //y2=2.08
r1089 (  38 41 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=46.99 //y=2.08 //x2=46.99 //y2=3.33
r1090 (  36 169 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=82.14 //y=4.44 //x2=82.14 //y2=4.44
r1091 (  34 159 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=78.44 //y=3.33 //x2=78.44 //y2=3.33
r1092 (  32 161 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=78.44 //y=4.44 //x2=78.44 //y2=4.44
r1093 (  30 151 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=65.86 //y=3.33 //x2=65.86 //y2=3.33
r1094 (  28 146 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=64.01 //y=3.33 //x2=64.01 //y2=3.33
r1095 (  26 117 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=62.53 //y=3.33 //x2=62.53 //y2=3.33
r1096 (  24 112 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=60.68 //y=3.33 //x2=60.68 //y2=3.33
r1097 (  22 75 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=55.13 //y=3.33 //x2=55.13 //y2=3.33
r1098 (  20 70 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=51.06 //y=3.33 //x2=51.06 //y2=3.33
r1099 (  18 41 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=46.99 //y=3.33 //x2=46.99 //y2=3.33
r1100 (  16 32 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=78.555 //y=4.44 //x2=78.44 //y2=4.44
r1101 (  15 36 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=82.025 //y=4.44 //x2=82.14 //y2=4.44
r1102 (  15 16 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=82.025 //y=4.44 //x2=78.555 //y2=4.44
r1103 (  14 30 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=65.975 //y=3.33 //x2=65.86 //y2=3.33
r1104 (  13 34 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=78.325 //y=3.33 //x2=78.44 //y2=3.33
r1105 (  13 14 ) resistor r=11.7844 //w=0.131 //l=12.35 //layer=m1 \
 //thickness=0.36 //x=78.325 //y=3.33 //x2=65.975 //y2=3.33
r1106 (  12 28 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=64.125 //y=3.33 //x2=64.01 //y2=3.33
r1107 (  11 30 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=65.745 //y=3.33 //x2=65.86 //y2=3.33
r1108 (  11 12 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 \
 //thickness=0.36 //x=65.745 //y=3.33 //x2=64.125 //y2=3.33
r1109 (  10 26 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=62.645 //y=3.33 //x2=62.53 //y2=3.33
r1110 (  9 28 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=63.895 //y=3.33 //x2=64.01 //y2=3.33
r1111 (  9 10 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=63.895 //y=3.33 //x2=62.645 //y2=3.33
r1112 (  8 24 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=60.795 //y=3.33 //x2=60.68 //y2=3.33
r1113 (  7 26 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=62.415 //y=3.33 //x2=62.53 //y2=3.33
r1114 (  7 8 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 \
 //thickness=0.36 //x=62.415 //y=3.33 //x2=60.795 //y2=3.33
r1115 (  6 22 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=55.245 //y=3.33 //x2=55.13 //y2=3.33
r1116 (  5 24 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=60.565 //y=3.33 //x2=60.68 //y2=3.33
r1117 (  5 6 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=60.565 //y=3.33 //x2=55.245 //y2=3.33
r1118 (  4 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=51.175 //y=3.33 //x2=51.06 //y2=3.33
r1119 (  3 22 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=55.015 //y=3.33 //x2=55.13 //y2=3.33
r1120 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=55.015 //y=3.33 //x2=51.175 //y2=3.33
r1121 (  2 18 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=47.105 //y=3.33 //x2=46.99 //y2=3.33
r1122 (  1 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=50.945 //y=3.33 //x2=51.06 //y2=3.33
r1123 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=50.945 //y=3.33 //x2=47.105 //y2=3.33
ends PM_TMRDFFRNQNX1\%noxref_17

subckt PM_TMRDFFRNQNX1\%noxref_18 ( 1 2 3 4 5 6 18 31 32 43 45 46 50 51 53 61 \
 65 69 72 73 74 75 76 77 78 79 80 84 85 86 91 93 96 97 98 99 100 105 107 109 \
 115 116 117 118 119 124 126 128 134 135 137 138 143 147 148 151 159 160 163 \
 171 173 174 )
c360 ( 174 0 ) capacitor c=0.0220235f //x=76.335 //y=5.02
c361 ( 173 0 ) capacitor c=0.0217503f //x=75.455 //y=5.02
c362 ( 171 0 ) capacitor c=0.00864721f //x=76.33 //y=0.905
c363 ( 163 0 ) capacitor c=0.0352016f //x=86.23 //y=4.705
c364 ( 160 0 ) capacitor c=0.0279733f //x=86.21 //y=1.915
c365 ( 159 0 ) capacitor c=0.0467621f //x=86.21 //y=2.08
c366 ( 151 0 ) capacitor c=0.03845f //x=79.59 //y=4.705
c367 ( 148 0 ) capacitor c=0.0300885f //x=79.55 //y=1.915
c368 ( 147 0 ) capacitor c=0.0520335f //x=79.55 //y=2.08
c369 ( 143 0 ) capacitor c=0.059212f //x=72.89 //y=4.7
c370 ( 138 0 ) capacitor c=0.0273931f //x=72.89 //y=1.915
c371 ( 137 0 ) capacitor c=0.0458323f //x=72.89 //y=2.08
c372 ( 135 0 ) capacitor c=0.0237734f //x=86.775 //y=1.255
c373 ( 134 0 ) capacitor c=0.0191782f //x=86.775 //y=0.905
c374 ( 128 0 ) capacitor c=0.0351663f //x=86.62 //y=1.405
c375 ( 126 0 ) capacitor c=0.0157803f //x=86.62 //y=0.75
c376 ( 124 0 ) capacitor c=0.0373879f //x=86.615 //y=4.795
c377 ( 119 0 ) capacitor c=0.0200628f //x=86.245 //y=1.56
c378 ( 118 0 ) capacitor c=0.0168575f //x=86.245 //y=1.255
c379 ( 117 0 ) capacitor c=0.0174993f //x=86.245 //y=0.905
c380 ( 116 0 ) capacitor c=0.0447087f //x=80.115 //y=1.25
c381 ( 115 0 ) capacitor c=0.019286f //x=80.115 //y=0.905
c382 ( 109 0 ) capacitor c=0.0187932f //x=79.96 //y=1.405
c383 ( 107 0 ) capacitor c=0.0157795f //x=79.96 //y=0.75
c384 ( 105 0 ) capacitor c=0.029531f //x=79.955 //y=4.795
c385 ( 100 0 ) capacitor c=0.0206178f //x=79.585 //y=1.56
c386 ( 99 0 ) capacitor c=0.016848f //x=79.585 //y=1.25
c387 ( 98 0 ) capacitor c=0.0174777f //x=79.585 //y=0.905
c388 ( 97 0 ) capacitor c=0.0432517f //x=73.41 //y=1.26
c389 ( 96 0 ) capacitor c=0.0200379f //x=73.41 //y=0.915
c390 ( 93 0 ) capacitor c=0.0158629f //x=73.255 //y=1.415
c391 ( 91 0 ) capacitor c=0.0157803f //x=73.255 //y=0.76
c392 ( 86 0 ) capacitor c=0.0218028f //x=72.88 //y=1.57
c393 ( 85 0 ) capacitor c=0.0207459f //x=72.88 //y=1.26
c394 ( 84 0 ) capacitor c=0.0194308f //x=72.88 //y=0.915
c395 ( 80 0 ) capacitor c=0.15325f //x=86.69 //y=6.025
c396 ( 79 0 ) capacitor c=0.110411f //x=86.25 //y=6.025
c397 ( 78 0 ) capacitor c=0.154236f //x=80.03 //y=6.025
c398 ( 77 0 ) capacitor c=0.110294f //x=79.59 //y=6.025
c399 ( 76 0 ) capacitor c=0.158794f //x=73.07 //y=6.02
c400 ( 75 0 ) capacitor c=0.110114f //x=72.63 //y=6.02
c401 ( 69 0 ) capacitor c=0.00501304f //x=86.23 //y=4.705
c402 ( 65 0 ) capacitor c=0.0024826f //x=76.48 //y=5.2
c403 ( 61 0 ) capacitor c=0.0899745f //x=86.21 //y=2.08
c404 ( 53 0 ) capacitor c=0.10473f //x=79.55 //y=2.08
c405 ( 51 0 ) capacitor c=0.00669947f //x=79.55 //y=4.54
c406 ( 50 0 ) capacitor c=0.106148f //x=76.96 //y=3.7
c407 ( 46 0 ) capacitor c=0.00468667f //x=76.605 //y=1.655
c408 ( 45 0 ) capacitor c=0.0131863f //x=76.875 //y=1.655
c409 ( 43 0 ) capacitor c=0.0141743f //x=76.875 //y=5.2
c410 ( 32 0 ) capacitor c=0.00265272f //x=75.685 //y=5.2
c411 ( 31 0 ) capacitor c=0.0150834f //x=76.395 //y=5.2
c412 ( 18 0 ) capacitor c=0.0870564f //x=72.89 //y=2.08
c413 ( 6 0 ) capacitor c=0.0101803f //x=79.665 //y=4.07
c414 ( 5 0 ) capacitor c=0.201218f //x=86.095 //y=4.07
c415 ( 4 0 ) capacitor c=0.00450722f //x=77.075 //y=3.7
c416 ( 3 0 ) capacitor c=0.0754105f //x=79.435 //y=3.7
c417 ( 2 0 ) capacitor c=0.00769527f //x=73.005 //y=3.7
c418 ( 1 0 ) capacitor c=0.0613342f //x=76.845 //y=3.7
r419 (  165 166 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=86.23 //y=4.795 //x2=86.23 //y2=4.87
r420 (  163 165 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=86.23 //y=4.705 //x2=86.23 //y2=4.795
r421 (  159 160 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=86.21 //y=2.08 //x2=86.21 //y2=1.915
r422 (  151 153 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=79.59 //y=4.705 //x2=79.59 //y2=4.795
r423 (  147 148 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=79.55 //y=2.08 //x2=79.55 //y2=1.915
r424 (  137 138 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=72.89 //y=2.08 //x2=72.89 //y2=1.915
r425 (  135 170 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=86.775 //y=1.255 //x2=86.775 //y2=1.367
r426 (  134 169 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=86.775 //y=0.905 //x2=86.735 //y2=0.75
r427 (  134 135 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=86.775 //y=0.905 //x2=86.775 //y2=1.255
r428 (  129 168 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=86.4 //y=1.405 //x2=86.285 //y2=1.405
r429 (  128 170 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=86.62 //y=1.405 //x2=86.775 //y2=1.367
r430 (  127 167 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=86.4 //y=0.75 //x2=86.285 //y2=0.75
r431 (  126 169 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=86.62 //y=0.75 //x2=86.735 //y2=0.75
r432 (  126 127 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=86.62 //y=0.75 //x2=86.4 //y2=0.75
r433 (  125 165 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=86.365 //y=4.795 //x2=86.23 //y2=4.795
r434 (  124 131 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=86.615 //y=4.795 //x2=86.69 //y2=4.87
r435 (  124 125 ) resistor r=128.191 //w=0.094 //l=0.25 //layer=ply \
 //thickness=0.18 //x=86.615 //y=4.795 //x2=86.365 //y2=4.795
r436 (  119 168 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=86.245 //y=1.56 //x2=86.285 //y2=1.405
r437 (  119 160 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=86.245 //y=1.56 //x2=86.245 //y2=1.915
r438 (  118 168 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=86.245 //y=1.255 //x2=86.285 //y2=1.405
r439 (  117 167 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=86.245 //y=0.905 //x2=86.285 //y2=0.75
r440 (  117 118 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=86.245 //y=0.905 //x2=86.245 //y2=1.255
r441 (  116 157 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.115 //y=1.25 //x2=80.075 //y2=1.405
r442 (  115 156 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.115 //y=0.905 //x2=80.075 //y2=0.75
r443 (  115 116 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=80.115 //y=0.905 //x2=80.115 //y2=1.25
r444 (  110 155 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=79.74 //y=1.405 //x2=79.625 //y2=1.405
r445 (  109 157 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=79.96 //y=1.405 //x2=80.075 //y2=1.405
r446 (  108 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=79.74 //y=0.75 //x2=79.625 //y2=0.75
r447 (  107 156 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=79.96 //y=0.75 //x2=80.075 //y2=0.75
r448 (  107 108 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=79.96 //y=0.75 //x2=79.74 //y2=0.75
r449 (  106 153 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=79.725 //y=4.795 //x2=79.59 //y2=4.795
r450 (  105 112 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=79.955 //y=4.795 //x2=80.03 //y2=4.87
r451 (  105 106 ) resistor r=117.936 //w=0.094 //l=0.23 //layer=ply \
 //thickness=0.18 //x=79.955 //y=4.795 //x2=79.725 //y2=4.795
r452 (  102 153 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=79.59 //y=4.87 //x2=79.59 //y2=4.795
r453 (  100 155 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.585 //y=1.56 //x2=79.625 //y2=1.405
r454 (  100 148 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=79.585 //y=1.56 //x2=79.585 //y2=1.915
r455 (  99 155 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.585 //y=1.25 //x2=79.625 //y2=1.405
r456 (  98 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.585 //y=0.905 //x2=79.625 //y2=0.75
r457 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=79.585 //y=0.905 //x2=79.585 //y2=1.25
r458 (  97 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=73.41 //y=1.26 //x2=73.37 //y2=1.415
r459 (  96 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=73.41 //y=0.915 //x2=73.37 //y2=0.76
r460 (  96 97 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=73.41 //y=0.915 //x2=73.41 //y2=1.26
r461 (  94 141 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.035 //y=1.415 //x2=72.92 //y2=1.415
r462 (  93 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.255 //y=1.415 //x2=73.37 //y2=1.415
r463 (  92 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.035 //y=0.76 //x2=72.92 //y2=0.76
r464 (  91 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=73.255 //y=0.76 //x2=73.37 //y2=0.76
r465 (  91 92 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=73.255 //y=0.76 //x2=73.035 //y2=0.76
r466 (  88 143 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=73.07 //y=4.865 //x2=72.89 //y2=4.7
r467 (  86 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.88 //y=1.57 //x2=72.92 //y2=1.415
r468 (  86 138 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=72.88 //y=1.57 //x2=72.88 //y2=1.915
r469 (  85 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.88 //y=1.26 //x2=72.92 //y2=1.415
r470 (  84 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.88 //y=0.915 //x2=72.92 //y2=0.76
r471 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=72.88 //y=0.915 //x2=72.88 //y2=1.26
r472 (  81 143 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=72.63 //y=4.865 //x2=72.89 //y2=4.7
r473 (  80 131 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=86.69 //y=6.025 //x2=86.69 //y2=4.87
r474 (  79 166 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=86.25 //y=6.025 //x2=86.25 //y2=4.87
r475 (  78 112 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=80.03 //y=6.025 //x2=80.03 //y2=4.87
r476 (  77 102 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=79.59 //y=6.025 //x2=79.59 //y2=4.87
r477 (  76 88 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=73.07 //y=6.02 //x2=73.07 //y2=4.865
r478 (  75 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=72.63 //y=6.02 //x2=72.63 //y2=4.865
r479 (  74 128 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=86.51 //y=1.405 //x2=86.62 //y2=1.405
r480 (  74 129 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=86.51 //y=1.405 //x2=86.4 //y2=1.405
r481 (  73 109 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=79.85 //y=1.405 //x2=79.96 //y2=1.405
r482 (  73 110 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=79.85 //y=1.405 //x2=79.74 //y2=1.405
r483 (  72 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=73.145 //y=1.415 //x2=73.255 //y2=1.415
r484 (  72 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=73.145 //y=1.415 //x2=73.035 //y2=1.415
r485 (  69 163 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=86.23 //y=4.705 //x2=86.23 //y2=4.705
r486 (  69 70 ) resistor r=10.3507 //w=0.207 //l=0.165 //layer=li \
 //thickness=0.1 //x=86.22 //y=4.705 //x2=86.22 //y2=4.54
r487 (  67 151 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=79.59 //y=4.705 //x2=79.59 //y2=4.705
r488 (  64 70 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=86.21 //y=4.07 //x2=86.21 //y2=4.54
r489 (  61 159 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=86.21 //y=2.08 //x2=86.21 //y2=2.08
r490 (  61 64 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=86.21 //y=2.08 //x2=86.21 //y2=4.07
r491 (  56 58 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=79.55 //y=3.7 //x2=79.55 //y2=4.07
r492 (  53 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=79.55 //y=2.08 //x2=79.55 //y2=2.08
r493 (  53 56 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=79.55 //y=2.08 //x2=79.55 //y2=3.7
r494 (  51 67 ) resistor r=11.2426 //w=0.191 //l=0.174714 //layer=li \
 //thickness=0.1 //x=79.55 //y=4.54 //x2=79.57 //y2=4.705
r495 (  51 58 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=79.55 //y=4.54 //x2=79.55 //y2=4.07
r496 (  48 50 ) resistor r=96.8556 //w=0.187 //l=1.415 //layer=li \
 //thickness=0.1 //x=76.96 //y=5.115 //x2=76.96 //y2=3.7
r497 (  47 50 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=76.96 //y=1.74 //x2=76.96 //y2=3.7
r498 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=76.875 //y=1.655 //x2=76.96 //y2=1.74
r499 (  45 46 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=76.875 //y=1.655 //x2=76.605 //y2=1.655
r500 (  44 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=76.565 //y=5.2 //x2=76.48 //y2=5.2
r501 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=76.875 //y=5.2 //x2=76.96 //y2=5.115
r502 (  43 44 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=76.875 //y=5.2 //x2=76.565 //y2=5.2
r503 (  39 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=76.52 //y=1.57 //x2=76.605 //y2=1.655
r504 (  39 171 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=76.52 //y=1.57 //x2=76.52 //y2=1
r505 (  33 65 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=76.48 //y=5.285 //x2=76.48 //y2=5.2
r506 (  33 174 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=76.48 //y=5.285 //x2=76.48 //y2=5.725
r507 (  31 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=76.395 //y=5.2 //x2=76.48 //y2=5.2
r508 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=76.395 //y=5.2 //x2=75.685 //y2=5.2
r509 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=75.6 //y=5.285 //x2=75.685 //y2=5.2
r510 (  25 173 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=75.6 //y=5.285 //x2=75.6 //y2=5.725
r511 (  23 143 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=72.89 //y=4.7 //x2=72.89 //y2=4.7
r512 (  21 23 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=72.89 //y=3.7 //x2=72.89 //y2=4.7
r513 (  18 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=72.89 //y=2.08 //x2=72.89 //y2=2.08
r514 (  18 21 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=72.89 //y=2.08 //x2=72.89 //y2=3.7
r515 (  16 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=86.21 //y=4.07 //x2=86.21 //y2=4.07
r516 (  14 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=79.55 //y=3.7 //x2=79.55 //y2=3.7
r517 (  12 58 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=79.55 //y=4.07 //x2=79.55 //y2=4.07
r518 (  10 50 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=76.96 //y=3.7 //x2=76.96 //y2=3.7
r519 (  8 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=72.89 //y=3.7 //x2=72.89 //y2=3.7
r520 (  6 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=79.665 //y=4.07 //x2=79.55 //y2=4.07
r521 (  5 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=86.095 //y=4.07 //x2=86.21 //y2=4.07
r522 (  5 6 ) resistor r=6.1355 //w=0.131 //l=6.43 //layer=m1 //thickness=0.36 \
 //x=86.095 //y=4.07 //x2=79.665 //y2=4.07
r523 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=77.075 //y=3.7 //x2=76.96 //y2=3.7
r524 (  3 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=79.435 //y=3.7 //x2=79.55 //y2=3.7
r525 (  3 4 ) resistor r=2.25191 //w=0.131 //l=2.36 //layer=m1 \
 //thickness=0.36 //x=79.435 //y=3.7 //x2=77.075 //y2=3.7
r526 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=73.005 //y=3.7 //x2=72.89 //y2=3.7
r527 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=76.845 //y=3.7 //x2=76.96 //y2=3.7
r528 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=76.845 //y=3.7 //x2=73.005 //y2=3.7
ends PM_TMRDFFRNQNX1\%noxref_18

subckt PM_TMRDFFRNQNX1\%noxref_19 ( 1 2 13 14 15 23 29 30 37 50 51 52 53 54 )
c91 ( 54 0 ) capacitor c=0.034295f //x=83.425 //y=5.025
c92 ( 53 0 ) capacitor c=0.0174957f //x=82.545 //y=5.025
c93 ( 51 0 ) capacitor c=0.0214849f //x=79.665 //y=5.025
c94 ( 50 0 ) capacitor c=0.0217161f //x=78.785 //y=5.025
c95 ( 49 0 ) capacitor c=0.00115294f //x=82.69 //y=6.91
c96 ( 37 0 ) capacitor c=0.0131238f //x=83.485 //y=6.91
c97 ( 30 0 ) capacitor c=0.00386507f //x=81.895 //y=6.91
c98 ( 29 0 ) capacitor c=0.00951687f //x=82.605 //y=6.91
c99 ( 23 0 ) capacitor c=0.0455351f //x=81.81 //y=5.21
c100 ( 15 0 ) capacitor c=0.00869404f //x=79.81 //y=5.295
c101 ( 14 0 ) capacitor c=0.00290434f //x=79.015 //y=5.21
c102 ( 13 0 ) capacitor c=0.0139202f //x=79.725 //y=5.21
c103 ( 2 0 ) capacitor c=0.0091252f //x=79.925 //y=5.21
c104 ( 1 0 ) capacitor c=0.0484159f //x=81.695 //y=5.21
r105 (  39 54 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=83.57 //y=6.825 //x2=83.57 //y2=6.74
r106 (  38 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.775 //y=6.91 //x2=82.69 //y2=6.91
r107 (  37 39 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=83.485 //y=6.91 //x2=83.57 //y2=6.825
r108 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=83.485 //y=6.91 //x2=82.775 //y2=6.91
r109 (  31 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.69 //y=6.825 //x2=82.69 //y2=6.91
r110 (  31 53 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.69 //y=6.825 //x2=82.69 //y2=6.74
r111 (  29 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.605 //y=6.91 //x2=82.69 //y2=6.91
r112 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=82.605 //y=6.91 //x2=81.895 //y2=6.91
r113 (  23 52 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=81.81 //y=5.21 //x2=81.81 //y2=6.06
r114 (  21 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=81.81 //y=6.825 //x2=81.895 //y2=6.91
r115 (  21 52 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.81 //y=6.825 //x2=81.81 //y2=6.74
r116 (  15 48 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=79.81 //y=5.295 //x2=79.81 //y2=5.17
r117 (  15 51 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=79.81 //y=5.295 //x2=79.81 //y2=6.06
r118 (  13 48 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=79.725 //y=5.21 //x2=79.81 //y2=5.17
r119 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=79.725 //y=5.21 //x2=79.015 //y2=5.21
r120 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=78.93 //y=5.295 //x2=79.015 //y2=5.21
r121 (  7 50 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=78.93 //y=5.295 //x2=78.93 //y2=5.72
r122 (  6 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=81.81 //y=5.21 //x2=81.81 //y2=5.21
r123 (  4 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=79.81 //y=5.21 //x2=79.81 //y2=5.21
r124 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=79.925 //y=5.21 //x2=79.81 //y2=5.21
r125 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=81.695 //y=5.21 //x2=81.81 //y2=5.21
r126 (  1 2 ) resistor r=1.68893 //w=0.131 //l=1.77 //layer=m1 \
 //thickness=0.36 //x=81.695 //y=5.21 //x2=79.925 //y2=5.21
ends PM_TMRDFFRNQNX1\%noxref_19

subckt PM_TMRDFFRNQNX1\%noxref_20 ( 1 2 3 4 5 6 18 31 32 43 45 46 50 52 61 67 \
 68 69 70 71 72 73 74 75 76 80 81 82 87 89 92 93 97 98 99 100 101 103 106 109 \
 110 111 112 113 114 115 116 120 122 125 126 127 128 133 134 139 151 158 160 \
 161 )
c493 ( 161 0 ) capacitor c=0.0220291f //x=24.535 //y=5.02
c494 ( 160 0 ) capacitor c=0.0217503f //x=23.655 //y=5.02
c495 ( 158 0 ) capacitor c=0.0084702f //x=24.53 //y=0.905
c496 ( 151 0 ) capacitor c=0.0583848f //x=85.1 //y=2.08
c497 ( 139 0 ) capacitor c=0.0587755f //x=21.09 //y=4.7
c498 ( 134 0 ) capacitor c=0.0273931f //x=21.09 //y=1.915
c499 ( 133 0 ) capacitor c=0.0456313f //x=21.09 //y=2.08
c500 ( 128 0 ) capacitor c=0.0316774f //x=85.805 //y=1.21
c501 ( 127 0 ) capacitor c=0.0187384f //x=85.805 //y=0.865
c502 ( 126 0 ) capacitor c=0.0590362f //x=85.445 //y=4.795
c503 ( 125 0 ) capacitor c=0.0296075f //x=85.735 //y=4.795
c504 ( 122 0 ) capacitor c=0.0157912f //x=85.65 //y=1.365
c505 ( 120 0 ) capacitor c=0.0149844f //x=85.65 //y=0.71
c506 ( 116 0 ) capacitor c=0.0302441f //x=85.275 //y=1.915
c507 ( 115 0 ) capacitor c=0.0234157f //x=85.275 //y=1.52
c508 ( 114 0 ) capacitor c=0.0234376f //x=85.275 //y=1.21
c509 ( 113 0 ) capacitor c=0.0199931f //x=85.275 //y=0.865
c510 ( 112 0 ) capacitor c=0.093437f //x=83.445 //y=1.915
c511 ( 111 0 ) capacitor c=0.0249466f //x=83.445 //y=1.56
c512 ( 110 0 ) capacitor c=0.0234397f //x=83.445 //y=1.25
c513 ( 109 0 ) capacitor c=0.0193195f //x=83.445 //y=0.905
c514 ( 106 0 ) capacitor c=0.0631944f //x=83.35 //y=4.87
c515 ( 103 0 ) capacitor c=0.0187941f //x=83.29 //y=1.405
c516 ( 101 0 ) capacitor c=0.0157803f //x=83.29 //y=0.75
c517 ( 100 0 ) capacitor c=0.010629f //x=82.985 //y=4.795
c518 ( 99 0 ) capacitor c=0.0194269f //x=83.275 //y=4.795
c519 ( 98 0 ) capacitor c=0.0365717f //x=82.915 //y=1.25
c520 ( 97 0 ) capacitor c=0.0175988f //x=82.915 //y=0.905
c521 ( 93 0 ) capacitor c=0.0432517f //x=21.61 //y=1.26
c522 ( 92 0 ) capacitor c=0.0200379f //x=21.61 //y=0.915
c523 ( 89 0 ) capacitor c=0.0148873f //x=21.455 //y=1.415
c524 ( 87 0 ) capacitor c=0.0157803f //x=21.455 //y=0.76
c525 ( 82 0 ) capacitor c=0.0218028f //x=21.08 //y=1.57
c526 ( 81 0 ) capacitor c=0.0207459f //x=21.08 //y=1.26
c527 ( 80 0 ) capacitor c=0.0194308f //x=21.08 //y=0.915
c528 ( 76 0 ) capacitor c=0.110622f //x=85.81 //y=6.025
c529 ( 75 0 ) capacitor c=0.154068f //x=85.37 //y=6.025
c530 ( 74 0 ) capacitor c=0.154291f //x=83.35 //y=6.025
c531 ( 73 0 ) capacitor c=0.110404f //x=82.91 //y=6.025
c532 ( 72 0 ) capacitor c=0.158794f //x=21.27 //y=6.02
c533 ( 71 0 ) capacitor c=0.110114f //x=20.83 //y=6.02
c534 ( 67 0 ) capacitor c=0.00211606f //x=24.68 //y=5.2
c535 ( 61 0 ) capacitor c=0.100881f //x=85.1 //y=2.08
c536 ( 52 0 ) capacitor c=0.105664f //x=83.62 //y=2.08
c537 ( 50 0 ) capacitor c=0.110129f //x=25.16 //y=2.96
c538 ( 46 0 ) capacitor c=0.00404073f //x=24.805 //y=1.655
c539 ( 45 0 ) capacitor c=0.0122201f //x=25.075 //y=1.655
c540 ( 43 0 ) capacitor c=0.0137995f //x=25.075 //y=5.2
c541 ( 32 0 ) capacitor c=0.00251635f //x=23.885 //y=5.2
c542 ( 31 0 ) capacitor c=0.0143649f //x=24.595 //y=5.2
c543 ( 18 0 ) capacitor c=0.0841327f //x=21.09 //y=2.08
c544 ( 6 0 ) capacitor c=0.0110448f //x=83.735 //y=2.08
c545 ( 5 0 ) capacitor c=0.0462526f //x=84.985 //y=2.08
c546 ( 4 0 ) capacitor c=0.00475948f //x=25.275 //y=2.96
c547 ( 3 0 ) capacitor c=1.08103f //x=83.505 //y=2.96
c548 ( 2 0 ) capacitor c=0.0130277f //x=21.205 //y=2.96
c549 ( 1 0 ) capacitor c=0.0776942f //x=25.045 //y=2.96
r550 (  133 134 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=21.09 //y=2.08 //x2=21.09 //y2=1.915
r551 (  128 157 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.805 //y=1.21 //x2=85.765 //y2=1.365
r552 (  127 156 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.805 //y=0.865 //x2=85.765 //y2=0.71
r553 (  127 128 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=85.805 //y=0.865 //x2=85.805 //y2=1.21
r554 (  125 129 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=85.735 //y=4.795 //x2=85.81 //y2=4.87
r555 (  125 126 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=85.735 //y=4.795 //x2=85.445 //y2=4.795
r556 (  123 155 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=85.43 //y=1.365 //x2=85.315 //y2=1.365
r557 (  122 157 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=85.65 //y=1.365 //x2=85.765 //y2=1.365
r558 (  121 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=85.43 //y=0.71 //x2=85.315 //y2=0.71
r559 (  120 156 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=85.65 //y=0.71 //x2=85.765 //y2=0.71
r560 (  120 121 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=85.65 //y=0.71 //x2=85.43 //y2=0.71
r561 (  117 126 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=85.37 //y=4.87 //x2=85.445 //y2=4.795
r562 (  117 153 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=85.37 //y=4.87 //x2=85.1 //y2=4.705
r563 (  116 151 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=85.275 //y=1.915 //x2=85.1 //y2=2.08
r564 (  115 155 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.275 //y=1.52 //x2=85.315 //y2=1.365
r565 (  115 116 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=85.275 //y=1.52 //x2=85.275 //y2=1.915
r566 (  114 155 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.275 //y=1.21 //x2=85.315 //y2=1.365
r567 (  113 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=85.275 //y=0.865 //x2=85.315 //y2=0.71
r568 (  113 114 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=85.275 //y=0.865 //x2=85.275 //y2=1.21
r569 (  112 147 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=83.445 //y=1.915 //x2=83.62 //y2=2.08
r570 (  111 145 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=83.445 //y=1.56 //x2=83.405 //y2=1.405
r571 (  111 112 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=83.445 //y=1.56 //x2=83.445 //y2=1.915
r572 (  110 145 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=83.445 //y=1.25 //x2=83.405 //y2=1.405
r573 (  109 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=83.445 //y=0.905 //x2=83.405 //y2=0.75
r574 (  109 110 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=83.445 //y=0.905 //x2=83.445 //y2=1.25
r575 (  106 149 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=83.35 //y=4.87 //x2=83.62 //y2=4.705
r576 (  104 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=83.07 //y=1.405 //x2=82.955 //y2=1.405
r577 (  103 145 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=83.29 //y=1.405 //x2=83.405 //y2=1.405
r578 (  102 142 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=83.07 //y=0.75 //x2=82.955 //y2=0.75
r579 (  101 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=83.29 //y=0.75 //x2=83.405 //y2=0.75
r580 (  101 102 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=83.29 //y=0.75 //x2=83.07 //y2=0.75
r581 (  99 106 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=83.275 //y=4.795 //x2=83.35 //y2=4.87
r582 (  99 100 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=83.275 //y=4.795 //x2=82.985 //y2=4.795
r583 (  98 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=82.915 //y=1.25 //x2=82.955 //y2=1.405
r584 (  97 142 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=82.915 //y=0.905 //x2=82.955 //y2=0.75
r585 (  97 98 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=82.915 //y=0.905 //x2=82.915 //y2=1.25
r586 (  94 100 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=82.91 //y=4.87 //x2=82.985 //y2=4.795
r587 (  93 141 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.61 //y=1.26 //x2=21.57 //y2=1.415
r588 (  92 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.61 //y=0.915 //x2=21.57 //y2=0.76
r589 (  92 93 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=21.61 //y=0.915 //x2=21.61 //y2=1.26
r590 (  90 137 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.235 //y=1.415 //x2=21.12 //y2=1.415
r591 (  89 141 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.455 //y=1.415 //x2=21.57 //y2=1.415
r592 (  88 136 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.235 //y=0.76 //x2=21.12 //y2=0.76
r593 (  87 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.455 //y=0.76 //x2=21.57 //y2=0.76
r594 (  87 88 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=21.455 //y=0.76 //x2=21.235 //y2=0.76
r595 (  84 139 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=21.27 //y=4.865 //x2=21.09 //y2=4.7
r596 (  82 137 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.08 //y=1.57 //x2=21.12 //y2=1.415
r597 (  82 134 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=21.08 //y=1.57 //x2=21.08 //y2=1.915
r598 (  81 137 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.08 //y=1.26 //x2=21.12 //y2=1.415
r599 (  80 136 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.08 //y=0.915 //x2=21.12 //y2=0.76
r600 (  80 81 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=21.08 //y=0.915 //x2=21.08 //y2=1.26
r601 (  77 139 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=20.83 //y=4.865 //x2=21.09 //y2=4.7
r602 (  76 129 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=85.81 //y=6.025 //x2=85.81 //y2=4.87
r603 (  75 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=85.37 //y=6.025 //x2=85.37 //y2=4.87
r604 (  74 106 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=83.35 //y=6.025 //x2=83.35 //y2=4.87
r605 (  73 94 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=82.91 //y=6.025 //x2=82.91 //y2=4.87
r606 (  72 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.27 //y=6.02 //x2=21.27 //y2=4.865
r607 (  71 77 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.83 //y=6.02 //x2=20.83 //y2=4.865
r608 (  70 122 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=85.54 //y=1.365 //x2=85.65 //y2=1.365
r609 (  70 123 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=85.54 //y=1.365 //x2=85.43 //y2=1.365
r610 (  69 103 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=83.18 //y=1.405 //x2=83.29 //y2=1.405
r611 (  69 104 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=83.18 //y=1.405 //x2=83.07 //y2=1.405
r612 (  68 89 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=21.345 //y=1.415 //x2=21.455 //y2=1.415
r613 (  68 90 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=21.345 //y=1.415 //x2=21.235 //y2=1.415
r614 (  65 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=85.1 //y=4.705 //x2=85.1 //y2=4.705
r615 (  61 151 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=85.1 //y=2.08 //x2=85.1 //y2=2.08
r616 (  61 65 ) resistor r=179.679 //w=0.187 //l=2.625 //layer=li \
 //thickness=0.1 //x=85.1 //y=2.08 //x2=85.1 //y2=4.705
r617 (  58 149 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=83.62 //y=4.705 //x2=83.62 //y2=4.705
r618 (  56 58 ) resistor r=119.444 //w=0.187 //l=1.745 //layer=li \
 //thickness=0.1 //x=83.62 //y=2.96 //x2=83.62 //y2=4.705
r619 (  52 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=83.62 //y=2.08 //x2=83.62 //y2=2.08
r620 (  52 56 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=83.62 //y=2.08 //x2=83.62 //y2=2.96
r621 (  48 50 ) resistor r=147.508 //w=0.187 //l=2.155 //layer=li \
 //thickness=0.1 //x=25.16 //y=5.115 //x2=25.16 //y2=2.96
r622 (  47 50 ) resistor r=83.508 //w=0.187 //l=1.22 //layer=li \
 //thickness=0.1 //x=25.16 //y=1.74 //x2=25.16 //y2=2.96
r623 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.075 //y=1.655 //x2=25.16 //y2=1.74
r624 (  45 46 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=25.075 //y=1.655 //x2=24.805 //y2=1.655
r625 (  44 67 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.765 //y=5.2 //x2=24.68 //y2=5.2
r626 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.075 //y=5.2 //x2=25.16 //y2=5.115
r627 (  43 44 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=25.075 //y=5.2 //x2=24.765 //y2=5.2
r628 (  39 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=24.72 //y=1.57 //x2=24.805 //y2=1.655
r629 (  39 158 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.72 //y=1.57 //x2=24.72 //y2=1
r630 (  33 67 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.68 //y=5.285 //x2=24.68 //y2=5.2
r631 (  33 161 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=24.68 //y=5.285 //x2=24.68 //y2=5.725
r632 (  31 67 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.595 //y=5.2 //x2=24.68 //y2=5.2
r633 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=24.595 //y=5.2 //x2=23.885 //y2=5.2
r634 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.8 //y=5.285 //x2=23.885 //y2=5.2
r635 (  25 160 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=23.8 //y=5.285 //x2=23.8 //y2=5.725
r636 (  23 139 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.09 //y=4.7 //x2=21.09 //y2=4.7
r637 (  21 23 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=21.09 //y=2.96 //x2=21.09 //y2=4.7
r638 (  18 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.09 //y=2.08 //x2=21.09 //y2=2.08
r639 (  18 21 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=21.09 //y=2.08 //x2=21.09 //y2=2.96
r640 (  16 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=85.1 //y=2.08 //x2=85.1 //y2=2.08
r641 (  14 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=83.62 //y=2.96 //x2=83.62 //y2=2.96
r642 (  12 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=83.62 //y=2.08 //x2=83.62 //y2=2.08
r643 (  10 50 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=25.16 //y=2.96 //x2=25.16 //y2=2.96
r644 (  8 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.09 //y=2.96 //x2=21.09 //y2=2.96
r645 (  6 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=83.735 //y=2.08 //x2=83.62 //y2=2.08
r646 (  5 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=84.985 //y=2.08 //x2=85.1 //y2=2.08
r647 (  5 6 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=84.985 //y=2.08 //x2=83.735 //y2=2.08
r648 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=25.275 //y=2.96 //x2=25.16 //y2=2.96
r649 (  3 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=83.505 //y=2.96 //x2=83.62 //y2=2.96
r650 (  3 4 ) resistor r=55.563 //w=0.131 //l=58.23 //layer=m1 \
 //thickness=0.36 //x=83.505 //y=2.96 //x2=25.275 //y2=2.96
r651 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.205 //y=2.96 //x2=21.09 //y2=2.96
r652 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=25.045 //y=2.96 //x2=25.16 //y2=2.96
r653 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=25.045 //y=2.96 //x2=21.205 //y2=2.96
ends PM_TMRDFFRNQNX1\%noxref_20

subckt PM_TMRDFFRNQNX1\%noxref_21 ( 1 2 13 14 15 21 27 28 35 46 47 48 49 50 )
c89 ( 50 0 ) capacitor c=0.0308836f //x=86.765 //y=5.025
c90 ( 49 0 ) capacitor c=0.0173945f //x=85.885 //y=5.025
c91 ( 47 0 ) capacitor c=0.0169278f //x=82.985 //y=5.025
c92 ( 46 0 ) capacitor c=0.0166762f //x=82.105 //y=5.025
c93 ( 45 0 ) capacitor c=0.00115294f //x=86.03 //y=6.91
c94 ( 35 0 ) capacitor c=0.0132983f //x=86.825 //y=6.91
c95 ( 28 0 ) capacitor c=0.00388794f //x=85.235 //y=6.91
c96 ( 27 0 ) capacitor c=0.00985708f //x=85.945 //y=6.91
c97 ( 21 0 ) capacitor c=0.0442221f //x=85.15 //y=5.21
c98 ( 15 0 ) capacitor c=0.0105083f //x=83.13 //y=5.295
c99 ( 14 0 ) capacitor c=0.00227812f //x=82.335 //y=5.21
c100 ( 13 0 ) capacitor c=0.0174384f //x=83.045 //y=5.21
c101 ( 2 0 ) capacitor c=0.00682032f //x=83.245 //y=5.21
c102 ( 1 0 ) capacitor c=0.0574911f //x=85.035 //y=5.21
r103 (  37 50 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=86.91 //y=6.825 //x2=86.91 //y2=6.74
r104 (  36 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=86.115 //y=6.91 //x2=86.03 //y2=6.91
r105 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=86.825 //y=6.91 //x2=86.91 //y2=6.825
r106 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=86.825 //y=6.91 //x2=86.115 //y2=6.91
r107 (  29 45 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=86.03 //y=6.825 //x2=86.03 //y2=6.91
r108 (  29 49 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=86.03 //y=6.825 //x2=86.03 //y2=6.74
r109 (  27 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=85.945 //y=6.91 //x2=86.03 //y2=6.91
r110 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=85.945 //y=6.91 //x2=85.235 //y2=6.91
r111 (  21 48 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=85.15 //y=5.21 //x2=85.15 //y2=6.06
r112 (  19 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=85.15 //y=6.825 //x2=85.235 //y2=6.91
r113 (  19 48 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=85.15 //y=6.825 //x2=85.15 //y2=6.74
r114 (  15 44 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=83.13 //y=5.295 //x2=83.13 //y2=5.17
r115 (  15 47 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=83.13 //y=5.295 //x2=83.13 //y2=6.06
r116 (  13 44 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=83.045 //y=5.21 //x2=83.13 //y2=5.17
r117 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=83.045 //y=5.21 //x2=82.335 //y2=5.21
r118 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=82.25 //y=5.295 //x2=82.335 //y2=5.21
r119 (  7 46 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=82.25 //y=5.295 //x2=82.25 //y2=5.72
r120 (  6 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=85.15 //y=5.21 //x2=85.15 //y2=5.21
r121 (  4 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=83.13 //y=5.21 //x2=83.13 //y2=5.21
r122 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=83.245 //y=5.21 //x2=83.13 //y2=5.21
r123 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=85.035 //y=5.21 //x2=85.15 //y2=5.21
r124 (  1 2 ) resistor r=1.70802 //w=0.131 //l=1.79 //layer=m1 \
 //thickness=0.36 //x=85.035 //y=5.21 //x2=83.245 //y2=5.21
ends PM_TMRDFFRNQNX1\%noxref_21

subckt PM_TMRDFFRNQNX1\%QN ( 1 2 3 4 11 12 13 14 15 16 17 18 31 32 45 47 48 63 \
 64 65 66 70 71 )
c169 ( 71 0 ) capacitor c=0.0167617f //x=86.325 //y=5.025
c170 ( 70 0 ) capacitor c=0.0164812f //x=85.445 //y=5.025
c171 ( 66 0 ) capacitor c=0.0108176f //x=86.32 //y=0.905
c172 ( 65 0 ) capacitor c=0.0131637f //x=82.99 //y=0.905
c173 ( 64 0 ) capacitor c=0.0131367f //x=79.66 //y=0.905
c174 ( 63 0 ) capacitor c=0.00421476f //x=86.47 //y=5.21
c175 ( 48 0 ) capacitor c=0.00775877f //x=86.595 //y=1.645
c176 ( 47 0 ) capacitor c=0.0165978f //x=86.865 //y=1.645
c177 ( 45 0 ) capacitor c=0.0160142f //x=86.865 //y=5.21
c178 ( 32 0 ) capacitor c=0.0029383f //x=85.675 //y=5.21
c179 ( 31 0 ) capacitor c=0.0155464f //x=86.385 //y=5.21
c180 ( 11 0 ) capacitor c=0.133166f //x=86.95 //y=2.22
c181 ( 4 0 ) capacitor c=0.00511584f //x=83.295 //y=1.18
c182 ( 3 0 ) capacitor c=0.0702096f //x=86.395 //y=1.18
c183 ( 2 0 ) capacitor c=0.0150174f //x=79.965 //y=1.18
c184 ( 1 0 ) capacitor c=0.0604206f //x=83.065 //y=1.18
r185 (  62 64 ) resistor r=13.3953 //w=0.172 //l=0.18 //layer=li \
 //thickness=0.1 //x=79.847 //y=1.18 //x2=79.847 //y2=1
r186 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=86.865 //y=1.645 //x2=86.95 //y2=1.73
r187 (  47 48 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=86.865 //y=1.645 //x2=86.595 //y2=1.645
r188 (  46 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=86.555 //y=5.21 //x2=86.47 //y2=5.21
r189 (  45 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=86.865 //y=5.21 //x2=86.95 //y2=5.125
r190 (  45 46 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=86.865 //y=5.21 //x2=86.555 //y2=5.21
r191 (  44 66 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=86.51 //y=1.18 //x2=86.51 //y2=1
r192 (  39 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=86.51 //y=1.56 //x2=86.595 //y2=1.645
r193 (  39 44 ) resistor r=26.0107 //w=0.187 //l=0.38 //layer=li \
 //thickness=0.1 //x=86.51 //y=1.56 //x2=86.51 //y2=1.18
r194 (  33 63 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=86.47 //y=5.295 //x2=86.47 //y2=5.21
r195 (  33 71 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=86.47 //y=5.295 //x2=86.47 //y2=5.72
r196 (  31 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=86.385 //y=5.21 //x2=86.47 //y2=5.21
r197 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=86.385 //y=5.21 //x2=85.675 //y2=5.21
r198 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=85.59 //y=5.295 //x2=85.675 //y2=5.21
r199 (  25 70 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=85.59 //y=5.295 //x2=85.59 //y2=5.72
r200 (  23 65 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=83.18 //y=1.18 //x2=83.18 //y2=1
r201 (  18 50 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=86.95 //y=4.81 //x2=86.95 //y2=5.125
r202 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=86.95 //y=4.44 //x2=86.95 //y2=4.81
r203 (  16 17 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=86.95 //y=4.07 //x2=86.95 //y2=4.44
r204 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=86.95 //y=3.7 //x2=86.95 //y2=4.07
r205 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=86.95 //y=3.33 //x2=86.95 //y2=3.7
r206 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=86.95 //y=2.96 //x2=86.95 //y2=3.33
r207 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=86.95 //y=2.59 //x2=86.95 //y2=2.96
r208 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=86.95 //y=2.22 //x2=86.95 //y2=2.59
r209 (  11 49 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=86.95 //y=2.22 //x2=86.95 //y2=1.73
r210 (  10 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=86.51 //y=1.18 //x2=86.51 //y2=1.18
r211 (  8 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=83.18 //y=1.18 //x2=83.18 //y2=1.18
r212 (  6 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=79.85 //y=1.18 //x2=79.85 //y2=1.18
r213 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=83.295 //y=1.18 //x2=83.18 //y2=1.18
r214 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=86.395 //y=1.18 //x2=86.51 //y2=1.18
r215 (  3 4 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=86.395 //y=1.18 //x2=83.295 //y2=1.18
r216 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=79.965 //y=1.18 //x2=79.85 //y2=1.18
r217 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=83.065 //y=1.18 //x2=83.18 //y2=1.18
r218 (  1 2 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=83.065 //y=1.18 //x2=79.965 //y2=1.18
ends PM_TMRDFFRNQNX1\%QN

subckt PM_TMRDFFRNQNX1\%noxref_23 ( 1 5 9 13 17 35 )
c46 ( 35 0 ) capacitor c=0.0703709f //x=0.455 //y=0.375
c47 ( 17 0 ) capacitor c=0.0221229f //x=2.445 //y=1.59
c48 ( 13 0 ) capacitor c=0.0156939f //x=2.445 //y=0.54
c49 ( 9 0 ) capacitor c=0.00678203f //x=1.56 //y=0.625
c50 ( 5 0 ) capacitor c=0.0206412f //x=1.475 //y=1.59
c51 ( 1 0 ) capacitor c=0.0109947f //x=0.59 //y=1.505
r52 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=1.59 //x2=1.56 //y2=1.63
r53 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=1.59 //x2=2.045 //y2=1.59
r54 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=1.59 //x2=2.53 //y2=1.59
r55 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=1.59 //x2=2.045 //y2=1.59
r56 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=0.54 //x2=1.56 //y2=0.5
r57 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=0.54 //x2=2.045 //y2=0.54
r58 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=0.54 //x2=2.53 //y2=0.54
r59 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=0.54 //x2=2.045 //y2=0.54
r60 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=1.63
r61 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=0.89
r62 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.5
r63 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.89
r64 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.675 //y=1.59 //x2=0.59 //y2=1.63
r65 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.675 //y=1.59 //x2=1.075 //y2=1.59
r66 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.475 //y=1.59 //x2=1.56 //y2=1.63
r67 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.475 //y=1.59 //x2=1.075 //y2=1.59
r68 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.59 //y=1.505 //x2=0.59 //y2=1.63
r69 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.59 //y=1.505 //x2=0.59 //y2=0.89
ends PM_TMRDFFRNQNX1\%noxref_23

subckt PM_TMRDFFRNQNX1\%noxref_24 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.043074f //x=2.965 //y=0.375
c53 ( 28 0 ) capacitor c=0.00465142f //x=1.86 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=3.1 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=4.07 //y=0.625
c56 ( 11 0 ) capacitor c=0.0149771f //x=3.985 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=3.1 //y=0.625
c58 ( 1 0 ) capacitor c=0.0251532f //x=3.015 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.185 //y=0.54 //x2=3.1 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.185 //y=0.54 //x2=3.585 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.985 //y=0.54 //x2=4.07 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.985 //y=0.54 //x2=3.585 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.135 //y=0.995 //x2=2.05 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=3.1 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=2.135 //y2=0.995
ends PM_TMRDFFRNQNX1\%noxref_24

subckt PM_TMRDFFRNQNX1\%noxref_25 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0686255f //x=5.265 //y=0.375
c53 ( 17 0 ) capacitor c=0.020294f //x=7.255 //y=1.59
c54 ( 13 0 ) capacitor c=0.0155578f //x=7.255 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=6.37 //y=0.625
c56 ( 5 0 ) capacitor c=0.0183576f //x=6.285 //y=1.59
c57 ( 1 0 ) capacitor c=0.00791969f //x=5.4 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.455 //y=1.59 //x2=6.37 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.455 //y=1.59 //x2=6.855 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.255 //y=1.59 //x2=7.34 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.255 //y=1.59 //x2=6.855 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.455 //y=0.54 //x2=6.37 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.455 //y=0.54 //x2=6.855 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.255 //y=0.54 //x2=7.34 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.255 //y=0.54 //x2=6.855 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=6.37 //y=1.505 //x2=6.37 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.37 //y=1.505 //x2=6.37 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.37 //y=0.625 //x2=6.37 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.37 //y=0.625 //x2=6.37 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.485 //y=1.59 //x2=5.4 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.485 //y=1.59 //x2=5.885 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.285 //y=1.59 //x2=6.37 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.285 //y=1.59 //x2=5.885 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=5.4 //y=1.505 //x2=5.4 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=5.4 //y=1.505 //x2=5.4 //y2=0.89
ends PM_TMRDFFRNQNX1\%noxref_25

subckt PM_TMRDFFRNQNX1\%noxref_26 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.041714f //x=7.775 //y=0.375
c54 ( 28 0 ) capacitor c=0.00462171f //x=6.67 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=7.91 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=8.88 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=8.795 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=7.91 //y=0.625
c59 ( 1 0 ) capacitor c=0.0227139f //x=7.825 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=8.88 //y=0.625 //x2=8.88 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=8.88 //y=0.625 //x2=8.88 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.995 //y=0.54 //x2=7.91 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.995 //y=0.54 //x2=8.395 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.795 //y=0.54 //x2=8.88 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.795 //y=0.54 //x2=8.395 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.91 //y=1.08 //x2=7.91 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=7.91 //y=1.08 //x2=7.91 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.91 //x2=7.91 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.91 //x2=7.91 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.625 //x2=7.91 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.625 //x2=7.91 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.945 //y=0.995 //x2=6.86 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.825 //y=0.995 //x2=7.91 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=7.825 //y=0.995 //x2=6.945 //y2=0.995
ends PM_TMRDFFRNQNX1\%noxref_26

subckt PM_TMRDFFRNQNX1\%noxref_27 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632682f //x=10.18 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=12.255 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=12.17 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=11.285 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=11.285 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=11.2 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=10.315 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=12.255 //y=0.615 //x2=12.255 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=12.255 //y=0.615 //x2=12.255 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.37 //y=0.53 //x2=11.285 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.37 //y=0.53 //x2=11.77 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.17 //y=0.53 //x2=12.255 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.17 //y=0.53 //x2=11.77 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=11.285 //y=1.495 //x2=11.285 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=11.285 //y=1.495 //x2=11.285 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=11.285 //y=0.615 //x2=11.285 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=11.285 //y=0.615 //x2=11.285 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.4 //y=1.58 //x2=10.315 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.4 //y=1.58 //x2=10.8 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.2 //y=1.58 //x2=11.285 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.2 //y=1.58 //x2=10.8 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=10.315 //y=1.495 //x2=10.315 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=10.315 //y=1.495 //x2=10.315 //y2=0.88
ends PM_TMRDFFRNQNX1\%noxref_27

subckt PM_TMRDFFRNQNX1\%noxref_28 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=13.405 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=15.395 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=15.395 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=14.51 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=14.425 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=13.54 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.595 //y=1.59 //x2=14.51 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.595 //y=1.59 //x2=14.995 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.395 //y=1.59 //x2=15.48 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.395 //y=1.59 //x2=14.995 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.595 //y=0.54 //x2=14.51 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.595 //y=0.54 //x2=14.995 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.395 //y=0.54 //x2=15.48 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.395 //y=0.54 //x2=14.995 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=14.51 //y=1.505 //x2=14.51 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=14.51 //y=1.505 //x2=14.51 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=14.51 //y=0.625 //x2=14.51 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=14.51 //y=0.625 //x2=14.51 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.625 //y=1.59 //x2=13.54 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.625 //y=1.59 //x2=14.025 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.425 //y=1.59 //x2=14.51 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.425 //y=1.59 //x2=14.025 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=13.54 //y=1.505 //x2=13.54 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=13.54 //y=1.505 //x2=13.54 //y2=0.89
ends PM_TMRDFFRNQNX1\%noxref_28

subckt PM_TMRDFFRNQNX1\%noxref_29 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0413887f //x=15.915 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=14.81 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=16.05 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=17.02 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=16.935 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=16.05 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=15.965 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=17.02 //y=0.625 //x2=17.02 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=17.02 //y=0.625 //x2=17.02 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.135 //y=0.54 //x2=16.05 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.135 //y=0.54 //x2=16.535 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.935 //y=0.54 //x2=17.02 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.935 //y=0.54 //x2=16.535 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=16.05 //y=1.08 //x2=16.05 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=16.05 //y=1.08 //x2=16.05 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=16.05 //y=0.91 //x2=16.05 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=16.05 //y=0.91 //x2=16.05 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=16.05 //y=0.625 //x2=16.05 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=16.05 //y=0.625 //x2=16.05 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.085 //y=0.995 //x2=15 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=15.965 //y=0.995 //x2=16.05 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=15.965 //y=0.995 //x2=15.085 //y2=0.995
ends PM_TMRDFFRNQNX1\%noxref_29

subckt PM_TMRDFFRNQNX1\%noxref_30 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=18.215 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=20.205 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=20.205 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=19.32 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=19.235 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=18.35 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.405 //y=1.59 //x2=19.32 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.405 //y=1.59 //x2=19.805 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.205 //y=1.59 //x2=20.29 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.205 //y=1.59 //x2=19.805 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.405 //y=0.54 //x2=19.32 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.405 //y=0.54 //x2=19.805 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.205 //y=0.54 //x2=20.29 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.205 //y=0.54 //x2=19.805 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=19.32 //y=1.505 //x2=19.32 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=19.32 //y=1.505 //x2=19.32 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=19.32 //y=0.625 //x2=19.32 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=19.32 //y=0.625 //x2=19.32 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.435 //y=1.59 //x2=18.35 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.435 //y=1.59 //x2=18.835 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.235 //y=1.59 //x2=19.32 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.235 //y=1.59 //x2=18.835 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=18.35 //y=1.505 //x2=18.35 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=18.35 //y=1.505 //x2=18.35 //y2=0.89
ends PM_TMRDFFRNQNX1\%noxref_30

subckt PM_TMRDFFRNQNX1\%noxref_31 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=20.725 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=19.62 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=20.86 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=21.83 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=21.745 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=20.86 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=20.775 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=21.83 //y=0.625 //x2=21.83 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=21.83 //y=0.625 //x2=21.83 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.945 //y=0.54 //x2=20.86 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.945 //y=0.54 //x2=21.345 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.745 //y=0.54 //x2=21.83 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.745 //y=0.54 //x2=21.345 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.86 //y=1.08 //x2=20.86 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=20.86 //y=1.08 //x2=20.86 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.86 //y=0.91 //x2=20.86 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=20.86 //y=0.91 //x2=20.86 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=20.86 //y=0.625 //x2=20.86 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=20.86 //y=0.625 //x2=20.86 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.895 //y=0.995 //x2=19.81 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.775 //y=0.995 //x2=20.86 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=20.775 //y=0.995 //x2=19.895 //y2=0.995
ends PM_TMRDFFRNQNX1\%noxref_31

subckt PM_TMRDFFRNQNX1\%noxref_32 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632682f //x=23.13 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=25.205 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=25.12 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=24.235 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=24.235 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=24.15 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=23.265 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=25.205 //y=0.615 //x2=25.205 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=25.205 //y=0.615 //x2=25.205 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=24.32 //y=0.53 //x2=24.235 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=24.32 //y=0.53 //x2=24.72 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.12 //y=0.53 //x2=25.205 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.12 //y=0.53 //x2=24.72 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=24.235 //y=1.495 //x2=24.235 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=24.235 //y=1.495 //x2=24.235 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=24.235 //y=0.615 //x2=24.235 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=24.235 //y=0.615 //x2=24.235 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.35 //y=1.58 //x2=23.265 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.35 //y=1.58 //x2=23.75 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=24.15 //y=1.58 //x2=24.235 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=24.15 //y=1.58 //x2=23.75 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=23.265 //y=1.495 //x2=23.265 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=23.265 //y=1.495 //x2=23.265 //y2=0.88
ends PM_TMRDFFRNQNX1\%noxref_32

subckt PM_TMRDFFRNQNX1\%noxref_33 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=26.355 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=28.345 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=28.345 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=27.46 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=27.375 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=26.49 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=27.545 //y=1.59 //x2=27.46 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=27.545 //y=1.59 //x2=27.945 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.345 //y=1.59 //x2=28.43 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=28.345 //y=1.59 //x2=27.945 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=27.545 //y=0.54 //x2=27.46 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=27.545 //y=0.54 //x2=27.945 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.345 //y=0.54 //x2=28.43 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=28.345 //y=0.54 //x2=27.945 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=27.46 //y=1.505 //x2=27.46 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=27.46 //y=1.505 //x2=27.46 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=27.46 //y=0.625 //x2=27.46 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=27.46 //y=0.625 //x2=27.46 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=26.575 //y=1.59 //x2=26.49 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.575 //y=1.59 //x2=26.975 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=27.375 //y=1.59 //x2=27.46 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=27.375 //y=1.59 //x2=26.975 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=26.49 //y=1.505 //x2=26.49 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=26.49 //y=1.505 //x2=26.49 //y2=0.89
ends PM_TMRDFFRNQNX1\%noxref_33

subckt PM_TMRDFFRNQNX1\%noxref_34 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=28.865 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=27.76 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=29 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=29.97 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=29.885 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=29 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=28.915 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=29.97 //y=0.625 //x2=29.97 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=29.97 //y=0.625 //x2=29.97 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=29.085 //y=0.54 //x2=29 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=29.085 //y=0.54 //x2=29.485 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=29.885 //y=0.54 //x2=29.97 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=29.885 //y=0.54 //x2=29.485 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=29 //y=1.08 //x2=29 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=29 //y=1.08 //x2=29 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=29 //y=0.91 //x2=29 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=29 //y=0.91 //x2=29 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=29 //y=0.625 //x2=29 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=29 //y=0.625 //x2=29 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.035 //y=0.995 //x2=27.95 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=28.915 //y=0.995 //x2=29 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=28.915 //y=0.995 //x2=28.035 //y2=0.995
ends PM_TMRDFFRNQNX1\%noxref_34

subckt PM_TMRDFFRNQNX1\%noxref_35 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=31.165 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=33.155 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=33.155 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=32.27 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=32.185 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=31.3 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=32.355 //y=1.59 //x2=32.27 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=32.355 //y=1.59 //x2=32.755 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.155 //y=1.59 //x2=33.24 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=33.155 //y=1.59 //x2=32.755 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=32.355 //y=0.54 //x2=32.27 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=32.355 //y=0.54 //x2=32.755 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.155 //y=0.54 //x2=33.24 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=33.155 //y=0.54 //x2=32.755 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=32.27 //y=1.505 //x2=32.27 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=32.27 //y=1.505 //x2=32.27 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=32.27 //y=0.625 //x2=32.27 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=32.27 //y=0.625 //x2=32.27 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=31.385 //y=1.59 //x2=31.3 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=31.385 //y=1.59 //x2=31.785 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=32.185 //y=1.59 //x2=32.27 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=32.185 //y=1.59 //x2=31.785 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=31.3 //y=1.505 //x2=31.3 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=31.3 //y=1.505 //x2=31.3 //y2=0.89
ends PM_TMRDFFRNQNX1\%noxref_35

subckt PM_TMRDFFRNQNX1\%noxref_36 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0413887f //x=33.675 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=32.57 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=33.81 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=34.78 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=34.695 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=33.81 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=33.725 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=34.78 //y=0.625 //x2=34.78 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=34.78 //y=0.625 //x2=34.78 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=33.895 //y=0.54 //x2=33.81 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=33.895 //y=0.54 //x2=34.295 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=34.695 //y=0.54 //x2=34.78 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=34.695 //y=0.54 //x2=34.295 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=33.81 //y=1.08 //x2=33.81 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=33.81 //y=1.08 //x2=33.81 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=33.81 //y=0.91 //x2=33.81 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=33.81 //y=0.91 //x2=33.81 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=33.81 //y=0.625 //x2=33.81 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=33.81 //y=0.625 //x2=33.81 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=32.845 //y=0.995 //x2=32.76 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=33.725 //y=0.995 //x2=33.81 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=33.725 //y=0.995 //x2=32.845 //y2=0.995
ends PM_TMRDFFRNQNX1\%noxref_36

subckt PM_TMRDFFRNQNX1\%noxref_37 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632682f //x=36.08 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=38.155 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=38.07 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=37.185 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=37.185 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=37.1 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=36.215 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=38.155 //y=0.615 //x2=38.155 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=38.155 //y=0.615 //x2=38.155 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=37.27 //y=0.53 //x2=37.185 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=37.27 //y=0.53 //x2=37.67 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=38.07 //y=0.53 //x2=38.155 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=38.07 //y=0.53 //x2=37.67 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=37.185 //y=1.495 //x2=37.185 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=37.185 //y=1.495 //x2=37.185 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=37.185 //y=0.615 //x2=37.185 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=37.185 //y=0.615 //x2=37.185 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=36.3 //y=1.58 //x2=36.215 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=36.3 //y=1.58 //x2=36.7 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=37.1 //y=1.58 //x2=37.185 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=37.1 //y=1.58 //x2=36.7 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=36.215 //y=1.495 //x2=36.215 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=36.215 //y=1.495 //x2=36.215 //y2=0.88
ends PM_TMRDFFRNQNX1\%noxref_37

subckt PM_TMRDFFRNQNX1\%noxref_38 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=39.305 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=41.295 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=41.295 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=40.41 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=40.325 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=39.44 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=40.495 //y=1.59 //x2=40.41 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=40.495 //y=1.59 //x2=40.895 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.295 //y=1.59 //x2=41.38 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=41.295 //y=1.59 //x2=40.895 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=40.495 //y=0.54 //x2=40.41 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=40.495 //y=0.54 //x2=40.895 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.295 //y=0.54 //x2=41.38 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=41.295 //y=0.54 //x2=40.895 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=40.41 //y=1.505 //x2=40.41 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=40.41 //y=1.505 //x2=40.41 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=40.41 //y=0.625 //x2=40.41 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=40.41 //y=0.625 //x2=40.41 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=39.525 //y=1.59 //x2=39.44 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=39.525 //y=1.59 //x2=39.925 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=40.325 //y=1.59 //x2=40.41 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=40.325 //y=1.59 //x2=39.925 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=39.44 //y=1.505 //x2=39.44 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=39.44 //y=1.505 //x2=39.44 //y2=0.89
ends PM_TMRDFFRNQNX1\%noxref_38

subckt PM_TMRDFFRNQNX1\%noxref_39 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0413887f //x=41.815 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=40.71 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=41.95 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=42.92 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=42.835 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=41.95 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=41.865 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=42.92 //y=0.625 //x2=42.92 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=42.92 //y=0.625 //x2=42.92 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=42.035 //y=0.54 //x2=41.95 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=42.035 //y=0.54 //x2=42.435 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=42.835 //y=0.54 //x2=42.92 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=42.835 //y=0.54 //x2=42.435 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=41.95 //y=1.08 //x2=41.95 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=41.95 //y=1.08 //x2=41.95 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=41.95 //y=0.91 //x2=41.95 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=41.95 //y=0.91 //x2=41.95 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=41.95 //y=0.625 //x2=41.95 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=41.95 //y=0.625 //x2=41.95 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.985 //y=0.995 //x2=40.9 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=41.865 //y=0.995 //x2=41.95 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=41.865 //y=0.995 //x2=40.985 //y2=0.995
ends PM_TMRDFFRNQNX1\%noxref_39

subckt PM_TMRDFFRNQNX1\%noxref_40 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=44.115 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=46.105 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=46.105 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=45.22 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=45.135 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=44.25 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=45.305 //y=1.59 //x2=45.22 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.305 //y=1.59 //x2=45.705 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.105 //y=1.59 //x2=46.19 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=46.105 //y=1.59 //x2=45.705 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=45.305 //y=0.54 //x2=45.22 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.305 //y=0.54 //x2=45.705 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.105 //y=0.54 //x2=46.19 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=46.105 //y=0.54 //x2=45.705 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=45.22 //y=1.505 //x2=45.22 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=45.22 //y=1.505 //x2=45.22 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=45.22 //y=0.625 //x2=45.22 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=45.22 //y=0.625 //x2=45.22 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=44.335 //y=1.59 //x2=44.25 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=44.335 //y=1.59 //x2=44.735 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=45.135 //y=1.59 //x2=45.22 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.135 //y=1.59 //x2=44.735 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=44.25 //y=1.505 //x2=44.25 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=44.25 //y=1.505 //x2=44.25 //y2=0.89
ends PM_TMRDFFRNQNX1\%noxref_40

subckt PM_TMRDFFRNQNX1\%noxref_41 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=46.625 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=45.52 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=46.76 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=47.73 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=47.645 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=46.76 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=46.675 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=47.73 //y=0.625 //x2=47.73 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=47.73 //y=0.625 //x2=47.73 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=46.845 //y=0.54 //x2=46.76 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=46.845 //y=0.54 //x2=47.245 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=47.645 //y=0.54 //x2=47.73 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=47.645 //y=0.54 //x2=47.245 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=46.76 //y=1.08 //x2=46.76 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=46.76 //y=1.08 //x2=46.76 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=46.76 //y=0.91 //x2=46.76 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=46.76 //y=0.91 //x2=46.76 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=46.76 //y=0.625 //x2=46.76 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=46.76 //y=0.625 //x2=46.76 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.795 //y=0.995 //x2=45.71 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=46.675 //y=0.995 //x2=46.76 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=46.675 //y=0.995 //x2=45.795 //y2=0.995
ends PM_TMRDFFRNQNX1\%noxref_41

subckt PM_TMRDFFRNQNX1\%noxref_42 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632682f //x=49.03 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=51.105 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=51.02 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=50.135 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=50.135 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=50.05 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=49.165 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=51.105 //y=0.615 //x2=51.105 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=51.105 //y=0.615 //x2=51.105 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=50.22 //y=0.53 //x2=50.135 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=50.22 //y=0.53 //x2=50.62 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=51.02 //y=0.53 //x2=51.105 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=51.02 //y=0.53 //x2=50.62 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=50.135 //y=1.495 //x2=50.135 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=50.135 //y=1.495 //x2=50.135 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=50.135 //y=0.615 //x2=50.135 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=50.135 //y=0.615 //x2=50.135 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=49.25 //y=1.58 //x2=49.165 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=49.25 //y=1.58 //x2=49.65 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=50.05 //y=1.58 //x2=50.135 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=50.05 //y=1.58 //x2=49.65 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=49.165 //y=1.495 //x2=49.165 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=49.165 //y=1.495 //x2=49.165 //y2=0.88
ends PM_TMRDFFRNQNX1\%noxref_42

subckt PM_TMRDFFRNQNX1\%noxref_43 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=52.255 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=54.245 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=54.245 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=53.36 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=53.275 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=52.39 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=53.445 //y=1.59 //x2=53.36 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=53.445 //y=1.59 //x2=53.845 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.245 //y=1.59 //x2=54.33 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.245 //y=1.59 //x2=53.845 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=53.445 //y=0.54 //x2=53.36 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=53.445 //y=0.54 //x2=53.845 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.245 //y=0.54 //x2=54.33 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.245 //y=0.54 //x2=53.845 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=53.36 //y=1.505 //x2=53.36 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=53.36 //y=1.505 //x2=53.36 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=53.36 //y=0.625 //x2=53.36 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=53.36 //y=0.625 //x2=53.36 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=52.475 //y=1.59 //x2=52.39 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=52.475 //y=1.59 //x2=52.875 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=53.275 //y=1.59 //x2=53.36 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=53.275 //y=1.59 //x2=52.875 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=52.39 //y=1.505 //x2=52.39 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=52.39 //y=1.505 //x2=52.39 //y2=0.89
ends PM_TMRDFFRNQNX1\%noxref_43

subckt PM_TMRDFFRNQNX1\%noxref_44 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=54.765 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=53.66 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=54.9 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=55.87 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=55.785 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=54.9 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=54.815 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=55.87 //y=0.625 //x2=55.87 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=55.87 //y=0.625 //x2=55.87 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=54.985 //y=0.54 //x2=54.9 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.985 //y=0.54 //x2=55.385 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=55.785 //y=0.54 //x2=55.87 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=55.785 //y=0.54 //x2=55.385 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=54.9 //y=1.08 //x2=54.9 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=54.9 //y=1.08 //x2=54.9 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=54.9 //y=0.91 //x2=54.9 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=54.9 //y=0.91 //x2=54.9 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=54.9 //y=0.625 //x2=54.9 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=54.9 //y=0.625 //x2=54.9 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.935 //y=0.995 //x2=53.85 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=54.815 //y=0.995 //x2=54.9 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=54.815 //y=0.995 //x2=53.935 //y2=0.995
ends PM_TMRDFFRNQNX1\%noxref_44

subckt PM_TMRDFFRNQNX1\%noxref_45 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=57.065 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=59.055 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=59.055 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=58.17 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=58.085 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=57.2 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=58.255 //y=1.59 //x2=58.17 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=58.255 //y=1.59 //x2=58.655 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.055 //y=1.59 //x2=59.14 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.055 //y=1.59 //x2=58.655 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=58.255 //y=0.54 //x2=58.17 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=58.255 //y=0.54 //x2=58.655 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.055 //y=0.54 //x2=59.14 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.055 //y=0.54 //x2=58.655 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=58.17 //y=1.505 //x2=58.17 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=58.17 //y=1.505 //x2=58.17 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=58.17 //y=0.625 //x2=58.17 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=58.17 //y=0.625 //x2=58.17 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=57.285 //y=1.59 //x2=57.2 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=57.285 //y=1.59 //x2=57.685 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=58.085 //y=1.59 //x2=58.17 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=58.085 //y=1.59 //x2=57.685 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=57.2 //y=1.505 //x2=57.2 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=57.2 //y=1.505 //x2=57.2 //y2=0.89
ends PM_TMRDFFRNQNX1\%noxref_45

subckt PM_TMRDFFRNQNX1\%noxref_46 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0413887f //x=59.575 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=58.47 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=59.71 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=60.68 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=60.595 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=59.71 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=59.625 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=60.68 //y=0.625 //x2=60.68 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=60.68 //y=0.625 //x2=60.68 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=59.795 //y=0.54 //x2=59.71 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.795 //y=0.54 //x2=60.195 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=60.595 //y=0.54 //x2=60.68 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=60.595 //y=0.54 //x2=60.195 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=59.71 //y=1.08 //x2=59.71 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=59.71 //y=1.08 //x2=59.71 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=59.71 //y=0.91 //x2=59.71 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=59.71 //y=0.91 //x2=59.71 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=59.71 //y=0.625 //x2=59.71 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=59.71 //y=0.625 //x2=59.71 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.745 //y=0.995 //x2=58.66 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=59.625 //y=0.995 //x2=59.71 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=59.625 //y=0.995 //x2=58.745 //y2=0.995
ends PM_TMRDFFRNQNX1\%noxref_46

subckt PM_TMRDFFRNQNX1\%noxref_47 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632682f //x=61.98 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=64.055 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=63.97 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=63.085 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=63.085 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=63 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=62.115 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=64.055 //y=0.615 //x2=64.055 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=64.055 //y=0.615 //x2=64.055 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=63.17 //y=0.53 //x2=63.085 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=63.17 //y=0.53 //x2=63.57 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=63.97 //y=0.53 //x2=64.055 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=63.97 //y=0.53 //x2=63.57 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=63.085 //y=1.495 //x2=63.085 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=63.085 //y=1.495 //x2=63.085 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=63.085 //y=0.615 //x2=63.085 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=63.085 //y=0.615 //x2=63.085 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=62.2 //y=1.58 //x2=62.115 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=62.2 //y=1.58 //x2=62.6 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=63 //y=1.58 //x2=63.085 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=63 //y=1.58 //x2=62.6 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=62.115 //y=1.495 //x2=62.115 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=62.115 //y=1.495 //x2=62.115 //y2=0.88
ends PM_TMRDFFRNQNX1\%noxref_47

subckt PM_TMRDFFRNQNX1\%noxref_48 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673029f //x=65.205 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=67.195 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=67.195 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=66.31 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=66.225 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=65.34 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=66.395 //y=1.59 //x2=66.31 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=66.395 //y=1.59 //x2=66.795 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.195 //y=1.59 //x2=67.28 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=67.195 //y=1.59 //x2=66.795 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=66.395 //y=0.54 //x2=66.31 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=66.395 //y=0.54 //x2=66.795 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.195 //y=0.54 //x2=67.28 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=67.195 //y=0.54 //x2=66.795 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=66.31 //y=1.505 //x2=66.31 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=66.31 //y=1.505 //x2=66.31 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=66.31 //y=0.625 //x2=66.31 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=66.31 //y=0.625 //x2=66.31 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=65.425 //y=1.59 //x2=65.34 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=65.425 //y=1.59 //x2=65.825 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=66.225 //y=1.59 //x2=66.31 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=66.225 //y=1.59 //x2=65.825 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=65.34 //y=1.505 //x2=65.34 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=65.34 //y=1.505 //x2=65.34 //y2=0.89
ends PM_TMRDFFRNQNX1\%noxref_48

subckt PM_TMRDFFRNQNX1\%noxref_49 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.0413887f //x=67.715 //y=0.375
c54 ( 28 0 ) capacitor c=0.0045748f //x=66.61 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=67.85 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=68.82 //y=0.625
c57 ( 11 0 ) capacitor c=0.0144218f //x=68.735 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=67.85 //y=0.625
c59 ( 1 0 ) capacitor c=0.0218888f //x=67.765 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=68.82 //y=0.625 //x2=68.82 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=68.82 //y=0.625 //x2=68.82 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=67.935 //y=0.54 //x2=67.85 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=67.935 //y=0.54 //x2=68.335 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=68.735 //y=0.54 //x2=68.82 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=68.735 //y=0.54 //x2=68.335 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=67.85 //y=1.08 //x2=67.85 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=67.85 //y=1.08 //x2=67.85 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=67.85 //y=0.91 //x2=67.85 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=67.85 //y=0.91 //x2=67.85 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=67.85 //y=0.625 //x2=67.85 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=67.85 //y=0.625 //x2=67.85 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.885 //y=0.995 //x2=66.8 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=67.765 //y=0.995 //x2=67.85 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=67.765 //y=0.995 //x2=66.885 //y2=0.995
ends PM_TMRDFFRNQNX1\%noxref_49

subckt PM_TMRDFFRNQNX1\%noxref_50 ( 1 5 9 13 17 35 )
c51 ( 35 0 ) capacitor c=0.0680259f //x=70.015 //y=0.375
c52 ( 17 0 ) capacitor c=0.0180446f //x=72.005 //y=1.59
c53 ( 13 0 ) capacitor c=0.0155283f //x=72.005 //y=0.54
c54 ( 9 0 ) capacitor c=0.00678203f //x=71.12 //y=0.625
c55 ( 5 0 ) capacitor c=0.0164013f //x=71.035 //y=1.59
c56 ( 1 0 ) capacitor c=0.00696517f //x=70.15 //y=1.505
r57 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=71.205 //y=1.59 //x2=71.12 //y2=1.63
r58 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=71.205 //y=1.59 //x2=71.605 //y2=1.59
r59 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.005 //y=1.59 //x2=72.09 //y2=1.59
r60 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=72.005 //y=1.59 //x2=71.605 //y2=1.59
r61 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=71.205 //y=0.54 //x2=71.12 //y2=0.5
r62 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=71.205 //y=0.54 //x2=71.605 //y2=0.54
r63 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.005 //y=0.54 //x2=72.09 //y2=0.54
r64 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=72.005 //y=0.54 //x2=71.605 //y2=0.54
r65 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=71.12 //y=1.505 //x2=71.12 //y2=1.63
r66 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=71.12 //y=1.505 //x2=71.12 //y2=0.89
r67 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=71.12 //y=0.625 //x2=71.12 //y2=0.5
r68 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=71.12 //y=0.625 //x2=71.12 //y2=0.89
r69 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=70.235 //y=1.59 //x2=70.15 //y2=1.63
r70 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=70.235 //y=1.59 //x2=70.635 //y2=1.59
r71 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=71.035 //y=1.59 //x2=71.12 //y2=1.63
r72 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=71.035 //y=1.59 //x2=70.635 //y2=1.59
r73 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=70.15 //y=1.505 //x2=70.15 //y2=1.63
r74 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=70.15 //y=1.505 //x2=70.15 //y2=0.89
ends PM_TMRDFFRNQNX1\%noxref_50

subckt PM_TMRDFFRNQNX1\%noxref_51 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0421963f //x=72.525 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=71.42 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=72.66 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=73.63 //y=0.625
c56 ( 11 0 ) capacitor c=0.014695f //x=73.545 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=72.66 //y=0.625
c58 ( 1 0 ) capacitor c=0.0234159f //x=72.575 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=73.63 //y=0.625 //x2=73.63 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=73.63 //y=0.625 //x2=73.63 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=72.745 //y=0.54 //x2=72.66 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=72.745 //y=0.54 //x2=73.145 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=73.545 //y=0.54 //x2=73.63 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=73.545 //y=0.54 //x2=73.145 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=72.66 //y=1.08 //x2=72.66 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=72.66 //y=1.08 //x2=72.66 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=72.66 //y=0.91 //x2=72.66 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=72.66 //y=0.91 //x2=72.66 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=72.66 //y=0.625 //x2=72.66 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=72.66 //y=0.625 //x2=72.66 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.695 //y=0.995 //x2=71.61 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=72.575 //y=0.995 //x2=72.66 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=72.575 //y=0.995 //x2=71.695 //y2=0.995
ends PM_TMRDFFRNQNX1\%noxref_51

subckt PM_TMRDFFRNQNX1\%noxref_52 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0634202f //x=74.93 //y=0.365
c52 ( 17 0 ) capacitor c=0.00722223f //x=77.005 //y=0.615
c53 ( 13 0 ) capacitor c=0.0147854f //x=76.92 //y=0.53
c54 ( 10 0 ) capacitor c=0.00638095f //x=76.035 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=76.035 //y=0.615
c56 ( 5 0 ) capacitor c=0.0189075f //x=75.95 //y=1.58
c57 ( 1 0 ) capacitor c=0.00798521f //x=75.065 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=77.005 //y=0.615 //x2=77.005 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=77.005 //y=0.615 //x2=77.005 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=76.12 //y=0.53 //x2=76.035 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=76.12 //y=0.53 //x2=76.52 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=76.92 //y=0.53 //x2=77.005 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=76.92 //y=0.53 //x2=76.52 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=76.035 //y=1.495 //x2=76.035 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=76.035 //y=1.495 //x2=76.035 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=76.035 //y=0.615 //x2=76.035 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=76.035 //y=0.615 //x2=76.035 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=75.15 //y=1.58 //x2=75.065 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=75.15 //y=1.58 //x2=75.55 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=75.95 //y=1.58 //x2=76.035 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=75.95 //y=1.58 //x2=75.55 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=75.065 //y=1.495 //x2=75.065 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=75.065 //y=1.495 //x2=75.065 //y2=0.88
ends PM_TMRDFFRNQNX1\%noxref_52

subckt PM_TMRDFFRNQNX1\%noxref_53 ( 1 5 9 10 13 17 29 )
c57 ( 29 0 ) capacitor c=0.0758145f //x=78.26 //y=0.365
c58 ( 17 0 ) capacitor c=0.0072249f //x=80.335 //y=0.615
c59 ( 13 0 ) capacitor c=0.0153682f //x=80.25 //y=0.53
c60 ( 10 0 ) capacitor c=0.00754305f //x=79.365 //y=1.495
c61 ( 9 0 ) capacitor c=0.006761f //x=79.365 //y=0.615
c62 ( 5 0 ) capacitor c=0.0213241f //x=79.28 //y=1.58
c63 ( 1 0 ) capacitor c=0.00492513f //x=78.395 //y=1.495
r64 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=80.335 //y=0.615 //x2=80.335 //y2=0.49
r65 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=80.335 //y=0.615 //x2=80.335 //y2=1.22
r66 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=79.45 //y=0.53 //x2=79.365 //y2=0.49
r67 (  14 29 ) resistor r=27.0374 //w=0.187 //l=0.395 //layer=li \
 //thickness=0.1 //x=79.45 //y=0.53 //x2=79.845 //y2=0.53
r68 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=80.25 //y=0.53 //x2=80.335 //y2=0.49
r69 (  13 29 ) resistor r=27.7219 //w=0.187 //l=0.405 //layer=li \
 //thickness=0.1 //x=80.25 //y=0.53 //x2=79.845 //y2=0.53
r70 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=79.365 //y=1.495 //x2=79.365 //y2=1.62
r71 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=79.365 //y=1.495 //x2=79.365 //y2=0.88
r72 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=79.365 //y=0.615 //x2=79.365 //y2=0.49
r73 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=79.365 //y=0.615 //x2=79.365 //y2=0.88
r74 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.48 //y=1.58 //x2=78.395 //y2=1.62
r75 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=78.48 //y=1.58 //x2=78.88 //y2=1.58
r76 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=79.28 //y=1.58 //x2=79.365 //y2=1.62
r77 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=79.28 //y=1.58 //x2=78.88 //y2=1.58
r78 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=78.395 //y=1.495 //x2=78.395 //y2=1.62
r79 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=78.395 //y=1.495 //x2=78.395 //y2=0.88
ends PM_TMRDFFRNQNX1\%noxref_53

subckt PM_TMRDFFRNQNX1\%noxref_54 ( 1 5 9 10 13 17 29 )
c55 ( 29 0 ) capacitor c=0.0723103f //x=81.59 //y=0.365
c56 ( 17 0 ) capacitor c=0.0072249f //x=83.665 //y=0.615
c57 ( 13 0 ) capacitor c=0.0155051f //x=83.58 //y=0.53
c58 ( 10 0 ) capacitor c=0.00876912f //x=82.695 //y=1.495
c59 ( 9 0 ) capacitor c=0.006761f //x=82.695 //y=0.615
c60 ( 5 0 ) capacitor c=0.0182818f //x=82.61 //y=1.58
c61 ( 1 0 ) capacitor c=0.00857722f //x=81.725 //y=1.495
r62 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=83.665 //y=0.615 //x2=83.665 //y2=0.49
r63 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=83.665 //y=0.615 //x2=83.665 //y2=1.22
r64 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=82.78 //y=0.53 //x2=82.695 //y2=0.49
r65 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=82.78 //y=0.53 //x2=83.18 //y2=0.53
r66 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=83.58 //y=0.53 //x2=83.665 //y2=0.49
r67 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=83.58 //y=0.53 //x2=83.18 //y2=0.53
r68 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=82.695 //y=1.495 //x2=82.695 //y2=1.62
r69 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=82.695 //y=1.495 //x2=82.695 //y2=0.88
r70 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=82.695 //y=0.615 //x2=82.695 //y2=0.49
r71 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=82.695 //y=0.615 //x2=82.695 //y2=0.88
r72 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=81.81 //y=1.58 //x2=81.725 //y2=1.62
r73 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=81.81 //y=1.58 //x2=82.21 //y2=1.58
r74 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=82.61 //y=1.58 //x2=82.695 //y2=1.62
r75 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=82.61 //y=1.58 //x2=82.21 //y2=1.58
r76 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=81.725 //y=1.495 //x2=81.725 //y2=1.62
r77 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=81.725 //y=1.495 //x2=81.725 //y2=0.88
ends PM_TMRDFFRNQNX1\%noxref_54

subckt PM_TMRDFFRNQNX1\%noxref_55 ( 1 5 9 10 13 17 29 )
c53 ( 29 0 ) capacitor c=0.0643725f //x=84.92 //y=0.365
c54 ( 17 0 ) capacitor c=0.00722228f //x=86.995 //y=0.615
c55 ( 13 0 ) capacitor c=0.0141607f //x=86.91 //y=0.53
c56 ( 10 0 ) capacitor c=0.00712138f //x=86.025 //y=1.495
c57 ( 9 0 ) capacitor c=0.006761f //x=86.025 //y=0.615
c58 ( 5 0 ) capacitor c=0.0233454f //x=85.94 //y=1.58
c59 ( 1 0 ) capacitor c=0.00481264f //x=85.055 //y=1.495
r60 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=86.995 //y=0.615 //x2=86.995 //y2=0.49
r61 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=86.995 //y=0.615 //x2=86.995 //y2=0.88
r62 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=86.11 //y=0.53 //x2=86.025 //y2=0.49
r63 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=86.11 //y=0.53 //x2=86.51 //y2=0.53
r64 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=86.91 //y=0.53 //x2=86.995 //y2=0.49
r65 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=86.91 //y=0.53 //x2=86.51 //y2=0.53
r66 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=86.025 //y=1.495 //x2=86.025 //y2=1.62
r67 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=86.025 //y=1.495 //x2=86.025 //y2=0.88
r68 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=86.025 //y=0.615 //x2=86.025 //y2=0.49
r69 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=86.025 //y=0.615 //x2=86.025 //y2=0.88
r70 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=85.14 //y=1.58 //x2=85.055 //y2=1.62
r71 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=85.14 //y=1.58 //x2=85.54 //y2=1.58
r72 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=85.94 //y=1.58 //x2=86.025 //y2=1.62
r73 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=85.94 //y=1.58 //x2=85.54 //y2=1.58
r74 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=85.055 //y=1.495 //x2=85.055 //y2=1.62
r75 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=85.055 //y=1.495 //x2=85.055 //y2=0.88
ends PM_TMRDFFRNQNX1\%noxref_55

