// File: pmos2.spi.pex
// Created: Tue Oct 15 16:00:16 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_PMOS2\%noxref_4 ( 1 2 6 )
c5 ( 7 0 ) capacitor c=0.0190444f //x=0.87 //y=-2.23
c6 ( 6 0 ) capacitor c=0.0437181f //x=1.16 //y=-2.23
c7 ( 2 0 ) capacitor c=0.168116f //x=1.235 //y=-1
c8 ( 1 0 ) capacitor c=0.168116f //x=0.795 //y=-1
r9 (  6 8 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.16 //y=-2.23 //x2=1.235 //y2=-2.155
r10 (  6 7 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.16 //y=-2.23 //x2=0.87 //y2=-2.23
r11 (  3 7 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=0.795 //y=-2.155 //x2=0.87 //y2=-2.23
r12 (  2 8 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.235 //y=-1 //x2=1.235 //y2=-2.155
r13 (  1 3 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=0.795 //y=-1 //x2=0.795 //y2=-2.155
ends PM_PMOS2\%noxref_4

