* SPICE3 file created from HA.ext - technology: sky130A

.subckt HA SUM COUT A B VDD GND
X0 SUM B a_1666_74 GND nshort w=3 l=0.15
X1 VDD B a_217_1004 VDD pshort w=2 l=0.15 M=2
X2 SUM a_1917_943 a_1685_1004 VDD pshort w=2 l=0.15 M=2
X3 GND A a_112_73 GND nshort w=3 l=0.15
X4 COUT a_217_1004 GND GND nshort w=3 l=0.15
X5 GND a_1917_943 a_2332_74 GND nshort w=3 l=0.15
X6 VDD A a_1685_1004 VDD pshort w=2 l=0.15 M=2
X7 VDD a_217_1004 COUT VDD pshort w=2 l=0.15 M=2
X8 a_1917_943 B GND GND nshort w=3 l=0.15
X9 VDD A a_1295_182 VDD pshort w=2 l=0.15 M=2
X10 a_2351_1004 B VDD VDD pshort w=2 l=0.15 M=2
X11 a_217_1004 A VDD VDD pshort w=2 l=0.15 M=2
X12 a_217_1004 B a_112_73 GND nshort w=3 l=0.15
X13 a_2351_1004 a_1295_182 SUM VDD pshort w=2 l=0.15 M=2
X14 VDD B a_1917_943 VDD pshort w=2 l=0.15 M=2
X15 SUM a_1295_182 a_2332_74 GND nshort w=3 l=0.15
X16 GND A a_1666_74 GND nshort w=3 l=0.15
X17 a_1295_182 A GND GND nshort w=3 l=0.15
C0 a_1917_943 B 2.85fF
C1 A B 2.08fF
C2 VDD GND 8.25fF
.ends
