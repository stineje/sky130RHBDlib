* SPICE3 file created from VOTER3X1.ext - technology: sky130A

.subckt VOTER3X1 Y A B C VDD GND
X0 GND B a_112_73 GND nshort w=3 l=0.15
X1 GND C a_1444_73 GND nshort w=3 l=0.15
X2 a_392_181 A a_1444_73 GND nshort w=3 l=0.15
X3 a_392_181 A a_881_1005 VDD pshort w=2 l=0.15 M=2
X4 VDD a_392_181 Y VDD pshort w=2 l=0.15 M=2
X5 VDD B a_217_1005 VDD pshort w=2 l=0.15 M=2
X6 a_881_1005 C a_217_1005 VDD pshort w=2 l=0.15 M=2
X7 VDD A a_217_1005 VDD pshort w=2 l=0.15 M=2
X8 a_392_181 A a_112_73 GND nshort w=3 l=0.15
X9 a_881_1005 B a_217_1005 VDD pshort w=2 l=0.15 M=2
X10 a_881_1005 C a_392_181 VDD pshort w=2 l=0.15 M=2
X11 a_392_181 C a_778_73 GND nshort w=3 l=0.15
X12 Y a_392_181 GND GND nshort w=3 l=0.15
X13 GND B a_778_73 GND nshort w=3 l=0.15
C0 VDD GND 6.15fF
.ends
