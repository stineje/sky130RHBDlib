// File: TMRDFFSNQX1.spi.pex
// Created: Tue Oct 15 15:52:45 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_TMRDFFSNQX1\%GND ( 1 143 147 150 155 163 169 179 185 195 201 207 215 \
 223 231 241 249 257 263 273 279 289 295 301 309 317 325 335 343 351 357 367 \
 373 383 389 395 403 411 419 429 437 445 451 457 465 476 481 485 498 501 504 \
 507 509 511 513 516 519 522 524 526 528 531 534 537 539 541 543 546 548 555 \
 562 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 \
 581 582 583 )
c1011 ( 583 0 ) capacitor c=0.0604367f //x=83.745 //y=0.37
c1012 ( 582 0 ) capacitor c=0.0215012f //x=80.91 //y=0.865
c1013 ( 581 0 ) capacitor c=0.0215012f //x=77.58 //y=0.865
c1014 ( 580 0 ) capacitor c=0.0207524f //x=74.25 //y=0.865
c1015 ( 579 0 ) capacitor c=0.0226075f //x=69.335 //y=0.875
c1016 ( 578 0 ) capacitor c=0.0207407f //x=66.11 //y=0.865
c1017 ( 577 0 ) capacitor c=0.0207407f //x=62.78 //y=0.865
c1018 ( 576 0 ) capacitor c=0.0225954f //x=57.865 //y=0.875
c1019 ( 575 0 ) capacitor c=0.0226075f //x=53.055 //y=0.875
c1020 ( 574 0 ) capacitor c=0.0207407f //x=49.83 //y=0.865
c1021 ( 573 0 ) capacitor c=0.0226075f //x=44.915 //y=0.875
c1022 ( 572 0 ) capacitor c=0.0207407f //x=41.69 //y=0.865
c1023 ( 571 0 ) capacitor c=0.0207407f //x=38.36 //y=0.865
c1024 ( 570 0 ) capacitor c=0.0225954f //x=33.445 //y=0.875
c1025 ( 569 0 ) capacitor c=0.0226075f //x=28.635 //y=0.875
c1026 ( 568 0 ) capacitor c=0.0207407f //x=25.41 //y=0.865
c1027 ( 567 0 ) capacitor c=0.0226075f //x=20.495 //y=0.875
c1028 ( 566 0 ) capacitor c=0.0207407f //x=17.27 //y=0.865
c1029 ( 565 0 ) capacitor c=0.0207407f //x=13.94 //y=0.865
c1030 ( 564 0 ) capacitor c=0.0226205f //x=9.025 //y=0.875
c1031 ( 563 0 ) capacitor c=0.0226323f //x=4.215 //y=0.875
c1032 ( 562 0 ) capacitor c=0.0207863f //x=0.99 //y=0.865
c1033 ( 555 0 ) capacitor c=0.234368f //x=84.85 //y=0
c1034 ( 548 0 ) capacitor c=0.101943f //x=83.25 //y=0
c1035 ( 547 0 ) capacitor c=0.00440095f //x=81.1 //y=0
c1036 ( 546 0 ) capacitor c=0.101477f //x=79.92 //y=0
c1037 ( 545 0 ) capacitor c=0.00440095f //x=77.7 //y=0
c1038 ( 543 0 ) capacitor c=0.116995f //x=76.59 //y=0
c1039 ( 542 0 ) capacitor c=0.00440095f //x=74.44 //y=0
c1040 ( 541 0 ) capacitor c=0.106826f //x=73.26 //y=0
c1041 ( 540 0 ) capacitor c=0.00440144f //x=69.525 //y=0
c1042 ( 539 0 ) capacitor c=0.104091f //x=68.45 //y=0
c1043 ( 538 0 ) capacitor c=0.00440095f //x=66.3 //y=0
c1044 ( 537 0 ) capacitor c=0.105123f //x=65.12 //y=0
c1045 ( 536 0 ) capacitor c=0.00440095f //x=62.9 //y=0
c1046 ( 534 0 ) capacitor c=0.108248f //x=61.79 //y=0
c1047 ( 533 0 ) capacitor c=0.00440144f //x=58.09 //y=0
c1048 ( 531 0 ) capacitor c=0.107229f //x=56.98 //y=0
c1049 ( 530 0 ) capacitor c=0.00440144f //x=53.28 //y=0
c1050 ( 528 0 ) capacitor c=0.104113f //x=52.17 //y=0
c1051 ( 527 0 ) capacitor c=0.00440095f //x=50.02 //y=0
c1052 ( 526 0 ) capacitor c=0.108351f //x=48.84 //y=0
c1053 ( 525 0 ) capacitor c=0.00440144f //x=45.105 //y=0
c1054 ( 524 0 ) capacitor c=0.10408f //x=44.03 //y=0
c1055 ( 523 0 ) capacitor c=0.00440095f //x=41.88 //y=0
c1056 ( 522 0 ) capacitor c=0.104882f //x=40.7 //y=0
c1057 ( 521 0 ) capacitor c=0.00440095f //x=38.48 //y=0
c1058 ( 519 0 ) capacitor c=0.108248f //x=37.37 //y=0
c1059 ( 518 0 ) capacitor c=0.00440144f //x=33.67 //y=0
c1060 ( 516 0 ) capacitor c=0.107229f //x=32.56 //y=0
c1061 ( 515 0 ) capacitor c=0.00440144f //x=28.86 //y=0
c1062 ( 513 0 ) capacitor c=0.104143f //x=27.75 //y=0
c1063 ( 512 0 ) capacitor c=0.00440095f //x=25.6 //y=0
c1064 ( 511 0 ) capacitor c=0.108018f //x=24.42 //y=0
c1065 ( 510 0 ) capacitor c=0.00440144f //x=20.685 //y=0
c1066 ( 509 0 ) capacitor c=0.104091f //x=19.61 //y=0
c1067 ( 508 0 ) capacitor c=0.00440095f //x=17.46 //y=0
c1068 ( 507 0 ) capacitor c=0.105123f //x=16.28 //y=0
c1069 ( 506 0 ) capacitor c=0.00440095f //x=14.06 //y=0
c1070 ( 504 0 ) capacitor c=0.108248f //x=12.95 //y=0
c1071 ( 503 0 ) capacitor c=0.00440144f //x=9.25 //y=0
c1072 ( 501 0 ) capacitor c=0.108235f //x=8.14 //y=0
c1073 ( 500 0 ) capacitor c=0.00440144f //x=4.44 //y=0
c1074 ( 498 0 ) capacitor c=0.105313f //x=3.33 //y=0
c1075 ( 497 0 ) capacitor c=0.00440095f //x=1.18 //y=0
c1076 ( 488 0 ) capacitor c=0.00583665f //x=84.85 //y=0.45
c1077 ( 485 0 ) capacitor c=0.00542558f //x=84.765 //y=0.535
c1078 ( 484 0 ) capacitor c=0.00479856f //x=84.365 //y=0.45
c1079 ( 481 0 ) capacitor c=0.00707849f //x=84.28 //y=0.535
c1080 ( 476 0 ) capacitor c=0.00588377f //x=83.88 //y=0.45
c1081 ( 473 0 ) capacitor c=0.0190475f //x=83.795 //y=0
c1082 ( 465 0 ) capacitor c=0.0749789f //x=83.08 //y=0
c1083 ( 457 0 ) capacitor c=0.0389876f //x=81.015 //y=0
c1084 ( 451 0 ) capacitor c=0.0716428f //x=79.75 //y=0
c1085 ( 445 0 ) capacitor c=0.0388276f //x=77.685 //y=0
c1086 ( 437 0 ) capacitor c=0.071962f //x=76.42 //y=0
c1087 ( 429 0 ) capacitor c=0.0391432f //x=74.355 //y=0
c1088 ( 419 0 ) capacitor c=0.133607f //x=73.09 //y=0
c1089 ( 411 0 ) capacitor c=0.0339325f //x=69.44 //y=0
c1090 ( 403 0 ) capacitor c=0.0718026f //x=68.28 //y=0
c1091 ( 395 0 ) capacitor c=0.0388888f //x=66.215 //y=0
c1092 ( 389 0 ) capacitor c=0.0718026f //x=64.95 //y=0
c1093 ( 383 0 ) capacitor c=0.0388888f //x=62.885 //y=0
c1094 ( 373 0 ) capacitor c=0.133362f //x=61.62 //y=0
c1095 ( 367 0 ) capacitor c=0.0339325f //x=57.97 //y=0
c1096 ( 357 0 ) capacitor c=0.133362f //x=56.81 //y=0
c1097 ( 351 0 ) capacitor c=0.0339325f //x=53.16 //y=0
c1098 ( 343 0 ) capacitor c=0.0718026f //x=52 //y=0
c1099 ( 335 0 ) capacitor c=0.0388888f //x=49.935 //y=0
c1100 ( 325 0 ) capacitor c=0.133362f //x=48.67 //y=0
c1101 ( 317 0 ) capacitor c=0.0339325f //x=45.02 //y=0
c1102 ( 309 0 ) capacitor c=0.0718026f //x=43.86 //y=0
c1103 ( 301 0 ) capacitor c=0.0388888f //x=41.795 //y=0
c1104 ( 295 0 ) capacitor c=0.0718026f //x=40.53 //y=0
c1105 ( 289 0 ) capacitor c=0.0388888f //x=38.465 //y=0
c1106 ( 279 0 ) capacitor c=0.133362f //x=37.2 //y=0
c1107 ( 273 0 ) capacitor c=0.0339325f //x=33.55 //y=0
c1108 ( 263 0 ) capacitor c=0.133362f //x=32.39 //y=0
c1109 ( 257 0 ) capacitor c=0.0339325f //x=28.74 //y=0
c1110 ( 249 0 ) capacitor c=0.0718026f //x=27.58 //y=0
c1111 ( 241 0 ) capacitor c=0.0388888f //x=25.515 //y=0
c1112 ( 231 0 ) capacitor c=0.133362f //x=24.25 //y=0
c1113 ( 223 0 ) capacitor c=0.0339325f //x=20.6 //y=0
c1114 ( 215 0 ) capacitor c=0.0718026f //x=19.44 //y=0
c1115 ( 207 0 ) capacitor c=0.0388888f //x=17.375 //y=0
c1116 ( 201 0 ) capacitor c=0.0718026f //x=16.11 //y=0
c1117 ( 195 0 ) capacitor c=0.0388888f //x=14.045 //y=0
c1118 ( 185 0 ) capacitor c=0.133404f //x=12.78 //y=0
c1119 ( 179 0 ) capacitor c=0.0339482f //x=9.13 //y=0
c1120 ( 169 0 ) capacitor c=0.133515f //x=7.97 //y=0
c1121 ( 163 0 ) capacitor c=0.0339482f //x=4.32 //y=0
c1122 ( 155 0 ) capacitor c=0.0720441f //x=3.16 //y=0
c1123 ( 150 0 ) capacitor c=0.179262f //x=0.74 //y=0
c1124 ( 147 0 ) capacitor c=0.0426751f //x=1.095 //y=0
c1125 ( 143 0 ) capacitor c=2.59091f //x=84.73 //y=0
r1126 (  554 555 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=84.73 //y=0 //x2=84.85 //y2=0
r1127 (  552 554 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=84.365 //y=0 //x2=84.73 //y2=0
r1128 (  551 552 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=83.99 //y=0 //x2=84.365 //y2=0
r1129 (  549 551 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=83.88 //y=0 //x2=83.99 //y2=0
r1130 (  489 583 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.85 //y=0.62 //x2=84.85 //y2=0.535
r1131 (  489 583 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=84.85 //y=0.62 //x2=84.85 //y2=1.225
r1132 (  488 583 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.85 //y=0.45 //x2=84.85 //y2=0.535
r1133 (  487 555 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=84.85 //y=0.17 //x2=84.85 //y2=0
r1134 (  487 488 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=84.85 //y=0.17 //x2=84.85 //y2=0.45
r1135 (  486 583 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.45 //y=0.535 //x2=84.365 //y2=0.535
r1136 (  485 583 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.765 //y=0.535 //x2=84.85 //y2=0.535
r1137 (  485 486 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=84.765 //y=0.535 //x2=84.45 //y2=0.535
r1138 (  484 583 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.365 //y=0.45 //x2=84.365 //y2=0.535
r1139 (  483 552 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=84.365 //y=0.17 //x2=84.365 //y2=0
r1140 (  483 484 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=84.365 //y=0.17 //x2=84.365 //y2=0.45
r1141 (  482 583 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=83.965 //y=0.535 //x2=83.88 //y2=0.535
r1142 (  481 583 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.28 //y=0.535 //x2=84.365 //y2=0.535
r1143 (  481 482 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=84.28 //y=0.535 //x2=83.965 //y2=0.535
r1144 (  477 583 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=83.88 //y=0.62 //x2=83.88 //y2=0.535
r1145 (  477 583 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=83.88 //y=0.62 //x2=83.88 //y2=1.225
r1146 (  476 583 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=83.88 //y=0.45 //x2=83.88 //y2=0.535
r1147 (  475 549 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=83.88 //y=0.17 //x2=83.88 //y2=0
r1148 (  475 476 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=83.88 //y=0.17 //x2=83.88 //y2=0.45
r1149 (  474 548 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=83.42 //y=0 //x2=83.25 //y2=0
r1150 (  473 549 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=83.795 //y=0 //x2=83.88 //y2=0
r1151 (  473 474 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=83.795 //y=0 //x2=83.42 //y2=0
r1152 (  468 470 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=81.4 //y=0 //x2=82.51 //y2=0
r1153 (  466 547 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.185 //y=0 //x2=81.1 //y2=0
r1154 (  466 468 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=81.185 //y=0 //x2=81.4 //y2=0
r1155 (  465 548 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=83.08 //y=0 //x2=83.25 //y2=0
r1156 (  465 470 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=83.08 //y=0 //x2=82.51 //y2=0
r1157 (  461 547 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=81.1 //y=0.17 //x2=81.1 //y2=0
r1158 (  461 582 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=81.1 //y=0.17 //x2=81.1 //y2=0.955
r1159 (  458 546 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=80.09 //y=0 //x2=79.92 //y2=0
r1160 (  458 460 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=80.09 //y=0 //x2=80.29 //y2=0
r1161 (  457 547 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.015 //y=0 //x2=81.1 //y2=0
r1162 (  457 460 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=81.015 //y=0 //x2=80.29 //y2=0
r1163 (  452 545 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=77.855 //y=0 //x2=77.77 //y2=0
r1164 (  452 454 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=77.855 //y=0 //x2=78.81 //y2=0
r1165 (  451 546 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=79.75 //y=0 //x2=79.92 //y2=0
r1166 (  451 454 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=79.75 //y=0 //x2=78.81 //y2=0
r1167 (  447 545 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=77.77 //y=0.17 //x2=77.77 //y2=0
r1168 (  447 581 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=77.77 //y=0.17 //x2=77.77 //y2=0.955
r1169 (  446 543 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.76 //y=0 //x2=76.59 //y2=0
r1170 (  445 545 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=77.685 //y=0 //x2=77.77 //y2=0
r1171 (  445 446 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=77.685 //y=0 //x2=76.76 //y2=0
r1172 (  440 442 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=75.11 //y=0 //x2=76.22 //y2=0
r1173 (  438 542 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.525 //y=0 //x2=74.44 //y2=0
r1174 (  438 440 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=74.525 //y=0 //x2=75.11 //y2=0
r1175 (  437 543 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.42 //y=0 //x2=76.59 //y2=0
r1176 (  437 442 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=76.42 //y=0 //x2=76.22 //y2=0
r1177 (  433 542 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=74.44 //y=0.17 //x2=74.44 //y2=0
r1178 (  433 580 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=74.44 //y=0.17 //x2=74.44 //y2=0.955
r1179 (  430 541 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.43 //y=0 //x2=73.26 //y2=0
r1180 (  430 432 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=73.43 //y=0 //x2=74 //y2=0
r1181 (  429 542 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.355 //y=0 //x2=74.44 //y2=0
r1182 (  429 432 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=74.355 //y=0 //x2=74 //y2=0
r1183 (  424 426 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=71.41 //y=0 //x2=72.52 //y2=0
r1184 (  422 424 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=70.3 //y=0 //x2=71.41 //y2=0
r1185 (  420 540 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.61 //y=0 //x2=69.525 //y2=0
r1186 (  420 422 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=69.61 //y=0 //x2=70.3 //y2=0
r1187 (  419 541 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.09 //y=0 //x2=73.26 //y2=0
r1188 (  419 426 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=73.09 //y=0 //x2=72.52 //y2=0
r1189 (  415 540 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=69.525 //y=0.17 //x2=69.525 //y2=0
r1190 (  415 579 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=69.525 //y=0.17 //x2=69.525 //y2=0.965
r1191 (  412 539 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.62 //y=0 //x2=68.45 //y2=0
r1192 (  412 414 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=68.62 //y=0 //x2=69.19 //y2=0
r1193 (  411 540 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.44 //y=0 //x2=69.525 //y2=0
r1194 (  411 414 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=69.44 //y=0 //x2=69.19 //y2=0
r1195 (  406 408 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=66.6 //y=0 //x2=67.71 //y2=0
r1196 (  404 538 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.385 //y=0 //x2=66.3 //y2=0
r1197 (  404 406 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=66.385 //y=0 //x2=66.6 //y2=0
r1198 (  403 539 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.28 //y=0 //x2=68.45 //y2=0
r1199 (  403 408 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=68.28 //y=0 //x2=67.71 //y2=0
r1200 (  399 538 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=66.3 //y=0.17 //x2=66.3 //y2=0
r1201 (  399 578 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=66.3 //y=0.17 //x2=66.3 //y2=0.955
r1202 (  396 537 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=65.29 //y=0 //x2=65.12 //y2=0
r1203 (  396 398 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=65.29 //y=0 //x2=65.49 //y2=0
r1204 (  395 538 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.215 //y=0 //x2=66.3 //y2=0
r1205 (  395 398 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=66.215 //y=0 //x2=65.49 //y2=0
r1206 (  390 536 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.055 //y=0 //x2=62.97 //y2=0
r1207 (  390 392 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=63.055 //y=0 //x2=64.01 //y2=0
r1208 (  389 537 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.95 //y=0 //x2=65.12 //y2=0
r1209 (  389 392 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=64.95 //y=0 //x2=64.01 //y2=0
r1210 (  385 536 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.97 //y=0.17 //x2=62.97 //y2=0
r1211 (  385 577 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=62.97 //y=0.17 //x2=62.97 //y2=0.955
r1212 (  384 534 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.96 //y=0 //x2=61.79 //y2=0
r1213 (  383 536 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.885 //y=0 //x2=62.97 //y2=0
r1214 (  383 384 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=62.885 //y=0 //x2=61.96 //y2=0
r1215 (  378 380 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=60.31 //y=0 //x2=61.42 //y2=0
r1216 (  376 378 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=59.2 //y=0 //x2=60.31 //y2=0
r1217 (  374 533 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.14 //y=0 //x2=58.055 //y2=0
r1218 (  374 376 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=58.14 //y=0 //x2=59.2 //y2=0
r1219 (  373 534 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.62 //y=0 //x2=61.79 //y2=0
r1220 (  373 380 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=61.62 //y=0 //x2=61.42 //y2=0
r1221 (  369 533 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.055 //y=0.17 //x2=58.055 //y2=0
r1222 (  369 576 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=58.055 //y=0.17 //x2=58.055 //y2=0.965
r1223 (  368 531 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.15 //y=0 //x2=56.98 //y2=0
r1224 (  367 533 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=57.97 //y=0 //x2=58.055 //y2=0
r1225 (  367 368 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=57.97 //y=0 //x2=57.15 //y2=0
r1226 (  362 364 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=55.5 //y=0 //x2=56.61 //y2=0
r1227 (  360 362 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=54.39 //y=0 //x2=55.5 //y2=0
r1228 (  358 530 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.33 //y=0 //x2=53.245 //y2=0
r1229 (  358 360 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=53.33 //y=0 //x2=54.39 //y2=0
r1230 (  357 531 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=56.81 //y=0 //x2=56.98 //y2=0
r1231 (  357 364 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=56.81 //y=0 //x2=56.61 //y2=0
r1232 (  353 530 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=53.245 //y=0.17 //x2=53.245 //y2=0
r1233 (  353 575 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=53.245 //y=0.17 //x2=53.245 //y2=0.965
r1234 (  352 528 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=52.34 //y=0 //x2=52.17 //y2=0
r1235 (  351 530 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.16 //y=0 //x2=53.245 //y2=0
r1236 (  351 352 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=53.16 //y=0 //x2=52.34 //y2=0
r1237 (  346 348 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=50.69 //y=0 //x2=51.8 //y2=0
r1238 (  344 527 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.105 //y=0 //x2=50.02 //y2=0
r1239 (  344 346 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=50.105 //y=0 //x2=50.69 //y2=0
r1240 (  343 528 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=52 //y=0 //x2=52.17 //y2=0
r1241 (  343 348 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=52 //y=0 //x2=51.8 //y2=0
r1242 (  339 527 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=50.02 //y=0.17 //x2=50.02 //y2=0
r1243 (  339 574 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=50.02 //y=0.17 //x2=50.02 //y2=0.955
r1244 (  336 526 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.01 //y=0 //x2=48.84 //y2=0
r1245 (  336 338 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=49.01 //y=0 //x2=49.58 //y2=0
r1246 (  335 527 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.935 //y=0 //x2=50.02 //y2=0
r1247 (  335 338 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=49.935 //y=0 //x2=49.58 //y2=0
r1248 (  330 332 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=46.99 //y=0 //x2=48.1 //y2=0
r1249 (  328 330 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=45.88 //y=0 //x2=46.99 //y2=0
r1250 (  326 525 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.19 //y=0 //x2=45.105 //y2=0
r1251 (  326 328 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=45.19 //y=0 //x2=45.88 //y2=0
r1252 (  325 526 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.67 //y=0 //x2=48.84 //y2=0
r1253 (  325 332 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=48.67 //y=0 //x2=48.1 //y2=0
r1254 (  321 525 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=45.105 //y=0.17 //x2=45.105 //y2=0
r1255 (  321 573 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=45.105 //y=0.17 //x2=45.105 //y2=0.965
r1256 (  318 524 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=44.2 //y=0 //x2=44.03 //y2=0
r1257 (  318 320 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=44.2 //y=0 //x2=44.77 //y2=0
r1258 (  317 525 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.02 //y=0 //x2=45.105 //y2=0
r1259 (  317 320 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=45.02 //y=0 //x2=44.77 //y2=0
r1260 (  312 314 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=42.18 //y=0 //x2=43.29 //y2=0
r1261 (  310 523 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.965 //y=0 //x2=41.88 //y2=0
r1262 (  310 312 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=41.965 //y=0 //x2=42.18 //y2=0
r1263 (  309 524 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.86 //y=0 //x2=44.03 //y2=0
r1264 (  309 314 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=43.86 //y=0 //x2=43.29 //y2=0
r1265 (  305 523 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=41.88 //y=0.17 //x2=41.88 //y2=0
r1266 (  305 572 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=41.88 //y=0.17 //x2=41.88 //y2=0.955
r1267 (  302 522 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.87 //y=0 //x2=40.7 //y2=0
r1268 (  302 304 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=40.87 //y=0 //x2=41.07 //y2=0
r1269 (  301 523 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.795 //y=0 //x2=41.88 //y2=0
r1270 (  301 304 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=41.795 //y=0 //x2=41.07 //y2=0
r1271 (  296 521 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.635 //y=0 //x2=38.55 //y2=0
r1272 (  296 298 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=38.635 //y=0 //x2=39.59 //y2=0
r1273 (  295 522 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.53 //y=0 //x2=40.7 //y2=0
r1274 (  295 298 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=40.53 //y=0 //x2=39.59 //y2=0
r1275 (  291 521 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.55 //y=0.17 //x2=38.55 //y2=0
r1276 (  291 571 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=38.55 //y=0.17 //x2=38.55 //y2=0.955
r1277 (  290 519 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.54 //y=0 //x2=37.37 //y2=0
r1278 (  289 521 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.465 //y=0 //x2=38.55 //y2=0
r1279 (  289 290 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=38.465 //y=0 //x2=37.54 //y2=0
r1280 (  284 286 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=35.89 //y=0 //x2=37 //y2=0
r1281 (  282 284 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=34.78 //y=0 //x2=35.89 //y2=0
r1282 (  280 518 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.72 //y=0 //x2=33.635 //y2=0
r1283 (  280 282 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=33.72 //y=0 //x2=34.78 //y2=0
r1284 (  279 519 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.2 //y=0 //x2=37.37 //y2=0
r1285 (  279 286 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=37.2 //y=0 //x2=37 //y2=0
r1286 (  275 518 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.635 //y=0.17 //x2=33.635 //y2=0
r1287 (  275 570 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=33.635 //y=0.17 //x2=33.635 //y2=0.965
r1288 (  274 516 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.73 //y=0 //x2=32.56 //y2=0
r1289 (  273 518 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.55 //y=0 //x2=33.635 //y2=0
r1290 (  273 274 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=33.55 //y=0 //x2=32.73 //y2=0
r1291 (  268 270 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=31.08 //y=0 //x2=32.19 //y2=0
r1292 (  266 268 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=29.97 //y=0 //x2=31.08 //y2=0
r1293 (  264 515 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.91 //y=0 //x2=28.825 //y2=0
r1294 (  264 266 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=28.91 //y=0 //x2=29.97 //y2=0
r1295 (  263 516 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.39 //y=0 //x2=32.56 //y2=0
r1296 (  263 270 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=32.39 //y=0 //x2=32.19 //y2=0
r1297 (  259 515 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=28.825 //y=0.17 //x2=28.825 //y2=0
r1298 (  259 569 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=28.825 //y=0.17 //x2=28.825 //y2=0.965
r1299 (  258 513 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.92 //y=0 //x2=27.75 //y2=0
r1300 (  257 515 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.74 //y=0 //x2=28.825 //y2=0
r1301 (  257 258 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=28.74 //y=0 //x2=27.92 //y2=0
r1302 (  252 254 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=26.27 //y=0 //x2=27.38 //y2=0
r1303 (  250 512 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.685 //y=0 //x2=25.6 //y2=0
r1304 (  250 252 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=25.685 //y=0 //x2=26.27 //y2=0
r1305 (  249 513 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.58 //y=0 //x2=27.75 //y2=0
r1306 (  249 254 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=27.58 //y=0 //x2=27.38 //y2=0
r1307 (  245 512 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.6 //y=0.17 //x2=25.6 //y2=0
r1308 (  245 568 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=25.6 //y=0.17 //x2=25.6 //y2=0.955
r1309 (  242 511 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.59 //y=0 //x2=24.42 //y2=0
r1310 (  242 244 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.59 //y=0 //x2=25.16 //y2=0
r1311 (  241 512 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.515 //y=0 //x2=25.6 //y2=0
r1312 (  241 244 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=25.515 //y=0 //x2=25.16 //y2=0
r1313 (  236 238 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=22.57 //y=0 //x2=23.68 //y2=0
r1314 (  234 236 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=21.46 //y=0 //x2=22.57 //y2=0
r1315 (  232 510 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.77 //y=0 //x2=20.685 //y2=0
r1316 (  232 234 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=20.77 //y=0 //x2=21.46 //y2=0
r1317 (  231 511 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.25 //y=0 //x2=24.42 //y2=0
r1318 (  231 238 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.25 //y=0 //x2=23.68 //y2=0
r1319 (  227 510 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.685 //y=0.17 //x2=20.685 //y2=0
r1320 (  227 567 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=20.685 //y=0.17 //x2=20.685 //y2=0.965
r1321 (  224 509 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.78 //y=0 //x2=19.61 //y2=0
r1322 (  224 226 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.78 //y=0 //x2=20.35 //y2=0
r1323 (  223 510 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.6 //y=0 //x2=20.685 //y2=0
r1324 (  223 226 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=20.6 //y=0 //x2=20.35 //y2=0
r1325 (  218 220 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=17.76 //y=0 //x2=18.87 //y2=0
r1326 (  216 508 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.545 //y=0 //x2=17.46 //y2=0
r1327 (  216 218 ) resistor r=7.70868 //w=0.357 //l=0.215 //layer=li \
 //thickness=0.1 //x=17.545 //y=0 //x2=17.76 //y2=0
r1328 (  215 509 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.44 //y=0 //x2=19.61 //y2=0
r1329 (  215 220 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.44 //y=0 //x2=18.87 //y2=0
r1330 (  211 508 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.46 //y=0.17 //x2=17.46 //y2=0
r1331 (  211 566 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=17.46 //y=0.17 //x2=17.46 //y2=0.955
r1332 (  208 507 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.45 //y=0 //x2=16.28 //y2=0
r1333 (  208 210 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=16.45 //y=0 //x2=16.65 //y2=0
r1334 (  207 508 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.375 //y=0 //x2=17.46 //y2=0
r1335 (  207 210 ) resistor r=25.9944 //w=0.357 //l=0.725 //layer=li \
 //thickness=0.1 //x=17.375 //y=0 //x2=16.65 //y2=0
r1336 (  202 506 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.215 //y=0 //x2=14.13 //y2=0
r1337 (  202 204 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=14.215 //y=0 //x2=15.17 //y2=0
r1338 (  201 507 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.11 //y=0 //x2=16.28 //y2=0
r1339 (  201 204 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=16.11 //y=0 //x2=15.17 //y2=0
r1340 (  197 506 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.13 //y=0.17 //x2=14.13 //y2=0
r1341 (  197 565 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=14.13 //y=0.17 //x2=14.13 //y2=0.955
r1342 (  196 504 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.12 //y=0 //x2=12.95 //y2=0
r1343 (  195 506 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.045 //y=0 //x2=14.13 //y2=0
r1344 (  195 196 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=14.045 //y=0 //x2=13.12 //y2=0
r1345 (  190 192 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=11.47 //y=0 //x2=12.58 //y2=0
r1346 (  188 190 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=10.36 //y=0 //x2=11.47 //y2=0
r1347 (  186 503 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.3 //y=0 //x2=9.215 //y2=0
r1348 (  186 188 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=9.3 //y=0 //x2=10.36 //y2=0
r1349 (  185 504 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.78 //y=0 //x2=12.95 //y2=0
r1350 (  185 192 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.78 //y=0 //x2=12.58 //y2=0
r1351 (  181 503 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.215 //y=0.17 //x2=9.215 //y2=0
r1352 (  181 564 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=9.215 //y=0.17 //x2=9.215 //y2=0.965
r1353 (  180 501 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=0 //x2=8.14 //y2=0
r1354 (  179 503 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.13 //y=0 //x2=9.215 //y2=0
r1355 (  179 180 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=9.13 //y=0 //x2=8.31 //y2=0
r1356 (  174 176 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r1357 (  172 174 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=5.55 //y=0 //x2=6.66 //y2=0
r1358 (  170 500 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.49 //y=0 //x2=4.405 //y2=0
r1359 (  170 172 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=4.49 //y=0 //x2=5.55 //y2=0
r1360 (  169 501 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=8.14 //y2=0
r1361 (  169 176 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=0 //x2=7.77 //y2=0
r1362 (  165 500 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.405 //y=0.17 //x2=4.405 //y2=0
r1363 (  165 563 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=4.405 //y=0.17 //x2=4.405 //y2=0.965
r1364 (  164 498 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=0 //x2=3.33 //y2=0
r1365 (  163 500 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.32 //y=0 //x2=4.405 //y2=0
r1366 (  163 164 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=4.32 //y=0 //x2=3.5 //y2=0
r1367 (  158 160 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r1368 (  156 497 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.18 //y2=0
r1369 (  156 158 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=1.265 //y=0 //x2=1.85 //y2=0
r1370 (  155 498 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=3.33 //y2=0
r1371 (  155 160 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=2.96 //y2=0
r1372 (  151 497 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r1373 (  151 562 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.955
r1374 (  147 497 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=1.18 //y2=0
r1375 (  147 150 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=1.095 //y=0 //x2=0.74 //y2=0
r1376 (  143 554 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=84.73 //y=0 //x2=84.73 //y2=0
r1377 (  141 551 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=83.99 //y=0 //x2=83.99 //y2=0
r1378 (  141 143 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=83.99 //y=0 //x2=84.73 //y2=0
r1379 (  139 470 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=82.51 //y=0 //x2=82.51 //y2=0
r1380 (  139 141 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=82.51 //y=0 //x2=83.99 //y2=0
r1381 (  137 468 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=81.4 //y=0 //x2=81.4 //y2=0
r1382 (  137 139 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=81.4 //y=0 //x2=82.51 //y2=0
r1383 (  135 460 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=80.29 //y=0 //x2=80.29 //y2=0
r1384 (  135 137 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=80.29 //y=0 //x2=81.4 //y2=0
r1385 (  133 454 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=78.81 //y=0 //x2=78.81 //y2=0
r1386 (  133 135 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=78.81 //y=0 //x2=80.29 //y2=0
r1387 (  131 545 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=77.7 //y=0 //x2=77.7 //y2=0
r1388 (  131 133 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=77.7 //y=0 //x2=78.81 //y2=0
r1389 (  129 442 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=76.22 //y=0 //x2=76.22 //y2=0
r1390 (  129 131 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=76.22 //y=0 //x2=77.7 //y2=0
r1391 (  127 440 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=75.11 //y=0 //x2=75.11 //y2=0
r1392 (  127 129 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=75.11 //y=0 //x2=76.22 //y2=0
r1393 (  125 432 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=74 //y=0 //x2=74 //y2=0
r1394 (  125 127 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=74 //y=0 //x2=75.11 //y2=0
r1395 (  123 426 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=72.52 //y=0 //x2=72.52 //y2=0
r1396 (  123 125 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=72.52 //y=0 //x2=74 //y2=0
r1397 (  121 424 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=71.41 //y=0 //x2=71.41 //y2=0
r1398 (  121 123 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=71.41 //y=0 //x2=72.52 //y2=0
r1399 (  119 422 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=70.3 //y=0 //x2=70.3 //y2=0
r1400 (  119 121 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=70.3 //y=0 //x2=71.41 //y2=0
r1401 (  117 414 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=69.19 //y=0 //x2=69.19 //y2=0
r1402 (  117 119 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=69.19 //y=0 //x2=70.3 //y2=0
r1403 (  115 408 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=67.71 //y=0 //x2=67.71 //y2=0
r1404 (  115 117 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=67.71 //y=0 //x2=69.19 //y2=0
r1405 (  113 406 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=66.6 //y=0 //x2=66.6 //y2=0
r1406 (  113 115 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=66.6 //y=0 //x2=67.71 //y2=0
r1407 (  111 398 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=65.49 //y=0 //x2=65.49 //y2=0
r1408 (  111 113 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=65.49 //y=0 //x2=66.6 //y2=0
r1409 (  109 392 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=64.01 //y=0 //x2=64.01 //y2=0
r1410 (  109 111 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=64.01 //y=0 //x2=65.49 //y2=0
r1411 (  107 536 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=62.9 //y=0 //x2=62.9 //y2=0
r1412 (  107 109 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=62.9 //y=0 //x2=64.01 //y2=0
r1413 (  105 380 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=61.42 //y=0 //x2=61.42 //y2=0
r1414 (  105 107 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=61.42 //y=0 //x2=62.9 //y2=0
r1415 (  103 378 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=60.31 //y=0 //x2=60.31 //y2=0
r1416 (  103 105 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=60.31 //y=0 //x2=61.42 //y2=0
r1417 (  101 376 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=59.2 //y=0 //x2=59.2 //y2=0
r1418 (  101 103 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=59.2 //y=0 //x2=60.31 //y2=0
r1419 (  99 533 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=58.09 //y=0 //x2=58.09 //y2=0
r1420 (  99 101 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=58.09 //y=0 //x2=59.2 //y2=0
r1421 (  97 364 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=56.61 //y=0 //x2=56.61 //y2=0
r1422 (  97 99 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=56.61 //y=0 //x2=58.09 //y2=0
r1423 (  95 362 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=55.5 //y=0 //x2=55.5 //y2=0
r1424 (  95 97 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=55.5 //y=0 //x2=56.61 //y2=0
r1425 (  93 360 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=54.39 //y=0 //x2=54.39 //y2=0
r1426 (  93 95 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=54.39 //y=0 //x2=55.5 //y2=0
r1427 (  91 530 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=53.28 //y=0 //x2=53.28 //y2=0
r1428 (  91 93 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=53.28 //y=0 //x2=54.39 //y2=0
r1429 (  89 348 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=51.8 //y=0 //x2=51.8 //y2=0
r1430 (  89 91 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=51.8 //y=0 //x2=53.28 //y2=0
r1431 (  87 346 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=50.69 //y=0 //x2=50.69 //y2=0
r1432 (  87 89 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=50.69 //y=0 //x2=51.8 //y2=0
r1433 (  85 338 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=49.58 //y=0 //x2=49.58 //y2=0
r1434 (  85 87 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=49.58 //y=0 //x2=50.69 //y2=0
r1435 (  83 332 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=48.1 //y=0 //x2=48.1 //y2=0
r1436 (  83 85 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=48.1 //y=0 //x2=49.58 //y2=0
r1437 (  81 330 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=46.99 //y=0 //x2=46.99 //y2=0
r1438 (  81 83 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=46.99 //y=0 //x2=48.1 //y2=0
r1439 (  79 328 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=45.88 //y=0 //x2=45.88 //y2=0
r1440 (  79 81 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=45.88 //y=0 //x2=46.99 //y2=0
r1441 (  77 320 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=44.77 //y=0 //x2=44.77 //y2=0
r1442 (  77 79 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=44.77 //y=0 //x2=45.88 //y2=0
r1443 (  75 314 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=43.29 //y=0 //x2=43.29 //y2=0
r1444 (  75 77 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=43.29 //y=0 //x2=44.77 //y2=0
r1445 (  72 312 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=42.18 //y=0 //x2=42.18 //y2=0
r1446 (  70 304 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=41.07 //y=0 //x2=41.07 //y2=0
r1447 (  70 72 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=41.07 //y=0 //x2=42.18 //y2=0
r1448 (  68 298 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=39.59 //y=0 //x2=39.59 //y2=0
r1449 (  68 70 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=39.59 //y=0 //x2=41.07 //y2=0
r1450 (  66 521 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=38.48 //y=0 //x2=38.48 //y2=0
r1451 (  66 68 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=38.48 //y=0 //x2=39.59 //y2=0
r1452 (  64 286 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37 //y=0 //x2=37 //y2=0
r1453 (  64 66 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=37 //y=0 //x2=38.48 //y2=0
r1454 (  62 284 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.89 //y=0 //x2=35.89 //y2=0
r1455 (  62 64 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=35.89 //y=0 //x2=37 //y2=0
r1456 (  60 282 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.78 //y=0 //x2=34.78 //y2=0
r1457 (  60 62 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=34.78 //y=0 //x2=35.89 //y2=0
r1458 (  58 518 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=33.67 //y=0 //x2=33.67 //y2=0
r1459 (  58 60 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=33.67 //y=0 //x2=34.78 //y2=0
r1460 (  56 270 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.19 //y=0 //x2=32.19 //y2=0
r1461 (  56 58 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=32.19 //y=0 //x2=33.67 //y2=0
r1462 (  54 268 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.08 //y=0 //x2=31.08 //y2=0
r1463 (  54 56 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.08 //y=0 //x2=32.19 //y2=0
r1464 (  52 266 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=29.97 //y=0 //x2=29.97 //y2=0
r1465 (  52 54 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=29.97 //y=0 //x2=31.08 //y2=0
r1466 (  50 515 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.86 //y=0 //x2=28.86 //y2=0
r1467 (  50 52 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=28.86 //y=0 //x2=29.97 //y2=0
r1468 (  48 254 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.38 //y=0 //x2=27.38 //y2=0
r1469 (  48 50 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=27.38 //y=0 //x2=28.86 //y2=0
r1470 (  46 252 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=26.27 //y=0 //x2=26.27 //y2=0
r1471 (  46 48 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=26.27 //y=0 //x2=27.38 //y2=0
r1472 (  44 244 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.16 //y=0 //x2=25.16 //y2=0
r1473 (  44 46 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=25.16 //y=0 //x2=26.27 //y2=0
r1474 (  42 238 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=0 //x2=23.68 //y2=0
r1475 (  42 44 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=23.68 //y=0 //x2=25.16 //y2=0
r1476 (  40 236 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.57 //y=0 //x2=22.57 //y2=0
r1477 (  40 42 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.57 //y=0 //x2=23.68 //y2=0
r1478 (  38 234 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.46 //y=0 //x2=21.46 //y2=0
r1479 (  38 40 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.46 //y=0 //x2=22.57 //y2=0
r1480 (  36 226 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=0 //x2=20.35 //y2=0
r1481 (  36 38 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=0 //x2=21.46 //y2=0
r1482 (  34 220 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.87 //y=0 //x2=18.87 //y2=0
r1483 (  34 36 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.87 //y=0 //x2=20.35 //y2=0
r1484 (  32 218 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=0 //x2=17.76 //y2=0
r1485 (  32 34 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=0 //x2=18.87 //y2=0
r1486 (  30 210 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=0 //x2=16.65 //y2=0
r1487 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=0 //x2=17.76 //y2=0
r1488 (  28 204 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=0 //x2=15.17 //y2=0
r1489 (  28 30 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=0 //x2=16.65 //y2=0
r1490 (  26 506 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=0 //x2=14.06 //y2=0
r1491 (  26 28 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=0 //x2=15.17 //y2=0
r1492 (  24 192 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=0 //x2=12.58 //y2=0
r1493 (  24 26 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=0 //x2=14.06 //y2=0
r1494 (  22 190 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=0 //x2=11.47 //y2=0
r1495 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=0 //x2=12.58 //y2=0
r1496 (  20 188 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r1497 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=0 //x2=11.47 //y2=0
r1498 (  18 503 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=0 //x2=9.25 //y2=0
r1499 (  18 20 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=0 //x2=10.36 //y2=0
r1500 (  16 176 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r1501 (  16 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=9.25 //y2=0
r1502 (  14 174 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r1503 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r1504 (  12 172 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r1505 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r1506 (  10 500 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r1507 (  10 12 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.55 //y2=0
r1508 (  8 160 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r1509 (  8 10 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.44 //y2=0
r1510 (  6 158 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r1511 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r1512 (  3 150 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r1513 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r1514 (  1 75 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=42.735 //y=0 //x2=43.29 //y2=0
r1515 (  1 72 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=42.735 //y=0 //x2=42.18 //y2=0
ends PM_TMRDFFSNQX1\%GND

subckt PM_TMRDFFSNQX1\%VDD ( 1 143 155 163 173 179 187 195 205 215 221 229 237 \
 247 257 263 271 281 291 295 305 315 323 327 337 347 355 365 371 379 387 397 \
 403 411 419 429 439 445 453 461 471 481 487 495 505 515 519 529 539 547 551 \
 561 571 579 589 595 603 611 621 627 635 643 653 663 669 677 685 695 705 711 \
 719 729 739 743 753 763 771 775 785 795 803 813 819 827 835 845 851 859 869 \
 877 890 893 899 905 909 914 919 924 930 936 940 945 950 955 961 967 971 976 \
 981 986 987 988 992 993 994 995 996 997 998 999 1000 1001 1002 1003 1004 1005 \
 1006 1007 1008 1009 1010 1011 1012 1013 1014 1015 1016 1017 1018 1019 1020 \
 1021 1022 1023 1024 1025 1026 1027 1028 1029 1030 1031 1032 1033 1034 1035 \
 1036 1037 1038 1039 1040 1041 1042 1043 1044 1045 1046 1047 1048 1049 1050 \
 1051 1052 1053 1054 1055 1056 1057 1058 1059 1060 )
c1105 ( 1060 0 ) capacitor c=0.0451925f //x=84.66 //y=5.02
c1106 ( 1059 0 ) capacitor c=0.0420333f //x=83.79 //y=5.02
c1107 ( 1058 0 ) capacitor c=0.0476806f //x=75.665 //y=5.025
c1108 ( 1057 0 ) capacitor c=0.0241714f //x=74.785 //y=5.025
c1109 ( 1056 0 ) capacitor c=0.0467094f //x=73.915 //y=5.025
c1110 ( 1055 0 ) capacitor c=0.0452179f //x=72.035 //y=5.02
c1111 ( 1054 0 ) capacitor c=0.024152f //x=71.155 //y=5.02
c1112 ( 1053 0 ) capacitor c=0.024152f //x=70.275 //y=5.02
c1113 ( 1052 0 ) capacitor c=0.0530764f //x=69.405 //y=5.02
c1114 ( 1051 0 ) capacitor c=0.0379509f //x=67.525 //y=5.02
c1115 ( 1050 0 ) capacitor c=0.0241088f //x=66.645 //y=5.02
c1116 ( 1049 0 ) capacitor c=0.0493657f //x=65.775 //y=5.02
c1117 ( 1048 0 ) capacitor c=0.0381505f //x=64.195 //y=5.02
c1118 ( 1047 0 ) capacitor c=0.0240074f //x=63.315 //y=5.02
c1119 ( 1046 0 ) capacitor c=0.049209f //x=62.445 //y=5.02
c1120 ( 1045 0 ) capacitor c=0.0452179f //x=60.565 //y=5.02
c1121 ( 1044 0 ) capacitor c=0.024152f //x=59.685 //y=5.02
c1122 ( 1043 0 ) capacitor c=0.024152f //x=58.805 //y=5.02
c1123 ( 1042 0 ) capacitor c=0.053132f //x=57.935 //y=5.02
c1124 ( 1041 0 ) capacitor c=0.0452179f //x=55.755 //y=5.02
c1125 ( 1040 0 ) capacitor c=0.024152f //x=54.875 //y=5.02
c1126 ( 1039 0 ) capacitor c=0.024152f //x=53.995 //y=5.02
c1127 ( 1038 0 ) capacitor c=0.0531894f //x=53.125 //y=5.02
c1128 ( 1037 0 ) capacitor c=0.0380679f //x=51.245 //y=5.02
c1129 ( 1036 0 ) capacitor c=0.024008f //x=50.365 //y=5.02
c1130 ( 1035 0 ) capacitor c=0.049209f //x=49.495 //y=5.02
c1131 ( 1034 0 ) capacitor c=0.0452179f //x=47.615 //y=5.02
c1132 ( 1033 0 ) capacitor c=0.024152f //x=46.735 //y=5.02
c1133 ( 1032 0 ) capacitor c=0.024152f //x=45.855 //y=5.02
c1134 ( 1031 0 ) capacitor c=0.0531894f //x=44.985 //y=5.02
c1135 ( 1030 0 ) capacitor c=0.0380679f //x=43.105 //y=5.02
c1136 ( 1029 0 ) capacitor c=0.024008f //x=42.225 //y=5.02
c1137 ( 1028 0 ) capacitor c=0.0490303f //x=41.355 //y=5.02
c1138 ( 1027 0 ) capacitor c=0.0380679f //x=39.775 //y=5.02
c1139 ( 1026 0 ) capacitor c=0.0240074f //x=38.895 //y=5.02
c1140 ( 1025 0 ) capacitor c=0.049209f //x=38.025 //y=5.02
c1141 ( 1024 0 ) capacitor c=0.0452179f //x=36.145 //y=5.02
c1142 ( 1023 0 ) capacitor c=0.024152f //x=35.265 //y=5.02
c1143 ( 1022 0 ) capacitor c=0.024152f //x=34.385 //y=5.02
c1144 ( 1021 0 ) capacitor c=0.053132f //x=33.515 //y=5.02
c1145 ( 1020 0 ) capacitor c=0.0452179f //x=31.335 //y=5.02
c1146 ( 1019 0 ) capacitor c=0.024152f //x=30.455 //y=5.02
c1147 ( 1018 0 ) capacitor c=0.024152f //x=29.575 //y=5.02
c1148 ( 1017 0 ) capacitor c=0.0531894f //x=28.705 //y=5.02
c1149 ( 1016 0 ) capacitor c=0.0380679f //x=26.825 //y=5.02
c1150 ( 1015 0 ) capacitor c=0.024008f //x=25.945 //y=5.02
c1151 ( 1014 0 ) capacitor c=0.049209f //x=25.075 //y=5.02
c1152 ( 1013 0 ) capacitor c=0.0452179f //x=23.195 //y=5.02
c1153 ( 1012 0 ) capacitor c=0.024152f //x=22.315 //y=5.02
c1154 ( 1011 0 ) capacitor c=0.024152f //x=21.435 //y=5.02
c1155 ( 1010 0 ) capacitor c=0.0531894f //x=20.565 //y=5.02
c1156 ( 1009 0 ) capacitor c=0.0380679f //x=18.685 //y=5.02
c1157 ( 1008 0 ) capacitor c=0.024008f //x=17.805 //y=5.02
c1158 ( 1007 0 ) capacitor c=0.0490303f //x=16.935 //y=5.02
c1159 ( 1006 0 ) capacitor c=0.0380679f //x=15.355 //y=5.02
c1160 ( 1005 0 ) capacitor c=0.0240074f //x=14.475 //y=5.02
c1161 ( 1004 0 ) capacitor c=0.049209f //x=13.605 //y=5.02
c1162 ( 1003 0 ) capacitor c=0.0452179f //x=11.725 //y=5.02
c1163 ( 1002 0 ) capacitor c=0.024152f //x=10.845 //y=5.02
c1164 ( 1001 0 ) capacitor c=0.024152f //x=9.965 //y=5.02
c1165 ( 1000 0 ) capacitor c=0.053132f //x=9.095 //y=5.02
c1166 ( 999 0 ) capacitor c=0.0452179f //x=6.915 //y=5.02
c1167 ( 998 0 ) capacitor c=0.024152f //x=6.035 //y=5.02
c1168 ( 997 0 ) capacitor c=0.02424f //x=5.155 //y=5.02
c1169 ( 996 0 ) capacitor c=0.0532367f //x=4.285 //y=5.02
c1170 ( 995 0 ) capacitor c=0.0381505f //x=2.405 //y=5.02
c1171 ( 994 0 ) capacitor c=0.0241853f //x=1.525 //y=5.02
c1172 ( 993 0 ) capacitor c=0.053196f //x=0.655 //y=5.02
c1173 ( 992 0 ) capacitor c=0.234643f //x=84.73 //y=7.4
c1174 ( 990 0 ) capacitor c=0.00591168f //x=83.99 //y=7.4
c1175 ( 988 0 ) capacitor c=0.107657f //x=83.25 //y=7.4
c1176 ( 987 0 ) capacitor c=0.113329f //x=79.92 //y=7.4
c1177 ( 986 0 ) capacitor c=0.121062f //x=76.59 //y=7.4
c1178 ( 985 0 ) capacitor c=0.00591168f //x=75.81 //y=7.4
c1179 ( 984 0 ) capacitor c=0.00591168f //x=74.93 //y=7.4
c1180 ( 983 0 ) capacitor c=0.00591168f //x=74 //y=7.4
c1181 ( 981 0 ) capacitor c=0.13666f //x=73.26 //y=7.4
c1182 ( 980 0 ) capacitor c=0.00591168f //x=72.18 //y=7.4
c1183 ( 979 0 ) capacitor c=0.00591168f //x=71.3 //y=7.4
c1184 ( 978 0 ) capacitor c=0.00591168f //x=70.42 //y=7.4
c1185 ( 977 0 ) capacitor c=0.00591168f //x=69.54 //y=7.4
c1186 ( 976 0 ) capacitor c=0.137467f //x=68.45 //y=7.4
c1187 ( 975 0 ) capacitor c=0.00591168f //x=67.71 //y=7.4
c1188 ( 973 0 ) capacitor c=0.00591168f //x=66.79 //y=7.4
c1189 ( 972 0 ) capacitor c=0.00591168f //x=65.91 //y=7.4
c1190 ( 971 0 ) capacitor c=0.115594f //x=65.12 //y=7.4
c1191 ( 970 0 ) capacitor c=0.00591168f //x=64.34 //y=7.4
c1192 ( 969 0 ) capacitor c=0.00591168f //x=63.46 //y=7.4
c1193 ( 968 0 ) capacitor c=0.00591168f //x=62.58 //y=7.4
c1194 ( 967 0 ) capacitor c=0.13452f //x=61.79 //y=7.4
c1195 ( 966 0 ) capacitor c=0.00591168f //x=60.71 //y=7.4
c1196 ( 965 0 ) capacitor c=0.00591168f //x=59.83 //y=7.4
c1197 ( 964 0 ) capacitor c=0.00591168f //x=58.95 //y=7.4
c1198 ( 963 0 ) capacitor c=0.00591168f //x=58.09 //y=7.4
c1199 ( 961 0 ) capacitor c=0.155082f //x=56.98 //y=7.4
c1200 ( 960 0 ) capacitor c=0.00591168f //x=55.9 //y=7.4
c1201 ( 959 0 ) capacitor c=0.00591168f //x=55.02 //y=7.4
c1202 ( 958 0 ) capacitor c=0.00591168f //x=54.14 //y=7.4
c1203 ( 957 0 ) capacitor c=0.00591168f //x=53.28 //y=7.4
c1204 ( 955 0 ) capacitor c=0.135216f //x=52.17 //y=7.4
c1205 ( 954 0 ) capacitor c=0.00591168f //x=51.39 //y=7.4
c1206 ( 953 0 ) capacitor c=0.00591168f //x=50.51 //y=7.4
c1207 ( 952 0 ) capacitor c=0.00591168f //x=49.58 //y=7.4
c1208 ( 950 0 ) capacitor c=0.138747f //x=48.84 //y=7.4
c1209 ( 949 0 ) capacitor c=0.00591168f //x=47.76 //y=7.4
c1210 ( 948 0 ) capacitor c=0.00591168f //x=46.88 //y=7.4
c1211 ( 947 0 ) capacitor c=0.00591168f //x=46 //y=7.4
c1212 ( 946 0 ) capacitor c=0.00591168f //x=45.12 //y=7.4
c1213 ( 945 0 ) capacitor c=0.135109f //x=44.03 //y=7.4
c1214 ( 944 0 ) capacitor c=0.00591168f //x=43.29 //y=7.4
c1215 ( 942 0 ) capacitor c=0.00591168f //x=42.37 //y=7.4
c1216 ( 941 0 ) capacitor c=0.00591168f //x=41.49 //y=7.4
c1217 ( 940 0 ) capacitor c=0.11432f //x=40.7 //y=7.4
c1218 ( 939 0 ) capacitor c=0.00591168f //x=39.92 //y=7.4
c1219 ( 938 0 ) capacitor c=0.00591168f //x=39.04 //y=7.4
c1220 ( 937 0 ) capacitor c=0.00591168f //x=38.16 //y=7.4
c1221 ( 936 0 ) capacitor c=0.13452f //x=37.37 //y=7.4
c1222 ( 935 0 ) capacitor c=0.00591168f //x=36.29 //y=7.4
c1223 ( 934 0 ) capacitor c=0.00591168f //x=35.41 //y=7.4
c1224 ( 933 0 ) capacitor c=0.00591168f //x=34.53 //y=7.4
c1225 ( 932 0 ) capacitor c=0.00591168f //x=33.67 //y=7.4
c1226 ( 930 0 ) capacitor c=0.155082f //x=32.56 //y=7.4
c1227 ( 929 0 ) capacitor c=0.00591168f //x=31.48 //y=7.4
c1228 ( 928 0 ) capacitor c=0.00591168f //x=30.6 //y=7.4
c1229 ( 927 0 ) capacitor c=0.00591168f //x=29.72 //y=7.4
c1230 ( 926 0 ) capacitor c=0.00591168f //x=28.86 //y=7.4
c1231 ( 924 0 ) capacitor c=0.135216f //x=27.75 //y=7.4
c1232 ( 923 0 ) capacitor c=0.00591168f //x=26.97 //y=7.4
c1233 ( 922 0 ) capacitor c=0.00591168f //x=26.09 //y=7.4
c1234 ( 921 0 ) capacitor c=0.00591168f //x=25.16 //y=7.4
c1235 ( 919 0 ) capacitor c=0.139023f //x=24.42 //y=7.4
c1236 ( 918 0 ) capacitor c=0.00591168f //x=23.34 //y=7.4
c1237 ( 917 0 ) capacitor c=0.00591168f //x=22.46 //y=7.4
c1238 ( 916 0 ) capacitor c=0.00591168f //x=21.58 //y=7.4
c1239 ( 915 0 ) capacitor c=0.00591168f //x=20.7 //y=7.4
c1240 ( 914 0 ) capacitor c=0.134951f //x=19.61 //y=7.4
c1241 ( 913 0 ) capacitor c=0.00591168f //x=18.87 //y=7.4
c1242 ( 911 0 ) capacitor c=0.00591168f //x=17.95 //y=7.4
c1243 ( 910 0 ) capacitor c=0.00591168f //x=17.07 //y=7.4
c1244 ( 909 0 ) capacitor c=0.11432f //x=16.28 //y=7.4
c1245 ( 908 0 ) capacitor c=0.00591168f //x=15.5 //y=7.4
c1246 ( 907 0 ) capacitor c=0.00591168f //x=14.62 //y=7.4
c1247 ( 906 0 ) capacitor c=0.00591168f //x=13.74 //y=7.4
c1248 ( 905 0 ) capacitor c=0.13452f //x=12.95 //y=7.4
c1249 ( 904 0 ) capacitor c=0.00591168f //x=11.87 //y=7.4
c1250 ( 903 0 ) capacitor c=0.00591168f //x=10.99 //y=7.4
c1251 ( 902 0 ) capacitor c=0.00591168f //x=10.11 //y=7.4
c1252 ( 901 0 ) capacitor c=0.00591168f //x=9.25 //y=7.4
c1253 ( 899 0 ) capacitor c=0.155082f //x=8.14 //y=7.4
c1254 ( 898 0 ) capacitor c=0.00591168f //x=7.06 //y=7.4
c1255 ( 897 0 ) capacitor c=0.00591168f //x=6.18 //y=7.4
c1256 ( 896 0 ) capacitor c=0.00591168f //x=5.3 //y=7.4
c1257 ( 895 0 ) capacitor c=0.00591168f //x=4.44 //y=7.4
c1258 ( 893 0 ) capacitor c=0.137297f //x=3.33 //y=7.4
c1259 ( 892 0 ) capacitor c=0.00591168f //x=2.55 //y=7.4
c1260 ( 891 0 ) capacitor c=0.00591168f //x=1.67 //y=7.4
c1261 ( 890 0 ) capacitor c=0.248311f //x=0.74 //y=7.4
c1262 ( 877 0 ) capacitor c=0.0287851f //x=84.72 //y=7.4
c1263 ( 869 0 ) capacitor c=0.0186283f //x=83.84 //y=7.4
c1264 ( 859 0 ) capacitor c=0.12108f //x=83.08 //y=7.4
c1265 ( 851 0 ) capacitor c=0.120978f //x=79.75 //y=7.4
c1266 ( 845 0 ) capacitor c=0.0236224f //x=76.42 //y=7.4
c1267 ( 835 0 ) capacitor c=0.028539f //x=75.725 //y=7.4
c1268 ( 827 0 ) capacitor c=0.0285075f //x=74.845 //y=7.4
c1269 ( 819 0 ) capacitor c=0.0240981f //x=73.965 //y=7.4
c1270 ( 813 0 ) capacitor c=0.0394633f //x=73.09 //y=7.4
c1271 ( 803 0 ) capacitor c=0.0288488f //x=72.095 //y=7.4
c1272 ( 795 0 ) capacitor c=0.0287514f //x=71.215 //y=7.4
c1273 ( 785 0 ) capacitor c=0.0284966f //x=70.335 //y=7.4
c1274 ( 775 0 ) capacitor c=0.0383672f //x=69.455 //y=7.4
c1275 ( 771 0 ) capacitor c=0.0237444f //x=68.28 //y=7.4
c1276 ( 763 0 ) capacitor c=0.0288357f //x=67.585 //y=7.4
c1277 ( 753 0 ) capacitor c=0.0291038f //x=66.705 //y=7.4
c1278 ( 743 0 ) capacitor c=0.0240981f //x=65.825 //y=7.4
c1279 ( 739 0 ) capacitor c=0.0236224f //x=64.95 //y=7.4
c1280 ( 729 0 ) capacitor c=0.0288598f //x=64.255 //y=7.4
c1281 ( 719 0 ) capacitor c=0.0288369f //x=63.375 //y=7.4
c1282 ( 711 0 ) capacitor c=0.0240981f //x=62.495 //y=7.4
c1283 ( 705 0 ) capacitor c=0.0394667f //x=61.62 //y=7.4
c1284 ( 695 0 ) capacitor c=0.0288488f //x=60.625 //y=7.4
c1285 ( 685 0 ) capacitor c=0.0287514f //x=59.745 //y=7.4
c1286 ( 677 0 ) capacitor c=0.0284966f //x=58.865 //y=7.4
c1287 ( 669 0 ) capacitor c=0.0383672f //x=57.985 //y=7.4
c1288 ( 663 0 ) capacitor c=0.0394667f //x=56.81 //y=7.4
c1289 ( 653 0 ) capacitor c=0.0288488f //x=55.815 //y=7.4
c1290 ( 643 0 ) capacitor c=0.0287505f //x=54.935 //y=7.4
c1291 ( 635 0 ) capacitor c=0.0284966f //x=54.055 //y=7.4
c1292 ( 627 0 ) capacitor c=0.0383672f //x=53.175 //y=7.4
c1293 ( 621 0 ) capacitor c=0.0236224f //x=52 //y=7.4
c1294 ( 611 0 ) capacitor c=0.0288359f //x=51.305 //y=7.4
c1295 ( 603 0 ) capacitor c=0.0288369f //x=50.425 //y=7.4
c1296 ( 595 0 ) capacitor c=0.0240981f //x=49.545 //y=7.4
c1297 ( 589 0 ) capacitor c=0.0394667f //x=48.67 //y=7.4
c1298 ( 579 0 ) capacitor c=0.0288488f //x=47.675 //y=7.4
c1299 ( 571 0 ) capacitor c=0.0287514f //x=46.795 //y=7.4
c1300 ( 561 0 ) capacitor c=0.0284966f //x=45.915 //y=7.4
c1301 ( 551 0 ) capacitor c=0.0383672f //x=45.035 //y=7.4
c1302 ( 547 0 ) capacitor c=0.0236224f //x=43.86 //y=7.4
c1303 ( 539 0 ) capacitor c=0.0288359f //x=43.165 //y=7.4
c1304 ( 529 0 ) capacitor c=0.0288369f //x=42.285 //y=7.4
c1305 ( 519 0 ) capacitor c=0.0240981f //x=41.405 //y=7.4
c1306 ( 515 0 ) capacitor c=0.0236224f //x=40.53 //y=7.4
c1307 ( 505 0 ) capacitor c=0.0288357f //x=39.835 //y=7.4
c1308 ( 495 0 ) capacitor c=0.0288369f //x=38.955 //y=7.4
c1309 ( 487 0 ) capacitor c=0.0240981f //x=38.075 //y=7.4
c1310 ( 481 0 ) capacitor c=0.0394667f //x=37.2 //y=7.4
c1311 ( 471 0 ) capacitor c=0.0288488f //x=36.205 //y=7.4
c1312 ( 461 0 ) capacitor c=0.0287514f //x=35.325 //y=7.4
c1313 ( 453 0 ) capacitor c=0.0284966f //x=34.445 //y=7.4
c1314 ( 445 0 ) capacitor c=0.0383672f //x=33.565 //y=7.4
c1315 ( 439 0 ) capacitor c=0.0394667f //x=32.39 //y=7.4
c1316 ( 429 0 ) capacitor c=0.0288488f //x=31.395 //y=7.4
c1317 ( 419 0 ) capacitor c=0.0287505f //x=30.515 //y=7.4
c1318 ( 411 0 ) capacitor c=0.0284966f //x=29.635 //y=7.4
c1319 ( 403 0 ) capacitor c=0.0383672f //x=28.755 //y=7.4
c1320 ( 397 0 ) capacitor c=0.0236224f //x=27.58 //y=7.4
c1321 ( 387 0 ) capacitor c=0.0288359f //x=26.885 //y=7.4
c1322 ( 379 0 ) capacitor c=0.0288369f //x=26.005 //y=7.4
c1323 ( 371 0 ) capacitor c=0.0240981f //x=25.125 //y=7.4
c1324 ( 365 0 ) capacitor c=0.0394667f //x=24.25 //y=7.4
c1325 ( 355 0 ) capacitor c=0.0288488f //x=23.255 //y=7.4
c1326 ( 347 0 ) capacitor c=0.0287514f //x=22.375 //y=7.4
c1327 ( 337 0 ) capacitor c=0.0284966f //x=21.495 //y=7.4
c1328 ( 327 0 ) capacitor c=0.0383672f //x=20.615 //y=7.4
c1329 ( 323 0 ) capacitor c=0.0236224f //x=19.44 //y=7.4
c1330 ( 315 0 ) capacitor c=0.0288359f //x=18.745 //y=7.4
c1331 ( 305 0 ) capacitor c=0.0288369f //x=17.865 //y=7.4
c1332 ( 295 0 ) capacitor c=0.0240981f //x=16.985 //y=7.4
c1333 ( 291 0 ) capacitor c=0.0236224f //x=16.11 //y=7.4
c1334 ( 281 0 ) capacitor c=0.0288357f //x=15.415 //y=7.4
c1335 ( 271 0 ) capacitor c=0.0288369f //x=14.535 //y=7.4
c1336 ( 263 0 ) capacitor c=0.0240981f //x=13.655 //y=7.4
c1337 ( 257 0 ) capacitor c=0.0394667f //x=12.78 //y=7.4
c1338 ( 247 0 ) capacitor c=0.0288488f //x=11.785 //y=7.4
c1339 ( 237 0 ) capacitor c=0.0287514f //x=10.905 //y=7.4
c1340 ( 229 0 ) capacitor c=0.0284966f //x=10.025 //y=7.4
c1341 ( 221 0 ) capacitor c=0.0383672f //x=9.145 //y=7.4
c1342 ( 215 0 ) capacitor c=0.0394667f //x=7.97 //y=7.4
c1343 ( 205 0 ) capacitor c=0.0288488f //x=6.975 //y=7.4
c1344 ( 195 0 ) capacitor c=0.0287505f //x=6.095 //y=7.4
c1345 ( 187 0 ) capacitor c=0.028511f //x=5.215 //y=7.4
c1346 ( 179 0 ) capacitor c=0.0383672f //x=4.335 //y=7.4
c1347 ( 173 0 ) capacitor c=0.0236224f //x=3.16 //y=7.4
c1348 ( 163 0 ) capacitor c=0.0288637f //x=2.465 //y=7.4
c1349 ( 155 0 ) capacitor c=0.0286367f //x=1.585 //y=7.4
c1350 ( 143 0 ) capacitor c=2.81857f //x=84.73 //y=7.4
r1351 (  879 992 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=84.805 //y=7.23 //x2=84.805 //y2=7.4
r1352 (  879 1060 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=84.805 //y=7.23 //x2=84.805 //y2=6.405
r1353 (  878 990 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.01 //y=7.4 //x2=83.925 //y2=7.4
r1354 (  877 992 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=84.72 //y=7.4 //x2=84.805 //y2=7.4
r1355 (  877 878 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=84.72 //y=7.4 //x2=84.01 //y2=7.4
r1356 (  871 990 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=83.925 //y=7.23 //x2=83.925 //y2=7.4
r1357 (  871 1059 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=83.925 //y=7.23 //x2=83.925 //y2=6.405
r1358 (  870 988 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=83.42 //y=7.4 //x2=83.25 //y2=7.4
r1359 (  869 990 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=83.84 //y=7.4 //x2=83.925 //y2=7.4
r1360 (  869 870 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=83.84 //y=7.4 //x2=83.42 //y2=7.4
r1361 (  864 866 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=81.4 //y=7.4 //x2=82.51 //y2=7.4
r1362 (  862 864 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=80.29 //y=7.4 //x2=81.4 //y2=7.4
r1363 (  860 987 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=80.09 //y=7.4 //x2=79.92 //y2=7.4
r1364 (  860 862 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=80.09 //y=7.4 //x2=80.29 //y2=7.4
r1365 (  859 988 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=83.08 //y=7.4 //x2=83.25 //y2=7.4
r1366 (  859 866 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=83.08 //y=7.4 //x2=82.51 //y2=7.4
r1367 (  854 856 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=77.7 //y=7.4 //x2=78.81 //y2=7.4
r1368 (  852 986 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.76 //y=7.4 //x2=76.59 //y2=7.4
r1369 (  852 854 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=76.76 //y=7.4 //x2=77.7 //y2=7.4
r1370 (  851 987 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=79.75 //y=7.4 //x2=79.92 //y2=7.4
r1371 (  851 856 ) resistor r=33.7031 //w=0.357 //l=0.94 //layer=li \
 //thickness=0.1 //x=79.75 //y=7.4 //x2=78.81 //y2=7.4
r1372 (  846 985 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.895 //y=7.4 //x2=75.81 //y2=7.4
r1373 (  846 848 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=75.895 //y=7.4 //x2=76.22 //y2=7.4
r1374 (  845 986 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=76.42 //y=7.4 //x2=76.59 //y2=7.4
r1375 (  845 848 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=76.42 //y=7.4 //x2=76.22 //y2=7.4
r1376 (  839 985 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=75.81 //y=7.23 //x2=75.81 //y2=7.4
r1377 (  839 1058 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=75.81 //y=7.23 //x2=75.81 //y2=6.4
r1378 (  836 984 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.015 //y=7.4 //x2=74.93 //y2=7.4
r1379 (  836 838 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=75.015 //y=7.4 //x2=75.11 //y2=7.4
r1380 (  835 985 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=75.725 //y=7.4 //x2=75.81 //y2=7.4
r1381 (  835 838 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=75.725 //y=7.4 //x2=75.11 //y2=7.4
r1382 (  829 984 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=74.93 //y=7.23 //x2=74.93 //y2=7.4
r1383 (  829 1057 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=74.93 //y=7.23 //x2=74.93 //y2=6.74
r1384 (  828 983 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.135 //y=7.4 //x2=74.05 //y2=7.4
r1385 (  827 984 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=74.845 //y=7.4 //x2=74.93 //y2=7.4
r1386 (  827 828 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=74.845 //y=7.4 //x2=74.135 //y2=7.4
r1387 (  821 983 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=74.05 //y=7.23 //x2=74.05 //y2=7.4
r1388 (  821 1056 ) resistor r=56.8128 //w=0.187 //l=0.83 //layer=li \
 //thickness=0.1 //x=74.05 //y=7.23 //x2=74.05 //y2=6.4
r1389 (  820 981 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.43 //y=7.4 //x2=73.26 //y2=7.4
r1390 (  819 983 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=73.965 //y=7.4 //x2=74.05 //y2=7.4
r1391 (  819 820 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=73.965 //y=7.4 //x2=73.43 //y2=7.4
r1392 (  814 980 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.265 //y=7.4 //x2=72.18 //y2=7.4
r1393 (  814 816 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=72.265 //y=7.4 //x2=72.52 //y2=7.4
r1394 (  813 981 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=73.09 //y=7.4 //x2=73.26 //y2=7.4
r1395 (  813 816 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=73.09 //y=7.4 //x2=72.52 //y2=7.4
r1396 (  807 980 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=72.18 //y=7.23 //x2=72.18 //y2=7.4
r1397 (  807 1055 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=72.18 //y=7.23 //x2=72.18 //y2=6.745
r1398 (  804 979 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.385 //y=7.4 //x2=71.3 //y2=7.4
r1399 (  804 806 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=71.385 //y=7.4 //x2=71.41 //y2=7.4
r1400 (  803 980 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=72.095 //y=7.4 //x2=72.18 //y2=7.4
r1401 (  803 806 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=72.095 //y=7.4 //x2=71.41 //y2=7.4
r1402 (  797 979 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=71.3 //y=7.23 //x2=71.3 //y2=7.4
r1403 (  797 1054 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=71.3 //y=7.23 //x2=71.3 //y2=6.745
r1404 (  796 978 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.505 //y=7.4 //x2=70.42 //y2=7.4
r1405 (  795 979 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.215 //y=7.4 //x2=71.3 //y2=7.4
r1406 (  795 796 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=71.215 //y=7.4 //x2=70.505 //y2=7.4
r1407 (  789 978 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=70.42 //y=7.23 //x2=70.42 //y2=7.4
r1408 (  789 1053 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=70.42 //y=7.23 //x2=70.42 //y2=6.745
r1409 (  786 977 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.625 //y=7.4 //x2=69.54 //y2=7.4
r1410 (  786 788 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=69.625 //y=7.4 //x2=70.3 //y2=7.4
r1411 (  785 978 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.335 //y=7.4 //x2=70.42 //y2=7.4
r1412 (  785 788 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=70.335 //y=7.4 //x2=70.3 //y2=7.4
r1413 (  779 977 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=69.54 //y=7.23 //x2=69.54 //y2=7.4
r1414 (  779 1052 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=69.54 //y=7.23 //x2=69.54 //y2=6.405
r1415 (  776 976 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.62 //y=7.4 //x2=68.45 //y2=7.4
r1416 (  776 778 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=68.62 //y=7.4 //x2=69.19 //y2=7.4
r1417 (  775 977 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=69.455 //y=7.4 //x2=69.54 //y2=7.4
r1418 (  775 778 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=69.455 //y=7.4 //x2=69.19 //y2=7.4
r1419 (  772 975 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.755 //y=7.4 //x2=67.67 //y2=7.4
r1420 (  771 976 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=68.28 //y=7.4 //x2=68.45 //y2=7.4
r1421 (  771 772 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=68.28 //y=7.4 //x2=67.755 //y2=7.4
r1422 (  765 975 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=67.67 //y=7.23 //x2=67.67 //y2=7.4
r1423 (  765 1051 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=67.67 //y=7.23 //x2=67.67 //y2=6.745
r1424 (  764 973 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.875 //y=7.4 //x2=66.79 //y2=7.4
r1425 (  763 975 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.585 //y=7.4 //x2=67.67 //y2=7.4
r1426 (  763 764 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=67.585 //y=7.4 //x2=66.875 //y2=7.4
r1427 (  757 973 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=66.79 //y=7.23 //x2=66.79 //y2=7.4
r1428 (  757 1050 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=66.79 //y=7.23 //x2=66.79 //y2=6.745
r1429 (  754 972 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.995 //y=7.4 //x2=65.91 //y2=7.4
r1430 (  754 756 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=65.995 //y=7.4 //x2=66.6 //y2=7.4
r1431 (  753 973 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=66.705 //y=7.4 //x2=66.79 //y2=7.4
r1432 (  753 756 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=66.705 //y=7.4 //x2=66.6 //y2=7.4
r1433 (  747 972 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=65.91 //y=7.23 //x2=65.91 //y2=7.4
r1434 (  747 1049 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=65.91 //y=7.23 //x2=65.91 //y2=6.405
r1435 (  744 971 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=65.29 //y=7.4 //x2=65.12 //y2=7.4
r1436 (  744 746 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=65.29 //y=7.4 //x2=65.49 //y2=7.4
r1437 (  743 972 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=65.825 //y=7.4 //x2=65.91 //y2=7.4
r1438 (  743 746 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=65.825 //y=7.4 //x2=65.49 //y2=7.4
r1439 (  740 970 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.425 //y=7.4 //x2=64.34 //y2=7.4
r1440 (  739 971 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.95 //y=7.4 //x2=65.12 //y2=7.4
r1441 (  739 740 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=64.95 //y=7.4 //x2=64.425 //y2=7.4
r1442 (  733 970 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=64.34 //y=7.23 //x2=64.34 //y2=7.4
r1443 (  733 1048 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=64.34 //y=7.23 //x2=64.34 //y2=6.745
r1444 (  730 969 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.545 //y=7.4 //x2=63.46 //y2=7.4
r1445 (  730 732 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=63.545 //y=7.4 //x2=64.01 //y2=7.4
r1446 (  729 970 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=64.255 //y=7.4 //x2=64.34 //y2=7.4
r1447 (  729 732 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=64.255 //y=7.4 //x2=64.01 //y2=7.4
r1448 (  723 969 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=63.46 //y=7.23 //x2=63.46 //y2=7.4
r1449 (  723 1047 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=63.46 //y=7.23 //x2=63.46 //y2=6.745
r1450 (  720 968 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.665 //y=7.4 //x2=62.58 //y2=7.4
r1451 (  720 722 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=62.665 //y=7.4 //x2=62.9 //y2=7.4
r1452 (  719 969 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.375 //y=7.4 //x2=63.46 //y2=7.4
r1453 (  719 722 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=63.375 //y=7.4 //x2=62.9 //y2=7.4
r1454 (  713 968 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=62.58 //y=7.23 //x2=62.58 //y2=7.4
r1455 (  713 1046 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=62.58 //y=7.23 //x2=62.58 //y2=6.405
r1456 (  712 967 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.96 //y=7.4 //x2=61.79 //y2=7.4
r1457 (  711 968 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=62.495 //y=7.4 //x2=62.58 //y2=7.4
r1458 (  711 712 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=62.495 //y=7.4 //x2=61.96 //y2=7.4
r1459 (  706 966 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.795 //y=7.4 //x2=60.71 //y2=7.4
r1460 (  706 708 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=60.795 //y=7.4 //x2=61.42 //y2=7.4
r1461 (  705 967 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=61.62 //y=7.4 //x2=61.79 //y2=7.4
r1462 (  705 708 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=61.62 //y=7.4 //x2=61.42 //y2=7.4
r1463 (  699 966 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=60.71 //y=7.23 //x2=60.71 //y2=7.4
r1464 (  699 1045 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=60.71 //y=7.23 //x2=60.71 //y2=6.745
r1465 (  696 965 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.915 //y=7.4 //x2=59.83 //y2=7.4
r1466 (  696 698 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=59.915 //y=7.4 //x2=60.31 //y2=7.4
r1467 (  695 966 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.625 //y=7.4 //x2=60.71 //y2=7.4
r1468 (  695 698 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=60.625 //y=7.4 //x2=60.31 //y2=7.4
r1469 (  689 965 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=59.83 //y=7.23 //x2=59.83 //y2=7.4
r1470 (  689 1044 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=59.83 //y=7.23 //x2=59.83 //y2=6.745
r1471 (  686 964 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.035 //y=7.4 //x2=58.95 //y2=7.4
r1472 (  686 688 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=59.035 //y=7.4 //x2=59.2 //y2=7.4
r1473 (  685 965 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.745 //y=7.4 //x2=59.83 //y2=7.4
r1474 (  685 688 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=59.745 //y=7.4 //x2=59.2 //y2=7.4
r1475 (  679 964 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.95 //y=7.23 //x2=58.95 //y2=7.4
r1476 (  679 1043 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=58.95 //y=7.23 //x2=58.95 //y2=6.745
r1477 (  678 963 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.155 //y=7.4 //x2=58.07 //y2=7.4
r1478 (  677 964 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=58.865 //y=7.4 //x2=58.95 //y2=7.4
r1479 (  677 678 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=58.865 //y=7.4 //x2=58.155 //y2=7.4
r1480 (  671 963 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=58.07 //y=7.23 //x2=58.07 //y2=7.4
r1481 (  671 1042 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=58.07 //y=7.23 //x2=58.07 //y2=6.405
r1482 (  670 961 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=57.15 //y=7.4 //x2=56.98 //y2=7.4
r1483 (  669 963 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=57.985 //y=7.4 //x2=58.07 //y2=7.4
r1484 (  669 670 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=57.985 //y=7.4 //x2=57.15 //y2=7.4
r1485 (  664 960 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.985 //y=7.4 //x2=55.9 //y2=7.4
r1486 (  664 666 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=55.985 //y=7.4 //x2=56.61 //y2=7.4
r1487 (  663 961 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=56.81 //y=7.4 //x2=56.98 //y2=7.4
r1488 (  663 666 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=56.81 //y=7.4 //x2=56.61 //y2=7.4
r1489 (  657 960 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=55.9 //y=7.23 //x2=55.9 //y2=7.4
r1490 (  657 1041 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=55.9 //y=7.23 //x2=55.9 //y2=6.745
r1491 (  654 959 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.105 //y=7.4 //x2=55.02 //y2=7.4
r1492 (  654 656 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=55.105 //y=7.4 //x2=55.5 //y2=7.4
r1493 (  653 960 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.815 //y=7.4 //x2=55.9 //y2=7.4
r1494 (  653 656 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=55.815 //y=7.4 //x2=55.5 //y2=7.4
r1495 (  647 959 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=55.02 //y=7.23 //x2=55.02 //y2=7.4
r1496 (  647 1040 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=55.02 //y=7.23 //x2=55.02 //y2=6.745
r1497 (  644 958 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.225 //y=7.4 //x2=54.14 //y2=7.4
r1498 (  644 646 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=54.225 //y=7.4 //x2=54.39 //y2=7.4
r1499 (  643 959 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.935 //y=7.4 //x2=55.02 //y2=7.4
r1500 (  643 646 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=54.935 //y=7.4 //x2=54.39 //y2=7.4
r1501 (  637 958 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=54.14 //y=7.23 //x2=54.14 //y2=7.4
r1502 (  637 1039 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=54.14 //y=7.23 //x2=54.14 //y2=6.745
r1503 (  636 957 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.345 //y=7.4 //x2=53.26 //y2=7.4
r1504 (  635 958 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.055 //y=7.4 //x2=54.14 //y2=7.4
r1505 (  635 636 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=54.055 //y=7.4 //x2=53.345 //y2=7.4
r1506 (  629 957 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=53.26 //y=7.23 //x2=53.26 //y2=7.4
r1507 (  629 1038 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=53.26 //y=7.23 //x2=53.26 //y2=6.405
r1508 (  628 955 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=52.34 //y=7.4 //x2=52.17 //y2=7.4
r1509 (  627 957 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=53.175 //y=7.4 //x2=53.26 //y2=7.4
r1510 (  627 628 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=53.175 //y=7.4 //x2=52.34 //y2=7.4
r1511 (  622 954 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.475 //y=7.4 //x2=51.39 //y2=7.4
r1512 (  622 624 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=51.475 //y=7.4 //x2=51.8 //y2=7.4
r1513 (  621 955 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=52 //y=7.4 //x2=52.17 //y2=7.4
r1514 (  621 624 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=52 //y=7.4 //x2=51.8 //y2=7.4
r1515 (  615 954 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=51.39 //y=7.23 //x2=51.39 //y2=7.4
r1516 (  615 1037 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=51.39 //y=7.23 //x2=51.39 //y2=6.745
r1517 (  612 953 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.595 //y=7.4 //x2=50.51 //y2=7.4
r1518 (  612 614 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=50.595 //y=7.4 //x2=50.69 //y2=7.4
r1519 (  611 954 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.305 //y=7.4 //x2=51.39 //y2=7.4
r1520 (  611 614 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=51.305 //y=7.4 //x2=50.69 //y2=7.4
r1521 (  605 953 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=50.51 //y=7.23 //x2=50.51 //y2=7.4
r1522 (  605 1036 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=50.51 //y=7.23 //x2=50.51 //y2=6.745
r1523 (  604 952 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.715 //y=7.4 //x2=49.63 //y2=7.4
r1524 (  603 953 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.425 //y=7.4 //x2=50.51 //y2=7.4
r1525 (  603 604 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=50.425 //y=7.4 //x2=49.715 //y2=7.4
r1526 (  597 952 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.63 //y=7.23 //x2=49.63 //y2=7.4
r1527 (  597 1035 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=49.63 //y=7.23 //x2=49.63 //y2=6.405
r1528 (  596 950 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=49.01 //y=7.4 //x2=48.84 //y2=7.4
r1529 (  595 952 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=49.545 //y=7.4 //x2=49.63 //y2=7.4
r1530 (  595 596 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=49.545 //y=7.4 //x2=49.01 //y2=7.4
r1531 (  590 949 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.845 //y=7.4 //x2=47.76 //y2=7.4
r1532 (  590 592 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=47.845 //y=7.4 //x2=48.1 //y2=7.4
r1533 (  589 950 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=48.67 //y=7.4 //x2=48.84 //y2=7.4
r1534 (  589 592 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=48.67 //y=7.4 //x2=48.1 //y2=7.4
r1535 (  583 949 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=47.76 //y=7.23 //x2=47.76 //y2=7.4
r1536 (  583 1034 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=47.76 //y=7.23 //x2=47.76 //y2=6.745
r1537 (  580 948 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.965 //y=7.4 //x2=46.88 //y2=7.4
r1538 (  580 582 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=46.965 //y=7.4 //x2=46.99 //y2=7.4
r1539 (  579 949 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.675 //y=7.4 //x2=47.76 //y2=7.4
r1540 (  579 582 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=47.675 //y=7.4 //x2=46.99 //y2=7.4
r1541 (  573 948 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=46.88 //y=7.23 //x2=46.88 //y2=7.4
r1542 (  573 1033 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.88 //y=7.23 //x2=46.88 //y2=6.745
r1543 (  572 947 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.085 //y=7.4 //x2=46 //y2=7.4
r1544 (  571 948 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.795 //y=7.4 //x2=46.88 //y2=7.4
r1545 (  571 572 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=46.795 //y=7.4 //x2=46.085 //y2=7.4
r1546 (  565 947 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=46 //y=7.23 //x2=46 //y2=7.4
r1547 (  565 1032 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46 //y=7.23 //x2=46 //y2=6.745
r1548 (  562 946 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.205 //y=7.4 //x2=45.12 //y2=7.4
r1549 (  562 564 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=45.205 //y=7.4 //x2=45.88 //y2=7.4
r1550 (  561 947 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.915 //y=7.4 //x2=46 //y2=7.4
r1551 (  561 564 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=45.915 //y=7.4 //x2=45.88 //y2=7.4
r1552 (  555 946 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=45.12 //y=7.23 //x2=45.12 //y2=7.4
r1553 (  555 1031 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=45.12 //y=7.23 //x2=45.12 //y2=6.405
r1554 (  552 945 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=44.2 //y=7.4 //x2=44.03 //y2=7.4
r1555 (  552 554 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=44.2 //y=7.4 //x2=44.77 //y2=7.4
r1556 (  551 946 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=45.035 //y=7.4 //x2=45.12 //y2=7.4
r1557 (  551 554 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=45.035 //y=7.4 //x2=44.77 //y2=7.4
r1558 (  548 944 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=43.335 //y=7.4 //x2=43.25 //y2=7.4
r1559 (  547 945 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.86 //y=7.4 //x2=44.03 //y2=7.4
r1560 (  547 548 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=43.86 //y=7.4 //x2=43.335 //y2=7.4
r1561 (  541 944 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=43.25 //y=7.23 //x2=43.25 //y2=7.4
r1562 (  541 1030 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=43.25 //y=7.23 //x2=43.25 //y2=6.745
r1563 (  540 942 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.455 //y=7.4 //x2=42.37 //y2=7.4
r1564 (  539 944 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=43.165 //y=7.4 //x2=43.25 //y2=7.4
r1565 (  539 540 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=43.165 //y=7.4 //x2=42.455 //y2=7.4
r1566 (  533 942 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=42.37 //y=7.23 //x2=42.37 //y2=7.4
r1567 (  533 1029 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=42.37 //y=7.23 //x2=42.37 //y2=6.745
r1568 (  530 941 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.575 //y=7.4 //x2=41.49 //y2=7.4
r1569 (  530 532 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=41.575 //y=7.4 //x2=42.18 //y2=7.4
r1570 (  529 942 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.285 //y=7.4 //x2=42.37 //y2=7.4
r1571 (  529 532 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=42.285 //y=7.4 //x2=42.18 //y2=7.4
r1572 (  523 941 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=41.49 //y=7.23 //x2=41.49 //y2=7.4
r1573 (  523 1028 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=41.49 //y=7.23 //x2=41.49 //y2=6.405
r1574 (  520 940 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.87 //y=7.4 //x2=40.7 //y2=7.4
r1575 (  520 522 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=40.87 //y=7.4 //x2=41.07 //y2=7.4
r1576 (  519 941 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=41.405 //y=7.4 //x2=41.49 //y2=7.4
r1577 (  519 522 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=41.405 //y=7.4 //x2=41.07 //y2=7.4
r1578 (  516 939 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=40.005 //y=7.4 //x2=39.92 //y2=7.4
r1579 (  515 940 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=40.53 //y=7.4 //x2=40.7 //y2=7.4
r1580 (  515 516 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=40.53 //y=7.4 //x2=40.005 //y2=7.4
r1581 (  509 939 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.92 //y=7.23 //x2=39.92 //y2=7.4
r1582 (  509 1027 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=39.92 //y=7.23 //x2=39.92 //y2=6.745
r1583 (  506 938 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.125 //y=7.4 //x2=39.04 //y2=7.4
r1584 (  506 508 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=39.125 //y=7.4 //x2=39.59 //y2=7.4
r1585 (  505 939 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.835 //y=7.4 //x2=39.92 //y2=7.4
r1586 (  505 508 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=39.835 //y=7.4 //x2=39.59 //y2=7.4
r1587 (  499 938 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=39.04 //y=7.23 //x2=39.04 //y2=7.4
r1588 (  499 1026 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=39.04 //y=7.23 //x2=39.04 //y2=6.745
r1589 (  496 937 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.245 //y=7.4 //x2=38.16 //y2=7.4
r1590 (  496 498 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=38.245 //y=7.4 //x2=38.48 //y2=7.4
r1591 (  495 938 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.955 //y=7.4 //x2=39.04 //y2=7.4
r1592 (  495 498 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=38.955 //y=7.4 //x2=38.48 //y2=7.4
r1593 (  489 937 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=38.16 //y=7.23 //x2=38.16 //y2=7.4
r1594 (  489 1025 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=38.16 //y=7.23 //x2=38.16 //y2=6.405
r1595 (  488 936 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.54 //y=7.4 //x2=37.37 //y2=7.4
r1596 (  487 937 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=38.075 //y=7.4 //x2=38.16 //y2=7.4
r1597 (  487 488 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=38.075 //y=7.4 //x2=37.54 //y2=7.4
r1598 (  482 935 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.375 //y=7.4 //x2=36.29 //y2=7.4
r1599 (  482 484 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=36.375 //y=7.4 //x2=37 //y2=7.4
r1600 (  481 936 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=37.2 //y=7.4 //x2=37.37 //y2=7.4
r1601 (  481 484 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=37.2 //y=7.4 //x2=37 //y2=7.4
r1602 (  475 935 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=36.29 //y=7.23 //x2=36.29 //y2=7.4
r1603 (  475 1024 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=36.29 //y=7.23 //x2=36.29 //y2=6.745
r1604 (  472 934 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.495 //y=7.4 //x2=35.41 //y2=7.4
r1605 (  472 474 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=35.495 //y=7.4 //x2=35.89 //y2=7.4
r1606 (  471 935 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=36.205 //y=7.4 //x2=36.29 //y2=7.4
r1607 (  471 474 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=36.205 //y=7.4 //x2=35.89 //y2=7.4
r1608 (  465 934 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=35.41 //y=7.23 //x2=35.41 //y2=7.4
r1609 (  465 1023 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=35.41 //y=7.23 //x2=35.41 //y2=6.745
r1610 (  462 933 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.615 //y=7.4 //x2=34.53 //y2=7.4
r1611 (  462 464 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=34.615 //y=7.4 //x2=34.78 //y2=7.4
r1612 (  461 934 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.325 //y=7.4 //x2=35.41 //y2=7.4
r1613 (  461 464 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=35.325 //y=7.4 //x2=34.78 //y2=7.4
r1614 (  455 933 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=34.53 //y=7.23 //x2=34.53 //y2=7.4
r1615 (  455 1022 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=34.53 //y=7.23 //x2=34.53 //y2=6.745
r1616 (  454 932 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.735 //y=7.4 //x2=33.65 //y2=7.4
r1617 (  453 933 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.445 //y=7.4 //x2=34.53 //y2=7.4
r1618 (  453 454 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=34.445 //y=7.4 //x2=33.735 //y2=7.4
r1619 (  447 932 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=33.65 //y=7.23 //x2=33.65 //y2=7.4
r1620 (  447 1021 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=33.65 //y=7.23 //x2=33.65 //y2=6.405
r1621 (  446 930 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.73 //y=7.4 //x2=32.56 //y2=7.4
r1622 (  445 932 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=33.565 //y=7.4 //x2=33.65 //y2=7.4
r1623 (  445 446 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=33.565 //y=7.4 //x2=32.73 //y2=7.4
r1624 (  440 929 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.565 //y=7.4 //x2=31.48 //y2=7.4
r1625 (  440 442 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=31.565 //y=7.4 //x2=32.19 //y2=7.4
r1626 (  439 930 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=32.39 //y=7.4 //x2=32.56 //y2=7.4
r1627 (  439 442 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=32.39 //y=7.4 //x2=32.19 //y2=7.4
r1628 (  433 929 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=31.48 //y=7.23 //x2=31.48 //y2=7.4
r1629 (  433 1020 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=31.48 //y=7.23 //x2=31.48 //y2=6.745
r1630 (  430 928 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.685 //y=7.4 //x2=30.6 //y2=7.4
r1631 (  430 432 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=30.685 //y=7.4 //x2=31.08 //y2=7.4
r1632 (  429 929 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.395 //y=7.4 //x2=31.48 //y2=7.4
r1633 (  429 432 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=31.395 //y=7.4 //x2=31.08 //y2=7.4
r1634 (  423 928 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=30.6 //y=7.23 //x2=30.6 //y2=7.4
r1635 (  423 1019 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=30.6 //y=7.23 //x2=30.6 //y2=6.745
r1636 (  420 927 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.805 //y=7.4 //x2=29.72 //y2=7.4
r1637 (  420 422 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=29.805 //y=7.4 //x2=29.97 //y2=7.4
r1638 (  419 928 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.515 //y=7.4 //x2=30.6 //y2=7.4
r1639 (  419 422 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=30.515 //y=7.4 //x2=29.97 //y2=7.4
r1640 (  413 927 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=29.72 //y=7.23 //x2=29.72 //y2=7.4
r1641 (  413 1018 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=29.72 //y=7.23 //x2=29.72 //y2=6.745
r1642 (  412 926 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.925 //y=7.4 //x2=28.84 //y2=7.4
r1643 (  411 927 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.635 //y=7.4 //x2=29.72 //y2=7.4
r1644 (  411 412 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=29.635 //y=7.4 //x2=28.925 //y2=7.4
r1645 (  405 926 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=28.84 //y=7.23 //x2=28.84 //y2=7.4
r1646 (  405 1017 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=28.84 //y=7.23 //x2=28.84 //y2=6.405
r1647 (  404 924 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.92 //y=7.4 //x2=27.75 //y2=7.4
r1648 (  403 926 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=28.755 //y=7.4 //x2=28.84 //y2=7.4
r1649 (  403 404 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=28.755 //y=7.4 //x2=27.92 //y2=7.4
r1650 (  398 923 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=27.055 //y=7.4 //x2=26.97 //y2=7.4
r1651 (  398 400 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=27.055 //y=7.4 //x2=27.38 //y2=7.4
r1652 (  397 924 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=27.58 //y=7.4 //x2=27.75 //y2=7.4
r1653 (  397 400 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=27.58 //y=7.4 //x2=27.38 //y2=7.4
r1654 (  391 923 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.97 //y=7.23 //x2=26.97 //y2=7.4
r1655 (  391 1016 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.97 //y=7.23 //x2=26.97 //y2=6.745
r1656 (  388 922 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.175 //y=7.4 //x2=26.09 //y2=7.4
r1657 (  388 390 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=26.175 //y=7.4 //x2=26.27 //y2=7.4
r1658 (  387 923 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.885 //y=7.4 //x2=26.97 //y2=7.4
r1659 (  387 390 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=26.885 //y=7.4 //x2=26.27 //y2=7.4
r1660 (  381 922 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=26.09 //y=7.23 //x2=26.09 //y2=7.4
r1661 (  381 1015 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=26.09 //y=7.23 //x2=26.09 //y2=6.745
r1662 (  380 921 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.295 //y=7.4 //x2=25.21 //y2=7.4
r1663 (  379 922 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.005 //y=7.4 //x2=26.09 //y2=7.4
r1664 (  379 380 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=26.005 //y=7.4 //x2=25.295 //y2=7.4
r1665 (  373 921 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.21 //y=7.23 //x2=25.21 //y2=7.4
r1666 (  373 1014 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=25.21 //y=7.23 //x2=25.21 //y2=6.405
r1667 (  372 919 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.59 //y=7.4 //x2=24.42 //y2=7.4
r1668 (  371 921 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.125 //y=7.4 //x2=25.21 //y2=7.4
r1669 (  371 372 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=25.125 //y=7.4 //x2=24.59 //y2=7.4
r1670 (  366 918 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.425 //y=7.4 //x2=23.34 //y2=7.4
r1671 (  366 368 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=23.425 //y=7.4 //x2=23.68 //y2=7.4
r1672 (  365 919 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.25 //y=7.4 //x2=24.42 //y2=7.4
r1673 (  365 368 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.25 //y=7.4 //x2=23.68 //y2=7.4
r1674 (  359 918 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.34 //y=7.23 //x2=23.34 //y2=7.4
r1675 (  359 1013 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=23.34 //y=7.23 //x2=23.34 //y2=6.745
r1676 (  356 917 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.545 //y=7.4 //x2=22.46 //y2=7.4
r1677 (  356 358 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=22.545 //y=7.4 //x2=22.57 //y2=7.4
r1678 (  355 918 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.255 //y=7.4 //x2=23.34 //y2=7.4
r1679 (  355 358 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=23.255 //y=7.4 //x2=22.57 //y2=7.4
r1680 (  349 917 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.46 //y=7.23 //x2=22.46 //y2=7.4
r1681 (  349 1012 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.46 //y=7.23 //x2=22.46 //y2=6.745
r1682 (  348 916 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.665 //y=7.4 //x2=21.58 //y2=7.4
r1683 (  347 917 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.375 //y=7.4 //x2=22.46 //y2=7.4
r1684 (  347 348 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.375 //y=7.4 //x2=21.665 //y2=7.4
r1685 (  341 916 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.58 //y=7.23 //x2=21.58 //y2=7.4
r1686 (  341 1011 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.58 //y=7.23 //x2=21.58 //y2=6.745
r1687 (  338 915 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.785 //y=7.4 //x2=20.7 //y2=7.4
r1688 (  338 340 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=20.785 //y=7.4 //x2=21.46 //y2=7.4
r1689 (  337 916 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.495 //y=7.4 //x2=21.58 //y2=7.4
r1690 (  337 340 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=21.495 //y=7.4 //x2=21.46 //y2=7.4
r1691 (  331 915 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.7 //y=7.23 //x2=20.7 //y2=7.4
r1692 (  331 1010 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=20.7 //y=7.23 //x2=20.7 //y2=6.405
r1693 (  328 914 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.78 //y=7.4 //x2=19.61 //y2=7.4
r1694 (  328 330 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=19.78 //y=7.4 //x2=20.35 //y2=7.4
r1695 (  327 915 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.615 //y=7.4 //x2=20.7 //y2=7.4
r1696 (  327 330 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=20.615 //y=7.4 //x2=20.35 //y2=7.4
r1697 (  324 913 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.915 //y=7.4 //x2=18.83 //y2=7.4
r1698 (  323 914 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.44 //y=7.4 //x2=19.61 //y2=7.4
r1699 (  323 324 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=19.44 //y=7.4 //x2=18.915 //y2=7.4
r1700 (  317 913 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.83 //y=7.23 //x2=18.83 //y2=7.4
r1701 (  317 1009 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=18.83 //y=7.23 //x2=18.83 //y2=6.745
r1702 (  316 911 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.035 //y=7.4 //x2=17.95 //y2=7.4
r1703 (  315 913 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.745 //y=7.4 //x2=18.83 //y2=7.4
r1704 (  315 316 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=18.745 //y=7.4 //x2=18.035 //y2=7.4
r1705 (  309 911 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.95 //y=7.23 //x2=17.95 //y2=7.4
r1706 (  309 1008 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=17.95 //y=7.23 //x2=17.95 //y2=6.745
r1707 (  306 910 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.155 //y=7.4 //x2=17.07 //y2=7.4
r1708 (  306 308 ) resistor r=21.6919 //w=0.357 //l=0.605 //layer=li \
 //thickness=0.1 //x=17.155 //y=7.4 //x2=17.76 //y2=7.4
r1709 (  305 911 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=17.865 //y=7.4 //x2=17.95 //y2=7.4
r1710 (  305 308 ) resistor r=3.76471 //w=0.357 //l=0.105 //layer=li \
 //thickness=0.1 //x=17.865 //y=7.4 //x2=17.76 //y2=7.4
r1711 (  299 910 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.07 //y=7.23 //x2=17.07 //y2=7.4
r1712 (  299 1007 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=17.07 //y=7.23 //x2=17.07 //y2=6.405
r1713 (  296 909 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.45 //y=7.4 //x2=16.28 //y2=7.4
r1714 (  296 298 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=16.45 //y=7.4 //x2=16.65 //y2=7.4
r1715 (  295 910 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.985 //y=7.4 //x2=17.07 //y2=7.4
r1716 (  295 298 ) resistor r=12.0112 //w=0.357 //l=0.335 //layer=li \
 //thickness=0.1 //x=16.985 //y=7.4 //x2=16.65 //y2=7.4
r1717 (  292 908 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.585 //y=7.4 //x2=15.5 //y2=7.4
r1718 (  291 909 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.11 //y=7.4 //x2=16.28 //y2=7.4
r1719 (  291 292 ) resistor r=18.8235 //w=0.357 //l=0.525 //layer=li \
 //thickness=0.1 //x=16.11 //y=7.4 //x2=15.585 //y2=7.4
r1720 (  285 908 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.5 //y=7.23 //x2=15.5 //y2=7.4
r1721 (  285 1006 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.5 //y=7.23 //x2=15.5 //y2=6.745
r1722 (  282 907 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.705 //y=7.4 //x2=14.62 //y2=7.4
r1723 (  282 284 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=14.705 //y=7.4 //x2=15.17 //y2=7.4
r1724 (  281 908 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.415 //y=7.4 //x2=15.5 //y2=7.4
r1725 (  281 284 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=15.415 //y=7.4 //x2=15.17 //y2=7.4
r1726 (  275 907 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.62 //y=7.23 //x2=14.62 //y2=7.4
r1727 (  275 1005 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.62 //y=7.23 //x2=14.62 //y2=6.745
r1728 (  272 906 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.825 //y=7.4 //x2=13.74 //y2=7.4
r1729 (  272 274 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=13.825 //y=7.4 //x2=14.06 //y2=7.4
r1730 (  271 907 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.535 //y=7.4 //x2=14.62 //y2=7.4
r1731 (  271 274 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=14.535 //y=7.4 //x2=14.06 //y2=7.4
r1732 (  265 906 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.74 //y=7.23 //x2=13.74 //y2=7.4
r1733 (  265 1004 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=13.74 //y=7.23 //x2=13.74 //y2=6.405
r1734 (  264 905 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.12 //y=7.4 //x2=12.95 //y2=7.4
r1735 (  263 906 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.655 //y=7.4 //x2=13.74 //y2=7.4
r1736 (  263 264 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=13.655 //y=7.4 //x2=13.12 //y2=7.4
r1737 (  258 904 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.955 //y=7.4 //x2=11.87 //y2=7.4
r1738 (  258 260 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=11.955 //y=7.4 //x2=12.58 //y2=7.4
r1739 (  257 905 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.78 //y=7.4 //x2=12.95 //y2=7.4
r1740 (  257 260 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.78 //y=7.4 //x2=12.58 //y2=7.4
r1741 (  251 904 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.87 //y=7.23 //x2=11.87 //y2=7.4
r1742 (  251 1003 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.87 //y=7.23 //x2=11.87 //y2=6.745
r1743 (  248 903 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.075 //y=7.4 //x2=10.99 //y2=7.4
r1744 (  248 250 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=11.075 //y=7.4 //x2=11.47 //y2=7.4
r1745 (  247 904 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.785 //y=7.4 //x2=11.87 //y2=7.4
r1746 (  247 250 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=11.785 //y=7.4 //x2=11.47 //y2=7.4
r1747 (  241 903 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.99 //y=7.23 //x2=10.99 //y2=7.4
r1748 (  241 1002 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.99 //y=7.23 //x2=10.99 //y2=6.745
r1749 (  238 902 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.195 //y=7.4 //x2=10.11 //y2=7.4
r1750 (  238 240 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=10.195 //y=7.4 //x2=10.36 //y2=7.4
r1751 (  237 903 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.905 //y=7.4 //x2=10.99 //y2=7.4
r1752 (  237 240 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=10.905 //y=7.4 //x2=10.36 //y2=7.4
r1753 (  231 902 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.11 //y=7.23 //x2=10.11 //y2=7.4
r1754 (  231 1001 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.11 //y=7.23 //x2=10.11 //y2=6.745
r1755 (  230 901 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.315 //y=7.4 //x2=9.23 //y2=7.4
r1756 (  229 902 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.025 //y=7.4 //x2=10.11 //y2=7.4
r1757 (  229 230 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.025 //y=7.4 //x2=9.315 //y2=7.4
r1758 (  223 901 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.23 //y=7.23 //x2=9.23 //y2=7.4
r1759 (  223 1000 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=9.23 //y=7.23 //x2=9.23 //y2=6.405
r1760 (  222 899 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.31 //y=7.4 //x2=8.14 //y2=7.4
r1761 (  221 901 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=9.145 //y=7.4 //x2=9.23 //y2=7.4
r1762 (  221 222 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=9.145 //y=7.4 //x2=8.31 //y2=7.4
r1763 (  216 898 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.145 //y=7.4 //x2=7.06 //y2=7.4
r1764 (  216 218 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=7.145 //y=7.4 //x2=7.77 //y2=7.4
r1765 (  215 899 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=8.14 //y2=7.4
r1766 (  215 218 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=7.97 //y=7.4 //x2=7.77 //y2=7.4
r1767 (  209 898 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.06 //y=7.23 //x2=7.06 //y2=7.4
r1768 (  209 999 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.06 //y=7.23 //x2=7.06 //y2=6.745
r1769 (  206 897 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.265 //y=7.4 //x2=6.18 //y2=7.4
r1770 (  206 208 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=6.265 //y=7.4 //x2=6.66 //y2=7.4
r1771 (  205 898 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.975 //y=7.4 //x2=7.06 //y2=7.4
r1772 (  205 208 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=6.975 //y=7.4 //x2=6.66 //y2=7.4
r1773 (  199 897 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.18 //y=7.23 //x2=6.18 //y2=7.4
r1774 (  199 998 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.18 //y=7.23 //x2=6.18 //y2=6.745
r1775 (  196 896 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.385 //y=7.4 //x2=5.3 //y2=7.4
r1776 (  196 198 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=5.385 //y=7.4 //x2=5.55 //y2=7.4
r1777 (  195 897 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.095 //y=7.4 //x2=6.18 //y2=7.4
r1778 (  195 198 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=6.095 //y=7.4 //x2=5.55 //y2=7.4
r1779 (  189 896 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.3 //y=7.23 //x2=5.3 //y2=7.4
r1780 (  189 997 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=5.3 //y=7.23 //x2=5.3 //y2=6.745
r1781 (  188 895 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.505 //y=7.4 //x2=4.42 //y2=7.4
r1782 (  187 896 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.215 //y=7.4 //x2=5.3 //y2=7.4
r1783 (  187 188 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=5.215 //y=7.4 //x2=4.505 //y2=7.4
r1784 (  181 895 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.42 //y=7.23 //x2=4.42 //y2=7.4
r1785 (  181 996 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=4.42 //y=7.23 //x2=4.42 //y2=6.405
r1786 (  180 893 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=7.4 //x2=3.33 //y2=7.4
r1787 (  179 895 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.335 //y=7.4 //x2=4.42 //y2=7.4
r1788 (  179 180 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=4.335 //y=7.4 //x2=3.5 //y2=7.4
r1789 (  174 892 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.55 //y2=7.4
r1790 (  174 176 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=2.635 //y=7.4 //x2=2.96 //y2=7.4
r1791 (  173 893 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=3.33 //y2=7.4
r1792 (  173 176 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=2.96 //y2=7.4
r1793 (  167 892 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=7.4
r1794 (  167 995 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.55 //y=7.23 //x2=2.55 //y2=6.745
r1795 (  164 891 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.67 //y2=7.4
r1796 (  164 166 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=1.755 //y=7.4 //x2=1.85 //y2=7.4
r1797 (  163 892 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=2.55 //y2=7.4
r1798 (  163 166 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=2.465 //y=7.4 //x2=1.85 //y2=7.4
r1799 (  157 891 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=7.4
r1800 (  157 994 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.67 //y=7.23 //x2=1.67 //y2=6.745
r1801 (  156 890 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.875 //y=7.4 //x2=0.79 //y2=7.4
r1802 (  155 891 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=1.67 //y2=7.4
r1803 (  155 156 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=1.585 //y=7.4 //x2=0.875 //y2=7.4
r1804 (  149 890 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=7.4
r1805 (  149 993 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=0.79 //y=7.23 //x2=0.79 //y2=6.405
r1806 (  143 992 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=84.73 //y=7.4 //x2=84.73 //y2=7.4
r1807 (  141 990 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=83.99 //y=7.4 //x2=83.99 //y2=7.4
r1808 (  141 143 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=83.99 //y=7.4 //x2=84.73 //y2=7.4
r1809 (  139 866 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=82.51 //y=7.4 //x2=82.51 //y2=7.4
r1810 (  139 141 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=82.51 //y=7.4 //x2=83.99 //y2=7.4
r1811 (  137 864 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=81.4 //y=7.4 //x2=81.4 //y2=7.4
r1812 (  137 139 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=81.4 //y=7.4 //x2=82.51 //y2=7.4
r1813 (  135 862 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=80.29 //y=7.4 //x2=80.29 //y2=7.4
r1814 (  135 137 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=80.29 //y=7.4 //x2=81.4 //y2=7.4
r1815 (  133 856 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=78.81 //y=7.4 //x2=78.81 //y2=7.4
r1816 (  133 135 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=78.81 //y=7.4 //x2=80.29 //y2=7.4
r1817 (  131 854 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=77.7 //y=7.4 //x2=77.7 //y2=7.4
r1818 (  131 133 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=77.7 //y=7.4 //x2=78.81 //y2=7.4
r1819 (  129 848 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=76.22 //y=7.4 //x2=76.22 //y2=7.4
r1820 (  129 131 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=76.22 //y=7.4 //x2=77.7 //y2=7.4
r1821 (  127 838 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=75.11 //y=7.4 //x2=75.11 //y2=7.4
r1822 (  127 129 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=75.11 //y=7.4 //x2=76.22 //y2=7.4
r1823 (  125 983 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=74 //y=7.4 //x2=74 //y2=7.4
r1824 (  125 127 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=74 //y=7.4 //x2=75.11 //y2=7.4
r1825 (  123 816 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=72.52 //y=7.4 //x2=72.52 //y2=7.4
r1826 (  123 125 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=72.52 //y=7.4 //x2=74 //y2=7.4
r1827 (  121 806 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=71.41 //y=7.4 //x2=71.41 //y2=7.4
r1828 (  121 123 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=71.41 //y=7.4 //x2=72.52 //y2=7.4
r1829 (  119 788 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=70.3 //y=7.4 //x2=70.3 //y2=7.4
r1830 (  119 121 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=70.3 //y=7.4 //x2=71.41 //y2=7.4
r1831 (  117 778 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=69.19 //y=7.4 //x2=69.19 //y2=7.4
r1832 (  117 119 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=69.19 //y=7.4 //x2=70.3 //y2=7.4
r1833 (  115 975 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=67.71 //y=7.4 //x2=67.71 //y2=7.4
r1834 (  115 117 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=67.71 //y=7.4 //x2=69.19 //y2=7.4
r1835 (  113 756 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=66.6 //y=7.4 //x2=66.6 //y2=7.4
r1836 (  113 115 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=66.6 //y=7.4 //x2=67.71 //y2=7.4
r1837 (  111 746 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=65.49 //y=7.4 //x2=65.49 //y2=7.4
r1838 (  111 113 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=65.49 //y=7.4 //x2=66.6 //y2=7.4
r1839 (  109 732 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=64.01 //y=7.4 //x2=64.01 //y2=7.4
r1840 (  109 111 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=64.01 //y=7.4 //x2=65.49 //y2=7.4
r1841 (  107 722 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=62.9 //y=7.4 //x2=62.9 //y2=7.4
r1842 (  107 109 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=62.9 //y=7.4 //x2=64.01 //y2=7.4
r1843 (  105 708 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=61.42 //y=7.4 //x2=61.42 //y2=7.4
r1844 (  105 107 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=61.42 //y=7.4 //x2=62.9 //y2=7.4
r1845 (  103 698 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=60.31 //y=7.4 //x2=60.31 //y2=7.4
r1846 (  103 105 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=60.31 //y=7.4 //x2=61.42 //y2=7.4
r1847 (  101 688 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=59.2 //y=7.4 //x2=59.2 //y2=7.4
r1848 (  101 103 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=59.2 //y=7.4 //x2=60.31 //y2=7.4
r1849 (  99 963 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=58.09 //y=7.4 //x2=58.09 //y2=7.4
r1850 (  99 101 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=58.09 //y=7.4 //x2=59.2 //y2=7.4
r1851 (  97 666 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=56.61 //y=7.4 //x2=56.61 //y2=7.4
r1852 (  97 99 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=56.61 //y=7.4 //x2=58.09 //y2=7.4
r1853 (  95 656 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=55.5 //y=7.4 //x2=55.5 //y2=7.4
r1854 (  95 97 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=55.5 //y=7.4 //x2=56.61 //y2=7.4
r1855 (  93 646 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=54.39 //y=7.4 //x2=54.39 //y2=7.4
r1856 (  93 95 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=54.39 //y=7.4 //x2=55.5 //y2=7.4
r1857 (  91 957 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=53.28 //y=7.4 //x2=53.28 //y2=7.4
r1858 (  91 93 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=53.28 //y=7.4 //x2=54.39 //y2=7.4
r1859 (  89 624 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=51.8 //y=7.4 //x2=51.8 //y2=7.4
r1860 (  89 91 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=51.8 //y=7.4 //x2=53.28 //y2=7.4
r1861 (  87 614 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=50.69 //y=7.4 //x2=50.69 //y2=7.4
r1862 (  87 89 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=50.69 //y=7.4 //x2=51.8 //y2=7.4
r1863 (  85 952 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=49.58 //y=7.4 //x2=49.58 //y2=7.4
r1864 (  85 87 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=49.58 //y=7.4 //x2=50.69 //y2=7.4
r1865 (  83 592 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=48.1 //y=7.4 //x2=48.1 //y2=7.4
r1866 (  83 85 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=48.1 //y=7.4 //x2=49.58 //y2=7.4
r1867 (  81 582 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=46.99 //y=7.4 //x2=46.99 //y2=7.4
r1868 (  81 83 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=46.99 //y=7.4 //x2=48.1 //y2=7.4
r1869 (  79 564 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=45.88 //y=7.4 //x2=45.88 //y2=7.4
r1870 (  79 81 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=45.88 //y=7.4 //x2=46.99 //y2=7.4
r1871 (  77 554 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=44.77 //y=7.4 //x2=44.77 //y2=7.4
r1872 (  77 79 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=44.77 //y=7.4 //x2=45.88 //y2=7.4
r1873 (  75 944 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=43.29 //y=7.4 //x2=43.29 //y2=7.4
r1874 (  75 77 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=43.29 //y=7.4 //x2=44.77 //y2=7.4
r1875 (  72 532 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=42.18 //y=7.4 //x2=42.18 //y2=7.4
r1876 (  70 522 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=41.07 //y=7.4 //x2=41.07 //y2=7.4
r1877 (  70 72 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=41.07 //y=7.4 //x2=42.18 //y2=7.4
r1878 (  68 508 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=39.59 //y=7.4 //x2=39.59 //y2=7.4
r1879 (  68 70 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=39.59 //y=7.4 //x2=41.07 //y2=7.4
r1880 (  66 498 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=38.48 //y=7.4 //x2=38.48 //y2=7.4
r1881 (  66 68 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=38.48 //y=7.4 //x2=39.59 //y2=7.4
r1882 (  64 484 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=37 //y=7.4 //x2=37 //y2=7.4
r1883 (  64 66 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=37 //y=7.4 //x2=38.48 //y2=7.4
r1884 (  62 474 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=35.89 //y=7.4 //x2=35.89 //y2=7.4
r1885 (  62 64 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=35.89 //y=7.4 //x2=37 //y2=7.4
r1886 (  60 464 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=34.78 //y=7.4 //x2=34.78 //y2=7.4
r1887 (  60 62 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=34.78 //y=7.4 //x2=35.89 //y2=7.4
r1888 (  58 932 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=33.67 //y=7.4 //x2=33.67 //y2=7.4
r1889 (  58 60 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=33.67 //y=7.4 //x2=34.78 //y2=7.4
r1890 (  56 442 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=32.19 //y=7.4 //x2=32.19 //y2=7.4
r1891 (  56 58 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=32.19 //y=7.4 //x2=33.67 //y2=7.4
r1892 (  54 432 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=31.08 //y=7.4 //x2=31.08 //y2=7.4
r1893 (  54 56 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=31.08 //y=7.4 //x2=32.19 //y2=7.4
r1894 (  52 422 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=29.97 //y=7.4 //x2=29.97 //y2=7.4
r1895 (  52 54 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=29.97 //y=7.4 //x2=31.08 //y2=7.4
r1896 (  50 926 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=28.86 //y=7.4 //x2=28.86 //y2=7.4
r1897 (  50 52 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=28.86 //y=7.4 //x2=29.97 //y2=7.4
r1898 (  48 400 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=27.38 //y=7.4 //x2=27.38 //y2=7.4
r1899 (  48 50 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=27.38 //y=7.4 //x2=28.86 //y2=7.4
r1900 (  46 390 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=26.27 //y=7.4 //x2=26.27 //y2=7.4
r1901 (  46 48 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=26.27 //y=7.4 //x2=27.38 //y2=7.4
r1902 (  44 921 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=25.16 //y=7.4 //x2=25.16 //y2=7.4
r1903 (  44 46 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=25.16 //y=7.4 //x2=26.27 //y2=7.4
r1904 (  42 368 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=7.4 //x2=23.68 //y2=7.4
r1905 (  42 44 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=23.68 //y=7.4 //x2=25.16 //y2=7.4
r1906 (  40 358 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.57 //y=7.4 //x2=22.57 //y2=7.4
r1907 (  40 42 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=22.57 //y=7.4 //x2=23.68 //y2=7.4
r1908 (  38 340 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.46 //y=7.4 //x2=21.46 //y2=7.4
r1909 (  38 40 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.46 //y=7.4 //x2=22.57 //y2=7.4
r1910 (  36 330 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=20.35 //y=7.4 //x2=20.35 //y2=7.4
r1911 (  36 38 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=20.35 //y=7.4 //x2=21.46 //y2=7.4
r1912 (  34 913 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.87 //y=7.4 //x2=18.87 //y2=7.4
r1913 (  34 36 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=18.87 //y=7.4 //x2=20.35 //y2=7.4
r1914 (  32 308 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.76 //y=7.4 //x2=17.76 //y2=7.4
r1915 (  32 34 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=17.76 //y=7.4 //x2=18.87 //y2=7.4
r1916 (  30 298 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.65 //y=7.4 //x2=16.65 //y2=7.4
r1917 (  30 32 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.65 //y=7.4 //x2=17.76 //y2=7.4
r1918 (  28 284 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=7.4 //x2=15.17 //y2=7.4
r1919 (  28 30 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=7.4 //x2=16.65 //y2=7.4
r1920 (  26 274 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=7.4 //x2=14.06 //y2=7.4
r1921 (  26 28 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=7.4 //x2=15.17 //y2=7.4
r1922 (  24 260 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=7.4 //x2=12.58 //y2=7.4
r1923 (  24 26 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=12.58 //y=7.4 //x2=14.06 //y2=7.4
r1924 (  22 250 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=7.4 //x2=11.47 //y2=7.4
r1925 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=7.4 //x2=12.58 //y2=7.4
r1926 (  20 240 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r1927 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=7.4 //x2=11.47 //y2=7.4
r1928 (  18 901 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=9.25 //y=7.4 //x2=9.25 //y2=7.4
r1929 (  18 20 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=9.25 //y=7.4 //x2=10.36 //y2=7.4
r1930 (  16 218 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=7.4 //x2=7.77 //y2=7.4
r1931 (  16 18 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=7.4 //x2=9.25 //y2=7.4
r1932 (  14 208 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r1933 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.4 //x2=7.77 //y2=7.4
r1934 (  12 198 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r1935 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.66 //y2=7.4
r1936 (  10 895 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r1937 (  10 12 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.55 //y2=7.4
r1938 (  8 176 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r1939 (  8 10 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.44 //y2=7.4
r1940 (  6 166 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r1941 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r1942 (  3 890 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r1943 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r1944 (  1 75 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=42.735 //y=7.4 //x2=43.29 //y2=7.4
r1945 (  1 72 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=42.735 //y=7.4 //x2=42.18 //y2=7.4
ends PM_TMRDFFSNQX1\%VDD

subckt PM_TMRDFFSNQX1\%noxref_3 ( 1 2 3 4 17 18 29 31 32 36 38 46 53 54 55 56 \
 57 58 59 60 61 62 63 64 66 72 73 74 75 79 80 81 82 83 85 91 92 93 94 114 116 \
 117 )
c244 ( 117 0 ) capacitor c=0.0220291f //x=1.965 //y=5.02
c245 ( 116 0 ) capacitor c=0.0217503f //x=1.085 //y=5.02
c246 ( 114 0 ) capacitor c=0.0084702f //x=1.96 //y=0.905
c247 ( 94 0 ) capacitor c=0.0556143f //x=9.525 //y=4.79
c248 ( 93 0 ) capacitor c=0.0293157f //x=9.815 //y=4.79
c249 ( 92 0 ) capacitor c=0.0347816f //x=9.48 //y=1.22
c250 ( 91 0 ) capacitor c=0.0187487f //x=9.48 //y=0.875
c251 ( 85 0 ) capacitor c=0.0137055f //x=9.325 //y=1.375
c252 ( 83 0 ) capacitor c=0.0149861f //x=9.325 //y=0.72
c253 ( 82 0 ) capacitor c=0.0965257f //x=8.95 //y=1.915
c254 ( 81 0 ) capacitor c=0.0229444f //x=8.95 //y=1.53
c255 ( 80 0 ) capacitor c=0.0234352f //x=8.95 //y=1.22
c256 ( 79 0 ) capacitor c=0.0198724f //x=8.95 //y=0.875
c257 ( 75 0 ) capacitor c=0.055995f //x=4.715 //y=4.79
c258 ( 74 0 ) capacitor c=0.0298189f //x=5.005 //y=4.79
c259 ( 73 0 ) capacitor c=0.0347816f //x=4.67 //y=1.22
c260 ( 72 0 ) capacitor c=0.0187487f //x=4.67 //y=0.875
c261 ( 66 0 ) capacitor c=0.0137055f //x=4.515 //y=1.375
c262 ( 64 0 ) capacitor c=0.0149861f //x=4.515 //y=0.72
c263 ( 63 0 ) capacitor c=0.0965245f //x=4.14 //y=1.915
c264 ( 62 0 ) capacitor c=0.0229444f //x=4.14 //y=1.53
c265 ( 61 0 ) capacitor c=0.0234352f //x=4.14 //y=1.22
c266 ( 60 0 ) capacitor c=0.0198724f //x=4.14 //y=0.875
c267 ( 59 0 ) capacitor c=0.110114f //x=9.89 //y=6.02
c268 ( 58 0 ) capacitor c=0.158956f //x=9.45 //y=6.02
c269 ( 57 0 ) capacitor c=0.110114f //x=5.08 //y=6.02
c270 ( 56 0 ) capacitor c=0.158956f //x=4.64 //y=6.02
c271 ( 53 0 ) capacitor c=0.0023043f //x=2.11 //y=5.2
c272 ( 46 0 ) capacitor c=0.100197f //x=9.25 //y=2.08
c273 ( 38 0 ) capacitor c=0.104868f //x=4.44 //y=2.08
c274 ( 36 0 ) capacitor c=0.110973f //x=2.59 //y=2.59
c275 ( 32 0 ) capacitor c=0.00468667f //x=2.235 //y=1.655
c276 ( 31 0 ) capacitor c=0.013082f //x=2.505 //y=1.655
c277 ( 29 0 ) capacitor c=0.0140934f //x=2.505 //y=5.2
c278 ( 18 0 ) capacitor c=0.00295092f //x=1.315 //y=5.2
c279 ( 17 0 ) capacitor c=0.0162034f //x=2.025 //y=5.2
c280 ( 4 0 ) capacitor c=0.00988709f //x=4.705 //y=2.59
c281 ( 3 0 ) capacitor c=0.110983f //x=9.135 //y=2.59
c282 ( 2 0 ) capacitor c=0.0138866f //x=2.705 //y=2.59
c283 ( 1 0 ) capacitor c=0.0386784f //x=4.295 //y=2.59
r284 (  93 95 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=9.815 //y=4.79 //x2=9.89 //y2=4.865
r285 (  93 94 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=9.815 //y=4.79 //x2=9.525 //y2=4.79
r286 (  92 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.48 //y=1.22 //x2=9.44 //y2=1.375
r287 (  91 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.48 //y=0.875 //x2=9.44 //y2=0.72
r288 (  91 92 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=9.48 //y=0.875 //x2=9.48 //y2=1.22
r289 (  88 94 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=9.45 //y=4.865 //x2=9.525 //y2=4.79
r290 (  88 111 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=9.45 //y=4.865 //x2=9.25 //y2=4.7
r291 (  86 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.105 //y=1.375 //x2=8.99 //y2=1.375
r292 (  85 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.325 //y=1.375 //x2=9.44 //y2=1.375
r293 (  84 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.105 //y=0.72 //x2=8.99 //y2=0.72
r294 (  83 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=9.325 //y=0.72 //x2=9.44 //y2=0.72
r295 (  83 84 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=9.325 //y=0.72 //x2=9.105 //y2=0.72
r296 (  82 109 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.915 //x2=9.25 //y2=2.08
r297 (  81 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.53 //x2=8.99 //y2=1.375
r298 (  81 82 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.53 //x2=8.95 //y2=1.915
r299 (  80 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.95 //y=1.22 //x2=8.99 //y2=1.375
r300 (  79 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.95 //y=0.875 //x2=8.99 //y2=0.72
r301 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.95 //y=0.875 //x2=8.95 //y2=1.22
r302 (  74 76 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.005 //y=4.79 //x2=5.08 //y2=4.865
r303 (  74 75 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=5.005 //y=4.79 //x2=4.715 //y2=4.79
r304 (  73 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.67 //y=1.22 //x2=4.63 //y2=1.375
r305 (  72 104 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.67 //y=0.875 //x2=4.63 //y2=0.72
r306 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.67 //y=0.875 //x2=4.67 //y2=1.22
r307 (  69 75 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.64 //y=4.865 //x2=4.715 //y2=4.79
r308 (  69 103 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=4.64 //y=4.865 //x2=4.44 //y2=4.7
r309 (  67 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.295 //y=1.375 //x2=4.18 //y2=1.375
r310 (  66 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.515 //y=1.375 //x2=4.63 //y2=1.375
r311 (  65 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.295 //y=0.72 //x2=4.18 //y2=0.72
r312 (  64 104 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.515 //y=0.72 //x2=4.63 //y2=0.72
r313 (  64 65 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.515 //y=0.72 //x2=4.295 //y2=0.72
r314 (  63 101 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.915 //x2=4.44 //y2=2.08
r315 (  62 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.53 //x2=4.18 //y2=1.375
r316 (  62 63 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.53 //x2=4.14 //y2=1.915
r317 (  61 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.14 //y=1.22 //x2=4.18 //y2=1.375
r318 (  60 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.14 //y=0.875 //x2=4.18 //y2=0.72
r319 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.14 //y=0.875 //x2=4.14 //y2=1.22
r320 (  59 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.89 //y=6.02 //x2=9.89 //y2=4.865
r321 (  58 88 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=9.45 //y=6.02 //x2=9.45 //y2=4.865
r322 (  57 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.08 //y=6.02 //x2=5.08 //y2=4.865
r323 (  56 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.64 //y=6.02 //x2=4.64 //y2=4.865
r324 (  55 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.215 //y=1.375 //x2=9.325 //y2=1.375
r325 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=9.215 //y=1.375 //x2=9.105 //y2=1.375
r326 (  54 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.405 //y=1.375 //x2=4.515 //y2=1.375
r327 (  54 67 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.405 //y=1.375 //x2=4.295 //y2=1.375
r328 (  51 111 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=4.7 //x2=9.25 //y2=4.7
r329 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=9.25 //y=2.59 //x2=9.25 //y2=4.7
r330 (  46 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=9.25 //y=2.08 //x2=9.25 //y2=2.08
r331 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=9.25 //y=2.08 //x2=9.25 //y2=2.59
r332 (  43 103 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=4.7 //x2=4.44 //y2=4.7
r333 (  41 43 ) resistor r=144.77 //w=0.187 //l=2.115 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.585 //x2=4.44 //y2=4.7
r334 (  38 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.44 //y=2.08 //x2=4.44 //y2=2.08
r335 (  38 41 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=4.44 //y=2.08 //x2=4.44 //y2=2.585
r336 (  34 36 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=2.59 //y=5.115 //x2=2.59 //y2=2.59
r337 (  33 36 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=2.59 //y=1.74 //x2=2.59 //y2=2.59
r338 (  31 33 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.59 //y2=1.74
r339 (  31 32 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.235 //y2=1.655
r340 (  30 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.195 //y=5.2 //x2=2.11 //y2=5.2
r341 (  29 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.59 //y2=5.115
r342 (  29 30 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.2 //x2=2.195 //y2=5.2
r343 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.235 //y2=1.655
r344 (  25 114 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r345 (  19 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.2
r346 (  19 117 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.285 //x2=2.11 //y2=5.725
r347 (  17 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=2.11 //y2=5.2
r348 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.025 //y=5.2 //x2=1.315 //y2=5.2
r349 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.315 //y2=5.2
r350 (  11 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=1.23 //y=5.285 //x2=1.23 //y2=5.725
r351 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=9.25 //y=2.59 //x2=9.25 //y2=2.59
r352 (  8 41 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.44 //y=2.585 //x2=4.44 //y2=2.585
r353 (  6 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.59 //y=2.59 //x2=2.59 //y2=2.59
r354 (  4 8 ) resistor r=0.164988 //w=0.206 //l=0.267488 //layer=m1 \
 //thickness=0.36 //x=4.705 //y=2.59 //x2=4.44 //y2=2.585
r355 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=9.135 //y=2.59 //x2=9.25 //y2=2.59
r356 (  3 4 ) resistor r=4.2271 //w=0.131 //l=4.43 //layer=m1 //thickness=0.36 \
 //x=9.135 //y=2.59 //x2=4.705 //y2=2.59
r357 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.705 //y=2.59 //x2=2.59 //y2=2.59
r358 (  1 8 ) resistor r=0.0921728 //w=0.206 //l=0.147479 //layer=m1 \
 //thickness=0.36 //x=4.295 //y=2.59 //x2=4.44 //y2=2.585
r359 (  1 2 ) resistor r=1.51718 //w=0.131 //l=1.59 //layer=m1 \
 //thickness=0.36 //x=4.295 //y=2.59 //x2=2.705 //y2=2.59
ends PM_TMRDFFSNQX1\%noxref_3

subckt PM_TMRDFFSNQX1\%noxref_4 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 \
 54 55 56 57 61 63 66 67 77 80 82 83 84 )
c164 ( 84 0 ) capacitor c=0.023087f //x=11.285 //y=5.02
c165 ( 83 0 ) capacitor c=0.023519f //x=10.405 //y=5.02
c166 ( 82 0 ) capacitor c=0.0224735f //x=9.525 //y=5.02
c167 ( 80 0 ) capacitor c=0.00872971f //x=11.535 //y=0.915
c168 ( 77 0 ) capacitor c=0.0588816f //x=14.06 //y=4.7
c169 ( 67 0 ) capacitor c=0.0318948f //x=14.395 //y=1.21
c170 ( 66 0 ) capacitor c=0.0187384f //x=14.395 //y=0.865
c171 ( 63 0 ) capacitor c=0.0141798f //x=14.24 //y=1.365
c172 ( 61 0 ) capacitor c=0.0149844f //x=14.24 //y=0.71
c173 ( 57 0 ) capacitor c=0.0813322f //x=13.865 //y=1.915
c174 ( 56 0 ) capacitor c=0.0229267f //x=13.865 //y=1.52
c175 ( 55 0 ) capacitor c=0.0234352f //x=13.865 //y=1.21
c176 ( 54 0 ) capacitor c=0.0199343f //x=13.865 //y=0.865
c177 ( 53 0 ) capacitor c=0.110275f //x=14.4 //y=6.02
c178 ( 52 0 ) capacitor c=0.154305f //x=13.96 //y=6.02
c179 ( 50 0 ) capacitor c=0.00106608f //x=11.43 //y=5.155
c180 ( 49 0 ) capacitor c=0.00207319f //x=10.55 //y=5.155
c181 ( 42 0 ) capacitor c=0.0869732f //x=14.06 //y=2.08
c182 ( 40 0 ) capacitor c=0.107064f //x=12.21 //y=2.59
c183 ( 36 0 ) capacitor c=0.00398962f //x=11.81 //y=1.665
c184 ( 35 0 ) capacitor c=0.0137288f //x=12.125 //y=1.665
c185 ( 29 0 ) capacitor c=0.0284988f //x=12.125 //y=5.155
c186 ( 21 0 ) capacitor c=0.0176454f //x=11.345 //y=5.155
c187 ( 14 0 ) capacitor c=0.00332903f //x=9.755 //y=5.155
c188 ( 13 0 ) capacitor c=0.0148427f //x=10.465 //y=5.155
c189 ( 2 0 ) capacitor c=0.00808366f //x=12.325 //y=2.59
c190 ( 1 0 ) capacitor c=0.0353429f //x=13.945 //y=2.59
r191 (  75 77 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=13.96 //y=4.7 //x2=14.06 //y2=4.7
r192 (  68 77 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=14.4 //y=4.865 //x2=14.06 //y2=4.7
r193 (  67 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.395 //y=1.21 //x2=14.355 //y2=1.365
r194 (  66 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.395 //y=0.865 //x2=14.355 //y2=0.71
r195 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.395 //y=0.865 //x2=14.395 //y2=1.21
r196 (  64 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.02 //y=1.365 //x2=13.905 //y2=1.365
r197 (  63 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.24 //y=1.365 //x2=14.355 //y2=1.365
r198 (  62 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.02 //y=0.71 //x2=13.905 //y2=0.71
r199 (  61 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.24 //y=0.71 //x2=14.355 //y2=0.71
r200 (  61 62 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=14.24 //y=0.71 //x2=14.02 //y2=0.71
r201 (  58 75 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=13.96 //y=4.865 //x2=13.96 //y2=4.7
r202 (  57 72 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.915 //x2=14.06 //y2=2.08
r203 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.52 //x2=13.905 //y2=1.365
r204 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.52 //x2=13.865 //y2=1.915
r205 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.865 //y=1.21 //x2=13.905 //y2=1.365
r206 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.865 //y=0.865 //x2=13.905 //y2=0.71
r207 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.865 //y=0.865 //x2=13.865 //y2=1.21
r208 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.4 //y=6.02 //x2=14.4 //y2=4.865
r209 (  52 58 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=13.96 //y=6.02 //x2=13.96 //y2=4.865
r210 (  51 63 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.13 //y=1.365 //x2=14.24 //y2=1.365
r211 (  51 64 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.13 //y=1.365 //x2=14.02 //y2=1.365
r212 (  47 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=4.7 //x2=14.06 //y2=4.7
r213 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=14.06 //y=2.59 //x2=14.06 //y2=4.7
r214 (  42 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=2.08 //x2=14.06 //y2=2.08
r215 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=14.06 //y=2.08 //x2=14.06 //y2=2.59
r216 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=12.21 //y=5.07 //x2=12.21 //y2=2.59
r217 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=12.21 //y=1.75 //x2=12.21 //y2=2.59
r218 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.125 //y=1.665 //x2=12.21 //y2=1.75
r219 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=12.125 //y=1.665 //x2=11.81 //y2=1.665
r220 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.725 //y=1.58 //x2=11.81 //y2=1.665
r221 (  31 80 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=11.725 //y=1.58 //x2=11.725 //y2=1.01
r222 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.515 //y=5.155 //x2=11.43 //y2=5.155
r223 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.125 //y=5.155 //x2=12.21 //y2=5.07
r224 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=12.125 //y=5.155 //x2=11.515 //y2=5.155
r225 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.43 //y=5.24 //x2=11.43 //y2=5.155
r226 (  23 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.43 //y=5.24 //x2=11.43 //y2=5.725
r227 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.635 //y=5.155 //x2=10.55 //y2=5.155
r228 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.345 //y=5.155 //x2=11.43 //y2=5.155
r229 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.345 //y=5.155 //x2=10.635 //y2=5.155
r230 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.55 //y=5.24 //x2=10.55 //y2=5.155
r231 (  15 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=10.55 //y=5.24 //x2=10.55 //y2=5.725
r232 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.465 //y=5.155 //x2=10.55 //y2=5.155
r233 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=10.465 //y=5.155 //x2=9.755 //y2=5.155
r234 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=9.67 //y=5.24 //x2=9.755 //y2=5.155
r235 (  7 82 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=9.67 //y=5.24 //x2=9.67 //y2=5.725
r236 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.06 //y=2.59 //x2=14.06 //y2=2.59
r237 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.21 //y=2.59 //x2=12.21 //y2=2.59
r238 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.325 //y=2.59 //x2=12.21 //y2=2.59
r239 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=2.59 //x2=14.06 //y2=2.59
r240 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=13.945 //y=2.59 //x2=12.325 //y2=2.59
ends PM_TMRDFFSNQX1\%noxref_4

subckt PM_TMRDFFSNQX1\%noxref_5 ( 1 2 3 4 11 13 23 24 31 39 45 46 50 52 61 62 \
 64 65 67 68 69 70 71 72 73 74 75 80 82 84 90 91 92 93 94 95 99 101 104 105 \
 110 111 114 128 131 133 134 135 )
c278 ( 135 0 ) capacitor c=0.023087f //x=6.475 //y=5.02
c279 ( 134 0 ) capacitor c=0.023519f //x=5.595 //y=5.02
c280 ( 133 0 ) capacitor c=0.0224735f //x=4.715 //y=5.02
c281 ( 131 0 ) capacitor c=0.00853354f //x=6.725 //y=0.915
c282 ( 128 0 ) capacitor c=0.0588816f //x=17.39 //y=4.7
c283 ( 114 0 ) capacitor c=0.0331534f //x=1.88 //y=4.7
c284 ( 111 0 ) capacitor c=0.0279499f //x=1.85 //y=1.915
c285 ( 110 0 ) capacitor c=0.0422587f //x=1.85 //y=2.08
c286 ( 105 0 ) capacitor c=0.0318948f //x=17.725 //y=1.21
c287 ( 104 0 ) capacitor c=0.0187384f //x=17.725 //y=0.865
c288 ( 101 0 ) capacitor c=0.0141798f //x=17.57 //y=1.365
c289 ( 99 0 ) capacitor c=0.0149844f //x=17.57 //y=0.71
c290 ( 95 0 ) capacitor c=0.0813322f //x=17.195 //y=1.915
c291 ( 94 0 ) capacitor c=0.0229267f //x=17.195 //y=1.52
c292 ( 93 0 ) capacitor c=0.0234352f //x=17.195 //y=1.21
c293 ( 92 0 ) capacitor c=0.0199343f //x=17.195 //y=0.865
c294 ( 91 0 ) capacitor c=0.0429696f //x=2.415 //y=1.25
c295 ( 90 0 ) capacitor c=0.0192208f //x=2.415 //y=0.905
c296 ( 84 0 ) capacitor c=0.0158629f //x=2.26 //y=1.405
c297 ( 82 0 ) capacitor c=0.0157803f //x=2.26 //y=0.75
c298 ( 80 0 ) capacitor c=0.0299681f //x=2.255 //y=4.79
c299 ( 75 0 ) capacitor c=0.0205163f //x=1.885 //y=1.56
c300 ( 74 0 ) capacitor c=0.0168481f //x=1.885 //y=1.25
c301 ( 73 0 ) capacitor c=0.0174783f //x=1.885 //y=0.905
c302 ( 72 0 ) capacitor c=0.110275f //x=17.73 //y=6.02
c303 ( 71 0 ) capacitor c=0.154305f //x=17.29 //y=6.02
c304 ( 70 0 ) capacitor c=0.15358f //x=2.33 //y=6.02
c305 ( 69 0 ) capacitor c=0.110281f //x=1.89 //y=6.02
c306 ( 65 0 ) capacitor c=0.0755336f //x=7.397 //y=3.905
c307 ( 64 0 ) capacitor c=0.0101843f //x=7.395 //y=4.07
c308 ( 62 0 ) capacitor c=0.00106608f //x=6.62 //y=5.155
c309 ( 61 0 ) capacitor c=0.00207162f //x=5.74 //y=5.155
c310 ( 52 0 ) capacitor c=0.0887144f //x=17.39 //y=2.08
c311 ( 50 0 ) capacitor c=0.0236247f //x=7.4 //y=5.07
c312 ( 46 0 ) capacitor c=0.00431225f //x=7 //y=1.665
c313 ( 45 0 ) capacitor c=0.0141453f //x=7.315 //y=1.665
c314 ( 39 0 ) capacitor c=0.0281378f //x=7.315 //y=5.155
c315 ( 31 0 ) capacitor c=0.0176454f //x=6.535 //y=5.155
c316 ( 24 0 ) capacitor c=0.00351598f //x=4.945 //y=5.155
c317 ( 23 0 ) capacitor c=0.0154196f //x=5.655 //y=5.155
c318 ( 13 0 ) capacitor c=0.0765924f //x=1.85 //y=2.08
c319 ( 11 0 ) capacitor c=0.00453889f //x=1.85 //y=4.535
c320 ( 4 0 ) capacitor c=0.00551102f //x=7.51 //y=4.07
c321 ( 3 0 ) capacitor c=0.143514f //x=17.275 //y=4.07
c322 ( 2 0 ) capacitor c=0.0165998f //x=1.965 //y=4.07
c323 ( 1 0 ) capacitor c=0.143583f //x=7.28 //y=4.07
r324 (  126 128 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=17.29 //y=4.7 //x2=17.39 //y2=4.7
r325 (  116 117 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.79 //x2=1.88 //y2=4.865
r326 (  114 116 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.88 //y=4.7 //x2=1.88 //y2=4.79
r327 (  110 111 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r328 (  106 128 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=17.73 //y=4.865 //x2=17.39 //y2=4.7
r329 (  105 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.725 //y=1.21 //x2=17.685 //y2=1.365
r330 (  104 129 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.725 //y=0.865 //x2=17.685 //y2=0.71
r331 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.725 //y=0.865 //x2=17.725 //y2=1.21
r332 (  102 125 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.35 //y=1.365 //x2=17.235 //y2=1.365
r333 (  101 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.57 //y=1.365 //x2=17.685 //y2=1.365
r334 (  100 124 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.35 //y=0.71 //x2=17.235 //y2=0.71
r335 (  99 129 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=17.57 //y=0.71 //x2=17.685 //y2=0.71
r336 (  99 100 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=17.57 //y=0.71 //x2=17.35 //y2=0.71
r337 (  96 126 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=17.29 //y=4.865 //x2=17.29 //y2=4.7
r338 (  95 123 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.915 //x2=17.39 //y2=2.08
r339 (  94 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.52 //x2=17.235 //y2=1.365
r340 (  94 95 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.52 //x2=17.195 //y2=1.915
r341 (  93 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.195 //y=1.21 //x2=17.235 //y2=1.365
r342 (  92 124 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=17.195 //y=0.865 //x2=17.235 //y2=0.71
r343 (  92 93 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=17.195 //y=0.865 //x2=17.195 //y2=1.21
r344 (  91 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.25 //x2=2.375 //y2=1.405
r345 (  90 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r346 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.25
r347 (  85 119 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r348 (  84 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.375 //y2=1.405
r349 (  83 118 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r350 (  82 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r351 (  82 83 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r352 (  81 116 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.015 //y=4.79 //x2=1.88 //y2=4.79
r353 (  80 87 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.33 //y2=4.865
r354 (  80 81 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.79 //x2=2.015 //y2=4.79
r355 (  75 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r356 (  75 111 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r357 (  74 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.25 //x2=1.925 //y2=1.405
r358 (  73 118 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r359 (  73 74 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.25
r360 (  72 106 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.73 //y=6.02 //x2=17.73 //y2=4.865
r361 (  71 96 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=17.29 //y=6.02 //x2=17.29 //y2=4.865
r362 (  70 87 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.02 //x2=2.33 //y2=4.865
r363 (  69 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.02 //x2=1.89 //y2=4.865
r364 (  68 101 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.46 //y=1.365 //x2=17.57 //y2=1.365
r365 (  68 102 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=17.46 //y=1.365 //x2=17.35 //y2=1.365
r366 (  67 84 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r367 (  67 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r368 (  64 66 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=7.397 //y=4.07 //x2=7.397 //y2=4.235
r369 (  64 65 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=7.397 //y=4.07 //x2=7.397 //y2=3.905
r370 (  60 114 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.88 //y=4.7 //x2=1.88 //y2=4.7
r371 (  57 128 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.39 //y=4.7 //x2=17.39 //y2=4.7
r372 (  55 57 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=17.39 //y=4.07 //x2=17.39 //y2=4.7
r373 (  52 123 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=17.39 //y=2.08 //x2=17.39 //y2=2.08
r374 (  52 55 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=17.39 //y=2.08 //x2=17.39 //y2=4.07
r375 (  50 66 ) resistor r=57.1551 //w=0.187 //l=0.835 //layer=li \
 //thickness=0.1 //x=7.4 //y=5.07 //x2=7.4 //y2=4.235
r376 (  47 65 ) resistor r=147.508 //w=0.187 //l=2.155 //layer=li \
 //thickness=0.1 //x=7.4 //y=1.75 //x2=7.4 //y2=3.905
r377 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.665 //x2=7.4 //y2=1.75
r378 (  45 46 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=7.315 //y=1.665 //x2=7 //y2=1.665
r379 (  41 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.915 //y=1.58 //x2=7 //y2=1.665
r380 (  41 131 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=6.915 //y=1.58 //x2=6.915 //y2=1.01
r381 (  40 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.705 //y=5.155 //x2=6.62 //y2=5.155
r382 (  39 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.155 //x2=7.4 //y2=5.07
r383 (  39 40 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=7.315 //y=5.155 //x2=6.705 //y2=5.155
r384 (  33 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.62 //y=5.24 //x2=6.62 //y2=5.155
r385 (  33 135 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.62 //y=5.24 //x2=6.62 //y2=5.725
r386 (  32 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.825 //y=5.155 //x2=5.74 //y2=5.155
r387 (  31 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.535 //y=5.155 //x2=6.62 //y2=5.155
r388 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=6.535 //y=5.155 //x2=5.825 //y2=5.155
r389 (  25 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.74 //y=5.24 //x2=5.74 //y2=5.155
r390 (  25 134 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=5.74 //y=5.24 //x2=5.74 //y2=5.725
r391 (  23 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.655 //y=5.155 //x2=5.74 //y2=5.155
r392 (  23 24 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=5.655 //y=5.155 //x2=4.945 //y2=5.155
r393 (  17 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.86 //y=5.24 //x2=4.945 //y2=5.155
r394 (  17 133 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.86 //y=5.24 //x2=4.86 //y2=5.725
r395 (  13 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r396 (  13 16 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=1.85 //y=2.08 //x2=1.85 //y2=4.07
r397 (  11 60 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.865 //y2=4.7
r398 (  11 16 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.535 //x2=1.85 //y2=4.07
r399 (  10 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.39 //y=4.07 //x2=17.39 //y2=4.07
r400 (  8 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=7.395 //y=4.07 //x2=7.395 //y2=4.07
r401 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.85 //y=4.07 //x2=1.85 //y2=4.07
r402 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.51 //y=4.07 //x2=7.395 //y2=4.07
r403 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.275 //y=4.07 //x2=17.39 //y2=4.07
r404 (  3 4 ) resistor r=9.31775 //w=0.131 //l=9.765 //layer=m1 \
 //thickness=0.36 //x=17.275 //y=4.07 //x2=7.51 //y2=4.07
r405 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.965 //y=4.07 //x2=1.85 //y2=4.07
r406 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=7.28 //y=4.07 //x2=7.395 //y2=4.07
r407 (  1 2 ) resistor r=5.07156 //w=0.131 //l=5.315 //layer=m1 \
 //thickness=0.36 //x=7.28 //y=4.07 //x2=1.965 //y2=4.07
ends PM_TMRDFFSNQX1\%noxref_5

subckt PM_TMRDFFSNQX1\%noxref_6 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 \
 47 48 49 51 57 58 59 60 72 74 75 )
c152 ( 75 0 ) capacitor c=0.0220291f //x=18.245 //y=5.02
c153 ( 74 0 ) capacitor c=0.0217503f //x=17.365 //y=5.02
c154 ( 72 0 ) capacitor c=0.0084702f //x=18.24 //y=0.905
c155 ( 60 0 ) capacitor c=0.0556143f //x=20.995 //y=4.79
c156 ( 59 0 ) capacitor c=0.0293157f //x=21.285 //y=4.79
c157 ( 58 0 ) capacitor c=0.0347816f //x=20.95 //y=1.22
c158 ( 57 0 ) capacitor c=0.0187487f //x=20.95 //y=0.875
c159 ( 51 0 ) capacitor c=0.0137055f //x=20.795 //y=1.375
c160 ( 49 0 ) capacitor c=0.0149861f //x=20.795 //y=0.72
c161 ( 48 0 ) capacitor c=0.096037f //x=20.42 //y=1.915
c162 ( 47 0 ) capacitor c=0.0228993f //x=20.42 //y=1.53
c163 ( 46 0 ) capacitor c=0.0234352f //x=20.42 //y=1.22
c164 ( 45 0 ) capacitor c=0.0198724f //x=20.42 //y=0.875
c165 ( 44 0 ) capacitor c=0.110114f //x=21.36 //y=6.02
c166 ( 43 0 ) capacitor c=0.158956f //x=20.92 //y=6.02
c167 ( 41 0 ) capacitor c=0.00211606f //x=18.39 //y=5.2
c168 ( 34 0 ) capacitor c=0.0963459f //x=20.72 //y=2.08
c169 ( 32 0 ) capacitor c=0.104321f //x=18.87 //y=4.07
c170 ( 28 0 ) capacitor c=0.00404073f //x=18.515 //y=1.655
c171 ( 27 0 ) capacitor c=0.0122201f //x=18.785 //y=1.655
c172 ( 25 0 ) capacitor c=0.0137995f //x=18.785 //y=5.2
c173 ( 14 0 ) capacitor c=0.00251459f //x=17.595 //y=5.2
c174 ( 13 0 ) capacitor c=0.0142423f //x=18.305 //y=5.2
c175 ( 2 0 ) capacitor c=0.00645515f //x=18.985 //y=4.07
c176 ( 1 0 ) capacitor c=0.0383007f //x=20.605 //y=4.07
r177 (  59 61 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=21.285 //y=4.79 //x2=21.36 //y2=4.865
r178 (  59 60 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=21.285 //y=4.79 //x2=20.995 //y2=4.79
r179 (  58 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.95 //y=1.22 //x2=20.91 //y2=1.375
r180 (  57 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.95 //y=0.875 //x2=20.91 //y2=0.72
r181 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.95 //y=0.875 //x2=20.95 //y2=1.22
r182 (  54 60 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.92 //y=4.865 //x2=20.995 //y2=4.79
r183 (  54 69 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=20.92 //y=4.865 //x2=20.72 //y2=4.7
r184 (  52 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.575 //y=1.375 //x2=20.46 //y2=1.375
r185 (  51 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.795 //y=1.375 //x2=20.91 //y2=1.375
r186 (  50 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.575 //y=0.72 //x2=20.46 //y2=0.72
r187 (  49 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=20.795 //y=0.72 //x2=20.91 //y2=0.72
r188 (  49 50 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=20.795 //y=0.72 //x2=20.575 //y2=0.72
r189 (  48 67 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.915 //x2=20.72 //y2=2.08
r190 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.53 //x2=20.46 //y2=1.375
r191 (  47 48 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.53 //x2=20.42 //y2=1.915
r192 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.42 //y=1.22 //x2=20.46 //y2=1.375
r193 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.42 //y=0.875 //x2=20.46 //y2=0.72
r194 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=20.42 //y=0.875 //x2=20.42 //y2=1.22
r195 (  44 61 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.36 //y=6.02 //x2=21.36 //y2=4.865
r196 (  43 54 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.92 //y=6.02 //x2=20.92 //y2=4.865
r197 (  42 51 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.685 //y=1.375 //x2=20.795 //y2=1.375
r198 (  42 52 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=20.685 //y=1.375 //x2=20.575 //y2=1.375
r199 (  39 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.72 //y=4.7 //x2=20.72 //y2=4.7
r200 (  37 39 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=20.72 //y=4.07 //x2=20.72 //y2=4.7
r201 (  34 67 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=20.72 //y=2.08 //x2=20.72 //y2=2.08
r202 (  34 37 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=20.72 //y=2.08 //x2=20.72 //y2=4.07
r203 (  30 32 ) resistor r=71.5294 //w=0.187 //l=1.045 //layer=li \
 //thickness=0.1 //x=18.87 //y=5.115 //x2=18.87 //y2=4.07
r204 (  29 32 ) resistor r=159.487 //w=0.187 //l=2.33 //layer=li \
 //thickness=0.1 //x=18.87 //y=1.74 //x2=18.87 //y2=4.07
r205 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.785 //y=1.655 //x2=18.87 //y2=1.74
r206 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=18.785 //y=1.655 //x2=18.515 //y2=1.655
r207 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.475 //y=5.2 //x2=18.39 //y2=5.2
r208 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.785 //y=5.2 //x2=18.87 //y2=5.115
r209 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=18.785 //y=5.2 //x2=18.475 //y2=5.2
r210 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=18.43 //y=1.57 //x2=18.515 //y2=1.655
r211 (  21 72 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=18.43 //y=1.57 //x2=18.43 //y2=1
r212 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.39 //y=5.285 //x2=18.39 //y2=5.2
r213 (  15 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=18.39 //y=5.285 //x2=18.39 //y2=5.725
r214 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.305 //y=5.2 //x2=18.39 //y2=5.2
r215 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=18.305 //y=5.2 //x2=17.595 //y2=5.2
r216 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=17.51 //y=5.285 //x2=17.595 //y2=5.2
r217 (  7 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=17.51 //y=5.285 //x2=17.51 //y2=5.725
r218 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=20.72 //y=4.07 //x2=20.72 //y2=4.07
r219 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.87 //y=4.07 //x2=18.87 //y2=4.07
r220 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.985 //y=4.07 //x2=18.87 //y2=4.07
r221 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=20.605 //y=4.07 //x2=20.72 //y2=4.07
r222 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=20.605 //y=4.07 //x2=18.985 //y2=4.07
ends PM_TMRDFFSNQX1\%noxref_6

subckt PM_TMRDFFSNQX1\%noxref_7 ( 1 2 3 4 5 6 16 24 37 38 49 51 52 56 58 65 66 \
 67 68 69 70 71 72 73 74 78 79 80 85 87 90 91 95 96 97 102 104 107 108 112 113 \
 114 119 121 124 125 127 128 133 137 138 143 147 148 153 156 158 159 )
c322 ( 159 0 ) capacitor c=0.0220291f //x=14.915 //y=5.02
c323 ( 158 0 ) capacitor c=0.0217503f //x=14.035 //y=5.02
c324 ( 156 0 ) capacitor c=0.00866655f //x=14.91 //y=0.905
c325 ( 153 0 ) capacitor c=0.0587755f //x=22.94 //y=4.7
c326 ( 148 0 ) capacitor c=0.0273931f //x=22.94 //y=1.915
c327 ( 147 0 ) capacitor c=0.0456313f //x=22.94 //y=2.08
c328 ( 143 0 ) capacitor c=0.0587755f //x=11.47 //y=4.7
c329 ( 138 0 ) capacitor c=0.0273931f //x=11.47 //y=1.915
c330 ( 137 0 ) capacitor c=0.0456313f //x=11.47 //y=2.08
c331 ( 133 0 ) capacitor c=0.058931f //x=6.66 //y=4.7
c332 ( 128 0 ) capacitor c=0.0267105f //x=6.66 //y=1.915
c333 ( 127 0 ) capacitor c=0.0457054f //x=6.66 //y=2.08
c334 ( 125 0 ) capacitor c=0.0432517f //x=23.46 //y=1.26
c335 ( 124 0 ) capacitor c=0.0200379f //x=23.46 //y=0.915
c336 ( 121 0 ) capacitor c=0.0148873f //x=23.305 //y=1.415
c337 ( 119 0 ) capacitor c=0.0157803f //x=23.305 //y=0.76
c338 ( 114 0 ) capacitor c=0.0218028f //x=22.93 //y=1.57
c339 ( 113 0 ) capacitor c=0.0207459f //x=22.93 //y=1.26
c340 ( 112 0 ) capacitor c=0.0194308f //x=22.93 //y=0.915
c341 ( 108 0 ) capacitor c=0.0432517f //x=11.99 //y=1.26
c342 ( 107 0 ) capacitor c=0.0200379f //x=11.99 //y=0.915
c343 ( 104 0 ) capacitor c=0.0148873f //x=11.835 //y=1.415
c344 ( 102 0 ) capacitor c=0.0157803f //x=11.835 //y=0.76
c345 ( 97 0 ) capacitor c=0.0218028f //x=11.46 //y=1.57
c346 ( 96 0 ) capacitor c=0.0207459f //x=11.46 //y=1.26
c347 ( 95 0 ) capacitor c=0.0194308f //x=11.46 //y=0.915
c348 ( 91 0 ) capacitor c=0.0432517f //x=7.18 //y=1.26
c349 ( 90 0 ) capacitor c=0.0200379f //x=7.18 //y=0.915
c350 ( 87 0 ) capacitor c=0.0158629f //x=7.025 //y=1.415
c351 ( 85 0 ) capacitor c=0.0157803f //x=7.025 //y=0.76
c352 ( 80 0 ) capacitor c=0.0218028f //x=6.65 //y=1.57
c353 ( 79 0 ) capacitor c=0.0207459f //x=6.65 //y=1.26
c354 ( 78 0 ) capacitor c=0.0194308f //x=6.65 //y=0.915
c355 ( 74 0 ) capacitor c=0.158794f //x=23.12 //y=6.02
c356 ( 73 0 ) capacitor c=0.110114f //x=22.68 //y=6.02
c357 ( 72 0 ) capacitor c=0.158794f //x=11.65 //y=6.02
c358 ( 71 0 ) capacitor c=0.110114f //x=11.21 //y=6.02
c359 ( 70 0 ) capacitor c=0.158048f //x=6.84 //y=6.02
c360 ( 69 0 ) capacitor c=0.110114f //x=6.4 //y=6.02
c361 ( 65 0 ) capacitor c=0.00211606f //x=15.06 //y=5.2
c362 ( 58 0 ) capacitor c=0.0839891f //x=22.94 //y=2.08
c363 ( 56 0 ) capacitor c=0.10649f //x=15.54 //y=3.7
c364 ( 52 0 ) capacitor c=0.00404073f //x=15.185 //y=1.655
c365 ( 51 0 ) capacitor c=0.0122201f //x=15.455 //y=1.655
c366 ( 49 0 ) capacitor c=0.0137522f //x=15.455 //y=5.2
c367 ( 38 0 ) capacitor c=0.00251635f //x=14.265 //y=5.2
c368 ( 37 0 ) capacitor c=0.0142529f //x=14.975 //y=5.2
c369 ( 24 0 ) capacitor c=0.0834768f //x=11.47 //y=2.08
c370 ( 16 0 ) capacitor c=0.0842778f //x=6.66 //y=2.08
c371 ( 6 0 ) capacitor c=0.0043044f //x=15.655 //y=3.7
c372 ( 5 0 ) capacitor c=0.13532f //x=22.825 //y=3.7
c373 ( 4 0 ) capacitor c=0.00443912f //x=11.585 //y=3.7
c374 ( 3 0 ) capacitor c=0.0668348f //x=15.425 //y=3.7
c375 ( 2 0 ) capacitor c=0.0143354f //x=6.775 //y=3.7
c376 ( 1 0 ) capacitor c=0.0815699f //x=11.355 //y=3.7
r377 (  147 148 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=22.94 //y=2.08 //x2=22.94 //y2=1.915
r378 (  137 138 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=11.47 //y=2.08 //x2=11.47 //y2=1.915
r379 (  127 128 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=6.66 //y=2.08 //x2=6.66 //y2=1.915
r380 (  125 155 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.46 //y=1.26 //x2=23.42 //y2=1.415
r381 (  124 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.46 //y=0.915 //x2=23.42 //y2=0.76
r382 (  124 125 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=23.46 //y=0.915 //x2=23.46 //y2=1.26
r383 (  122 151 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.085 //y=1.415 //x2=22.97 //y2=1.415
r384 (  121 155 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.305 //y=1.415 //x2=23.42 //y2=1.415
r385 (  120 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.085 //y=0.76 //x2=22.97 //y2=0.76
r386 (  119 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.305 //y=0.76 //x2=23.42 //y2=0.76
r387 (  119 120 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=23.305 //y=0.76 //x2=23.085 //y2=0.76
r388 (  116 153 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=23.12 //y=4.865 //x2=22.94 //y2=4.7
r389 (  114 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.93 //y=1.57 //x2=22.97 //y2=1.415
r390 (  114 148 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.93 //y=1.57 //x2=22.93 //y2=1.915
r391 (  113 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.93 //y=1.26 //x2=22.97 //y2=1.415
r392 (  112 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=22.93 //y=0.915 //x2=22.97 //y2=0.76
r393 (  112 113 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=22.93 //y=0.915 //x2=22.93 //y2=1.26
r394 (  109 153 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=22.68 //y=4.865 //x2=22.94 //y2=4.7
r395 (  108 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.99 //y=1.26 //x2=11.95 //y2=1.415
r396 (  107 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.99 //y=0.915 //x2=11.95 //y2=0.76
r397 (  107 108 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.99 //y=0.915 //x2=11.99 //y2=1.26
r398 (  105 141 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.615 //y=1.415 //x2=11.5 //y2=1.415
r399 (  104 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.835 //y=1.415 //x2=11.95 //y2=1.415
r400 (  103 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.615 //y=0.76 //x2=11.5 //y2=0.76
r401 (  102 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.835 //y=0.76 //x2=11.95 //y2=0.76
r402 (  102 103 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=11.835 //y=0.76 //x2=11.615 //y2=0.76
r403 (  99 143 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=11.65 //y=4.865 //x2=11.47 //y2=4.7
r404 (  97 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.46 //y=1.57 //x2=11.5 //y2=1.415
r405 (  97 138 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.46 //y=1.57 //x2=11.46 //y2=1.915
r406 (  96 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.46 //y=1.26 //x2=11.5 //y2=1.415
r407 (  95 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.46 //y=0.915 //x2=11.5 //y2=0.76
r408 (  95 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.46 //y=0.915 //x2=11.46 //y2=1.26
r409 (  92 143 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=11.21 //y=4.865 //x2=11.47 //y2=4.7
r410 (  91 135 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.18 //y=1.26 //x2=7.14 //y2=1.415
r411 (  90 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.18 //y=0.915 //x2=7.14 //y2=0.76
r412 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=7.18 //y=0.915 //x2=7.18 //y2=1.26
r413 (  88 131 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.805 //y=1.415 //x2=6.69 //y2=1.415
r414 (  87 135 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.025 //y=1.415 //x2=7.14 //y2=1.415
r415 (  86 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.805 //y=0.76 //x2=6.69 //y2=0.76
r416 (  85 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=7.025 //y=0.76 //x2=7.14 //y2=0.76
r417 (  85 86 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=7.025 //y=0.76 //x2=6.805 //y2=0.76
r418 (  82 133 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=6.84 //y=4.865 //x2=6.66 //y2=4.7
r419 (  80 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.65 //y=1.57 //x2=6.69 //y2=1.415
r420 (  80 128 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.65 //y=1.57 //x2=6.65 //y2=1.915
r421 (  79 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.65 //y=1.26 //x2=6.69 //y2=1.415
r422 (  78 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.65 //y=0.915 //x2=6.69 //y2=0.76
r423 (  78 79 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.65 //y=0.915 //x2=6.65 //y2=1.26
r424 (  75 133 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=6.4 //y=4.865 //x2=6.66 //y2=4.7
r425 (  74 116 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=23.12 //y=6.02 //x2=23.12 //y2=4.865
r426 (  73 109 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.68 //y=6.02 //x2=22.68 //y2=4.865
r427 (  72 99 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.65 //y=6.02 //x2=11.65 //y2=4.865
r428 (  71 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.21 //y=6.02 //x2=11.21 //y2=4.865
r429 (  70 82 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.84 //y=6.02 //x2=6.84 //y2=4.865
r430 (  69 75 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.4 //y=6.02 //x2=6.4 //y2=4.865
r431 (  68 121 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.195 //y=1.415 //x2=23.305 //y2=1.415
r432 (  68 122 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.195 //y=1.415 //x2=23.085 //y2=1.415
r433 (  67 104 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.725 //y=1.415 //x2=11.835 //y2=1.415
r434 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.725 //y=1.415 //x2=11.615 //y2=1.415
r435 (  66 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.915 //y=1.415 //x2=7.025 //y2=1.415
r436 (  66 88 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=6.915 //y=1.415 //x2=6.805 //y2=1.415
r437 (  63 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.94 //y=4.7 //x2=22.94 //y2=4.7
r438 (  61 63 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=22.94 //y=3.7 //x2=22.94 //y2=4.7
r439 (  58 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=22.94 //y=2.08 //x2=22.94 //y2=2.08
r440 (  58 61 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=22.94 //y=2.08 //x2=22.94 //y2=3.7
r441 (  54 56 ) resistor r=96.8556 //w=0.187 //l=1.415 //layer=li \
 //thickness=0.1 //x=15.54 //y=5.115 //x2=15.54 //y2=3.7
r442 (  53 56 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=15.54 //y=1.74 //x2=15.54 //y2=3.7
r443 (  51 53 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.455 //y=1.655 //x2=15.54 //y2=1.74
r444 (  51 52 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=15.455 //y=1.655 //x2=15.185 //y2=1.655
r445 (  50 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.145 //y=5.2 //x2=15.06 //y2=5.2
r446 (  49 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.455 //y=5.2 //x2=15.54 //y2=5.115
r447 (  49 50 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=15.455 //y=5.2 //x2=15.145 //y2=5.2
r448 (  45 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=15.1 //y=1.57 //x2=15.185 //y2=1.655
r449 (  45 156 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=15.1 //y=1.57 //x2=15.1 //y2=1
r450 (  39 65 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.06 //y=5.285 //x2=15.06 //y2=5.2
r451 (  39 159 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=15.06 //y=5.285 //x2=15.06 //y2=5.725
r452 (  37 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.975 //y=5.2 //x2=15.06 //y2=5.2
r453 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=14.975 //y=5.2 //x2=14.265 //y2=5.2
r454 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.18 //y=5.285 //x2=14.265 //y2=5.2
r455 (  31 158 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=14.18 //y=5.285 //x2=14.18 //y2=5.725
r456 (  29 143 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.47 //y=4.7 //x2=11.47 //y2=4.7
r457 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=11.47 //y=3.7 //x2=11.47 //y2=4.7
r458 (  24 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.47 //y=2.08 //x2=11.47 //y2=2.08
r459 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=11.47 //y=2.08 //x2=11.47 //y2=3.7
r460 (  21 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=4.7 //x2=6.66 //y2=4.7
r461 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=6.66 //y=3.7 //x2=6.66 //y2=4.7
r462 (  16 127 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=6.66 //y=2.08 //x2=6.66 //y2=2.08
r463 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=6.66 //y=2.08 //x2=6.66 //y2=3.7
r464 (  14 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=22.94 //y=3.7 //x2=22.94 //y2=3.7
r465 (  12 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.54 //y=3.7 //x2=15.54 //y2=3.7
r466 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.47 //y=3.7 //x2=11.47 //y2=3.7
r467 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=6.66 //y=3.7 //x2=6.66 //y2=3.7
r468 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.655 //y=3.7 //x2=15.54 //y2=3.7
r469 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=22.825 //y=3.7 //x2=22.94 //y2=3.7
r470 (  5 6 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=22.825 //y=3.7 //x2=15.655 //y2=3.7
r471 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.585 //y=3.7 //x2=11.47 //y2=3.7
r472 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.425 //y=3.7 //x2=15.54 //y2=3.7
r473 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=15.425 //y=3.7 //x2=11.585 //y2=3.7
r474 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.775 //y=3.7 //x2=6.66 //y2=3.7
r475 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.355 //y=3.7 //x2=11.47 //y2=3.7
r476 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=11.355 //y=3.7 //x2=6.775 //y2=3.7
ends PM_TMRDFFSNQX1\%noxref_7

subckt PM_TMRDFFSNQX1\%noxref_8 ( 1 2 3 4 17 18 29 31 32 36 38 46 53 54 55 56 \
 57 58 59 60 61 62 63 64 66 72 73 74 75 79 80 81 82 83 85 91 92 93 94 114 116 \
 117 )
c232 ( 117 0 ) capacitor c=0.0220291f //x=26.385 //y=5.02
c233 ( 116 0 ) capacitor c=0.0217503f //x=25.505 //y=5.02
c234 ( 114 0 ) capacitor c=0.0084702f //x=26.38 //y=0.905
c235 ( 94 0 ) capacitor c=0.0556143f //x=33.945 //y=4.79
c236 ( 93 0 ) capacitor c=0.0293157f //x=34.235 //y=4.79
c237 ( 92 0 ) capacitor c=0.0347816f //x=33.9 //y=1.22
c238 ( 91 0 ) capacitor c=0.0187487f //x=33.9 //y=0.875
c239 ( 85 0 ) capacitor c=0.0137055f //x=33.745 //y=1.375
c240 ( 83 0 ) capacitor c=0.0149861f //x=33.745 //y=0.72
c241 ( 82 0 ) capacitor c=0.096037f //x=33.37 //y=1.915
c242 ( 81 0 ) capacitor c=0.0228993f //x=33.37 //y=1.53
c243 ( 80 0 ) capacitor c=0.0234352f //x=33.37 //y=1.22
c244 ( 79 0 ) capacitor c=0.0198724f //x=33.37 //y=0.875
c245 ( 75 0 ) capacitor c=0.0557698f //x=29.135 //y=4.79
c246 ( 74 0 ) capacitor c=0.0293157f //x=29.425 //y=4.79
c247 ( 73 0 ) capacitor c=0.0347816f //x=29.09 //y=1.22
c248 ( 72 0 ) capacitor c=0.0187487f //x=29.09 //y=0.875
c249 ( 66 0 ) capacitor c=0.0137055f //x=28.935 //y=1.375
c250 ( 64 0 ) capacitor c=0.0149861f //x=28.935 //y=0.72
c251 ( 63 0 ) capacitor c=0.096037f //x=28.56 //y=1.915
c252 ( 62 0 ) capacitor c=0.0228993f //x=28.56 //y=1.53
c253 ( 61 0 ) capacitor c=0.0234352f //x=28.56 //y=1.22
c254 ( 60 0 ) capacitor c=0.0198724f //x=28.56 //y=0.875
c255 ( 59 0 ) capacitor c=0.110114f //x=34.31 //y=6.02
c256 ( 58 0 ) capacitor c=0.158956f //x=33.87 //y=6.02
c257 ( 57 0 ) capacitor c=0.110114f //x=29.5 //y=6.02
c258 ( 56 0 ) capacitor c=0.158956f //x=29.06 //y=6.02
c259 ( 53 0 ) capacitor c=0.00211606f //x=26.53 //y=5.2
c260 ( 46 0 ) capacitor c=0.0943831f //x=33.67 //y=2.08
c261 ( 38 0 ) capacitor c=0.0969522f //x=28.86 //y=2.08
c262 ( 36 0 ) capacitor c=0.105101f //x=27.01 //y=2.59
c263 ( 32 0 ) capacitor c=0.00404073f //x=26.655 //y=1.655
c264 ( 31 0 ) capacitor c=0.0122201f //x=26.925 //y=1.655
c265 ( 29 0 ) capacitor c=0.0137995f //x=26.925 //y=5.2
c266 ( 18 0 ) capacitor c=0.00251635f //x=25.735 //y=5.2
c267 ( 17 0 ) capacitor c=0.0143649f //x=26.445 //y=5.2
c268 ( 4 0 ) capacitor c=0.00673266f //x=29.125 //y=2.59
c269 ( 3 0 ) capacitor c=0.0686809f //x=33.555 //y=2.59
c270 ( 2 0 ) capacitor c=0.0121637f //x=27.125 //y=2.59
c271 ( 1 0 ) capacitor c=0.0230071f //x=28.715 //y=2.59
r272 (  93 95 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=34.235 //y=4.79 //x2=34.31 //y2=4.865
r273 (  93 94 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=34.235 //y=4.79 //x2=33.945 //y2=4.79
r274 (  92 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.9 //y=1.22 //x2=33.86 //y2=1.375
r275 (  91 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.9 //y=0.875 //x2=33.86 //y2=0.72
r276 (  91 92 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=33.9 //y=0.875 //x2=33.9 //y2=1.22
r277 (  88 94 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=33.87 //y=4.865 //x2=33.945 //y2=4.79
r278 (  88 111 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=33.87 //y=4.865 //x2=33.67 //y2=4.7
r279 (  86 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=33.525 //y=1.375 //x2=33.41 //y2=1.375
r280 (  85 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=33.745 //y=1.375 //x2=33.86 //y2=1.375
r281 (  84 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=33.525 //y=0.72 //x2=33.41 //y2=0.72
r282 (  83 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=33.745 //y=0.72 //x2=33.86 //y2=0.72
r283 (  83 84 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=33.745 //y=0.72 //x2=33.525 //y2=0.72
r284 (  82 109 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=33.37 //y=1.915 //x2=33.67 //y2=2.08
r285 (  81 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.37 //y=1.53 //x2=33.41 //y2=1.375
r286 (  81 82 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=33.37 //y=1.53 //x2=33.37 //y2=1.915
r287 (  80 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.37 //y=1.22 //x2=33.41 //y2=1.375
r288 (  79 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=33.37 //y=0.875 //x2=33.41 //y2=0.72
r289 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=33.37 //y=0.875 //x2=33.37 //y2=1.22
r290 (  74 76 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=29.425 //y=4.79 //x2=29.5 //y2=4.865
r291 (  74 75 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=29.425 //y=4.79 //x2=29.135 //y2=4.79
r292 (  73 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.09 //y=1.22 //x2=29.05 //y2=1.375
r293 (  72 104 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.09 //y=0.875 //x2=29.05 //y2=0.72
r294 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=29.09 //y=0.875 //x2=29.09 //y2=1.22
r295 (  69 75 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=29.06 //y=4.865 //x2=29.135 //y2=4.79
r296 (  69 103 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=29.06 //y=4.865 //x2=28.86 //y2=4.7
r297 (  67 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.715 //y=1.375 //x2=28.6 //y2=1.375
r298 (  66 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.935 //y=1.375 //x2=29.05 //y2=1.375
r299 (  65 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.715 //y=0.72 //x2=28.6 //y2=0.72
r300 (  64 104 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=28.935 //y=0.72 //x2=29.05 //y2=0.72
r301 (  64 65 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=28.935 //y=0.72 //x2=28.715 //y2=0.72
r302 (  63 101 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=28.56 //y=1.915 //x2=28.86 //y2=2.08
r303 (  62 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.56 //y=1.53 //x2=28.6 //y2=1.375
r304 (  62 63 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=28.56 //y=1.53 //x2=28.56 //y2=1.915
r305 (  61 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.56 //y=1.22 //x2=28.6 //y2=1.375
r306 (  60 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=28.56 //y=0.875 //x2=28.6 //y2=0.72
r307 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=28.56 //y=0.875 //x2=28.56 //y2=1.22
r308 (  59 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=34.31 //y=6.02 //x2=34.31 //y2=4.865
r309 (  58 88 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=33.87 //y=6.02 //x2=33.87 //y2=4.865
r310 (  57 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=29.5 //y=6.02 //x2=29.5 //y2=4.865
r311 (  56 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=29.06 //y=6.02 //x2=29.06 //y2=4.865
r312 (  55 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=33.635 //y=1.375 //x2=33.745 //y2=1.375
r313 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=33.635 //y=1.375 //x2=33.525 //y2=1.375
r314 (  54 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=28.825 //y=1.375 //x2=28.935 //y2=1.375
r315 (  54 67 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=28.825 //y=1.375 //x2=28.715 //y2=1.375
r316 (  51 111 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=33.67 //y=4.7 //x2=33.67 //y2=4.7
r317 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=33.67 //y=2.59 //x2=33.67 //y2=4.7
r318 (  46 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=33.67 //y=2.08 //x2=33.67 //y2=2.08
r319 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=33.67 //y=2.08 //x2=33.67 //y2=2.59
r320 (  43 103 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=28.86 //y=4.7 //x2=28.86 //y2=4.7
r321 (  41 43 ) resistor r=144.77 //w=0.187 //l=2.115 //layer=li \
 //thickness=0.1 //x=28.86 //y=2.585 //x2=28.86 //y2=4.7
r322 (  38 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=28.86 //y=2.08 //x2=28.86 //y2=2.08
r323 (  38 41 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=28.86 //y=2.08 //x2=28.86 //y2=2.585
r324 (  34 36 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=27.01 //y=5.115 //x2=27.01 //y2=2.59
r325 (  33 36 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=27.01 //y=1.74 //x2=27.01 //y2=2.59
r326 (  31 33 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=26.925 //y=1.655 //x2=27.01 //y2=1.74
r327 (  31 32 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=26.925 //y=1.655 //x2=26.655 //y2=1.655
r328 (  30 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.615 //y=5.2 //x2=26.53 //y2=5.2
r329 (  29 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=26.925 //y=5.2 //x2=27.01 //y2=5.115
r330 (  29 30 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=26.925 //y=5.2 //x2=26.615 //y2=5.2
r331 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=26.57 //y=1.57 //x2=26.655 //y2=1.655
r332 (  25 114 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=26.57 //y=1.57 //x2=26.57 //y2=1
r333 (  19 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.53 //y=5.285 //x2=26.53 //y2=5.2
r334 (  19 117 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=26.53 //y=5.285 //x2=26.53 //y2=5.725
r335 (  17 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=26.445 //y=5.2 //x2=26.53 //y2=5.2
r336 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=26.445 //y=5.2 //x2=25.735 //y2=5.2
r337 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.65 //y=5.285 //x2=25.735 //y2=5.2
r338 (  11 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=25.65 //y=5.285 //x2=25.65 //y2=5.725
r339 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=33.67 //y=2.59 //x2=33.67 //y2=2.59
r340 (  8 41 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=28.86 //y=2.585 //x2=28.86 //y2=2.585
r341 (  6 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=27.01 //y=2.59 //x2=27.01 //y2=2.59
r342 (  4 8 ) resistor r=0.164988 //w=0.206 //l=0.267488 //layer=m1 \
 //thickness=0.36 //x=29.125 //y=2.59 //x2=28.86 //y2=2.585
r343 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=33.555 //y=2.59 //x2=33.67 //y2=2.59
r344 (  3 4 ) resistor r=4.2271 //w=0.131 //l=4.43 //layer=m1 //thickness=0.36 \
 //x=33.555 //y=2.59 //x2=29.125 //y2=2.59
r345 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=27.125 //y=2.59 //x2=27.01 //y2=2.59
r346 (  1 8 ) resistor r=0.0921728 //w=0.206 //l=0.147479 //layer=m1 \
 //thickness=0.36 //x=28.715 //y=2.59 //x2=28.86 //y2=2.585
r347 (  1 2 ) resistor r=1.51718 //w=0.131 //l=1.59 //layer=m1 \
 //thickness=0.36 //x=28.715 //y=2.59 //x2=27.125 //y2=2.59
ends PM_TMRDFFSNQX1\%noxref_8

subckt PM_TMRDFFSNQX1\%noxref_9 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 \
 54 55 56 57 61 63 66 67 77 80 82 83 84 )
c166 ( 84 0 ) capacitor c=0.023087f //x=35.705 //y=5.02
c167 ( 83 0 ) capacitor c=0.023519f //x=34.825 //y=5.02
c168 ( 82 0 ) capacitor c=0.0224735f //x=33.945 //y=5.02
c169 ( 80 0 ) capacitor c=0.00872971f //x=35.955 //y=0.915
c170 ( 77 0 ) capacitor c=0.0588816f //x=38.48 //y=4.7
c171 ( 67 0 ) capacitor c=0.0318948f //x=38.815 //y=1.21
c172 ( 66 0 ) capacitor c=0.0187384f //x=38.815 //y=0.865
c173 ( 63 0 ) capacitor c=0.0141798f //x=38.66 //y=1.365
c174 ( 61 0 ) capacitor c=0.0149844f //x=38.66 //y=0.71
c175 ( 57 0 ) capacitor c=0.0813322f //x=38.285 //y=1.915
c176 ( 56 0 ) capacitor c=0.0229267f //x=38.285 //y=1.52
c177 ( 55 0 ) capacitor c=0.0234352f //x=38.285 //y=1.21
c178 ( 54 0 ) capacitor c=0.0199343f //x=38.285 //y=0.865
c179 ( 53 0 ) capacitor c=0.110275f //x=38.82 //y=6.02
c180 ( 52 0 ) capacitor c=0.154305f //x=38.38 //y=6.02
c181 ( 50 0 ) capacitor c=0.00106608f //x=35.85 //y=5.155
c182 ( 49 0 ) capacitor c=0.00207319f //x=34.97 //y=5.155
c183 ( 42 0 ) capacitor c=0.0839295f //x=38.48 //y=2.08
c184 ( 40 0 ) capacitor c=0.10402f //x=36.63 //y=2.59
c185 ( 36 0 ) capacitor c=0.00398962f //x=36.23 //y=1.665
c186 ( 35 0 ) capacitor c=0.0137288f //x=36.545 //y=1.665
c187 ( 29 0 ) capacitor c=0.0284988f //x=36.545 //y=5.155
c188 ( 21 0 ) capacitor c=0.0176454f //x=35.765 //y=5.155
c189 ( 14 0 ) capacitor c=0.00332903f //x=34.175 //y=5.155
c190 ( 13 0 ) capacitor c=0.0148427f //x=34.885 //y=5.155
c191 ( 2 0 ) capacitor c=0.00808366f //x=36.745 //y=2.59
c192 ( 1 0 ) capacitor c=0.0353429f //x=38.365 //y=2.59
r193 (  75 77 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=38.38 //y=4.7 //x2=38.48 //y2=4.7
r194 (  68 77 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=38.82 //y=4.865 //x2=38.48 //y2=4.7
r195 (  67 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.815 //y=1.21 //x2=38.775 //y2=1.365
r196 (  66 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.815 //y=0.865 //x2=38.775 //y2=0.71
r197 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=38.815 //y=0.865 //x2=38.815 //y2=1.21
r198 (  64 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=38.44 //y=1.365 //x2=38.325 //y2=1.365
r199 (  63 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=38.66 //y=1.365 //x2=38.775 //y2=1.365
r200 (  62 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=38.44 //y=0.71 //x2=38.325 //y2=0.71
r201 (  61 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=38.66 //y=0.71 //x2=38.775 //y2=0.71
r202 (  61 62 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=38.66 //y=0.71 //x2=38.44 //y2=0.71
r203 (  58 75 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=38.38 //y=4.865 //x2=38.38 //y2=4.7
r204 (  57 72 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=38.285 //y=1.915 //x2=38.48 //y2=2.08
r205 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.285 //y=1.52 //x2=38.325 //y2=1.365
r206 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=38.285 //y=1.52 //x2=38.285 //y2=1.915
r207 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.285 //y=1.21 //x2=38.325 //y2=1.365
r208 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=38.285 //y=0.865 //x2=38.325 //y2=0.71
r209 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=38.285 //y=0.865 //x2=38.285 //y2=1.21
r210 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=38.82 //y=6.02 //x2=38.82 //y2=4.865
r211 (  52 58 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=38.38 //y=6.02 //x2=38.38 //y2=4.865
r212 (  51 63 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=38.55 //y=1.365 //x2=38.66 //y2=1.365
r213 (  51 64 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=38.55 //y=1.365 //x2=38.44 //y2=1.365
r214 (  47 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=38.48 //y=4.7 //x2=38.48 //y2=4.7
r215 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=38.48 //y=2.59 //x2=38.48 //y2=4.7
r216 (  42 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=38.48 //y=2.08 //x2=38.48 //y2=2.08
r217 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=38.48 //y=2.08 //x2=38.48 //y2=2.59
r218 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=36.63 //y=5.07 //x2=36.63 //y2=2.59
r219 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=36.63 //y=1.75 //x2=36.63 //y2=2.59
r220 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=36.545 //y=1.665 //x2=36.63 //y2=1.75
r221 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=36.545 //y=1.665 //x2=36.23 //y2=1.665
r222 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=36.145 //y=1.58 //x2=36.23 //y2=1.665
r223 (  31 80 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=36.145 //y=1.58 //x2=36.145 //y2=1.01
r224 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.935 //y=5.155 //x2=35.85 //y2=5.155
r225 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=36.545 //y=5.155 //x2=36.63 //y2=5.07
r226 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=36.545 //y=5.155 //x2=35.935 //y2=5.155
r227 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.85 //y=5.24 //x2=35.85 //y2=5.155
r228 (  23 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=35.85 //y=5.24 //x2=35.85 //y2=5.725
r229 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.055 //y=5.155 //x2=34.97 //y2=5.155
r230 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.765 //y=5.155 //x2=35.85 //y2=5.155
r231 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=35.765 //y=5.155 //x2=35.055 //y2=5.155
r232 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.97 //y=5.24 //x2=34.97 //y2=5.155
r233 (  15 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=34.97 //y=5.24 //x2=34.97 //y2=5.725
r234 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.885 //y=5.155 //x2=34.97 //y2=5.155
r235 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=34.885 //y=5.155 //x2=34.175 //y2=5.155
r236 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=34.09 //y=5.24 //x2=34.175 //y2=5.155
r237 (  7 82 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=34.09 //y=5.24 //x2=34.09 //y2=5.725
r238 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=38.48 //y=2.59 //x2=38.48 //y2=2.59
r239 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=36.63 //y=2.59 //x2=36.63 //y2=2.59
r240 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=36.745 //y=2.59 //x2=36.63 //y2=2.59
r241 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=38.365 //y=2.59 //x2=38.48 //y2=2.59
r242 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=38.365 //y=2.59 //x2=36.745 //y2=2.59
ends PM_TMRDFFSNQX1\%noxref_9

subckt PM_TMRDFFSNQX1\%noxref_10 ( 1 2 3 4 11 13 23 24 31 39 45 46 50 52 61 62 \
 64 65 67 68 69 70 71 72 73 74 75 80 82 84 90 91 92 93 94 95 99 101 104 105 \
 110 111 114 128 131 133 134 135 )
c281 ( 135 0 ) capacitor c=0.023087f //x=30.895 //y=5.02
c282 ( 134 0 ) capacitor c=0.023519f //x=30.015 //y=5.02
c283 ( 133 0 ) capacitor c=0.0224735f //x=29.135 //y=5.02
c284 ( 131 0 ) capacitor c=0.00853354f //x=31.145 //y=0.915
c285 ( 128 0 ) capacitor c=0.0588816f //x=41.81 //y=4.7
c286 ( 114 0 ) capacitor c=0.0331095f //x=26.3 //y=4.7
c287 ( 111 0 ) capacitor c=0.0279499f //x=26.27 //y=1.915
c288 ( 110 0 ) capacitor c=0.0421676f //x=26.27 //y=2.08
c289 ( 105 0 ) capacitor c=0.0318948f //x=42.145 //y=1.21
c290 ( 104 0 ) capacitor c=0.0187384f //x=42.145 //y=0.865
c291 ( 101 0 ) capacitor c=0.0141798f //x=41.99 //y=1.365
c292 ( 99 0 ) capacitor c=0.0149844f //x=41.99 //y=0.71
c293 ( 95 0 ) capacitor c=0.0813322f //x=41.615 //y=1.915
c294 ( 94 0 ) capacitor c=0.0229267f //x=41.615 //y=1.52
c295 ( 93 0 ) capacitor c=0.0234352f //x=41.615 //y=1.21
c296 ( 92 0 ) capacitor c=0.0199343f //x=41.615 //y=0.865
c297 ( 91 0 ) capacitor c=0.0429696f //x=26.835 //y=1.25
c298 ( 90 0 ) capacitor c=0.0192208f //x=26.835 //y=0.905
c299 ( 84 0 ) capacitor c=0.0148884f //x=26.68 //y=1.405
c300 ( 82 0 ) capacitor c=0.0157803f //x=26.68 //y=0.75
c301 ( 80 0 ) capacitor c=0.0295235f //x=26.675 //y=4.79
c302 ( 75 0 ) capacitor c=0.0205163f //x=26.305 //y=1.56
c303 ( 74 0 ) capacitor c=0.0168481f //x=26.305 //y=1.25
c304 ( 73 0 ) capacitor c=0.0174783f //x=26.305 //y=0.905
c305 ( 72 0 ) capacitor c=0.110275f //x=42.15 //y=6.02
c306 ( 71 0 ) capacitor c=0.154305f //x=41.71 //y=6.02
c307 ( 70 0 ) capacitor c=0.15358f //x=26.75 //y=6.02
c308 ( 69 0 ) capacitor c=0.110281f //x=26.31 //y=6.02
c309 ( 65 0 ) capacitor c=0.0715637f //x=31.817 //y=3.905
c310 ( 64 0 ) capacitor c=0.0101843f //x=31.815 //y=4.07
c311 ( 62 0 ) capacitor c=0.00106608f //x=31.04 //y=5.155
c312 ( 61 0 ) capacitor c=0.00207162f //x=30.16 //y=5.155
c313 ( 52 0 ) capacitor c=0.0857541f //x=41.81 //y=2.08
c314 ( 50 0 ) capacitor c=0.0236247f //x=31.82 //y=5.07
c315 ( 46 0 ) capacitor c=0.00398962f //x=31.42 //y=1.665
c316 ( 45 0 ) capacitor c=0.0135805f //x=31.735 //y=1.665
c317 ( 39 0 ) capacitor c=0.0281378f //x=31.735 //y=5.155
c318 ( 31 0 ) capacitor c=0.0176454f //x=30.955 //y=5.155
c319 ( 24 0 ) capacitor c=0.00332903f //x=29.365 //y=5.155
c320 ( 23 0 ) capacitor c=0.014837f //x=30.075 //y=5.155
c321 ( 13 0 ) capacitor c=0.0705158f //x=26.27 //y=2.08
c322 ( 11 0 ) capacitor c=0.00453889f //x=26.27 //y=4.535
c323 ( 4 0 ) capacitor c=0.00551102f //x=31.93 //y=4.07
c324 ( 3 0 ) capacitor c=0.141703f //x=41.695 //y=4.07
c325 ( 2 0 ) capacitor c=0.0142462f //x=26.385 //y=4.07
c326 ( 1 0 ) capacitor c=0.0882171f //x=31.7 //y=4.07
r327 (  126 128 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=41.71 //y=4.7 //x2=41.81 //y2=4.7
r328 (  116 117 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=26.3 //y=4.79 //x2=26.3 //y2=4.865
r329 (  114 116 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=26.3 //y=4.7 //x2=26.3 //y2=4.79
r330 (  110 111 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=26.27 //y=2.08 //x2=26.27 //y2=1.915
r331 (  106 128 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=42.15 //y=4.865 //x2=41.81 //y2=4.7
r332 (  105 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.145 //y=1.21 //x2=42.105 //y2=1.365
r333 (  104 129 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.145 //y=0.865 //x2=42.105 //y2=0.71
r334 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=42.145 //y=0.865 //x2=42.145 //y2=1.21
r335 (  102 125 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.77 //y=1.365 //x2=41.655 //y2=1.365
r336 (  101 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.99 //y=1.365 //x2=42.105 //y2=1.365
r337 (  100 124 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.77 //y=0.71 //x2=41.655 //y2=0.71
r338 (  99 129 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=41.99 //y=0.71 //x2=42.105 //y2=0.71
r339 (  99 100 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=41.99 //y=0.71 //x2=41.77 //y2=0.71
r340 (  96 126 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=41.71 //y=4.865 //x2=41.71 //y2=4.7
r341 (  95 123 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=41.615 //y=1.915 //x2=41.81 //y2=2.08
r342 (  94 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.615 //y=1.52 //x2=41.655 //y2=1.365
r343 (  94 95 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=41.615 //y=1.52 //x2=41.615 //y2=1.915
r344 (  93 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.615 //y=1.21 //x2=41.655 //y2=1.365
r345 (  92 124 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=41.615 //y=0.865 //x2=41.655 //y2=0.71
r346 (  92 93 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=41.615 //y=0.865 //x2=41.615 //y2=1.21
r347 (  91 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.835 //y=1.25 //x2=26.795 //y2=1.405
r348 (  90 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.835 //y=0.905 //x2=26.795 //y2=0.75
r349 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=26.835 //y=0.905 //x2=26.835 //y2=1.25
r350 (  85 119 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.46 //y=1.405 //x2=26.345 //y2=1.405
r351 (  84 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.68 //y=1.405 //x2=26.795 //y2=1.405
r352 (  83 118 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.46 //y=0.75 //x2=26.345 //y2=0.75
r353 (  82 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=26.68 //y=0.75 //x2=26.795 //y2=0.75
r354 (  82 83 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=26.68 //y=0.75 //x2=26.46 //y2=0.75
r355 (  81 116 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=26.435 //y=4.79 //x2=26.3 //y2=4.79
r356 (  80 87 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=26.675 //y=4.79 //x2=26.75 //y2=4.865
r357 (  80 81 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=26.675 //y=4.79 //x2=26.435 //y2=4.79
r358 (  75 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.305 //y=1.56 //x2=26.345 //y2=1.405
r359 (  75 111 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=26.305 //y=1.56 //x2=26.305 //y2=1.915
r360 (  74 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.305 //y=1.25 //x2=26.345 //y2=1.405
r361 (  73 118 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=26.305 //y=0.905 //x2=26.345 //y2=0.75
r362 (  73 74 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=26.305 //y=0.905 //x2=26.305 //y2=1.25
r363 (  72 106 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=42.15 //y=6.02 //x2=42.15 //y2=4.865
r364 (  71 96 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=41.71 //y=6.02 //x2=41.71 //y2=4.865
r365 (  70 87 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.75 //y=6.02 //x2=26.75 //y2=4.865
r366 (  69 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=26.31 //y=6.02 //x2=26.31 //y2=4.865
r367 (  68 101 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=41.88 //y=1.365 //x2=41.99 //y2=1.365
r368 (  68 102 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=41.88 //y=1.365 //x2=41.77 //y2=1.365
r369 (  67 84 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=26.57 //y=1.405 //x2=26.68 //y2=1.405
r370 (  67 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=26.57 //y=1.405 //x2=26.46 //y2=1.405
r371 (  64 66 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=31.817 //y=4.07 //x2=31.817 //y2=4.235
r372 (  64 65 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=31.817 //y=4.07 //x2=31.817 //y2=3.905
r373 (  60 114 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.3 //y=4.7 //x2=26.3 //y2=4.7
r374 (  57 128 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=41.81 //y=4.7 //x2=41.81 //y2=4.7
r375 (  55 57 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=41.81 //y=4.07 //x2=41.81 //y2=4.7
r376 (  52 123 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=41.81 //y=2.08 //x2=41.81 //y2=2.08
r377 (  52 55 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=41.81 //y=2.08 //x2=41.81 //y2=4.07
r378 (  50 66 ) resistor r=57.1551 //w=0.187 //l=0.835 //layer=li \
 //thickness=0.1 //x=31.82 //y=5.07 //x2=31.82 //y2=4.235
r379 (  47 65 ) resistor r=147.508 //w=0.187 //l=2.155 //layer=li \
 //thickness=0.1 //x=31.82 //y=1.75 //x2=31.82 //y2=3.905
r380 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=31.735 //y=1.665 //x2=31.82 //y2=1.75
r381 (  45 46 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=31.735 //y=1.665 //x2=31.42 //y2=1.665
r382 (  41 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=31.335 //y=1.58 //x2=31.42 //y2=1.665
r383 (  41 131 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=31.335 //y=1.58 //x2=31.335 //y2=1.01
r384 (  40 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.125 //y=5.155 //x2=31.04 //y2=5.155
r385 (  39 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=31.735 //y=5.155 //x2=31.82 //y2=5.07
r386 (  39 40 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=31.735 //y=5.155 //x2=31.125 //y2=5.155
r387 (  33 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=31.04 //y=5.24 //x2=31.04 //y2=5.155
r388 (  33 135 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=31.04 //y=5.24 //x2=31.04 //y2=5.725
r389 (  32 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.245 //y=5.155 //x2=30.16 //y2=5.155
r390 (  31 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.955 //y=5.155 //x2=31.04 //y2=5.155
r391 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=30.955 //y=5.155 //x2=30.245 //y2=5.155
r392 (  25 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.16 //y=5.24 //x2=30.16 //y2=5.155
r393 (  25 134 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=30.16 //y=5.24 //x2=30.16 //y2=5.725
r394 (  23 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.075 //y=5.155 //x2=30.16 //y2=5.155
r395 (  23 24 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=30.075 //y=5.155 //x2=29.365 //y2=5.155
r396 (  17 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=29.28 //y=5.24 //x2=29.365 //y2=5.155
r397 (  17 133 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=29.28 //y=5.24 //x2=29.28 //y2=5.725
r398 (  13 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=26.27 //y=2.08 //x2=26.27 //y2=2.08
r399 (  13 16 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=26.27 //y=2.08 //x2=26.27 //y2=4.07
r400 (  11 60 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=26.27 //y=4.535 //x2=26.285 //y2=4.7
r401 (  11 16 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=26.27 //y=4.535 //x2=26.27 //y2=4.07
r402 (  10 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=41.81 //y=4.07 //x2=41.81 //y2=4.07
r403 (  8 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=31.815 //y=4.07 //x2=31.815 //y2=4.07
r404 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=26.27 //y=4.07 //x2=26.27 //y2=4.07
r405 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.93 //y=4.07 //x2=31.815 //y2=4.07
r406 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=41.695 //y=4.07 //x2=41.81 //y2=4.07
r407 (  3 4 ) resistor r=9.31775 //w=0.131 //l=9.765 //layer=m1 \
 //thickness=0.36 //x=41.695 //y=4.07 //x2=31.93 //y2=4.07
r408 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=26.385 //y=4.07 //x2=26.27 //y2=4.07
r409 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.7 //y=4.07 //x2=31.815 //y2=4.07
r410 (  1 2 ) resistor r=5.07156 //w=0.131 //l=5.315 //layer=m1 \
 //thickness=0.36 //x=31.7 //y=4.07 //x2=26.385 //y2=4.07
ends PM_TMRDFFSNQX1\%noxref_10

subckt PM_TMRDFFSNQX1\%noxref_11 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 \
 47 48 49 51 57 58 59 60 72 74 75 )
c155 ( 75 0 ) capacitor c=0.0220291f //x=42.665 //y=5.02
c156 ( 74 0 ) capacitor c=0.0217503f //x=41.785 //y=5.02
c157 ( 72 0 ) capacitor c=0.0084702f //x=42.66 //y=0.905
c158 ( 60 0 ) capacitor c=0.0556143f //x=45.415 //y=4.79
c159 ( 59 0 ) capacitor c=0.0293157f //x=45.705 //y=4.79
c160 ( 58 0 ) capacitor c=0.0347816f //x=45.37 //y=1.22
c161 ( 57 0 ) capacitor c=0.0187487f //x=45.37 //y=0.875
c162 ( 51 0 ) capacitor c=0.0137055f //x=45.215 //y=1.375
c163 ( 49 0 ) capacitor c=0.0149861f //x=45.215 //y=0.72
c164 ( 48 0 ) capacitor c=0.096037f //x=44.84 //y=1.915
c165 ( 47 0 ) capacitor c=0.0228993f //x=44.84 //y=1.53
c166 ( 46 0 ) capacitor c=0.0234352f //x=44.84 //y=1.22
c167 ( 45 0 ) capacitor c=0.0198724f //x=44.84 //y=0.875
c168 ( 44 0 ) capacitor c=0.110114f //x=45.78 //y=6.02
c169 ( 43 0 ) capacitor c=0.158956f //x=45.34 //y=6.02
c170 ( 41 0 ) capacitor c=0.00211606f //x=42.81 //y=5.2
c171 ( 34 0 ) capacitor c=0.0944841f //x=45.14 //y=2.08
c172 ( 32 0 ) capacitor c=0.10219f //x=43.29 //y=2.59
c173 ( 28 0 ) capacitor c=0.00404073f //x=42.935 //y=1.655
c174 ( 27 0 ) capacitor c=0.0122201f //x=43.205 //y=1.655
c175 ( 25 0 ) capacitor c=0.0137995f //x=43.205 //y=5.2
c176 ( 14 0 ) capacitor c=0.00251459f //x=42.015 //y=5.2
c177 ( 13 0 ) capacitor c=0.0143649f //x=42.725 //y=5.2
c178 ( 2 0 ) capacitor c=0.0115544f //x=43.405 //y=2.59
c179 ( 1 0 ) capacitor c=0.0317176f //x=45.025 //y=2.59
r180 (  59 61 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=45.705 //y=4.79 //x2=45.78 //y2=4.865
r181 (  59 60 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=45.705 //y=4.79 //x2=45.415 //y2=4.79
r182 (  58 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.37 //y=1.22 //x2=45.33 //y2=1.375
r183 (  57 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.37 //y=0.875 //x2=45.33 //y2=0.72
r184 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=45.37 //y=0.875 //x2=45.37 //y2=1.22
r185 (  54 60 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=45.34 //y=4.865 //x2=45.415 //y2=4.79
r186 (  54 69 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=45.34 //y=4.865 //x2=45.14 //y2=4.7
r187 (  52 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.995 //y=1.375 //x2=44.88 //y2=1.375
r188 (  51 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.215 //y=1.375 //x2=45.33 //y2=1.375
r189 (  50 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=44.995 //y=0.72 //x2=44.88 //y2=0.72
r190 (  49 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.215 //y=0.72 //x2=45.33 //y2=0.72
r191 (  49 50 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=45.215 //y=0.72 //x2=44.995 //y2=0.72
r192 (  48 67 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=44.84 //y=1.915 //x2=45.14 //y2=2.08
r193 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.84 //y=1.53 //x2=44.88 //y2=1.375
r194 (  47 48 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=44.84 //y=1.53 //x2=44.84 //y2=1.915
r195 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.84 //y=1.22 //x2=44.88 //y2=1.375
r196 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=44.84 //y=0.875 //x2=44.88 //y2=0.72
r197 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=44.84 //y=0.875 //x2=44.84 //y2=1.22
r198 (  44 61 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.78 //y=6.02 //x2=45.78 //y2=4.865
r199 (  43 54 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=45.34 //y=6.02 //x2=45.34 //y2=4.865
r200 (  42 51 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=45.105 //y=1.375 //x2=45.215 //y2=1.375
r201 (  42 52 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=45.105 //y=1.375 //x2=44.995 //y2=1.375
r202 (  39 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=45.14 //y=4.7 //x2=45.14 //y2=4.7
r203 (  37 39 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=45.14 //y=2.59 //x2=45.14 //y2=4.7
r204 (  34 67 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=45.14 //y=2.08 //x2=45.14 //y2=2.08
r205 (  34 37 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=45.14 //y=2.08 //x2=45.14 //y2=2.59
r206 (  30 32 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=43.29 //y=5.115 //x2=43.29 //y2=2.59
r207 (  29 32 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=43.29 //y=1.74 //x2=43.29 //y2=2.59
r208 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=43.205 //y=1.655 //x2=43.29 //y2=1.74
r209 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=43.205 //y=1.655 //x2=42.935 //y2=1.655
r210 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.895 //y=5.2 //x2=42.81 //y2=5.2
r211 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=43.205 //y=5.2 //x2=43.29 //y2=5.115
r212 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=43.205 //y=5.2 //x2=42.895 //y2=5.2
r213 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=42.85 //y=1.57 //x2=42.935 //y2=1.655
r214 (  21 72 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=42.85 //y=1.57 //x2=42.85 //y2=1
r215 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.81 //y=5.285 //x2=42.81 //y2=5.2
r216 (  15 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=42.81 //y=5.285 //x2=42.81 //y2=5.725
r217 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=42.725 //y=5.2 //x2=42.81 //y2=5.2
r218 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=42.725 //y=5.2 //x2=42.015 //y2=5.2
r219 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=41.93 //y=5.285 //x2=42.015 //y2=5.2
r220 (  7 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=41.93 //y=5.285 //x2=41.93 //y2=5.725
r221 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=45.14 //y=2.59 //x2=45.14 //y2=2.59
r222 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=43.29 //y=2.59 //x2=43.29 //y2=2.59
r223 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=43.405 //y=2.59 //x2=43.29 //y2=2.59
r224 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=45.025 //y=2.59 //x2=45.14 //y2=2.59
r225 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=45.025 //y=2.59 //x2=43.405 //y2=2.59
ends PM_TMRDFFSNQX1\%noxref_11

subckt PM_TMRDFFSNQX1\%noxref_12 ( 1 2 3 4 5 6 16 24 37 38 49 51 52 56 58 65 \
 66 67 68 69 70 71 72 73 74 78 79 80 85 87 90 91 95 96 97 102 104 107 108 112 \
 113 114 119 121 124 125 127 128 133 137 138 143 147 148 153 156 158 159 )
c322 ( 159 0 ) capacitor c=0.0220291f //x=39.335 //y=5.02
c323 ( 158 0 ) capacitor c=0.0217503f //x=38.455 //y=5.02
c324 ( 156 0 ) capacitor c=0.00866655f //x=39.33 //y=0.905
c325 ( 153 0 ) capacitor c=0.0587755f //x=47.36 //y=4.7
c326 ( 148 0 ) capacitor c=0.0273931f //x=47.36 //y=1.915
c327 ( 147 0 ) capacitor c=0.0456313f //x=47.36 //y=2.08
c328 ( 143 0 ) capacitor c=0.0587755f //x=35.89 //y=4.7
c329 ( 138 0 ) capacitor c=0.0273931f //x=35.89 //y=1.915
c330 ( 137 0 ) capacitor c=0.0456313f //x=35.89 //y=2.08
c331 ( 133 0 ) capacitor c=0.058931f //x=31.08 //y=4.7
c332 ( 128 0 ) capacitor c=0.0267105f //x=31.08 //y=1.915
c333 ( 127 0 ) capacitor c=0.0456313f //x=31.08 //y=2.08
c334 ( 125 0 ) capacitor c=0.0432517f //x=47.88 //y=1.26
c335 ( 124 0 ) capacitor c=0.0200379f //x=47.88 //y=0.915
c336 ( 121 0 ) capacitor c=0.0148873f //x=47.725 //y=1.415
c337 ( 119 0 ) capacitor c=0.0157803f //x=47.725 //y=0.76
c338 ( 114 0 ) capacitor c=0.0218028f //x=47.35 //y=1.57
c339 ( 113 0 ) capacitor c=0.0207459f //x=47.35 //y=1.26
c340 ( 112 0 ) capacitor c=0.0194308f //x=47.35 //y=0.915
c341 ( 108 0 ) capacitor c=0.0432517f //x=36.41 //y=1.26
c342 ( 107 0 ) capacitor c=0.0200379f //x=36.41 //y=0.915
c343 ( 104 0 ) capacitor c=0.0148873f //x=36.255 //y=1.415
c344 ( 102 0 ) capacitor c=0.0157803f //x=36.255 //y=0.76
c345 ( 97 0 ) capacitor c=0.0218028f //x=35.88 //y=1.57
c346 ( 96 0 ) capacitor c=0.0207459f //x=35.88 //y=1.26
c347 ( 95 0 ) capacitor c=0.0194308f //x=35.88 //y=0.915
c348 ( 91 0 ) capacitor c=0.0432517f //x=31.6 //y=1.26
c349 ( 90 0 ) capacitor c=0.0200379f //x=31.6 //y=0.915
c350 ( 87 0 ) capacitor c=0.0148873f //x=31.445 //y=1.415
c351 ( 85 0 ) capacitor c=0.0157803f //x=31.445 //y=0.76
c352 ( 80 0 ) capacitor c=0.0218028f //x=31.07 //y=1.57
c353 ( 79 0 ) capacitor c=0.0207459f //x=31.07 //y=1.26
c354 ( 78 0 ) capacitor c=0.0194308f //x=31.07 //y=0.915
c355 ( 74 0 ) capacitor c=0.158794f //x=47.54 //y=6.02
c356 ( 73 0 ) capacitor c=0.110114f //x=47.1 //y=6.02
c357 ( 72 0 ) capacitor c=0.158794f //x=36.07 //y=6.02
c358 ( 71 0 ) capacitor c=0.110114f //x=35.63 //y=6.02
c359 ( 70 0 ) capacitor c=0.158048f //x=31.26 //y=6.02
c360 ( 69 0 ) capacitor c=0.110114f //x=30.82 //y=6.02
c361 ( 65 0 ) capacitor c=0.00211606f //x=39.48 //y=5.2
c362 ( 58 0 ) capacitor c=0.0808586f //x=47.36 //y=2.08
c363 ( 56 0 ) capacitor c=0.103614f //x=39.96 //y=3.7
c364 ( 52 0 ) capacitor c=0.00404073f //x=39.605 //y=1.655
c365 ( 51 0 ) capacitor c=0.0122201f //x=39.875 //y=1.655
c366 ( 49 0 ) capacitor c=0.0137522f //x=39.875 //y=5.2
c367 ( 38 0 ) capacitor c=0.00251635f //x=38.685 //y=5.2
c368 ( 37 0 ) capacitor c=0.0142529f //x=39.395 //y=5.2
c369 ( 24 0 ) capacitor c=0.0811636f //x=35.89 //y=2.08
c370 ( 16 0 ) capacitor c=0.0796434f //x=31.08 //y=2.08
c371 ( 6 0 ) capacitor c=0.00405261f //x=40.075 //y=3.7
c372 ( 5 0 ) capacitor c=0.120326f //x=47.245 //y=3.7
c373 ( 4 0 ) capacitor c=0.00412452f //x=36.005 //y=3.7
c374 ( 3 0 ) capacitor c=0.0546427f //x=39.845 //y=3.7
c375 ( 2 0 ) capacitor c=0.0138772f //x=31.195 //y=3.7
c376 ( 1 0 ) capacitor c=0.0670382f //x=35.775 //y=3.7
r377 (  147 148 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=47.36 //y=2.08 //x2=47.36 //y2=1.915
r378 (  137 138 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=35.89 //y=2.08 //x2=35.89 //y2=1.915
r379 (  127 128 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=31.08 //y=2.08 //x2=31.08 //y2=1.915
r380 (  125 155 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.88 //y=1.26 //x2=47.84 //y2=1.415
r381 (  124 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.88 //y=0.915 //x2=47.84 //y2=0.76
r382 (  124 125 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=47.88 //y=0.915 //x2=47.88 //y2=1.26
r383 (  122 151 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=47.505 //y=1.415 //x2=47.39 //y2=1.415
r384 (  121 155 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=47.725 //y=1.415 //x2=47.84 //y2=1.415
r385 (  120 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=47.505 //y=0.76 //x2=47.39 //y2=0.76
r386 (  119 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=47.725 //y=0.76 //x2=47.84 //y2=0.76
r387 (  119 120 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=47.725 //y=0.76 //x2=47.505 //y2=0.76
r388 (  116 153 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=47.54 //y=4.865 //x2=47.36 //y2=4.7
r389 (  114 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.35 //y=1.57 //x2=47.39 //y2=1.415
r390 (  114 148 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=47.35 //y=1.57 //x2=47.35 //y2=1.915
r391 (  113 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.35 //y=1.26 //x2=47.39 //y2=1.415
r392 (  112 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=47.35 //y=0.915 //x2=47.39 //y2=0.76
r393 (  112 113 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=47.35 //y=0.915 //x2=47.35 //y2=1.26
r394 (  109 153 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=47.1 //y=4.865 //x2=47.36 //y2=4.7
r395 (  108 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.41 //y=1.26 //x2=36.37 //y2=1.415
r396 (  107 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=36.41 //y=0.915 //x2=36.37 //y2=0.76
r397 (  107 108 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=36.41 //y=0.915 //x2=36.41 //y2=1.26
r398 (  105 141 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=36.035 //y=1.415 //x2=35.92 //y2=1.415
r399 (  104 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=36.255 //y=1.415 //x2=36.37 //y2=1.415
r400 (  103 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=36.035 //y=0.76 //x2=35.92 //y2=0.76
r401 (  102 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=36.255 //y=0.76 //x2=36.37 //y2=0.76
r402 (  102 103 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=36.255 //y=0.76 //x2=36.035 //y2=0.76
r403 (  99 143 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=36.07 //y=4.865 //x2=35.89 //y2=4.7
r404 (  97 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.88 //y=1.57 //x2=35.92 //y2=1.415
r405 (  97 138 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=35.88 //y=1.57 //x2=35.88 //y2=1.915
r406 (  96 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.88 //y=1.26 //x2=35.92 //y2=1.415
r407 (  95 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=35.88 //y=0.915 //x2=35.92 //y2=0.76
r408 (  95 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=35.88 //y=0.915 //x2=35.88 //y2=1.26
r409 (  92 143 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=35.63 //y=4.865 //x2=35.89 //y2=4.7
r410 (  91 135 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.6 //y=1.26 //x2=31.56 //y2=1.415
r411 (  90 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.6 //y=0.915 //x2=31.56 //y2=0.76
r412 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=31.6 //y=0.915 //x2=31.6 //y2=1.26
r413 (  88 131 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.225 //y=1.415 //x2=31.11 //y2=1.415
r414 (  87 135 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.445 //y=1.415 //x2=31.56 //y2=1.415
r415 (  86 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.225 //y=0.76 //x2=31.11 //y2=0.76
r416 (  85 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=31.445 //y=0.76 //x2=31.56 //y2=0.76
r417 (  85 86 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=31.445 //y=0.76 //x2=31.225 //y2=0.76
r418 (  82 133 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=31.26 //y=4.865 //x2=31.08 //y2=4.7
r419 (  80 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.07 //y=1.57 //x2=31.11 //y2=1.415
r420 (  80 128 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=31.07 //y=1.57 //x2=31.07 //y2=1.915
r421 (  79 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.07 //y=1.26 //x2=31.11 //y2=1.415
r422 (  78 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=31.07 //y=0.915 //x2=31.11 //y2=0.76
r423 (  78 79 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=31.07 //y=0.915 //x2=31.07 //y2=1.26
r424 (  75 133 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=30.82 //y=4.865 //x2=31.08 //y2=4.7
r425 (  74 116 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=47.54 //y=6.02 //x2=47.54 //y2=4.865
r426 (  73 109 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=47.1 //y=6.02 //x2=47.1 //y2=4.865
r427 (  72 99 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=36.07 //y=6.02 //x2=36.07 //y2=4.865
r428 (  71 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=35.63 //y=6.02 //x2=35.63 //y2=4.865
r429 (  70 82 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=31.26 //y=6.02 //x2=31.26 //y2=4.865
r430 (  69 75 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=30.82 //y=6.02 //x2=30.82 //y2=4.865
r431 (  68 121 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=47.615 //y=1.415 //x2=47.725 //y2=1.415
r432 (  68 122 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=47.615 //y=1.415 //x2=47.505 //y2=1.415
r433 (  67 104 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=36.145 //y=1.415 //x2=36.255 //y2=1.415
r434 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=36.145 //y=1.415 //x2=36.035 //y2=1.415
r435 (  66 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=31.335 //y=1.415 //x2=31.445 //y2=1.415
r436 (  66 88 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=31.335 //y=1.415 //x2=31.225 //y2=1.415
r437 (  63 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=47.36 //y=4.7 //x2=47.36 //y2=4.7
r438 (  61 63 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=47.36 //y=3.7 //x2=47.36 //y2=4.7
r439 (  58 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=47.36 //y=2.08 //x2=47.36 //y2=2.08
r440 (  58 61 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=47.36 //y=2.08 //x2=47.36 //y2=3.7
r441 (  54 56 ) resistor r=96.8556 //w=0.187 //l=1.415 //layer=li \
 //thickness=0.1 //x=39.96 //y=5.115 //x2=39.96 //y2=3.7
r442 (  53 56 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=39.96 //y=1.74 //x2=39.96 //y2=3.7
r443 (  51 53 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=39.875 //y=1.655 //x2=39.96 //y2=1.74
r444 (  51 52 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=39.875 //y=1.655 //x2=39.605 //y2=1.655
r445 (  50 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.565 //y=5.2 //x2=39.48 //y2=5.2
r446 (  49 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=39.875 //y=5.2 //x2=39.96 //y2=5.115
r447 (  49 50 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=39.875 //y=5.2 //x2=39.565 //y2=5.2
r448 (  45 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=39.52 //y=1.57 //x2=39.605 //y2=1.655
r449 (  45 156 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=39.52 //y=1.57 //x2=39.52 //y2=1
r450 (  39 65 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.48 //y=5.285 //x2=39.48 //y2=5.2
r451 (  39 159 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=39.48 //y=5.285 //x2=39.48 //y2=5.725
r452 (  37 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=39.395 //y=5.2 //x2=39.48 //y2=5.2
r453 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=39.395 //y=5.2 //x2=38.685 //y2=5.2
r454 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=38.6 //y=5.285 //x2=38.685 //y2=5.2
r455 (  31 158 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=38.6 //y=5.285 //x2=38.6 //y2=5.725
r456 (  29 143 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=35.89 //y=4.7 //x2=35.89 //y2=4.7
r457 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=35.89 //y=3.7 //x2=35.89 //y2=4.7
r458 (  24 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=35.89 //y=2.08 //x2=35.89 //y2=2.08
r459 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=35.89 //y=2.08 //x2=35.89 //y2=3.7
r460 (  21 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.08 //y=4.7 //x2=31.08 //y2=4.7
r461 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=31.08 //y=3.7 //x2=31.08 //y2=4.7
r462 (  16 127 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=31.08 //y=2.08 //x2=31.08 //y2=2.08
r463 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=31.08 //y=2.08 //x2=31.08 //y2=3.7
r464 (  14 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=47.36 //y=3.7 //x2=47.36 //y2=3.7
r465 (  12 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=39.96 //y=3.7 //x2=39.96 //y2=3.7
r466 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=35.89 //y=3.7 //x2=35.89 //y2=3.7
r467 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=31.08 //y=3.7 //x2=31.08 //y2=3.7
r468 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=40.075 //y=3.7 //x2=39.96 //y2=3.7
r469 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=47.245 //y=3.7 //x2=47.36 //y2=3.7
r470 (  5 6 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=47.245 //y=3.7 //x2=40.075 //y2=3.7
r471 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=36.005 //y=3.7 //x2=35.89 //y2=3.7
r472 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=39.845 //y=3.7 //x2=39.96 //y2=3.7
r473 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=39.845 //y=3.7 //x2=36.005 //y2=3.7
r474 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=31.195 //y=3.7 //x2=31.08 //y2=3.7
r475 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=35.775 //y=3.7 //x2=35.89 //y2=3.7
r476 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=35.775 //y=3.7 //x2=31.195 //y2=3.7
ends PM_TMRDFFSNQX1\%noxref_12

subckt PM_TMRDFFSNQX1\%noxref_13 ( 1 2 3 4 6 7 8 9 10 23 25 35 36 43 51 57 58 \
 62 65 67 75 81 82 86 89 90 91 92 93 94 95 96 97 98 99 100 105 107 109 115 116 \
 117 118 119 124 126 128 134 135 136 137 138 143 145 147 153 154 156 157 160 \
 169 170 173 181 182 185 193 195 196 197 )
c467 ( 197 0 ) capacitor c=0.023087f //x=47.175 //y=5.02
c468 ( 196 0 ) capacitor c=0.023519f //x=46.295 //y=5.02
c469 ( 195 0 ) capacitor c=0.0224735f //x=45.415 //y=5.02
c470 ( 193 0 ) capacitor c=0.00872971f //x=47.425 //y=0.915
c471 ( 185 0 ) capacitor c=0.0352016f //x=81.79 //y=4.705
c472 ( 182 0 ) capacitor c=0.0279733f //x=81.77 //y=1.915
c473 ( 181 0 ) capacitor c=0.0467621f //x=81.77 //y=2.08
c474 ( 173 0 ) capacitor c=0.03845f //x=75.15 //y=4.705
c475 ( 170 0 ) capacitor c=0.0300885f //x=75.11 //y=1.915
c476 ( 169 0 ) capacitor c=0.0520257f //x=75.11 //y=2.08
c477 ( 160 0 ) capacitor c=0.0331095f //x=42.58 //y=4.7
c478 ( 157 0 ) capacitor c=0.0279499f //x=42.55 //y=1.915
c479 ( 156 0 ) capacitor c=0.0421676f //x=42.55 //y=2.08
c480 ( 154 0 ) capacitor c=0.0237734f //x=82.335 //y=1.255
c481 ( 153 0 ) capacitor c=0.0191782f //x=82.335 //y=0.905
c482 ( 147 0 ) capacitor c=0.0351663f //x=82.18 //y=1.405
c483 ( 145 0 ) capacitor c=0.0157803f //x=82.18 //y=0.75
c484 ( 143 0 ) capacitor c=0.0374703f //x=82.175 //y=4.795
c485 ( 138 0 ) capacitor c=0.0200628f //x=81.805 //y=1.56
c486 ( 137 0 ) capacitor c=0.0168575f //x=81.805 //y=1.255
c487 ( 136 0 ) capacitor c=0.0174993f //x=81.805 //y=0.905
c488 ( 135 0 ) capacitor c=0.0447087f //x=75.675 //y=1.25
c489 ( 134 0 ) capacitor c=0.019286f //x=75.675 //y=0.905
c490 ( 128 0 ) capacitor c=0.0187932f //x=75.52 //y=1.405
c491 ( 126 0 ) capacitor c=0.0157795f //x=75.52 //y=0.75
c492 ( 124 0 ) capacitor c=0.029531f //x=75.515 //y=4.795
c493 ( 119 0 ) capacitor c=0.0206178f //x=75.145 //y=1.56
c494 ( 118 0 ) capacitor c=0.016848f //x=75.145 //y=1.25
c495 ( 117 0 ) capacitor c=0.0174777f //x=75.145 //y=0.905
c496 ( 116 0 ) capacitor c=0.0429696f //x=43.115 //y=1.25
c497 ( 115 0 ) capacitor c=0.0192208f //x=43.115 //y=0.905
c498 ( 109 0 ) capacitor c=0.0148884f //x=42.96 //y=1.405
c499 ( 107 0 ) capacitor c=0.0157803f //x=42.96 //y=0.75
c500 ( 105 0 ) capacitor c=0.0295235f //x=42.955 //y=4.79
c501 ( 100 0 ) capacitor c=0.0205163f //x=42.585 //y=1.56
c502 ( 99 0 ) capacitor c=0.0168481f //x=42.585 //y=1.25
c503 ( 98 0 ) capacitor c=0.0174783f //x=42.585 //y=0.905
c504 ( 97 0 ) capacitor c=0.15325f //x=82.25 //y=6.025
c505 ( 96 0 ) capacitor c=0.110411f //x=81.81 //y=6.025
c506 ( 95 0 ) capacitor c=0.154236f //x=75.59 //y=6.025
c507 ( 94 0 ) capacitor c=0.110294f //x=75.15 //y=6.025
c508 ( 93 0 ) capacitor c=0.15358f //x=43.03 //y=6.02
c509 ( 92 0 ) capacitor c=0.110281f //x=42.59 //y=6.02
c510 ( 86 0 ) capacitor c=0.00501304f //x=81.79 //y=4.705
c511 ( 82 0 ) capacitor c=0.00106608f //x=47.32 //y=5.155
c512 ( 81 0 ) capacitor c=0.00207319f //x=46.44 //y=5.155
c513 ( 75 0 ) capacitor c=0.0901308f //x=81.77 //y=2.08
c514 ( 67 0 ) capacitor c=0.104623f //x=75.11 //y=2.08
c515 ( 65 0 ) capacitor c=0.00669947f //x=75.11 //y=4.54
c516 ( 62 0 ) capacitor c=0.106131f //x=48.1 //y=2.59
c517 ( 58 0 ) capacitor c=0.00398962f //x=47.7 //y=1.665
c518 ( 57 0 ) capacitor c=0.0137288f //x=48.015 //y=1.665
c519 ( 51 0 ) capacitor c=0.0284988f //x=48.015 //y=5.155
c520 ( 43 0 ) capacitor c=0.0176454f //x=47.235 //y=5.155
c521 ( 36 0 ) capacitor c=0.00332903f //x=45.645 //y=5.155
c522 ( 35 0 ) capacitor c=0.0148427f //x=46.355 //y=5.155
c523 ( 25 0 ) capacitor c=0.0689632f //x=42.55 //y=2.08
c524 ( 23 0 ) capacitor c=0.00453889f //x=42.55 //y=4.535
c525 ( 10 0 ) capacitor c=0.0144297f //x=75.225 //y=4.07
c526 ( 9 0 ) capacitor c=0.181505f //x=81.655 //y=4.07
c527 ( 8 0 ) capacitor c=1.21334e-19 //x=50.775 //y=2.96
c528 ( 7 0 ) capacitor c=0.431437f //x=74.995 //y=2.96
c529 ( 4 0 ) capacitor c=0.00871105f //x=48.215 //y=2.59
c530 ( 3 0 ) capacitor c=0.0344714f //x=50.605 //y=2.59
c531 ( 2 0 ) capacitor c=0.00621861f //x=42.665 //y=4.07
c532 ( 1 0 ) capacitor c=0.0841928f //x=47.985 //y=4.07
r533 (  187 188 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=81.79 //y=4.795 //x2=81.79 //y2=4.87
r534 (  185 187 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=81.79 //y=4.705 //x2=81.79 //y2=4.795
r535 (  181 182 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=81.77 //y=2.08 //x2=81.77 //y2=1.915
r536 (  173 175 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=75.15 //y=4.705 //x2=75.15 //y2=4.795
r537 (  169 170 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=75.11 //y=2.08 //x2=75.11 //y2=1.915
r538 (  162 163 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=42.58 //y=4.79 //x2=42.58 //y2=4.865
r539 (  160 162 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=42.58 //y=4.7 //x2=42.58 //y2=4.79
r540 (  156 157 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=42.55 //y=2.08 //x2=42.55 //y2=1.915
r541 (  154 192 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=82.335 //y=1.255 //x2=82.335 //y2=1.367
r542 (  153 191 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=82.335 //y=0.905 //x2=82.295 //y2=0.75
r543 (  153 154 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=82.335 //y=0.905 //x2=82.335 //y2=1.255
r544 (  148 190 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=81.96 //y=1.405 //x2=81.845 //y2=1.405
r545 (  147 192 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=82.18 //y=1.405 //x2=82.335 //y2=1.367
r546 (  146 189 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=81.96 //y=0.75 //x2=81.845 //y2=0.75
r547 (  145 191 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=82.18 //y=0.75 //x2=82.295 //y2=0.75
r548 (  145 146 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=82.18 //y=0.75 //x2=81.96 //y2=0.75
r549 (  144 187 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=81.925 //y=4.795 //x2=81.79 //y2=4.795
r550 (  143 150 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=82.175 //y=4.795 //x2=82.25 //y2=4.87
r551 (  143 144 ) resistor r=128.191 //w=0.094 //l=0.25 //layer=ply \
 //thickness=0.18 //x=82.175 //y=4.795 //x2=81.925 //y2=4.795
r552 (  138 190 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=81.805 //y=1.56 //x2=81.845 //y2=1.405
r553 (  138 182 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=81.805 //y=1.56 //x2=81.805 //y2=1.915
r554 (  137 190 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=81.805 //y=1.255 //x2=81.845 //y2=1.405
r555 (  136 189 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=81.805 //y=0.905 //x2=81.845 //y2=0.75
r556 (  136 137 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=81.805 //y=0.905 //x2=81.805 //y2=1.255
r557 (  135 179 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.675 //y=1.25 //x2=75.635 //y2=1.405
r558 (  134 178 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.675 //y=0.905 //x2=75.635 //y2=0.75
r559 (  134 135 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=75.675 //y=0.905 //x2=75.675 //y2=1.25
r560 (  129 177 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.3 //y=1.405 //x2=75.185 //y2=1.405
r561 (  128 179 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.52 //y=1.405 //x2=75.635 //y2=1.405
r562 (  127 176 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.3 //y=0.75 //x2=75.185 //y2=0.75
r563 (  126 178 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=75.52 //y=0.75 //x2=75.635 //y2=0.75
r564 (  126 127 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=75.52 //y=0.75 //x2=75.3 //y2=0.75
r565 (  125 175 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=75.285 //y=4.795 //x2=75.15 //y2=4.795
r566 (  124 131 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=75.515 //y=4.795 //x2=75.59 //y2=4.87
r567 (  124 125 ) resistor r=117.936 //w=0.094 //l=0.23 //layer=ply \
 //thickness=0.18 //x=75.515 //y=4.795 //x2=75.285 //y2=4.795
r568 (  121 175 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=75.15 //y=4.87 //x2=75.15 //y2=4.795
r569 (  119 177 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.145 //y=1.56 //x2=75.185 //y2=1.405
r570 (  119 170 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=75.145 //y=1.56 //x2=75.145 //y2=1.915
r571 (  118 177 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.145 //y=1.25 //x2=75.185 //y2=1.405
r572 (  117 176 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=75.145 //y=0.905 //x2=75.185 //y2=0.75
r573 (  117 118 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=75.145 //y=0.905 //x2=75.145 //y2=1.25
r574 (  116 167 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=43.115 //y=1.25 //x2=43.075 //y2=1.405
r575 (  115 166 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=43.115 //y=0.905 //x2=43.075 //y2=0.75
r576 (  115 116 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=43.115 //y=0.905 //x2=43.115 //y2=1.25
r577 (  110 165 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.74 //y=1.405 //x2=42.625 //y2=1.405
r578 (  109 167 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.96 //y=1.405 //x2=43.075 //y2=1.405
r579 (  108 164 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.74 //y=0.75 //x2=42.625 //y2=0.75
r580 (  107 166 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=42.96 //y=0.75 //x2=43.075 //y2=0.75
r581 (  107 108 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=42.96 //y=0.75 //x2=42.74 //y2=0.75
r582 (  106 162 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=42.715 //y=4.79 //x2=42.58 //y2=4.79
r583 (  105 112 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=42.955 //y=4.79 //x2=43.03 //y2=4.865
r584 (  105 106 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=42.955 //y=4.79 //x2=42.715 //y2=4.79
r585 (  100 165 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.585 //y=1.56 //x2=42.625 //y2=1.405
r586 (  100 157 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=42.585 //y=1.56 //x2=42.585 //y2=1.915
r587 (  99 165 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.585 //y=1.25 //x2=42.625 //y2=1.405
r588 (  98 164 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=42.585 //y=0.905 //x2=42.625 //y2=0.75
r589 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=42.585 //y=0.905 //x2=42.585 //y2=1.25
r590 (  97 150 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=82.25 //y=6.025 //x2=82.25 //y2=4.87
r591 (  96 188 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=81.81 //y=6.025 //x2=81.81 //y2=4.87
r592 (  95 131 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=75.59 //y=6.025 //x2=75.59 //y2=4.87
r593 (  94 121 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=75.15 //y=6.025 //x2=75.15 //y2=4.87
r594 (  93 112 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=43.03 //y=6.02 //x2=43.03 //y2=4.865
r595 (  92 163 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=42.59 //y=6.02 //x2=42.59 //y2=4.865
r596 (  91 147 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=82.07 //y=1.405 //x2=82.18 //y2=1.405
r597 (  91 148 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=82.07 //y=1.405 //x2=81.96 //y2=1.405
r598 (  90 128 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=75.41 //y=1.405 //x2=75.52 //y2=1.405
r599 (  90 129 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=75.41 //y=1.405 //x2=75.3 //y2=1.405
r600 (  89 109 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=42.85 //y=1.405 //x2=42.96 //y2=1.405
r601 (  89 110 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=42.85 //y=1.405 //x2=42.74 //y2=1.405
r602 (  86 185 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=81.79 //y=4.705 //x2=81.79 //y2=4.705
r603 (  86 87 ) resistor r=10.3507 //w=0.207 //l=0.165 //layer=li \
 //thickness=0.1 //x=81.78 //y=4.705 //x2=81.78 //y2=4.54
r604 (  84 173 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=75.15 //y=4.705 //x2=75.15 //y2=4.705
r605 (  80 160 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=42.58 //y=4.7 //x2=42.58 //y2=4.7
r606 (  78 87 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=81.77 //y=4.07 //x2=81.77 //y2=4.54
r607 (  75 181 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=81.77 //y=2.08 //x2=81.77 //y2=2.08
r608 (  75 78 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=81.77 //y=2.08 //x2=81.77 //y2=4.07
r609 (  70 72 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=75.11 //y=2.96 //x2=75.11 //y2=4.07
r610 (  67 169 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=75.11 //y=2.08 //x2=75.11 //y2=2.08
r611 (  67 70 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=75.11 //y=2.08 //x2=75.11 //y2=2.96
r612 (  65 84 ) resistor r=11.2426 //w=0.191 //l=0.174714 //layer=li \
 //thickness=0.1 //x=75.11 //y=4.54 //x2=75.13 //y2=4.705
r613 (  65 72 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=75.11 //y=4.54 //x2=75.11 //y2=4.07
r614 (  62 64 ) resistor r=101.305 //w=0.187 //l=1.48 //layer=li \
 //thickness=0.1 //x=48.1 //y=2.59 //x2=48.1 //y2=4.07
r615 (  60 64 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=48.1 //y=5.07 //x2=48.1 //y2=4.07
r616 (  59 62 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=48.1 //y=1.75 //x2=48.1 //y2=2.59
r617 (  57 59 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=48.015 //y=1.665 //x2=48.1 //y2=1.75
r618 (  57 58 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=48.015 //y=1.665 //x2=47.7 //y2=1.665
r619 (  53 58 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=47.615 //y=1.58 //x2=47.7 //y2=1.665
r620 (  53 193 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=47.615 //y=1.58 //x2=47.615 //y2=1.01
r621 (  52 82 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.405 //y=5.155 //x2=47.32 //y2=5.155
r622 (  51 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=48.015 //y=5.155 //x2=48.1 //y2=5.07
r623 (  51 52 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=48.015 //y=5.155 //x2=47.405 //y2=5.155
r624 (  45 82 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.32 //y=5.24 //x2=47.32 //y2=5.155
r625 (  45 197 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=47.32 //y=5.24 //x2=47.32 //y2=5.725
r626 (  44 81 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.525 //y=5.155 //x2=46.44 //y2=5.155
r627 (  43 82 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=47.235 //y=5.155 //x2=47.32 //y2=5.155
r628 (  43 44 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=47.235 //y=5.155 //x2=46.525 //y2=5.155
r629 (  37 81 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.44 //y=5.24 //x2=46.44 //y2=5.155
r630 (  37 196 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=46.44 //y=5.24 //x2=46.44 //y2=5.725
r631 (  35 81 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.355 //y=5.155 //x2=46.44 //y2=5.155
r632 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=46.355 //y=5.155 //x2=45.645 //y2=5.155
r633 (  29 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=45.56 //y=5.24 //x2=45.645 //y2=5.155
r634 (  29 195 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=45.56 //y=5.24 //x2=45.56 //y2=5.725
r635 (  25 156 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=42.55 //y=2.08 //x2=42.55 //y2=2.08
r636 (  25 28 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=42.55 //y=2.08 //x2=42.55 //y2=4.07
r637 (  23 80 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=42.55 //y=4.535 //x2=42.565 //y2=4.7
r638 (  23 28 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=42.55 //y=4.535 //x2=42.55 //y2=4.07
r639 (  22 78 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=81.77 //y=4.07 //x2=81.77 //y2=4.07
r640 (  20 70 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=75.11 //y=2.96 //x2=75.11 //y2=2.96
r641 (  18 72 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=75.11 //y=4.07 //x2=75.11 //y2=4.07
r642 (  16 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=48.1 //y=4.07 //x2=48.1 //y2=4.07
r643 (  14 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=48.1 //y=2.59 //x2=48.1 //y2=2.59
r644 (  12 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=42.55 //y=4.07 //x2=42.55 //y2=4.07
r645 (  10 18 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=75.225 //y=4.07 //x2=75.11 //y2=4.07
r646 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=81.655 //y=4.07 //x2=81.77 //y2=4.07
r647 (  9 10 ) resistor r=6.1355 //w=0.131 //l=6.43 //layer=m1 \
 //thickness=0.36 //x=81.655 //y=4.07 //x2=75.225 //y2=4.07
r648 (  7 20 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=74.995 //y=2.96 //x2=75.11 //y2=2.96
r649 (  7 8 ) resistor r=23.1107 //w=0.131 //l=24.22 //layer=m1 \
 //thickness=0.36 //x=74.995 //y=2.96 //x2=50.775 //y2=2.96
r650 (  6 8 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=50.69 //y=2.875 //x2=50.775 //y2=2.96
r651 (  5 6 ) resistor r=0.19084 //w=0.131 //l=0.2 //layer=m1 //thickness=0.36 \
 //x=50.69 //y=2.675 //x2=50.69 //y2=2.875
r652 (  4 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=48.215 //y=2.59 //x2=48.1 //y2=2.59
r653 (  3 5 ) resistor r=0.0698411 //w=0.17 //l=0.120208 //layer=m1 \
 //thickness=0.36 //x=50.605 //y=2.59 //x2=50.69 //y2=2.675
r654 (  3 4 ) resistor r=2.28053 //w=0.131 //l=2.39 //layer=m1 \
 //thickness=0.36 //x=50.605 //y=2.59 //x2=48.215 //y2=2.59
r655 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=42.665 //y=4.07 //x2=42.55 //y2=4.07
r656 (  1 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=47.985 //y=4.07 //x2=48.1 //y2=4.07
r657 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=47.985 //y=4.07 //x2=42.665 //y2=4.07
ends PM_TMRDFFSNQX1\%noxref_13

subckt PM_TMRDFFSNQX1\%D ( 1 2 3 4 11 12 13 14 15 16 17 18 19 20 21 22 23 25 \
 38 49 58 59 60 61 62 63 64 65 66 67 68 69 70 74 76 79 80 84 85 86 87 91 93 96 \
 97 101 102 103 104 108 110 113 114 124 133 142 )
c321 ( 142 0 ) capacitor c=0.0588816f //x=49.95 //y=4.7
c322 ( 133 0 ) capacitor c=0.0588816f //x=25.53 //y=4.7
c323 ( 124 0 ) capacitor c=0.0667949f //x=1.11 //y=4.7
c324 ( 114 0 ) capacitor c=0.0318948f //x=50.285 //y=1.21
c325 ( 113 0 ) capacitor c=0.0187384f //x=50.285 //y=0.865
c326 ( 110 0 ) capacitor c=0.0141798f //x=50.13 //y=1.365
c327 ( 108 0 ) capacitor c=0.0149844f //x=50.13 //y=0.71
c328 ( 104 0 ) capacitor c=0.0813322f //x=49.755 //y=1.915
c329 ( 103 0 ) capacitor c=0.0229267f //x=49.755 //y=1.52
c330 ( 102 0 ) capacitor c=0.0234352f //x=49.755 //y=1.21
c331 ( 101 0 ) capacitor c=0.0199343f //x=49.755 //y=0.865
c332 ( 97 0 ) capacitor c=0.0318948f //x=25.865 //y=1.21
c333 ( 96 0 ) capacitor c=0.0187384f //x=25.865 //y=0.865
c334 ( 93 0 ) capacitor c=0.0141798f //x=25.71 //y=1.365
c335 ( 91 0 ) capacitor c=0.0149844f //x=25.71 //y=0.71
c336 ( 87 0 ) capacitor c=0.0813322f //x=25.335 //y=1.915
c337 ( 86 0 ) capacitor c=0.0229267f //x=25.335 //y=1.52
c338 ( 85 0 ) capacitor c=0.0234352f //x=25.335 //y=1.21
c339 ( 84 0 ) capacitor c=0.0199343f //x=25.335 //y=0.865
c340 ( 80 0 ) capacitor c=0.0318948f //x=1.445 //y=1.21
c341 ( 79 0 ) capacitor c=0.0187384f //x=1.445 //y=0.865
c342 ( 76 0 ) capacitor c=0.0141798f //x=1.29 //y=1.365
c343 ( 74 0 ) capacitor c=0.0149844f //x=1.29 //y=0.71
c344 ( 70 0 ) capacitor c=0.0844059f //x=0.915 //y=1.915
c345 ( 69 0 ) capacitor c=0.0229722f //x=0.915 //y=1.52
c346 ( 68 0 ) capacitor c=0.0234352f //x=0.915 //y=1.21
c347 ( 67 0 ) capacitor c=0.0199343f //x=0.915 //y=0.865
c348 ( 66 0 ) capacitor c=0.110275f //x=50.29 //y=6.02
c349 ( 65 0 ) capacitor c=0.154305f //x=49.85 //y=6.02
c350 ( 64 0 ) capacitor c=0.110275f //x=25.87 //y=6.02
c351 ( 63 0 ) capacitor c=0.154305f //x=25.43 //y=6.02
c352 ( 62 0 ) capacitor c=0.110275f //x=1.45 //y=6.02
c353 ( 61 0 ) capacitor c=0.154305f //x=1.01 //y=6.02
c354 ( 49 0 ) capacitor c=0.0876359f //x=49.95 //y=2.08
c355 ( 38 0 ) capacitor c=0.0903622f //x=25.53 //y=2.08
c356 ( 25 0 ) capacitor c=0.111725f //x=1.11 //y=2.08
c357 ( 4 0 ) capacitor c=0.00583987f //x=25.645 //y=2.96
c358 ( 3 0 ) capacitor c=0.373149f //x=49.835 //y=2.96
c359 ( 2 0 ) capacitor c=0.0150814f //x=1.225 //y=2.96
c360 ( 1 0 ) capacitor c=0.470661f //x=25.415 //y=2.96
r361 (  140 142 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=49.85 //y=4.7 //x2=49.95 //y2=4.7
r362 (  131 133 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=25.43 //y=4.7 //x2=25.53 //y2=4.7
r363 (  122 124 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.7 //x2=1.11 //y2=4.7
r364 (  115 142 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=50.29 //y=4.865 //x2=49.95 //y2=4.7
r365 (  114 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.285 //y=1.21 //x2=50.245 //y2=1.365
r366 (  113 143 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.285 //y=0.865 //x2=50.245 //y2=0.71
r367 (  113 114 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=50.285 //y=0.865 //x2=50.285 //y2=1.21
r368 (  111 139 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.91 //y=1.365 //x2=49.795 //y2=1.365
r369 (  110 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.13 //y=1.365 //x2=50.245 //y2=1.365
r370 (  109 138 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=49.91 //y=0.71 //x2=49.795 //y2=0.71
r371 (  108 143 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.13 //y=0.71 //x2=50.245 //y2=0.71
r372 (  108 109 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=50.13 //y=0.71 //x2=49.91 //y2=0.71
r373 (  105 140 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=49.85 //y=4.865 //x2=49.85 //y2=4.7
r374 (  104 137 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=49.755 //y=1.915 //x2=49.95 //y2=2.08
r375 (  103 139 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.755 //y=1.52 //x2=49.795 //y2=1.365
r376 (  103 104 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=49.755 //y=1.52 //x2=49.755 //y2=1.915
r377 (  102 139 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.755 //y=1.21 //x2=49.795 //y2=1.365
r378 (  101 138 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=49.755 //y=0.865 //x2=49.795 //y2=0.71
r379 (  101 102 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=49.755 //y=0.865 //x2=49.755 //y2=1.21
r380 (  98 133 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=25.87 //y=4.865 //x2=25.53 //y2=4.7
r381 (  97 135 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.865 //y=1.21 //x2=25.825 //y2=1.365
r382 (  96 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.865 //y=0.865 //x2=25.825 //y2=0.71
r383 (  96 97 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=25.865 //y=0.865 //x2=25.865 //y2=1.21
r384 (  94 130 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.49 //y=1.365 //x2=25.375 //y2=1.365
r385 (  93 135 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.71 //y=1.365 //x2=25.825 //y2=1.365
r386 (  92 129 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.49 //y=0.71 //x2=25.375 //y2=0.71
r387 (  91 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=25.71 //y=0.71 //x2=25.825 //y2=0.71
r388 (  91 92 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=25.71 //y=0.71 //x2=25.49 //y2=0.71
r389 (  88 131 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=25.43 //y=4.865 //x2=25.43 //y2=4.7
r390 (  87 128 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=25.335 //y=1.915 //x2=25.53 //y2=2.08
r391 (  86 130 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.335 //y=1.52 //x2=25.375 //y2=1.365
r392 (  86 87 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=25.335 //y=1.52 //x2=25.335 //y2=1.915
r393 (  85 130 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.335 //y=1.21 //x2=25.375 //y2=1.365
r394 (  84 129 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=25.335 //y=0.865 //x2=25.375 //y2=0.71
r395 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=25.335 //y=0.865 //x2=25.335 //y2=1.21
r396 (  81 124 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=1.45 //y=4.865 //x2=1.11 //y2=4.7
r397 (  80 126 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.21 //x2=1.405 //y2=1.365
r398 (  79 125 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.405 //y2=0.71
r399 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.865 //x2=1.445 //y2=1.21
r400 (  77 121 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.365 //x2=0.955 //y2=1.365
r401 (  76 126 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.365 //x2=1.405 //y2=1.365
r402 (  75 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.71 //x2=0.955 //y2=0.71
r403 (  74 125 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.405 //y2=0.71
r404 (  74 75 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.71 //x2=1.07 //y2=0.71
r405 (  71 122 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.01 //y=4.865 //x2=1.01 //y2=4.7
r406 (  70 119 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r407 (  69 121 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.955 //y2=1.365
r408 (  69 70 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.52 //x2=0.915 //y2=1.915
r409 (  68 121 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.21 //x2=0.955 //y2=1.365
r410 (  67 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.955 //y2=0.71
r411 (  67 68 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.865 //x2=0.915 //y2=1.21
r412 (  66 115 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=50.29 //y=6.02 //x2=50.29 //y2=4.865
r413 (  65 105 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=49.85 //y=6.02 //x2=49.85 //y2=4.865
r414 (  64 98 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=25.87 //y=6.02 //x2=25.87 //y2=4.865
r415 (  63 88 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=25.43 //y=6.02 //x2=25.43 //y2=4.865
r416 (  62 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.02 //x2=1.45 //y2=4.865
r417 (  61 71 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.02 //x2=1.01 //y2=4.865
r418 (  60 110 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=50.02 //y=1.365 //x2=50.13 //y2=1.365
r419 (  60 111 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=50.02 //y=1.365 //x2=49.91 //y2=1.365
r420 (  59 93 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.6 //y=1.365 //x2=25.71 //y2=1.365
r421 (  59 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=25.6 //y=1.365 //x2=25.49 //y2=1.365
r422 (  58 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.29 //y2=1.365
r423 (  58 77 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.365 //x2=1.07 //y2=1.365
r424 (  56 142 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=49.95 //y=4.7 //x2=49.95 //y2=4.7
r425 (  49 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=49.95 //y=2.08 //x2=49.95 //y2=2.08
r426 (  46 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=25.53 //y=4.7 //x2=25.53 //y2=4.7
r427 (  38 128 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=25.53 //y=2.08 //x2=25.53 //y2=2.08
r428 (  35 124 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r429 (  25 119 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r430 (  23 56 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=49.95 //y=4.07 //x2=49.95 //y2=4.7
r431 (  22 23 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=49.95 //y=3.7 //x2=49.95 //y2=4.07
r432 (  21 22 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=49.95 //y=2.96 //x2=49.95 //y2=3.7
r433 (  21 49 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li \
 //thickness=0.1 //x=49.95 //y=2.96 //x2=49.95 //y2=2.08
r434 (  20 46 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=25.53 //y=4.07 //x2=25.53 //y2=4.7
r435 (  19 20 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=25.53 //y=3.7 //x2=25.53 //y2=4.07
r436 (  18 19 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=25.53 //y=2.96 //x2=25.53 //y2=3.7
r437 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=25.53 //y=2.59 //x2=25.53 //y2=2.96
r438 (  17 38 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=25.53 //y=2.59 //x2=25.53 //y2=2.08
r439 (  16 35 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.44 //x2=1.11 //y2=4.7
r440 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.07 //x2=1.11 //y2=4.44
r441 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=3.7 //x2=1.11 //y2=4.07
r442 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=3.33 //x2=1.11 //y2=3.7
r443 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.96 //x2=1.11 //y2=3.33
r444 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.59 //x2=1.11 //y2=2.96
r445 (  11 25 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.59 //x2=1.11 //y2=2.08
r446 (  10 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=49.95 //y=2.96 //x2=49.95 //y2=2.96
r447 (  8 18 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=25.53 //y=2.96 //x2=25.53 //y2=2.96
r448 (  6 12 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.11 //y=2.96 //x2=1.11 //y2=2.96
r449 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=25.645 //y=2.96 //x2=25.53 //y2=2.96
r450 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=49.835 //y=2.96 //x2=49.95 //y2=2.96
r451 (  3 4 ) resistor r=23.0821 //w=0.131 //l=24.19 //layer=m1 \
 //thickness=0.36 //x=49.835 //y=2.96 //x2=25.645 //y2=2.96
r452 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.225 //y=2.96 //x2=1.11 //y2=2.96
r453 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=25.415 //y=2.96 //x2=25.53 //y2=2.96
r454 (  1 2 ) resistor r=23.0821 //w=0.131 //l=24.19 //layer=m1 \
 //thickness=0.36 //x=25.415 //y=2.96 //x2=1.225 //y2=2.96
ends PM_TMRDFFSNQX1\%D

subckt PM_TMRDFFSNQX1\%noxref_15 ( 1 2 3 4 17 18 29 31 32 36 38 46 53 54 55 56 \
 57 58 59 60 61 62 63 64 66 72 73 74 75 79 80 81 82 83 85 91 92 93 94 114 116 \
 117 )
c237 ( 117 0 ) capacitor c=0.0220291f //x=50.805 //y=5.02
c238 ( 116 0 ) capacitor c=0.0217503f //x=49.925 //y=5.02
c239 ( 114 0 ) capacitor c=0.0084702f //x=50.8 //y=0.905
c240 ( 94 0 ) capacitor c=0.0556143f //x=58.365 //y=4.79
c241 ( 93 0 ) capacitor c=0.0293157f //x=58.655 //y=4.79
c242 ( 92 0 ) capacitor c=0.0347816f //x=58.32 //y=1.22
c243 ( 91 0 ) capacitor c=0.0187487f //x=58.32 //y=0.875
c244 ( 85 0 ) capacitor c=0.0137055f //x=58.165 //y=1.375
c245 ( 83 0 ) capacitor c=0.0149861f //x=58.165 //y=0.72
c246 ( 82 0 ) capacitor c=0.096037f //x=57.79 //y=1.915
c247 ( 81 0 ) capacitor c=0.0228993f //x=57.79 //y=1.53
c248 ( 80 0 ) capacitor c=0.0234352f //x=57.79 //y=1.22
c249 ( 79 0 ) capacitor c=0.0198724f //x=57.79 //y=0.875
c250 ( 75 0 ) capacitor c=0.0557698f //x=53.555 //y=4.79
c251 ( 74 0 ) capacitor c=0.0293157f //x=53.845 //y=4.79
c252 ( 73 0 ) capacitor c=0.0347816f //x=53.51 //y=1.22
c253 ( 72 0 ) capacitor c=0.0187487f //x=53.51 //y=0.875
c254 ( 66 0 ) capacitor c=0.0137055f //x=53.355 //y=1.375
c255 ( 64 0 ) capacitor c=0.0149861f //x=53.355 //y=0.72
c256 ( 63 0 ) capacitor c=0.096037f //x=52.98 //y=1.915
c257 ( 62 0 ) capacitor c=0.0228993f //x=52.98 //y=1.53
c258 ( 61 0 ) capacitor c=0.0234352f //x=52.98 //y=1.22
c259 ( 60 0 ) capacitor c=0.0198724f //x=52.98 //y=0.875
c260 ( 59 0 ) capacitor c=0.110114f //x=58.73 //y=6.02
c261 ( 58 0 ) capacitor c=0.158956f //x=58.29 //y=6.02
c262 ( 57 0 ) capacitor c=0.110114f //x=53.92 //y=6.02
c263 ( 56 0 ) capacitor c=0.158956f //x=53.48 //y=6.02
c264 ( 53 0 ) capacitor c=0.00211606f //x=50.95 //y=5.2
c265 ( 46 0 ) capacitor c=0.0943831f //x=58.09 //y=2.08
c266 ( 38 0 ) capacitor c=0.0969368f //x=53.28 //y=2.08
c267 ( 36 0 ) capacitor c=0.104747f //x=51.43 //y=2.59
c268 ( 32 0 ) capacitor c=0.00404073f //x=51.075 //y=1.655
c269 ( 31 0 ) capacitor c=0.0122201f //x=51.345 //y=1.655
c270 ( 29 0 ) capacitor c=0.0137995f //x=51.345 //y=5.2
c271 ( 18 0 ) capacitor c=0.00251635f //x=50.155 //y=5.2
c272 ( 17 0 ) capacitor c=0.0143649f //x=50.865 //y=5.2
c273 ( 4 0 ) capacitor c=0.00673266f //x=53.545 //y=2.59
c274 ( 3 0 ) capacitor c=0.0686809f //x=57.975 //y=2.59
c275 ( 2 0 ) capacitor c=0.00515785f //x=51.545 //y=2.59
c276 ( 1 0 ) capacitor c=0.0230071f //x=53.135 //y=2.59
r277 (  93 95 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=58.655 //y=4.79 //x2=58.73 //y2=4.865
r278 (  93 94 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=58.655 //y=4.79 //x2=58.365 //y2=4.79
r279 (  92 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.32 //y=1.22 //x2=58.28 //y2=1.375
r280 (  91 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.32 //y=0.875 //x2=58.28 //y2=0.72
r281 (  91 92 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=58.32 //y=0.875 //x2=58.32 //y2=1.22
r282 (  88 94 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=58.29 //y=4.865 //x2=58.365 //y2=4.79
r283 (  88 111 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=58.29 //y=4.865 //x2=58.09 //y2=4.7
r284 (  86 107 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=57.945 //y=1.375 //x2=57.83 //y2=1.375
r285 (  85 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.165 //y=1.375 //x2=58.28 //y2=1.375
r286 (  84 106 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=57.945 //y=0.72 //x2=57.83 //y2=0.72
r287 (  83 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.165 //y=0.72 //x2=58.28 //y2=0.72
r288 (  83 84 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=58.165 //y=0.72 //x2=57.945 //y2=0.72
r289 (  82 109 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=57.79 //y=1.915 //x2=58.09 //y2=2.08
r290 (  81 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=57.79 //y=1.53 //x2=57.83 //y2=1.375
r291 (  81 82 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=57.79 //y=1.53 //x2=57.79 //y2=1.915
r292 (  80 107 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=57.79 //y=1.22 //x2=57.83 //y2=1.375
r293 (  79 106 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=57.79 //y=0.875 //x2=57.83 //y2=0.72
r294 (  79 80 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=57.79 //y=0.875 //x2=57.79 //y2=1.22
r295 (  74 76 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=53.845 //y=4.79 //x2=53.92 //y2=4.865
r296 (  74 75 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=53.845 //y=4.79 //x2=53.555 //y2=4.79
r297 (  73 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.51 //y=1.22 //x2=53.47 //y2=1.375
r298 (  72 104 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.51 //y=0.875 //x2=53.47 //y2=0.72
r299 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=53.51 //y=0.875 //x2=53.51 //y2=1.22
r300 (  69 75 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=53.48 //y=4.865 //x2=53.555 //y2=4.79
r301 (  69 103 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=53.48 //y=4.865 //x2=53.28 //y2=4.7
r302 (  67 99 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.135 //y=1.375 //x2=53.02 //y2=1.375
r303 (  66 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.355 //y=1.375 //x2=53.47 //y2=1.375
r304 (  65 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.135 //y=0.72 //x2=53.02 //y2=0.72
r305 (  64 104 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=53.355 //y=0.72 //x2=53.47 //y2=0.72
r306 (  64 65 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=53.355 //y=0.72 //x2=53.135 //y2=0.72
r307 (  63 101 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=52.98 //y=1.915 //x2=53.28 //y2=2.08
r308 (  62 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.98 //y=1.53 //x2=53.02 //y2=1.375
r309 (  62 63 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=52.98 //y=1.53 //x2=52.98 //y2=1.915
r310 (  61 99 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.98 //y=1.22 //x2=53.02 //y2=1.375
r311 (  60 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=52.98 //y=0.875 //x2=53.02 //y2=0.72
r312 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=52.98 //y=0.875 //x2=52.98 //y2=1.22
r313 (  59 95 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=58.73 //y=6.02 //x2=58.73 //y2=4.865
r314 (  58 88 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=58.29 //y=6.02 //x2=58.29 //y2=4.865
r315 (  57 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=53.92 //y=6.02 //x2=53.92 //y2=4.865
r316 (  56 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=53.48 //y=6.02 //x2=53.48 //y2=4.865
r317 (  55 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=58.055 //y=1.375 //x2=58.165 //y2=1.375
r318 (  55 86 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=58.055 //y=1.375 //x2=57.945 //y2=1.375
r319 (  54 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=53.245 //y=1.375 //x2=53.355 //y2=1.375
r320 (  54 67 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=53.245 //y=1.375 //x2=53.135 //y2=1.375
r321 (  51 111 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=58.09 //y=4.7 //x2=58.09 //y2=4.7
r322 (  49 51 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=58.09 //y=2.59 //x2=58.09 //y2=4.7
r323 (  46 109 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=58.09 //y=2.08 //x2=58.09 //y2=2.08
r324 (  46 49 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=58.09 //y=2.08 //x2=58.09 //y2=2.59
r325 (  43 103 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=53.28 //y=4.7 //x2=53.28 //y2=4.7
r326 (  41 43 ) resistor r=144.77 //w=0.187 //l=2.115 //layer=li \
 //thickness=0.1 //x=53.28 //y=2.585 //x2=53.28 //y2=4.7
r327 (  38 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=53.28 //y=2.08 //x2=53.28 //y2=2.08
r328 (  38 41 ) resistor r=34.5668 //w=0.187 //l=0.505 //layer=li \
 //thickness=0.1 //x=53.28 //y=2.08 //x2=53.28 //y2=2.585
r329 (  34 36 ) resistor r=172.834 //w=0.187 //l=2.525 //layer=li \
 //thickness=0.1 //x=51.43 //y=5.115 //x2=51.43 //y2=2.59
r330 (  33 36 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=51.43 //y=1.74 //x2=51.43 //y2=2.59
r331 (  31 33 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=51.345 //y=1.655 //x2=51.43 //y2=1.74
r332 (  31 32 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=51.345 //y=1.655 //x2=51.075 //y2=1.655
r333 (  30 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=51.035 //y=5.2 //x2=50.95 //y2=5.2
r334 (  29 34 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=51.345 //y=5.2 //x2=51.43 //y2=5.115
r335 (  29 30 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=51.345 //y=5.2 //x2=51.035 //y2=5.2
r336 (  25 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=50.99 //y=1.57 //x2=51.075 //y2=1.655
r337 (  25 114 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=50.99 //y=1.57 //x2=50.99 //y2=1
r338 (  19 53 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.95 //y=5.285 //x2=50.95 //y2=5.2
r339 (  19 117 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=50.95 //y=5.285 //x2=50.95 //y2=5.725
r340 (  17 53 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=50.865 //y=5.2 //x2=50.95 //y2=5.2
r341 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=50.865 //y=5.2 //x2=50.155 //y2=5.2
r342 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=50.07 //y=5.285 //x2=50.155 //y2=5.2
r343 (  11 116 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=50.07 //y=5.285 //x2=50.07 //y2=5.725
r344 (  10 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=58.09 //y=2.59 //x2=58.09 //y2=2.59
r345 (  8 41 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=53.28 //y=2.585 //x2=53.28 //y2=2.585
r346 (  6 36 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=51.43 //y=2.59 //x2=51.43 //y2=2.59
r347 (  4 8 ) resistor r=0.164988 //w=0.206 //l=0.267488 //layer=m1 \
 //thickness=0.36 //x=53.545 //y=2.59 //x2=53.28 //y2=2.585
r348 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=57.975 //y=2.59 //x2=58.09 //y2=2.59
r349 (  3 4 ) resistor r=4.2271 //w=0.131 //l=4.43 //layer=m1 //thickness=0.36 \
 //x=57.975 //y=2.59 //x2=53.545 //y2=2.59
r350 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=51.545 //y=2.59 //x2=51.43 //y2=2.59
r351 (  1 8 ) resistor r=0.0921728 //w=0.206 //l=0.147479 //layer=m1 \
 //thickness=0.36 //x=53.135 //y=2.59 //x2=53.28 //y2=2.585
r352 (  1 2 ) resistor r=1.51718 //w=0.131 //l=1.59 //layer=m1 \
 //thickness=0.36 //x=53.135 //y=2.59 //x2=51.545 //y2=2.59
ends PM_TMRDFFSNQX1\%noxref_15

subckt PM_TMRDFFSNQX1\%noxref_16 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 \
 54 55 56 57 61 63 66 67 77 80 82 83 84 )
c164 ( 84 0 ) capacitor c=0.023087f //x=60.125 //y=5.02
c165 ( 83 0 ) capacitor c=0.023519f //x=59.245 //y=5.02
c166 ( 82 0 ) capacitor c=0.0224735f //x=58.365 //y=5.02
c167 ( 80 0 ) capacitor c=0.00872971f //x=60.375 //y=0.915
c168 ( 77 0 ) capacitor c=0.0588816f //x=62.9 //y=4.7
c169 ( 67 0 ) capacitor c=0.0318948f //x=63.235 //y=1.21
c170 ( 66 0 ) capacitor c=0.0187384f //x=63.235 //y=0.865
c171 ( 63 0 ) capacitor c=0.0141798f //x=63.08 //y=1.365
c172 ( 61 0 ) capacitor c=0.0149844f //x=63.08 //y=0.71
c173 ( 57 0 ) capacitor c=0.0813322f //x=62.705 //y=1.915
c174 ( 56 0 ) capacitor c=0.0229267f //x=62.705 //y=1.52
c175 ( 55 0 ) capacitor c=0.0234352f //x=62.705 //y=1.21
c176 ( 54 0 ) capacitor c=0.0199343f //x=62.705 //y=0.865
c177 ( 53 0 ) capacitor c=0.110275f //x=63.24 //y=6.02
c178 ( 52 0 ) capacitor c=0.154305f //x=62.8 //y=6.02
c179 ( 50 0 ) capacitor c=0.00106608f //x=60.27 //y=5.155
c180 ( 49 0 ) capacitor c=0.00207319f //x=59.39 //y=5.155
c181 ( 42 0 ) capacitor c=0.0839295f //x=62.9 //y=2.08
c182 ( 40 0 ) capacitor c=0.10402f //x=61.05 //y=2.59
c183 ( 36 0 ) capacitor c=0.00398962f //x=60.65 //y=1.665
c184 ( 35 0 ) capacitor c=0.0137288f //x=60.965 //y=1.665
c185 ( 29 0 ) capacitor c=0.0284988f //x=60.965 //y=5.155
c186 ( 21 0 ) capacitor c=0.0176454f //x=60.185 //y=5.155
c187 ( 14 0 ) capacitor c=0.00332903f //x=58.595 //y=5.155
c188 ( 13 0 ) capacitor c=0.0148427f //x=59.305 //y=5.155
c189 ( 2 0 ) capacitor c=0.00808366f //x=61.165 //y=2.59
c190 ( 1 0 ) capacitor c=0.0353429f //x=62.785 //y=2.59
r191 (  75 77 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=62.8 //y=4.7 //x2=62.9 //y2=4.7
r192 (  68 77 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=63.24 //y=4.865 //x2=62.9 //y2=4.7
r193 (  67 79 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.235 //y=1.21 //x2=63.195 //y2=1.365
r194 (  66 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.235 //y=0.865 //x2=63.195 //y2=0.71
r195 (  66 67 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=63.235 //y=0.865 //x2=63.235 //y2=1.21
r196 (  64 74 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=62.86 //y=1.365 //x2=62.745 //y2=1.365
r197 (  63 79 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.08 //y=1.365 //x2=63.195 //y2=1.365
r198 (  62 73 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=62.86 //y=0.71 //x2=62.745 //y2=0.71
r199 (  61 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.08 //y=0.71 //x2=63.195 //y2=0.71
r200 (  61 62 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=63.08 //y=0.71 //x2=62.86 //y2=0.71
r201 (  58 75 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=62.8 //y=4.865 //x2=62.8 //y2=4.7
r202 (  57 72 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=62.705 //y=1.915 //x2=62.9 //y2=2.08
r203 (  56 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.705 //y=1.52 //x2=62.745 //y2=1.365
r204 (  56 57 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=62.705 //y=1.52 //x2=62.705 //y2=1.915
r205 (  55 74 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.705 //y=1.21 //x2=62.745 //y2=1.365
r206 (  54 73 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=62.705 //y=0.865 //x2=62.745 //y2=0.71
r207 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=62.705 //y=0.865 //x2=62.705 //y2=1.21
r208 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=63.24 //y=6.02 //x2=63.24 //y2=4.865
r209 (  52 58 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=62.8 //y=6.02 //x2=62.8 //y2=4.865
r210 (  51 63 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=62.97 //y=1.365 //x2=63.08 //y2=1.365
r211 (  51 64 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=62.97 //y=1.365 //x2=62.86 //y2=1.365
r212 (  47 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=62.9 //y=4.7 //x2=62.9 //y2=4.7
r213 (  45 47 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=62.9 //y=2.59 //x2=62.9 //y2=4.7
r214 (  42 72 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=62.9 //y=2.08 //x2=62.9 //y2=2.08
r215 (  42 45 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=62.9 //y=2.08 //x2=62.9 //y2=2.59
r216 (  38 40 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=61.05 //y=5.07 //x2=61.05 //y2=2.59
r217 (  37 40 ) resistor r=57.4973 //w=0.187 //l=0.84 //layer=li \
 //thickness=0.1 //x=61.05 //y=1.75 //x2=61.05 //y2=2.59
r218 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=60.965 //y=1.665 //x2=61.05 //y2=1.75
r219 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=60.965 //y=1.665 //x2=60.65 //y2=1.665
r220 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=60.565 //y=1.58 //x2=60.65 //y2=1.665
r221 (  31 80 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=60.565 //y=1.58 //x2=60.565 //y2=1.01
r222 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.355 //y=5.155 //x2=60.27 //y2=5.155
r223 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=60.965 //y=5.155 //x2=61.05 //y2=5.07
r224 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=60.965 //y=5.155 //x2=60.355 //y2=5.155
r225 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.27 //y=5.24 //x2=60.27 //y2=5.155
r226 (  23 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=60.27 //y=5.24 //x2=60.27 //y2=5.725
r227 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.475 //y=5.155 //x2=59.39 //y2=5.155
r228 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=60.185 //y=5.155 //x2=60.27 //y2=5.155
r229 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=60.185 //y=5.155 //x2=59.475 //y2=5.155
r230 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.39 //y=5.24 //x2=59.39 //y2=5.155
r231 (  15 83 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=59.39 //y=5.24 //x2=59.39 //y2=5.725
r232 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.305 //y=5.155 //x2=59.39 //y2=5.155
r233 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=59.305 //y=5.155 //x2=58.595 //y2=5.155
r234 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=58.51 //y=5.24 //x2=58.595 //y2=5.155
r235 (  7 82 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=58.51 //y=5.24 //x2=58.51 //y2=5.725
r236 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=62.9 //y=2.59 //x2=62.9 //y2=2.59
r237 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=61.05 //y=2.59 //x2=61.05 //y2=2.59
r238 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=61.165 //y=2.59 //x2=61.05 //y2=2.59
r239 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=62.785 //y=2.59 //x2=62.9 //y2=2.59
r240 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=62.785 //y=2.59 //x2=61.165 //y2=2.59
ends PM_TMRDFFSNQX1\%noxref_16

subckt PM_TMRDFFSNQX1\%CLK ( 1 2 3 4 5 6 7 8 9 10 23 24 25 26 27 28 29 30 31 \
 32 33 34 35 36 37 39 49 51 58 66 68 74 82 84 95 96 97 98 99 100 101 102 103 \
 104 105 106 107 108 109 110 111 112 113 114 115 117 123 124 125 126 127 132 \
 133 134 139 141 143 149 150 151 152 153 155 161 162 163 164 165 170 171 172 \
 177 179 181 187 188 189 190 191 193 199 200 201 202 203 208 209 210 215 217 \
 219 225 226 230 239 240 243 254 263 264 267 278 287 288 291 )
c755 ( 291 0 ) capacitor c=0.0331838f //x=63.67 //y=4.7
c756 ( 288 0 ) capacitor c=0.0279499f //x=63.64 //y=1.915
c757 ( 287 0 ) capacitor c=0.0421676f //x=63.64 //y=2.08
c758 ( 278 0 ) capacitor c=0.0334842f //x=54.39 //y=4.7
c759 ( 267 0 ) capacitor c=0.0331706f //x=39.25 //y=4.7
c760 ( 264 0 ) capacitor c=0.0279499f //x=39.22 //y=1.915
c761 ( 263 0 ) capacitor c=0.0421676f //x=39.22 //y=2.08
c762 ( 254 0 ) capacitor c=0.0334842f //x=29.97 //y=4.7
c763 ( 243 0 ) capacitor c=0.0331706f //x=14.83 //y=4.7
c764 ( 240 0 ) capacitor c=0.0279499f //x=14.8 //y=1.915
c765 ( 239 0 ) capacitor c=0.0421676f //x=14.8 //y=2.08
c766 ( 230 0 ) capacitor c=0.0334842f //x=5.55 //y=4.7
c767 ( 226 0 ) capacitor c=0.0429696f //x=64.205 //y=1.25
c768 ( 225 0 ) capacitor c=0.0192208f //x=64.205 //y=0.905
c769 ( 219 0 ) capacitor c=0.0148884f //x=64.05 //y=1.405
c770 ( 217 0 ) capacitor c=0.0157803f //x=64.05 //y=0.75
c771 ( 215 0 ) capacitor c=0.0299681f //x=64.045 //y=4.79
c772 ( 210 0 ) capacitor c=0.0205163f //x=63.675 //y=1.56
c773 ( 209 0 ) capacitor c=0.0168481f //x=63.675 //y=1.25
c774 ( 208 0 ) capacitor c=0.0174783f //x=63.675 //y=0.905
c775 ( 203 0 ) capacitor c=0.0245352f //x=54.725 //y=4.79
c776 ( 202 0 ) capacitor c=0.0825763f //x=54.48 //y=1.915
c777 ( 201 0 ) capacitor c=0.0170266f //x=54.48 //y=1.45
c778 ( 200 0 ) capacitor c=0.018609f //x=54.48 //y=1.22
c779 ( 199 0 ) capacitor c=0.0187309f //x=54.48 //y=0.91
c780 ( 193 0 ) capacitor c=0.014725f //x=54.325 //y=1.375
c781 ( 191 0 ) capacitor c=0.0146567f //x=54.325 //y=0.755
c782 ( 190 0 ) capacitor c=0.0335408f //x=53.955 //y=1.22
c783 ( 189 0 ) capacitor c=0.0173761f //x=53.955 //y=0.91
c784 ( 188 0 ) capacitor c=0.0429696f //x=39.785 //y=1.25
c785 ( 187 0 ) capacitor c=0.0192208f //x=39.785 //y=0.905
c786 ( 181 0 ) capacitor c=0.0148884f //x=39.63 //y=1.405
c787 ( 179 0 ) capacitor c=0.0157803f //x=39.63 //y=0.75
c788 ( 177 0 ) capacitor c=0.0295235f //x=39.625 //y=4.79
c789 ( 172 0 ) capacitor c=0.0205163f //x=39.255 //y=1.56
c790 ( 171 0 ) capacitor c=0.0168481f //x=39.255 //y=1.25
c791 ( 170 0 ) capacitor c=0.0174783f //x=39.255 //y=0.905
c792 ( 165 0 ) capacitor c=0.0245352f //x=30.305 //y=4.79
c793 ( 164 0 ) capacitor c=0.0825763f //x=30.06 //y=1.915
c794 ( 163 0 ) capacitor c=0.0170266f //x=30.06 //y=1.45
c795 ( 162 0 ) capacitor c=0.018609f //x=30.06 //y=1.22
c796 ( 161 0 ) capacitor c=0.0187309f //x=30.06 //y=0.91
c797 ( 155 0 ) capacitor c=0.014725f //x=29.905 //y=1.375
c798 ( 153 0 ) capacitor c=0.0146567f //x=29.905 //y=0.755
c799 ( 152 0 ) capacitor c=0.0335408f //x=29.535 //y=1.22
c800 ( 151 0 ) capacitor c=0.0173761f //x=29.535 //y=0.91
c801 ( 150 0 ) capacitor c=0.0429696f //x=15.365 //y=1.25
c802 ( 149 0 ) capacitor c=0.0192208f //x=15.365 //y=0.905
c803 ( 143 0 ) capacitor c=0.0148884f //x=15.21 //y=1.405
c804 ( 141 0 ) capacitor c=0.0157803f //x=15.21 //y=0.75
c805 ( 139 0 ) capacitor c=0.0295235f //x=15.205 //y=4.79
c806 ( 134 0 ) capacitor c=0.0205163f //x=14.835 //y=1.56
c807 ( 133 0 ) capacitor c=0.0168481f //x=14.835 //y=1.25
c808 ( 132 0 ) capacitor c=0.0174783f //x=14.835 //y=0.905
c809 ( 127 0 ) capacitor c=0.0245352f //x=5.885 //y=4.79
c810 ( 126 0 ) capacitor c=0.0826403f //x=5.64 //y=1.915
c811 ( 125 0 ) capacitor c=0.0170266f //x=5.64 //y=1.45
c812 ( 124 0 ) capacitor c=0.018609f //x=5.64 //y=1.22
c813 ( 123 0 ) capacitor c=0.0187309f //x=5.64 //y=0.91
c814 ( 117 0 ) capacitor c=0.014725f //x=5.485 //y=1.375
c815 ( 115 0 ) capacitor c=0.0146567f //x=5.485 //y=0.755
c816 ( 114 0 ) capacitor c=0.0335408f //x=5.115 //y=1.22
c817 ( 113 0 ) capacitor c=0.0173761f //x=5.115 //y=0.91
c818 ( 112 0 ) capacitor c=0.15358f //x=64.12 //y=6.02
c819 ( 111 0 ) capacitor c=0.110281f //x=63.68 //y=6.02
c820 ( 110 0 ) capacitor c=0.110114f //x=54.8 //y=6.02
c821 ( 109 0 ) capacitor c=0.11012f //x=54.36 //y=6.02
c822 ( 108 0 ) capacitor c=0.15358f //x=39.7 //y=6.02
c823 ( 107 0 ) capacitor c=0.110281f //x=39.26 //y=6.02
c824 ( 106 0 ) capacitor c=0.110114f //x=30.38 //y=6.02
c825 ( 105 0 ) capacitor c=0.11012f //x=29.94 //y=6.02
c826 ( 104 0 ) capacitor c=0.15358f //x=15.28 //y=6.02
c827 ( 103 0 ) capacitor c=0.110281f //x=14.84 //y=6.02
c828 ( 102 0 ) capacitor c=0.110114f //x=5.96 //y=6.02
c829 ( 101 0 ) capacitor c=0.11012f //x=5.52 //y=6.02
c830 ( 84 0 ) capacitor c=0.0691208f //x=63.64 //y=2.08
c831 ( 82 0 ) capacitor c=0.00369614f //x=63.64 //y=4.535
c832 ( 74 0 ) capacitor c=0.0900341f //x=54.39 //y=2.08
c833 ( 68 0 ) capacitor c=0.0687295f //x=39.22 //y=2.08
c834 ( 66 0 ) capacitor c=0.00369614f //x=39.22 //y=4.535
c835 ( 58 0 ) capacitor c=0.0900341f //x=29.97 //y=2.08
c836 ( 51 0 ) capacitor c=0.0706177f //x=14.8 //y=2.08
c837 ( 49 0 ) capacitor c=0.00369614f //x=14.8 //y=4.535
c838 ( 39 0 ) capacitor c=0.0953538f //x=5.55 //y=2.08
c839 ( 10 0 ) capacitor c=0.00697397f //x=54.505 //y=4.44
c840 ( 9 0 ) capacitor c=0.213217f //x=63.525 //y=4.44
c841 ( 8 0 ) capacitor c=0.00680508f //x=39.335 //y=4.44
c842 ( 7 0 ) capacitor c=0.354845f //x=54.275 //y=4.44
c843 ( 6 0 ) capacitor c=0.00697397f //x=30.085 //y=4.44
c844 ( 5 0 ) capacitor c=0.201328f //x=39.105 //y=4.44
c845 ( 4 0 ) capacitor c=0.00680508f //x=14.915 //y=4.44
c846 ( 3 0 ) capacitor c=0.368123f //x=29.855 //y=4.44
c847 ( 2 0 ) capacitor c=0.0154455f //x=5.665 //y=4.44
c848 ( 1 0 ) capacitor c=0.201328f //x=14.685 //y=4.44
r849 (  293 294 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=63.67 //y=4.79 //x2=63.67 //y2=4.865
r850 (  291 293 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=63.67 //y=4.7 //x2=63.67 //y2=4.79
r851 (  287 288 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=63.64 //y=2.08 //x2=63.64 //y2=1.915
r852 (  280 281 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=54.39 //y=4.79 //x2=54.39 //y2=4.865
r853 (  278 280 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=54.39 //y=4.7 //x2=54.39 //y2=4.79
r854 (  269 270 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=39.25 //y=4.79 //x2=39.25 //y2=4.865
r855 (  267 269 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=39.25 //y=4.7 //x2=39.25 //y2=4.79
r856 (  263 264 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=39.22 //y=2.08 //x2=39.22 //y2=1.915
r857 (  256 257 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=29.97 //y=4.79 //x2=29.97 //y2=4.865
r858 (  254 256 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=29.97 //y=4.7 //x2=29.97 //y2=4.79
r859 (  245 246 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=14.83 //y=4.79 //x2=14.83 //y2=4.865
r860 (  243 245 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=14.83 //y=4.7 //x2=14.83 //y2=4.79
r861 (  239 240 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=14.8 //y=2.08 //x2=14.8 //y2=1.915
r862 (  232 233 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=5.55 //y=4.79 //x2=5.55 //y2=4.865
r863 (  230 232 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=5.55 //y=4.7 //x2=5.55 //y2=4.79
r864 (  226 298 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=64.205 //y=1.25 //x2=64.165 //y2=1.405
r865 (  225 297 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=64.205 //y=0.905 //x2=64.165 //y2=0.75
r866 (  225 226 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=64.205 //y=0.905 //x2=64.205 //y2=1.25
r867 (  220 296 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.83 //y=1.405 //x2=63.715 //y2=1.405
r868 (  219 298 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=64.05 //y=1.405 //x2=64.165 //y2=1.405
r869 (  218 295 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=63.83 //y=0.75 //x2=63.715 //y2=0.75
r870 (  217 297 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=64.05 //y=0.75 //x2=64.165 //y2=0.75
r871 (  217 218 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=64.05 //y=0.75 //x2=63.83 //y2=0.75
r872 (  216 293 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=63.805 //y=4.79 //x2=63.67 //y2=4.79
r873 (  215 222 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=64.045 //y=4.79 //x2=64.12 //y2=4.865
r874 (  215 216 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=64.045 //y=4.79 //x2=63.805 //y2=4.79
r875 (  210 296 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.675 //y=1.56 //x2=63.715 //y2=1.405
r876 (  210 288 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=63.675 //y=1.56 //x2=63.675 //y2=1.915
r877 (  209 296 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.675 //y=1.25 //x2=63.715 //y2=1.405
r878 (  208 295 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=63.675 //y=0.905 //x2=63.715 //y2=0.75
r879 (  208 209 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=63.675 //y=0.905 //x2=63.675 //y2=1.25
r880 (  204 280 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=54.525 //y=4.79 //x2=54.39 //y2=4.79
r881 (  203 205 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=54.725 //y=4.79 //x2=54.8 //y2=4.865
r882 (  203 204 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=54.725 //y=4.79 //x2=54.525 //y2=4.79
r883 (  202 285 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=54.48 //y=1.915 //x2=54.405 //y2=2.08
r884 (  201 283 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=54.48 //y=1.45 //x2=54.44 //y2=1.375
r885 (  201 202 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=54.48 //y=1.45 //x2=54.48 //y2=1.915
r886 (  200 283 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.48 //y=1.22 //x2=54.44 //y2=1.375
r887 (  199 282 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=54.48 //y=0.91 //x2=54.44 //y2=0.755
r888 (  199 200 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=54.48 //y=0.91 //x2=54.48 //y2=1.22
r889 (  194 276 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.11 //y=1.375 //x2=53.995 //y2=1.375
r890 (  193 283 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.325 //y=1.375 //x2=54.44 //y2=1.375
r891 (  192 275 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.11 //y=0.755 //x2=53.995 //y2=0.755
r892 (  191 282 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=54.325 //y=0.755 //x2=54.44 //y2=0.755
r893 (  191 192 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=54.325 //y=0.755 //x2=54.11 //y2=0.755
r894 (  190 276 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.955 //y=1.22 //x2=53.995 //y2=1.375
r895 (  189 275 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=53.955 //y=0.91 //x2=53.995 //y2=0.755
r896 (  189 190 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=53.955 //y=0.91 //x2=53.955 //y2=1.22
r897 (  188 274 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.785 //y=1.25 //x2=39.745 //y2=1.405
r898 (  187 273 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.785 //y=0.905 //x2=39.745 //y2=0.75
r899 (  187 188 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=39.785 //y=0.905 //x2=39.785 //y2=1.25
r900 (  182 272 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.41 //y=1.405 //x2=39.295 //y2=1.405
r901 (  181 274 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.63 //y=1.405 //x2=39.745 //y2=1.405
r902 (  180 271 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.41 //y=0.75 //x2=39.295 //y2=0.75
r903 (  179 273 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=39.63 //y=0.75 //x2=39.745 //y2=0.75
r904 (  179 180 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=39.63 //y=0.75 //x2=39.41 //y2=0.75
r905 (  178 269 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=39.385 //y=4.79 //x2=39.25 //y2=4.79
r906 (  177 184 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=39.625 //y=4.79 //x2=39.7 //y2=4.865
r907 (  177 178 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=39.625 //y=4.79 //x2=39.385 //y2=4.79
r908 (  172 272 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.255 //y=1.56 //x2=39.295 //y2=1.405
r909 (  172 264 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=39.255 //y=1.56 //x2=39.255 //y2=1.915
r910 (  171 272 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.255 //y=1.25 //x2=39.295 //y2=1.405
r911 (  170 271 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=39.255 //y=0.905 //x2=39.295 //y2=0.75
r912 (  170 171 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=39.255 //y=0.905 //x2=39.255 //y2=1.25
r913 (  166 256 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=30.105 //y=4.79 //x2=29.97 //y2=4.79
r914 (  165 167 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=30.305 //y=4.79 //x2=30.38 //y2=4.865
r915 (  165 166 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=30.305 //y=4.79 //x2=30.105 //y2=4.79
r916 (  164 261 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=30.06 //y=1.915 //x2=29.985 //y2=2.08
r917 (  163 259 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=30.06 //y=1.45 //x2=30.02 //y2=1.375
r918 (  163 164 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=30.06 //y=1.45 //x2=30.06 //y2=1.915
r919 (  162 259 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.06 //y=1.22 //x2=30.02 //y2=1.375
r920 (  161 258 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=30.06 //y=0.91 //x2=30.02 //y2=0.755
r921 (  161 162 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=30.06 //y=0.91 //x2=30.06 //y2=1.22
r922 (  156 252 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.69 //y=1.375 //x2=29.575 //y2=1.375
r923 (  155 259 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.905 //y=1.375 //x2=30.02 //y2=1.375
r924 (  154 251 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.69 //y=0.755 //x2=29.575 //y2=0.755
r925 (  153 258 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=29.905 //y=0.755 //x2=30.02 //y2=0.755
r926 (  153 154 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=29.905 //y=0.755 //x2=29.69 //y2=0.755
r927 (  152 252 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.535 //y=1.22 //x2=29.575 //y2=1.375
r928 (  151 251 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=29.535 //y=0.91 //x2=29.575 //y2=0.755
r929 (  151 152 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=29.535 //y=0.91 //x2=29.535 //y2=1.22
r930 (  150 250 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.365 //y=1.25 //x2=15.325 //y2=1.405
r931 (  149 249 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.365 //y=0.905 //x2=15.325 //y2=0.75
r932 (  149 150 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=15.365 //y=0.905 //x2=15.365 //y2=1.25
r933 (  144 248 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.99 //y=1.405 //x2=14.875 //y2=1.405
r934 (  143 250 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.21 //y=1.405 //x2=15.325 //y2=1.405
r935 (  142 247 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.99 //y=0.75 //x2=14.875 //y2=0.75
r936 (  141 249 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.21 //y=0.75 //x2=15.325 //y2=0.75
r937 (  141 142 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=15.21 //y=0.75 //x2=14.99 //y2=0.75
r938 (  140 245 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=14.965 //y=4.79 //x2=14.83 //y2=4.79
r939 (  139 146 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.205 //y=4.79 //x2=15.28 //y2=4.865
r940 (  139 140 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=15.205 //y=4.79 //x2=14.965 //y2=4.79
r941 (  134 248 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.835 //y=1.56 //x2=14.875 //y2=1.405
r942 (  134 240 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=14.835 //y=1.56 //x2=14.835 //y2=1.915
r943 (  133 248 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.835 //y=1.25 //x2=14.875 //y2=1.405
r944 (  132 247 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.835 //y=0.905 //x2=14.875 //y2=0.75
r945 (  132 133 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.835 //y=0.905 //x2=14.835 //y2=1.25
r946 (  128 232 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=5.685 //y=4.79 //x2=5.55 //y2=4.79
r947 (  127 129 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.885 //y=4.79 //x2=5.96 //y2=4.865
r948 (  127 128 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=5.885 //y=4.79 //x2=5.685 //y2=4.79
r949 (  126 237 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.915 //x2=5.565 //y2=2.08
r950 (  125 235 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.45 //x2=5.6 //y2=1.375
r951 (  125 126 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.45 //x2=5.64 //y2=1.915
r952 (  124 235 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.64 //y=1.22 //x2=5.6 //y2=1.375
r953 (  123 234 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.64 //y=0.91 //x2=5.6 //y2=0.755
r954 (  123 124 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=5.64 //y=0.91 //x2=5.64 //y2=1.22
r955 (  118 228 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.27 //y=1.375 //x2=5.155 //y2=1.375
r956 (  117 235 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.485 //y=1.375 //x2=5.6 //y2=1.375
r957 (  116 227 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.27 //y=0.755 //x2=5.155 //y2=0.755
r958 (  115 234 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.485 //y=0.755 //x2=5.6 //y2=0.755
r959 (  115 116 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=5.485 //y=0.755 //x2=5.27 //y2=0.755
r960 (  114 228 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.115 //y=1.22 //x2=5.155 //y2=1.375
r961 (  113 227 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.115 //y=0.91 //x2=5.155 //y2=0.755
r962 (  113 114 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=5.115 //y=0.91 //x2=5.115 //y2=1.22
r963 (  112 222 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=64.12 //y=6.02 //x2=64.12 //y2=4.865
r964 (  111 294 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=63.68 //y=6.02 //x2=63.68 //y2=4.865
r965 (  110 205 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=54.8 //y=6.02 //x2=54.8 //y2=4.865
r966 (  109 281 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=54.36 //y=6.02 //x2=54.36 //y2=4.865
r967 (  108 184 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=39.7 //y=6.02 //x2=39.7 //y2=4.865
r968 (  107 270 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=39.26 //y=6.02 //x2=39.26 //y2=4.865
r969 (  106 167 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=30.38 //y=6.02 //x2=30.38 //y2=4.865
r970 (  105 257 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=29.94 //y=6.02 //x2=29.94 //y2=4.865
r971 (  104 146 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.28 //y=6.02 //x2=15.28 //y2=4.865
r972 (  103 246 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.84 //y=6.02 //x2=14.84 //y2=4.865
r973 (  102 129 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.96 //y=6.02 //x2=5.96 //y2=4.865
r974 (  101 233 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.52 //y=6.02 //x2=5.52 //y2=4.865
r975 (  100 219 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=63.94 //y=1.405 //x2=64.05 //y2=1.405
r976 (  100 220 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=63.94 //y=1.405 //x2=63.83 //y2=1.405
r977 (  99 193 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=54.217 //y=1.375 //x2=54.325 //y2=1.375
r978 (  99 194 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=54.217 //y=1.375 //x2=54.11 //y2=1.375
r979 (  98 181 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=39.52 //y=1.405 //x2=39.63 //y2=1.405
r980 (  98 182 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=39.52 //y=1.405 //x2=39.41 //y2=1.405
r981 (  97 155 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=29.797 //y=1.375 //x2=29.905 //y2=1.375
r982 (  97 156 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=29.797 //y=1.375 //x2=29.69 //y2=1.375
r983 (  96 143 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.1 //y=1.405 //x2=15.21 //y2=1.405
r984 (  96 144 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=15.1 //y=1.405 //x2=14.99 //y2=1.405
r985 (  95 117 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=5.377 //y=1.375 //x2=5.485 //y2=1.375
r986 (  95 118 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=5.377 //y=1.375 //x2=5.27 //y2=1.375
r987 (  94 291 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=63.67 //y=4.7 //x2=63.67 //y2=4.7
r988 (  92 267 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=39.25 //y=4.7 //x2=39.25 //y2=4.7
r989 (  90 243 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.83 //y=4.7 //x2=14.83 //y2=4.7
r990 (  84 287 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=63.64 //y=2.08 //x2=63.64 //y2=2.08
r991 (  82 94 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=63.64 //y=4.535 //x2=63.655 //y2=4.7
r992 (  80 278 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=54.39 //y=4.7 //x2=54.39 //y2=4.7
r993 (  74 285 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=54.39 //y=2.08 //x2=54.39 //y2=2.08
r994 (  68 263 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=39.22 //y=2.08 //x2=39.22 //y2=2.08
r995 (  66 92 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=39.22 //y=4.535 //x2=39.235 //y2=4.7
r996 (  64 254 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=29.97 //y=4.7 //x2=29.97 //y2=4.7
r997 (  58 261 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=29.97 //y=2.08 //x2=29.97 //y2=2.08
r998 (  51 239 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.8 //y=2.08 //x2=14.8 //y2=2.08
r999 (  49 90 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=14.8 //y=4.535 //x2=14.815 //y2=4.7
r1000 (  47 230 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.55 //y=4.7 //x2=5.55 //y2=4.7
r1001 (  39 237 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.55 //y=2.08 //x2=5.55 //y2=2.08
r1002 (  37 82 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=63.64 //y=4.44 //x2=63.64 //y2=4.535
r1003 (  36 37 ) resistor r=126.631 //w=0.187 //l=1.85 //layer=li \
 //thickness=0.1 //x=63.64 //y=2.59 //x2=63.64 //y2=4.44
r1004 (  36 84 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=63.64 //y=2.59 //x2=63.64 //y2=2.08
r1005 (  35 80 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=54.39 //y=4.44 //x2=54.39 //y2=4.7
r1006 (  34 35 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=54.39 //y=3.7 //x2=54.39 //y2=4.44
r1007 (  34 74 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=54.39 //y=3.7 //x2=54.39 //y2=2.08
r1008 (  33 66 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=39.22 //y=4.44 //x2=39.22 //y2=4.535
r1009 (  32 33 ) resistor r=126.631 //w=0.187 //l=1.85 //layer=li \
 //thickness=0.1 //x=39.22 //y=2.59 //x2=39.22 //y2=4.44
r1010 (  32 68 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=39.22 //y=2.59 //x2=39.22 //y2=2.08
r1011 (  31 64 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=29.97 //y=4.44 //x2=29.97 //y2=4.7
r1012 (  30 31 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=29.97 //y=3.7 //x2=29.97 //y2=4.44
r1013 (  30 58 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=29.97 //y=3.7 //x2=29.97 //y2=2.08
r1014 (  29 49 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=14.8 //y=4.44 //x2=14.8 //y2=4.535
r1015 (  28 29 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=14.8 //y=3.33 //x2=14.8 //y2=4.44
r1016 (  27 28 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=14.8 //y=2.59 //x2=14.8 //y2=3.33
r1017 (  27 51 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=14.8 //y=2.59 //x2=14.8 //y2=2.08
r1018 (  26 47 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=5.55 //y=4.44 //x2=5.55 //y2=4.7
r1019 (  25 26 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=5.55 //y=3.7 //x2=5.55 //y2=4.44
r1020 (  24 25 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=5.55 //y=3.33 //x2=5.55 //y2=3.7
r1021 (  23 24 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=5.55 //y=2.22 //x2=5.55 //y2=3.33
r1022 (  23 39 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=5.55 //y=2.22 //x2=5.55 //y2=2.08
r1023 (  22 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=63.64 //y=4.44 //x2=63.64 //y2=4.44
r1024 (  20 35 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=54.39 //y=4.44 //x2=54.39 //y2=4.44
r1025 (  18 33 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=39.22 //y=4.44 //x2=39.22 //y2=4.44
r1026 (  16 31 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=29.97 //y=4.44 //x2=29.97 //y2=4.44
r1027 (  14 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.8 //y=4.44 //x2=14.8 //y2=4.44
r1028 (  12 26 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.55 //y=4.44 //x2=5.55 //y2=4.44
r1029 (  10 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=54.505 //y=4.44 //x2=54.39 //y2=4.44
r1030 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=63.525 //y=4.44 //x2=63.64 //y2=4.44
r1031 (  9 10 ) resistor r=8.60687 //w=0.131 //l=9.02 //layer=m1 \
 //thickness=0.36 //x=63.525 //y=4.44 //x2=54.505 //y2=4.44
r1032 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=39.335 //y=4.44 //x2=39.22 //y2=4.44
r1033 (  7 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=54.275 //y=4.44 //x2=54.39 //y2=4.44
r1034 (  7 8 ) resistor r=14.2557 //w=0.131 //l=14.94 //layer=m1 \
 //thickness=0.36 //x=54.275 //y=4.44 //x2=39.335 //y2=4.44
r1035 (  6 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=30.085 //y=4.44 //x2=29.97 //y2=4.44
r1036 (  5 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=39.105 //y=4.44 //x2=39.22 //y2=4.44
r1037 (  5 6 ) resistor r=8.60687 //w=0.131 //l=9.02 //layer=m1 \
 //thickness=0.36 //x=39.105 //y=4.44 //x2=30.085 //y2=4.44
r1038 (  4 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=14.915 //y=4.44 //x2=14.8 //y2=4.44
r1039 (  3 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=29.855 //y=4.44 //x2=29.97 //y2=4.44
r1040 (  3 4 ) resistor r=14.2557 //w=0.131 //l=14.94 //layer=m1 \
 //thickness=0.36 //x=29.855 //y=4.44 //x2=14.915 //y2=4.44
r1041 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.665 //y=4.44 //x2=5.55 //y2=4.44
r1042 (  1 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=14.685 //y=4.44 //x2=14.8 //y2=4.44
r1043 (  1 2 ) resistor r=8.60687 //w=0.131 //l=9.02 //layer=m1 \
 //thickness=0.36 //x=14.685 //y=4.44 //x2=5.665 //y2=4.44
ends PM_TMRDFFSNQX1\%CLK

subckt PM_TMRDFFSNQX1\%noxref_18 ( 1 2 3 4 11 13 23 24 31 39 45 46 50 52 61 62 \
 64 65 67 68 69 70 71 72 73 74 75 80 82 84 90 91 92 93 94 95 99 101 104 105 \
 110 111 114 128 131 133 134 135 )
c291 ( 135 0 ) capacitor c=0.023087f //x=55.315 //y=5.02
c292 ( 134 0 ) capacitor c=0.023519f //x=54.435 //y=5.02
c293 ( 133 0 ) capacitor c=0.0224735f //x=53.555 //y=5.02
c294 ( 131 0 ) capacitor c=0.00853354f //x=55.565 //y=0.915
c295 ( 128 0 ) capacitor c=0.0597793f //x=66.23 //y=4.7
c296 ( 114 0 ) capacitor c=0.0331095f //x=50.72 //y=4.7
c297 ( 111 0 ) capacitor c=0.0279499f //x=50.69 //y=1.915
c298 ( 110 0 ) capacitor c=0.0421676f //x=50.69 //y=2.08
c299 ( 105 0 ) capacitor c=0.0318948f //x=66.565 //y=1.21
c300 ( 104 0 ) capacitor c=0.0187384f //x=66.565 //y=0.865
c301 ( 101 0 ) capacitor c=0.0141798f //x=66.41 //y=1.365
c302 ( 99 0 ) capacitor c=0.0149844f //x=66.41 //y=0.71
c303 ( 95 0 ) capacitor c=0.0813322f //x=66.035 //y=1.915
c304 ( 94 0 ) capacitor c=0.0229267f //x=66.035 //y=1.52
c305 ( 93 0 ) capacitor c=0.0234352f //x=66.035 //y=1.21
c306 ( 92 0 ) capacitor c=0.0199343f //x=66.035 //y=0.865
c307 ( 91 0 ) capacitor c=0.0429696f //x=51.255 //y=1.25
c308 ( 90 0 ) capacitor c=0.0192208f //x=51.255 //y=0.905
c309 ( 84 0 ) capacitor c=0.0148884f //x=51.1 //y=1.405
c310 ( 82 0 ) capacitor c=0.0157803f //x=51.1 //y=0.75
c311 ( 80 0 ) capacitor c=0.0295235f //x=51.095 //y=4.79
c312 ( 75 0 ) capacitor c=0.0205163f //x=50.725 //y=1.56
c313 ( 74 0 ) capacitor c=0.0168481f //x=50.725 //y=1.25
c314 ( 73 0 ) capacitor c=0.0174783f //x=50.725 //y=0.905
c315 ( 72 0 ) capacitor c=0.110141f //x=66.57 //y=6.02
c316 ( 71 0 ) capacitor c=0.154305f //x=66.13 //y=6.02
c317 ( 70 0 ) capacitor c=0.15358f //x=51.17 //y=6.02
c318 ( 69 0 ) capacitor c=0.110281f //x=50.73 //y=6.02
c319 ( 65 0 ) capacitor c=0.0715637f //x=56.237 //y=3.905
c320 ( 64 0 ) capacitor c=0.0101843f //x=56.235 //y=4.07
c321 ( 62 0 ) capacitor c=0.00106608f //x=55.46 //y=5.155
c322 ( 61 0 ) capacitor c=0.00207162f //x=54.58 //y=5.155
c323 ( 52 0 ) capacitor c=0.0873188f //x=66.23 //y=2.08
c324 ( 50 0 ) capacitor c=0.0236247f //x=56.24 //y=5.07
c325 ( 46 0 ) capacitor c=0.00398962f //x=55.84 //y=1.665
c326 ( 45 0 ) capacitor c=0.0135805f //x=56.155 //y=1.665
c327 ( 39 0 ) capacitor c=0.0281378f //x=56.155 //y=5.155
c328 ( 31 0 ) capacitor c=0.0176454f //x=55.375 //y=5.155
c329 ( 24 0 ) capacitor c=0.00332903f //x=53.785 //y=5.155
c330 ( 23 0 ) capacitor c=0.014837f //x=54.495 //y=5.155
c331 ( 13 0 ) capacitor c=0.0676912f //x=50.69 //y=2.08
c332 ( 11 0 ) capacitor c=0.00453889f //x=50.69 //y=4.535
c333 ( 4 0 ) capacitor c=0.00551102f //x=56.35 //y=4.07
c334 ( 3 0 ) capacitor c=0.180782f //x=66.115 //y=4.07
c335 ( 2 0 ) capacitor c=0.0100678f //x=50.805 //y=4.07
c336 ( 1 0 ) capacitor c=0.0882171f //x=56.12 //y=4.07
r337 (  126 128 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=66.13 //y=4.7 //x2=66.23 //y2=4.7
r338 (  116 117 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=50.72 //y=4.79 //x2=50.72 //y2=4.865
r339 (  114 116 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=50.72 //y=4.7 //x2=50.72 //y2=4.79
r340 (  110 111 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=50.69 //y=2.08 //x2=50.69 //y2=1.915
r341 (  106 128 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=66.57 //y=4.865 //x2=66.23 //y2=4.7
r342 (  105 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.565 //y=1.21 //x2=66.525 //y2=1.365
r343 (  104 129 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.565 //y=0.865 //x2=66.525 //y2=0.71
r344 (  104 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=66.565 //y=0.865 //x2=66.565 //y2=1.21
r345 (  102 125 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.19 //y=1.365 //x2=66.075 //y2=1.365
r346 (  101 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.41 //y=1.365 //x2=66.525 //y2=1.365
r347 (  100 124 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.19 //y=0.71 //x2=66.075 //y2=0.71
r348 (  99 129 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=66.41 //y=0.71 //x2=66.525 //y2=0.71
r349 (  99 100 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=66.41 //y=0.71 //x2=66.19 //y2=0.71
r350 (  96 126 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=66.13 //y=4.865 //x2=66.13 //y2=4.7
r351 (  95 123 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=66.035 //y=1.915 //x2=66.23 //y2=2.08
r352 (  94 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.035 //y=1.52 //x2=66.075 //y2=1.365
r353 (  94 95 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=66.035 //y=1.52 //x2=66.035 //y2=1.915
r354 (  93 125 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.035 //y=1.21 //x2=66.075 //y2=1.365
r355 (  92 124 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=66.035 //y=0.865 //x2=66.075 //y2=0.71
r356 (  92 93 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=66.035 //y=0.865 //x2=66.035 //y2=1.21
r357 (  91 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.255 //y=1.25 //x2=51.215 //y2=1.405
r358 (  90 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=51.255 //y=0.905 //x2=51.215 //y2=0.75
r359 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=51.255 //y=0.905 //x2=51.255 //y2=1.25
r360 (  85 119 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.88 //y=1.405 //x2=50.765 //y2=1.405
r361 (  84 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=51.1 //y=1.405 //x2=51.215 //y2=1.405
r362 (  83 118 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=50.88 //y=0.75 //x2=50.765 //y2=0.75
r363 (  82 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=51.1 //y=0.75 //x2=51.215 //y2=0.75
r364 (  82 83 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=51.1 //y=0.75 //x2=50.88 //y2=0.75
r365 (  81 116 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=50.855 //y=4.79 //x2=50.72 //y2=4.79
r366 (  80 87 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=51.095 //y=4.79 //x2=51.17 //y2=4.865
r367 (  80 81 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=51.095 //y=4.79 //x2=50.855 //y2=4.79
r368 (  75 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.725 //y=1.56 //x2=50.765 //y2=1.405
r369 (  75 111 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=50.725 //y=1.56 //x2=50.725 //y2=1.915
r370 (  74 119 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.725 //y=1.25 //x2=50.765 //y2=1.405
r371 (  73 118 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=50.725 //y=0.905 //x2=50.765 //y2=0.75
r372 (  73 74 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=50.725 //y=0.905 //x2=50.725 //y2=1.25
r373 (  72 106 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=66.57 //y=6.02 //x2=66.57 //y2=4.865
r374 (  71 96 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=66.13 //y=6.02 //x2=66.13 //y2=4.865
r375 (  70 87 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=51.17 //y=6.02 //x2=51.17 //y2=4.865
r376 (  69 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=50.73 //y=6.02 //x2=50.73 //y2=4.865
r377 (  68 101 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=66.3 //y=1.365 //x2=66.41 //y2=1.365
r378 (  68 102 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=66.3 //y=1.365 //x2=66.19 //y2=1.365
r379 (  67 84 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=50.99 //y=1.405 //x2=51.1 //y2=1.405
r380 (  67 85 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=50.99 //y=1.405 //x2=50.88 //y2=1.405
r381 (  64 66 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=56.237 //y=4.07 //x2=56.237 //y2=4.235
r382 (  64 65 ) resistor r=11 //w=0.192 //l=0.165 //layer=li //thickness=0.1 \
 //x=56.237 //y=4.07 //x2=56.237 //y2=3.905
r383 (  60 114 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=50.72 //y=4.7 //x2=50.72 //y2=4.7
r384 (  57 128 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=66.23 //y=4.7 //x2=66.23 //y2=4.7
r385 (  55 57 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=66.23 //y=4.07 //x2=66.23 //y2=4.7
r386 (  52 123 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=66.23 //y=2.08 //x2=66.23 //y2=2.08
r387 (  52 55 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=66.23 //y=2.08 //x2=66.23 //y2=4.07
r388 (  50 66 ) resistor r=57.1551 //w=0.187 //l=0.835 //layer=li \
 //thickness=0.1 //x=56.24 //y=5.07 //x2=56.24 //y2=4.235
r389 (  47 65 ) resistor r=147.508 //w=0.187 //l=2.155 //layer=li \
 //thickness=0.1 //x=56.24 //y=1.75 //x2=56.24 //y2=3.905
r390 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.155 //y=1.665 //x2=56.24 //y2=1.75
r391 (  45 46 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=56.155 //y=1.665 //x2=55.84 //y2=1.665
r392 (  41 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=55.755 //y=1.58 //x2=55.84 //y2=1.665
r393 (  41 131 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=55.755 //y=1.58 //x2=55.755 //y2=1.01
r394 (  40 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.545 //y=5.155 //x2=55.46 //y2=5.155
r395 (  39 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=56.155 //y=5.155 //x2=56.24 //y2=5.07
r396 (  39 40 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=56.155 //y=5.155 //x2=55.545 //y2=5.155
r397 (  33 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.46 //y=5.24 //x2=55.46 //y2=5.155
r398 (  33 135 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=55.46 //y=5.24 //x2=55.46 //y2=5.725
r399 (  32 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.665 //y=5.155 //x2=54.58 //y2=5.155
r400 (  31 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=55.375 //y=5.155 //x2=55.46 //y2=5.155
r401 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=55.375 //y=5.155 //x2=54.665 //y2=5.155
r402 (  25 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.58 //y=5.24 //x2=54.58 //y2=5.155
r403 (  25 134 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=54.58 //y=5.24 //x2=54.58 //y2=5.725
r404 (  23 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.495 //y=5.155 //x2=54.58 //y2=5.155
r405 (  23 24 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=54.495 //y=5.155 //x2=53.785 //y2=5.155
r406 (  17 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=53.7 //y=5.24 //x2=53.785 //y2=5.155
r407 (  17 133 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=53.7 //y=5.24 //x2=53.7 //y2=5.725
r408 (  13 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=50.69 //y=2.08 //x2=50.69 //y2=2.08
r409 (  13 16 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=50.69 //y=2.08 //x2=50.69 //y2=4.07
r410 (  11 60 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=50.69 //y=4.535 //x2=50.705 //y2=4.7
r411 (  11 16 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=50.69 //y=4.535 //x2=50.69 //y2=4.07
r412 (  10 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=66.23 //y=4.07 //x2=66.23 //y2=4.07
r413 (  8 64 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=56.235 //y=4.07 //x2=56.235 //y2=4.07
r414 (  6 16 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=50.69 //y=4.07 //x2=50.69 //y2=4.07
r415 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=56.35 //y=4.07 //x2=56.235 //y2=4.07
r416 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=66.115 //y=4.07 //x2=66.23 //y2=4.07
r417 (  3 4 ) resistor r=9.31775 //w=0.131 //l=9.765 //layer=m1 \
 //thickness=0.36 //x=66.115 //y=4.07 //x2=56.35 //y2=4.07
r418 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=50.805 //y=4.07 //x2=50.69 //y2=4.07
r419 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=56.12 //y=4.07 //x2=56.235 //y2=4.07
r420 (  1 2 ) resistor r=5.07156 //w=0.131 //l=5.315 //layer=m1 \
 //thickness=0.36 //x=56.12 //y=4.07 //x2=50.805 //y2=4.07
ends PM_TMRDFFSNQX1\%noxref_18

subckt PM_TMRDFFSNQX1\%noxref_19 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 \
 47 48 49 51 57 58 59 60 72 74 75 )
c165 ( 75 0 ) capacitor c=0.0220291f //x=67.085 //y=5.02
c166 ( 74 0 ) capacitor c=0.0217503f //x=66.205 //y=5.02
c167 ( 72 0 ) capacitor c=0.0084702f //x=67.08 //y=0.905
c168 ( 60 0 ) capacitor c=0.0546771f //x=69.835 //y=4.79
c169 ( 59 0 ) capacitor c=0.0293157f //x=70.125 //y=4.79
c170 ( 58 0 ) capacitor c=0.0347816f //x=69.79 //y=1.22
c171 ( 57 0 ) capacitor c=0.0187487f //x=69.79 //y=0.875
c172 ( 51 0 ) capacitor c=0.0137055f //x=69.635 //y=1.375
c173 ( 49 0 ) capacitor c=0.0149861f //x=69.635 //y=0.72
c174 ( 48 0 ) capacitor c=0.096037f //x=69.26 //y=1.915
c175 ( 47 0 ) capacitor c=0.0228993f //x=69.26 //y=1.53
c176 ( 46 0 ) capacitor c=0.0234352f //x=69.26 //y=1.22
c177 ( 45 0 ) capacitor c=0.0198724f //x=69.26 //y=0.875
c178 ( 44 0 ) capacitor c=0.110114f //x=70.2 //y=6.02
c179 ( 43 0 ) capacitor c=0.15724f //x=69.76 //y=6.02
c180 ( 41 0 ) capacitor c=0.00211606f //x=67.23 //y=5.2
c181 ( 34 0 ) capacitor c=0.101814f //x=69.56 //y=2.08
c182 ( 32 0 ) capacitor c=0.107182f //x=67.71 //y=4.81
c183 ( 28 0 ) capacitor c=0.00404073f //x=67.355 //y=1.655
c184 ( 27 0 ) capacitor c=0.0122201f //x=67.625 //y=1.655
c185 ( 25 0 ) capacitor c=0.0136983f //x=67.625 //y=5.2
c186 ( 14 0 ) capacitor c=0.00272496f //x=66.435 //y=5.2
c187 ( 13 0 ) capacitor c=0.0151328f //x=67.145 //y=5.2
c188 ( 2 0 ) capacitor c=0.0137738f //x=67.825 //y=4.81
c189 ( 1 0 ) capacitor c=0.0535064f //x=69.445 //y=4.81
r190 (  59 61 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=70.125 //y=4.79 //x2=70.2 //y2=4.865
r191 (  59 60 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=70.125 //y=4.79 //x2=69.835 //y2=4.79
r192 (  58 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.79 //y=1.22 //x2=69.75 //y2=1.375
r193 (  57 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.79 //y=0.875 //x2=69.75 //y2=0.72
r194 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=69.79 //y=0.875 //x2=69.79 //y2=1.22
r195 (  54 60 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=69.76 //y=4.865 //x2=69.835 //y2=4.79
r196 (  54 69 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=69.76 //y=4.865 //x2=69.56 //y2=4.7
r197 (  52 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.415 //y=1.375 //x2=69.3 //y2=1.375
r198 (  51 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.635 //y=1.375 //x2=69.75 //y2=1.375
r199 (  50 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.415 //y=0.72 //x2=69.3 //y2=0.72
r200 (  49 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=69.635 //y=0.72 //x2=69.75 //y2=0.72
r201 (  49 50 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=69.635 //y=0.72 //x2=69.415 //y2=0.72
r202 (  48 67 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=69.26 //y=1.915 //x2=69.56 //y2=2.08
r203 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.26 //y=1.53 //x2=69.3 //y2=1.375
r204 (  47 48 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=69.26 //y=1.53 //x2=69.26 //y2=1.915
r205 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.26 //y=1.22 //x2=69.3 //y2=1.375
r206 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=69.26 //y=0.875 //x2=69.3 //y2=0.72
r207 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=69.26 //y=0.875 //x2=69.26 //y2=1.22
r208 (  44 61 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=70.2 //y=6.02 //x2=70.2 //y2=4.865
r209 (  43 54 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=69.76 //y=6.02 //x2=69.76 //y2=4.865
r210 (  42 51 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=69.525 //y=1.375 //x2=69.635 //y2=1.375
r211 (  42 52 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=69.525 //y=1.375 //x2=69.415 //y2=1.375
r212 (  37 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=69.56 //y=4.7 //x2=69.56 //y2=4.7
r213 (  37 39 ) resistor r=7.52941 //w=0.187 //l=0.11 //layer=li \
 //thickness=0.1 //x=69.56 //y=4.7 //x2=69.56 //y2=4.81
r214 (  34 67 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=69.56 //y=2.08 //x2=69.56 //y2=2.08
r215 (  34 37 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li \
 //thickness=0.1 //x=69.56 //y=2.08 //x2=69.56 //y2=4.7
r216 (  30 32 ) resistor r=20.877 //w=0.187 //l=0.305 //layer=li \
 //thickness=0.1 //x=67.71 //y=5.115 //x2=67.71 //y2=4.81
r217 (  29 32 ) resistor r=210.139 //w=0.187 //l=3.07 //layer=li \
 //thickness=0.1 //x=67.71 //y=1.74 //x2=67.71 //y2=4.81
r218 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=67.625 //y=1.655 //x2=67.71 //y2=1.74
r219 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=67.625 //y=1.655 //x2=67.355 //y2=1.655
r220 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.315 //y=5.2 //x2=67.23 //y2=5.2
r221 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=67.625 //y=5.2 //x2=67.71 //y2=5.115
r222 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=67.625 //y=5.2 //x2=67.315 //y2=5.2
r223 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=67.27 //y=1.57 //x2=67.355 //y2=1.655
r224 (  21 72 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=67.27 //y=1.57 //x2=67.27 //y2=1
r225 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.23 //y=5.285 //x2=67.23 //y2=5.2
r226 (  15 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=67.23 //y=5.285 //x2=67.23 //y2=5.725
r227 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=67.145 //y=5.2 //x2=67.23 //y2=5.2
r228 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=67.145 //y=5.2 //x2=66.435 //y2=5.2
r229 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=66.35 //y=5.285 //x2=66.435 //y2=5.2
r230 (  7 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=66.35 //y=5.285 //x2=66.35 //y2=5.725
r231 (  6 39 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=69.56 //y=4.81 //x2=69.56 //y2=4.81
r232 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=67.71 //y=4.81 //x2=67.71 //y2=4.81
r233 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=67.825 //y=4.81 //x2=67.71 //y2=4.81
r234 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=69.445 //y=4.81 //x2=69.56 //y2=4.81
r235 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=69.445 //y=4.81 //x2=67.825 //y2=4.81
ends PM_TMRDFFSNQX1\%noxref_19

subckt PM_TMRDFFSNQX1\%SN ( 1 2 3 4 5 6 7 8 9 10 23 24 25 26 27 28 29 30 31 32 \
 34 44 54 62 70 79 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 \
 104 105 106 108 114 115 116 117 118 123 124 125 127 133 134 135 136 137 142 \
 143 144 146 152 153 154 155 156 161 162 163 165 171 172 173 174 175 180 181 \
 182 184 190 191 192 193 194 199 200 201 203 209 210 211 212 213 221 232 243 \
 254 265 276 )
c815 ( 276 0 ) capacitor c=0.0335551f //x=70.67 //y=4.7
c816 ( 265 0 ) capacitor c=0.0335551f //x=59.2 //y=4.7
c817 ( 254 0 ) capacitor c=0.0335551f //x=46.25 //y=4.7
c818 ( 243 0 ) capacitor c=0.0335551f //x=34.78 //y=4.7
c819 ( 232 0 ) capacitor c=0.0335551f //x=21.83 //y=4.7
c820 ( 221 0 ) capacitor c=0.0335551f //x=10.36 //y=4.7
c821 ( 213 0 ) capacitor c=0.0245352f //x=71.005 //y=4.79
c822 ( 212 0 ) capacitor c=0.0827272f //x=70.76 //y=1.915
c823 ( 211 0 ) capacitor c=0.0170266f //x=70.76 //y=1.45
c824 ( 210 0 ) capacitor c=0.018609f //x=70.76 //y=1.22
c825 ( 209 0 ) capacitor c=0.0187309f //x=70.76 //y=0.91
c826 ( 203 0 ) capacitor c=0.014725f //x=70.605 //y=1.375
c827 ( 201 0 ) capacitor c=0.0146567f //x=70.605 //y=0.755
c828 ( 200 0 ) capacitor c=0.0335408f //x=70.235 //y=1.22
c829 ( 199 0 ) capacitor c=0.0173761f //x=70.235 //y=0.91
c830 ( 194 0 ) capacitor c=0.0245352f //x=59.535 //y=4.79
c831 ( 193 0 ) capacitor c=0.0825033f //x=59.29 //y=1.915
c832 ( 192 0 ) capacitor c=0.0170266f //x=59.29 //y=1.45
c833 ( 191 0 ) capacitor c=0.018609f //x=59.29 //y=1.22
c834 ( 190 0 ) capacitor c=0.0187309f //x=59.29 //y=0.91
c835 ( 184 0 ) capacitor c=0.014725f //x=59.135 //y=1.375
c836 ( 182 0 ) capacitor c=0.0146567f //x=59.135 //y=0.755
c837 ( 181 0 ) capacitor c=0.0335408f //x=58.765 //y=1.22
c838 ( 180 0 ) capacitor c=0.0173761f //x=58.765 //y=0.91
c839 ( 175 0 ) capacitor c=0.0245352f //x=46.585 //y=4.79
c840 ( 174 0 ) capacitor c=0.0825033f //x=46.34 //y=1.915
c841 ( 173 0 ) capacitor c=0.0170266f //x=46.34 //y=1.45
c842 ( 172 0 ) capacitor c=0.018609f //x=46.34 //y=1.22
c843 ( 171 0 ) capacitor c=0.0187309f //x=46.34 //y=0.91
c844 ( 165 0 ) capacitor c=0.014725f //x=46.185 //y=1.375
c845 ( 163 0 ) capacitor c=0.0146567f //x=46.185 //y=0.755
c846 ( 162 0 ) capacitor c=0.0335408f //x=45.815 //y=1.22
c847 ( 161 0 ) capacitor c=0.0173761f //x=45.815 //y=0.91
c848 ( 156 0 ) capacitor c=0.0245352f //x=35.115 //y=4.79
c849 ( 155 0 ) capacitor c=0.0825033f //x=34.87 //y=1.915
c850 ( 154 0 ) capacitor c=0.0170266f //x=34.87 //y=1.45
c851 ( 153 0 ) capacitor c=0.018609f //x=34.87 //y=1.22
c852 ( 152 0 ) capacitor c=0.0187309f //x=34.87 //y=0.91
c853 ( 146 0 ) capacitor c=0.014725f //x=34.715 //y=1.375
c854 ( 144 0 ) capacitor c=0.0146567f //x=34.715 //y=0.755
c855 ( 143 0 ) capacitor c=0.0335408f //x=34.345 //y=1.22
c856 ( 142 0 ) capacitor c=0.0173761f //x=34.345 //y=0.91
c857 ( 137 0 ) capacitor c=0.0245352f //x=22.165 //y=4.79
c858 ( 136 0 ) capacitor c=0.0825033f //x=21.92 //y=1.915
c859 ( 135 0 ) capacitor c=0.0170266f //x=21.92 //y=1.45
c860 ( 134 0 ) capacitor c=0.018609f //x=21.92 //y=1.22
c861 ( 133 0 ) capacitor c=0.0187309f //x=21.92 //y=0.91
c862 ( 127 0 ) capacitor c=0.014725f //x=21.765 //y=1.375
c863 ( 125 0 ) capacitor c=0.0146567f //x=21.765 //y=0.755
c864 ( 124 0 ) capacitor c=0.0335408f //x=21.395 //y=1.22
c865 ( 123 0 ) capacitor c=0.0173761f //x=21.395 //y=0.91
c866 ( 118 0 ) capacitor c=0.0245352f //x=10.695 //y=4.79
c867 ( 117 0 ) capacitor c=0.0826756f //x=10.45 //y=1.915
c868 ( 116 0 ) capacitor c=0.0170266f //x=10.45 //y=1.45
c869 ( 115 0 ) capacitor c=0.018609f //x=10.45 //y=1.22
c870 ( 114 0 ) capacitor c=0.0187309f //x=10.45 //y=0.91
c871 ( 108 0 ) capacitor c=0.014725f //x=10.295 //y=1.375
c872 ( 106 0 ) capacitor c=0.0146567f //x=10.295 //y=0.755
c873 ( 105 0 ) capacitor c=0.0335408f //x=9.925 //y=1.22
c874 ( 104 0 ) capacitor c=0.0173761f //x=9.925 //y=0.91
c875 ( 103 0 ) capacitor c=0.110114f //x=71.08 //y=6.02
c876 ( 102 0 ) capacitor c=0.109821f //x=70.64 //y=6.02
c877 ( 101 0 ) capacitor c=0.110114f //x=59.61 //y=6.02
c878 ( 100 0 ) capacitor c=0.11012f //x=59.17 //y=6.02
c879 ( 99 0 ) capacitor c=0.110114f //x=46.66 //y=6.02
c880 ( 98 0 ) capacitor c=0.11012f //x=46.22 //y=6.02
c881 ( 97 0 ) capacitor c=0.110114f //x=35.19 //y=6.02
c882 ( 96 0 ) capacitor c=0.11012f //x=34.75 //y=6.02
c883 ( 95 0 ) capacitor c=0.110114f //x=22.24 //y=6.02
c884 ( 94 0 ) capacitor c=0.11012f //x=21.8 //y=6.02
c885 ( 93 0 ) capacitor c=0.110114f //x=10.77 //y=6.02
c886 ( 92 0 ) capacitor c=0.11012f //x=10.33 //y=6.02
c887 ( 79 0 ) capacitor c=0.0933884f //x=70.67 //y=2.08
c888 ( 70 0 ) capacitor c=0.0895052f //x=59.2 //y=2.08
c889 ( 62 0 ) capacitor c=0.0894348f //x=46.25 //y=2.08
c890 ( 54 0 ) capacitor c=0.0895052f //x=34.78 //y=2.08
c891 ( 44 0 ) capacitor c=0.0925216f //x=21.83 //y=2.08
c892 ( 34 0 ) capacitor c=0.0921487f //x=10.36 //y=2.08
c893 ( 10 0 ) capacitor c=0.00692137f //x=59.315 //y=2.22
c894 ( 9 0 ) capacitor c=0.263609f //x=70.555 //y=2.22
c895 ( 8 0 ) capacitor c=0.00692137f //x=46.365 //y=2.22
c896 ( 7 0 ) capacitor c=0.257357f //x=59.085 //y=2.22
c897 ( 6 0 ) capacitor c=0.00692137f //x=34.895 //y=2.22
c898 ( 5 0 ) capacitor c=0.240835f //x=46.135 //y=2.22
c899 ( 4 0 ) capacitor c=0.00692137f //x=21.945 //y=2.22
c900 ( 3 0 ) capacitor c=0.266406f //x=34.665 //y=2.22
c901 ( 2 0 ) capacitor c=0.0154797f //x=10.475 //y=2.22
c902 ( 1 0 ) capacitor c=0.248273f //x=21.715 //y=2.22
r903 (  278 279 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=70.67 //y=4.79 //x2=70.67 //y2=4.865
r904 (  276 278 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=70.67 //y=4.7 //x2=70.67 //y2=4.79
r905 (  267 268 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=59.2 //y=4.79 //x2=59.2 //y2=4.865
r906 (  265 267 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=59.2 //y=4.7 //x2=59.2 //y2=4.79
r907 (  256 257 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=46.25 //y=4.79 //x2=46.25 //y2=4.865
r908 (  254 256 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=46.25 //y=4.7 //x2=46.25 //y2=4.79
r909 (  245 246 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=34.78 //y=4.79 //x2=34.78 //y2=4.865
r910 (  243 245 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=34.78 //y=4.7 //x2=34.78 //y2=4.79
r911 (  234 235 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=21.83 //y=4.79 //x2=21.83 //y2=4.865
r912 (  232 234 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=21.83 //y=4.7 //x2=21.83 //y2=4.79
r913 (  223 224 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=10.36 //y=4.79 //x2=10.36 //y2=4.865
r914 (  221 223 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=10.36 //y=4.7 //x2=10.36 //y2=4.79
r915 (  214 278 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=70.805 //y=4.79 //x2=70.67 //y2=4.79
r916 (  213 215 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=71.005 //y=4.79 //x2=71.08 //y2=4.865
r917 (  213 214 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=71.005 //y=4.79 //x2=70.805 //y2=4.79
r918 (  212 283 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=70.76 //y=1.915 //x2=70.685 //y2=2.08
r919 (  211 281 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=70.76 //y=1.45 //x2=70.72 //y2=1.375
r920 (  211 212 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=70.76 //y=1.45 //x2=70.76 //y2=1.915
r921 (  210 281 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.76 //y=1.22 //x2=70.72 //y2=1.375
r922 (  209 280 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.76 //y=0.91 //x2=70.72 //y2=0.755
r923 (  209 210 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=70.76 //y=0.91 //x2=70.76 //y2=1.22
r924 (  204 274 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.39 //y=1.375 //x2=70.275 //y2=1.375
r925 (  203 281 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.605 //y=1.375 //x2=70.72 //y2=1.375
r926 (  202 273 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.39 //y=0.755 //x2=70.275 //y2=0.755
r927 (  201 280 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=70.605 //y=0.755 //x2=70.72 //y2=0.755
r928 (  201 202 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=70.605 //y=0.755 //x2=70.39 //y2=0.755
r929 (  200 274 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.235 //y=1.22 //x2=70.275 //y2=1.375
r930 (  199 273 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=70.235 //y=0.91 //x2=70.275 //y2=0.755
r931 (  199 200 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=70.235 //y=0.91 //x2=70.235 //y2=1.22
r932 (  195 267 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=59.335 //y=4.79 //x2=59.2 //y2=4.79
r933 (  194 196 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=59.535 //y=4.79 //x2=59.61 //y2=4.865
r934 (  194 195 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=59.535 //y=4.79 //x2=59.335 //y2=4.79
r935 (  193 272 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=59.29 //y=1.915 //x2=59.215 //y2=2.08
r936 (  192 270 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=59.29 //y=1.45 //x2=59.25 //y2=1.375
r937 (  192 193 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=59.29 //y=1.45 //x2=59.29 //y2=1.915
r938 (  191 270 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.29 //y=1.22 //x2=59.25 //y2=1.375
r939 (  190 269 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=59.29 //y=0.91 //x2=59.25 //y2=0.755
r940 (  190 191 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=59.29 //y=0.91 //x2=59.29 //y2=1.22
r941 (  185 263 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.92 //y=1.375 //x2=58.805 //y2=1.375
r942 (  184 270 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.135 //y=1.375 //x2=59.25 //y2=1.375
r943 (  183 262 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=58.92 //y=0.755 //x2=58.805 //y2=0.755
r944 (  182 269 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=59.135 //y=0.755 //x2=59.25 //y2=0.755
r945 (  182 183 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=59.135 //y=0.755 //x2=58.92 //y2=0.755
r946 (  181 263 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.765 //y=1.22 //x2=58.805 //y2=1.375
r947 (  180 262 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=58.765 //y=0.91 //x2=58.805 //y2=0.755
r948 (  180 181 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=58.765 //y=0.91 //x2=58.765 //y2=1.22
r949 (  176 256 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=46.385 //y=4.79 //x2=46.25 //y2=4.79
r950 (  175 177 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=46.585 //y=4.79 //x2=46.66 //y2=4.865
r951 (  175 176 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=46.585 //y=4.79 //x2=46.385 //y2=4.79
r952 (  174 261 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=46.34 //y=1.915 //x2=46.265 //y2=2.08
r953 (  173 259 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=46.34 //y=1.45 //x2=46.3 //y2=1.375
r954 (  173 174 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=46.34 //y=1.45 //x2=46.34 //y2=1.915
r955 (  172 259 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.34 //y=1.22 //x2=46.3 //y2=1.375
r956 (  171 258 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=46.34 //y=0.91 //x2=46.3 //y2=0.755
r957 (  171 172 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=46.34 //y=0.91 //x2=46.34 //y2=1.22
r958 (  166 252 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.97 //y=1.375 //x2=45.855 //y2=1.375
r959 (  165 259 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.185 //y=1.375 //x2=46.3 //y2=1.375
r960 (  164 251 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=45.97 //y=0.755 //x2=45.855 //y2=0.755
r961 (  163 258 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=46.185 //y=0.755 //x2=46.3 //y2=0.755
r962 (  163 164 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=46.185 //y=0.755 //x2=45.97 //y2=0.755
r963 (  162 252 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.815 //y=1.22 //x2=45.855 //y2=1.375
r964 (  161 251 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=45.815 //y=0.91 //x2=45.855 //y2=0.755
r965 (  161 162 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=45.815 //y=0.91 //x2=45.815 //y2=1.22
r966 (  157 245 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=34.915 //y=4.79 //x2=34.78 //y2=4.79
r967 (  156 158 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=35.115 //y=4.79 //x2=35.19 //y2=4.865
r968 (  156 157 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=35.115 //y=4.79 //x2=34.915 //y2=4.79
r969 (  155 250 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=34.87 //y=1.915 //x2=34.795 //y2=2.08
r970 (  154 248 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=34.87 //y=1.45 //x2=34.83 //y2=1.375
r971 (  154 155 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=34.87 //y=1.45 //x2=34.87 //y2=1.915
r972 (  153 248 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.87 //y=1.22 //x2=34.83 //y2=1.375
r973 (  152 247 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.87 //y=0.91 //x2=34.83 //y2=0.755
r974 (  152 153 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=34.87 //y=0.91 //x2=34.87 //y2=1.22
r975 (  147 241 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.5 //y=1.375 //x2=34.385 //y2=1.375
r976 (  146 248 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.715 //y=1.375 //x2=34.83 //y2=1.375
r977 (  145 240 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.5 //y=0.755 //x2=34.385 //y2=0.755
r978 (  144 247 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=34.715 //y=0.755 //x2=34.83 //y2=0.755
r979 (  144 145 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=34.715 //y=0.755 //x2=34.5 //y2=0.755
r980 (  143 241 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.345 //y=1.22 //x2=34.385 //y2=1.375
r981 (  142 240 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=34.345 //y=0.91 //x2=34.385 //y2=0.755
r982 (  142 143 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=34.345 //y=0.91 //x2=34.345 //y2=1.22
r983 (  138 234 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=21.965 //y=4.79 //x2=21.83 //y2=4.79
r984 (  137 139 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=22.165 //y=4.79 //x2=22.24 //y2=4.865
r985 (  137 138 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=22.165 //y=4.79 //x2=21.965 //y2=4.79
r986 (  136 239 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.915 //x2=21.845 //y2=2.08
r987 (  135 237 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.45 //x2=21.88 //y2=1.375
r988 (  135 136 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.45 //x2=21.92 //y2=1.915
r989 (  134 237 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.92 //y=1.22 //x2=21.88 //y2=1.375
r990 (  133 236 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.92 //y=0.91 //x2=21.88 //y2=0.755
r991 (  133 134 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.92 //y=0.91 //x2=21.92 //y2=1.22
r992 (  128 230 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.55 //y=1.375 //x2=21.435 //y2=1.375
r993 (  127 237 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.765 //y=1.375 //x2=21.88 //y2=1.375
r994 (  126 229 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.55 //y=0.755 //x2=21.435 //y2=0.755
r995 (  125 236 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.765 //y=0.755 //x2=21.88 //y2=0.755
r996 (  125 126 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=21.765 //y=0.755 //x2=21.55 //y2=0.755
r997 (  124 230 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.395 //y=1.22 //x2=21.435 //y2=1.375
r998 (  123 229 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.91 //x2=21.435 //y2=0.755
r999 (  123 124 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=21.395 //y=0.91 //x2=21.395 //y2=1.22
r1000 (  119 223 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=10.495 //y=4.79 //x2=10.36 //y2=4.79
r1001 (  118 120 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=10.695 //y=4.79 //x2=10.77 //y2=4.865
r1002 (  118 119 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=10.695 //y=4.79 //x2=10.495 //y2=4.79
r1003 (  117 228 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.915 //x2=10.375 //y2=2.08
r1004 (  116 226 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.45 //x2=10.41 //y2=1.375
r1005 (  116 117 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.45 //x2=10.45 //y2=1.915
r1006 (  115 226 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.45 //y=1.22 //x2=10.41 //y2=1.375
r1007 (  114 225 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.45 //y=0.91 //x2=10.41 //y2=0.755
r1008 (  114 115 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=10.45 //y=0.91 //x2=10.45 //y2=1.22
r1009 (  109 219 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.08 //y=1.375 //x2=9.965 //y2=1.375
r1010 (  108 226 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.295 //y=1.375 //x2=10.41 //y2=1.375
r1011 (  107 218 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.08 //y=0.755 //x2=9.965 //y2=0.755
r1012 (  106 225 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.295 //y=0.755 //x2=10.41 //y2=0.755
r1013 (  106 107 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=10.295 //y=0.755 //x2=10.08 //y2=0.755
r1014 (  105 219 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.925 //y=1.22 //x2=9.965 //y2=1.375
r1015 (  104 218 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=9.925 //y=0.91 //x2=9.965 //y2=0.755
r1016 (  104 105 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=9.925 //y=0.91 //x2=9.925 //y2=1.22
r1017 (  103 215 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=71.08 //y=6.02 //x2=71.08 //y2=4.865
r1018 (  102 279 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=70.64 //y=6.02 //x2=70.64 //y2=4.865
r1019 (  101 196 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.61 //y=6.02 //x2=59.61 //y2=4.865
r1020 (  100 268 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=59.17 //y=6.02 //x2=59.17 //y2=4.865
r1021 (  99 177 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=46.66 //y=6.02 //x2=46.66 //y2=4.865
r1022 (  98 257 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=46.22 //y=6.02 //x2=46.22 //y2=4.865
r1023 (  97 158 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=35.19 //y=6.02 //x2=35.19 //y2=4.865
r1024 (  96 246 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=34.75 //y=6.02 //x2=34.75 //y2=4.865
r1025 (  95 139 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=22.24 //y=6.02 //x2=22.24 //y2=4.865
r1026 (  94 235 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.8 //y=6.02 //x2=21.8 //y2=4.865
r1027 (  93 120 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.77 //y=6.02 //x2=10.77 //y2=4.865
r1028 (  92 224 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.33 //y=6.02 //x2=10.33 //y2=4.865
r1029 (  91 203 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=70.497 //y=1.375 //x2=70.605 //y2=1.375
r1030 (  91 204 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=70.497 //y=1.375 //x2=70.39 //y2=1.375
r1031 (  90 184 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=59.027 //y=1.375 //x2=59.135 //y2=1.375
r1032 (  90 185 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=59.027 //y=1.375 //x2=58.92 //y2=1.375
r1033 (  89 165 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=46.077 //y=1.375 //x2=46.185 //y2=1.375
r1034 (  89 166 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=46.077 //y=1.375 //x2=45.97 //y2=1.375
r1035 (  88 146 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=34.607 //y=1.375 //x2=34.715 //y2=1.375
r1036 (  88 147 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=34.607 //y=1.375 //x2=34.5 //y2=1.375
r1037 (  87 127 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=21.657 //y=1.375 //x2=21.765 //y2=1.375
r1038 (  87 128 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=21.657 //y=1.375 //x2=21.55 //y2=1.375
r1039 (  86 108 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=10.187 //y=1.375 //x2=10.295 //y2=1.375
r1040 (  86 109 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=10.187 //y=1.375 //x2=10.08 //y2=1.375
r1041 (  84 276 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=70.67 //y=4.7 //x2=70.67 //y2=4.7
r1042 (  79 283 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=70.67 //y=2.08 //x2=70.67 //y2=2.08
r1043 (  76 265 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=59.2 //y=4.7 //x2=59.2 //y2=4.7
r1044 (  70 272 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=59.2 //y=2.08 //x2=59.2 //y2=2.08
r1045 (  67 254 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=46.25 //y=4.7 //x2=46.25 //y2=4.7
r1046 (  65 67 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=46.25 //y=2.22 //x2=46.25 //y2=4.7
r1047 (  62 261 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=46.25 //y=2.08 //x2=46.25 //y2=2.08
r1048 (  62 65 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=46.25 //y=2.08 //x2=46.25 //y2=2.22
r1049 (  59 243 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.78 //y=4.7 //x2=34.78 //y2=4.7
r1050 (  54 250 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=34.78 //y=2.08 //x2=34.78 //y2=2.08
r1051 (  51 232 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.83 //y=4.7 //x2=21.83 //y2=4.7
r1052 (  44 239 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.83 //y=2.08 //x2=21.83 //y2=2.08
r1053 (  41 221 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.36 //y=4.7 //x2=10.36 //y2=4.7
r1054 (  34 228 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.36 //y=2.08 //x2=10.36 //y2=2.08
r1055 (  32 84 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=70.67 //y=2.22 //x2=70.67 //y2=4.7
r1056 (  32 79 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=70.67 //y=2.22 //x2=70.67 //y2=2.08
r1057 (  31 76 ) resistor r=144.428 //w=0.187 //l=2.11 //layer=li \
 //thickness=0.1 //x=59.2 //y=2.59 //x2=59.2 //y2=4.7
r1058 (  30 31 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=59.2 //y=2.22 //x2=59.2 //y2=2.59
r1059 (  30 70 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=59.2 //y=2.22 //x2=59.2 //y2=2.08
r1060 (  29 59 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=34.78 //y=2.22 //x2=34.78 //y2=4.7
r1061 (  29 54 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=34.78 //y=2.22 //x2=34.78 //y2=2.08
r1062 (  28 51 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=21.83 //y=4.07 //x2=21.83 //y2=4.7
r1063 (  27 28 ) resistor r=101.305 //w=0.187 //l=1.48 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.59 //x2=21.83 //y2=4.07
r1064 (  26 27 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.22 //x2=21.83 //y2=2.59
r1065 (  26 44 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.22 //x2=21.83 //y2=2.08
r1066 (  25 41 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=10.36 //y=3.33 //x2=10.36 //y2=4.7
r1067 (  24 25 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.59 //x2=10.36 //y2=3.33
r1068 (  23 24 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.22 //x2=10.36 //y2=2.59
r1069 (  23 34 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=10.36 //y=2.22 //x2=10.36 //y2=2.08
r1070 (  22 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=70.67 //y=2.22 //x2=70.67 //y2=2.22
r1071 (  20 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=59.2 //y=2.22 //x2=59.2 //y2=2.22
r1072 (  18 65 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=46.25 //y=2.22 //x2=46.25 //y2=2.22
r1073 (  16 29 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=34.78 //y=2.22 //x2=34.78 //y2=2.22
r1074 (  14 26 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.83 //y=2.22 //x2=21.83 //y2=2.22
r1075 (  12 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.36 //y=2.22 //x2=10.36 //y2=2.22
r1076 (  10 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=59.315 //y=2.22 //x2=59.2 //y2=2.22
r1077 (  9 22 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=70.555 //y=2.22 //x2=70.67 //y2=2.22
r1078 (  9 10 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=70.555 //y=2.22 //x2=59.315 //y2=2.22
r1079 (  8 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=46.365 //y=2.22 //x2=46.25 //y2=2.22
r1080 (  7 20 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=59.085 //y=2.22 //x2=59.2 //y2=2.22
r1081 (  7 8 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=59.085 //y=2.22 //x2=46.365 //y2=2.22
r1082 (  6 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.895 //y=2.22 //x2=34.78 //y2=2.22
r1083 (  5 18 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=46.135 //y=2.22 //x2=46.25 //y2=2.22
r1084 (  5 6 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=46.135 //y=2.22 //x2=34.895 //y2=2.22
r1085 (  4 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.945 //y=2.22 //x2=21.83 //y2=2.22
r1086 (  3 16 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=34.665 //y=2.22 //x2=34.78 //y2=2.22
r1087 (  3 4 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=34.665 //y=2.22 //x2=21.945 //y2=2.22
r1088 (  2 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.475 //y=2.22 //x2=10.36 //y2=2.22
r1089 (  1 14 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.715 //y=2.22 //x2=21.83 //y2=2.22
r1090 (  1 2 ) resistor r=10.7252 //w=0.131 //l=11.24 //layer=m1 \
 //thickness=0.36 //x=21.715 //y=2.22 //x2=10.475 //y2=2.22
ends PM_TMRDFFSNQX1\%SN

subckt PM_TMRDFFSNQX1\%noxref_21 ( 1 2 3 4 5 6 16 24 37 38 49 51 52 56 58 65 \
 66 67 68 69 70 71 72 73 74 78 79 80 85 87 90 91 95 96 97 102 104 107 108 112 \
 113 114 119 121 124 125 127 128 133 137 138 143 147 148 153 156 158 159 )
c321 ( 159 0 ) capacitor c=0.0220291f //x=63.755 //y=5.02
c322 ( 158 0 ) capacitor c=0.0217503f //x=62.875 //y=5.02
c323 ( 156 0 ) capacitor c=0.00866655f //x=63.75 //y=0.905
c324 ( 153 0 ) capacitor c=0.0587755f //x=71.78 //y=4.7
c325 ( 148 0 ) capacitor c=0.0273931f //x=71.78 //y=1.915
c326 ( 147 0 ) capacitor c=0.0458323f //x=71.78 //y=2.08
c327 ( 143 0 ) capacitor c=0.0587755f //x=60.31 //y=4.7
c328 ( 138 0 ) capacitor c=0.0273931f //x=60.31 //y=1.915
c329 ( 137 0 ) capacitor c=0.0456313f //x=60.31 //y=2.08
c330 ( 133 0 ) capacitor c=0.058931f //x=55.5 //y=4.7
c331 ( 128 0 ) capacitor c=0.0267105f //x=55.5 //y=1.915
c332 ( 127 0 ) capacitor c=0.0456313f //x=55.5 //y=2.08
c333 ( 125 0 ) capacitor c=0.0432517f //x=72.3 //y=1.26
c334 ( 124 0 ) capacitor c=0.0200379f //x=72.3 //y=0.915
c335 ( 121 0 ) capacitor c=0.0158629f //x=72.145 //y=1.415
c336 ( 119 0 ) capacitor c=0.0157803f //x=72.145 //y=0.76
c337 ( 114 0 ) capacitor c=0.0218028f //x=71.77 //y=1.57
c338 ( 113 0 ) capacitor c=0.0207459f //x=71.77 //y=1.26
c339 ( 112 0 ) capacitor c=0.0194308f //x=71.77 //y=0.915
c340 ( 108 0 ) capacitor c=0.0432517f //x=60.83 //y=1.26
c341 ( 107 0 ) capacitor c=0.0200379f //x=60.83 //y=0.915
c342 ( 104 0 ) capacitor c=0.0148873f //x=60.675 //y=1.415
c343 ( 102 0 ) capacitor c=0.0157803f //x=60.675 //y=0.76
c344 ( 97 0 ) capacitor c=0.0218028f //x=60.3 //y=1.57
c345 ( 96 0 ) capacitor c=0.0207459f //x=60.3 //y=1.26
c346 ( 95 0 ) capacitor c=0.0194308f //x=60.3 //y=0.915
c347 ( 91 0 ) capacitor c=0.0432517f //x=56.02 //y=1.26
c348 ( 90 0 ) capacitor c=0.0200379f //x=56.02 //y=0.915
c349 ( 87 0 ) capacitor c=0.0148873f //x=55.865 //y=1.415
c350 ( 85 0 ) capacitor c=0.0157803f //x=55.865 //y=0.76
c351 ( 80 0 ) capacitor c=0.0218028f //x=55.49 //y=1.57
c352 ( 79 0 ) capacitor c=0.0207459f //x=55.49 //y=1.26
c353 ( 78 0 ) capacitor c=0.0194308f //x=55.49 //y=0.915
c354 ( 74 0 ) capacitor c=0.158794f //x=71.96 //y=6.02
c355 ( 73 0 ) capacitor c=0.110114f //x=71.52 //y=6.02
c356 ( 72 0 ) capacitor c=0.158794f //x=60.49 //y=6.02
c357 ( 71 0 ) capacitor c=0.110114f //x=60.05 //y=6.02
c358 ( 70 0 ) capacitor c=0.158048f //x=55.68 //y=6.02
c359 ( 69 0 ) capacitor c=0.110114f //x=55.24 //y=6.02
c360 ( 65 0 ) capacitor c=0.0023043f //x=63.9 //y=5.2
c361 ( 58 0 ) capacitor c=0.08651f //x=71.78 //y=2.08
c362 ( 56 0 ) capacitor c=0.104743f //x=64.38 //y=3.7
c363 ( 52 0 ) capacitor c=0.00404073f //x=64.025 //y=1.655
c364 ( 51 0 ) capacitor c=0.0122201f //x=64.295 //y=1.655
c365 ( 49 0 ) capacitor c=0.0140462f //x=64.295 //y=5.2
c366 ( 38 0 ) capacitor c=0.00251635f //x=63.105 //y=5.2
c367 ( 37 0 ) capacitor c=0.0143111f //x=63.815 //y=5.2
c368 ( 24 0 ) capacitor c=0.0811636f //x=60.31 //y=2.08
c369 ( 16 0 ) capacitor c=0.0796434f //x=55.5 //y=2.08
c370 ( 6 0 ) capacitor c=0.00405261f //x=64.495 //y=3.7
c371 ( 5 0 ) capacitor c=0.139723f //x=71.665 //y=3.7
c372 ( 4 0 ) capacitor c=0.00412452f //x=60.425 //y=3.7
c373 ( 3 0 ) capacitor c=0.0546427f //x=64.265 //y=3.7
c374 ( 2 0 ) capacitor c=0.0138772f //x=55.615 //y=3.7
c375 ( 1 0 ) capacitor c=0.0670382f //x=60.195 //y=3.7
r376 (  147 148 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=71.78 //y=2.08 //x2=71.78 //y2=1.915
r377 (  137 138 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=60.31 //y=2.08 //x2=60.31 //y2=1.915
r378 (  127 128 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=55.5 //y=2.08 //x2=55.5 //y2=1.915
r379 (  125 155 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.3 //y=1.26 //x2=72.26 //y2=1.415
r380 (  124 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=72.3 //y=0.915 //x2=72.26 //y2=0.76
r381 (  124 125 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=72.3 //y=0.915 //x2=72.3 //y2=1.26
r382 (  122 151 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=71.925 //y=1.415 //x2=71.81 //y2=1.415
r383 (  121 155 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=72.145 //y=1.415 //x2=72.26 //y2=1.415
r384 (  120 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=71.925 //y=0.76 //x2=71.81 //y2=0.76
r385 (  119 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=72.145 //y=0.76 //x2=72.26 //y2=0.76
r386 (  119 120 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=72.145 //y=0.76 //x2=71.925 //y2=0.76
r387 (  116 153 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=71.96 //y=4.865 //x2=71.78 //y2=4.7
r388 (  114 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.77 //y=1.57 //x2=71.81 //y2=1.415
r389 (  114 148 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=71.77 //y=1.57 //x2=71.77 //y2=1.915
r390 (  113 151 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.77 //y=1.26 //x2=71.81 //y2=1.415
r391 (  112 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=71.77 //y=0.915 //x2=71.81 //y2=0.76
r392 (  112 113 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=71.77 //y=0.915 //x2=71.77 //y2=1.26
r393 (  109 153 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=71.52 //y=4.865 //x2=71.78 //y2=4.7
r394 (  108 145 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.83 //y=1.26 //x2=60.79 //y2=1.415
r395 (  107 144 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.83 //y=0.915 //x2=60.79 //y2=0.76
r396 (  107 108 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=60.83 //y=0.915 //x2=60.83 //y2=1.26
r397 (  105 141 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=60.455 //y=1.415 //x2=60.34 //y2=1.415
r398 (  104 145 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=60.675 //y=1.415 //x2=60.79 //y2=1.415
r399 (  103 140 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=60.455 //y=0.76 //x2=60.34 //y2=0.76
r400 (  102 144 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=60.675 //y=0.76 //x2=60.79 //y2=0.76
r401 (  102 103 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=60.675 //y=0.76 //x2=60.455 //y2=0.76
r402 (  99 143 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=60.49 //y=4.865 //x2=60.31 //y2=4.7
r403 (  97 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.3 //y=1.57 //x2=60.34 //y2=1.415
r404 (  97 138 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=60.3 //y=1.57 //x2=60.3 //y2=1.915
r405 (  96 141 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.3 //y=1.26 //x2=60.34 //y2=1.415
r406 (  95 140 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=60.3 //y=0.915 //x2=60.34 //y2=0.76
r407 (  95 96 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=60.3 //y=0.915 //x2=60.3 //y2=1.26
r408 (  92 143 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=60.05 //y=4.865 //x2=60.31 //y2=4.7
r409 (  91 135 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.02 //y=1.26 //x2=55.98 //y2=1.415
r410 (  90 134 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=56.02 //y=0.915 //x2=55.98 //y2=0.76
r411 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=56.02 //y=0.915 //x2=56.02 //y2=1.26
r412 (  88 131 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.645 //y=1.415 //x2=55.53 //y2=1.415
r413 (  87 135 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.865 //y=1.415 //x2=55.98 //y2=1.415
r414 (  86 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.645 //y=0.76 //x2=55.53 //y2=0.76
r415 (  85 134 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=55.865 //y=0.76 //x2=55.98 //y2=0.76
r416 (  85 86 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=55.865 //y=0.76 //x2=55.645 //y2=0.76
r417 (  82 133 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=55.68 //y=4.865 //x2=55.5 //y2=4.7
r418 (  80 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.49 //y=1.57 //x2=55.53 //y2=1.415
r419 (  80 128 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=55.49 //y=1.57 //x2=55.49 //y2=1.915
r420 (  79 131 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.49 //y=1.26 //x2=55.53 //y2=1.415
r421 (  78 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=55.49 //y=0.915 //x2=55.53 //y2=0.76
r422 (  78 79 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=55.49 //y=0.915 //x2=55.49 //y2=1.26
r423 (  75 133 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=55.24 //y=4.865 //x2=55.5 //y2=4.7
r424 (  74 116 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=71.96 //y=6.02 //x2=71.96 //y2=4.865
r425 (  73 109 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=71.52 //y=6.02 //x2=71.52 //y2=4.865
r426 (  72 99 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=60.49 //y=6.02 //x2=60.49 //y2=4.865
r427 (  71 92 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=60.05 //y=6.02 //x2=60.05 //y2=4.865
r428 (  70 82 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.68 //y=6.02 //x2=55.68 //y2=4.865
r429 (  69 75 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=55.24 //y=6.02 //x2=55.24 //y2=4.865
r430 (  68 121 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=72.035 //y=1.415 //x2=72.145 //y2=1.415
r431 (  68 122 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=72.035 //y=1.415 //x2=71.925 //y2=1.415
r432 (  67 104 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=60.565 //y=1.415 //x2=60.675 //y2=1.415
r433 (  67 105 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=60.565 //y=1.415 //x2=60.455 //y2=1.415
r434 (  66 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=55.755 //y=1.415 //x2=55.865 //y2=1.415
r435 (  66 88 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=55.755 //y=1.415 //x2=55.645 //y2=1.415
r436 (  63 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=71.78 //y=4.7 //x2=71.78 //y2=4.7
r437 (  61 63 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=71.78 //y=3.7 //x2=71.78 //y2=4.7
r438 (  58 147 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=71.78 //y=2.08 //x2=71.78 //y2=2.08
r439 (  58 61 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=71.78 //y=2.08 //x2=71.78 //y2=3.7
r440 (  54 56 ) resistor r=96.8556 //w=0.187 //l=1.415 //layer=li \
 //thickness=0.1 //x=64.38 //y=5.115 //x2=64.38 //y2=3.7
r441 (  53 56 ) resistor r=134.16 //w=0.187 //l=1.96 //layer=li \
 //thickness=0.1 //x=64.38 //y=1.74 //x2=64.38 //y2=3.7
r442 (  51 53 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=64.295 //y=1.655 //x2=64.38 //y2=1.74
r443 (  51 52 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=64.295 //y=1.655 //x2=64.025 //y2=1.655
r444 (  50 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.985 //y=5.2 //x2=63.9 //y2=5.2
r445 (  49 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=64.295 //y=5.2 //x2=64.38 //y2=5.115
r446 (  49 50 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=64.295 //y=5.2 //x2=63.985 //y2=5.2
r447 (  45 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=63.94 //y=1.57 //x2=64.025 //y2=1.655
r448 (  45 156 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=63.94 //y=1.57 //x2=63.94 //y2=1
r449 (  39 65 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.9 //y=5.285 //x2=63.9 //y2=5.2
r450 (  39 159 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=63.9 //y=5.285 //x2=63.9 //y2=5.725
r451 (  37 65 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=63.815 //y=5.2 //x2=63.9 //y2=5.2
r452 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=63.815 //y=5.2 //x2=63.105 //y2=5.2
r453 (  31 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=63.02 //y=5.285 //x2=63.105 //y2=5.2
r454 (  31 158 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=63.02 //y=5.285 //x2=63.02 //y2=5.725
r455 (  29 143 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=60.31 //y=4.7 //x2=60.31 //y2=4.7
r456 (  27 29 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=60.31 //y=3.7 //x2=60.31 //y2=4.7
r457 (  24 137 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=60.31 //y=2.08 //x2=60.31 //y2=2.08
r458 (  24 27 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=60.31 //y=2.08 //x2=60.31 //y2=3.7
r459 (  21 133 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=55.5 //y=4.7 //x2=55.5 //y2=4.7
r460 (  19 21 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=55.5 //y=3.7 //x2=55.5 //y2=4.7
r461 (  16 127 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=55.5 //y=2.08 //x2=55.5 //y2=2.08
r462 (  16 19 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=55.5 //y=2.08 //x2=55.5 //y2=3.7
r463 (  14 61 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=71.78 //y=3.7 //x2=71.78 //y2=3.7
r464 (  12 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=64.38 //y=3.7 //x2=64.38 //y2=3.7
r465 (  10 27 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=60.31 //y=3.7 //x2=60.31 //y2=3.7
r466 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=55.5 //y=3.7 //x2=55.5 //y2=3.7
r467 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=64.495 //y=3.7 //x2=64.38 //y2=3.7
r468 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=71.665 //y=3.7 //x2=71.78 //y2=3.7
r469 (  5 6 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=71.665 //y=3.7 //x2=64.495 //y2=3.7
r470 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=60.425 //y=3.7 //x2=60.31 //y2=3.7
r471 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=64.265 //y=3.7 //x2=64.38 //y2=3.7
r472 (  3 4 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=64.265 //y=3.7 //x2=60.425 //y2=3.7
r473 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=55.615 //y=3.7 //x2=55.5 //y2=3.7
r474 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=60.195 //y=3.7 //x2=60.31 //y2=3.7
r475 (  1 2 ) resistor r=4.37023 //w=0.131 //l=4.58 //layer=m1 \
 //thickness=0.36 //x=60.195 //y=3.7 //x2=55.615 //y2=3.7
ends PM_TMRDFFSNQX1\%noxref_21

subckt PM_TMRDFFSNQX1\%noxref_22 ( 1 2 13 14 15 23 29 30 37 50 51 52 53 54 )
c91 ( 54 0 ) capacitor c=0.034295f //x=78.985 //y=5.025
c92 ( 53 0 ) capacitor c=0.0174957f //x=78.105 //y=5.025
c93 ( 51 0 ) capacitor c=0.0214849f //x=75.225 //y=5.025
c94 ( 50 0 ) capacitor c=0.0217161f //x=74.345 //y=5.025
c95 ( 49 0 ) capacitor c=0.00115294f //x=78.25 //y=6.91
c96 ( 37 0 ) capacitor c=0.0131238f //x=79.045 //y=6.91
c97 ( 30 0 ) capacitor c=0.00386507f //x=77.455 //y=6.91
c98 ( 29 0 ) capacitor c=0.00951687f //x=78.165 //y=6.91
c99 ( 23 0 ) capacitor c=0.0455351f //x=77.37 //y=5.21
c100 ( 15 0 ) capacitor c=0.00871244f //x=75.37 //y=5.295
c101 ( 14 0 ) capacitor c=0.00290434f //x=74.575 //y=5.21
c102 ( 13 0 ) capacitor c=0.0139202f //x=75.285 //y=5.21
c103 ( 2 0 ) capacitor c=0.0091252f //x=75.485 //y=5.21
c104 ( 1 0 ) capacitor c=0.0484159f //x=77.255 //y=5.21
r105 (  39 54 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=79.13 //y=6.825 //x2=79.13 //y2=6.74
r106 (  38 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.335 //y=6.91 //x2=78.25 //y2=6.91
r107 (  37 39 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=79.045 //y=6.91 //x2=79.13 //y2=6.825
r108 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=79.045 //y=6.91 //x2=78.335 //y2=6.91
r109 (  31 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.25 //y=6.825 //x2=78.25 //y2=6.91
r110 (  31 53 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.25 //y=6.825 //x2=78.25 //y2=6.74
r111 (  29 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=78.165 //y=6.91 //x2=78.25 //y2=6.91
r112 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=78.165 //y=6.91 //x2=77.455 //y2=6.91
r113 (  23 52 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=77.37 //y=5.21 //x2=77.37 //y2=6.06
r114 (  21 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=77.37 //y=6.825 //x2=77.455 //y2=6.91
r115 (  21 52 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=77.37 //y=6.825 //x2=77.37 //y2=6.74
r116 (  15 48 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=75.37 //y=5.295 //x2=75.37 //y2=5.17
r117 (  15 51 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=75.37 //y=5.295 //x2=75.37 //y2=6.06
r118 (  13 48 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=75.285 //y=5.21 //x2=75.37 //y2=5.17
r119 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=75.285 //y=5.21 //x2=74.575 //y2=5.21
r120 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=74.49 //y=5.295 //x2=74.575 //y2=5.21
r121 (  7 50 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=74.49 //y=5.295 //x2=74.49 //y2=5.72
r122 (  6 23 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=77.37 //y=5.21 //x2=77.37 //y2=5.21
r123 (  4 48 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=75.37 //y=5.21 //x2=75.37 //y2=5.21
r124 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=75.485 //y=5.21 //x2=75.37 //y2=5.21
r125 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=77.255 //y=5.21 //x2=77.37 //y2=5.21
r126 (  1 2 ) resistor r=1.68893 //w=0.131 //l=1.77 //layer=m1 \
 //thickness=0.36 //x=77.255 //y=5.21 //x2=75.485 //y2=5.21
ends PM_TMRDFFSNQX1\%noxref_22

subckt PM_TMRDFFSNQX1\%noxref_23 ( 1 2 3 4 5 6 15 17 27 28 35 43 49 50 54 56 \
 64 73 74 75 76 77 78 79 80 81 82 83 84 85 86 91 93 95 101 102 103 104 105 106 \
 110 112 115 116 117 118 122 123 124 125 129 131 137 138 140 141 144 153 166 \
 169 171 172 173 )
c364 ( 173 0 ) capacitor c=0.023087f //x=71.595 //y=5.02
c365 ( 172 0 ) capacitor c=0.023519f //x=70.715 //y=5.02
c366 ( 171 0 ) capacitor c=0.0224735f //x=69.835 //y=5.02
c367 ( 169 0 ) capacitor c=0.0087111f //x=71.845 //y=0.915
c368 ( 166 0 ) capacitor c=0.0655948f //x=77.7 //y=4.705
c369 ( 153 0 ) capacitor c=0.0545009f //x=74 //y=2.08
c370 ( 144 0 ) capacitor c=0.0331706f //x=67 //y=4.7
c371 ( 141 0 ) capacitor c=0.0279499f //x=66.97 //y=1.915
c372 ( 140 0 ) capacitor c=0.0421676f //x=66.97 //y=2.08
c373 ( 138 0 ) capacitor c=0.0342409f //x=78.035 //y=1.21
c374 ( 137 0 ) capacitor c=0.0187384f //x=78.035 //y=0.865
c375 ( 131 0 ) capacitor c=0.0141797f //x=77.88 //y=1.365
c376 ( 129 0 ) capacitor c=0.0149844f //x=77.88 //y=0.71
c377 ( 125 0 ) capacitor c=0.10193f //x=77.505 //y=1.915
c378 ( 124 0 ) capacitor c=0.0225105f //x=77.505 //y=1.52
c379 ( 123 0 ) capacitor c=0.0234376f //x=77.505 //y=1.21
c380 ( 122 0 ) capacitor c=0.0199343f //x=77.505 //y=0.865
c381 ( 118 0 ) capacitor c=0.0318948f //x=74.705 //y=1.21
c382 ( 117 0 ) capacitor c=0.0187384f //x=74.705 //y=0.865
c383 ( 116 0 ) capacitor c=0.0607141f //x=74.345 //y=4.795
c384 ( 115 0 ) capacitor c=0.0292043f //x=74.635 //y=4.795
c385 ( 112 0 ) capacitor c=0.0157913f //x=74.55 //y=1.365
c386 ( 110 0 ) capacitor c=0.0149844f //x=74.55 //y=0.71
c387 ( 106 0 ) capacitor c=0.0302441f //x=74.175 //y=1.915
c388 ( 105 0 ) capacitor c=0.0238107f //x=74.175 //y=1.52
c389 ( 104 0 ) capacitor c=0.0234352f //x=74.175 //y=1.21
c390 ( 103 0 ) capacitor c=0.0199931f //x=74.175 //y=0.865
c391 ( 102 0 ) capacitor c=0.0429696f //x=67.535 //y=1.25
c392 ( 101 0 ) capacitor c=0.0192208f //x=67.535 //y=0.905
c393 ( 95 0 ) capacitor c=0.0148884f //x=67.38 //y=1.405
c394 ( 93 0 ) capacitor c=0.0157803f //x=67.38 //y=0.75
c395 ( 91 0 ) capacitor c=0.0295235f //x=67.375 //y=4.79
c396 ( 86 0 ) capacitor c=0.0205163f //x=67.005 //y=1.56
c397 ( 85 0 ) capacitor c=0.0168481f //x=67.005 //y=1.25
c398 ( 84 0 ) capacitor c=0.0174783f //x=67.005 //y=0.905
c399 ( 83 0 ) capacitor c=0.110336f //x=78.03 //y=6.025
c400 ( 82 0 ) capacitor c=0.154049f //x=77.59 //y=6.025
c401 ( 81 0 ) capacitor c=0.110003f //x=74.71 //y=6.025
c402 ( 80 0 ) capacitor c=0.15424f //x=74.27 //y=6.025
c403 ( 79 0 ) capacitor c=0.15358f //x=67.45 //y=6.02
c404 ( 78 0 ) capacitor c=0.110281f //x=67.01 //y=6.02
c405 ( 74 0 ) capacitor c=0.00106608f //x=71.74 //y=5.155
c406 ( 73 0 ) capacitor c=0.00207319f //x=70.86 //y=5.155
c407 ( 64 0 ) capacitor c=0.117496f //x=77.7 //y=2.08
c408 ( 56 0 ) capacitor c=0.0977815f //x=74 //y=2.08
c409 ( 54 0 ) capacitor c=0.107824f //x=72.52 //y=4.44
c410 ( 50 0 ) capacitor c=0.00463522f //x=72.12 //y=1.665
c411 ( 49 0 ) capacitor c=0.0148737f //x=72.435 //y=1.665
c412 ( 43 0 ) capacitor c=0.0281823f //x=72.435 //y=5.155
c413 ( 35 0 ) capacitor c=0.0176454f //x=71.655 //y=5.155
c414 ( 28 0 ) capacitor c=0.00332903f //x=70.065 //y=5.155
c415 ( 27 0 ) capacitor c=0.0148427f //x=70.775 //y=5.155
c416 ( 17 0 ) capacitor c=0.0713479f //x=66.97 //y=2.08
c417 ( 15 0 ) capacitor c=0.00369614f //x=66.97 //y=4.535
c418 ( 6 0 ) capacitor c=0.00522811f //x=74.115 //y=4.44
c419 ( 5 0 ) capacitor c=0.085624f //x=77.585 //y=4.44
c420 ( 4 0 ) capacitor c=0.0060226f //x=72.635 //y=4.44
c421 ( 3 0 ) capacitor c=0.0410264f //x=73.885 //y=4.44
c422 ( 2 0 ) capacitor c=0.0120792f //x=67.085 //y=4.44
c423 ( 1 0 ) capacitor c=0.11349f //x=72.405 //y=4.44
r424 (  164 166 ) resistor r=22.7554 //w=0.233 //l=0.11 //layer=ply \
 //thickness=0.18 //x=77.59 //y=4.705 //x2=77.7 //y2=4.705
r425 (  146 147 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=67 //y=4.79 //x2=67 //y2=4.865
r426 (  144 146 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=67 //y=4.7 //x2=67 //y2=4.79
r427 (  140 141 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=66.97 //y=2.08 //x2=66.97 //y2=1.915
r428 (  138 168 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.035 //y=1.21 //x2=77.995 //y2=1.365
r429 (  137 167 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.035 //y=0.865 //x2=77.995 //y2=0.71
r430 (  137 138 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=78.035 //y=0.865 //x2=78.035 //y2=1.21
r431 (  134 166 ) resistor r=68.2661 //w=0.233 //l=0.404166 //layer=ply \
 //thickness=0.18 //x=78.03 //y=4.87 //x2=77.7 //y2=4.705
r432 (  132 163 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=77.66 //y=1.365 //x2=77.545 //y2=1.365
r433 (  131 168 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=77.88 //y=1.365 //x2=77.995 //y2=1.365
r434 (  130 162 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=77.66 //y=0.71 //x2=77.545 //y2=0.71
r435 (  129 167 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=77.88 //y=0.71 //x2=77.995 //y2=0.71
r436 (  129 130 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=77.88 //y=0.71 //x2=77.66 //y2=0.71
r437 (  126 164 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=77.59 //y=4.87 //x2=77.59 //y2=4.705
r438 (  125 161 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=77.505 //y=1.915 //x2=77.7 //y2=2.08
r439 (  124 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=77.505 //y=1.52 //x2=77.545 //y2=1.365
r440 (  124 125 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=77.505 //y=1.52 //x2=77.505 //y2=1.915
r441 (  123 163 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=77.505 //y=1.21 //x2=77.545 //y2=1.365
r442 (  122 162 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=77.505 //y=0.865 //x2=77.545 //y2=0.71
r443 (  122 123 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=77.505 //y=0.865 //x2=77.505 //y2=1.21
r444 (  118 159 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.705 //y=1.21 //x2=74.665 //y2=1.365
r445 (  117 158 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.705 //y=0.865 //x2=74.665 //y2=0.71
r446 (  117 118 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=74.705 //y=0.865 //x2=74.705 //y2=1.21
r447 (  115 119 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=74.635 //y=4.795 //x2=74.71 //y2=4.87
r448 (  115 116 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=74.635 //y=4.795 //x2=74.345 //y2=4.795
r449 (  113 157 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.33 //y=1.365 //x2=74.215 //y2=1.365
r450 (  112 159 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.55 //y=1.365 //x2=74.665 //y2=1.365
r451 (  111 156 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.33 //y=0.71 //x2=74.215 //y2=0.71
r452 (  110 158 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=74.55 //y=0.71 //x2=74.665 //y2=0.71
r453 (  110 111 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=74.55 //y=0.71 //x2=74.33 //y2=0.71
r454 (  107 116 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=74.27 //y=4.87 //x2=74.345 //y2=4.795
r455 (  107 155 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=74.27 //y=4.87 //x2=74 //y2=4.705
r456 (  106 153 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=74.175 //y=1.915 //x2=74 //y2=2.08
r457 (  105 157 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.175 //y=1.52 //x2=74.215 //y2=1.365
r458 (  105 106 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=74.175 //y=1.52 //x2=74.175 //y2=1.915
r459 (  104 157 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.175 //y=1.21 //x2=74.215 //y2=1.365
r460 (  103 156 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=74.175 //y=0.865 //x2=74.215 //y2=0.71
r461 (  103 104 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=74.175 //y=0.865 //x2=74.175 //y2=1.21
r462 (  102 151 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=67.535 //y=1.25 //x2=67.495 //y2=1.405
r463 (  101 150 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=67.535 //y=0.905 //x2=67.495 //y2=0.75
r464 (  101 102 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=67.535 //y=0.905 //x2=67.535 //y2=1.25
r465 (  96 149 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=67.16 //y=1.405 //x2=67.045 //y2=1.405
r466 (  95 151 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=67.38 //y=1.405 //x2=67.495 //y2=1.405
r467 (  94 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=67.16 //y=0.75 //x2=67.045 //y2=0.75
r468 (  93 150 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=67.38 //y=0.75 //x2=67.495 //y2=0.75
r469 (  93 94 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=67.38 //y=0.75 //x2=67.16 //y2=0.75
r470 (  92 146 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=67.135 //y=4.79 //x2=67 //y2=4.79
r471 (  91 98 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=67.375 //y=4.79 //x2=67.45 //y2=4.865
r472 (  91 92 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=67.375 //y=4.79 //x2=67.135 //y2=4.79
r473 (  86 149 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=67.005 //y=1.56 //x2=67.045 //y2=1.405
r474 (  86 141 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=67.005 //y=1.56 //x2=67.005 //y2=1.915
r475 (  85 149 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=67.005 //y=1.25 //x2=67.045 //y2=1.405
r476 (  84 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=67.005 //y=0.905 //x2=67.045 //y2=0.75
r477 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=67.005 //y=0.905 //x2=67.005 //y2=1.25
r478 (  83 134 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=78.03 //y=6.025 //x2=78.03 //y2=4.87
r479 (  82 126 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=77.59 //y=6.025 //x2=77.59 //y2=4.87
r480 (  81 119 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=74.71 //y=6.025 //x2=74.71 //y2=4.87
r481 (  80 107 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=74.27 //y=6.025 //x2=74.27 //y2=4.87
r482 (  79 98 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=67.45 //y=6.02 //x2=67.45 //y2=4.865
r483 (  78 147 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=67.01 //y=6.02 //x2=67.01 //y2=4.865
r484 (  77 131 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=77.77 //y=1.365 //x2=77.88 //y2=1.365
r485 (  77 132 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=77.77 //y=1.365 //x2=77.66 //y2=1.365
r486 (  76 112 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=74.44 //y=1.365 //x2=74.55 //y2=1.365
r487 (  76 113 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=74.44 //y=1.365 //x2=74.33 //y2=1.365
r488 (  75 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=67.27 //y=1.405 //x2=67.38 //y2=1.405
r489 (  75 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=67.27 //y=1.405 //x2=67.16 //y2=1.405
r490 (  72 144 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=67 //y=4.7 //x2=67 //y2=4.7
r491 (  69 166 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=77.7 //y=4.705 //x2=77.7 //y2=4.705
r492 (  67 69 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=77.7 //y=4.44 //x2=77.7 //y2=4.705
r493 (  64 161 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=77.7 //y=2.08 //x2=77.7 //y2=2.08
r494 (  64 67 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=77.7 //y=2.08 //x2=77.7 //y2=4.44
r495 (  61 155 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=74 //y=4.705 //x2=74 //y2=4.705
r496 (  59 61 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=74 //y=4.44 //x2=74 //y2=4.705
r497 (  56 153 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=74 //y=2.08 //x2=74 //y2=2.08
r498 (  56 59 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=74 //y=2.08 //x2=74 //y2=4.44
r499 (  52 54 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=72.52 //y=5.07 //x2=72.52 //y2=4.44
r500 (  51 54 ) resistor r=184.128 //w=0.187 //l=2.69 //layer=li \
 //thickness=0.1 //x=72.52 //y=1.75 //x2=72.52 //y2=4.44
r501 (  49 51 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=72.435 //y=1.665 //x2=72.52 //y2=1.75
r502 (  49 50 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=72.435 //y=1.665 //x2=72.12 //y2=1.665
r503 (  45 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=72.035 //y=1.58 //x2=72.12 //y2=1.665
r504 (  45 169 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=72.035 //y=1.58 //x2=72.035 //y2=1.01
r505 (  44 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.825 //y=5.155 //x2=71.74 //y2=5.155
r506 (  43 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=72.435 //y=5.155 //x2=72.52 //y2=5.07
r507 (  43 44 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=72.435 //y=5.155 //x2=71.825 //y2=5.155
r508 (  37 74 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.74 //y=5.24 //x2=71.74 //y2=5.155
r509 (  37 173 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=71.74 //y=5.24 //x2=71.74 //y2=5.725
r510 (  36 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.945 //y=5.155 //x2=70.86 //y2=5.155
r511 (  35 74 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=71.655 //y=5.155 //x2=71.74 //y2=5.155
r512 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=71.655 //y=5.155 //x2=70.945 //y2=5.155
r513 (  29 73 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.86 //y=5.24 //x2=70.86 //y2=5.155
r514 (  29 172 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=70.86 //y=5.24 //x2=70.86 //y2=5.725
r515 (  27 73 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.775 //y=5.155 //x2=70.86 //y2=5.155
r516 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=70.775 //y=5.155 //x2=70.065 //y2=5.155
r517 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=69.98 //y=5.24 //x2=70.065 //y2=5.155
r518 (  21 171 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=69.98 //y=5.24 //x2=69.98 //y2=5.725
r519 (  17 140 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=66.97 //y=2.08 //x2=66.97 //y2=2.08
r520 (  17 20 ) resistor r=161.54 //w=0.187 //l=2.36 //layer=li \
 //thickness=0.1 //x=66.97 //y=2.08 //x2=66.97 //y2=4.44
r521 (  15 72 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=66.97 //y=4.535 //x2=66.985 //y2=4.7
r522 (  15 20 ) resistor r=6.50267 //w=0.187 //l=0.095 //layer=li \
 //thickness=0.1 //x=66.97 //y=4.535 //x2=66.97 //y2=4.44
r523 (  14 67 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=77.7 //y=4.44 //x2=77.7 //y2=4.44
r524 (  12 59 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 //x=74 \
 //y=4.44 //x2=74 //y2=4.44
r525 (  10 54 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=72.52 //y=4.44 //x2=72.52 //y2=4.44
r526 (  8 20 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=66.97 //y=4.44 //x2=66.97 //y2=4.44
r527 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=74.115 //y=4.44 //x2=74 //y2=4.44
r528 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=77.585 //y=4.44 //x2=77.7 //y2=4.44
r529 (  5 6 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=77.585 //y=4.44 //x2=74.115 //y2=4.44
r530 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=72.635 //y=4.44 //x2=72.52 //y2=4.44
r531 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=73.885 //y=4.44 //x2=74 //y2=4.44
r532 (  3 4 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=73.885 //y=4.44 //x2=72.635 //y2=4.44
r533 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=67.085 //y=4.44 //x2=66.97 //y2=4.44
r534 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=72.405 //y=4.44 //x2=72.52 //y2=4.44
r535 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=72.405 //y=4.44 //x2=67.085 //y2=4.44
ends PM_TMRDFFSNQX1\%noxref_23

subckt PM_TMRDFFSNQX1\%noxref_24 ( 1 2 3 4 5 6 17 19 29 30 37 45 51 52 56 58 \
 67 75 76 77 78 79 80 81 82 83 84 85 86 87 88 93 95 97 103 104 108 109 110 111 \
 112 114 117 120 121 122 123 124 125 126 127 131 133 136 137 138 139 144 145 \
 148 165 172 174 175 176 )
c474 ( 176 0 ) capacitor c=0.023087f //x=22.755 //y=5.02
c475 ( 175 0 ) capacitor c=0.023519f //x=21.875 //y=5.02
c476 ( 174 0 ) capacitor c=0.0224735f //x=20.995 //y=5.02
c477 ( 172 0 ) capacitor c=0.00872971f //x=23.005 //y=0.915
c478 ( 165 0 ) capacitor c=0.0583848f //x=80.66 //y=2.08
c479 ( 148 0 ) capacitor c=0.0331095f //x=18.16 //y=4.7
c480 ( 145 0 ) capacitor c=0.0279499f //x=18.13 //y=1.915
c481 ( 144 0 ) capacitor c=0.0421676f //x=18.13 //y=2.08
c482 ( 139 0 ) capacitor c=0.0316774f //x=81.365 //y=1.21
c483 ( 138 0 ) capacitor c=0.0187384f //x=81.365 //y=0.865
c484 ( 137 0 ) capacitor c=0.0590362f //x=81.005 //y=4.795
c485 ( 136 0 ) capacitor c=0.0296075f //x=81.295 //y=4.795
c486 ( 133 0 ) capacitor c=0.0157912f //x=81.21 //y=1.365
c487 ( 131 0 ) capacitor c=0.0149844f //x=81.21 //y=0.71
c488 ( 127 0 ) capacitor c=0.0302441f //x=80.835 //y=1.915
c489 ( 126 0 ) capacitor c=0.0234157f //x=80.835 //y=1.52
c490 ( 125 0 ) capacitor c=0.0234376f //x=80.835 //y=1.21
c491 ( 124 0 ) capacitor c=0.0199931f //x=80.835 //y=0.865
c492 ( 123 0 ) capacitor c=0.0962905f //x=79.005 //y=1.915
c493 ( 122 0 ) capacitor c=0.0249466f //x=79.005 //y=1.56
c494 ( 121 0 ) capacitor c=0.0234397f //x=79.005 //y=1.25
c495 ( 120 0 ) capacitor c=0.0193195f //x=79.005 //y=0.905
c496 ( 117 0 ) capacitor c=0.0631944f //x=78.91 //y=4.87
c497 ( 114 0 ) capacitor c=0.0187941f //x=78.85 //y=1.405
c498 ( 112 0 ) capacitor c=0.0157803f //x=78.85 //y=0.75
c499 ( 111 0 ) capacitor c=0.010629f //x=78.545 //y=4.795
c500 ( 110 0 ) capacitor c=0.0194269f //x=78.835 //y=4.795
c501 ( 109 0 ) capacitor c=0.0365717f //x=78.475 //y=1.25
c502 ( 108 0 ) capacitor c=0.0175988f //x=78.475 //y=0.905
c503 ( 104 0 ) capacitor c=0.0429696f //x=18.695 //y=1.25
c504 ( 103 0 ) capacitor c=0.0192208f //x=18.695 //y=0.905
c505 ( 97 0 ) capacitor c=0.0148884f //x=18.54 //y=1.405
c506 ( 95 0 ) capacitor c=0.0157803f //x=18.54 //y=0.75
c507 ( 93 0 ) capacitor c=0.0295235f //x=18.535 //y=4.79
c508 ( 88 0 ) capacitor c=0.0205163f //x=18.165 //y=1.56
c509 ( 87 0 ) capacitor c=0.0168481f //x=18.165 //y=1.25
c510 ( 86 0 ) capacitor c=0.0174783f //x=18.165 //y=0.905
c511 ( 85 0 ) capacitor c=0.110622f //x=81.37 //y=6.025
c512 ( 84 0 ) capacitor c=0.154068f //x=80.93 //y=6.025
c513 ( 83 0 ) capacitor c=0.154291f //x=78.91 //y=6.025
c514 ( 82 0 ) capacitor c=0.110404f //x=78.47 //y=6.025
c515 ( 81 0 ) capacitor c=0.15358f //x=18.61 //y=6.02
c516 ( 80 0 ) capacitor c=0.110281f //x=18.17 //y=6.02
c517 ( 76 0 ) capacitor c=0.00106608f //x=22.9 //y=5.155
c518 ( 75 0 ) capacitor c=0.00207319f //x=22.02 //y=5.155
c519 ( 67 0 ) capacitor c=0.100881f //x=80.66 //y=2.08
c520 ( 58 0 ) capacitor c=0.105667f //x=79.18 //y=2.08
c521 ( 56 0 ) capacitor c=0.110278f //x=23.68 //y=3.33
c522 ( 52 0 ) capacitor c=0.00398962f //x=23.28 //y=1.665
c523 ( 51 0 ) capacitor c=0.0137288f //x=23.595 //y=1.665
c524 ( 45 0 ) capacitor c=0.0284988f //x=23.595 //y=5.155
c525 ( 37 0 ) capacitor c=0.0176454f //x=22.815 //y=5.155
c526 ( 30 0 ) capacitor c=0.00332903f //x=21.225 //y=5.155
c527 ( 29 0 ) capacitor c=0.0148427f //x=21.935 //y=5.155
c528 ( 19 0 ) capacitor c=0.0698389f //x=18.13 //y=2.08
c529 ( 17 0 ) capacitor c=0.00453889f //x=18.13 //y=4.535
c530 ( 6 0 ) capacitor c=0.0112698f //x=79.295 //y=2.08
c531 ( 5 0 ) capacitor c=0.0463273f //x=80.545 //y=2.08
c532 ( 4 0 ) capacitor c=0.00605889f //x=23.795 //y=3.33
c533 ( 3 0 ) capacitor c=0.948787f //x=79.065 //y=3.33
c534 ( 2 0 ) capacitor c=0.0137368f //x=18.245 //y=3.33
c535 ( 1 0 ) capacitor c=0.0790615f //x=23.565 //y=3.33
r536 (  150 151 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=18.16 //y=4.79 //x2=18.16 //y2=4.865
r537 (  148 150 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=18.16 //y=4.7 //x2=18.16 //y2=4.79
r538 (  144 145 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=18.13 //y=2.08 //x2=18.13 //y2=1.915
r539 (  139 171 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=81.365 //y=1.21 //x2=81.325 //y2=1.365
r540 (  138 170 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=81.365 //y=0.865 //x2=81.325 //y2=0.71
r541 (  138 139 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=81.365 //y=0.865 //x2=81.365 //y2=1.21
r542 (  136 140 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=81.295 //y=4.795 //x2=81.37 //y2=4.87
r543 (  136 137 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=81.295 //y=4.795 //x2=81.005 //y2=4.795
r544 (  134 169 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=80.99 //y=1.365 //x2=80.875 //y2=1.365
r545 (  133 171 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=81.21 //y=1.365 //x2=81.325 //y2=1.365
r546 (  132 168 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=80.99 //y=0.71 //x2=80.875 //y2=0.71
r547 (  131 170 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=81.21 //y=0.71 //x2=81.325 //y2=0.71
r548 (  131 132 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=81.21 //y=0.71 //x2=80.99 //y2=0.71
r549 (  128 137 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=80.93 //y=4.87 //x2=81.005 //y2=4.795
r550 (  128 167 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=80.93 //y=4.87 //x2=80.66 //y2=4.705
r551 (  127 165 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=80.835 //y=1.915 //x2=80.66 //y2=2.08
r552 (  126 169 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.835 //y=1.52 //x2=80.875 //y2=1.365
r553 (  126 127 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=80.835 //y=1.52 //x2=80.835 //y2=1.915
r554 (  125 169 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.835 //y=1.21 //x2=80.875 //y2=1.365
r555 (  124 168 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=80.835 //y=0.865 //x2=80.875 //y2=0.71
r556 (  124 125 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=80.835 //y=0.865 //x2=80.835 //y2=1.21
r557 (  123 161 ) resistor r=30.4513 //w=0.277 //l=0.243926 //layer=ply \
 //thickness=0.18 //x=79.005 //y=1.915 //x2=79.18 //y2=2.08
r558 (  122 159 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.005 //y=1.56 //x2=78.965 //y2=1.405
r559 (  122 123 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=79.005 //y=1.56 //x2=79.005 //y2=1.915
r560 (  121 159 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.005 //y=1.25 //x2=78.965 //y2=1.405
r561 (  120 158 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=79.005 //y=0.905 //x2=78.965 //y2=0.75
r562 (  120 121 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=79.005 //y=0.905 //x2=79.005 //y2=1.25
r563 (  117 163 ) resistor r=51.6429 //w=0.252 //l=0.34271 //layer=ply \
 //thickness=0.18 //x=78.91 //y=4.87 //x2=79.18 //y2=4.705
r564 (  115 157 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.63 //y=1.405 //x2=78.515 //y2=1.405
r565 (  114 159 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.85 //y=1.405 //x2=78.965 //y2=1.405
r566 (  113 156 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.63 //y=0.75 //x2=78.515 //y2=0.75
r567 (  112 158 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=78.85 //y=0.75 //x2=78.965 //y2=0.75
r568 (  112 113 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=78.85 //y=0.75 //x2=78.63 //y2=0.75
r569 (  110 117 ) resistor r=22.1787 //w=0.252 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=78.835 //y=4.795 //x2=78.91 //y2=4.87
r570 (  110 111 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=78.835 //y=4.795 //x2=78.545 //y2=4.795
r571 (  109 157 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.475 //y=1.25 //x2=78.515 //y2=1.405
r572 (  108 156 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=78.475 //y=0.905 //x2=78.515 //y2=0.75
r573 (  108 109 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=78.475 //y=0.905 //x2=78.475 //y2=1.25
r574 (  105 111 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=78.47 //y=4.87 //x2=78.545 //y2=4.795
r575 (  104 155 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.695 //y=1.25 //x2=18.655 //y2=1.405
r576 (  103 154 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.695 //y=0.905 //x2=18.655 //y2=0.75
r577 (  103 104 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.695 //y=0.905 //x2=18.695 //y2=1.25
r578 (  98 153 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.32 //y=1.405 //x2=18.205 //y2=1.405
r579 (  97 155 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.54 //y=1.405 //x2=18.655 //y2=1.405
r580 (  96 152 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.32 //y=0.75 //x2=18.205 //y2=0.75
r581 (  95 154 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.54 //y=0.75 //x2=18.655 //y2=0.75
r582 (  95 96 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=18.54 //y=0.75 //x2=18.32 //y2=0.75
r583 (  94 150 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=18.295 //y=4.79 //x2=18.16 //y2=4.79
r584 (  93 100 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=18.535 //y=4.79 //x2=18.61 //y2=4.865
r585 (  93 94 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=18.535 //y=4.79 //x2=18.295 //y2=4.79
r586 (  88 153 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.165 //y=1.56 //x2=18.205 //y2=1.405
r587 (  88 145 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=18.165 //y=1.56 //x2=18.165 //y2=1.915
r588 (  87 153 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.165 //y=1.25 //x2=18.205 //y2=1.405
r589 (  86 152 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.165 //y=0.905 //x2=18.205 //y2=0.75
r590 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.165 //y=0.905 //x2=18.165 //y2=1.25
r591 (  85 140 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=81.37 //y=6.025 //x2=81.37 //y2=4.87
r592 (  84 128 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=80.93 //y=6.025 //x2=80.93 //y2=4.87
r593 (  83 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=78.91 //y=6.025 //x2=78.91 //y2=4.87
r594 (  82 105 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=78.47 //y=6.025 //x2=78.47 //y2=4.87
r595 (  81 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.61 //y=6.02 //x2=18.61 //y2=4.865
r596 (  80 151 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=18.17 //y=6.02 //x2=18.17 //y2=4.865
r597 (  79 133 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=81.1 //y=1.365 //x2=81.21 //y2=1.365
r598 (  79 134 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=81.1 //y=1.365 //x2=80.99 //y2=1.365
r599 (  78 114 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=78.74 //y=1.405 //x2=78.85 //y2=1.405
r600 (  78 115 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=78.74 //y=1.405 //x2=78.63 //y2=1.405
r601 (  77 97 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.43 //y=1.405 //x2=18.54 //y2=1.405
r602 (  77 98 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.43 //y=1.405 //x2=18.32 //y2=1.405
r603 (  74 148 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.16 //y=4.7 //x2=18.16 //y2=4.7
r604 (  71 167 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=80.66 //y=4.705 //x2=80.66 //y2=4.705
r605 (  67 165 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=80.66 //y=2.08 //x2=80.66 //y2=2.08
r606 (  67 71 ) resistor r=179.679 //w=0.187 //l=2.625 //layer=li \
 //thickness=0.1 //x=80.66 //y=2.08 //x2=80.66 //y2=4.705
r607 (  64 163 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=79.18 //y=4.705 //x2=79.18 //y2=4.705
r608 (  62 64 ) resistor r=94.1176 //w=0.187 //l=1.375 //layer=li \
 //thickness=0.1 //x=79.18 //y=3.33 //x2=79.18 //y2=4.705
r609 (  58 161 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=79.18 //y=2.08 //x2=79.18 //y2=2.08
r610 (  58 62 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=79.18 //y=2.08 //x2=79.18 //y2=3.33
r611 (  54 56 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=23.68 //y=5.07 //x2=23.68 //y2=3.33
r612 (  53 56 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=23.68 //y=1.75 //x2=23.68 //y2=3.33
r613 (  51 53 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.595 //y=1.665 //x2=23.68 //y2=1.75
r614 (  51 52 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=23.595 //y=1.665 //x2=23.28 //y2=1.665
r615 (  47 52 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.195 //y=1.58 //x2=23.28 //y2=1.665
r616 (  47 172 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=23.195 //y=1.58 //x2=23.195 //y2=1.01
r617 (  46 76 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.985 //y=5.155 //x2=22.9 //y2=5.155
r618 (  45 54 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.595 //y=5.155 //x2=23.68 //y2=5.07
r619 (  45 46 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=23.595 //y=5.155 //x2=22.985 //y2=5.155
r620 (  39 76 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.9 //y=5.24 //x2=22.9 //y2=5.155
r621 (  39 176 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.9 //y=5.24 //x2=22.9 //y2=5.725
r622 (  38 75 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.105 //y=5.155 //x2=22.02 //y2=5.155
r623 (  37 76 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.815 //y=5.155 //x2=22.9 //y2=5.155
r624 (  37 38 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=22.815 //y=5.155 //x2=22.105 //y2=5.155
r625 (  31 75 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.02 //y=5.24 //x2=22.02 //y2=5.155
r626 (  31 175 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=22.02 //y=5.24 //x2=22.02 //y2=5.725
r627 (  29 75 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.935 //y=5.155 //x2=22.02 //y2=5.155
r628 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=21.935 //y=5.155 //x2=21.225 //y2=5.155
r629 (  23 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.14 //y=5.24 //x2=21.225 //y2=5.155
r630 (  23 174 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.14 //y=5.24 //x2=21.14 //y2=5.725
r631 (  19 144 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.13 //y=2.08 //x2=18.13 //y2=2.08
r632 (  19 22 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=18.13 //y=2.08 //x2=18.13 //y2=3.33
r633 (  17 74 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=18.13 //y=4.535 //x2=18.145 //y2=4.7
r634 (  17 22 ) resistor r=82.4813 //w=0.187 //l=1.205 //layer=li \
 //thickness=0.1 //x=18.13 //y=4.535 //x2=18.13 //y2=3.33
r635 (  16 67 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=80.66 //y=2.08 //x2=80.66 //y2=2.08
r636 (  14 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=79.18 //y=3.33 //x2=79.18 //y2=3.33
r637 (  12 58 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=79.18 //y=2.08 //x2=79.18 //y2=2.08
r638 (  10 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=23.68 //y=3.33 //x2=23.68 //y2=3.33
r639 (  8 22 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.13 //y=3.33 //x2=18.13 //y2=3.33
r640 (  6 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=79.295 //y=2.08 //x2=79.18 //y2=2.08
r641 (  5 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=80.545 //y=2.08 //x2=80.66 //y2=2.08
r642 (  5 6 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=80.545 //y=2.08 //x2=79.295 //y2=2.08
r643 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.795 //y=3.33 //x2=23.68 //y2=3.33
r644 (  3 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=79.065 //y=3.33 //x2=79.18 //y2=3.33
r645 (  3 4 ) resistor r=52.7385 //w=0.131 //l=55.27 //layer=m1 \
 //thickness=0.36 //x=79.065 //y=3.33 //x2=23.795 //y2=3.33
r646 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.245 //y=3.33 //x2=18.13 //y2=3.33
r647 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.565 //y=3.33 //x2=23.68 //y2=3.33
r648 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=23.565 //y=3.33 //x2=18.245 //y2=3.33
ends PM_TMRDFFSNQX1\%noxref_24

subckt PM_TMRDFFSNQX1\%noxref_25 ( 1 2 13 14 15 21 27 28 35 46 47 48 49 50 )
c90 ( 50 0 ) capacitor c=0.0306574f //x=82.325 //y=5.025
c91 ( 49 0 ) capacitor c=0.0173945f //x=81.445 //y=5.025
c92 ( 47 0 ) capacitor c=0.0169278f //x=78.545 //y=5.025
c93 ( 46 0 ) capacitor c=0.0166762f //x=77.665 //y=5.025
c94 ( 45 0 ) capacitor c=0.00115294f //x=81.59 //y=6.91
c95 ( 35 0 ) capacitor c=0.0132983f //x=82.385 //y=6.91
c96 ( 28 0 ) capacitor c=0.00388794f //x=80.795 //y=6.91
c97 ( 27 0 ) capacitor c=0.00985708f //x=81.505 //y=6.91
c98 ( 21 0 ) capacitor c=0.0442221f //x=80.71 //y=5.21
c99 ( 15 0 ) capacitor c=0.0105083f //x=78.69 //y=5.295
c100 ( 14 0 ) capacitor c=0.00227812f //x=77.895 //y=5.21
c101 ( 13 0 ) capacitor c=0.0174384f //x=78.605 //y=5.21
c102 ( 2 0 ) capacitor c=0.00682032f //x=78.805 //y=5.21
c103 ( 1 0 ) capacitor c=0.0573196f //x=80.595 //y=5.21
r104 (  37 50 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.47 //y=6.825 //x2=82.47 //y2=6.74
r105 (  36 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.675 //y=6.91 //x2=81.59 //y2=6.91
r106 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=82.385 //y=6.91 //x2=82.47 //y2=6.825
r107 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=82.385 //y=6.91 //x2=81.675 //y2=6.91
r108 (  29 45 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.59 //y=6.825 //x2=81.59 //y2=6.91
r109 (  29 49 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.59 //y=6.825 //x2=81.59 //y2=6.74
r110 (  27 45 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.505 //y=6.91 //x2=81.59 //y2=6.91
r111 (  27 28 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=81.505 //y=6.91 //x2=80.795 //y2=6.91
r112 (  21 48 ) resistor r=58.1818 //w=0.187 //l=0.85 //layer=li \
 //thickness=0.1 //x=80.71 //y=5.21 //x2=80.71 //y2=6.06
r113 (  19 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=80.71 //y=6.825 //x2=80.795 //y2=6.91
r114 (  19 48 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=80.71 //y=6.825 //x2=80.71 //y2=6.74
r115 (  15 44 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=78.69 //y=5.295 //x2=78.69 //y2=5.17
r116 (  15 47 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=78.69 //y=5.295 //x2=78.69 //y2=6.06
r117 (  13 44 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.605 //y=5.21 //x2=78.69 //y2=5.17
r118 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=78.605 //y=5.21 //x2=77.895 //y2=5.21
r119 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=77.81 //y=5.295 //x2=77.895 //y2=5.21
r120 (  7 46 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=77.81 //y=5.295 //x2=77.81 //y2=5.72
r121 (  6 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=80.71 //y=5.21 //x2=80.71 //y2=5.21
r122 (  4 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=78.69 //y=5.21 //x2=78.69 //y2=5.21
r123 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=78.805 //y=5.21 //x2=78.69 //y2=5.21
r124 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=80.595 //y=5.21 //x2=80.71 //y2=5.21
r125 (  1 2 ) resistor r=1.70802 //w=0.131 //l=1.79 //layer=m1 \
 //thickness=0.36 //x=80.595 //y=5.21 //x2=78.805 //y2=5.21
ends PM_TMRDFFSNQX1\%noxref_25

subckt PM_TMRDFFSNQX1\%noxref_26 ( 1 2 3 4 5 6 29 30 43 45 46 50 52 63 64 65 \
 66 67 68 69 70 74 75 76 78 84 85 87 95 96 97 101 102 )
c240 ( 102 0 ) capacitor c=0.0167617f //x=81.885 //y=5.025
c241 ( 101 0 ) capacitor c=0.0164812f //x=81.005 //y=5.025
c242 ( 97 0 ) capacitor c=0.0110092f //x=81.88 //y=0.905
c243 ( 96 0 ) capacitor c=0.0131637f //x=78.55 //y=0.905
c244 ( 95 0 ) capacitor c=0.0131367f //x=75.22 //y=0.905
c245 ( 87 0 ) capacitor c=0.0537799f //x=83.99 //y=2.085
c246 ( 85 0 ) capacitor c=0.0435629f //x=84.63 //y=1.255
c247 ( 84 0 ) capacitor c=0.0200386f //x=84.63 //y=0.91
c248 ( 78 0 ) capacitor c=0.0152946f //x=84.475 //y=1.41
c249 ( 76 0 ) capacitor c=0.0157804f //x=84.475 //y=0.755
c250 ( 75 0 ) capacitor c=0.05065f //x=84.22 //y=4.79
c251 ( 74 0 ) capacitor c=0.0322983f //x=84.51 //y=4.79
c252 ( 70 0 ) capacitor c=0.0290017f //x=84.1 //y=1.92
c253 ( 69 0 ) capacitor c=0.0250027f //x=84.1 //y=1.565
c254 ( 68 0 ) capacitor c=0.0234316f //x=84.1 //y=1.255
c255 ( 67 0 ) capacitor c=0.0200596f //x=84.1 //y=0.91
c256 ( 66 0 ) capacitor c=0.154218f //x=84.585 //y=6.02
c257 ( 65 0 ) capacitor c=0.154243f //x=84.145 //y=6.02
c258 ( 63 0 ) capacitor c=0.00421476f //x=82.03 //y=5.21
c259 ( 52 0 ) capacitor c=0.0942569f //x=83.99 //y=2.085
c260 ( 50 0 ) capacitor c=0.112965f //x=82.51 //y=4.07
c261 ( 46 0 ) capacitor c=0.00775877f //x=82.155 //y=1.645
c262 ( 45 0 ) capacitor c=0.0161066f //x=82.425 //y=1.645
c263 ( 43 0 ) capacitor c=0.0151634f //x=82.425 //y=5.21
c264 ( 30 0 ) capacitor c=0.0029383f //x=81.235 //y=5.21
c265 ( 29 0 ) capacitor c=0.0155464f //x=81.945 //y=5.21
c266 ( 6 0 ) capacitor c=0.00867855f //x=82.625 //y=4.07
c267 ( 5 0 ) capacitor c=0.0786471f //x=83.875 //y=4.07
c268 ( 4 0 ) capacitor c=0.0054338f //x=78.855 //y=1.18
c269 ( 3 0 ) capacitor c=0.0704773f //x=81.955 //y=1.18
c270 ( 2 0 ) capacitor c=0.0153777f //x=75.525 //y=1.18
c271 ( 1 0 ) capacitor c=0.0651236f //x=78.625 //y=1.18
r272 (  87 88 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=83.99 //y=2.085 //x2=84.1 //y2=2.085
r273 (  85 94 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=84.63 //y=1.255 //x2=84.59 //y2=1.41
r274 (  84 93 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=84.63 //y=0.91 //x2=84.59 //y2=0.755
r275 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=84.63 //y=0.91 //x2=84.63 //y2=1.255
r276 (  79 92 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=84.255 //y=1.41 //x2=84.14 //y2=1.41
r277 (  78 94 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=84.475 //y=1.41 //x2=84.59 //y2=1.41
r278 (  77 91 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=84.255 //y=0.755 //x2=84.14 //y2=0.755
r279 (  76 93 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=84.475 //y=0.755 //x2=84.59 //y2=0.755
r280 (  76 77 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=84.475 //y=0.755 //x2=84.255 //y2=0.755
r281 (  74 81 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=84.51 //y=4.79 //x2=84.585 //y2=4.865
r282 (  74 75 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=84.51 //y=4.79 //x2=84.22 //y2=4.79
r283 (  71 75 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=84.145 //y=4.865 //x2=84.22 //y2=4.79
r284 (  71 90 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=84.145 //y=4.865 //x2=83.99 //y2=4.7
r285 (  70 88 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=84.1 //y=1.92 //x2=84.1 //y2=2.085
r286 (  69 92 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=84.1 //y=1.565 //x2=84.14 //y2=1.41
r287 (  69 70 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=84.1 //y=1.565 //x2=84.1 //y2=1.92
r288 (  68 92 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=84.1 //y=1.255 //x2=84.14 //y2=1.41
r289 (  67 91 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=84.1 //y=0.91 //x2=84.14 //y2=0.755
r290 (  67 68 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=84.1 //y=0.91 //x2=84.1 //y2=1.255
r291 (  66 81 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=84.585 //y=6.02 //x2=84.585 //y2=4.865
r292 (  65 71 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=84.145 //y=6.02 //x2=84.145 //y2=4.865
r293 (  64 78 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=84.365 //y=1.41 //x2=84.475 //y2=1.41
r294 (  64 79 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=84.365 //y=1.41 //x2=84.255 //y2=1.41
r295 (  62 95 ) resistor r=13.3953 //w=0.172 //l=0.18 //layer=li \
 //thickness=0.1 //x=75.407 //y=1.18 //x2=75.407 //y2=1
r296 (  57 90 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=83.99 //y=4.7 //x2=83.99 //y2=4.7
r297 (  55 57 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=83.99 //y=4.07 //x2=83.99 //y2=4.7
r298 (  52 87 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=83.99 //y=2.085 //x2=83.99 //y2=2.085
r299 (  52 55 ) resistor r=135.872 //w=0.187 //l=1.985 //layer=li \
 //thickness=0.1 //x=83.99 //y=2.085 //x2=83.99 //y2=4.07
r300 (  48 50 ) resistor r=72.2139 //w=0.187 //l=1.055 //layer=li \
 //thickness=0.1 //x=82.51 //y=5.125 //x2=82.51 //y2=4.07
r301 (  47 50 ) resistor r=160.171 //w=0.187 //l=2.34 //layer=li \
 //thickness=0.1 //x=82.51 //y=1.73 //x2=82.51 //y2=4.07
r302 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=82.425 //y=1.645 //x2=82.51 //y2=1.73
r303 (  45 46 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=82.425 //y=1.645 //x2=82.155 //y2=1.645
r304 (  44 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.115 //y=5.21 //x2=82.03 //y2=5.21
r305 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=82.425 //y=5.21 //x2=82.51 //y2=5.125
r306 (  43 44 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=82.425 //y=5.21 //x2=82.115 //y2=5.21
r307 (  42 97 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=82.07 //y=1.18 //x2=82.07 //y2=1
r308 (  37 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=82.07 //y=1.56 //x2=82.155 //y2=1.645
r309 (  37 42 ) resistor r=26.0107 //w=0.187 //l=0.38 //layer=li \
 //thickness=0.1 //x=82.07 //y=1.56 //x2=82.07 //y2=1.18
r310 (  31 63 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=82.03 //y=5.295 //x2=82.03 //y2=5.21
r311 (  31 102 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=82.03 //y=5.295 //x2=82.03 //y2=5.72
r312 (  29 63 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=81.945 //y=5.21 //x2=82.03 //y2=5.21
r313 (  29 30 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=81.945 //y=5.21 //x2=81.235 //y2=5.21
r314 (  23 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=81.15 //y=5.295 //x2=81.235 //y2=5.21
r315 (  23 101 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=81.15 //y=5.295 //x2=81.15 //y2=5.72
r316 (  21 96 ) resistor r=12.3209 //w=0.187 //l=0.18 //layer=li \
 //thickness=0.1 //x=78.74 //y=1.18 //x2=78.74 //y2=1
r317 (  16 55 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=83.99 //y=4.07 //x2=83.99 //y2=4.07
r318 (  14 50 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=82.51 //y=4.07 //x2=82.51 //y2=4.07
r319 (  12 42 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=82.07 //y=1.18 //x2=82.07 //y2=1.18
r320 (  10 21 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=78.74 //y=1.18 //x2=78.74 //y2=1.18
r321 (  8 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=75.41 //y=1.18 //x2=75.41 //y2=1.18
r322 (  6 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=82.625 //y=4.07 //x2=82.51 //y2=4.07
r323 (  5 16 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=83.875 //y=4.07 //x2=83.99 //y2=4.07
r324 (  5 6 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=83.875 //y=4.07 //x2=82.625 //y2=4.07
r325 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=78.855 //y=1.18 //x2=78.74 //y2=1.18
r326 (  3 12 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=81.955 //y=1.18 //x2=82.07 //y2=1.18
r327 (  3 4 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=81.955 //y=1.18 //x2=78.855 //y2=1.18
r328 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=75.525 //y=1.18 //x2=75.41 //y2=1.18
r329 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=78.625 //y=1.18 //x2=78.74 //y2=1.18
r330 (  1 2 ) resistor r=2.95802 //w=0.131 //l=3.1 //layer=m1 //thickness=0.36 \
 //x=78.625 //y=1.18 //x2=75.525 //y2=1.18
ends PM_TMRDFFSNQX1\%noxref_26

subckt PM_TMRDFFSNQX1\%noxref_27 ( 1 5 9 10 13 17 29 )
c50 ( 29 0 ) capacitor c=0.0632971f //x=0.56 //y=0.365
c51 ( 17 0 ) capacitor c=0.0072343f //x=2.635 //y=0.615
c52 ( 13 0 ) capacitor c=0.0147753f //x=2.55 //y=0.53
c53 ( 10 0 ) capacitor c=0.00638095f //x=1.665 //y=1.495
c54 ( 9 0 ) capacitor c=0.006761f //x=1.665 //y=0.615
c55 ( 5 0 ) capacitor c=0.02021f //x=1.58 //y=1.58
c56 ( 1 0 ) capacitor c=0.0113547f //x=0.695 //y=1.495
r57 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.49
r58 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r59 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.75 //y=0.53 //x2=1.665 //y2=0.49
r60 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=2.15 //y2=0.53
r61 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.49
r62 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.55 //y=0.53 //x2=2.15 //y2=0.53
r63 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=1.62
r64 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.665 //y=1.495 //x2=1.665 //y2=0.88
r65 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.49
r66 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r67 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.78 //y=1.58 //x2=0.695 //y2=1.62
r68 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.78 //y=1.58 //x2=1.18 //y2=1.58
r69 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.58 //y=1.58 //x2=1.665 //y2=1.62
r70 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.58 //y=1.58 //x2=1.18 //y2=1.58
r71 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.695 //y=1.495 //x2=0.695 //y2=1.62
r72 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.695 //y=1.495 //x2=0.695 //y2=0.88
ends PM_TMRDFFSNQX1\%noxref_27

subckt PM_TMRDFFSNQX1\%noxref_28 ( 1 5 9 13 17 35 )
c51 ( 35 0 ) capacitor c=0.0680128f //x=3.785 //y=0.375
c52 ( 17 0 ) capacitor c=0.018806f //x=5.775 //y=1.59
c53 ( 13 0 ) capacitor c=0.0155484f //x=5.775 //y=0.54
c54 ( 9 0 ) capacitor c=0.00678203f //x=4.89 //y=0.625
c55 ( 5 0 ) capacitor c=0.017077f //x=4.805 //y=1.59
c56 ( 1 0 ) capacitor c=0.00729042f //x=3.92 //y=1.505
r57 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.975 //y=1.59 //x2=4.89 //y2=1.63
r58 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.975 //y=1.59 //x2=5.375 //y2=1.59
r59 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.775 //y=1.59 //x2=5.86 //y2=1.59
r60 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.775 //y=1.59 //x2=5.375 //y2=1.59
r61 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.975 //y=0.54 //x2=4.89 //y2=0.5
r62 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.975 //y=0.54 //x2=5.375 //y2=0.54
r63 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.775 //y=0.54 //x2=5.86 //y2=0.54
r64 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.775 //y=0.54 //x2=5.375 //y2=0.54
r65 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.89 //y=1.505 //x2=4.89 //y2=1.63
r66 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=4.89 //y=1.505 //x2=4.89 //y2=0.89
r67 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=4.89 //y=0.625 //x2=4.89 //y2=0.5
r68 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=4.89 //y=0.625 //x2=4.89 //y2=0.89
r69 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.005 //y=1.59 //x2=3.92 //y2=1.63
r70 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.005 //y=1.59 //x2=4.405 //y2=1.59
r71 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=4.805 //y=1.59 //x2=4.89 //y2=1.63
r72 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=4.805 //y=1.59 //x2=4.405 //y2=1.59
r73 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.92 //y=1.505 //x2=3.92 //y2=1.63
r74 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=3.92 //y=1.505 //x2=3.92 //y2=0.89
ends PM_TMRDFFSNQX1\%noxref_28

subckt PM_TMRDFFSNQX1\%noxref_29 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.041888f //x=6.295 //y=0.375
c53 ( 28 0 ) capacitor c=0.00460056f //x=5.19 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=6.43 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=7.4 //y=0.625
c56 ( 11 0 ) capacitor c=0.0145763f //x=7.315 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=6.43 //y=0.625
c58 ( 1 0 ) capacitor c=0.022715f //x=6.345 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=7.4 //y=0.625 //x2=7.4 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=7.4 //y=0.625 //x2=7.4 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.515 //y=0.54 //x2=6.43 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.515 //y=0.54 //x2=6.915 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.315 //y=0.54 //x2=7.4 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.315 //y=0.54 //x2=6.915 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=6.43 //y=1.08 //x2=6.43 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=6.43 //y=1.08 //x2=6.43 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.91 //x2=6.43 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.91 //x2=6.43 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.625 //x2=6.43 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.43 //y=0.625 //x2=6.43 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.465 //y=0.995 //x2=5.38 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=6.345 //y=0.995 //x2=6.43 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=6.345 //y=0.995 //x2=5.465 //y2=0.995
ends PM_TMRDFFSNQX1\%noxref_29

subckt PM_TMRDFFSNQX1\%noxref_30 ( 1 5 9 13 17 35 )
c53 ( 35 0 ) capacitor c=0.0679545f //x=8.595 //y=0.375
c54 ( 17 0 ) capacitor c=0.0193993f //x=10.585 //y=1.59
c55 ( 13 0 ) capacitor c=0.0155066f //x=10.585 //y=0.54
c56 ( 9 0 ) capacitor c=0.00678203f //x=9.7 //y=0.625
c57 ( 5 0 ) capacitor c=0.0174845f //x=9.615 //y=1.59
c58 ( 1 0 ) capacitor c=0.00729042f //x=8.73 //y=1.505
r59 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.785 //y=1.59 //x2=9.7 //y2=1.63
r60 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.785 //y=1.59 //x2=10.185 //y2=1.59
r61 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.585 //y=1.59 //x2=10.67 //y2=1.59
r62 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.585 //y=1.59 //x2=10.185 //y2=1.59
r63 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.785 //y=0.54 //x2=9.7 //y2=0.5
r64 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.785 //y=0.54 //x2=10.185 //y2=0.54
r65 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.585 //y=0.54 //x2=10.67 //y2=0.54
r66 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.585 //y=0.54 //x2=10.185 //y2=0.54
r67 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=9.7 //y=1.505 //x2=9.7 //y2=1.63
r68 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=9.7 //y=1.505 //x2=9.7 //y2=0.89
r69 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=9.7 //y=0.625 //x2=9.7 //y2=0.5
r70 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=9.7 //y=0.625 //x2=9.7 //y2=0.89
r71 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.815 //y=1.59 //x2=8.73 //y2=1.63
r72 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.815 //y=1.59 //x2=9.215 //y2=1.59
r73 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=9.615 //y=1.59 //x2=9.7 //y2=1.63
r74 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=9.615 //y=1.59 //x2=9.215 //y2=1.59
r75 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=8.73 //y=1.505 //x2=8.73 //y2=1.63
r76 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=8.73 //y=1.505 //x2=8.73 //y2=0.89
ends PM_TMRDFFSNQX1\%noxref_30

subckt PM_TMRDFFSNQX1\%noxref_31 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=11.105 //y=0.375
c53 ( 28 0 ) capacitor c=0.00460343f //x=10 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=11.24 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=12.21 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=12.125 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=11.24 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=11.155 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=12.21 //y=0.625 //x2=12.21 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=12.21 //y=0.625 //x2=12.21 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.325 //y=0.54 //x2=11.24 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.325 //y=0.54 //x2=11.725 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.125 //y=0.54 //x2=12.21 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.125 //y=0.54 //x2=11.725 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.24 //y=1.08 //x2=11.24 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=11.24 //y=1.08 //x2=11.24 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.91 //x2=11.24 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.91 //x2=11.24 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.625 //x2=11.24 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=11.24 //y=0.625 //x2=11.24 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.275 //y=0.995 //x2=10.19 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=11.155 //y=0.995 //x2=11.24 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=11.155 //y=0.995 //x2=10.275 //y2=0.995
ends PM_TMRDFFSNQX1\%noxref_31

subckt PM_TMRDFFSNQX1\%noxref_32 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632682f //x=13.51 //y=0.365
c52 ( 17 0 ) capacitor c=0.00722223f //x=15.585 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=15.5 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=14.615 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=14.615 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=14.53 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=13.645 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=15.585 //y=0.615 //x2=15.585 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=15.585 //y=0.615 //x2=15.585 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.7 //y=0.53 //x2=14.615 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.7 //y=0.53 //x2=15.1 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=15.5 //y=0.53 //x2=15.585 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.5 //y=0.53 //x2=15.1 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=14.615 //y=1.495 //x2=14.615 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=14.615 //y=1.495 //x2=14.615 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=14.615 //y=0.615 //x2=14.615 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=14.615 //y=0.615 //x2=14.615 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.73 //y=1.58 //x2=13.645 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.73 //y=1.58 //x2=14.13 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.53 //y=1.58 //x2=14.615 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.53 //y=1.58 //x2=14.13 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=13.645 //y=1.495 //x2=13.645 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=13.645 //y=1.495 //x2=13.645 //y2=0.88
ends PM_TMRDFFSNQX1\%noxref_32

subckt PM_TMRDFFSNQX1\%noxref_33 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632684f //x=16.84 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=18.915 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=18.83 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=17.945 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=17.945 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=17.86 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=16.975 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=18.915 //y=0.615 //x2=18.915 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=18.915 //y=0.615 //x2=18.915 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.03 //y=0.53 //x2=17.945 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.03 //y=0.53 //x2=18.43 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.83 //y=0.53 //x2=18.915 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.83 //y=0.53 //x2=18.43 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=17.945 //y=1.495 //x2=17.945 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=17.945 //y=1.495 //x2=17.945 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=17.945 //y=0.615 //x2=17.945 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=17.945 //y=0.615 //x2=17.945 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.06 //y=1.58 //x2=16.975 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.06 //y=1.58 //x2=17.46 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=17.86 //y=1.58 //x2=17.945 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=17.86 //y=1.58 //x2=17.46 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=16.975 //y=1.495 //x2=16.975 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=16.975 //y=1.495 //x2=16.975 //y2=0.88
ends PM_TMRDFFSNQX1\%noxref_33

subckt PM_TMRDFFSNQX1\%noxref_34 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=20.065 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=22.055 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=22.055 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=21.17 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=21.085 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=20.2 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.255 //y=1.59 //x2=21.17 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.255 //y=1.59 //x2=21.655 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.055 //y=1.59 //x2=22.14 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.055 //y=1.59 //x2=21.655 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.255 //y=0.54 //x2=21.17 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.255 //y=0.54 //x2=21.655 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=22.055 //y=0.54 //x2=22.14 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.055 //y=0.54 //x2=21.655 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=21.17 //y=1.505 //x2=21.17 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=21.17 //y=1.505 //x2=21.17 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=21.17 //y=0.625 //x2=21.17 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=21.17 //y=0.625 //x2=21.17 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.285 //y=1.59 //x2=20.2 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.285 //y=1.59 //x2=20.685 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.085 //y=1.59 //x2=21.17 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.085 //y=1.59 //x2=20.685 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=20.2 //y=1.505 //x2=20.2 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=20.2 //y=1.505 //x2=20.2 //y2=0.89
ends PM_TMRDFFSNQX1\%noxref_34

subckt PM_TMRDFFSNQX1\%noxref_35 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0413887f //x=22.575 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=21.47 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=22.71 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=23.68 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=23.595 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=22.71 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=22.625 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=23.68 //y=0.625 //x2=23.68 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=23.68 //y=0.625 //x2=23.68 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=22.795 //y=0.54 //x2=22.71 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=22.795 //y=0.54 //x2=23.195 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.595 //y=0.54 //x2=23.68 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.595 //y=0.54 //x2=23.195 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.71 //y=1.08 //x2=22.71 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=22.71 //y=1.08 //x2=22.71 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.91 //x2=22.71 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.91 //x2=22.71 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.625 //x2=22.71 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=22.71 //y=0.625 //x2=22.71 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.745 //y=0.995 //x2=21.66 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=22.625 //y=0.995 //x2=22.71 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=22.625 //y=0.995 //x2=21.745 //y2=0.995
ends PM_TMRDFFSNQX1\%noxref_35

subckt PM_TMRDFFSNQX1\%noxref_36 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0633518f //x=24.98 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=27.055 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=26.97 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=26.085 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=26.085 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=26 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=25.115 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=27.055 //y=0.615 //x2=27.055 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=27.055 //y=0.615 //x2=27.055 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=26.17 //y=0.53 //x2=26.085 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.17 //y=0.53 //x2=26.57 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=26.97 //y=0.53 //x2=27.055 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26.97 //y=0.53 //x2=26.57 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=26.085 //y=1.495 //x2=26.085 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=26.085 //y=1.495 //x2=26.085 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=26.085 //y=0.615 //x2=26.085 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=26.085 //y=0.615 //x2=26.085 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.2 //y=1.58 //x2=25.115 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.2 //y=1.58 //x2=25.6 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=26 //y=1.58 //x2=26.085 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=26 //y=1.58 //x2=25.6 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=25.115 //y=1.495 //x2=25.115 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=25.115 //y=1.495 //x2=25.115 //y2=0.88
ends PM_TMRDFFSNQX1\%noxref_36

subckt PM_TMRDFFSNQX1\%noxref_37 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673195f //x=28.205 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=30.195 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=30.195 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=29.31 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=29.225 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=28.34 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=29.395 //y=1.59 //x2=29.31 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=29.395 //y=1.59 //x2=29.795 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.195 //y=1.59 //x2=30.28 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.195 //y=1.59 //x2=29.795 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=29.395 //y=0.54 //x2=29.31 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=29.395 //y=0.54 //x2=29.795 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=30.195 //y=0.54 //x2=30.28 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.195 //y=0.54 //x2=29.795 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=29.31 //y=1.505 //x2=29.31 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=29.31 //y=1.505 //x2=29.31 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=29.31 //y=0.625 //x2=29.31 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=29.31 //y=0.625 //x2=29.31 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=28.425 //y=1.59 //x2=28.34 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=28.425 //y=1.59 //x2=28.825 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=29.225 //y=1.59 //x2=29.31 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=29.225 //y=1.59 //x2=28.825 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=28.34 //y=1.505 //x2=28.34 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=28.34 //y=1.505 //x2=28.34 //y2=0.89
ends PM_TMRDFFSNQX1\%noxref_37

subckt PM_TMRDFFSNQX1\%noxref_38 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414739f //x=30.715 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=29.61 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=30.85 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=31.82 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=31.735 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=30.85 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=30.765 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=31.82 //y=0.625 //x2=31.82 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=31.82 //y=0.625 //x2=31.82 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=30.935 //y=0.54 //x2=30.85 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=30.935 //y=0.54 //x2=31.335 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=31.735 //y=0.54 //x2=31.82 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=31.735 //y=0.54 //x2=31.335 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=30.85 //y=1.08 //x2=30.85 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=30.85 //y=1.08 //x2=30.85 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=30.85 //y=0.91 //x2=30.85 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=30.85 //y=0.91 //x2=30.85 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=30.85 //y=0.625 //x2=30.85 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=30.85 //y=0.625 //x2=30.85 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=29.885 //y=0.995 //x2=29.8 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=30.765 //y=0.995 //x2=30.85 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=30.765 //y=0.995 //x2=29.885 //y2=0.995
ends PM_TMRDFFSNQX1\%noxref_38

subckt PM_TMRDFFSNQX1\%noxref_39 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=33.015 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=35.005 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=35.005 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=34.12 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=34.035 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=33.15 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=34.205 //y=1.59 //x2=34.12 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=34.205 //y=1.59 //x2=34.605 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.005 //y=1.59 //x2=35.09 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.005 //y=1.59 //x2=34.605 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=34.205 //y=0.54 //x2=34.12 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=34.205 //y=0.54 //x2=34.605 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=35.005 //y=0.54 //x2=35.09 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.005 //y=0.54 //x2=34.605 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=34.12 //y=1.505 //x2=34.12 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=34.12 //y=1.505 //x2=34.12 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=34.12 //y=0.625 //x2=34.12 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=34.12 //y=0.625 //x2=34.12 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=33.235 //y=1.59 //x2=33.15 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=33.235 //y=1.59 //x2=33.635 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=34.035 //y=1.59 //x2=34.12 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=34.035 //y=1.59 //x2=33.635 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=33.15 //y=1.505 //x2=33.15 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=33.15 //y=1.505 //x2=33.15 //y2=0.89
ends PM_TMRDFFSNQX1\%noxref_39

subckt PM_TMRDFFSNQX1\%noxref_40 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=35.525 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=34.42 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=35.66 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=36.63 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=36.545 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=35.66 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=35.575 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=36.63 //y=0.625 //x2=36.63 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=36.63 //y=0.625 //x2=36.63 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=35.745 //y=0.54 //x2=35.66 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=35.745 //y=0.54 //x2=36.145 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=36.545 //y=0.54 //x2=36.63 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=36.545 //y=0.54 //x2=36.145 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=35.66 //y=1.08 //x2=35.66 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=35.66 //y=1.08 //x2=35.66 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=35.66 //y=0.91 //x2=35.66 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=35.66 //y=0.91 //x2=35.66 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=35.66 //y=0.625 //x2=35.66 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=35.66 //y=0.625 //x2=35.66 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=34.695 //y=0.995 //x2=34.61 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=35.575 //y=0.995 //x2=35.66 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=35.575 //y=0.995 //x2=34.695 //y2=0.995
ends PM_TMRDFFSNQX1\%noxref_40

subckt PM_TMRDFFSNQX1\%noxref_41 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632682f //x=37.93 //y=0.365
c52 ( 17 0 ) capacitor c=0.00722223f //x=40.005 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=39.92 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=39.035 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=39.035 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=38.95 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=38.065 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=40.005 //y=0.615 //x2=40.005 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=40.005 //y=0.615 //x2=40.005 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=39.12 //y=0.53 //x2=39.035 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=39.12 //y=0.53 //x2=39.52 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=39.92 //y=0.53 //x2=40.005 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=39.92 //y=0.53 //x2=39.52 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=39.035 //y=1.495 //x2=39.035 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=39.035 //y=1.495 //x2=39.035 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=39.035 //y=0.615 //x2=39.035 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=39.035 //y=0.615 //x2=39.035 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=38.15 //y=1.58 //x2=38.065 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=38.15 //y=1.58 //x2=38.55 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=38.95 //y=1.58 //x2=39.035 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=38.95 //y=1.58 //x2=38.55 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=38.065 //y=1.495 //x2=38.065 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=38.065 //y=1.495 //x2=38.065 //y2=0.88
ends PM_TMRDFFSNQX1\%noxref_41

subckt PM_TMRDFFSNQX1\%noxref_42 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.063352f //x=41.26 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=43.335 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=43.25 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=42.365 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=42.365 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=42.28 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=41.395 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=43.335 //y=0.615 //x2=43.335 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=43.335 //y=0.615 //x2=43.335 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=42.45 //y=0.53 //x2=42.365 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=42.45 //y=0.53 //x2=42.85 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=43.25 //y=0.53 //x2=43.335 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=43.25 //y=0.53 //x2=42.85 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=42.365 //y=1.495 //x2=42.365 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=42.365 //y=1.495 //x2=42.365 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=42.365 //y=0.615 //x2=42.365 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=42.365 //y=0.615 //x2=42.365 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=41.48 //y=1.58 //x2=41.395 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=41.48 //y=1.58 //x2=41.88 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=42.28 //y=1.58 //x2=42.365 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=42.28 //y=1.58 //x2=41.88 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=41.395 //y=1.495 //x2=41.395 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=41.395 //y=1.495 //x2=41.395 //y2=0.88
ends PM_TMRDFFSNQX1\%noxref_42

subckt PM_TMRDFFSNQX1\%noxref_43 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=44.485 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=46.475 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=46.475 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=45.59 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=45.505 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=44.62 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=45.675 //y=1.59 //x2=45.59 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.675 //y=1.59 //x2=46.075 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.475 //y=1.59 //x2=46.56 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=46.475 //y=1.59 //x2=46.075 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=45.675 //y=0.54 //x2=45.59 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.675 //y=0.54 //x2=46.075 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.475 //y=0.54 //x2=46.56 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=46.475 //y=0.54 //x2=46.075 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=45.59 //y=1.505 //x2=45.59 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=45.59 //y=1.505 //x2=45.59 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=45.59 //y=0.625 //x2=45.59 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=45.59 //y=0.625 //x2=45.59 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=44.705 //y=1.59 //x2=44.62 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=44.705 //y=1.59 //x2=45.105 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=45.505 //y=1.59 //x2=45.59 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=45.505 //y=1.59 //x2=45.105 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=44.62 //y=1.505 //x2=44.62 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=44.62 //y=1.505 //x2=44.62 //y2=0.89
ends PM_TMRDFFSNQX1\%noxref_43

subckt PM_TMRDFFSNQX1\%noxref_44 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=46.995 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=45.89 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=47.13 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=48.1 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=48.015 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=47.13 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=47.045 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=48.1 //y=0.625 //x2=48.1 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=48.1 //y=0.625 //x2=48.1 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=47.215 //y=0.54 //x2=47.13 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=47.215 //y=0.54 //x2=47.615 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=48.015 //y=0.54 //x2=48.1 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=48.015 //y=0.54 //x2=47.615 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=47.13 //y=1.08 //x2=47.13 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=47.13 //y=1.08 //x2=47.13 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=47.13 //y=0.91 //x2=47.13 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=47.13 //y=0.91 //x2=47.13 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=47.13 //y=0.625 //x2=47.13 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=47.13 //y=0.625 //x2=47.13 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=46.165 //y=0.995 //x2=46.08 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=47.045 //y=0.995 //x2=47.13 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=47.045 //y=0.995 //x2=46.165 //y2=0.995
ends PM_TMRDFFSNQX1\%noxref_44

subckt PM_TMRDFFSNQX1\%noxref_45 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0633518f //x=49.4 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=51.475 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=51.39 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=50.505 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=50.505 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=50.42 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=49.535 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=51.475 //y=0.615 //x2=51.475 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=51.475 //y=0.615 //x2=51.475 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=50.59 //y=0.53 //x2=50.505 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=50.59 //y=0.53 //x2=50.99 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=51.39 //y=0.53 //x2=51.475 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=51.39 //y=0.53 //x2=50.99 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=50.505 //y=1.495 //x2=50.505 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=50.505 //y=1.495 //x2=50.505 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=50.505 //y=0.615 //x2=50.505 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=50.505 //y=0.615 //x2=50.505 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=49.62 //y=1.58 //x2=49.535 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=49.62 //y=1.58 //x2=50.02 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=50.42 //y=1.58 //x2=50.505 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=50.42 //y=1.58 //x2=50.02 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=49.535 //y=1.495 //x2=49.535 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=49.535 //y=1.495 //x2=49.535 //y2=0.88
ends PM_TMRDFFSNQX1\%noxref_45

subckt PM_TMRDFFSNQX1\%noxref_46 ( 1 5 9 13 17 35 )
c49 ( 35 0 ) capacitor c=0.0673195f //x=52.625 //y=0.375
c50 ( 17 0 ) capacitor c=0.0178317f //x=54.615 //y=1.59
c51 ( 13 0 ) capacitor c=0.0154936f //x=54.615 //y=0.54
c52 ( 9 0 ) capacitor c=0.00678203f //x=53.73 //y=0.625
c53 ( 5 0 ) capacitor c=0.0164013f //x=53.645 //y=1.59
c54 ( 1 0 ) capacitor c=0.00696517f //x=52.76 //y=1.505
r55 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=53.815 //y=1.59 //x2=53.73 //y2=1.63
r56 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=53.815 //y=1.59 //x2=54.215 //y2=1.59
r57 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.615 //y=1.59 //x2=54.7 //y2=1.59
r58 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.615 //y=1.59 //x2=54.215 //y2=1.59
r59 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=53.815 //y=0.54 //x2=53.73 //y2=0.5
r60 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=53.815 //y=0.54 //x2=54.215 //y2=0.54
r61 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.615 //y=0.54 //x2=54.7 //y2=0.54
r62 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=54.615 //y=0.54 //x2=54.215 //y2=0.54
r63 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=53.73 //y=1.505 //x2=53.73 //y2=1.63
r64 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=53.73 //y=1.505 //x2=53.73 //y2=0.89
r65 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=53.73 //y=0.625 //x2=53.73 //y2=0.5
r66 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=53.73 //y=0.625 //x2=53.73 //y2=0.89
r67 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=52.845 //y=1.59 //x2=52.76 //y2=1.63
r68 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=52.845 //y=1.59 //x2=53.245 //y2=1.59
r69 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=53.645 //y=1.59 //x2=53.73 //y2=1.63
r70 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=53.645 //y=1.59 //x2=53.245 //y2=1.59
r71 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=52.76 //y=1.505 //x2=52.76 //y2=1.63
r72 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=52.76 //y=1.505 //x2=52.76 //y2=0.89
ends PM_TMRDFFSNQX1\%noxref_46

subckt PM_TMRDFFSNQX1\%noxref_47 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414739f //x=55.135 //y=0.375
c53 ( 28 0 ) capacitor c=0.0045748f //x=54.03 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=55.27 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=56.24 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=56.155 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=55.27 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218888f //x=55.185 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=56.24 //y=0.625 //x2=56.24 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=56.24 //y=0.625 //x2=56.24 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=55.355 //y=0.54 //x2=55.27 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=55.355 //y=0.54 //x2=55.755 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=56.155 //y=0.54 //x2=56.24 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=56.155 //y=0.54 //x2=55.755 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=55.27 //y=1.08 //x2=55.27 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=55.27 //y=1.08 //x2=55.27 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=55.27 //y=0.91 //x2=55.27 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=55.27 //y=0.91 //x2=55.27 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=55.27 //y=0.625 //x2=55.27 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=55.27 //y=0.625 //x2=55.27 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=54.305 //y=0.995 //x2=54.22 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=55.185 //y=0.995 //x2=55.27 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=55.185 //y=0.995 //x2=54.305 //y2=0.995
ends PM_TMRDFFSNQX1\%noxref_47

subckt PM_TMRDFFSNQX1\%noxref_48 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0673029f //x=57.435 //y=0.375
c53 ( 17 0 ) capacitor c=0.0178286f //x=59.425 //y=1.59
c54 ( 13 0 ) capacitor c=0.0154917f //x=59.425 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=58.54 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=58.455 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=57.57 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=58.625 //y=1.59 //x2=58.54 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=58.625 //y=1.59 //x2=59.025 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.425 //y=1.59 //x2=59.51 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.425 //y=1.59 //x2=59.025 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=58.625 //y=0.54 //x2=58.54 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=58.625 //y=0.54 //x2=59.025 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.425 //y=0.54 //x2=59.51 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=59.425 //y=0.54 //x2=59.025 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=58.54 //y=1.505 //x2=58.54 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=58.54 //y=1.505 //x2=58.54 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=58.54 //y=0.625 //x2=58.54 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=58.54 //y=0.625 //x2=58.54 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=57.655 //y=1.59 //x2=57.57 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=57.655 //y=1.59 //x2=58.055 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=58.455 //y=1.59 //x2=58.54 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=58.455 //y=1.59 //x2=58.055 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=57.57 //y=1.505 //x2=57.57 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=57.57 //y=1.505 //x2=57.57 //y2=0.89
ends PM_TMRDFFSNQX1\%noxref_48

subckt PM_TMRDFFSNQX1\%noxref_49 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0414744f //x=59.945 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=58.84 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=60.08 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=61.05 //y=0.625
c56 ( 11 0 ) capacitor c=0.0144274f //x=60.965 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=60.08 //y=0.625
c58 ( 1 0 ) capacitor c=0.0218873f //x=59.995 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=61.05 //y=0.625 //x2=61.05 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=61.05 //y=0.625 //x2=61.05 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=60.165 //y=0.54 //x2=60.08 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=60.165 //y=0.54 //x2=60.565 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=60.965 //y=0.54 //x2=61.05 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=60.965 //y=0.54 //x2=60.565 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=60.08 //y=1.08 //x2=60.08 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=60.08 //y=1.08 //x2=60.08 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=60.08 //y=0.91 //x2=60.08 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=60.08 //y=0.91 //x2=60.08 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=60.08 //y=0.625 //x2=60.08 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=60.08 //y=0.625 //x2=60.08 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=59.115 //y=0.995 //x2=59.03 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=59.995 //y=0.995 //x2=60.08 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=59.995 //y=0.995 //x2=59.115 //y2=0.995
ends PM_TMRDFFSNQX1\%noxref_49

subckt PM_TMRDFFSNQX1\%noxref_50 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632682f //x=62.35 //y=0.365
c52 ( 17 0 ) capacitor c=0.00722223f //x=64.425 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=64.34 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=63.455 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=63.455 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=63.37 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=62.485 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=64.425 //y=0.615 //x2=64.425 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=64.425 //y=0.615 //x2=64.425 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=63.54 //y=0.53 //x2=63.455 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=63.54 //y=0.53 //x2=63.94 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=64.34 //y=0.53 //x2=64.425 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=64.34 //y=0.53 //x2=63.94 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=63.455 //y=1.495 //x2=63.455 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=63.455 //y=1.495 //x2=63.455 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=63.455 //y=0.615 //x2=63.455 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=63.455 //y=0.615 //x2=63.455 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=62.57 //y=1.58 //x2=62.485 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=62.57 //y=1.58 //x2=62.97 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=63.37 //y=1.58 //x2=63.455 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=63.37 //y=1.58 //x2=62.97 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=62.485 //y=1.495 //x2=62.485 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=62.485 //y=1.495 //x2=62.485 //y2=0.88
ends PM_TMRDFFSNQX1\%noxref_50

subckt PM_TMRDFFSNQX1\%noxref_51 ( 1 5 9 10 13 17 29 )
c51 ( 29 0 ) capacitor c=0.0632684f //x=65.68 //y=0.365
c52 ( 17 0 ) capacitor c=0.0072343f //x=67.755 //y=0.615
c53 ( 13 0 ) capacitor c=0.0145084f //x=67.67 //y=0.53
c54 ( 10 0 ) capacitor c=0.00582081f //x=66.785 //y=1.495
c55 ( 9 0 ) capacitor c=0.006761f //x=66.785 //y=0.615
c56 ( 5 0 ) capacitor c=0.0173046f //x=66.7 //y=1.58
c57 ( 1 0 ) capacitor c=0.00733328f //x=65.815 //y=1.495
r58 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=67.755 //y=0.615 //x2=67.755 //y2=0.49
r59 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=67.755 //y=0.615 //x2=67.755 //y2=0.88
r60 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=66.87 //y=0.53 //x2=66.785 //y2=0.49
r61 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=66.87 //y=0.53 //x2=67.27 //y2=0.53
r62 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=67.67 //y=0.53 //x2=67.755 //y2=0.49
r63 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=67.67 //y=0.53 //x2=67.27 //y2=0.53
r64 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=66.785 //y=1.495 //x2=66.785 //y2=1.62
r65 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=66.785 //y=1.495 //x2=66.785 //y2=0.88
r66 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=66.785 //y=0.615 //x2=66.785 //y2=0.49
r67 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=66.785 //y=0.615 //x2=66.785 //y2=0.88
r68 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=65.9 //y=1.58 //x2=65.815 //y2=1.62
r69 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=65.9 //y=1.58 //x2=66.3 //y2=1.58
r70 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=66.7 //y=1.58 //x2=66.785 //y2=1.62
r71 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=66.7 //y=1.58 //x2=66.3 //y2=1.58
r72 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=65.815 //y=1.495 //x2=65.815 //y2=1.62
r73 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=65.815 //y=1.495 //x2=65.815 //y2=0.88
ends PM_TMRDFFSNQX1\%noxref_51

subckt PM_TMRDFFSNQX1\%noxref_52 ( 1 5 9 13 17 35 )
c51 ( 35 0 ) capacitor c=0.0680259f //x=68.905 //y=0.375
c52 ( 17 0 ) capacitor c=0.0180446f //x=70.895 //y=1.59
c53 ( 13 0 ) capacitor c=0.0155283f //x=70.895 //y=0.54
c54 ( 9 0 ) capacitor c=0.00678203f //x=70.01 //y=0.625
c55 ( 5 0 ) capacitor c=0.0164013f //x=69.925 //y=1.59
c56 ( 1 0 ) capacitor c=0.00696517f //x=69.04 //y=1.505
r57 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=70.095 //y=1.59 //x2=70.01 //y2=1.63
r58 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=70.095 //y=1.59 //x2=70.495 //y2=1.59
r59 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.895 //y=1.59 //x2=70.98 //y2=1.59
r60 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=70.895 //y=1.59 //x2=70.495 //y2=1.59
r61 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=70.095 //y=0.54 //x2=70.01 //y2=0.5
r62 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=70.095 //y=0.54 //x2=70.495 //y2=0.54
r63 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.895 //y=0.54 //x2=70.98 //y2=0.54
r64 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=70.895 //y=0.54 //x2=70.495 //y2=0.54
r65 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=70.01 //y=1.505 //x2=70.01 //y2=1.63
r66 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=70.01 //y=1.505 //x2=70.01 //y2=0.89
r67 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=70.01 //y=0.625 //x2=70.01 //y2=0.5
r68 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=70.01 //y=0.625 //x2=70.01 //y2=0.89
r69 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=69.125 //y=1.59 //x2=69.04 //y2=1.63
r70 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=69.125 //y=1.59 //x2=69.525 //y2=1.59
r71 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=69.925 //y=1.59 //x2=70.01 //y2=1.63
r72 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=69.925 //y=1.59 //x2=69.525 //y2=1.59
r73 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=69.04 //y=1.505 //x2=69.04 //y2=1.63
r74 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=69.04 //y=1.505 //x2=69.04 //y2=0.89
ends PM_TMRDFFSNQX1\%noxref_52

subckt PM_TMRDFFSNQX1\%noxref_53 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.042068f //x=71.415 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=70.31 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=71.55 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=72.52 //y=0.625
c56 ( 11 0 ) capacitor c=0.014695f //x=72.435 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=71.55 //y=0.625
c58 ( 1 0 ) capacitor c=0.0234159f //x=71.465 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=72.52 //y=0.625 //x2=72.52 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=72.52 //y=0.625 //x2=72.52 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=71.635 //y=0.54 //x2=71.55 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=71.635 //y=0.54 //x2=72.035 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=72.435 //y=0.54 //x2=72.52 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=72.435 //y=0.54 //x2=72.035 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=71.55 //y=1.08 //x2=71.55 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=71.55 //y=1.08 //x2=71.55 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=71.55 //y=0.91 //x2=71.55 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=71.55 //y=0.91 //x2=71.55 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=71.55 //y=0.625 //x2=71.55 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=71.55 //y=0.625 //x2=71.55 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=70.585 //y=0.995 //x2=70.5 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=71.465 //y=0.995 //x2=71.55 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=71.465 //y=0.995 //x2=70.585 //y2=0.995
ends PM_TMRDFFSNQX1\%noxref_53

subckt PM_TMRDFFSNQX1\%noxref_54 ( 1 5 9 10 13 17 29 )
c57 ( 29 0 ) capacitor c=0.0761166f //x=73.82 //y=0.365
c58 ( 17 0 ) capacitor c=0.0072249f //x=75.895 //y=0.615
c59 ( 13 0 ) capacitor c=0.0154142f //x=75.81 //y=0.53
c60 ( 10 0 ) capacitor c=0.00754234f //x=74.925 //y=1.495
c61 ( 9 0 ) capacitor c=0.006761f //x=74.925 //y=0.615
c62 ( 5 0 ) capacitor c=0.0213241f //x=74.84 //y=1.58
c63 ( 1 0 ) capacitor c=0.00492513f //x=73.955 //y=1.495
r64 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=75.895 //y=0.615 //x2=75.895 //y2=0.49
r65 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=75.895 //y=0.615 //x2=75.895 //y2=1.22
r66 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=75.01 //y=0.53 //x2=74.925 //y2=0.49
r67 (  14 29 ) resistor r=27.0374 //w=0.187 //l=0.395 //layer=li \
 //thickness=0.1 //x=75.01 //y=0.53 //x2=75.405 //y2=0.53
r68 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=75.81 //y=0.53 //x2=75.895 //y2=0.49
r69 (  13 29 ) resistor r=27.7219 //w=0.187 //l=0.405 //layer=li \
 //thickness=0.1 //x=75.81 //y=0.53 //x2=75.405 //y2=0.53
r70 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=74.925 //y=1.495 //x2=74.925 //y2=1.62
r71 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=74.925 //y=1.495 //x2=74.925 //y2=0.88
r72 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=74.925 //y=0.615 //x2=74.925 //y2=0.49
r73 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=74.925 //y=0.615 //x2=74.925 //y2=0.88
r74 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=74.04 //y=1.58 //x2=73.955 //y2=1.62
r75 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=74.04 //y=1.58 //x2=74.44 //y2=1.58
r76 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=74.84 //y=1.58 //x2=74.925 //y2=1.62
r77 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=74.84 //y=1.58 //x2=74.44 //y2=1.58
r78 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=73.955 //y=1.495 //x2=73.955 //y2=1.62
r79 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=73.955 //y=1.495 //x2=73.955 //y2=0.88
ends PM_TMRDFFSNQX1\%noxref_54

subckt PM_TMRDFFSNQX1\%noxref_55 ( 1 5 9 10 13 17 29 )
c55 ( 29 0 ) capacitor c=0.0723103f //x=77.15 //y=0.365
c56 ( 17 0 ) capacitor c=0.0072249f //x=79.225 //y=0.615
c57 ( 13 0 ) capacitor c=0.0155051f //x=79.14 //y=0.53
c58 ( 10 0 ) capacitor c=0.00907139f //x=78.255 //y=1.495
c59 ( 9 0 ) capacitor c=0.006761f //x=78.255 //y=0.615
c60 ( 5 0 ) capacitor c=0.019003f //x=78.17 //y=1.58
c61 ( 1 0 ) capacitor c=0.00885385f //x=77.285 //y=1.495
r62 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=79.225 //y=0.615 //x2=79.225 //y2=0.49
r63 (  17 29 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=79.225 //y=0.615 //x2=79.225 //y2=1.22
r64 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.34 //y=0.53 //x2=78.255 //y2=0.49
r65 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=78.34 //y=0.53 //x2=78.74 //y2=0.53
r66 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=79.14 //y=0.53 //x2=79.225 //y2=0.49
r67 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=79.14 //y=0.53 //x2=78.74 //y2=0.53
r68 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=78.255 //y=1.495 //x2=78.255 //y2=1.62
r69 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=78.255 //y=1.495 //x2=78.255 //y2=0.88
r70 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=78.255 //y=0.615 //x2=78.255 //y2=0.49
r71 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=78.255 //y=0.615 //x2=78.255 //y2=0.88
r72 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=77.37 //y=1.58 //x2=77.285 //y2=1.62
r73 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=77.37 //y=1.58 //x2=77.77 //y2=1.58
r74 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=78.17 //y=1.58 //x2=78.255 //y2=1.62
r75 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=78.17 //y=1.58 //x2=77.77 //y2=1.58
r76 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=77.285 //y=1.495 //x2=77.285 //y2=1.62
r77 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=77.285 //y=1.495 //x2=77.285 //y2=0.88
ends PM_TMRDFFSNQX1\%noxref_55

subckt PM_TMRDFFSNQX1\%noxref_56 ( 1 5 9 10 13 17 29 )
c56 ( 29 0 ) capacitor c=0.0637832f //x=80.48 //y=0.365
c57 ( 17 0 ) capacitor c=0.00722228f //x=82.555 //y=0.615
c58 ( 13 0 ) capacitor c=0.0141607f //x=82.47 //y=0.53
c59 ( 10 0 ) capacitor c=0.00712138f //x=81.585 //y=1.495
c60 ( 9 0 ) capacitor c=0.006761f //x=81.585 //y=0.615
c61 ( 5 0 ) capacitor c=0.0233454f //x=81.5 //y=1.58
c62 ( 1 0 ) capacitor c=0.00481264f //x=80.615 //y=1.495
r63 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=82.555 //y=0.615 //x2=82.555 //y2=0.49
r64 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=82.555 //y=0.615 //x2=82.555 //y2=0.88
r65 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=81.67 //y=0.53 //x2=81.585 //y2=0.49
r66 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=81.67 //y=0.53 //x2=82.07 //y2=0.53
r67 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=82.47 //y=0.53 //x2=82.555 //y2=0.49
r68 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=82.47 //y=0.53 //x2=82.07 //y2=0.53
r69 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=81.585 //y=1.495 //x2=81.585 //y2=1.62
r70 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=81.585 //y=1.495 //x2=81.585 //y2=0.88
r71 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=81.585 //y=0.615 //x2=81.585 //y2=0.49
r72 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=81.585 //y=0.615 //x2=81.585 //y2=0.88
r73 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=80.7 //y=1.58 //x2=80.615 //y2=1.62
r74 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=80.7 //y=1.58 //x2=81.1 //y2=1.58
r75 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=81.5 //y=1.58 //x2=81.585 //y2=1.62
r76 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=81.5 //y=1.58 //x2=81.1 //y2=1.58
r77 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=80.615 //y=1.495 //x2=80.615 //y2=1.62
r78 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=80.615 //y=1.495 //x2=80.615 //y2=0.88
ends PM_TMRDFFSNQX1\%noxref_56

subckt PM_TMRDFFSNQX1\%Q ( 1 2 3 4 5 6 7 18 19 20 21 31 33 )
c44 ( 33 0 ) capacitor c=0.028734f //x=84.22 //y=5.02
c45 ( 31 0 ) capacitor c=0.0172744f //x=84.175 //y=0.91
c46 ( 21 0 ) capacitor c=0.00575887f //x=84.45 //y=4.58
c47 ( 20 0 ) capacitor c=0.0136889f //x=84.645 //y=4.58
c48 ( 19 0 ) capacitor c=0.00636159f //x=84.445 //y=2.08
c49 ( 18 0 ) capacitor c=0.0140707f //x=84.645 //y=2.08
c50 ( 1 0 ) capacitor c=0.105613f //x=84.73 //y=2.22
r51 (  20 23 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=84.645 //y=4.58 //x2=84.73 //y2=4.495
r52 (  20 21 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=84.645 //y=4.58 //x2=84.45 //y2=4.58
r53 (  18 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=84.645 //y=2.08 //x2=84.73 //y2=2.165
r54 (  18 19 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=84.645 //y=2.08 //x2=84.445 //y2=2.08
r55 (  12 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=84.365 //y=4.665 //x2=84.45 //y2=4.58
r56 (  12 33 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=84.365 //y=4.665 //x2=84.365 //y2=5.725
r57 (  8 19 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=84.36 //y=1.995 //x2=84.445 //y2=2.08
r58 (  8 31 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=84.36 //y=1.995 //x2=84.36 //y2=1.005
r59 (  7 23 ) resistor r=3.76471 //w=0.187 //l=0.055 //layer=li \
 //thickness=0.1 //x=84.73 //y=4.44 //x2=84.73 //y2=4.495
r60 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=84.73 //y=4.07 //x2=84.73 //y2=4.44
r61 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=84.73 //y=3.7 //x2=84.73 //y2=4.07
r62 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=84.73 //y=3.33 //x2=84.73 //y2=3.7
r63 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=84.73 //y=2.96 //x2=84.73 //y2=3.33
r64 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=84.73 //y=2.59 //x2=84.73 //y2=2.96
r65 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=84.73 //y=2.22 //x2=84.73 //y2=2.59
r66 (  1 22 ) resistor r=3.76471 //w=0.187 //l=0.055 //layer=li \
 //thickness=0.1 //x=84.73 //y=2.22 //x2=84.73 //y2=2.165
ends PM_TMRDFFSNQX1\%Q

