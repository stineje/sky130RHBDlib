magic
tech sky130A
magscale 1 2
timestamp 1669564312
<< nwell >>
rect -87 786 531 1550
<< pwell >>
rect -34 -34 34 544
rect 57 -17 91 17
rect 410 -34 478 544
<< nmos >>
rect 155 296 185 349
tri 185 296 201 312 sw
rect 155 266 261 296
tri 261 266 291 296 sw
rect 155 165 185 266
tri 185 250 201 266 nw
tri 245 250 261 266 ne
tri 185 165 201 181 sw
tri 245 165 261 181 se
rect 261 165 291 266
tri 155 135 185 165 ne
rect 185 135 261 165
tri 261 135 291 165 nw
<< pmos >>
rect 163 1004 193 1404
rect 251 1004 281 1404
<< ndiff >>
rect 99 333 155 349
rect 99 299 109 333
rect 143 299 155 333
rect 99 261 155 299
rect 185 333 345 349
rect 185 312 303 333
tri 185 296 201 312 ne
rect 201 299 303 312
rect 337 299 345 333
rect 201 296 345 299
tri 261 266 291 296 ne
rect 99 227 109 261
rect 143 227 155 261
rect 99 193 155 227
rect 99 159 109 193
rect 143 159 155 193
tri 185 250 201 266 se
rect 201 250 245 266
tri 245 250 261 266 sw
rect 185 217 261 250
rect 185 183 205 217
rect 239 183 261 217
rect 185 181 261 183
tri 185 165 201 181 ne
rect 201 165 245 181
tri 245 165 261 181 nw
rect 291 261 345 296
rect 291 227 303 261
rect 337 227 345 261
rect 291 193 345 227
rect 99 135 155 159
tri 155 135 185 165 sw
tri 261 135 291 165 se
rect 291 159 303 193
rect 337 159 345 193
rect 291 135 345 159
rect 99 123 345 135
rect 99 89 109 123
rect 143 89 205 123
rect 239 89 303 123
rect 337 89 345 123
rect 99 73 345 89
<< pdiff >>
rect 107 1366 163 1404
rect 107 1332 117 1366
rect 151 1332 163 1366
rect 107 1298 163 1332
rect 107 1264 117 1298
rect 151 1264 163 1298
rect 107 1230 163 1264
rect 107 1196 117 1230
rect 151 1196 163 1230
rect 107 1162 163 1196
rect 107 1128 117 1162
rect 151 1128 163 1162
rect 107 1094 163 1128
rect 107 1060 117 1094
rect 151 1060 163 1094
rect 107 1004 163 1060
rect 193 1366 251 1404
rect 193 1332 205 1366
rect 239 1332 251 1366
rect 193 1298 251 1332
rect 193 1264 205 1298
rect 239 1264 251 1298
rect 193 1230 251 1264
rect 193 1196 205 1230
rect 239 1196 251 1230
rect 193 1162 251 1196
rect 193 1128 205 1162
rect 239 1128 251 1162
rect 193 1094 251 1128
rect 193 1060 205 1094
rect 239 1060 251 1094
rect 193 1004 251 1060
rect 281 1366 335 1404
rect 281 1332 293 1366
rect 327 1332 335 1366
rect 281 1298 335 1332
rect 281 1264 293 1298
rect 327 1264 335 1298
rect 281 1230 335 1264
rect 281 1196 293 1230
rect 327 1196 335 1230
rect 281 1162 335 1196
rect 281 1128 293 1162
rect 327 1128 335 1162
rect 281 1094 335 1128
rect 281 1060 293 1094
rect 327 1060 335 1094
rect 281 1004 335 1060
<< ndiffc >>
rect 109 299 143 333
rect 303 299 337 333
rect 109 227 143 261
rect 109 159 143 193
rect 205 183 239 217
rect 303 227 337 261
rect 303 159 337 193
rect 109 89 143 123
rect 205 89 239 123
rect 303 89 337 123
<< pdiffc >>
rect 117 1332 151 1366
rect 117 1264 151 1298
rect 117 1196 151 1230
rect 117 1128 151 1162
rect 117 1060 151 1094
rect 205 1332 239 1366
rect 205 1264 239 1298
rect 205 1196 239 1230
rect 205 1128 239 1162
rect 205 1060 239 1094
rect 293 1332 327 1366
rect 293 1264 327 1298
rect 293 1196 327 1230
rect 293 1128 327 1162
rect 293 1060 327 1094
<< psubdiff >>
rect -34 482 478 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 410 461 478 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 410 427 427 461
rect 461 427 478 461
rect -34 313 34 353
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 410 313 478 353
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect -34 17 34 57
rect 410 57 427 91
rect 461 57 478 91
rect 410 17 478 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 478 17
rect -34 -34 478 -17
<< nsubdiff >>
rect -34 1497 478 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 478 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 410 1423 478 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 410 979 478 1019
rect 410 945 427 979
rect 461 945 478 979
rect -34 871 -17 905
rect 17 884 34 905
rect 410 905 478 945
rect 410 884 427 905
rect 17 871 427 884
rect 461 871 478 905
rect -34 822 478 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 427 427 461 461
rect 427 353 461 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 427 279 461 313
rect 427 205 461 239
rect 427 131 461 165
rect 427 57 461 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 427 1389 461 1423
rect 427 1315 461 1349
rect 427 1241 461 1275
rect 427 1167 461 1201
rect 427 1093 461 1127
rect 427 1019 461 1053
rect -17 945 17 979
rect 427 945 461 979
rect -17 871 17 905
rect 427 871 461 905
<< poly >>
rect 163 1404 193 1430
rect 251 1404 281 1430
rect 163 973 193 1004
rect 251 973 281 1004
rect 121 957 281 973
rect 121 923 131 957
rect 165 943 281 957
rect 165 923 175 943
rect 121 907 175 923
rect 121 433 175 449
rect 121 399 131 433
rect 165 413 175 433
rect 165 399 185 413
rect 121 383 185 399
rect 155 349 185 383
<< polycont >>
rect 131 923 165 957
rect 131 399 165 433
<< locali >>
rect -34 1497 478 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 478 1497
rect -34 1446 478 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 117 1366 151 1446
rect 117 1298 151 1332
rect 117 1230 151 1264
rect 117 1162 151 1196
rect 117 1094 151 1128
rect 117 1016 151 1060
rect 205 1366 239 1404
rect 205 1298 239 1332
rect 205 1230 239 1264
rect 205 1162 239 1196
rect 205 1094 239 1128
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 131 957 165 973
rect 205 957 239 1060
rect 293 1366 327 1446
rect 293 1298 327 1332
rect 293 1230 327 1264
rect 293 1162 327 1196
rect 293 1094 327 1128
rect 293 1016 327 1060
rect 410 1423 478 1446
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect 165 923 239 957
rect 410 979 478 1019
rect 410 945 427 979
rect 461 945 478 979
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 131 433 165 923
rect 410 905 478 945
rect 410 871 427 905
rect 461 871 478 905
rect 410 822 478 871
rect 131 383 165 399
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect -34 34 34 57
rect 109 333 143 349
rect 109 261 143 299
rect 109 193 143 227
rect 205 217 239 609
rect 410 461 478 544
rect 410 427 427 461
rect 461 427 478 461
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect 205 167 239 183
rect 303 333 337 349
rect 303 261 337 299
rect 303 193 337 227
rect 109 123 143 159
rect 303 123 337 159
rect 143 89 205 123
rect 239 89 303 123
rect 109 34 143 89
rect 205 34 239 89
rect 303 34 337 89
rect 410 313 478 353
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect 410 57 427 91
rect 461 57 478 91
rect 410 34 478 57
rect -34 17 478 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 478 17
rect -34 -34 478 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
<< metal1 >>
rect -34 1497 478 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 478 1497
rect -34 1446 478 1463
rect -34 17 478 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 478 17
rect -34 -34 478 -17
<< labels >>
rlabel metal1 205 575 239 609 1 YN
port 1 n
rlabel metal1 205 501 239 535 1 YN
port 2 n
rlabel metal1 205 427 239 461 1 YN
port 3 n
rlabel metal1 -34 1446 478 1514 1 VPWR
port 4 n
rlabel metal1 -34 -34 478 34 1 VGND
port 5 n
rlabel nwell 57 1463 91 1497 1 VPB
port 6 n
rlabel pwell 57 -17 91 17 1 VNB
port 7 n
<< end >>
