* SPICE3 file created from TMRDFFSNRNQX1.ext - technology: sky130A

.subckt TMRDFFSNRNQX1 Q D CLK SN RN VDD GND
X0 GND D dffsnrnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X1 dffsnrnx1_pcell_0/m1_831_501# dffsnrnx1_pcell_0/m1_716_649# dffsnrnx1_pcell_0/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X2 dffsnrnx1_pcell_0/nand3x1_pcell_0/li_393_182# RN dffsnrnx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X3 VDD D dffsnrnx1_pcell_0/m1_831_501# VDD pshort w=2 l=0.15
X4 VDD RN dffsnrnx1_pcell_0/m1_831_501# VDD pshort w=2 l=0.15
X5 VDD dffsnrnx1_pcell_0/m1_716_649# dffsnrnx1_pcell_0/m1_831_501# VDD pshort w=2 l=0.15
X6 GND dffsnrnx1_pcell_0/m1_831_501# dffsnrnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X7 dffsnrnx1_pcell_0/m1_716_649# dffsnrnx1_pcell_0/m1_1660_723# dffsnrnx1_pcell_0/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X8 dffsnrnx1_pcell_0/nand3x1_pcell_1/li_393_182# CLK dffsnrnx1_pcell_0/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X9 VDD dffsnrnx1_pcell_0/m1_831_501# dffsnrnx1_pcell_0/m1_716_649# VDD pshort w=2 l=0.15
X10 VDD CLK dffsnrnx1_pcell_0/m1_716_649# VDD pshort w=2 l=0.15
X11 VDD dffsnrnx1_pcell_0/m1_1660_723# dffsnrnx1_pcell_0/m1_716_649# VDD pshort w=2 l=0.15
X12 GND dffsnrnx1_pcell_0/m1_831_501# dffsnrnx1_pcell_0/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X13 dffsnrnx1_pcell_0/m1_2757_501# dffsnrnx1_pcell_0/m1_1660_723# dffsnrnx1_pcell_0/nand3x1_pcell_2/li_393_182# GND nshort w=3 l=0.15
X14 dffsnrnx1_pcell_0/nand3x1_pcell_2/li_393_182# SN dffsnrnx1_pcell_0/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X15 VDD dffsnrnx1_pcell_0/m1_831_501# dffsnrnx1_pcell_0/m1_2757_501# VDD pshort w=2 l=0.15
X16 VDD SN dffsnrnx1_pcell_0/m1_2757_501# VDD pshort w=2 l=0.15
X17 VDD dffsnrnx1_pcell_0/m1_1660_723# dffsnrnx1_pcell_0/m1_2757_501# VDD pshort w=2 l=0.15
X18 GND dffsnrnx1_pcell_0/m1_2757_501# dffsnrnx1_pcell_0/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X19 dffsnrnx1_pcell_0/m1_1660_723# RN dffsnrnx1_pcell_0/nand3x1_pcell_3/li_393_182# GND nshort w=3 l=0.15
X20 dffsnrnx1_pcell_0/nand3x1_pcell_3/li_393_182# CLK dffsnrnx1_pcell_0/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X21 VDD dffsnrnx1_pcell_0/m1_2757_501# dffsnrnx1_pcell_0/m1_1660_723# VDD pshort w=2 l=0.15
X22 VDD CLK dffsnrnx1_pcell_0/m1_1660_723# VDD pshort w=2 l=0.15
X23 VDD RN dffsnrnx1_pcell_0/m1_1660_723# VDD pshort w=2 l=0.15
X24 GND dffsnrnx1_pcell_0/m1_716_649# dffsnrnx1_pcell_0/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X25 m1_4715_501# m1_5643_945# dffsnrnx1_pcell_0/nand3x1_pcell_4/li_393_182# GND nshort w=3 l=0.15
X26 dffsnrnx1_pcell_0/nand3x1_pcell_4/li_393_182# RN dffsnrnx1_pcell_0/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X27 VDD dffsnrnx1_pcell_0/m1_716_649# m1_4715_501# VDD pshort w=2 l=0.15
X28 VDD RN m1_4715_501# VDD pshort w=2 l=0.15
X29 VDD m1_5643_945# m1_4715_501# VDD pshort w=2 l=0.15
X30 GND m1_4715_501# dffsnrnx1_pcell_0/nand3x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X31 m1_5643_945# dffsnrnx1_pcell_0/m1_1660_723# dffsnrnx1_pcell_0/nand3x1_pcell_5/li_393_182# GND nshort w=3 l=0.15
X32 dffsnrnx1_pcell_0/nand3x1_pcell_5/li_393_182# SN dffsnrnx1_pcell_0/nand3x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X33 VDD m1_4715_501# m1_5643_945# VDD pshort w=2 l=0.15
X34 VDD SN m1_5643_945# VDD pshort w=2 l=0.15
X35 VDD dffsnrnx1_pcell_0/m1_1660_723# m1_5643_945# VDD pshort w=2 l=0.15
X36 GND D dffsnrnx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X37 dffsnrnx1_pcell_1/m1_831_501# dffsnrnx1_pcell_1/m1_716_649# dffsnrnx1_pcell_1/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X38 dffsnrnx1_pcell_1/nand3x1_pcell_0/li_393_182# RN dffsnrnx1_pcell_1/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X39 VDD D dffsnrnx1_pcell_1/m1_831_501# VDD pshort w=2 l=0.15
X40 VDD RN dffsnrnx1_pcell_1/m1_831_501# VDD pshort w=2 l=0.15
X41 VDD dffsnrnx1_pcell_1/m1_716_649# dffsnrnx1_pcell_1/m1_831_501# VDD pshort w=2 l=0.15
X42 GND dffsnrnx1_pcell_1/m1_831_501# dffsnrnx1_pcell_1/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X43 dffsnrnx1_pcell_1/m1_716_649# dffsnrnx1_pcell_1/m1_1660_723# dffsnrnx1_pcell_1/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X44 dffsnrnx1_pcell_1/nand3x1_pcell_1/li_393_182# CLK dffsnrnx1_pcell_1/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X45 VDD dffsnrnx1_pcell_1/m1_831_501# dffsnrnx1_pcell_1/m1_716_649# VDD pshort w=2 l=0.15
X46 VDD CLK dffsnrnx1_pcell_1/m1_716_649# VDD pshort w=2 l=0.15
X47 VDD dffsnrnx1_pcell_1/m1_1660_723# dffsnrnx1_pcell_1/m1_716_649# VDD pshort w=2 l=0.15
X48 GND dffsnrnx1_pcell_1/m1_831_501# dffsnrnx1_pcell_1/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X49 dffsnrnx1_pcell_1/m1_2757_501# dffsnrnx1_pcell_1/m1_1660_723# dffsnrnx1_pcell_1/nand3x1_pcell_2/li_393_182# GND nshort w=3 l=0.15
X50 dffsnrnx1_pcell_1/nand3x1_pcell_2/li_393_182# SN dffsnrnx1_pcell_1/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X51 VDD dffsnrnx1_pcell_1/m1_831_501# dffsnrnx1_pcell_1/m1_2757_501# VDD pshort w=2 l=0.15
X52 VDD SN dffsnrnx1_pcell_1/m1_2757_501# VDD pshort w=2 l=0.15
X53 VDD dffsnrnx1_pcell_1/m1_1660_723# dffsnrnx1_pcell_1/m1_2757_501# VDD pshort w=2 l=0.15
X54 GND dffsnrnx1_pcell_1/m1_2757_501# dffsnrnx1_pcell_1/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X55 dffsnrnx1_pcell_1/m1_1660_723# RN dffsnrnx1_pcell_1/nand3x1_pcell_3/li_393_182# GND nshort w=3 l=0.15
X56 dffsnrnx1_pcell_1/nand3x1_pcell_3/li_393_182# CLK dffsnrnx1_pcell_1/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X57 VDD dffsnrnx1_pcell_1/m1_2757_501# dffsnrnx1_pcell_1/m1_1660_723# VDD pshort w=2 l=0.15
X58 VDD CLK dffsnrnx1_pcell_1/m1_1660_723# VDD pshort w=2 l=0.15
X59 VDD RN dffsnrnx1_pcell_1/m1_1660_723# VDD pshort w=2 l=0.15
X60 GND dffsnrnx1_pcell_1/m1_716_649# dffsnrnx1_pcell_1/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X61 m1_10487_501# m1_11449_723# dffsnrnx1_pcell_1/nand3x1_pcell_4/li_393_182# GND nshort w=3 l=0.15
X62 dffsnrnx1_pcell_1/nand3x1_pcell_4/li_393_182# RN dffsnrnx1_pcell_1/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X63 VDD dffsnrnx1_pcell_1/m1_716_649# m1_10487_501# VDD pshort w=2 l=0.15
X64 VDD RN m1_10487_501# VDD pshort w=2 l=0.15
X65 VDD m1_11449_723# m1_10487_501# VDD pshort w=2 l=0.15
X66 GND m1_10487_501# dffsnrnx1_pcell_1/nand3x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X67 m1_11449_723# dffsnrnx1_pcell_1/m1_1660_723# dffsnrnx1_pcell_1/nand3x1_pcell_5/li_393_182# GND nshort w=3 l=0.15
X68 dffsnrnx1_pcell_1/nand3x1_pcell_5/li_393_182# SN dffsnrnx1_pcell_1/nand3x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X69 VDD m1_10487_501# m1_11449_723# VDD pshort w=2 l=0.15
X70 VDD SN m1_11449_723# VDD pshort w=2 l=0.15
X71 VDD dffsnrnx1_pcell_1/m1_1660_723# m1_11449_723# VDD pshort w=2 l=0.15
X72 GND D dffsnrnx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X73 dffsnrnx1_pcell_2/m1_831_501# dffsnrnx1_pcell_2/m1_716_649# dffsnrnx1_pcell_2/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X74 dffsnrnx1_pcell_2/nand3x1_pcell_0/li_393_182# RN dffsnrnx1_pcell_2/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X75 VDD D dffsnrnx1_pcell_2/m1_831_501# VDD pshort w=2 l=0.15
X76 VDD RN dffsnrnx1_pcell_2/m1_831_501# VDD pshort w=2 l=0.15
X77 VDD dffsnrnx1_pcell_2/m1_716_649# dffsnrnx1_pcell_2/m1_831_501# VDD pshort w=2 l=0.15
X78 GND dffsnrnx1_pcell_2/m1_831_501# dffsnrnx1_pcell_2/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X79 dffsnrnx1_pcell_2/m1_716_649# dffsnrnx1_pcell_2/m1_1660_723# dffsnrnx1_pcell_2/nand3x1_pcell_1/li_393_182# GND nshort w=3 l=0.15
X80 dffsnrnx1_pcell_2/nand3x1_pcell_1/li_393_182# CLK dffsnrnx1_pcell_2/nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X81 VDD dffsnrnx1_pcell_2/m1_831_501# dffsnrnx1_pcell_2/m1_716_649# VDD pshort w=2 l=0.15
X82 VDD CLK dffsnrnx1_pcell_2/m1_716_649# VDD pshort w=2 l=0.15
X83 VDD dffsnrnx1_pcell_2/m1_1660_723# dffsnrnx1_pcell_2/m1_716_649# VDD pshort w=2 l=0.15
X84 GND dffsnrnx1_pcell_2/m1_831_501# dffsnrnx1_pcell_2/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X85 dffsnrnx1_pcell_2/m1_2757_501# dffsnrnx1_pcell_2/m1_1660_723# dffsnrnx1_pcell_2/nand3x1_pcell_2/li_393_182# GND nshort w=3 l=0.15
X86 dffsnrnx1_pcell_2/nand3x1_pcell_2/li_393_182# SN dffsnrnx1_pcell_2/nand3x1_pcell_2/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X87 VDD dffsnrnx1_pcell_2/m1_831_501# dffsnrnx1_pcell_2/m1_2757_501# VDD pshort w=2 l=0.15
X88 VDD SN dffsnrnx1_pcell_2/m1_2757_501# VDD pshort w=2 l=0.15
X89 VDD dffsnrnx1_pcell_2/m1_1660_723# dffsnrnx1_pcell_2/m1_2757_501# VDD pshort w=2 l=0.15
X90 GND dffsnrnx1_pcell_2/m1_2757_501# dffsnrnx1_pcell_2/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X91 dffsnrnx1_pcell_2/m1_1660_723# RN dffsnrnx1_pcell_2/nand3x1_pcell_3/li_393_182# GND nshort w=3 l=0.15
X92 dffsnrnx1_pcell_2/nand3x1_pcell_3/li_393_182# CLK dffsnrnx1_pcell_2/nand3x1_pcell_3/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X93 VDD dffsnrnx1_pcell_2/m1_2757_501# dffsnrnx1_pcell_2/m1_1660_723# VDD pshort w=2 l=0.15
X94 VDD CLK dffsnrnx1_pcell_2/m1_1660_723# VDD pshort w=2 l=0.15
X95 VDD RN dffsnrnx1_pcell_2/m1_1660_723# VDD pshort w=2 l=0.15
X96 GND dffsnrnx1_pcell_2/m1_716_649# dffsnrnx1_pcell_2/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X97 m1_16259_501# m1_16111_427# dffsnrnx1_pcell_2/nand3x1_pcell_4/li_393_182# GND nshort w=3 l=0.15
X98 dffsnrnx1_pcell_2/nand3x1_pcell_4/li_393_182# RN dffsnrnx1_pcell_2/nand3x1_pcell_4/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X99 VDD dffsnrnx1_pcell_2/m1_716_649# m1_16259_501# VDD pshort w=2 l=0.15
X100 VDD RN m1_16259_501# VDD pshort w=2 l=0.15
X101 VDD m1_16111_427# m1_16259_501# VDD pshort w=2 l=0.15
X102 GND m1_16259_501# dffsnrnx1_pcell_2/nand3x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X103 m1_16111_427# dffsnrnx1_pcell_2/m1_1660_723# dffsnrnx1_pcell_2/nand3x1_pcell_5/li_393_182# GND nshort w=3 l=0.15
X104 dffsnrnx1_pcell_2/nand3x1_pcell_5/li_393_182# SN dffsnrnx1_pcell_2/nand3x1_pcell_5/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X105 VDD m1_16259_501# m1_16111_427# VDD pshort w=2 l=0.15
X106 VDD SN m1_16111_427# VDD pshort w=2 l=0.15
X107 VDD dffsnrnx1_pcell_2/m1_1660_723# m1_16111_427# VDD pshort w=2 l=0.15
X108 GND m1_5643_945# voter3x1_pcell_0/votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X109 GND m1_5643_945# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X110 GND m1_16111_427# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X111 voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# m1_5643_945# VDD VDD pshort w=2 l=0.15
X112 voter3x1_pcell_0/m1_1867_797# m1_16111_427# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_1/a_0_0# GND nshort w=3 l=0.15
X113 voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# m1_11449_723# VDD VDD pshort w=2 l=0.15
X114 voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# m1_16111_427# voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X115 voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# m1_5643_945# voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# VDD pshort w=2 l=0.15
X116 voter3x1_pcell_0/m1_1867_797# m1_16111_427# voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X117 voter3x1_pcell_0/m1_1867_797# m1_11449_723# voter3x1_pcell_0/votern3x1_pcell_0/a_893_1059# VDD pshort w=2 l=0.15
X118 voter3x1_pcell_0/m1_1867_797# m1_11449_723# voter3x1_pcell_0/votern3x1_pcell_0/nmos_top_0/a_0_0# GND nshort w=3 l=0.15
X119 voter3x1_pcell_0/m1_1867_797# m1_11449_723# voter3x1_pcell_0/votern3x1_pcell_0/nmos_bottom_2/a_0_0# GND nshort w=3 l=0.15
X120 Q voter3x1_pcell_0/m1_1867_797# GND GND nshort w=3 l=0.15
X121 VDD voter3x1_pcell_0/m1_1867_797# Q VDD pshort w=2 l=0.15
C0 SN dffsnrnx1_pcell_2/m1_716_649# 3.98fF
C1 D CLK 11.68fF
C2 VDD RN 2.54fF
C3 SN CLK 2.43fF
C4 m1_5643_945# CLK 10.85fF
C5 SN m1_11449_723# 2.80fF
C6 D VDD 5.91fF
C7 m1_5643_945# m1_11449_723# 5.28fF
C8 D RN 2.05fF
C9 dffsnrnx1_pcell_2/m1_716_649# m1_11449_723# 2.04fF
C10 dffsnrnx1_pcell_2/m1_716_649# dffsnrnx1_pcell_2/m1_1660_723# 3.19fF
C11 dffsnrnx1_pcell_1/m1_716_649# dffsnrnx1_pcell_1/m1_1660_723# 3.19fF
C12 m1_5643_945# VDD 6.87fF
C13 SN RN 5.64fF
C14 m1_11449_723# CLK 3.10fF
C15 dffsnrnx1_pcell_1/m1_716_649# SN 3.98fF
C16 voter3x1_pcell_0/votern3x1_pcell_0/a_805_1331# VDD 2.05fF
C17 VDD CLK 7.14fF
C18 D dffsnrnx1_pcell_1/m1_1660_723# 4.46fF
C19 RN CLK 2.23fF
C20 dffsnrnx1_pcell_2/m1_1660_723# m1_11449_723# 4.46fF
C21 D SN 2.38fF
C22 D m1_5643_945# 3.08fF
C23 dffsnrnx1_pcell_0/m1_1660_723# D 4.47fF
C24 dffsnrnx1_pcell_0/m1_716_649# SN 2.04fF
C25 VDD m1_11449_723# 4.03fF
C26 dffsnrnx1_pcell_0/m1_1660_723# dffsnrnx1_pcell_0/m1_716_649# 3.19fF
C27 m1_5643_945# SN 5.30fF
C28 VDD GND 3.02fF
.ends
