magic
tech sky130A
magscale 1 2
timestamp 1669215543
<< nwell >>
rect 87 885 136 1550
rect 31 823 190 885
rect 87 786 136 823
<< pwell >>
rect -34 -34 256 544
<< psubdiff >>
rect 34 482 188 544
rect 34 -17 94 17
rect 128 -17 188 17
rect 34 -34 188 -17
<< nsubdiff >>
rect 34 1497 188 1514
rect 34 1463 94 1497
rect 128 1463 188 1497
rect 34 822 188 884
<< psubdiffcont >>
rect 94 -17 128 17
<< nsubdiffcont >>
rect 94 1463 128 1497
<< locali >>
rect 34 1497 188 1514
rect 34 1463 94 1497
rect 128 1463 188 1497
rect 34 1446 188 1463
rect 34 17 188 34
rect 34 -17 94 17
rect 128 -17 188 17
rect 34 -34 188 -17
<< metal1 >>
rect 34 1446 188 1514
rect -34 -34 256 34
use diff_ring_side  diff_ring_side_0 pcells
timestamp 1652319726
transform 1 0 0 0 1 0
box -87 -34 87 1550
use diff_ring_side  diff_ring_side_1
timestamp 1652319726
transform 1 0 222 0 1 0
box -87 -34 87 1550
<< labels >>
rlabel metal1 -34 1446 256 1514 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 -34 -34 256 34 1 GND
port 2 nsew ground bidirectional abutment
<< properties >>
string LEFclass CORE SPACER
string LEFsite unitrh
string FIXED_BBOX 0 0 222 1480
string LEFsymmetry X Y R90
<< end >>
