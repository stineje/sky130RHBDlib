* SPICE3 file created from XNOR2X1.ext - technology: sky130A

.subckt XNOR2X1 Y A B VDD GND
X0 Y B a_575_1004 VDD pshort w=2 l=0.15 M=2
X1 a_1241_1004 a_185_182 Y VDD pshort w=2 l=0.15 M=2
X2 VDD B a_806_165 VDD pshort w=2 l=0.15 M=2
X3 a_185_182 A GND GND nshort w=3 l=0.15
X4 Y a_806_165 a_556_73 GND nshort w=3 l=0.15
X5 VDD A a_575_1004 VDD pshort w=2 l=0.15 M=2
X6 VDD A a_185_182 VDD pshort w=2 l=0.15 M=2
X7 a_806_165 B GND GND nshort w=3 l=0.15
X8 VDD a_806_165 a_1241_1004 VDD pshort w=2 l=0.15 M=2
X9 GND B a_1222_73 GND nshort w=3 l=0.15
X10 GND A a_556_73 GND nshort w=3 l=0.15
X11 Y a_185_182 a_1222_73 GND nshort w=3 l=0.15
C0 B a_806_165 2.21fF
C1 VDD GND 5.63fF
.ends
