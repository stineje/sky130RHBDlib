magic
tech sky130A
magscale 1 2
timestamp 1645210163
use sky130_fd_io__top_gpio_pad  sky130_fd_io__top_gpio_pad_0
timestamp 1645210163
transform 1 0 0 0 1 0
box 960 18991 14040 34071
use sky130_fd_io__com_bus_hookup  sky130_fd_io__com_bus_hookup_0
timestamp 1645210163
transform 1 0 0 0 1 0
box 0 -142 15000 39451
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 27722820
string GDS_START 27722714
<< end >>
