* SPICE3 file created from AOI3X1.ext - technology: sky130A

.subckt AOI3X1 YN A B C VDD GND
M1000 YN.t3 C.t0 a_797_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 YN a_217_1050.t6 GND.t2 nshort w=-1.605u l=1.765u
+  ad=0.3582p pd=3.15u as=0p ps=0u
M1002 GND A.t1 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=2.1157p pd=14.51u as=0p ps=0u
M1003 VDD.t5 a_217_1050.t5 a_797_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VDD.t2 A.t0 a_217_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VDD.t0 B.t0 a_217_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 YN C.t2 GND.t1 nshort w=-1.83u l=2.06u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_217_1050.t1 A.t2 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_797_1051.t1 C.t1 YN.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_797_1051.t3 a_217_1050.t7 VDD.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 YN C GND GND nshort w=3u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_217_1050.t4 B.t2 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 YN VDD 0.25fF
C1 C VDD 0.07fF
C2 B A 0.27fF
C3 YN C 0.26fF
C4 VDD A 0.08fF
C5 B VDD 0.07fF
R0 C.n0 C.t1 470.752
R1 C.n0 C.t0 384.527
R2 C.n1 C.t2 241.172
R3 C.n1 C.n0 110.173
R4 C.n2 C.n1 76
R5 C.n2 C 0.046
R6 a_797_1051.t0 a_797_1051.n0 101.66
R7 a_797_1051.n0 a_797_1051.t1 101.659
R8 a_797_1051.n0 a_797_1051.t2 14.294
R9 a_797_1051.n0 a_797_1051.t3 14.282
R10 YN.n8 YN.n7 188.74
R11 YN.n8 YN.n0 138.783
R12 YN.n7 YN.n6 133.539
R13 YN.n3 YN.n1 80.526
R14 YN.n9 YN.n8 76
R15 YN.n7 YN.n3 48.405
R16 YN.n3 YN.n2 30
R17 YN.n6 YN.n5 22.578
R18 YN.n0 YN.t2 14.282
R19 YN.n0 YN.t3 14.282
R20 YN.n6 YN.n4 8.58
R21 YN.n9 YN 0.046
R22 a_217_1050.n4 a_217_1050.t7 486.819
R23 a_217_1050.n4 a_217_1050.t5 384.527
R24 a_217_1050.n6 a_217_1050.n3 232.158
R25 a_217_1050.n5 a_217_1050.t6 197.395
R26 a_217_1050.n5 a_217_1050.n4 186.206
R27 a_217_1050.n6 a_217_1050.n5 153.315
R28 a_217_1050.n8 a_217_1050.n6 130.933
R29 a_217_1050.n3 a_217_1050.n2 76.002
R30 a_217_1050.n8 a_217_1050.n7 30
R31 a_217_1050.n9 a_217_1050.n0 24.383
R32 a_217_1050.n9 a_217_1050.n8 23.684
R33 a_217_1050.n1 a_217_1050.t0 14.282
R34 a_217_1050.n1 a_217_1050.t4 14.282
R35 a_217_1050.n2 a_217_1050.t2 14.282
R36 a_217_1050.n2 a_217_1050.t1 14.282
R37 a_217_1050.n3 a_217_1050.n1 12.85
R38 VDD.n134 VDD.n132 144.705
R39 VDD.n40 VDD.n39 76
R40 VDD.n47 VDD.n46 76
R41 VDD.n51 VDD.n50 76
R42 VDD.n77 VDD.n76 76
R43 VDD.n136 VDD.n135 76
R44 VDD.n131 VDD.n130 76
R45 VDD.n126 VDD.n125 76
R46 VDD.n121 VDD.n120 76
R47 VDD.n115 VDD.n114 76
R48 VDD.n110 VDD.n109 76
R49 VDD.n105 VDD.n104 76
R50 VDD.n100 VDD.n99 76
R51 VDD.n101 VDD.t1 55.106
R52 VDD.n127 VDD.t0 55.106
R53 VDD.n42 VDD.n41 41.183
R54 VDD.n117 VDD.n116 40.824
R55 VDD.n67 VDD.n66 36.774
R56 VDD.n123 VDD.n122 36.608
R57 VDD.n34 VDD.n33 34.942
R58 VDD.n44 VDD.n43 32.032
R59 VDD.n107 VDD.n106 32.032
R60 VDD.n99 VDD.n96 21.841
R61 VDD.n23 VDD.n20 21.841
R62 VDD.n116 VDD.t3 14.282
R63 VDD.n116 VDD.t2 14.282
R64 VDD.n41 VDD.t4 14.282
R65 VDD.n41 VDD.t5 14.282
R66 VDD.n96 VDD.n79 14.167
R67 VDD.n79 VDD.n78 14.167
R68 VDD.n72 VDD.n53 14.167
R69 VDD.n53 VDD.n52 14.167
R70 VDD.n20 VDD.n19 14.167
R71 VDD.n19 VDD.n17 14.167
R72 VDD.n32 VDD.n29 14.167
R73 VDD.n29 VDD.n28 14.167
R74 VDD.n76 VDD.n73 14.167
R75 VDD.n23 VDD.n22 13.653
R76 VDD.n22 VDD.n21 13.653
R77 VDD.n32 VDD.n31 13.653
R78 VDD.n31 VDD.n30 13.653
R79 VDD.n29 VDD.n25 13.653
R80 VDD.n25 VDD.n24 13.653
R81 VDD.n28 VDD.n27 13.653
R82 VDD.n27 VDD.n26 13.653
R83 VDD.n39 VDD.n38 13.653
R84 VDD.n38 VDD.n37 13.653
R85 VDD.n46 VDD.n45 13.653
R86 VDD.n45 VDD.n44 13.653
R87 VDD.n50 VDD.n49 13.653
R88 VDD.n49 VDD.n48 13.653
R89 VDD.n76 VDD.n75 13.653
R90 VDD.n75 VDD.n74 13.653
R91 VDD.n135 VDD.n134 13.653
R92 VDD.n134 VDD.n133 13.653
R93 VDD.n130 VDD.n129 13.653
R94 VDD.n129 VDD.n128 13.653
R95 VDD.n125 VDD.n124 13.653
R96 VDD.n124 VDD.n123 13.653
R97 VDD.n120 VDD.n119 13.653
R98 VDD.n119 VDD.n118 13.653
R99 VDD.n114 VDD.n113 13.653
R100 VDD.n113 VDD.n112 13.653
R101 VDD.n109 VDD.n108 13.653
R102 VDD.n108 VDD.n107 13.653
R103 VDD.n104 VDD.n103 13.653
R104 VDD.n103 VDD.n102 13.653
R105 VDD.n99 VDD.n98 13.653
R106 VDD.n98 VDD.n97 13.653
R107 VDD.n4 VDD.n2 12.915
R108 VDD.n4 VDD.n3 12.66
R109 VDD.n10 VDD.n9 12.343
R110 VDD.n12 VDD.n11 12.343
R111 VDD.n10 VDD.n7 12.343
R112 VDD.n120 VDD.n117 8.658
R113 VDD.n73 VDD.n72 7.674
R114 VDD.n57 VDD.n56 7.5
R115 VDD.n60 VDD.n59 7.5
R116 VDD.n62 VDD.n61 7.5
R117 VDD.n65 VDD.n64 7.5
R118 VDD.n72 VDD.n71 7.5
R119 VDD.n91 VDD.n90 7.5
R120 VDD.n85 VDD.n84 7.5
R121 VDD.n87 VDD.n86 7.5
R122 VDD.n93 VDD.n83 7.5
R123 VDD.n93 VDD.n81 7.5
R124 VDD.n96 VDD.n95 7.5
R125 VDD.n20 VDD.n16 7.5
R126 VDD.n2 VDD.n1 7.5
R127 VDD.n9 VDD.n8 7.5
R128 VDD.n7 VDD.n6 7.5
R129 VDD.n19 VDD.n18 7.5
R130 VDD.n14 VDD.n0 7.5
R131 VDD.n94 VDD.n80 6.772
R132 VDD.n92 VDD.n89 6.772
R133 VDD.n88 VDD.n85 6.772
R134 VDD.n88 VDD.n87 6.772
R135 VDD.n92 VDD.n91 6.772
R136 VDD.n95 VDD.n94 6.772
R137 VDD.n71 VDD.n70 6.772
R138 VDD.n58 VDD.n55 6.772
R139 VDD.n63 VDD.n60 6.772
R140 VDD.n68 VDD.n65 6.772
R141 VDD.n68 VDD.n67 6.772
R142 VDD.n63 VDD.n62 6.772
R143 VDD.n58 VDD.n57 6.772
R144 VDD.n70 VDD.n54 6.772
R145 VDD.n33 VDD.n23 6.487
R146 VDD.n33 VDD.n32 6.475
R147 VDD.n16 VDD.n15 6.458
R148 VDD.n83 VDD.n82 6.202
R149 VDD.n46 VDD.n42 5.903
R150 VDD.n37 VDD.n36 4.576
R151 VDD.n112 VDD.n111 4.576
R152 VDD.n104 VDD.n101 2.754
R153 VDD.n130 VDD.n127 2.361
R154 VDD.n14 VDD.n5 1.329
R155 VDD.n14 VDD.n10 1.329
R156 VDD.n14 VDD.n12 1.329
R157 VDD.n14 VDD.n13 1.329
R158 VDD.n15 VDD.n14 0.696
R159 VDD.n14 VDD.n4 0.696
R160 VDD.n93 VDD.n92 0.365
R161 VDD.n93 VDD.n88 0.365
R162 VDD.n94 VDD.n93 0.365
R163 VDD.n69 VDD.n68 0.365
R164 VDD.n69 VDD.n63 0.365
R165 VDD.n69 VDD.n58 0.365
R166 VDD.n70 VDD.n69 0.365
R167 VDD.n100 VDD 0.207
R168 VDD.n40 VDD.n35 0.181
R169 VDD.n121 VDD.n115 0.181
R170 VDD.n35 VDD.n34 0.145
R171 VDD.n47 VDD.n40 0.145
R172 VDD.n51 VDD.n47 0.145
R173 VDD.n77 VDD.n51 0.145
R174 VDD VDD.n77 0.145
R175 VDD VDD.n136 0.145
R176 VDD.n136 VDD.n131 0.145
R177 VDD.n131 VDD.n126 0.145
R178 VDD.n126 VDD.n121 0.145
R179 VDD.n115 VDD.n110 0.145
R180 VDD.n110 VDD.n105 0.145
R181 VDD.n105 VDD.n100 0.145
R182 A.n0 A.t0 480.392
R183 A.n0 A.t2 403.272
R184 A.n1 A.t1 230.374
R185 A.n1 A.n0 151.553
R186 A.n2 A.n1 76
R187 A.n2 A 0.046
R188 GND.n39 GND.n38 219.745
R189 GND.n39 GND.n37 85.529
R190 GND.n8 GND.n1 76.145
R191 GND.n45 GND.n44 76
R192 GND.n8 GND.n7 76
R193 GND.n14 GND.n13 76
R194 GND.n17 GND.n16 76
R195 GND.n23 GND.n22 76
R196 GND.n28 GND.n27 76
R197 GND.n35 GND.n34 76
R198 GND.n42 GND.n41 76
R199 GND.n71 GND.n70 76
R200 GND.n68 GND.n67 76
R201 GND.n65 GND.n64 76
R202 GND.n62 GND.n61 76
R203 GND.n59 GND.n58 76
R204 GND.n56 GND.n55 76
R205 GND.n48 GND.n47 76
R206 GND.n53 GND.n52 63.835
R207 GND.n52 GND.n51 28.421
R208 GND.n52 GND.n50 25.263
R209 GND.n50 GND.n49 24.383
R210 GND.n25 GND.n24 19.735
R211 GND.n20 GND.n19 19.735
R212 GND.n12 GND.n11 19.735
R213 GND.n5 GND.n4 19.735
R214 GND.n33 GND.n32 19.735
R215 GND.n11 GND.t1 19.724
R216 GND.n24 GND.t2 19.724
R217 GND.n41 GND.n40 14.167
R218 GND.n47 GND.n46 13.653
R219 GND.n55 GND.n54 13.653
R220 GND.n58 GND.n57 13.653
R221 GND.n61 GND.n60 13.653
R222 GND.n64 GND.n63 13.653
R223 GND.n67 GND.n66 13.653
R224 GND.n70 GND.n69 13.653
R225 GND.n41 GND.n36 13.653
R226 GND.n34 GND.n29 13.653
R227 GND.n27 GND.n26 13.653
R228 GND.n22 GND.n21 13.653
R229 GND.n16 GND.n15 13.653
R230 GND.n13 GND.n9 13.653
R231 GND.n7 GND.n6 13.653
R232 GND.n32 GND.n31 12.837
R233 GND.n4 GND.n3 11.605
R234 GND.n3 GND.n2 9.809
R235 GND.n22 GND.n20 8.854
R236 GND.n31 GND.n30 7.566
R237 GND.n40 GND.n39 7.312
R238 GND.t1 GND.n10 7.04
R239 GND.n19 GND.n18 5.774
R240 GND.n13 GND.n12 3.935
R241 GND.n27 GND.n25 3.935
R242 GND.n55 GND.n53 3.935
R243 GND.n7 GND.n5 0.983
R244 GND.n34 GND.n33 0.983
R245 GND.n1 GND.n0 0.596
R246 GND.n44 GND.n43 0.596
R247 GND.n45 GND 0.207
R248 GND.n23 GND.n17 0.181
R249 GND.n62 GND.n59 0.181
R250 GND.n14 GND.n8 0.145
R251 GND.n17 GND.n14 0.145
R252 GND.n28 GND.n23 0.145
R253 GND.n35 GND.n28 0.145
R254 GND.n42 GND.n35 0.145
R255 GND GND.n42 0.145
R256 GND GND.n71 0.145
R257 GND.n71 GND.n68 0.145
R258 GND.n68 GND.n65 0.145
R259 GND.n65 GND.n62 0.145
R260 GND.n59 GND.n56 0.145
R261 GND.n56 GND.n48 0.145
R262 GND.n48 GND.n45 0.145
R263 a_112_101.t0 a_112_101.n1 34.62
R264 a_112_101.t0 a_112_101.n0 8.137
R265 a_112_101.t0 a_112_101.n2 4.69
R266 B.n0 B.t0 472.359
R267 B.n0 B.t2 384.527
R268 B.n1 B.t1 214.619
R269 B.n1 B.n0 136.613
R270 B.n2 B.n1 76
R271 B.n2 B 0.046
C6 VDD GND 5.71fF
C7 a_112_101.n0 GND 0.05fF
C8 a_112_101.n1 GND 0.12fF
C9 a_112_101.n2 GND 0.04fF
C10 VDD.n0 GND 0.14fF
C11 VDD.n1 GND 0.02fF
C12 VDD.n2 GND 0.02fF
C13 VDD.n3 GND 0.04fF
C14 VDD.n4 GND 0.01fF
C15 VDD.n6 GND 0.02fF
C16 VDD.n7 GND 0.02fF
C17 VDD.n8 GND 0.02fF
C18 VDD.n9 GND 0.02fF
C19 VDD.n11 GND 0.02fF
C20 VDD.n14 GND 0.43fF
C21 VDD.n16 GND 0.03fF
C22 VDD.n17 GND 0.02fF
C23 VDD.n18 GND 0.02fF
C24 VDD.n19 GND 0.02fF
C25 VDD.n20 GND 0.03fF
C26 VDD.n21 GND 0.26fF
C27 VDD.n22 GND 0.02fF
C28 VDD.n23 GND 0.03fF
C29 VDD.n24 GND 0.26fF
C30 VDD.n25 GND 0.01fF
C31 VDD.n26 GND 0.28fF
C32 VDD.n27 GND 0.01fF
C33 VDD.n28 GND 0.02fF
C34 VDD.n29 GND 0.02fF
C35 VDD.n30 GND 0.26fF
C36 VDD.n31 GND 0.01fF
C37 VDD.n32 GND 0.02fF
C38 VDD.n33 GND 0.00fF
C39 VDD.n34 GND 0.08fF
C40 VDD.n35 GND 0.02fF
C41 VDD.n36 GND 0.16fF
C42 VDD.n37 GND 0.13fF
C43 VDD.n38 GND 0.01fF
C44 VDD.n39 GND 0.02fF
C45 VDD.n40 GND 0.02fF
C46 VDD.n41 GND 0.10fF
C47 VDD.n42 GND 0.02fF
C48 VDD.n43 GND 0.13fF
C49 VDD.n44 GND 0.15fF
C50 VDD.n45 GND 0.01fF
C51 VDD.n46 GND 0.02fF
C52 VDD.n47 GND 0.02fF
C53 VDD.n48 GND 0.23fF
C54 VDD.n49 GND 0.01fF
C55 VDD.n50 GND 0.02fF
C56 VDD.n51 GND 0.02fF
C57 VDD.n52 GND 0.02fF
C58 VDD.n53 GND 0.02fF
C59 VDD.n54 GND 0.02fF
C60 VDD.n55 GND 0.02fF
C61 VDD.n56 GND 0.02fF
C62 VDD.n57 GND 0.02fF
C63 VDD.n59 GND 0.02fF
C64 VDD.n60 GND 0.02fF
C65 VDD.n61 GND 0.02fF
C66 VDD.n62 GND 0.02fF
C67 VDD.n64 GND 0.03fF
C68 VDD.n65 GND 0.02fF
C69 VDD.n66 GND 0.21fF
C70 VDD.n67 GND 0.04fF
C71 VDD.n69 GND 0.26fF
C72 VDD.n71 GND 0.02fF
C73 VDD.n72 GND 0.02fF
C74 VDD.n73 GND 0.03fF
C75 VDD.n74 GND 0.26fF
C76 VDD.n75 GND 0.01fF
C77 VDD.n76 GND 0.02fF
C78 VDD.n77 GND 0.02fF
C79 VDD.n78 GND 0.02fF
C80 VDD.n79 GND 0.02fF
C81 VDD.n80 GND 0.02fF
C82 VDD.n81 GND 0.14fF
C83 VDD.n82 GND 0.03fF
C84 VDD.n83 GND 0.02fF
C85 VDD.n84 GND 0.02fF
C86 VDD.n85 GND 0.02fF
C87 VDD.n86 GND 0.02fF
C88 VDD.n87 GND 0.02fF
C89 VDD.n89 GND 0.02fF
C90 VDD.n90 GND 0.02fF
C91 VDD.n91 GND 0.02fF
C92 VDD.n93 GND 0.43fF
C93 VDD.n95 GND 0.03fF
C94 VDD.n96 GND 0.03fF
C95 VDD.n97 GND 0.26fF
C96 VDD.n98 GND 0.02fF
C97 VDD.n99 GND 0.03fF
C98 VDD.n100 GND 0.03fF
C99 VDD.n101 GND 0.06fF
C100 VDD.n102 GND 0.23fF
C101 VDD.n103 GND 0.01fF
C102 VDD.n104 GND 0.01fF
C103 VDD.n105 GND 0.02fF
C104 VDD.n106 GND 0.13fF
C105 VDD.n107 GND 0.15fF
C106 VDD.n108 GND 0.01fF
C107 VDD.n109 GND 0.02fF
C108 VDD.n110 GND 0.02fF
C109 VDD.n111 GND 0.16fF
C110 VDD.n112 GND 0.13fF
C111 VDD.n113 GND 0.01fF
C112 VDD.n114 GND 0.02fF
C113 VDD.n115 GND 0.02fF
C114 VDD.n116 GND 0.10fF
C115 VDD.n117 GND 0.02fF
C116 VDD.n118 GND 0.28fF
C117 VDD.n119 GND 0.01fF
C118 VDD.n120 GND 0.02fF
C119 VDD.n121 GND 0.02fF
C120 VDD.n122 GND 0.13fF
C121 VDD.n123 GND 0.16fF
C122 VDD.n124 GND 0.01fF
C123 VDD.n125 GND 0.02fF
C124 VDD.n126 GND 0.02fF
C125 VDD.n127 GND 0.05fF
C126 VDD.n128 GND 0.23fF
C127 VDD.n129 GND 0.01fF
C128 VDD.n130 GND 0.01fF
C129 VDD.n131 GND 0.02fF
C130 VDD.n132 GND 0.02fF
C131 VDD.n133 GND 0.26fF
C132 VDD.n134 GND 0.01fF
C133 VDD.n135 GND 0.02fF
C134 VDD.n136 GND 0.02fF
C135 a_217_1050.n0 GND 0.03fF
C136 a_217_1050.n1 GND 0.42fF
C137 a_217_1050.n2 GND 0.50fF
C138 a_217_1050.n3 GND 0.32fF
C139 a_217_1050.n4 GND 0.36fF
C140 a_217_1050.n5 GND 0.45fF
C141 a_217_1050.n6 GND 0.48fF
C142 a_217_1050.n7 GND 0.03fF
C143 a_217_1050.n8 GND 0.16fF
C144 a_217_1050.n9 GND 0.04fF
C145 YN.n0 GND 0.64fF
C146 YN.n1 GND 0.06fF
C147 YN.n2 GND 0.03fF
C148 YN.n3 GND 0.13fF
C149 YN.n4 GND 0.04fF
C150 YN.n5 GND 0.05fF
C151 YN.n6 GND 0.19fF
C152 YN.n7 GND 0.45fF
C153 YN.n8 GND 0.39fF
C154 YN.n9 GND 0.01fF
C155 a_797_1051.n0 GND 0.52fF
.ends
