magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 530 157 735 203
rect 1 21 735 157
rect 30 -17 64 21
<< locali >>
rect 122 265 156 492
rect 651 432 719 493
rect 122 199 225 265
rect 300 199 381 323
rect 653 299 719 432
rect 483 153 551 265
rect 674 165 719 299
rect 651 51 719 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 27 165 79 425
rect 191 343 241 527
rect 331 363 449 416
rect 511 369 577 527
rect 415 333 449 363
rect 415 299 619 333
rect 415 165 449 299
rect 585 265 619 299
rect 27 131 449 165
rect 585 199 640 265
rect 27 51 79 131
rect 331 128 449 131
rect 175 17 241 97
rect 331 51 397 128
rect 509 17 576 94
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 122 199 225 265 6 A
port 1 nsew signal input
rlabel locali s 122 265 156 492 6 A
port 1 nsew signal input
rlabel locali s 300 199 381 323 6 B
port 2 nsew signal input
rlabel locali s 483 153 551 265 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 735 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 530 157 735 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 651 51 719 165 6 X
port 8 nsew signal output
rlabel locali s 674 165 719 299 6 X
port 8 nsew signal output
rlabel locali s 653 299 719 432 6 X
port 8 nsew signal output
rlabel locali s 651 432 719 493 6 X
port 8 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 736 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1663022
string GDS_START 1656898
<< end >>
