* SPICE3 file created from BUFX1.ext - technology: sky130A

.subckt BUFX1 Y A VDD GND
M1000 a_185_209.t0 A.t1 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 Y a_185_209.t3 GND.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1002 VDD.t1 a_185_209.t4 Y.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD.t2 A.t2 a_185_209.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y.t0 a_185_209.t5 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 A VDD 0.12fF
C1 VDD Y 0.79fF
R0 A.n0 A.t2 512.525
R1 A.n0 A.t1 371.139
R2 A.n1 A.t0 210.434
R3 A.n1 A.n0 173.2
R4 A.n2 A.n1 76
R5 A.n2 A 0.046
R6 GND.n28 GND.n27 219.745
R7 GND.n28 GND.n26 85.529
R8 GND.n9 GND.n1 76.145
R9 GND.n34 GND.n33 76
R10 GND.n9 GND.n8 76
R11 GND.n17 GND.n16 76
R12 GND.n24 GND.n23 76
R13 GND.n31 GND.n30 76
R14 GND.n62 GND.n61 76
R15 GND.n59 GND.n58 76
R16 GND.n51 GND.n50 76
R17 GND.n43 GND.n42 76
R18 GND.n39 GND.t1 39.412
R19 GND.n5 GND.n4 35.01
R20 GND.n55 GND.n54 35.01
R21 GND.n3 GND.n2 29.127
R22 GND.n12 GND.t0 20.794
R23 GND.n6 GND.n5 19.735
R24 GND.n14 GND.n13 19.735
R25 GND.n22 GND.n21 19.735
R26 GND.n56 GND.n55 19.735
R27 GND.n48 GND.n47 19.735
R28 GND.n41 GND.n40 19.735
R29 GND.n5 GND.n3 19.017
R30 GND.n55 GND.n53 19.017
R31 GND.n39 GND.n38 17.185
R32 GND.n30 GND.n29 14.167
R33 GND.n42 GND.n35 13.653
R34 GND.n50 GND.n49 13.653
R35 GND.n58 GND.n57 13.653
R36 GND.n61 GND.n60 13.653
R37 GND.n30 GND.n25 13.653
R38 GND.n23 GND.n18 13.653
R39 GND.n16 GND.n15 13.653
R40 GND.n8 GND.n7 13.653
R41 GND.n21 GND.n20 12.837
R42 GND.n20 GND.n19 7.566
R43 GND.n53 GND.n52 7.5
R44 GND.n46 GND.n45 7.5
R45 GND.n29 GND.n28 7.312
R46 GND.n40 GND.n39 6.139
R47 GND.n11 GND.n10 4.551
R48 GND.n37 GND.n36 4.551
R49 GND.n8 GND.n6 3.935
R50 GND.n58 GND.n56 3.935
R51 GND.n23 GND.n22 3.541
R52 GND.n42 GND.n41 3.541
R53 GND.t0 GND.n11 2.238
R54 GND.t1 GND.n37 2.238
R55 GND.n45 GND.n44 1.935
R56 GND.n1 GND.n0 0.596
R57 GND.n33 GND.n32 0.596
R58 GND.n13 GND.n12 0.358
R59 GND.n47 GND.n46 0.358
R60 GND.n34 GND 0.207
R61 GND.n16 GND.n14 0.196
R62 GND.n50 GND.n48 0.196
R63 GND.n17 GND.n9 0.157
R64 GND.n24 GND.n17 0.157
R65 GND.n59 GND.n51 0.157
R66 GND.n51 GND.n43 0.157
R67 GND.n31 GND.n24 0.145
R68 GND GND.n31 0.145
R69 GND GND.n62 0.145
R70 GND.n62 GND.n59 0.145
R71 GND.n43 GND.n34 0.145
R72 a_185_209.n1 a_185_209.t4 512.525
R73 a_185_209.n1 a_185_209.t5 371.139
R74 a_185_209.n3 a_185_209.n0 237.113
R75 a_185_209.n2 a_185_209.n1 226.306
R76 a_185_209.n2 a_185_209.t3 157.328
R77 a_185_209.n3 a_185_209.n2 153.043
R78 a_185_209.n5 a_185_209.n3 132.431
R79 a_185_209.n5 a_185_209.n4 15.218
R80 a_185_209.n0 a_185_209.t1 14.282
R81 a_185_209.n0 a_185_209.t0 14.282
R82 a_185_209.n6 a_185_209.n5 12.014
R83 VDD.n107 VDD.n105 144.705
R84 VDD.n26 VDD.n25 77.792
R85 VDD.n36 VDD.n35 77.792
R86 VDD.n101 VDD.n100 77.792
R87 VDD.n90 VDD.n89 77.792
R88 VDD.n29 VDD.n23 76.145
R89 VDD.n29 VDD.n28 76
R90 VDD.n33 VDD.n32 76
R91 VDD.n39 VDD.n38 76
R92 VDD.n65 VDD.n64 76
R93 VDD.n109 VDD.n108 76
R94 VDD.n104 VDD.n103 76
R95 VDD.n98 VDD.n97 76
R96 VDD.n94 VDD.n93 76
R97 VDD.n88 VDD.n87 76
R98 VDD.n92 VDD.t3 55.106
R99 VDD.n99 VDD.t2 55.106
R100 VDD.n34 VDD.t0 55.106
R101 VDD.n24 VDD.t1 55.106
R102 VDD.n57 VDD.n56 36.774
R103 VDD.n87 VDD.n84 21.841
R104 VDD.n23 VDD.n20 21.841
R105 VDD.n84 VDD.n67 14.167
R106 VDD.n67 VDD.n66 14.167
R107 VDD.n62 VDD.n43 14.167
R108 VDD.n43 VDD.n42 14.167
R109 VDD.n20 VDD.n19 14.167
R110 VDD.n19 VDD.n17 14.167
R111 VDD.n64 VDD.n63 14.167
R112 VDD.n23 VDD.n22 13.653
R113 VDD.n22 VDD.n21 13.653
R114 VDD.n28 VDD.n27 13.653
R115 VDD.n27 VDD.n26 13.653
R116 VDD.n32 VDD.n31 13.653
R117 VDD.n31 VDD.n30 13.653
R118 VDD.n38 VDD.n37 13.653
R119 VDD.n37 VDD.n36 13.653
R120 VDD.n64 VDD.n41 13.653
R121 VDD.n41 VDD.n40 13.653
R122 VDD.n108 VDD.n107 13.653
R123 VDD.n107 VDD.n106 13.653
R124 VDD.n103 VDD.n102 13.653
R125 VDD.n102 VDD.n101 13.653
R126 VDD.n97 VDD.n96 13.653
R127 VDD.n96 VDD.n95 13.653
R128 VDD.n93 VDD.n91 13.653
R129 VDD.n91 VDD.n90 13.653
R130 VDD.n87 VDD.n86 13.653
R131 VDD.n86 VDD.n85 13.653
R132 VDD.n4 VDD.n2 12.915
R133 VDD.n4 VDD.n3 12.66
R134 VDD.n13 VDD.n12 12.343
R135 VDD.n11 VDD.n10 12.343
R136 VDD.n8 VDD.n7 12.343
R137 VDD.n63 VDD.n62 7.674
R138 VDD.n47 VDD.n46 7.5
R139 VDD.n50 VDD.n49 7.5
R140 VDD.n52 VDD.n51 7.5
R141 VDD.n55 VDD.n54 7.5
R142 VDD.n62 VDD.n61 7.5
R143 VDD.n79 VDD.n78 7.5
R144 VDD.n73 VDD.n72 7.5
R145 VDD.n75 VDD.n74 7.5
R146 VDD.n81 VDD.n71 7.5
R147 VDD.n81 VDD.n69 7.5
R148 VDD.n84 VDD.n83 7.5
R149 VDD.n20 VDD.n16 7.5
R150 VDD.n2 VDD.n1 7.5
R151 VDD.n7 VDD.n6 7.5
R152 VDD.n10 VDD.n9 7.5
R153 VDD.n19 VDD.n18 7.5
R154 VDD.n14 VDD.n0 7.5
R155 VDD.n82 VDD.n68 6.772
R156 VDD.n80 VDD.n77 6.772
R157 VDD.n76 VDD.n73 6.772
R158 VDD.n76 VDD.n75 6.772
R159 VDD.n80 VDD.n79 6.772
R160 VDD.n83 VDD.n82 6.772
R161 VDD.n61 VDD.n60 6.772
R162 VDD.n48 VDD.n45 6.772
R163 VDD.n53 VDD.n50 6.772
R164 VDD.n58 VDD.n55 6.772
R165 VDD.n58 VDD.n57 6.772
R166 VDD.n53 VDD.n52 6.772
R167 VDD.n48 VDD.n47 6.772
R168 VDD.n60 VDD.n44 6.772
R169 VDD.n16 VDD.n15 6.458
R170 VDD.n71 VDD.n70 6.202
R171 VDD.n28 VDD.n24 1.967
R172 VDD.n38 VDD.n34 1.967
R173 VDD.n103 VDD.n99 1.967
R174 VDD.n93 VDD.n92 1.967
R175 VDD.n14 VDD.n5 1.329
R176 VDD.n14 VDD.n8 1.329
R177 VDD.n14 VDD.n11 1.329
R178 VDD.n14 VDD.n13 1.329
R179 VDD.n15 VDD.n14 0.696
R180 VDD.n14 VDD.n4 0.696
R181 VDD.n81 VDD.n80 0.365
R182 VDD.n81 VDD.n76 0.365
R183 VDD.n82 VDD.n81 0.365
R184 VDD.n59 VDD.n58 0.365
R185 VDD.n59 VDD.n53 0.365
R186 VDD.n59 VDD.n48 0.365
R187 VDD.n60 VDD.n59 0.365
R188 VDD.n88 VDD 0.207
R189 VDD.n33 VDD.n29 0.157
R190 VDD.n39 VDD.n33 0.157
R191 VDD.n104 VDD.n98 0.157
R192 VDD.n98 VDD.n94 0.157
R193 VDD.n65 VDD.n39 0.145
R194 VDD VDD.n65 0.145
R195 VDD VDD.n109 0.145
R196 VDD.n109 VDD.n104 0.145
R197 VDD.n94 VDD.n88 0.145
R198 Y.n2 Y.n1 200.754
R199 Y.n2 Y.n0 184.007
R200 Y.n3 Y.n2 76
R201 Y.n0 Y.t1 14.282
R202 Y.n0 Y.t0 14.282
R203 Y.n3 Y 0.046
C2 VDD GND 4.29fF
C3 Y.n0 GND 0.80fF
C4 Y.n1 GND 0.37fF
C5 Y.n2 GND 0.50fF
C6 Y.n3 GND 0.01fF
C7 VDD.n0 GND 0.10fF
C8 VDD.n1 GND 0.02fF
C9 VDD.n2 GND 0.02fF
C10 VDD.n3 GND 0.04fF
C11 VDD.n4 GND 0.01fF
C12 VDD.n6 GND 0.02fF
C13 VDD.n7 GND 0.02fF
C14 VDD.n9 GND 0.02fF
C15 VDD.n10 GND 0.02fF
C16 VDD.n12 GND 0.02fF
C17 VDD.n14 GND 0.40fF
C18 VDD.n16 GND 0.03fF
C19 VDD.n17 GND 0.02fF
C20 VDD.n18 GND 0.02fF
C21 VDD.n19 GND 0.02fF
C22 VDD.n20 GND 0.03fF
C23 VDD.n21 GND 0.24fF
C24 VDD.n22 GND 0.02fF
C25 VDD.n23 GND 0.03fF
C26 VDD.n24 GND 0.05fF
C27 VDD.n25 GND 0.13fF
C28 VDD.n26 GND 0.18fF
C29 VDD.n27 GND 0.01fF
C30 VDD.n28 GND 0.01fF
C31 VDD.n29 GND 0.06fF
C32 VDD.n30 GND 0.15fF
C33 VDD.n31 GND 0.01fF
C34 VDD.n32 GND 0.02fF
C35 VDD.n33 GND 0.02fF
C36 VDD.n34 GND 0.05fF
C37 VDD.n35 GND 0.13fF
C38 VDD.n36 GND 0.18fF
C39 VDD.n37 GND 0.01fF
C40 VDD.n38 GND 0.01fF
C41 VDD.n39 GND 0.02fF
C42 VDD.n40 GND 0.24fF
C43 VDD.n41 GND 0.01fF
C44 VDD.n42 GND 0.02fF
C45 VDD.n43 GND 0.02fF
C46 VDD.n44 GND 0.02fF
C47 VDD.n45 GND 0.02fF
C48 VDD.n46 GND 0.02fF
C49 VDD.n47 GND 0.02fF
C50 VDD.n49 GND 0.02fF
C51 VDD.n50 GND 0.02fF
C52 VDD.n51 GND 0.02fF
C53 VDD.n52 GND 0.02fF
C54 VDD.n54 GND 0.03fF
C55 VDD.n55 GND 0.02fF
C56 VDD.n56 GND 0.13fF
C57 VDD.n57 GND 0.03fF
C58 VDD.n59 GND 0.24fF
C59 VDD.n61 GND 0.02fF
C60 VDD.n62 GND 0.02fF
C61 VDD.n63 GND 0.03fF
C62 VDD.n64 GND 0.02fF
C63 VDD.n65 GND 0.02fF
C64 VDD.n66 GND 0.02fF
C65 VDD.n67 GND 0.02fF
C66 VDD.n68 GND 0.02fF
C67 VDD.n69 GND 0.10fF
C68 VDD.n70 GND 0.03fF
C69 VDD.n71 GND 0.02fF
C70 VDD.n72 GND 0.02fF
C71 VDD.n73 GND 0.02fF
C72 VDD.n74 GND 0.02fF
C73 VDD.n75 GND 0.02fF
C74 VDD.n77 GND 0.02fF
C75 VDD.n78 GND 0.02fF
C76 VDD.n79 GND 0.02fF
C77 VDD.n81 GND 0.40fF
C78 VDD.n83 GND 0.03fF
C79 VDD.n84 GND 0.03fF
C80 VDD.n85 GND 0.24fF
C81 VDD.n86 GND 0.02fF
C82 VDD.n87 GND 0.03fF
C83 VDD.n88 GND 0.02fF
C84 VDD.n89 GND 0.13fF
C85 VDD.n90 GND 0.18fF
C86 VDD.n91 GND 0.01fF
C87 VDD.n92 GND 0.05fF
C88 VDD.n93 GND 0.01fF
C89 VDD.n94 GND 0.02fF
C90 VDD.n95 GND 0.15fF
C91 VDD.n96 GND 0.01fF
C92 VDD.n97 GND 0.02fF
C93 VDD.n98 GND 0.02fF
C94 VDD.n99 GND 0.05fF
C95 VDD.n100 GND 0.13fF
C96 VDD.n101 GND 0.18fF
C97 VDD.n102 GND 0.01fF
C98 VDD.n103 GND 0.01fF
C99 VDD.n104 GND 0.02fF
C100 VDD.n105 GND 0.02fF
C101 VDD.n106 GND 0.24fF
C102 VDD.n107 GND 0.01fF
C103 VDD.n108 GND 0.02fF
C104 VDD.n109 GND 0.02fF
C105 a_185_209.n0 GND 0.67fF
C106 a_185_209.n1 GND 0.36fF
C107 a_185_209.n2 GND 0.47fF
C108 a_185_209.n3 GND 0.49fF
C109 a_185_209.n4 GND 0.07fF
C110 a_185_209.n5 GND 0.15fF
C111 a_185_209.n6 GND 0.04fF
.ends
