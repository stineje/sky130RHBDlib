* SPICE3 file created from DFFQX1.ext - technology: sky130A

.subckt DFFQX1 Q D CLK VDD GND
X0 GND dffx1_pcell_0/m1_2165_649# dffx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 ad=1.0746e+12p pd=9.42e+06u as=0p ps=0u w=3.01e+06u l=150000u
X1 dffx1_pcell_0/m1_258_797# CLK dffx1_pcell_0/nand2x1_pcell_2/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X2 VDD dffx1_pcell_0/m1_2165_649# dffx1_pcell_0/m1_258_797# VDD sky130_fd_pr__pfet_01v8 ad=1.58435e+13p pd=8.669e+07u as=-0p ps=0u w=2e+06u l=150000u M=2
X3 VDD CLK dffx1_pcell_0/m1_258_797# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=2e+06u l=150000u M=2
X4 GND dffx1_pcell_0/m1_833_723# dffx1_pcell_0/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X5 m1_3531_649# Q dffx1_pcell_0/nand2x1_pcell_3/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X6 VDD dffx1_pcell_0/m1_833_723# m1_3531_649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=2e+06u l=150000u M=2
X7 VDD Q m1_3531_649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=2e+06u l=150000u M=2
X8 GND m1_3531_649# dffx1_pcell_0/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X9 Q dffx1_pcell_0/m1_258_797# dffx1_pcell_0/nand2x1_pcell_4/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 ad=1.791e+11p pd=1.57e+06u as=0p ps=0u w=3.01e+06u l=150000u
X10 VDD m1_3531_649# Q VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-5.7875e+10p ps=9.165e+06u w=2e+06u l=150000u M=2
X11 VDD dffx1_pcell_0/m1_258_797# Q VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=2e+06u l=150000u M=2
X12 GND dffx1_pcell_0/m1_258_797# dffx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X13 dffx1_pcell_0/m1_833_723# dffx1_pcell_0/m1_685_649# dffx1_pcell_0/nand3x1_pcell_0/li_393_182# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X14 dffx1_pcell_0/nand3x1_pcell_0/li_393_182# CLK dffx1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X15 VDD dffx1_pcell_0/m1_258_797# dffx1_pcell_0/m1_833_723# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=2e+06u l=150000u M=2
X16 VDD CLK dffx1_pcell_0/m1_833_723# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=2e+06u l=150000u M=2
X17 VDD dffx1_pcell_0/m1_685_649# dffx1_pcell_0/m1_833_723# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=2e+06u l=150000u M=2
X18 GND dffx1_pcell_0/m1_833_723# dffx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X19 dffx1_pcell_0/m1_685_649# D dffx1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X20 VDD dffx1_pcell_0/m1_833_723# dffx1_pcell_0/m1_685_649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=2e+06u l=150000u M=2
X21 VDD D dffx1_pcell_0/m1_685_649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=2e+06u l=150000u M=2
X22 GND dffx1_pcell_0/m1_685_649# dffx1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X23 dffx1_pcell_0/m1_2165_649# dffx1_pcell_0/m1_258_797# dffx1_pcell_0/nand2x1_pcell_1/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X24 VDD dffx1_pcell_0/m1_685_649# dffx1_pcell_0/m1_2165_649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=2e+06u l=150000u M=2
X25 VDD dffx1_pcell_0/m1_258_797# dffx1_pcell_0/m1_2165_649# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=2e+06u l=150000u M=2
C0 dffx1_pcell_0/m1_258_797# VDD 3.17fF
C1 VDD dffx1_pcell_0/m1_833_723# 2.30fF
C2 dffx1_pcell_0/m1_258_797# CLK 2.96fF
C3 dffx1_pcell_0/m1_258_797# dffx1_pcell_0/m1_833_723# 3.01fF
.ends
