* SPICE3 file created from INVX1.ext - technology: sky130A

.subckt INVX1 Y A VPB VNB
M1000 VPB.t1 a_121_384# a_185_182.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_185_182.t0 a_121_384# VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u

R0 a_185_182.n3 a_185_182.n1 355.848
R1 a_185_182.n3 a_185_182.n2 30
R2 a_185_182.n4 a_185_182.n0 24.383
R3 a_185_182.n4 a_185_182.n3 23.684
R4 a_185_182.n1 a_185_182.t2 14.282
R5 a_185_182.n1 a_185_182.t0 14.282
R6 VPB VPB.n62 126.832
R7 VPB.n52 VPB.n51 76
R8 VPB.n44 VPB.n15 76
R9 VPB.n55 VPB.n54 76
R10 VPB.n46 VPB.n45 68.979
R11 VPB.n42 VPB.n41 64.528
R12 VPB.n14 VPB.t0 55.106
R13 VPB.n40 VPB.t1 55.106
R14 VPB.n59 VPB.n55 20.452
R15 VPB.n39 VPB.n36 20.452
R16 VPB.n39 VPB.n38 13.653
R17 VPB.n38 VPB.n37 13.653
R18 VPB.n44 VPB.n43 13.653
R19 VPB.n43 VPB.n42 13.653
R20 VPB.n51 VPB.n50 13.653
R21 VPB.n50 VPB.n49 13.653
R22 VPB.n48 VPB.n47 13.653
R23 VPB.n47 VPB.n46 13.653
R24 VPB.n55 VPB.n0 13.653
R25 VPB VPB.n0 13.653
R26 VPB.n59 VPB.n58 13.276
R27 VPB.n58 VPB.n56 13.276
R28 VPB.n51 VPB.n44 13.276
R29 VPB.n51 VPB.n48 13.276
R30 VPB.n36 VPB.n18 13.276
R31 VPB.n18 VPB.n16 13.276
R32 VPB.n23 VPB.n21 12.796
R33 VPB.n23 VPB.n22 12.564
R34 VPB.n31 VPB.n30 12.198
R35 VPB.n27 VPB.n26 12.198
R36 VPB.n31 VPB.n28 12.198
R37 VPB.n55 VPB.n14 10.944
R38 VPB.n40 VPB.n39 10.585
R39 VPB.n36 VPB.n35 7.5
R40 VPB.n21 VPB.n20 7.5
R41 VPB.n26 VPB.n25 7.5
R42 VPB.n30 VPB.n29 7.5
R43 VPB.n18 VPB.n17 7.5
R44 VPB.n33 VPB.n19 7.5
R45 VPB.n58 VPB.n57 7.5
R46 VPB.n12 VPB.n11 7.5
R47 VPB.n6 VPB.n5 7.5
R48 VPB.n8 VPB.n7 7.5
R49 VPB.n2 VPB.n1 7.5
R50 VPB.n60 VPB.n59 7.5
R51 VPB.n13 VPB.n10 6.729
R52 VPB.n9 VPB.n6 6.729
R53 VPB.n4 VPB.n2 6.729
R54 VPB.n4 VPB.n3 6.728
R55 VPB.n9 VPB.n8 6.728
R56 VPB.n13 VPB.n12 6.728
R57 VPB.n61 VPB.n60 6.728
R58 VPB.n35 VPB.n34 6.398
R59 VPB.n44 VPB.n40 2.691
R60 VPB.n48 VPB.n14 2.332
R61 VPB.n33 VPB.n24 1.402
R62 VPB.n33 VPB.n27 1.402
R63 VPB.n33 VPB.n31 1.402
R64 VPB.n33 VPB.n32 1.402
R65 VPB.n34 VPB.n33 0.735
R66 VPB.n33 VPB.n23 0.735
R67 VPB.n62 VPB.n13 0.387
R68 VPB.n62 VPB.n9 0.387
R69 VPB.n62 VPB.n4 0.387
R70 VPB.n62 VPB.n61 0.387
R71 VPB.n54 VPB 0.198
R72 VPB.n52 VPB.n15 0.136
R73 VPB.n53 VPB.n52 0.136
R74 VPB.n54 VPB.n53 0.136
R75 VNB VNB.n62 300.778
R76 VNB.n38 VNB.n11 76
R77 VNB.n46 VNB.n45 76
R78 VNB.n49 VNB.n48 76
R79 VNB.n44 VNB.n43 49.896
R80 VNB.n16 VNB.n15 35.01
R81 VNB.t0 VNB.n6 32.601
R82 VNB.n34 VNB.n31 20.452
R83 VNB.n50 VNB.n49 20.452
R84 VNB.n35 VNB.n16 20.094
R85 VNB.n39 VNB.n13 20.094
R86 VNB.n10 VNB.n9 20.094
R87 VNB.n16 VNB.n14 19.017
R88 VNB.n8 VNB.t0 17.353
R89 VNB.n38 VNB.n37 13.653
R90 VNB.n37 VNB.n36 13.653
R91 VNB.n45 VNB.n44 13.653
R92 VNB.n42 VNB.n41 13.653
R93 VNB.n41 VNB.n40 13.653
R94 VNB.n49 VNB.n0 13.653
R95 VNB VNB.n0 13.653
R96 VNB.n34 VNB.n33 13.653
R97 VNB.n33 VNB.n32 13.653
R98 VNB.n57 VNB.n54 13.577
R99 VNB.n19 VNB.n17 13.276
R100 VNB.n31 VNB.n19 13.276
R101 VNB.n45 VNB.n42 13.276
R102 VNB.n3 VNB.n1 13.276
R103 VNB.n50 VNB.n3 13.276
R104 VNB.n39 VNB.n38 13.097
R105 VNB.n9 VNB.n8 12.837
R106 VNB.n49 VNB.n10 9.329
R107 VNB.n35 VNB.n34 8.97
R108 VNB.n8 VNB.n7 7.566
R109 VNB.n59 VNB.n58 7.5
R110 VNB.n51 VNB.n50 7.5
R111 VNB.n3 VNB.n2 7.5
R112 VNB.n56 VNB.n55 7.5
R113 VNB.n25 VNB.n24 7.5
R114 VNB.n21 VNB.n20 7.5
R115 VNB.n19 VNB.n18 7.5
R116 VNB.n31 VNB.n30 7.5
R117 VNB.n61 VNB.n59 7.011
R118 VNB.n27 VNB.n25 7.011
R119 VNB.n23 VNB.n21 7.011
R120 VNB.n30 VNB.n29 7.01
R121 VNB.n23 VNB.n22 7.01
R122 VNB.n27 VNB.n26 7.01
R123 VNB.n61 VNB.n60 7.01
R124 VNB.n57 VNB.n56 6.788
R125 VNB.n52 VNB.n51 6.788
R126 VNB.n5 VNB.n4 4.551
R127 VNB.n38 VNB.n35 4.305
R128 VNB.n42 VNB.n10 3.947
R129 VNB.t0 VNB.n5 2.238
R130 VNB.n62 VNB.n53 0.921
R131 VNB.n62 VNB.n57 0.476
R132 VNB.n62 VNB.n52 0.475
R133 VNB.n13 VNB.n12 0.358
R134 VNB.n28 VNB.n23 0.246
R135 VNB.n29 VNB.n28 0.246
R136 VNB.n28 VNB.n27 0.246
R137 VNB.n62 VNB.n61 0.246
R138 VNB.n48 VNB 0.198
R139 VNB.n45 VNB.n39 0.179
R140 VNB.n46 VNB.n11 0.136
R141 VNB.n47 VNB.n46 0.136
R142 VNB.n48 VNB.n47 0.136




























































.ends
