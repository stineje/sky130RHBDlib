magic
tech sky130A
magscale 1 2
timestamp 1669201007
<< nwell >>
rect -87 786 2529 1550
<< pwell >>
rect -34 -34 2476 544
<< nmos >>
rect 155 297 185 350
tri 185 297 201 313 sw
rect 155 267 261 297
tri 261 267 291 297 sw
rect 155 166 185 267
tri 185 251 201 267 nw
tri 245 251 261 267 ne
tri 185 166 201 182 sw
tri 245 166 261 182 se
rect 261 166 291 267
tri 155 136 185 166 ne
rect 185 136 261 166
tri 261 136 291 166 nw
rect 612 288 642 349
tri 642 288 658 304 sw
rect 806 296 836 349
tri 836 296 852 312 sw
rect 612 258 718 288
tri 718 258 748 288 sw
rect 806 266 912 296
tri 912 266 942 296 sw
rect 612 157 642 258
tri 642 242 658 258 nw
tri 702 242 718 258 ne
tri 642 157 658 173 sw
tri 702 157 718 173 se
rect 718 157 748 258
rect 806 165 836 266
tri 836 250 852 266 nw
tri 896 250 912 266 ne
tri 836 165 852 181 sw
tri 896 165 912 181 se
rect 912 165 942 266
tri 612 127 642 157 ne
rect 642 127 718 157
tri 718 127 748 157 nw
tri 806 135 836 165 ne
rect 836 135 912 165
tri 912 135 942 165 nw
rect 1278 288 1308 349
tri 1308 288 1324 304 sw
rect 1472 296 1502 349
tri 1502 296 1518 312 sw
rect 1278 258 1384 288
tri 1384 258 1414 288 sw
rect 1472 266 1578 296
tri 1578 266 1608 296 sw
rect 1278 157 1308 258
tri 1308 242 1324 258 nw
tri 1368 242 1384 258 ne
tri 1308 157 1324 173 sw
tri 1368 157 1384 173 se
rect 1384 157 1414 258
rect 1472 165 1502 266
tri 1502 250 1518 266 nw
tri 1562 250 1578 266 ne
tri 1502 165 1518 181 sw
tri 1562 165 1578 181 se
rect 1578 165 1608 266
tri 1278 127 1308 157 ne
rect 1308 127 1384 157
tri 1384 127 1414 157 nw
tri 1472 135 1502 165 ne
rect 1502 135 1578 165
tri 1578 135 1608 165 nw
rect 1944 288 1974 349
tri 1974 288 1990 304 sw
rect 2138 296 2168 349
tri 2168 296 2184 312 sw
rect 1944 258 2050 288
tri 2050 258 2080 288 sw
rect 2138 266 2244 296
tri 2244 266 2274 296 sw
rect 1944 157 1974 258
tri 1974 242 1990 258 nw
tri 2034 242 2050 258 ne
tri 1974 157 1990 173 sw
tri 2034 157 2050 173 se
rect 2050 157 2080 258
rect 2138 165 2168 266
tri 2168 250 2184 266 nw
tri 2228 250 2244 266 ne
tri 2168 165 2184 181 sw
tri 2228 165 2244 181 se
rect 2244 165 2274 266
tri 1944 127 1974 157 ne
rect 1974 127 2050 157
tri 2050 127 2080 157 nw
tri 2138 135 2168 165 ne
rect 2168 135 2244 165
tri 2244 135 2274 165 nw
<< pmos >>
rect 164 1004 194 1404
rect 252 1004 282 1404
rect 631 1004 661 1404
rect 719 1004 749 1404
rect 807 1004 837 1404
rect 895 1004 925 1404
rect 1297 1004 1327 1404
rect 1385 1004 1415 1404
rect 1473 1004 1503 1404
rect 1561 1004 1591 1404
rect 1963 1004 1993 1404
rect 2051 1004 2081 1404
rect 2139 1004 2169 1404
rect 2227 1004 2257 1404
<< ndiff >>
rect 99 334 155 350
rect 99 300 109 334
rect 143 300 155 334
rect 99 262 155 300
rect 185 334 345 350
rect 185 313 303 334
tri 185 297 201 313 ne
rect 201 300 303 313
rect 337 300 345 334
rect 201 297 345 300
tri 261 267 291 297 ne
rect 99 228 109 262
rect 143 228 155 262
rect 99 194 155 228
rect 99 160 109 194
rect 143 160 155 194
tri 185 251 201 267 se
rect 201 251 245 267
tri 245 251 261 267 sw
rect 185 218 261 251
rect 185 184 205 218
rect 239 184 261 218
rect 185 182 261 184
tri 185 166 201 182 ne
rect 201 166 245 182
tri 245 166 261 182 nw
rect 291 262 345 297
rect 291 228 303 262
rect 337 228 345 262
rect 291 194 345 228
rect 99 136 155 160
tri 155 136 185 166 sw
tri 261 136 291 166 se
rect 291 160 303 194
rect 337 160 345 194
rect 291 136 345 160
rect 99 124 345 136
rect 99 90 109 124
rect 143 90 205 124
rect 239 90 303 124
rect 337 90 345 124
rect 99 74 345 90
rect 556 333 612 349
rect 556 299 566 333
rect 600 299 612 333
rect 556 261 612 299
rect 642 333 806 349
rect 642 304 663 333
tri 642 288 658 304 ne
rect 658 299 663 304
rect 697 299 760 333
rect 794 299 806 333
rect 658 288 806 299
rect 836 312 998 349
tri 836 296 852 312 ne
rect 852 296 998 312
rect 556 227 566 261
rect 600 227 612 261
tri 718 258 748 288 ne
rect 748 261 806 288
tri 912 266 942 296 ne
rect 556 193 612 227
rect 556 159 566 193
rect 600 159 612 193
rect 556 127 612 159
tri 642 242 658 258 se
rect 658 242 702 258
tri 702 242 718 258 sw
rect 642 208 718 242
rect 642 174 663 208
rect 697 174 718 208
rect 642 173 718 174
tri 642 157 658 173 ne
rect 658 157 702 173
tri 702 157 718 173 nw
rect 748 227 760 261
rect 794 227 806 261
rect 748 193 806 227
rect 748 159 760 193
rect 794 159 806 193
tri 836 250 852 266 se
rect 852 250 896 266
tri 896 250 912 266 sw
rect 836 217 912 250
rect 836 183 857 217
rect 891 183 912 217
rect 836 181 912 183
tri 836 165 852 181 ne
rect 852 165 896 181
tri 896 165 912 181 nw
rect 942 261 998 296
rect 942 227 954 261
rect 988 227 998 261
rect 942 193 998 227
tri 612 127 642 157 sw
tri 718 127 748 157 se
rect 748 135 806 159
tri 806 135 836 165 sw
tri 912 135 942 165 se
rect 942 159 954 193
rect 988 159 998 193
rect 942 135 998 159
rect 748 127 998 135
rect 556 123 998 127
rect 556 89 566 123
rect 600 89 760 123
rect 794 89 857 123
rect 891 89 954 123
rect 988 89 998 123
rect 556 73 998 89
rect 1222 333 1278 349
rect 1222 299 1232 333
rect 1266 299 1278 333
rect 1222 261 1278 299
rect 1308 333 1472 349
rect 1308 304 1329 333
tri 1308 288 1324 304 ne
rect 1324 299 1329 304
rect 1363 299 1426 333
rect 1460 299 1472 333
rect 1324 288 1472 299
rect 1502 312 1664 349
tri 1502 296 1518 312 ne
rect 1518 296 1664 312
rect 1222 227 1232 261
rect 1266 227 1278 261
tri 1384 258 1414 288 ne
rect 1414 261 1472 288
tri 1578 266 1608 296 ne
rect 1222 193 1278 227
rect 1222 159 1232 193
rect 1266 159 1278 193
rect 1222 127 1278 159
tri 1308 242 1324 258 se
rect 1324 242 1368 258
tri 1368 242 1384 258 sw
rect 1308 208 1384 242
rect 1308 174 1329 208
rect 1363 174 1384 208
rect 1308 173 1384 174
tri 1308 157 1324 173 ne
rect 1324 157 1368 173
tri 1368 157 1384 173 nw
rect 1414 227 1426 261
rect 1460 227 1472 261
rect 1414 193 1472 227
rect 1414 159 1426 193
rect 1460 159 1472 193
tri 1502 250 1518 266 se
rect 1518 250 1562 266
tri 1562 250 1578 266 sw
rect 1502 217 1578 250
rect 1502 183 1523 217
rect 1557 183 1578 217
rect 1502 181 1578 183
tri 1502 165 1518 181 ne
rect 1518 165 1562 181
tri 1562 165 1578 181 nw
rect 1608 261 1664 296
rect 1608 227 1620 261
rect 1654 227 1664 261
rect 1608 193 1664 227
tri 1278 127 1308 157 sw
tri 1384 127 1414 157 se
rect 1414 135 1472 159
tri 1472 135 1502 165 sw
tri 1578 135 1608 165 se
rect 1608 159 1620 193
rect 1654 159 1664 193
rect 1608 135 1664 159
rect 1414 127 1664 135
rect 1222 123 1664 127
rect 1222 89 1232 123
rect 1266 89 1426 123
rect 1460 89 1523 123
rect 1557 89 1620 123
rect 1654 89 1664 123
rect 1222 73 1664 89
rect 1888 333 1944 349
rect 1888 299 1898 333
rect 1932 299 1944 333
rect 1888 261 1944 299
rect 1974 333 2138 349
rect 1974 304 1995 333
tri 1974 288 1990 304 ne
rect 1990 299 1995 304
rect 2029 299 2092 333
rect 2126 299 2138 333
rect 1990 288 2138 299
rect 2168 312 2330 349
tri 2168 296 2184 312 ne
rect 2184 296 2330 312
rect 1888 227 1898 261
rect 1932 227 1944 261
tri 2050 258 2080 288 ne
rect 2080 261 2138 288
tri 2244 266 2274 296 ne
rect 1888 193 1944 227
rect 1888 159 1898 193
rect 1932 159 1944 193
rect 1888 127 1944 159
tri 1974 242 1990 258 se
rect 1990 242 2034 258
tri 2034 242 2050 258 sw
rect 1974 208 2050 242
rect 1974 174 1995 208
rect 2029 174 2050 208
rect 1974 173 2050 174
tri 1974 157 1990 173 ne
rect 1990 157 2034 173
tri 2034 157 2050 173 nw
rect 2080 227 2092 261
rect 2126 227 2138 261
rect 2080 193 2138 227
rect 2080 159 2092 193
rect 2126 159 2138 193
tri 2168 250 2184 266 se
rect 2184 250 2228 266
tri 2228 250 2244 266 sw
rect 2168 217 2244 250
rect 2168 183 2189 217
rect 2223 183 2244 217
rect 2168 181 2244 183
tri 2168 165 2184 181 ne
rect 2184 165 2228 181
tri 2228 165 2244 181 nw
rect 2274 261 2330 296
rect 2274 227 2286 261
rect 2320 227 2330 261
rect 2274 193 2330 227
tri 1944 127 1974 157 sw
tri 2050 127 2080 157 se
rect 2080 135 2138 159
tri 2138 135 2168 165 sw
tri 2244 135 2274 165 se
rect 2274 159 2286 193
rect 2320 159 2330 193
rect 2274 135 2330 159
rect 2080 127 2330 135
rect 1888 123 2330 127
rect 1888 89 1898 123
rect 1932 89 2092 123
rect 2126 89 2189 123
rect 2223 89 2286 123
rect 2320 89 2330 123
rect 1888 73 2330 89
<< pdiff >>
rect 108 1366 164 1404
rect 108 1332 118 1366
rect 152 1332 164 1366
rect 108 1298 164 1332
rect 108 1264 118 1298
rect 152 1264 164 1298
rect 108 1230 164 1264
rect 108 1196 118 1230
rect 152 1196 164 1230
rect 108 1162 164 1196
rect 108 1128 118 1162
rect 152 1128 164 1162
rect 108 1093 164 1128
rect 108 1059 118 1093
rect 152 1059 164 1093
rect 108 1004 164 1059
rect 194 1366 252 1404
rect 194 1332 206 1366
rect 240 1332 252 1366
rect 194 1298 252 1332
rect 194 1264 206 1298
rect 240 1264 252 1298
rect 194 1230 252 1264
rect 194 1196 206 1230
rect 240 1196 252 1230
rect 194 1162 252 1196
rect 194 1128 206 1162
rect 240 1128 252 1162
rect 194 1093 252 1128
rect 194 1059 206 1093
rect 240 1059 252 1093
rect 194 1004 252 1059
rect 282 1366 336 1404
rect 282 1332 294 1366
rect 328 1332 336 1366
rect 282 1298 336 1332
rect 282 1264 294 1298
rect 328 1264 336 1298
rect 282 1230 336 1264
rect 282 1196 294 1230
rect 328 1196 336 1230
rect 282 1162 336 1196
rect 282 1128 294 1162
rect 328 1128 336 1162
rect 282 1093 336 1128
rect 282 1059 294 1093
rect 328 1059 336 1093
rect 282 1004 336 1059
rect 575 1366 631 1404
rect 575 1332 585 1366
rect 619 1332 631 1366
rect 575 1298 631 1332
rect 575 1264 585 1298
rect 619 1264 631 1298
rect 575 1230 631 1264
rect 575 1196 585 1230
rect 619 1196 631 1230
rect 575 1162 631 1196
rect 575 1128 585 1162
rect 619 1128 631 1162
rect 575 1093 631 1128
rect 575 1059 585 1093
rect 619 1059 631 1093
rect 575 1004 631 1059
rect 661 1366 719 1404
rect 661 1332 673 1366
rect 707 1332 719 1366
rect 661 1298 719 1332
rect 661 1264 673 1298
rect 707 1264 719 1298
rect 661 1230 719 1264
rect 661 1196 673 1230
rect 707 1196 719 1230
rect 661 1162 719 1196
rect 661 1128 673 1162
rect 707 1128 719 1162
rect 661 1093 719 1128
rect 661 1059 673 1093
rect 707 1059 719 1093
rect 661 1004 719 1059
rect 749 1366 807 1404
rect 749 1332 761 1366
rect 795 1332 807 1366
rect 749 1298 807 1332
rect 749 1264 761 1298
rect 795 1264 807 1298
rect 749 1230 807 1264
rect 749 1196 761 1230
rect 795 1196 807 1230
rect 749 1162 807 1196
rect 749 1128 761 1162
rect 795 1128 807 1162
rect 749 1004 807 1128
rect 837 1366 895 1404
rect 837 1332 849 1366
rect 883 1332 895 1366
rect 837 1298 895 1332
rect 837 1264 849 1298
rect 883 1264 895 1298
rect 837 1230 895 1264
rect 837 1196 849 1230
rect 883 1196 895 1230
rect 837 1162 895 1196
rect 837 1128 849 1162
rect 883 1128 895 1162
rect 837 1093 895 1128
rect 837 1059 849 1093
rect 883 1059 895 1093
rect 837 1004 895 1059
rect 925 1366 979 1404
rect 925 1332 937 1366
rect 971 1332 979 1366
rect 925 1298 979 1332
rect 925 1264 937 1298
rect 971 1264 979 1298
rect 925 1230 979 1264
rect 925 1196 937 1230
rect 971 1196 979 1230
rect 925 1162 979 1196
rect 925 1128 937 1162
rect 971 1128 979 1162
rect 925 1004 979 1128
rect 1241 1366 1297 1404
rect 1241 1332 1251 1366
rect 1285 1332 1297 1366
rect 1241 1298 1297 1332
rect 1241 1264 1251 1298
rect 1285 1264 1297 1298
rect 1241 1230 1297 1264
rect 1241 1196 1251 1230
rect 1285 1196 1297 1230
rect 1241 1162 1297 1196
rect 1241 1128 1251 1162
rect 1285 1128 1297 1162
rect 1241 1093 1297 1128
rect 1241 1059 1251 1093
rect 1285 1059 1297 1093
rect 1241 1004 1297 1059
rect 1327 1366 1385 1404
rect 1327 1332 1339 1366
rect 1373 1332 1385 1366
rect 1327 1298 1385 1332
rect 1327 1264 1339 1298
rect 1373 1264 1385 1298
rect 1327 1230 1385 1264
rect 1327 1196 1339 1230
rect 1373 1196 1385 1230
rect 1327 1162 1385 1196
rect 1327 1128 1339 1162
rect 1373 1128 1385 1162
rect 1327 1093 1385 1128
rect 1327 1059 1339 1093
rect 1373 1059 1385 1093
rect 1327 1004 1385 1059
rect 1415 1366 1473 1404
rect 1415 1332 1427 1366
rect 1461 1332 1473 1366
rect 1415 1298 1473 1332
rect 1415 1264 1427 1298
rect 1461 1264 1473 1298
rect 1415 1230 1473 1264
rect 1415 1196 1427 1230
rect 1461 1196 1473 1230
rect 1415 1162 1473 1196
rect 1415 1128 1427 1162
rect 1461 1128 1473 1162
rect 1415 1004 1473 1128
rect 1503 1366 1561 1404
rect 1503 1332 1515 1366
rect 1549 1332 1561 1366
rect 1503 1298 1561 1332
rect 1503 1264 1515 1298
rect 1549 1264 1561 1298
rect 1503 1230 1561 1264
rect 1503 1196 1515 1230
rect 1549 1196 1561 1230
rect 1503 1162 1561 1196
rect 1503 1128 1515 1162
rect 1549 1128 1561 1162
rect 1503 1093 1561 1128
rect 1503 1059 1515 1093
rect 1549 1059 1561 1093
rect 1503 1004 1561 1059
rect 1591 1366 1645 1404
rect 1591 1332 1603 1366
rect 1637 1332 1645 1366
rect 1591 1298 1645 1332
rect 1591 1264 1603 1298
rect 1637 1264 1645 1298
rect 1591 1230 1645 1264
rect 1591 1196 1603 1230
rect 1637 1196 1645 1230
rect 1591 1162 1645 1196
rect 1591 1128 1603 1162
rect 1637 1128 1645 1162
rect 1591 1004 1645 1128
rect 1907 1366 1963 1404
rect 1907 1332 1917 1366
rect 1951 1332 1963 1366
rect 1907 1298 1963 1332
rect 1907 1264 1917 1298
rect 1951 1264 1963 1298
rect 1907 1230 1963 1264
rect 1907 1196 1917 1230
rect 1951 1196 1963 1230
rect 1907 1162 1963 1196
rect 1907 1128 1917 1162
rect 1951 1128 1963 1162
rect 1907 1093 1963 1128
rect 1907 1059 1917 1093
rect 1951 1059 1963 1093
rect 1907 1004 1963 1059
rect 1993 1366 2051 1404
rect 1993 1332 2005 1366
rect 2039 1332 2051 1366
rect 1993 1298 2051 1332
rect 1993 1264 2005 1298
rect 2039 1264 2051 1298
rect 1993 1230 2051 1264
rect 1993 1196 2005 1230
rect 2039 1196 2051 1230
rect 1993 1162 2051 1196
rect 1993 1128 2005 1162
rect 2039 1128 2051 1162
rect 1993 1093 2051 1128
rect 1993 1059 2005 1093
rect 2039 1059 2051 1093
rect 1993 1004 2051 1059
rect 2081 1366 2139 1404
rect 2081 1332 2093 1366
rect 2127 1332 2139 1366
rect 2081 1298 2139 1332
rect 2081 1264 2093 1298
rect 2127 1264 2139 1298
rect 2081 1230 2139 1264
rect 2081 1196 2093 1230
rect 2127 1196 2139 1230
rect 2081 1162 2139 1196
rect 2081 1128 2093 1162
rect 2127 1128 2139 1162
rect 2081 1004 2139 1128
rect 2169 1366 2227 1404
rect 2169 1332 2181 1366
rect 2215 1332 2227 1366
rect 2169 1298 2227 1332
rect 2169 1264 2181 1298
rect 2215 1264 2227 1298
rect 2169 1230 2227 1264
rect 2169 1196 2181 1230
rect 2215 1196 2227 1230
rect 2169 1162 2227 1196
rect 2169 1128 2181 1162
rect 2215 1128 2227 1162
rect 2169 1093 2227 1128
rect 2169 1059 2181 1093
rect 2215 1059 2227 1093
rect 2169 1004 2227 1059
rect 2257 1366 2311 1404
rect 2257 1332 2269 1366
rect 2303 1332 2311 1366
rect 2257 1298 2311 1332
rect 2257 1264 2269 1298
rect 2303 1264 2311 1298
rect 2257 1230 2311 1264
rect 2257 1196 2269 1230
rect 2303 1196 2311 1230
rect 2257 1162 2311 1196
rect 2257 1128 2269 1162
rect 2303 1128 2311 1162
rect 2257 1004 2311 1128
<< ndiffc >>
rect 109 300 143 334
rect 303 300 337 334
rect 109 228 143 262
rect 109 160 143 194
rect 205 184 239 218
rect 303 228 337 262
rect 303 160 337 194
rect 109 90 143 124
rect 205 90 239 124
rect 303 90 337 124
rect 566 299 600 333
rect 663 299 697 333
rect 760 299 794 333
rect 566 227 600 261
rect 566 159 600 193
rect 663 174 697 208
rect 760 227 794 261
rect 760 159 794 193
rect 857 183 891 217
rect 954 227 988 261
rect 954 159 988 193
rect 566 89 600 123
rect 760 89 794 123
rect 857 89 891 123
rect 954 89 988 123
rect 1232 299 1266 333
rect 1329 299 1363 333
rect 1426 299 1460 333
rect 1232 227 1266 261
rect 1232 159 1266 193
rect 1329 174 1363 208
rect 1426 227 1460 261
rect 1426 159 1460 193
rect 1523 183 1557 217
rect 1620 227 1654 261
rect 1620 159 1654 193
rect 1232 89 1266 123
rect 1426 89 1460 123
rect 1523 89 1557 123
rect 1620 89 1654 123
rect 1898 299 1932 333
rect 1995 299 2029 333
rect 2092 299 2126 333
rect 1898 227 1932 261
rect 1898 159 1932 193
rect 1995 174 2029 208
rect 2092 227 2126 261
rect 2092 159 2126 193
rect 2189 183 2223 217
rect 2286 227 2320 261
rect 2286 159 2320 193
rect 1898 89 1932 123
rect 2092 89 2126 123
rect 2189 89 2223 123
rect 2286 89 2320 123
<< pdiffc >>
rect 118 1332 152 1366
rect 118 1264 152 1298
rect 118 1196 152 1230
rect 118 1128 152 1162
rect 118 1059 152 1093
rect 206 1332 240 1366
rect 206 1264 240 1298
rect 206 1196 240 1230
rect 206 1128 240 1162
rect 206 1059 240 1093
rect 294 1332 328 1366
rect 294 1264 328 1298
rect 294 1196 328 1230
rect 294 1128 328 1162
rect 294 1059 328 1093
rect 585 1332 619 1366
rect 585 1264 619 1298
rect 585 1196 619 1230
rect 585 1128 619 1162
rect 585 1059 619 1093
rect 673 1332 707 1366
rect 673 1264 707 1298
rect 673 1196 707 1230
rect 673 1128 707 1162
rect 673 1059 707 1093
rect 761 1332 795 1366
rect 761 1264 795 1298
rect 761 1196 795 1230
rect 761 1128 795 1162
rect 849 1332 883 1366
rect 849 1264 883 1298
rect 849 1196 883 1230
rect 849 1128 883 1162
rect 849 1059 883 1093
rect 937 1332 971 1366
rect 937 1264 971 1298
rect 937 1196 971 1230
rect 937 1128 971 1162
rect 1251 1332 1285 1366
rect 1251 1264 1285 1298
rect 1251 1196 1285 1230
rect 1251 1128 1285 1162
rect 1251 1059 1285 1093
rect 1339 1332 1373 1366
rect 1339 1264 1373 1298
rect 1339 1196 1373 1230
rect 1339 1128 1373 1162
rect 1339 1059 1373 1093
rect 1427 1332 1461 1366
rect 1427 1264 1461 1298
rect 1427 1196 1461 1230
rect 1427 1128 1461 1162
rect 1515 1332 1549 1366
rect 1515 1264 1549 1298
rect 1515 1196 1549 1230
rect 1515 1128 1549 1162
rect 1515 1059 1549 1093
rect 1603 1332 1637 1366
rect 1603 1264 1637 1298
rect 1603 1196 1637 1230
rect 1603 1128 1637 1162
rect 1917 1332 1951 1366
rect 1917 1264 1951 1298
rect 1917 1196 1951 1230
rect 1917 1128 1951 1162
rect 1917 1059 1951 1093
rect 2005 1332 2039 1366
rect 2005 1264 2039 1298
rect 2005 1196 2039 1230
rect 2005 1128 2039 1162
rect 2005 1059 2039 1093
rect 2093 1332 2127 1366
rect 2093 1264 2127 1298
rect 2093 1196 2127 1230
rect 2093 1128 2127 1162
rect 2181 1332 2215 1366
rect 2181 1264 2215 1298
rect 2181 1196 2215 1230
rect 2181 1128 2215 1162
rect 2181 1059 2215 1093
rect 2269 1332 2303 1366
rect 2269 1264 2303 1298
rect 2269 1196 2303 1230
rect 2269 1128 2303 1162
<< psubdiff >>
rect -34 482 2476 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 410 461 478 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 410 427 427 461
rect 461 427 478 461
rect 1076 461 1144 482
rect -34 313 34 353
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 410 313 478 353
rect 1076 427 1093 461
rect 1127 427 1144 461
rect 1742 461 1810 482
rect 1076 387 1144 427
rect 1076 353 1093 387
rect 1127 353 1144 387
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect -34 17 34 57
rect 410 57 427 91
rect 461 57 478 91
rect 1076 313 1144 353
rect 1742 427 1759 461
rect 1793 427 1810 461
rect 2408 461 2476 482
rect 1742 387 1810 427
rect 1742 353 1759 387
rect 1793 353 1810 387
rect 1076 279 1093 313
rect 1127 279 1144 313
rect 1076 239 1144 279
rect 1076 205 1093 239
rect 1127 205 1144 239
rect 1076 165 1144 205
rect 1076 131 1093 165
rect 1127 131 1144 165
rect 1076 91 1144 131
rect 410 17 478 57
rect 1076 57 1093 91
rect 1127 57 1144 91
rect 1742 313 1810 353
rect 2408 427 2425 461
rect 2459 427 2476 461
rect 2408 387 2476 427
rect 2408 353 2425 387
rect 2459 353 2476 387
rect 1742 279 1759 313
rect 1793 279 1810 313
rect 1742 239 1810 279
rect 1742 205 1759 239
rect 1793 205 1810 239
rect 1742 165 1810 205
rect 1742 131 1759 165
rect 1793 131 1810 165
rect 1742 91 1810 131
rect 1076 17 1144 57
rect 1742 57 1759 91
rect 1793 57 1810 91
rect 2408 313 2476 353
rect 2408 279 2425 313
rect 2459 279 2476 313
rect 2408 239 2476 279
rect 2408 205 2425 239
rect 2459 205 2476 239
rect 2408 165 2476 205
rect 2408 131 2425 165
rect 2459 131 2476 165
rect 2408 91 2476 131
rect 1742 17 1810 57
rect 2408 57 2425 91
rect 2459 57 2476 91
rect 2408 17 2476 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2476 17
rect -34 -34 2476 -17
<< nsubdiff >>
rect -34 1497 2476 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2476 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 410 1423 478 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 1076 1423 1144 1463
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 410 979 478 1019
rect 1076 1389 1093 1423
rect 1127 1389 1144 1423
rect 1742 1423 1810 1463
rect 1076 1349 1144 1389
rect 1076 1315 1093 1349
rect 1127 1315 1144 1349
rect 1076 1275 1144 1315
rect 1076 1241 1093 1275
rect 1127 1241 1144 1275
rect 1076 1201 1144 1241
rect 1076 1167 1093 1201
rect 1127 1167 1144 1201
rect 1076 1127 1144 1167
rect 1076 1093 1093 1127
rect 1127 1093 1144 1127
rect 1076 1053 1144 1093
rect 1076 1019 1093 1053
rect 1127 1019 1144 1053
rect 410 945 427 979
rect 461 945 478 979
rect -34 871 -17 905
rect 17 884 34 905
rect 410 905 478 945
rect 1076 979 1144 1019
rect 1742 1389 1759 1423
rect 1793 1389 1810 1423
rect 2408 1423 2476 1463
rect 1742 1349 1810 1389
rect 1742 1315 1759 1349
rect 1793 1315 1810 1349
rect 1742 1275 1810 1315
rect 1742 1241 1759 1275
rect 1793 1241 1810 1275
rect 1742 1201 1810 1241
rect 1742 1167 1759 1201
rect 1793 1167 1810 1201
rect 1742 1127 1810 1167
rect 1742 1093 1759 1127
rect 1793 1093 1810 1127
rect 1742 1053 1810 1093
rect 1742 1019 1759 1053
rect 1793 1019 1810 1053
rect 1076 945 1093 979
rect 1127 945 1144 979
rect 410 884 427 905
rect 17 871 427 884
rect 461 884 478 905
rect 1076 905 1144 945
rect 1742 979 1810 1019
rect 2408 1389 2425 1423
rect 2459 1389 2476 1423
rect 2408 1349 2476 1389
rect 2408 1315 2425 1349
rect 2459 1315 2476 1349
rect 2408 1275 2476 1315
rect 2408 1241 2425 1275
rect 2459 1241 2476 1275
rect 2408 1201 2476 1241
rect 2408 1167 2425 1201
rect 2459 1167 2476 1201
rect 2408 1127 2476 1167
rect 2408 1093 2425 1127
rect 2459 1093 2476 1127
rect 2408 1053 2476 1093
rect 2408 1019 2425 1053
rect 2459 1019 2476 1053
rect 1742 945 1759 979
rect 1793 945 1810 979
rect 1076 884 1093 905
rect 461 871 1093 884
rect 1127 884 1144 905
rect 1742 905 1810 945
rect 2408 979 2476 1019
rect 2408 945 2425 979
rect 2459 945 2476 979
rect 1742 884 1759 905
rect 1127 871 1759 884
rect 1793 884 1810 905
rect 2408 905 2476 945
rect 2408 884 2425 905
rect 1793 871 2425 884
rect 2459 871 2476 905
rect -34 822 2476 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 427 427 461 461
rect 427 353 461 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1093 427 1127 461
rect 1093 353 1127 387
rect 427 279 461 313
rect 427 205 461 239
rect 427 131 461 165
rect 427 57 461 91
rect 1759 427 1793 461
rect 1759 353 1793 387
rect 1093 279 1127 313
rect 1093 205 1127 239
rect 1093 131 1127 165
rect 1093 57 1127 91
rect 2425 427 2459 461
rect 2425 353 2459 387
rect 1759 279 1793 313
rect 1759 205 1793 239
rect 1759 131 1793 165
rect 1759 57 1793 91
rect 2425 279 2459 313
rect 2425 205 2459 239
rect 2425 131 2459 165
rect 2425 57 2459 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 427 1389 461 1423
rect 427 1315 461 1349
rect 427 1241 461 1275
rect 427 1167 461 1201
rect 427 1093 461 1127
rect 427 1019 461 1053
rect -17 945 17 979
rect 1093 1389 1127 1423
rect 1093 1315 1127 1349
rect 1093 1241 1127 1275
rect 1093 1167 1127 1201
rect 1093 1093 1127 1127
rect 1093 1019 1127 1053
rect 427 945 461 979
rect -17 871 17 905
rect 1759 1389 1793 1423
rect 1759 1315 1793 1349
rect 1759 1241 1793 1275
rect 1759 1167 1793 1201
rect 1759 1093 1793 1127
rect 1759 1019 1793 1053
rect 1093 945 1127 979
rect 427 871 461 905
rect 2425 1389 2459 1423
rect 2425 1315 2459 1349
rect 2425 1241 2459 1275
rect 2425 1167 2459 1201
rect 2425 1093 2459 1127
rect 2425 1019 2459 1053
rect 1759 945 1793 979
rect 1093 871 1127 905
rect 2425 945 2459 979
rect 1759 871 1793 905
rect 2425 871 2459 905
<< poly >>
rect 164 1404 194 1430
rect 252 1404 282 1430
rect 631 1404 661 1430
rect 719 1404 749 1430
rect 807 1404 837 1430
rect 895 1404 925 1430
rect 164 973 194 1004
rect 252 973 282 1004
rect 121 957 282 973
rect 121 923 131 957
rect 165 943 282 957
rect 1297 1404 1327 1430
rect 1385 1404 1415 1430
rect 1473 1404 1503 1430
rect 1561 1404 1591 1430
rect 165 923 175 943
rect 121 907 175 923
rect 631 973 661 1004
rect 719 973 749 1004
rect 807 973 837 1004
rect 895 973 925 1004
rect 631 957 749 973
rect 631 943 649 957
rect 639 923 649 943
rect 683 943 749 957
rect 793 957 925 973
rect 683 923 693 943
rect 639 907 693 923
rect 793 923 803 957
rect 837 943 925 957
rect 1963 1404 1993 1430
rect 2051 1404 2081 1430
rect 2139 1404 2169 1430
rect 2227 1404 2257 1430
rect 837 923 847 943
rect 793 907 847 923
rect 1297 973 1327 1004
rect 1385 973 1415 1004
rect 1473 973 1503 1004
rect 1561 973 1591 1004
rect 1297 957 1415 973
rect 1297 943 1315 957
rect 1305 923 1315 943
rect 1349 943 1415 957
rect 1459 957 1591 973
rect 1349 923 1359 943
rect 1305 907 1359 923
rect 1459 923 1469 957
rect 1503 943 1591 957
rect 1503 923 1513 943
rect 1459 907 1513 923
rect 1963 973 1993 1004
rect 2051 973 2081 1004
rect 2139 973 2169 1004
rect 2227 973 2257 1004
rect 1963 957 2081 973
rect 1963 943 1981 957
rect 1971 923 1981 943
rect 2015 943 2081 957
rect 2125 957 2257 973
rect 2015 923 2025 943
rect 1971 907 2025 923
rect 2125 923 2135 957
rect 2169 943 2257 957
rect 2169 923 2179 943
rect 2125 907 2179 923
rect 121 434 175 450
rect 121 400 131 434
rect 165 413 175 434
rect 165 400 185 413
rect 121 384 185 400
rect 155 350 185 384
rect 639 433 693 449
rect 639 413 649 433
rect 612 399 649 413
rect 683 399 693 433
rect 612 383 693 399
rect 787 433 841 449
rect 787 399 797 433
rect 831 399 841 433
rect 787 383 841 399
rect 1305 433 1359 449
rect 1305 413 1315 433
rect 612 349 642 383
rect 806 349 836 383
rect 1278 399 1315 413
rect 1349 399 1359 433
rect 1278 383 1359 399
rect 1453 433 1507 449
rect 1453 399 1463 433
rect 1497 399 1507 433
rect 1453 383 1507 399
rect 1971 433 2025 449
rect 1971 413 1981 433
rect 1278 349 1308 383
rect 1472 349 1502 383
rect 1944 399 1981 413
rect 2015 399 2025 433
rect 1944 383 2025 399
rect 2119 433 2173 449
rect 2119 399 2129 433
rect 2163 399 2173 433
rect 2119 383 2173 399
rect 1944 349 1974 383
rect 2138 349 2168 383
<< polycont >>
rect 131 923 165 957
rect 649 923 683 957
rect 803 923 837 957
rect 1315 923 1349 957
rect 1469 923 1503 957
rect 1981 923 2015 957
rect 2135 923 2169 957
rect 131 400 165 434
rect 649 399 683 433
rect 797 399 831 433
rect 1315 399 1349 433
rect 1463 399 1497 433
rect 1981 399 2015 433
rect 2129 399 2163 433
<< locali >>
rect -34 1497 2476 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2476 1497
rect -34 1446 2476 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 118 1366 152 1446
rect 118 1298 152 1332
rect 118 1230 152 1264
rect 118 1162 152 1196
rect 118 1093 152 1128
rect 118 1037 152 1059
rect 206 1366 240 1404
rect 206 1298 240 1332
rect 206 1230 240 1264
rect 206 1162 240 1196
rect 206 1093 240 1128
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 131 957 165 973
rect 131 609 165 923
rect 206 933 240 1059
rect 294 1366 328 1446
rect 294 1298 328 1332
rect 294 1230 328 1264
rect 294 1162 328 1196
rect 294 1093 328 1128
rect 294 1037 328 1059
rect 410 1423 478 1446
rect 410 1389 427 1423
rect 461 1389 478 1423
rect 410 1349 478 1389
rect 410 1315 427 1349
rect 461 1315 478 1349
rect 410 1275 478 1315
rect 410 1241 427 1275
rect 461 1241 478 1275
rect 410 1201 478 1241
rect 410 1167 427 1201
rect 461 1167 478 1201
rect 410 1127 478 1167
rect 410 1093 427 1127
rect 461 1093 478 1127
rect 410 1053 478 1093
rect 410 1019 427 1053
rect 461 1019 478 1053
rect 585 1366 619 1446
rect 585 1298 619 1332
rect 585 1230 619 1264
rect 585 1162 619 1196
rect 585 1093 619 1128
rect 585 1027 619 1059
rect 673 1366 707 1404
rect 673 1298 707 1332
rect 673 1230 707 1264
rect 673 1162 707 1196
rect 673 1093 707 1128
rect 761 1366 795 1446
rect 761 1298 795 1332
rect 761 1230 795 1264
rect 761 1162 795 1196
rect 761 1111 795 1128
rect 849 1366 883 1404
rect 849 1298 883 1332
rect 849 1230 883 1264
rect 849 1162 883 1196
rect 673 1057 707 1059
rect 849 1093 883 1128
rect 937 1366 971 1446
rect 937 1298 971 1332
rect 937 1230 971 1264
rect 937 1162 971 1196
rect 937 1111 971 1128
rect 1076 1423 1144 1446
rect 1076 1389 1093 1423
rect 1127 1389 1144 1423
rect 1076 1349 1144 1389
rect 1076 1315 1093 1349
rect 1127 1315 1144 1349
rect 1076 1275 1144 1315
rect 1076 1241 1093 1275
rect 1127 1241 1144 1275
rect 1076 1201 1144 1241
rect 1076 1167 1093 1201
rect 1127 1167 1144 1201
rect 1076 1127 1144 1167
rect 849 1057 883 1059
rect 1076 1093 1093 1127
rect 1127 1093 1144 1127
rect 673 1023 979 1057
rect 410 979 478 1019
rect 410 945 427 979
rect 461 945 478 979
rect 206 899 313 933
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 131 434 165 575
rect 279 683 313 899
rect 410 905 478 945
rect 410 871 427 905
rect 461 871 478 905
rect 410 822 478 871
rect 649 957 683 973
rect 803 957 837 973
rect 279 433 313 649
rect 649 609 683 923
rect 131 384 165 400
rect 205 399 313 433
rect 410 461 478 544
rect 410 427 427 461
rect 461 427 478 461
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect -34 34 34 57
rect 109 334 143 350
rect 109 262 143 300
rect 109 194 143 228
rect 205 218 239 399
rect 410 387 478 427
rect 410 353 427 387
rect 461 353 478 387
rect 649 433 683 575
rect 649 383 683 399
rect 797 923 803 942
rect 797 907 837 923
rect 797 433 831 907
rect 797 383 831 399
rect 945 609 979 1023
rect 1076 1053 1144 1093
rect 1076 1019 1093 1053
rect 1127 1019 1144 1053
rect 1251 1366 1285 1446
rect 1251 1298 1285 1332
rect 1251 1230 1285 1264
rect 1251 1162 1285 1196
rect 1251 1093 1285 1128
rect 1251 1027 1285 1059
rect 1339 1366 1373 1404
rect 1339 1298 1373 1332
rect 1339 1230 1373 1264
rect 1339 1162 1373 1196
rect 1339 1093 1373 1128
rect 1427 1366 1461 1446
rect 1427 1298 1461 1332
rect 1427 1230 1461 1264
rect 1427 1162 1461 1196
rect 1427 1111 1461 1128
rect 1515 1366 1549 1404
rect 1515 1298 1549 1332
rect 1515 1230 1549 1264
rect 1515 1162 1549 1196
rect 1339 1057 1373 1059
rect 1515 1093 1549 1128
rect 1603 1366 1637 1446
rect 1603 1298 1637 1332
rect 1603 1230 1637 1264
rect 1603 1162 1637 1196
rect 1603 1111 1637 1128
rect 1742 1423 1810 1446
rect 1742 1389 1759 1423
rect 1793 1389 1810 1423
rect 1742 1349 1810 1389
rect 1742 1315 1759 1349
rect 1793 1315 1810 1349
rect 1742 1275 1810 1315
rect 1742 1241 1759 1275
rect 1793 1241 1810 1275
rect 1742 1201 1810 1241
rect 1742 1167 1759 1201
rect 1793 1167 1810 1201
rect 1742 1127 1810 1167
rect 1515 1057 1549 1059
rect 1742 1093 1759 1127
rect 1793 1093 1810 1127
rect 1339 1023 1645 1057
rect 1076 979 1144 1019
rect 1076 945 1093 979
rect 1127 945 1144 979
rect 1076 905 1144 945
rect 1076 871 1093 905
rect 1127 871 1144 905
rect 1076 822 1144 871
rect 1315 957 1349 973
rect 1469 957 1503 973
rect 205 168 239 184
rect 303 334 337 350
rect 303 262 337 300
rect 303 194 337 228
rect 109 124 143 160
rect 303 124 337 160
rect 143 90 205 124
rect 239 90 303 124
rect 109 34 143 90
rect 206 34 240 90
rect 303 34 337 90
rect 410 313 478 353
rect 410 279 427 313
rect 461 279 478 313
rect 410 239 478 279
rect 410 205 427 239
rect 461 205 478 239
rect 410 165 478 205
rect 410 131 427 165
rect 461 131 478 165
rect 410 91 478 131
rect 410 57 427 91
rect 461 57 478 91
rect 566 333 600 349
rect 760 333 794 349
rect 945 348 979 575
rect 1315 683 1349 923
rect 600 299 663 333
rect 697 299 760 333
rect 566 261 600 299
rect 566 193 600 227
rect 760 261 794 299
rect 566 123 600 159
rect 566 73 600 89
rect 663 208 697 224
rect 410 34 478 57
rect 663 34 697 174
rect 760 193 794 227
rect 857 314 979 348
rect 1076 461 1144 544
rect 1076 427 1093 461
rect 1127 427 1144 461
rect 1076 387 1144 427
rect 1076 353 1093 387
rect 1127 353 1144 387
rect 1315 433 1349 649
rect 1315 383 1349 399
rect 1463 923 1469 942
rect 1463 907 1503 923
rect 1463 433 1497 907
rect 1463 383 1497 399
rect 1611 683 1645 1023
rect 1742 1053 1810 1093
rect 1742 1019 1759 1053
rect 1793 1019 1810 1053
rect 1917 1366 1951 1446
rect 1917 1298 1951 1332
rect 1917 1230 1951 1264
rect 1917 1162 1951 1196
rect 1917 1093 1951 1128
rect 1917 1027 1951 1059
rect 2005 1366 2039 1404
rect 2005 1298 2039 1332
rect 2005 1230 2039 1264
rect 2005 1162 2039 1196
rect 2005 1093 2039 1128
rect 2093 1366 2127 1446
rect 2093 1298 2127 1332
rect 2093 1230 2127 1264
rect 2093 1162 2127 1196
rect 2093 1111 2127 1128
rect 2181 1366 2215 1404
rect 2181 1298 2215 1332
rect 2181 1230 2215 1264
rect 2181 1162 2215 1196
rect 2005 1057 2039 1059
rect 2181 1093 2215 1128
rect 2269 1366 2303 1446
rect 2269 1298 2303 1332
rect 2269 1230 2303 1264
rect 2269 1162 2303 1196
rect 2269 1111 2303 1128
rect 2408 1423 2476 1446
rect 2408 1389 2425 1423
rect 2459 1389 2476 1423
rect 2408 1349 2476 1389
rect 2408 1315 2425 1349
rect 2459 1315 2476 1349
rect 2408 1275 2476 1315
rect 2408 1241 2425 1275
rect 2459 1241 2476 1275
rect 2408 1201 2476 1241
rect 2408 1167 2425 1201
rect 2459 1167 2476 1201
rect 2408 1127 2476 1167
rect 2181 1057 2215 1059
rect 2408 1093 2425 1127
rect 2459 1093 2476 1127
rect 2005 1023 2311 1057
rect 1742 979 1810 1019
rect 1742 945 1759 979
rect 1793 945 1810 979
rect 1742 905 1810 945
rect 1742 871 1759 905
rect 1793 871 1810 905
rect 1742 822 1810 871
rect 1981 957 2015 973
rect 2135 957 2169 973
rect 857 217 891 314
rect 1076 313 1144 353
rect 1076 279 1093 313
rect 1127 279 1144 313
rect 857 167 891 183
rect 954 261 988 277
rect 954 193 988 227
rect 760 123 794 159
rect 954 123 988 159
rect 794 89 857 123
rect 891 89 954 123
rect 760 73 794 89
rect 954 73 988 89
rect 1076 239 1144 279
rect 1076 205 1093 239
rect 1127 205 1144 239
rect 1076 165 1144 205
rect 1076 131 1093 165
rect 1127 131 1144 165
rect 1076 91 1144 131
rect 1076 57 1093 91
rect 1127 57 1144 91
rect 1232 333 1266 349
rect 1426 333 1460 349
rect 1611 348 1645 649
rect 1981 609 2015 923
rect 1266 299 1329 333
rect 1363 299 1426 333
rect 1232 261 1266 299
rect 1232 193 1266 227
rect 1426 261 1460 299
rect 1232 123 1266 159
rect 1232 73 1266 89
rect 1329 208 1363 224
rect 1076 34 1144 57
rect 1329 34 1363 174
rect 1426 193 1460 227
rect 1523 314 1645 348
rect 1742 461 1810 544
rect 1742 427 1759 461
rect 1793 427 1810 461
rect 1742 387 1810 427
rect 1742 353 1759 387
rect 1793 353 1810 387
rect 1981 433 2015 575
rect 1981 383 2015 399
rect 2129 923 2135 942
rect 2129 907 2169 923
rect 2129 683 2163 907
rect 2129 433 2163 649
rect 2129 383 2163 399
rect 1523 217 1557 314
rect 1742 313 1810 353
rect 1742 279 1759 313
rect 1793 279 1810 313
rect 1523 167 1557 183
rect 1620 261 1654 277
rect 1620 193 1654 227
rect 1426 123 1460 159
rect 1620 123 1654 159
rect 1460 89 1523 123
rect 1557 89 1620 123
rect 1426 73 1460 89
rect 1620 73 1654 89
rect 1742 239 1810 279
rect 1742 205 1759 239
rect 1793 205 1810 239
rect 1742 165 1810 205
rect 1742 131 1759 165
rect 1793 131 1810 165
rect 1742 91 1810 131
rect 1742 57 1759 91
rect 1793 57 1810 91
rect 1898 333 1932 349
rect 2092 333 2126 349
rect 2277 348 2311 1023
rect 2408 1053 2476 1093
rect 2408 1019 2425 1053
rect 2459 1019 2476 1053
rect 2408 979 2476 1019
rect 2408 945 2425 979
rect 2459 945 2476 979
rect 2408 905 2476 945
rect 2408 871 2425 905
rect 2459 871 2476 905
rect 2408 822 2476 871
rect 1932 299 1995 333
rect 2029 299 2092 333
rect 1898 261 1932 299
rect 1898 193 1932 227
rect 2092 261 2126 299
rect 1898 123 1932 159
rect 1898 73 1932 89
rect 1995 208 2029 224
rect 1742 34 1810 57
rect 1995 34 2029 174
rect 2092 193 2126 227
rect 2189 314 2311 348
rect 2408 461 2476 544
rect 2408 427 2425 461
rect 2459 427 2476 461
rect 2408 387 2476 427
rect 2408 353 2425 387
rect 2459 353 2476 387
rect 2189 217 2223 314
rect 2408 313 2476 353
rect 2408 279 2425 313
rect 2459 279 2476 313
rect 2189 167 2223 183
rect 2286 261 2320 277
rect 2286 193 2320 227
rect 2092 123 2126 159
rect 2286 123 2320 159
rect 2126 89 2189 123
rect 2223 89 2286 123
rect 2092 73 2126 89
rect 2286 73 2320 89
rect 2408 239 2476 279
rect 2408 205 2425 239
rect 2459 205 2476 239
rect 2408 165 2476 205
rect 2408 131 2425 165
rect 2459 131 2476 165
rect 2408 91 2476 131
rect 2408 57 2425 91
rect 2459 57 2476 91
rect 2408 34 2476 57
rect -34 17 2476 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2476 17
rect -34 -34 2476 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 649 1463 683 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1611 1463 1645 1497
rect 1685 1463 1719 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 131 575 165 609
rect 279 649 313 683
rect 649 575 683 609
rect 945 575 979 609
rect 1315 649 1349 683
rect 1611 649 1645 683
rect 1981 575 2015 609
rect 2129 649 2163 683
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 649 -17 683 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1611 -17 1645 17
rect 1685 -17 1719 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
<< metal1 >>
rect -34 1497 2476 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 649 1497
rect 683 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1611 1497
rect 1645 1463 1685 1497
rect 1719 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2476 1497
rect -34 1446 2476 1463
rect 273 683 319 689
rect 1309 683 1355 689
rect 1605 683 1651 689
rect 2123 683 2169 689
rect 267 649 279 683
rect 313 649 1315 683
rect 1349 649 1361 683
rect 1599 649 1611 683
rect 1645 649 2129 683
rect 2163 649 2175 683
rect 273 643 319 649
rect 1309 643 1355 649
rect 1605 643 1651 649
rect 2123 643 2169 649
rect 125 609 171 615
rect 643 609 689 615
rect 939 609 985 615
rect 1975 609 2021 615
rect 119 575 131 609
rect 165 575 649 609
rect 683 575 695 609
rect 933 575 945 609
rect 979 575 1981 609
rect 2015 575 2027 609
rect 125 569 171 575
rect 643 569 689 575
rect 939 569 985 575
rect 1975 569 2021 575
rect -34 17 2476 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 501 17
rect 535 -17 575 17
rect 609 -17 649 17
rect 683 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1611 17
rect 1645 -17 1685 17
rect 1719 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2476 17
rect -34 -34 2476 -17
<< labels >>
rlabel metal1 2277 649 2311 683 1 Y
port 1 n
rlabel metal1 2277 723 2311 757 1 Y
port 2 n
rlabel metal1 2277 797 2311 831 1 Y
port 3 n
rlabel metal1 2277 871 2311 905 1 Y
port 4 n
rlabel metal1 2277 945 2311 979 1 Y
port 5 n
rlabel metal1 2277 575 2311 609 1 Y
port 6 n
rlabel metal1 2277 501 2311 535 1 Y
port 7 n
rlabel metal1 2277 427 2311 461 1 Y
port 8 n
rlabel metal1 797 723 831 757 1 A0
port 9 n
rlabel metal1 797 797 831 831 1 A0
port 10 n
rlabel metal1 797 871 831 905 1 A0
port 11 n
rlabel metal1 797 575 831 609 1 A0
port 12 n
rlabel metal1 797 501 831 535 1 A0
port 13 n
rlabel metal1 797 427 831 461 1 A0
port 14 n
rlabel metal1 1463 723 1497 757 1 A1
port 15 n
rlabel metal1 1463 649 1497 683 1 A1
port 16 n
rlabel metal1 1463 501 1497 535 1 A1
port 17 n
rlabel metal1 1463 427 1497 461 1 A1
port 18 n
rlabel metal1 1463 871 1497 905 1 A1
port 19 n
rlabel metal1 1463 797 1497 831 1 A1
port 20 n
rlabel metal1 131 575 165 609 1 S
port 21 n
rlabel metal1 131 649 165 683 1 S
port 22 n
rlabel metal1 131 723 165 757 1 S
port 23 n
rlabel metal1 131 797 165 831 1 S
port 24 n
rlabel metal1 131 871 165 905 1 S
port 25 n
rlabel metal1 131 501 165 535 1 S
port 26 n
rlabel metal1 131 427 165 461 1 S
port 27 n
rlabel metal1 649 871 683 905 1 S
port 28 n
rlabel metal1 649 797 683 831 1 S
port 29 n
rlabel metal1 649 723 683 757 1 S
port 30 n
rlabel metal1 649 575 683 609 1 S
port 31 n
rlabel metal1 649 501 683 535 1 S
port 32 n
rlabel metal1 649 427 683 461 1 S
port 33 n
rlabel metal1 -34 1446 2476 1514 1 VPWR
port 34 n
rlabel metal1 -34 -34 2476 34 1 VGND
port 35 n
rlabel nwell 57 1463 91 1497 1 VPB
port 36 n
rlabel pwell 57 -17 91 17 1 VNB
port 37 n
<< end >>
