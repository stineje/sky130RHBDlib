magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 98 157 367 203
rect 1 21 367 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 174 47 204 177
rect 258 47 288 177
<< scpmoshvt >>
rect 79 361 109 489
rect 174 297 204 497
rect 258 297 288 497
<< ndiff >>
rect 124 131 174 177
rect 27 106 79 131
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 93 174 131
rect 109 59 128 93
rect 162 59 174 93
rect 109 47 174 59
rect 204 123 258 177
rect 204 89 214 123
rect 248 89 258 123
rect 204 47 258 89
rect 288 165 341 177
rect 288 131 298 165
rect 332 131 341 165
rect 288 97 341 131
rect 288 63 298 97
rect 332 63 341 97
rect 288 47 341 63
<< pdiff >>
rect 124 489 174 497
rect 27 477 79 489
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 361 79 375
rect 109 477 174 489
rect 109 443 128 477
rect 162 443 174 477
rect 109 409 174 443
rect 109 375 128 409
rect 162 375 174 409
rect 109 361 174 375
rect 124 297 174 361
rect 204 461 258 497
rect 204 427 214 461
rect 248 427 258 461
rect 204 380 258 427
rect 204 346 214 380
rect 248 346 258 380
rect 204 297 258 346
rect 288 485 341 497
rect 288 451 298 485
rect 332 451 341 485
rect 288 417 341 451
rect 288 383 298 417
rect 332 383 341 417
rect 288 349 341 383
rect 288 315 298 349
rect 332 315 341 349
rect 288 297 341 315
<< ndiffc >>
rect 35 72 69 106
rect 128 59 162 93
rect 214 89 248 123
rect 298 131 332 165
rect 298 63 332 97
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 128 443 162 477
rect 128 375 162 409
rect 214 427 248 461
rect 214 346 248 380
rect 298 451 332 485
rect 298 383 332 417
rect 298 315 332 349
<< poly >>
rect 79 489 109 515
rect 174 497 204 523
rect 258 497 288 523
rect 79 265 109 361
rect 174 265 204 297
rect 258 265 288 297
rect 27 249 109 265
rect 27 215 37 249
rect 71 215 109 249
rect 27 199 109 215
rect 151 249 288 265
rect 151 215 161 249
rect 195 215 288 249
rect 151 199 288 215
rect 79 131 109 199
rect 174 177 204 199
rect 258 177 288 199
rect 79 21 109 47
rect 174 21 204 47
rect 258 21 288 47
<< polycont >>
rect 37 215 71 249
rect 161 215 195 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 35 477 69 493
rect 35 409 69 443
rect 112 477 178 527
rect 112 443 128 477
rect 162 443 178 477
rect 112 409 178 443
rect 112 375 128 409
rect 162 375 178 409
rect 212 461 263 493
rect 212 427 214 461
rect 248 427 263 461
rect 212 380 263 427
rect 35 341 69 375
rect 212 346 214 380
rect 248 346 263 380
rect 35 307 178 341
rect 212 312 263 346
rect 17 249 88 271
rect 17 215 37 249
rect 71 215 88 249
rect 17 197 88 215
rect 144 265 178 307
rect 144 249 195 265
rect 144 215 161 249
rect 144 199 195 215
rect 144 161 178 199
rect 229 166 263 312
rect 298 485 350 527
rect 332 451 350 485
rect 298 417 350 451
rect 332 383 350 417
rect 298 349 350 383
rect 332 315 350 349
rect 298 297 350 315
rect 35 127 178 161
rect 35 106 69 127
rect 212 123 263 166
rect 35 51 69 72
rect 112 59 128 93
rect 162 59 178 93
rect 112 17 178 59
rect 212 89 214 123
rect 248 89 263 123
rect 212 51 263 89
rect 298 165 350 185
rect 332 131 350 165
rect 298 97 350 131
rect 332 63 350 97
rect 298 17 350 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel locali s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel locali s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel locali s 212 85 246 119 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 212 357 246 391 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 212 425 246 459 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 buf_2
rlabel metal1 s 0 -48 368 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 368 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 368 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 3092062
string GDS_START 3087626
string path 0.000 13.600 9.200 13.600 
<< end >>
