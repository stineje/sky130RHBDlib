** sch_path: /home/rjridle/OpenRadHardSCL/sky130A/libs.tech/xschem/sky130_stdcells/fa_1.sym
.subckt fa_1

.ends
.end
