* SPICE3 file created from NAND2X1.ext - technology: sky130A

.subckt NAND2X1 Y A B VPB VNB
M1000 VNB a_168_157# a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1001 VPB.t1 a_168_157# a_217_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPB.t3 a_343_383# a_217_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_217_1004.t0 a_168_157# VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_217_1004.t3 a_343_383# VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VPB a_168_157# 0.08fF
C1 a_343_383# VPB 0.07fF
C2 a_343_383# a_168_157# 0.26fF
R0 a_217_1004.n5 a_217_1004.n3 356.633
R1 a_217_1004.n3 a_217_1004.n2 76.002
R2 a_217_1004.n5 a_217_1004.n4 30
R3 a_217_1004.n6 a_217_1004.n0 24.383
R4 a_217_1004.n6 a_217_1004.n5 23.684
R5 a_217_1004.n1 a_217_1004.t2 14.282
R6 a_217_1004.n1 a_217_1004.t3 14.282
R7 a_217_1004.n2 a_217_1004.t1 14.282
R8 a_217_1004.n2 a_217_1004.t0 14.282
R9 a_217_1004.n3 a_217_1004.n1 12.85
R10 VPB VPB.n78 126.832
R11 VPB.n71 VPB.n70 76
R12 VPB.n42 VPB.t0 55.106
R13 VPB.n60 VPB.t3 55.106
R14 VPB.n57 VPB.n56 48.952
R15 VPB.n44 VPB.n43 44.502
R16 VPB.n51 VPB.n41 40.824
R17 VPB.n65 VPB.n64 35.118
R18 VPB.n75 VPB.n71 20.452
R19 VPB.n40 VPB.n37 20.452
R20 VPB.n53 VPB.n52 17.801
R21 VPB.n41 VPB.t2 14.282
R22 VPB.n41 VPB.t1 14.282
R23 VPB.n40 VPB.n39 13.653
R24 VPB.n39 VPB.n38 13.653
R25 VPB.n63 VPB.n62 13.653
R26 VPB.n62 VPB.n61 13.653
R27 VPB.n59 VPB.n58 13.653
R28 VPB.n58 VPB.n57 13.653
R29 VPB.n55 VPB.n54 13.653
R30 VPB.n54 VPB.n53 13.653
R31 VPB.n50 VPB.n49 13.653
R32 VPB.n49 VPB.n48 13.653
R33 VPB.n46 VPB.n45 13.653
R34 VPB.n45 VPB.n44 13.653
R35 VPB.n16 VPB.n15 13.653
R36 VPB.n15 VPB.n14 13.653
R37 VPB.n71 VPB.n0 13.653
R38 VPB VPB.n0 13.653
R39 VPB.n48 VPB.n47 13.35
R40 VPB.n75 VPB.n74 13.276
R41 VPB.n74 VPB.n72 13.276
R42 VPB.n59 VPB.n55 13.276
R43 VPB.n50 VPB.n46 13.276
R44 VPB.n71 VPB.n16 13.276
R45 VPB.n37 VPB.n19 13.276
R46 VPB.n19 VPB.n17 13.276
R47 VPB.n24 VPB.n22 12.796
R48 VPB.n24 VPB.n23 12.564
R49 VPB.n30 VPB.n29 12.198
R50 VPB.n32 VPB.n31 12.198
R51 VPB.n30 VPB.n27 12.198
R52 VPB.n60 VPB.n59 11.841
R53 VPB.n46 VPB.n42 11.482
R54 VPB.n37 VPB.n36 7.5
R55 VPB.n22 VPB.n21 7.5
R56 VPB.n29 VPB.n28 7.5
R57 VPB.n27 VPB.n26 7.5
R58 VPB.n19 VPB.n18 7.5
R59 VPB.n34 VPB.n20 7.5
R60 VPB.n74 VPB.n73 7.5
R61 VPB.n12 VPB.n11 7.5
R62 VPB.n6 VPB.n5 7.5
R63 VPB.n8 VPB.n7 7.5
R64 VPB.n2 VPB.n1 7.5
R65 VPB.n76 VPB.n75 7.5
R66 VPB.n51 VPB.n50 6.817
R67 VPB.n13 VPB.n10 6.729
R68 VPB.n9 VPB.n6 6.729
R69 VPB.n4 VPB.n2 6.729
R70 VPB.n4 VPB.n3 6.728
R71 VPB.n9 VPB.n8 6.728
R72 VPB.n13 VPB.n12 6.728
R73 VPB.n77 VPB.n76 6.728
R74 VPB.n55 VPB.n51 6.458
R75 VPB.n36 VPB.n35 6.398
R76 VPB.n64 VPB.n40 6.112
R77 VPB.n64 VPB.n63 6.101
R78 VPB.n42 VPB.n16 1.794
R79 VPB.n63 VPB.n60 1.435
R80 VPB.n34 VPB.n25 1.402
R81 VPB.n34 VPB.n30 1.402
R82 VPB.n34 VPB.n32 1.402
R83 VPB.n34 VPB.n33 1.402
R84 VPB.n35 VPB.n34 0.735
R85 VPB.n34 VPB.n24 0.735
R86 VPB.n78 VPB.n13 0.387
R87 VPB.n78 VPB.n9 0.387
R88 VPB.n78 VPB.n4 0.387
R89 VPB.n78 VPB.n77 0.387
R90 VPB.n70 VPB 0.198
R91 VPB.n66 VPB.n65 0.136
R92 VPB.n68 VPB.n67 0.136
R93 VPB.n69 VPB.n68 0.136
R94 VPB.n70 VPB.n69 0.136
R95 VPB VPB.n66 0.068
R96 VPB.n67 VPB 0.068
R97 a_112_73.n10 a_112_73.n9 93.333
R98 a_112_73.n2 a_112_73.n1 41.622
R99 a_112_73.n13 a_112_73.n12 26.667
R100 a_112_73.n6 a_112_73.n5 24.977
R101 a_112_73.t0 a_112_73.n2 21.209
R102 a_112_73.t0 a_112_73.n3 11.595
R103 a_112_73.t1 a_112_73.n8 8.137
R104 a_112_73.t0 a_112_73.n0 6.109
R105 a_112_73.t1 a_112_73.n7 4.864
R106 a_112_73.t0 a_112_73.n4 3.871
R107 a_112_73.t0 a_112_73.n13 2.535
R108 a_112_73.n13 a_112_73.t1 1.145
R109 a_112_73.n7 a_112_73.n6 1.13
R110 a_112_73.t1 a_112_73.n11 0.804
R111 a_112_73.n11 a_112_73.n10 0.136
R112 VNB VNB.n62 300.778
R113 VNB.n29 VNB.n25 84.842
R114 VNB.n49 VNB.n48 76
R115 VNB.n27 VNB.n26 36.678
R116 VNB.n43 VNB.n42 35.118
R117 VNB.n24 VNB.n21 20.452
R118 VNB.n50 VNB.n49 20.452
R119 VNB.n41 VNB.n40 13.653
R120 VNB.n40 VNB.n39 13.653
R121 VNB.n38 VNB.n37 13.653
R122 VNB.n37 VNB.n36 13.653
R123 VNB.n35 VNB.n34 13.653
R124 VNB.n34 VNB.n33 13.653
R125 VNB.n32 VNB.n31 13.653
R126 VNB.n31 VNB.n30 13.653
R127 VNB.n28 VNB.n27 13.653
R128 VNB.n6 VNB.n5 13.653
R129 VNB.n5 VNB.n4 13.653
R130 VNB.n49 VNB.n0 13.653
R131 VNB VNB.n0 13.653
R132 VNB.n24 VNB.n23 13.653
R133 VNB.n23 VNB.n22 13.653
R134 VNB.n57 VNB.n54 13.577
R135 VNB.n9 VNB.n7 13.276
R136 VNB.n21 VNB.n9 13.276
R137 VNB.n41 VNB.n38 13.276
R138 VNB.n38 VNB.n35 13.276
R139 VNB.n35 VNB.n32 13.276
R140 VNB.n28 VNB.n6 13.276
R141 VNB.n49 VNB.n6 13.276
R142 VNB.n3 VNB.n1 13.276
R143 VNB.n50 VNB.n3 13.276
R144 VNB.n32 VNB.n29 10.764
R145 VNB.n59 VNB.n58 7.5
R146 VNB.n51 VNB.n50 7.5
R147 VNB.n3 VNB.n2 7.5
R148 VNB.n56 VNB.n55 7.5
R149 VNB.n15 VNB.n14 7.5
R150 VNB.n11 VNB.n10 7.5
R151 VNB.n9 VNB.n8 7.5
R152 VNB.n21 VNB.n20 7.5
R153 VNB.n61 VNB.n59 7.011
R154 VNB.n17 VNB.n15 7.011
R155 VNB.n13 VNB.n11 7.011
R156 VNB.n20 VNB.n19 7.01
R157 VNB.n13 VNB.n12 7.01
R158 VNB.n17 VNB.n16 7.01
R159 VNB.n61 VNB.n60 7.01
R160 VNB.n57 VNB.n56 6.788
R161 VNB.n52 VNB.n51 6.788
R162 VNB.n42 VNB.n24 6.111
R163 VNB.n42 VNB.n41 6.1
R164 VNB.n29 VNB.n28 2.511
R165 VNB.n62 VNB.n53 0.921
R166 VNB.n62 VNB.n57 0.476
R167 VNB.n62 VNB.n52 0.475
R168 VNB.n18 VNB.n13 0.246
R169 VNB.n19 VNB.n18 0.246
R170 VNB.n18 VNB.n17 0.246
R171 VNB.n62 VNB.n61 0.246
R172 VNB.n48 VNB 0.198
R173 VNB.n44 VNB.n43 0.136
R174 VNB.n46 VNB.n45 0.136
R175 VNB.n47 VNB.n46 0.136
R176 VNB.n48 VNB.n47 0.136
R177 VNB VNB.n44 0.068
R178 VNB.n45 VNB 0.068
C3 VPB VNB 3.66fF
C4 a_112_73.n0 VNB 0.02fF
C5 a_112_73.n1 VNB 0.09fF
C6 a_112_73.n2 VNB 0.07fF
C7 a_112_73.n3 VNB 0.05fF
C8 a_112_73.n4 VNB 0.00fF
C9 a_112_73.n5 VNB 0.04fF
C10 a_112_73.n6 VNB 0.05fF
C11 a_112_73.n7 VNB 0.02fF
C12 a_112_73.n8 VNB 0.05fF
C13 a_112_73.n9 VNB 0.02fF
C14 a_112_73.n10 VNB 0.07fF
C15 a_112_73.n11 VNB 0.16fF
C16 a_112_73.t1 VNB 0.22fF
C17 a_112_73.n12 VNB 0.08fF
C18 a_112_73.n13 VNB 0.00fF
C19 VPB.n0 VNB 0.03fF
C20 VPB.n1 VNB 0.03fF
C21 VPB.n2 VNB 0.02fF
C22 VPB.n3 VNB 0.13fF
C23 VPB.n5 VNB 0.02fF
C24 VPB.n6 VNB 0.02fF
C25 VPB.n7 VNB 0.02fF
C26 VPB.n8 VNB 0.02fF
C27 VPB.n10 VNB 0.02fF
C28 VPB.n11 VNB 0.02fF
C29 VPB.n12 VNB 0.02fF
C30 VPB.n14 VNB 0.22fF
C31 VPB.n15 VNB 0.02fF
C32 VPB.n16 VNB 0.01fF
C33 VPB.n17 VNB 0.02fF
C34 VPB.n18 VNB 0.02fF
C35 VPB.n19 VNB 0.02fF
C36 VPB.n20 VNB 0.13fF
C37 VPB.n21 VNB 0.02fF
C38 VPB.n22 VNB 0.02fF
C39 VPB.n23 VNB 0.04fF
C40 VPB.n24 VNB 0.01fF
C41 VPB.n26 VNB 0.02fF
C42 VPB.n27 VNB 0.02fF
C43 VPB.n28 VNB 0.02fF
C44 VPB.n29 VNB 0.02fF
C45 VPB.n31 VNB 0.02fF
C46 VPB.n34 VNB 0.42fF
C47 VPB.n36 VNB 0.03fF
C48 VPB.n37 VNB 0.04fF
C49 VPB.n38 VNB 0.25fF
C50 VPB.n39 VNB 0.03fF
C51 VPB.n40 VNB 0.03fF
C52 VPB.n41 VNB 0.09fF
C53 VPB.n42 VNB 0.05fF
C54 VPB.n43 VNB 0.13fF
C55 VPB.n44 VNB 0.15fF
C56 VPB.n45 VNB 0.02fF
C57 VPB.n46 VNB 0.02fF
C58 VPB.n47 VNB 0.13fF
C59 VPB.n48 VNB 0.14fF
C60 VPB.n49 VNB 0.02fF
C61 VPB.n50 VNB 0.02fF
C62 VPB.n51 VNB 0.02fF
C63 VPB.n52 VNB 0.13fF
C64 VPB.n53 VNB 0.14fF
C65 VPB.n54 VNB 0.02fF
C66 VPB.n55 VNB 0.02fF
C67 VPB.n56 VNB 0.13fF
C68 VPB.n57 VNB 0.15fF
C69 VPB.n58 VNB 0.02fF
C70 VPB.n59 VNB 0.02fF
C71 VPB.n60 VNB 0.05fF
C72 VPB.n61 VNB 0.21fF
C73 VPB.n62 VNB 0.02fF
C74 VPB.n63 VNB 0.01fF
C75 VPB.n64 VNB 0.00fF
C76 VPB.n65 VNB 0.09fF
C77 VPB.n66 VNB 0.02fF
C78 VPB.n67 VNB 0.02fF
C79 VPB.n68 VNB 0.02fF
C80 VPB.n69 VNB 0.02fF
C81 VPB.n70 VNB 0.03fF
C82 VPB.n71 VNB 0.03fF
C83 VPB.n72 VNB 0.02fF
C84 VPB.n73 VNB 0.02fF
C85 VPB.n74 VNB 0.02fF
C86 VPB.n75 VNB 0.04fF
C87 VPB.n76 VNB 0.03fF
C88 VPB.n78 VNB 0.39fF
C89 a_217_1004.n0 VNB 0.04fF
C90 a_217_1004.n1 VNB 0.47fF
C91 a_217_1004.n2 VNB 0.55fF
C92 a_217_1004.n3 VNB 0.48fF
C93 a_217_1004.n4 VNB 0.03fF
C94 a_217_1004.n5 VNB 0.41fF
C95 a_217_1004.n6 VNB 0.05fF
.ends
