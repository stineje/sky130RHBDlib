* SPICE3 file created from AO3X1.ext - technology: sky130A

.subckt AO3X1 Y A B C VDD VSS
X0 VDD A a_223_1051 VDD sky130_fd_pr__pfet_01v8 ad=2.78p pd=2.278u as=0p ps=0u w=2u l=0.15u M=2
X1 a_223_1051 a_653_990 C VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.8p ps=4.58u w=2u l=0.15u M=2
X2 C B a_108_101 VSS sky130_fd_pr__nfet_01v8 ad=1.3277p pd=9.77u as=0p ps=0u w=3u l=0.15u
X3 Y C VDD VDD sky130_fd_pr__pfet_01v8 ad=5.8p pd=4.58u as=0p ps=0u w=2u l=0.15u M=2
X4 a_223_1051 B VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2u l=0.15u M=2
X5 Y C VSS VSS sky130_fd_pr__nfet_01v8 ad=1.791p pd=1.57u as=1.499p ps=1.124u w=3u l=0.15u
X6 VSS A a_108_101 VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
X7 VSS a_653_990 C VSS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=3u l=0.15u
C0 a_223_1051 VDD 2.28fF
C1 VDD VSS 2.67fF
.ends
