// File: TMRDFFSNRNQNX1.spi.TMRDFFSNRNQNX1.pxi
// Created: Tue Oct 15 15:53:00 2024
// 
simulator lang=spectre
x_PM_TMRDFFSNRNQNX1\%GND ( GND N_GND_c_89_p N_GND_c_208_p N_GND_c_1_p \
 N_GND_c_215_p N_GND_c_31_p N_GND_c_38_p N_GND_c_41_p N_GND_c_48_p \
 N_GND_c_57_p N_GND_c_64_p N_GND_c_73_p N_GND_c_80_p N_GND_c_94_p \
 N_GND_c_101_p N_GND_c_218_p N_GND_c_225_p N_GND_c_141_p N_GND_c_148_p \
 N_GND_c_151_p N_GND_c_158_p N_GND_c_167_p N_GND_c_174_p N_GND_c_181_p \
 N_GND_c_188_p N_GND_c_347_p N_GND_c_348_p N_GND_c_228_p N_GND_c_235_p \
 N_GND_c_246_p N_GND_c_253_p N_GND_c_256_p N_GND_c_263_p N_GND_c_272_p \
 N_GND_c_279_p N_GND_c_292_p N_GND_c_299_p N_GND_c_416_p N_GND_c_422_p \
 N_GND_c_104_p N_GND_c_111_p N_GND_c_114_p N_GND_c_120_p N_GND_c_448_p \
 N_GND_c_2_p N_GND_c_3_p N_GND_c_4_p N_GND_c_5_p N_GND_c_6_p N_GND_c_7_p \
 N_GND_c_8_p N_GND_c_9_p N_GND_c_10_p N_GND_c_11_p N_GND_c_12_p N_GND_c_13_p \
 N_GND_c_14_p N_GND_c_15_p N_GND_c_16_p N_GND_c_17_p N_GND_c_18_p N_GND_c_19_p \
 N_GND_c_20_p N_GND_c_21_p N_GND_c_22_p N_GND_M0_noxref_d N_GND_M3_noxref_d \
 N_GND_M6_noxref_d N_GND_M9_noxref_d N_GND_M12_noxref_d N_GND_M15_noxref_d \
 N_GND_M18_noxref_d N_GND_M21_noxref_d N_GND_M24_noxref_d N_GND_M27_noxref_d \
 N_GND_M30_noxref_d N_GND_M33_noxref_d N_GND_M36_noxref_d N_GND_M39_noxref_d \
 N_GND_M42_noxref_d N_GND_M45_noxref_d N_GND_M48_noxref_d N_GND_M51_noxref_d \
 N_GND_M54_noxref_d N_GND_M56_noxref_d N_GND_M58_noxref_d )  \
 PM_TMRDFFSNRNQNX1\%GND
x_PM_TMRDFFSNRNQNX1\%VDD ( VDD N_VDD_c_1085_p N_VDD_c_1658_p N_VDD_c_1063_n \
 N_VDD_c_1086_p N_VDD_c_1087_p N_VDD_c_1093_p N_VDD_c_1097_p N_VDD_c_1648_p \
 N_VDD_c_1106_p N_VDD_c_1175_p N_VDD_c_1181_p N_VDD_c_1185_p N_VDD_c_1784_p \
 N_VDD_c_1110_p N_VDD_c_1135_p N_VDD_c_1141_p N_VDD_c_1145_p N_VDD_c_1787_p \
 N_VDD_c_1151_p N_VDD_c_1358_p N_VDD_c_1364_p N_VDD_c_1368_p N_VDD_c_1796_p \
 N_VDD_c_1195_p N_VDD_c_1300_p N_VDD_c_1306_p N_VDD_c_1217_p N_VDD_c_1218_p \
 N_VDD_c_1219_p N_VDD_c_1402_p N_VDD_c_1380_p N_VDD_c_1220_p N_VDD_c_1221_p \
 N_VDD_c_1222_p N_VDD_c_1436_p N_VDD_c_1442_p N_VDD_c_1223_p N_VDD_c_1224_p \
 N_VDD_c_1225_p N_VDD_c_1524_p N_VDD_c_1530_p N_VDD_c_1226_p N_VDD_c_1227_p \
 N_VDD_c_1228_p N_VDD_c_1484_p N_VDD_c_1490_p N_VDD_c_1229_p N_VDD_c_1230_p \
 N_VDD_c_1231_p N_VDD_c_1569_p N_VDD_c_1575_p N_VDD_c_1232_p N_VDD_c_1233_p \
 N_VDD_c_1234_p N_VDD_c_1920_p N_VDD_c_1626_p N_VDD_c_1235_p N_VDD_c_1236_p \
 N_VDD_c_1237_p N_VDD_c_1613_p N_VDD_c_1591_p N_VDD_c_1238_p N_VDD_c_1239_p \
 N_VDD_c_1240_p N_VDD_c_1697_p N_VDD_c_1703_p N_VDD_c_1241_p N_VDD_c_1242_p \
 N_VDD_c_1243_p N_VDD_c_1836_p N_VDD_c_1853_p N_VDD_c_1244_p N_VDD_c_1245_p \
 N_VDD_c_1246_p N_VDD_c_1745_p N_VDD_c_1751_p N_VDD_c_1247_p N_VDD_c_1248_p \
 N_VDD_c_1249_p N_VDD_c_1840_p N_VDD_c_1928_p N_VDD_c_1276_p N_VDD_c_1277_p \
 N_VDD_c_1278_p N_VDD_c_1932_p N_VDD_c_2030_p N_VDD_c_1279_p N_VDD_c_1280_p \
 N_VDD_c_1281_p N_VDD_c_1964_p N_VDD_c_1994_p N_VDD_c_1282_p N_VDD_c_1283_p \
 N_VDD_c_1290_p N_VDD_c_2050_p N_VDD_c_2051_p N_VDD_c_1331_p N_VDD_c_1064_n \
 N_VDD_c_1065_n N_VDD_c_1066_n N_VDD_c_1067_n N_VDD_c_1068_n N_VDD_c_1069_n \
 N_VDD_c_1070_n N_VDD_c_1071_n N_VDD_c_1072_n N_VDD_c_1073_n N_VDD_c_1074_n \
 N_VDD_c_1075_n N_VDD_c_1076_n N_VDD_c_1077_n N_VDD_c_1078_n N_VDD_c_1079_n \
 N_VDD_c_1080_n N_VDD_c_1081_n N_VDD_c_1082_n N_VDD_c_1083_n N_VDD_c_1084_n \
 N_VDD_M60_noxref_s N_VDD_M61_noxref_d N_VDD_M63_noxref_d N_VDD_M65_noxref_d \
 N_VDD_M66_noxref_s N_VDD_M67_noxref_d N_VDD_M69_noxref_d N_VDD_M71_noxref_d \
 N_VDD_M72_noxref_s N_VDD_M73_noxref_d N_VDD_M75_noxref_d N_VDD_M77_noxref_d \
 N_VDD_M78_noxref_s N_VDD_M79_noxref_d N_VDD_M81_noxref_d N_VDD_M83_noxref_d \
 N_VDD_M84_noxref_s N_VDD_M85_noxref_d N_VDD_M87_noxref_d N_VDD_M89_noxref_d \
 N_VDD_M90_noxref_s N_VDD_M91_noxref_d N_VDD_M93_noxref_d N_VDD_M95_noxref_d \
 N_VDD_M96_noxref_s N_VDD_M97_noxref_d N_VDD_M99_noxref_d N_VDD_M101_noxref_d \
 N_VDD_M102_noxref_s N_VDD_M103_noxref_d N_VDD_M105_noxref_d \
 N_VDD_M107_noxref_d N_VDD_M108_noxref_s N_VDD_M109_noxref_d \
 N_VDD_M111_noxref_d N_VDD_M113_noxref_d N_VDD_M114_noxref_s \
 N_VDD_M115_noxref_d N_VDD_M117_noxref_d N_VDD_M119_noxref_d \
 N_VDD_M120_noxref_s N_VDD_M121_noxref_d N_VDD_M123_noxref_d \
 N_VDD_M125_noxref_d N_VDD_M126_noxref_s N_VDD_M127_noxref_d \
 N_VDD_M129_noxref_d N_VDD_M131_noxref_d N_VDD_M132_noxref_s \
 N_VDD_M133_noxref_d N_VDD_M135_noxref_d N_VDD_M137_noxref_d \
 N_VDD_M138_noxref_s N_VDD_M139_noxref_d N_VDD_M141_noxref_d \
 N_VDD_M143_noxref_d N_VDD_M144_noxref_s N_VDD_M145_noxref_d \
 N_VDD_M147_noxref_d N_VDD_M149_noxref_d N_VDD_M150_noxref_s \
 N_VDD_M151_noxref_d N_VDD_M153_noxref_d N_VDD_M155_noxref_d \
 N_VDD_M156_noxref_s N_VDD_M157_noxref_d N_VDD_M159_noxref_d \
 N_VDD_M161_noxref_d N_VDD_M162_noxref_s N_VDD_M163_noxref_d \
 N_VDD_M165_noxref_d N_VDD_M167_noxref_d N_VDD_M168_noxref_s \
 N_VDD_M169_noxref_d N_VDD_M171_noxref_d )  PM_TMRDFFSNRNQNX1\%VDD
x_PM_TMRDFFSNRNQNX1\%noxref_3 ( N_noxref_3_c_2221_n N_noxref_3_c_2222_n \
 N_noxref_3_c_2223_n N_noxref_3_c_2224_n N_noxref_3_c_2250_n \
 N_noxref_3_c_2254_n N_noxref_3_c_2256_n N_noxref_3_c_2260_n \
 N_noxref_3_c_2225_n N_noxref_3_c_2396_p N_noxref_3_c_2226_n \
 N_noxref_3_c_2227_n N_noxref_3_c_2228_n N_noxref_3_c_2408_p \
 N_noxref_3_c_2317_p N_noxref_3_M3_noxref_g N_noxref_3_M6_noxref_g \
 N_noxref_3_M66_noxref_g N_noxref_3_M67_noxref_g N_noxref_3_M72_noxref_g \
 N_noxref_3_M73_noxref_g N_noxref_3_c_2229_n N_noxref_3_c_2231_n \
 N_noxref_3_c_2232_n N_noxref_3_c_2233_n N_noxref_3_c_2234_n \
 N_noxref_3_c_2235_n N_noxref_3_c_2236_n N_noxref_3_c_2238_n \
 N_noxref_3_c_2321_p N_noxref_3_c_2279_n N_noxref_3_c_2239_n \
 N_noxref_3_c_2241_n N_noxref_3_c_2242_n N_noxref_3_c_2243_n \
 N_noxref_3_c_2244_n N_noxref_3_c_2245_n N_noxref_3_c_2246_n \
 N_noxref_3_c_2248_n N_noxref_3_c_2301_p N_noxref_3_c_2281_n \
 N_noxref_3_M2_noxref_d N_noxref_3_M60_noxref_d N_noxref_3_M62_noxref_d \
 N_noxref_3_M64_noxref_d )  PM_TMRDFFSNRNQNX1\%noxref_3
x_PM_TMRDFFSNRNQNX1\%noxref_4 ( N_noxref_4_c_2461_n N_noxref_4_c_2462_n \
 N_noxref_4_c_2477_n N_noxref_4_c_2481_n N_noxref_4_c_2483_n \
 N_noxref_4_c_2487_n N_noxref_4_c_2463_n N_noxref_4_c_2590_p \
 N_noxref_4_c_2464_n N_noxref_4_c_2465_n N_noxref_4_c_2605_p \
 N_noxref_4_c_2532_p N_noxref_4_M9_noxref_g N_noxref_4_M78_noxref_g \
 N_noxref_4_M79_noxref_g N_noxref_4_c_2466_n N_noxref_4_c_2468_n \
 N_noxref_4_c_2469_n N_noxref_4_c_2470_n N_noxref_4_c_2471_n \
 N_noxref_4_c_2472_n N_noxref_4_c_2473_n N_noxref_4_c_2475_n \
 N_noxref_4_c_2536_p N_noxref_4_c_2499_n N_noxref_4_M8_noxref_d \
 N_noxref_4_M72_noxref_d N_noxref_4_M74_noxref_d N_noxref_4_M76_noxref_d )  \
 PM_TMRDFFSNRNQNX1\%noxref_4
x_PM_TMRDFFSNRNQNX1\%noxref_5 ( N_noxref_5_c_2626_n N_noxref_5_c_2692_n \
 N_noxref_5_c_2627_n N_noxref_5_c_2695_n N_noxref_5_c_2628_n \
 N_noxref_5_c_2643_n N_noxref_5_c_2647_n N_noxref_5_c_2649_n \
 N_noxref_5_c_2653_n N_noxref_5_c_2629_n N_noxref_5_c_2809_p \
 N_noxref_5_c_2657_n N_noxref_5_c_2630_n N_noxref_5_c_2789_p \
 N_noxref_5_c_2751_p N_noxref_5_M2_noxref_g N_noxref_5_M12_noxref_g \
 N_noxref_5_M64_noxref_g N_noxref_5_M65_noxref_g N_noxref_5_M84_noxref_g \
 N_noxref_5_M85_noxref_g N_noxref_5_c_2711_n N_noxref_5_c_2712_n \
 N_noxref_5_c_2713_n N_noxref_5_c_2714_n N_noxref_5_c_2715_n \
 N_noxref_5_c_2717_n N_noxref_5_c_2718_n N_noxref_5_c_2631_n \
 N_noxref_5_c_2633_n N_noxref_5_c_2634_n N_noxref_5_c_2635_n \
 N_noxref_5_c_2636_n N_noxref_5_c_2637_n N_noxref_5_c_2638_n \
 N_noxref_5_c_2640_n N_noxref_5_c_2734_p N_noxref_5_c_2669_n \
 N_noxref_5_c_2720_n N_noxref_5_c_2721_n N_noxref_5_c_2723_n \
 N_noxref_5_M5_noxref_d N_noxref_5_M66_noxref_d N_noxref_5_M68_noxref_d \
 N_noxref_5_M70_noxref_d )  PM_TMRDFFSNRNQNX1\%noxref_5
x_PM_TMRDFFSNRNQNX1\%noxref_6 ( N_noxref_6_c_2893_n N_noxref_6_c_2894_n \
 N_noxref_6_c_2934_n N_noxref_6_c_2990_n N_noxref_6_c_3219_p \
 N_noxref_6_c_2993_n N_noxref_6_c_3220_p N_noxref_6_c_3007_n \
 N_noxref_6_c_3012_n N_noxref_6_c_3016_n N_noxref_6_c_3020_n \
 N_noxref_6_c_3022_n N_noxref_6_c_3026_n N_noxref_6_c_2895_n \
 N_noxref_6_c_3255_p N_noxref_6_c_2896_n N_noxref_6_c_2897_n \
 N_noxref_6_c_2898_n N_noxref_6_c_2901_n N_noxref_6_c_3282_p \
 N_noxref_6_c_3093_p N_noxref_6_M15_noxref_g N_noxref_6_M54_noxref_g \
 N_noxref_6_M56_noxref_g N_noxref_6_M90_noxref_g N_noxref_6_M91_noxref_g \
 N_noxref_6_M168_noxref_g N_noxref_6_M169_noxref_g N_noxref_6_M172_noxref_g \
 N_noxref_6_M173_noxref_g N_noxref_6_c_2903_n N_noxref_6_c_2905_n \
 N_noxref_6_c_2906_n N_noxref_6_c_2907_n N_noxref_6_c_2908_n \
 N_noxref_6_c_2909_n N_noxref_6_c_2910_n N_noxref_6_c_2912_n \
 N_noxref_6_c_3098_p N_noxref_6_c_3052_n N_noxref_6_c_2913_n \
 N_noxref_6_c_2915_n N_noxref_6_c_2916_n N_noxref_6_c_2917_n \
 N_noxref_6_c_2918_n N_noxref_6_c_2919_n N_noxref_6_c_3381_p \
 N_noxref_6_c_3054_n N_noxref_6_c_2920_n N_noxref_6_c_2922_n \
 N_noxref_6_c_2923_n N_noxref_6_c_2925_n N_noxref_6_c_3416_p \
 N_noxref_6_c_2926_n N_noxref_6_c_2927_n N_noxref_6_c_2928_n \
 N_noxref_6_c_2929_n N_noxref_6_c_2931_n N_noxref_6_c_2932_n \
 N_noxref_6_c_3056_n N_noxref_6_M14_noxref_d N_noxref_6_M84_noxref_d \
 N_noxref_6_M86_noxref_d N_noxref_6_M88_noxref_d )  PM_TMRDFFSNRNQNX1\%noxref_6
x_PM_TMRDFFSNRNQNX1\%noxref_7 ( N_noxref_7_c_3577_n N_noxref_7_c_3579_n \
 N_noxref_7_c_3584_n N_noxref_7_c_3586_n N_noxref_7_c_3623_n \
 N_noxref_7_c_3625_n N_noxref_7_c_3527_n N_noxref_7_c_3528_n \
 N_noxref_7_c_3534_n N_noxref_7_c_3538_n N_noxref_7_c_3540_n \
 N_noxref_7_c_3544_n N_noxref_7_c_3529_n N_noxref_7_c_3751_p \
 N_noxref_7_c_3548_n N_noxref_7_c_3530_n N_noxref_7_c_3714_p \
 N_noxref_7_c_3762_p N_noxref_7_M5_noxref_g N_noxref_7_M8_noxref_g \
 N_noxref_7_M17_noxref_g N_noxref_7_M70_noxref_g N_noxref_7_M71_noxref_g \
 N_noxref_7_M76_noxref_g N_noxref_7_M77_noxref_g N_noxref_7_M94_noxref_g \
 N_noxref_7_M95_noxref_g N_noxref_7_c_3638_n N_noxref_7_c_3639_n \
 N_noxref_7_c_3640_n N_noxref_7_c_3641_n N_noxref_7_c_3642_n \
 N_noxref_7_c_3644_n N_noxref_7_c_3645_n N_noxref_7_c_3599_n \
 N_noxref_7_c_3600_n N_noxref_7_c_3601_n N_noxref_7_c_3602_n \
 N_noxref_7_c_3603_n N_noxref_7_c_3605_n N_noxref_7_c_3606_n \
 N_noxref_7_c_3677_p N_noxref_7_c_3678_p N_noxref_7_c_3679_p \
 N_noxref_7_c_3680_p N_noxref_7_c_3668_p N_noxref_7_c_3682_p \
 N_noxref_7_c_3669_p N_noxref_7_c_3647_n N_noxref_7_c_3648_n \
 N_noxref_7_c_3650_n N_noxref_7_c_3608_n N_noxref_7_c_3609_n \
 N_noxref_7_c_3611_n N_noxref_7_c_3672_p N_noxref_7_c_3673_p \
 N_noxref_7_c_3660_n N_noxref_7_M11_noxref_d N_noxref_7_M78_noxref_d \
 N_noxref_7_M80_noxref_d N_noxref_7_M82_noxref_d )  PM_TMRDFFSNRNQNX1\%noxref_7
x_PM_TMRDFFSNRNQNX1\%noxref_8 ( N_noxref_8_c_3906_n N_noxref_8_c_3904_n \
 N_noxref_8_c_3866_n N_noxref_8_c_3870_n N_noxref_8_c_3874_n \
 N_noxref_8_c_3876_n N_noxref_8_c_3880_n N_noxref_8_c_3867_n \
 N_noxref_8_c_3986_p N_noxref_8_c_3884_n N_noxref_8_c_4022_p \
 N_noxref_8_c_3958_n N_noxref_8_M14_noxref_g N_noxref_8_M88_noxref_g \
 N_noxref_8_M89_noxref_g N_noxref_8_c_3927_n N_noxref_8_c_3928_n \
 N_noxref_8_c_3929_n N_noxref_8_c_3930_n N_noxref_8_c_3931_n \
 N_noxref_8_c_3933_n N_noxref_8_c_3934_n N_noxref_8_c_3936_n \
 N_noxref_8_c_3937_n N_noxref_8_c_3939_n N_noxref_8_M17_noxref_d \
 N_noxref_8_M90_noxref_d N_noxref_8_M92_noxref_d N_noxref_8_M94_noxref_d )  \
 PM_TMRDFFSNRNQNX1\%noxref_8
x_PM_TMRDFFSNRNQNX1\%noxref_9 ( N_noxref_9_c_4042_n N_noxref_9_c_4043_n \
 N_noxref_9_c_4044_n N_noxref_9_c_4045_n N_noxref_9_c_4071_n \
 N_noxref_9_c_4075_n N_noxref_9_c_4077_n N_noxref_9_c_4081_n \
 N_noxref_9_c_4046_n N_noxref_9_c_4223_p N_noxref_9_c_4047_n \
 N_noxref_9_c_4048_n N_noxref_9_c_4049_n N_noxref_9_c_4235_p \
 N_noxref_9_c_4151_p N_noxref_9_M21_noxref_g N_noxref_9_M24_noxref_g \
 N_noxref_9_M102_noxref_g N_noxref_9_M103_noxref_g N_noxref_9_M108_noxref_g \
 N_noxref_9_M109_noxref_g N_noxref_9_c_4050_n N_noxref_9_c_4052_n \
 N_noxref_9_c_4053_n N_noxref_9_c_4054_n N_noxref_9_c_4055_n \
 N_noxref_9_c_4056_n N_noxref_9_c_4057_n N_noxref_9_c_4059_n \
 N_noxref_9_c_4127_n N_noxref_9_c_4100_n N_noxref_9_c_4060_n \
 N_noxref_9_c_4062_n N_noxref_9_c_4063_n N_noxref_9_c_4064_n \
 N_noxref_9_c_4065_n N_noxref_9_c_4066_n N_noxref_9_c_4067_n \
 N_noxref_9_c_4069_n N_noxref_9_c_4129_n N_noxref_9_c_4102_n \
 N_noxref_9_M20_noxref_d N_noxref_9_M96_noxref_d N_noxref_9_M98_noxref_d \
 N_noxref_9_M100_noxref_d )  PM_TMRDFFSNRNQNX1\%noxref_9
x_PM_TMRDFFSNRNQNX1\%noxref_10 ( N_noxref_10_c_4295_n N_noxref_10_c_4296_n \
 N_noxref_10_c_4311_n N_noxref_10_c_4315_n N_noxref_10_c_4317_n \
 N_noxref_10_c_4321_n N_noxref_10_c_4297_n N_noxref_10_c_4428_p \
 N_noxref_10_c_4298_n N_noxref_10_c_4299_n N_noxref_10_c_4443_p \
 N_noxref_10_c_4373_p N_noxref_10_M27_noxref_g N_noxref_10_M114_noxref_g \
 N_noxref_10_M115_noxref_g N_noxref_10_c_4300_n N_noxref_10_c_4302_n \
 N_noxref_10_c_4303_n N_noxref_10_c_4304_n N_noxref_10_c_4305_n \
 N_noxref_10_c_4306_n N_noxref_10_c_4307_n N_noxref_10_c_4309_n \
 N_noxref_10_c_4355_n N_noxref_10_c_4333_n N_noxref_10_M26_noxref_d \
 N_noxref_10_M108_noxref_d N_noxref_10_M110_noxref_d N_noxref_10_M112_noxref_d \
 )  PM_TMRDFFSNRNQNX1\%noxref_10
x_PM_TMRDFFSNRNQNX1\%noxref_11 ( N_noxref_11_c_4534_n N_noxref_11_c_4533_n \
 N_noxref_11_c_4541_n N_noxref_11_c_4543_n N_noxref_11_c_4464_n \
 N_noxref_11_c_4479_n N_noxref_11_c_4483_n N_noxref_11_c_4485_n \
 N_noxref_11_c_4489_n N_noxref_11_c_4465_n N_noxref_11_c_4650_p \
 N_noxref_11_c_4493_n N_noxref_11_c_4466_n N_noxref_11_c_4644_p \
 N_noxref_11_c_4595_p N_noxref_11_M20_noxref_g N_noxref_11_M30_noxref_g \
 N_noxref_11_M100_noxref_g N_noxref_11_M101_noxref_g N_noxref_11_M120_noxref_g \
 N_noxref_11_M121_noxref_g N_noxref_11_c_4559_n N_noxref_11_c_4560_n \
 N_noxref_11_c_4561_n N_noxref_11_c_4562_n N_noxref_11_c_4563_n \
 N_noxref_11_c_4565_n N_noxref_11_c_4566_n N_noxref_11_c_4467_n \
 N_noxref_11_c_4469_n N_noxref_11_c_4470_n N_noxref_11_c_4471_n \
 N_noxref_11_c_4472_n N_noxref_11_c_4473_n N_noxref_11_c_4474_n \
 N_noxref_11_c_4476_n N_noxref_11_c_4530_n N_noxref_11_c_4505_n \
 N_noxref_11_c_4568_n N_noxref_11_c_4569_n N_noxref_11_c_4532_n \
 N_noxref_11_M23_noxref_d N_noxref_11_M102_noxref_d N_noxref_11_M104_noxref_d \
 N_noxref_11_M106_noxref_d )  PM_TMRDFFSNRNQNX1\%noxref_11
x_PM_TMRDFFSNRNQNX1\%noxref_12 ( N_noxref_12_c_4809_n N_noxref_12_c_4849_n \
 N_noxref_12_c_4814_n N_noxref_12_c_4816_n N_noxref_12_c_4853_n \
 N_noxref_12_c_4855_n N_noxref_12_c_4745_n N_noxref_12_c_4746_n \
 N_noxref_12_c_4752_n N_noxref_12_c_4756_n N_noxref_12_c_4758_n \
 N_noxref_12_c_4762_n N_noxref_12_c_4747_n N_noxref_12_c_4968_p \
 N_noxref_12_c_4766_n N_noxref_12_c_4748_n N_noxref_12_c_4957_p \
 N_noxref_12_c_4979_p N_noxref_12_M23_noxref_g N_noxref_12_M26_noxref_g \
 N_noxref_12_M35_noxref_g N_noxref_12_M106_noxref_g N_noxref_12_M107_noxref_g \
 N_noxref_12_M112_noxref_g N_noxref_12_M113_noxref_g N_noxref_12_M130_noxref_g \
 N_noxref_12_M131_noxref_g N_noxref_12_c_4868_n N_noxref_12_c_4869_n \
 N_noxref_12_c_4870_n N_noxref_12_c_4871_n N_noxref_12_c_4872_n \
 N_noxref_12_c_4874_n N_noxref_12_c_4875_n N_noxref_12_c_4829_n \
 N_noxref_12_c_4830_n N_noxref_12_c_4831_n N_noxref_12_c_4832_n \
 N_noxref_12_c_4833_n N_noxref_12_c_4835_n N_noxref_12_c_4836_n \
 N_noxref_12_c_4899_p N_noxref_12_c_4900_p N_noxref_12_c_4901_p \
 N_noxref_12_c_4902_p N_noxref_12_c_4890_p N_noxref_12_c_4904_p \
 N_noxref_12_c_4891_p N_noxref_12_c_4877_n N_noxref_12_c_4878_n \
 N_noxref_12_c_4806_n N_noxref_12_c_4838_n N_noxref_12_c_4839_n \
 N_noxref_12_c_4807_n N_noxref_12_c_4894_p N_noxref_12_c_4895_p \
 N_noxref_12_c_4808_n N_noxref_12_M29_noxref_d N_noxref_12_M114_noxref_d \
 N_noxref_12_M116_noxref_d N_noxref_12_M118_noxref_d )  \
 PM_TMRDFFSNRNQNX1\%noxref_12
x_PM_TMRDFFSNRNQNX1\%noxref_13 ( N_noxref_13_c_5099_n N_noxref_13_c_5149_n \
 N_noxref_13_c_5101_n N_noxref_13_c_5106_n N_noxref_13_c_5110_n \
 N_noxref_13_c_5112_n N_noxref_13_c_5116_n N_noxref_13_c_5102_n \
 N_noxref_13_c_5183_p N_noxref_13_c_5103_n N_noxref_13_c_5219_p \
 N_noxref_13_c_5161_n N_noxref_13_M32_noxref_g N_noxref_13_M124_noxref_g \
 N_noxref_13_M125_noxref_g N_noxref_13_c_5197_p N_noxref_13_c_5198_p \
 N_noxref_13_c_5199_p N_noxref_13_c_5252_p N_noxref_13_c_5185_p \
 N_noxref_13_c_5254_p N_noxref_13_c_5234_p N_noxref_13_c_5186_p \
 N_noxref_13_c_5202_p N_noxref_13_c_5145_n N_noxref_13_M35_noxref_d \
 N_noxref_13_M126_noxref_d N_noxref_13_M128_noxref_d N_noxref_13_M130_noxref_d \
 )  PM_TMRDFFSNRNQNX1\%noxref_13
x_PM_TMRDFFSNRNQNX1\%D ( N_D_c_5277_n N_D_c_5278_n N_D_c_5328_n N_D_c_5334_n D \
 D D D D D D D D D D D D D N_D_c_5279_n N_D_c_5280_n N_D_c_5281_n \
 N_D_M0_noxref_g N_D_M18_noxref_g N_D_M36_noxref_g N_D_M60_noxref_g \
 N_D_M61_noxref_g N_D_M96_noxref_g N_D_M97_noxref_g N_D_M132_noxref_g \
 N_D_M133_noxref_g N_D_c_5282_n N_D_c_5284_n N_D_c_5285_n N_D_c_5286_n \
 N_D_c_5287_n N_D_c_5288_n N_D_c_5289_n N_D_c_5291_n N_D_c_5376_n N_D_c_5356_n \
 N_D_c_5292_n N_D_c_5294_n N_D_c_5295_n N_D_c_5296_n N_D_c_5297_n N_D_c_5298_n \
 N_D_c_5299_n N_D_c_5301_n N_D_c_5400_n N_D_c_5358_n N_D_c_5302_n N_D_c_5304_n \
 N_D_c_5305_n N_D_c_5306_n N_D_c_5307_n N_D_c_5308_n N_D_c_5309_n N_D_c_5311_n \
 N_D_c_5402_n N_D_c_5360_n )  PM_TMRDFFSNRNQNX1\%D
x_PM_TMRDFFSNRNQNX1\%noxref_15 ( N_noxref_15_c_5619_n N_noxref_15_c_5620_n \
 N_noxref_15_c_5621_n N_noxref_15_c_5622_n N_noxref_15_c_5648_n \
 N_noxref_15_c_5652_n N_noxref_15_c_5654_n N_noxref_15_c_5658_n \
 N_noxref_15_c_5623_n N_noxref_15_c_5792_p N_noxref_15_c_5624_n \
 N_noxref_15_c_5625_n N_noxref_15_c_5626_n N_noxref_15_c_5804_p \
 N_noxref_15_c_5761_p N_noxref_15_M39_noxref_g N_noxref_15_M42_noxref_g \
 N_noxref_15_M138_noxref_g N_noxref_15_M139_noxref_g N_noxref_15_M144_noxref_g \
 N_noxref_15_M145_noxref_g N_noxref_15_c_5627_n N_noxref_15_c_5629_n \
 N_noxref_15_c_5630_n N_noxref_15_c_5631_n N_noxref_15_c_5632_n \
 N_noxref_15_c_5633_n N_noxref_15_c_5634_n N_noxref_15_c_5636_n \
 N_noxref_15_c_5704_n N_noxref_15_c_5677_n N_noxref_15_c_5637_n \
 N_noxref_15_c_5639_n N_noxref_15_c_5640_n N_noxref_15_c_5641_n \
 N_noxref_15_c_5642_n N_noxref_15_c_5643_n N_noxref_15_c_5644_n \
 N_noxref_15_c_5646_n N_noxref_15_c_5706_n N_noxref_15_c_5679_n \
 N_noxref_15_M38_noxref_d N_noxref_15_M132_noxref_d N_noxref_15_M134_noxref_d \
 N_noxref_15_M136_noxref_d )  PM_TMRDFFSNRNQNX1\%noxref_15
x_PM_TMRDFFSNRNQNX1\%noxref_16 ( N_noxref_16_c_5872_n N_noxref_16_c_5873_n \
 N_noxref_16_c_5888_n N_noxref_16_c_5892_n N_noxref_16_c_5894_n \
 N_noxref_16_c_5898_n N_noxref_16_c_5874_n N_noxref_16_c_5971_p \
 N_noxref_16_c_5875_n N_noxref_16_c_5876_n N_noxref_16_c_5986_p \
 N_noxref_16_c_5994_p N_noxref_16_M45_noxref_g N_noxref_16_M150_noxref_g \
 N_noxref_16_M151_noxref_g N_noxref_16_c_5877_n N_noxref_16_c_5879_n \
 N_noxref_16_c_5880_n N_noxref_16_c_5881_n N_noxref_16_c_5882_n \
 N_noxref_16_c_5883_n N_noxref_16_c_5884_n N_noxref_16_c_5886_n \
 N_noxref_16_c_5932_n N_noxref_16_c_5910_n N_noxref_16_M44_noxref_d \
 N_noxref_16_M144_noxref_d N_noxref_16_M146_noxref_d N_noxref_16_M148_noxref_d \
 )  PM_TMRDFFSNRNQNX1\%noxref_16
x_PM_TMRDFFSNRNQNX1\%CLK ( N_CLK_c_6046_n N_CLK_c_6057_n N_CLK_c_6058_n \
 N_CLK_c_6067_n N_CLK_c_6068_n N_CLK_c_6190_n N_CLK_c_6070_n N_CLK_c_6192_n \
 N_CLK_c_6074_n N_CLK_c_6196_n CLK CLK CLK CLK CLK CLK CLK CLK CLK CLK CLK CLK \
 N_CLK_c_6040_n N_CLK_c_6041_n N_CLK_c_6042_n N_CLK_c_6043_n N_CLK_c_6044_n \
 N_CLK_c_6045_n N_CLK_M4_noxref_g N_CLK_M10_noxref_g N_CLK_M22_noxref_g \
 N_CLK_M28_noxref_g N_CLK_M40_noxref_g N_CLK_M46_noxref_g N_CLK_M68_noxref_g \
 N_CLK_M69_noxref_g N_CLK_M80_noxref_g N_CLK_M81_noxref_g N_CLK_M104_noxref_g \
 N_CLK_M105_noxref_g N_CLK_M116_noxref_g N_CLK_M117_noxref_g \
 N_CLK_M140_noxref_g N_CLK_M141_noxref_g N_CLK_M152_noxref_g \
 N_CLK_M153_noxref_g N_CLK_c_6121_n N_CLK_c_6124_n N_CLK_c_6635_p \
 N_CLK_c_6642_p N_CLK_c_6126_n N_CLK_c_6127_n N_CLK_c_6128_n N_CLK_c_6129_n \
 N_CLK_c_6179_n N_CLK_c_6150_n N_CLK_c_6153_n N_CLK_c_6655_p N_CLK_c_6662_p \
 N_CLK_c_6155_n N_CLK_c_6156_n N_CLK_c_6157_n N_CLK_c_6158_n N_CLK_c_6261_n \
 N_CLK_c_6285_n N_CLK_c_6288_n N_CLK_c_6675_p N_CLK_c_6682_p N_CLK_c_6290_n \
 N_CLK_c_6291_n N_CLK_c_6292_n N_CLK_c_6293_n N_CLK_c_6211_n N_CLK_c_6311_n \
 N_CLK_c_6314_n N_CLK_c_6695_p N_CLK_c_6702_p N_CLK_c_6316_n N_CLK_c_6317_n \
 N_CLK_c_6318_n N_CLK_c_6319_n N_CLK_c_6212_n N_CLK_c_6421_n N_CLK_c_6424_n \
 N_CLK_c_6715_p N_CLK_c_6722_p N_CLK_c_6426_n N_CLK_c_6427_n N_CLK_c_6428_n \
 N_CLK_c_6429_n N_CLK_c_6213_n N_CLK_c_6446_n N_CLK_c_6449_n N_CLK_c_6735_p \
 N_CLK_c_6742_p N_CLK_c_6451_n N_CLK_c_6452_n N_CLK_c_6453_n N_CLK_c_6454_n \
 N_CLK_c_6214_n N_CLK_c_6131_n N_CLK_c_6160_n N_CLK_c_6215_n N_CLK_c_6216_n \
 N_CLK_c_6217_n N_CLK_c_6218_n )  PM_TMRDFFSNRNQNX1\%CLK
x_PM_TMRDFFSNRNQNX1\%noxref_18 ( N_noxref_18_c_6814_n N_noxref_18_c_6820_n \
 N_noxref_18_c_6821_n N_noxref_18_c_6823_n N_noxref_18_c_6747_n \
 N_noxref_18_c_6762_n N_noxref_18_c_6766_n N_noxref_18_c_6768_n \
 N_noxref_18_c_6772_n N_noxref_18_c_6748_n N_noxref_18_c_6881_p \
 N_noxref_18_c_6776_n N_noxref_18_c_6749_n N_noxref_18_c_6873_n \
 N_noxref_18_c_6956_p N_noxref_18_M38_noxref_g N_noxref_18_M48_noxref_g \
 N_noxref_18_M136_noxref_g N_noxref_18_M137_noxref_g N_noxref_18_M156_noxref_g \
 N_noxref_18_M157_noxref_g N_noxref_18_c_6839_n N_noxref_18_c_6840_n \
 N_noxref_18_c_6841_n N_noxref_18_c_6842_n N_noxref_18_c_6843_n \
 N_noxref_18_c_6845_n N_noxref_18_c_6846_n N_noxref_18_c_6750_n \
 N_noxref_18_c_6752_n N_noxref_18_c_6753_n N_noxref_18_c_6754_n \
 N_noxref_18_c_6755_n N_noxref_18_c_6756_n N_noxref_18_c_6757_n \
 N_noxref_18_c_6759_n N_noxref_18_c_6900_p N_noxref_18_c_6788_n \
 N_noxref_18_c_6848_n N_noxref_18_c_6849_n N_noxref_18_c_6812_n \
 N_noxref_18_M41_noxref_d N_noxref_18_M138_noxref_d N_noxref_18_M140_noxref_d \
 N_noxref_18_M142_noxref_d )  PM_TMRDFFSNRNQNX1\%noxref_18
x_PM_TMRDFFSNRNQNX1\%RN ( N_RN_c_7021_n N_RN_c_7032_n N_RN_c_7033_n \
 N_RN_c_7037_n N_RN_c_7038_n N_RN_c_7045_n N_RN_c_7046_n N_RN_c_7057_n \
 N_RN_c_7058_n N_RN_c_7062_n N_RN_c_7063_n N_RN_c_7070_n N_RN_c_7071_n \
 N_RN_c_7082_n N_RN_c_7083_n N_RN_c_7087_n RN RN RN RN RN RN RN RN RN RN RN RN \
 RN RN RN RN RN RN RN RN RN RN RN RN RN RN RN RN RN N_RN_c_7088_n \
 N_RN_c_7089_n N_RN_c_7090_n N_RN_c_7091_n N_RN_c_7092_n N_RN_c_7093_n \
 N_RN_c_7094_n N_RN_c_7095_n N_RN_c_7096_n N_RN_M1_noxref_g N_RN_M11_noxref_g \
 N_RN_M13_noxref_g N_RN_M19_noxref_g N_RN_M29_noxref_g N_RN_M31_noxref_g \
 N_RN_M37_noxref_g N_RN_M47_noxref_g N_RN_M49_noxref_g N_RN_M62_noxref_g \
 N_RN_M63_noxref_g N_RN_M82_noxref_g N_RN_M83_noxref_g N_RN_M86_noxref_g \
 N_RN_M87_noxref_g N_RN_M98_noxref_g N_RN_M99_noxref_g N_RN_M118_noxref_g \
 N_RN_M119_noxref_g N_RN_M122_noxref_g N_RN_M123_noxref_g N_RN_M134_noxref_g \
 N_RN_M135_noxref_g N_RN_M154_noxref_g N_RN_M155_noxref_g N_RN_M158_noxref_g \
 N_RN_M159_noxref_g N_RN_c_7528_n N_RN_c_7531_n N_RN_c_7864_p N_RN_c_7872_p \
 N_RN_c_7204_n N_RN_c_7205_n N_RN_c_7206_n N_RN_c_7207_n N_RN_c_7161_n \
 N_RN_c_7295_n N_RN_c_7296_n N_RN_c_7297_n N_RN_c_7298_n N_RN_c_7299_n \
 N_RN_c_7301_n N_RN_c_7302_n N_RN_c_7211_n N_RN_c_7214_n N_RN_c_7925_p \
 N_RN_c_7933_p N_RN_c_7216_n N_RN_c_7217_n N_RN_c_7218_n N_RN_c_7219_n \
 N_RN_c_7255_n N_RN_c_7539_n N_RN_c_7542_n N_RN_c_7962_p N_RN_c_7970_p \
 N_RN_c_7394_n N_RN_c_7395_n N_RN_c_7396_n N_RN_c_7397_n N_RN_c_7256_n \
 N_RN_c_7441_n N_RN_c_7442_n N_RN_c_7443_n N_RN_c_7444_n N_RN_c_7445_n \
 N_RN_c_7447_n N_RN_c_7448_n N_RN_c_7401_n N_RN_c_7404_n N_RN_c_8023_p \
 N_RN_c_8031_p N_RN_c_7406_n N_RN_c_7407_n N_RN_c_7408_n N_RN_c_7409_n \
 N_RN_c_7257_n N_RN_c_7549_n N_RN_c_7552_n N_RN_c_8060_p N_RN_c_8068_p \
 N_RN_c_7554_n N_RN_c_7555_n N_RN_c_7556_n N_RN_c_7557_n N_RN_c_7258_n \
 N_RN_c_7649_n N_RN_c_7650_n N_RN_c_7651_n N_RN_c_7800_p N_RN_c_7781_p \
 N_RN_c_7802_p N_RN_c_7782_p N_RN_c_7714_n N_RN_c_7717_n N_RN_c_8117_p \
 N_RN_c_8124_p N_RN_c_7719_n N_RN_c_7720_n N_RN_c_7721_n N_RN_c_7722_n \
 N_RN_c_7259_n N_RN_c_7162_n N_RN_c_7304_n N_RN_c_7305_n N_RN_c_7307_n \
 N_RN_c_7223_n N_RN_c_7261_n N_RN_c_7450_n N_RN_c_7451_n N_RN_c_7262_n \
 N_RN_c_7263_n N_RN_c_7264_n N_RN_c_7670_n N_RN_c_7672_n N_RN_c_7265_n \
 N_RN_c_7268_n )  PM_TMRDFFSNRNQNX1\%RN
x_PM_TMRDFFSNRNQNX1\%SN ( N_SN_c_8129_n N_SN_c_8183_n N_SN_c_8132_n \
 N_SN_c_8226_n N_SN_c_8135_n N_SN_c_8340_n N_SN_c_8138_n N_SN_c_8399_n \
 N_SN_c_8141_n N_SN_c_8468_n SN SN SN SN SN SN SN SN SN N_SN_c_8145_n \
 N_SN_c_8146_n N_SN_c_8147_n N_SN_c_8148_n N_SN_c_8149_n N_SN_c_8150_n \
 N_SN_M7_noxref_g N_SN_M16_noxref_g N_SN_M25_noxref_g N_SN_M34_noxref_g \
 N_SN_M43_noxref_g N_SN_M52_noxref_g N_SN_M74_noxref_g N_SN_M75_noxref_g \
 N_SN_M92_noxref_g N_SN_M93_noxref_g N_SN_M110_noxref_g N_SN_M111_noxref_g \
 N_SN_M128_noxref_g N_SN_M129_noxref_g N_SN_M146_noxref_g N_SN_M147_noxref_g \
 N_SN_M164_noxref_g N_SN_M165_noxref_g N_SN_c_8192_n N_SN_c_8195_n \
 N_SN_c_8712_p N_SN_c_8719_p N_SN_c_8197_n N_SN_c_8198_n N_SN_c_8199_n \
 N_SN_c_8200_n N_SN_c_8215_n N_SN_c_8249_n N_SN_c_8252_n N_SN_c_8732_p \
 N_SN_c_8739_p N_SN_c_8254_n N_SN_c_8255_n N_SN_c_8256_n N_SN_c_8257_n \
 N_SN_c_8259_n N_SN_c_8349_n N_SN_c_8352_n N_SN_c_8752_p N_SN_c_8759_p \
 N_SN_c_8354_n N_SN_c_8355_n N_SN_c_8356_n N_SN_c_8357_n N_SN_c_8260_n \
 N_SN_c_8690_p N_SN_c_8692_p N_SN_c_8772_p N_SN_c_8779_p N_SN_c_8423_n \
 N_SN_c_8424_n N_SN_c_8425_n N_SN_c_8426_n N_SN_c_8261_n N_SN_c_8477_n \
 N_SN_c_8480_n N_SN_c_8792_p N_SN_c_8799_p N_SN_c_8482_n N_SN_c_8483_n \
 N_SN_c_8484_n N_SN_c_8485_n N_SN_c_8262_n N_SN_c_8653_p N_SN_c_8655_p \
 N_SN_c_8816_p N_SN_c_8823_p N_SN_c_8609_p N_SN_c_8610_p N_SN_c_8611_p \
 N_SN_c_8598_p N_SN_c_8263_n N_SN_c_8202_n N_SN_c_8264_n N_SN_c_8268_n \
 N_SN_c_8269_n N_SN_c_8270_n N_SN_c_8271_n )  PM_TMRDFFSNRNQNX1\%SN
x_PM_TMRDFFSNRNQNX1\%noxref_21 ( N_noxref_21_c_8898_n N_noxref_21_c_8935_n \
 N_noxref_21_c_8878_n N_noxref_21_c_8905_n N_noxref_21_c_8880_n \
 N_noxref_21_c_8881_n N_noxref_21_c_8828_n N_noxref_21_c_8829_n \
 N_noxref_21_c_8835_n N_noxref_21_c_8839_n N_noxref_21_c_8841_n \
 N_noxref_21_c_8845_n N_noxref_21_c_8830_n N_noxref_21_c_9017_n \
 N_noxref_21_c_8849_n N_noxref_21_c_8831_n N_noxref_21_c_8951_n \
 N_noxref_21_c_9025_n N_noxref_21_M41_noxref_g N_noxref_21_M44_noxref_g \
 N_noxref_21_M53_noxref_g N_noxref_21_M142_noxref_g N_noxref_21_M143_noxref_g \
 N_noxref_21_M148_noxref_g N_noxref_21_M149_noxref_g N_noxref_21_M166_noxref_g \
 N_noxref_21_M167_noxref_g N_noxref_21_c_8955_n N_noxref_21_c_8956_n \
 N_noxref_21_c_8957_n N_noxref_21_c_8994_n N_noxref_21_c_8995_n \
 N_noxref_21_c_8997_n N_noxref_21_c_8998_n N_noxref_21_c_8918_n \
 N_noxref_21_c_8919_n N_noxref_21_c_8920_n N_noxref_21_c_8921_n \
 N_noxref_21_c_8922_n N_noxref_21_c_8924_n N_noxref_21_c_8925_n \
 N_noxref_21_c_9072_n N_noxref_21_c_9073_n N_noxref_21_c_9074_n \
 N_noxref_21_c_9106_p N_noxref_21_c_9094_p N_noxref_21_c_9108_p \
 N_noxref_21_c_9095_p N_noxref_21_c_8958_n N_noxref_21_c_8960_n \
 N_noxref_21_c_8895_n N_noxref_21_c_8927_n N_noxref_21_c_8928_n \
 N_noxref_21_c_8896_n N_noxref_21_c_9081_n N_noxref_21_c_9083_n \
 N_noxref_21_c_8897_n N_noxref_21_M47_noxref_d N_noxref_21_M150_noxref_d \
 N_noxref_21_M152_noxref_d N_noxref_21_M154_noxref_d )  \
 PM_TMRDFFSNRNQNX1\%noxref_21
x_PM_TMRDFFSNRNQNX1\%noxref_22 ( N_noxref_22_c_9171_n N_noxref_22_c_9174_n \
 N_noxref_22_c_9175_n N_noxref_22_c_9180_n N_noxref_22_c_9184_n \
 N_noxref_22_c_9186_n N_noxref_22_c_9190_n N_noxref_22_c_9176_n \
 N_noxref_22_c_9285_p N_noxref_22_c_9177_n N_noxref_22_c_9251_n \
 N_noxref_22_c_9268_n N_noxref_22_M50_noxref_g N_noxref_22_M160_noxref_g \
 N_noxref_22_M161_noxref_g N_noxref_22_c_9232_n N_noxref_22_c_9233_n \
 N_noxref_22_c_9234_n N_noxref_22_c_9312_p N_noxref_22_c_9292_p \
 N_noxref_22_c_9314_p N_noxref_22_c_9293_p N_noxref_22_c_9235_n \
 N_noxref_22_c_9238_n N_noxref_22_c_9222_n N_noxref_22_M53_noxref_d \
 N_noxref_22_M162_noxref_d N_noxref_22_M164_noxref_d N_noxref_22_M166_noxref_d \
 )  PM_TMRDFFSNRNQNX1\%noxref_22
x_PM_TMRDFFSNRNQNX1\%noxref_23 ( N_noxref_23_c_9342_n N_noxref_23_c_9348_n \
 N_noxref_23_c_9353_n N_noxref_23_c_9357_n N_noxref_23_c_9359_n \
 N_noxref_23_c_9362_n N_noxref_23_c_9388_n N_noxref_23_c_9364_n \
 N_noxref_23_c_9395_p N_noxref_23_M168_noxref_d N_noxref_23_M170_noxref_d \
 N_noxref_23_M172_noxref_s N_noxref_23_M173_noxref_d N_noxref_23_M175_noxref_d \
 )  PM_TMRDFFSNRNQNX1\%noxref_23
x_PM_TMRDFFSNRNQNX1\%noxref_24 ( N_noxref_24_c_9433_n N_noxref_24_c_9437_n \
 N_noxref_24_c_9440_n N_noxref_24_c_9446_n N_noxref_24_c_9448_n \
 N_noxref_24_c_9449_n N_noxref_24_c_9478_n N_noxref_24_c_9482_n \
 N_noxref_24_c_9484_n N_noxref_24_c_9488_n N_noxref_24_c_9450_n \
 N_noxref_24_c_9630_n N_noxref_24_c_9451_n N_noxref_24_c_9452_n \
 N_noxref_24_c_9453_n N_noxref_24_c_9455_n N_noxref_24_c_9574_n \
 N_noxref_24_c_9639_n N_noxref_24_M51_noxref_g N_noxref_24_M57_noxref_g \
 N_noxref_24_M58_noxref_g N_noxref_24_M162_noxref_g N_noxref_24_M163_noxref_g \
 N_noxref_24_M174_noxref_g N_noxref_24_M175_noxref_g N_noxref_24_M176_noxref_g \
 N_noxref_24_M177_noxref_g N_noxref_24_c_9456_n N_noxref_24_c_9458_n \
 N_noxref_24_c_9459_n N_noxref_24_c_9460_n N_noxref_24_c_9461_n \
 N_noxref_24_c_9462_n N_noxref_24_c_9463_n N_noxref_24_c_9465_n \
 N_noxref_24_c_9604_n N_noxref_24_c_9509_n N_noxref_24_c_9550_n \
 N_noxref_24_c_9553_n N_noxref_24_c_9675_p N_noxref_24_c_9555_n \
 N_noxref_24_c_9742_p N_noxref_24_c_9743_p N_noxref_24_c_9511_n \
 N_noxref_24_c_9559_n N_noxref_24_c_9560_n N_noxref_24_c_9561_n \
 N_noxref_24_c_9466_n N_noxref_24_c_9467_n N_noxref_24_c_9469_n \
 N_noxref_24_c_9709_p N_noxref_24_c_9470_n N_noxref_24_c_9471_n \
 N_noxref_24_c_9472_n N_noxref_24_c_9699_p N_noxref_24_c_9512_n \
 N_noxref_24_c_9473_n N_noxref_24_c_9475_n N_noxref_24_c_9476_n \
 N_noxref_24_M50_noxref_d N_noxref_24_M156_noxref_d N_noxref_24_M158_noxref_d \
 N_noxref_24_M160_noxref_d )  PM_TMRDFFSNRNQNX1\%noxref_24
x_PM_TMRDFFSNRNQNX1\%noxref_25 ( N_noxref_25_c_9823_n N_noxref_25_c_9827_n \
 N_noxref_25_c_9838_n N_noxref_25_c_9829_n N_noxref_25_c_9830_n \
 N_noxref_25_c_9831_n N_noxref_25_c_9882_n N_noxref_25_c_9833_n \
 N_noxref_25_c_9893_p N_noxref_25_M172_noxref_d N_noxref_25_M174_noxref_d \
 N_noxref_25_M176_noxref_s N_noxref_25_M177_noxref_d N_noxref_25_M179_noxref_d \
 )  PM_TMRDFFSNRNQNX1\%noxref_25
x_PM_TMRDFFSNRNQNX1\%noxref_26 ( N_noxref_26_c_10048_n N_noxref_26_c_10043_n \
 N_noxref_26_c_10050_n N_noxref_26_c_10052_n N_noxref_26_c_10053_n \
 N_noxref_26_c_9933_n N_noxref_26_c_10055_n N_noxref_26_c_10119_n \
 N_noxref_26_c_9912_n N_noxref_26_c_10001_n N_noxref_26_c_9913_n \
 N_noxref_26_c_9943_n N_noxref_26_c_9944_n N_noxref_26_c_9948_n \
 N_noxref_26_c_9950_n N_noxref_26_c_9954_n N_noxref_26_c_9915_n \
 N_noxref_26_c_10146_n N_noxref_26_c_9958_n N_noxref_26_c_9916_n \
 N_noxref_26_c_9962_n N_noxref_26_c_9917_n N_noxref_26_c_9919_n \
 N_noxref_26_c_10150_n N_noxref_26_c_10083_n N_noxref_26_c_10237_n \
 N_noxref_26_M33_noxref_g N_noxref_26_M55_noxref_g N_noxref_26_M59_noxref_g \
 N_noxref_26_M126_noxref_g N_noxref_26_M127_noxref_g N_noxref_26_M170_noxref_g \
 N_noxref_26_M171_noxref_g N_noxref_26_M178_noxref_g N_noxref_26_M179_noxref_g \
 N_noxref_26_c_9921_n N_noxref_26_c_9923_n N_noxref_26_c_9924_n \
 N_noxref_26_c_9925_n N_noxref_26_c_9926_n N_noxref_26_c_9927_n \
 N_noxref_26_c_9928_n N_noxref_26_c_9930_n N_noxref_26_c_10024_n \
 N_noxref_26_c_9977_n N_noxref_26_c_10026_n N_noxref_26_c_10029_n \
 N_noxref_26_c_10031_n N_noxref_26_c_9979_n N_noxref_26_c_10280_p \
 N_noxref_26_c_10242_n N_noxref_26_c_10035_n N_noxref_26_c_10036_n \
 N_noxref_26_c_10243_n N_noxref_26_c_10246_n N_noxref_26_c_10247_n \
 N_noxref_26_c_10305_p N_noxref_26_c_10288_p N_noxref_26_c_10250_n \
 N_noxref_26_c_10251_n N_noxref_26_c_10252_n N_noxref_26_c_9931_n \
 N_noxref_26_c_10355_p N_noxref_26_c_9980_n N_noxref_26_c_10254_n \
 N_noxref_26_c_10301_p N_noxref_26_c_10257_n N_noxref_26_M32_noxref_d \
 N_noxref_26_M120_noxref_d N_noxref_26_M122_noxref_d N_noxref_26_M124_noxref_d \
 )  PM_TMRDFFSNRNQNX1\%noxref_26
x_PM_TMRDFFSNRNQNX1\%Q ( Q N_Q_c_10368_n N_Q_c_10375_n N_Q_c_10376_n \
 N_Q_c_10382_n N_Q_c_10433_n N_Q_c_10397_n N_Q_c_10398_n N_Q_c_10383_n \
 N_Q_c_10492_n N_Q_c_10384_n N_Q_c_10500_n N_Q_M55_noxref_d N_Q_M57_noxref_d \
 N_Q_M59_noxref_d N_Q_M176_noxref_d N_Q_M178_noxref_d )  PM_TMRDFFSNRNQNX1\%Q
x_PM_TMRDFFSNRNQNX1\%noxref_28 ( N_noxref_28_c_10558_n N_noxref_28_c_10542_n \
 N_noxref_28_c_10546_n N_noxref_28_c_10549_n N_noxref_28_c_10566_n \
 N_noxref_28_M0_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_28
x_PM_TMRDFFSNRNQNX1\%noxref_29 ( N_noxref_29_c_10591_n N_noxref_29_c_10593_n \
 N_noxref_29_c_10596_n N_noxref_29_c_10598_n N_noxref_29_c_10606_n \
 N_noxref_29_M1_noxref_d N_noxref_29_M2_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_29
x_PM_TMRDFFSNRNQNX1\%noxref_30 ( N_noxref_30_c_10658_n N_noxref_30_c_10643_n \
 N_noxref_30_c_10647_n N_noxref_30_c_10650_n N_noxref_30_c_10673_n \
 N_noxref_30_M3_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_30
x_PM_TMRDFFSNRNQNX1\%noxref_31 ( N_noxref_31_c_10692_n N_noxref_31_c_10694_n \
 N_noxref_31_c_10697_n N_noxref_31_c_10699_n N_noxref_31_c_10707_n \
 N_noxref_31_M4_noxref_d N_noxref_31_M5_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_31
x_PM_TMRDFFSNRNQNX1\%noxref_32 ( N_noxref_32_c_10759_n N_noxref_32_c_10744_n \
 N_noxref_32_c_10748_n N_noxref_32_c_10751_n N_noxref_32_c_10774_n \
 N_noxref_32_M6_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_32
x_PM_TMRDFFSNRNQNX1\%noxref_33 ( N_noxref_33_c_10793_n N_noxref_33_c_10795_n \
 N_noxref_33_c_10798_n N_noxref_33_c_10800_n N_noxref_33_c_10808_n \
 N_noxref_33_M7_noxref_d N_noxref_33_M8_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_33
x_PM_TMRDFFSNRNQNX1\%noxref_34 ( N_noxref_34_c_10860_n N_noxref_34_c_10845_n \
 N_noxref_34_c_10849_n N_noxref_34_c_10852_n N_noxref_34_c_10875_n \
 N_noxref_34_M9_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_34
x_PM_TMRDFFSNRNQNX1\%noxref_35 ( N_noxref_35_c_10894_n N_noxref_35_c_10896_n \
 N_noxref_35_c_10899_n N_noxref_35_c_10901_n N_noxref_35_c_10909_n \
 N_noxref_35_M10_noxref_d N_noxref_35_M11_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_35
x_PM_TMRDFFSNRNQNX1\%noxref_36 ( N_noxref_36_c_10962_n N_noxref_36_c_10947_n \
 N_noxref_36_c_10951_n N_noxref_36_c_10954_n N_noxref_36_c_10979_n \
 N_noxref_36_M12_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_36
x_PM_TMRDFFSNRNQNX1\%noxref_37 ( N_noxref_37_c_10999_n N_noxref_37_c_11001_n \
 N_noxref_37_c_11004_n N_noxref_37_c_11006_n N_noxref_37_c_11014_n \
 N_noxref_37_M13_noxref_d N_noxref_37_M14_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_37
x_PM_TMRDFFSNRNQNX1\%noxref_38 ( N_noxref_38_c_11066_n N_noxref_38_c_11051_n \
 N_noxref_38_c_11055_n N_noxref_38_c_11058_n N_noxref_38_c_11081_n \
 N_noxref_38_M15_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_38
x_PM_TMRDFFSNRNQNX1\%noxref_39 ( N_noxref_39_c_11100_n N_noxref_39_c_11102_n \
 N_noxref_39_c_11105_n N_noxref_39_c_11107_n N_noxref_39_c_11117_n \
 N_noxref_39_M16_noxref_d N_noxref_39_M17_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_39
x_PM_TMRDFFSNRNQNX1\%noxref_40 ( N_noxref_40_c_11167_n N_noxref_40_c_11152_n \
 N_noxref_40_c_11156_n N_noxref_40_c_11159_n N_noxref_40_c_11184_n \
 N_noxref_40_M18_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_40
x_PM_TMRDFFSNRNQNX1\%noxref_41 ( N_noxref_41_c_11204_n N_noxref_41_c_11206_n \
 N_noxref_41_c_11209_n N_noxref_41_c_11211_n N_noxref_41_c_11219_n \
 N_noxref_41_M19_noxref_d N_noxref_41_M20_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_41
x_PM_TMRDFFSNRNQNX1\%noxref_42 ( N_noxref_42_c_11271_n N_noxref_42_c_11256_n \
 N_noxref_42_c_11260_n N_noxref_42_c_11263_n N_noxref_42_c_11286_n \
 N_noxref_42_M21_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_42
x_PM_TMRDFFSNRNQNX1\%noxref_43 ( N_noxref_43_c_11305_n N_noxref_43_c_11307_n \
 N_noxref_43_c_11310_n N_noxref_43_c_11312_n N_noxref_43_c_11320_n \
 N_noxref_43_M22_noxref_d N_noxref_43_M23_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_43
x_PM_TMRDFFSNRNQNX1\%noxref_44 ( N_noxref_44_c_11372_n N_noxref_44_c_11357_n \
 N_noxref_44_c_11361_n N_noxref_44_c_11364_n N_noxref_44_c_11387_n \
 N_noxref_44_M24_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_44
x_PM_TMRDFFSNRNQNX1\%noxref_45 ( N_noxref_45_c_11406_n N_noxref_45_c_11408_n \
 N_noxref_45_c_11411_n N_noxref_45_c_11413_n N_noxref_45_c_11421_n \
 N_noxref_45_M25_noxref_d N_noxref_45_M26_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_45
x_PM_TMRDFFSNRNQNX1\%noxref_46 ( N_noxref_46_c_11473_n N_noxref_46_c_11458_n \
 N_noxref_46_c_11462_n N_noxref_46_c_11465_n N_noxref_46_c_11488_n \
 N_noxref_46_M27_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_46
x_PM_TMRDFFSNRNQNX1\%noxref_47 ( N_noxref_47_c_11507_n N_noxref_47_c_11509_n \
 N_noxref_47_c_11512_n N_noxref_47_c_11514_n N_noxref_47_c_11522_n \
 N_noxref_47_M28_noxref_d N_noxref_47_M29_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_47
x_PM_TMRDFFSNRNQNX1\%noxref_48 ( N_noxref_48_c_11575_n N_noxref_48_c_11560_n \
 N_noxref_48_c_11564_n N_noxref_48_c_11567_n N_noxref_48_c_11591_n \
 N_noxref_48_M30_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_48
x_PM_TMRDFFSNRNQNX1\%noxref_49 ( N_noxref_49_c_11612_n N_noxref_49_c_11614_n \
 N_noxref_49_c_11617_n N_noxref_49_c_11619_n N_noxref_49_c_11629_n \
 N_noxref_49_M31_noxref_d N_noxref_49_M32_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_49
x_PM_TMRDFFSNRNQNX1\%noxref_50 ( N_noxref_50_c_11680_n N_noxref_50_c_11664_n \
 N_noxref_50_c_11668_n N_noxref_50_c_11671_n N_noxref_50_c_11682_n \
 N_noxref_50_M33_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_50
x_PM_TMRDFFSNRNQNX1\%noxref_51 ( N_noxref_51_c_11713_n N_noxref_51_c_11715_n \
 N_noxref_51_c_11718_n N_noxref_51_c_11720_n N_noxref_51_c_11730_n \
 N_noxref_51_M34_noxref_d N_noxref_51_M35_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_51
x_PM_TMRDFFSNRNQNX1\%noxref_52 ( N_noxref_52_c_11780_n N_noxref_52_c_11765_n \
 N_noxref_52_c_11769_n N_noxref_52_c_11772_n N_noxref_52_c_11797_n \
 N_noxref_52_M36_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_52
x_PM_TMRDFFSNRNQNX1\%noxref_53 ( N_noxref_53_c_11817_n N_noxref_53_c_11819_n \
 N_noxref_53_c_11822_n N_noxref_53_c_11824_n N_noxref_53_c_11832_n \
 N_noxref_53_M37_noxref_d N_noxref_53_M38_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_53
x_PM_TMRDFFSNRNQNX1\%noxref_54 ( N_noxref_54_c_11884_n N_noxref_54_c_11869_n \
 N_noxref_54_c_11873_n N_noxref_54_c_11876_n N_noxref_54_c_11898_n \
 N_noxref_54_M39_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_54
x_PM_TMRDFFSNRNQNX1\%noxref_55 ( N_noxref_55_c_11918_n N_noxref_55_c_11920_n \
 N_noxref_55_c_11923_n N_noxref_55_c_11925_n N_noxref_55_c_11945_n \
 N_noxref_55_M40_noxref_d N_noxref_55_M41_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_55
x_PM_TMRDFFSNRNQNX1\%noxref_56 ( N_noxref_56_c_11985_n N_noxref_56_c_11970_n \
 N_noxref_56_c_11974_n N_noxref_56_c_11977_n N_noxref_56_c_12000_n \
 N_noxref_56_M42_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_56
x_PM_TMRDFFSNRNQNX1\%noxref_57 ( N_noxref_57_c_12019_n N_noxref_57_c_12021_n \
 N_noxref_57_c_12024_n N_noxref_57_c_12026_n N_noxref_57_c_12034_n \
 N_noxref_57_M43_noxref_d N_noxref_57_M44_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_57
x_PM_TMRDFFSNRNQNX1\%noxref_58 ( N_noxref_58_c_12086_n N_noxref_58_c_12071_n \
 N_noxref_58_c_12075_n N_noxref_58_c_12078_n N_noxref_58_c_12100_n \
 N_noxref_58_M45_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_58
x_PM_TMRDFFSNRNQNX1\%noxref_59 ( N_noxref_59_c_12120_n N_noxref_59_c_12122_n \
 N_noxref_59_c_12125_n N_noxref_59_c_12127_n N_noxref_59_c_12152_n \
 N_noxref_59_M46_noxref_d N_noxref_59_M47_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_59
x_PM_TMRDFFSNRNQNX1\%noxref_60 ( N_noxref_60_c_12188_n N_noxref_60_c_12173_n \
 N_noxref_60_c_12177_n N_noxref_60_c_12180_n N_noxref_60_c_12202_n \
 N_noxref_60_M48_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_60
x_PM_TMRDFFSNRNQNX1\%noxref_61 ( N_noxref_61_c_12224_n N_noxref_61_c_12226_n \
 N_noxref_61_c_12229_n N_noxref_61_c_12231_n N_noxref_61_c_12257_n \
 N_noxref_61_M49_noxref_d N_noxref_61_M50_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_61
x_PM_TMRDFFSNRNQNX1\%noxref_62 ( N_noxref_62_c_12302_n N_noxref_62_c_12278_n \
 N_noxref_62_c_12282_n N_noxref_62_c_12285_n N_noxref_62_c_12295_n \
 N_noxref_62_M51_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_62
x_PM_TMRDFFSNRNQNX1\%noxref_63 ( N_noxref_63_c_12329_n N_noxref_63_c_12331_n \
 N_noxref_63_c_12334_n N_noxref_63_c_12336_n N_noxref_63_c_12358_n \
 N_noxref_63_M52_noxref_d N_noxref_63_M53_noxref_s )  \
 PM_TMRDFFSNRNQNX1\%noxref_63
x_PM_TMRDFFSNRNQNX1\%noxref_64 ( N_noxref_64_c_12399_n N_noxref_64_c_12381_n \
 N_noxref_64_c_12385_n N_noxref_64_c_12388_n N_noxref_64_c_12389_n \
 N_noxref_64_c_12391_n N_noxref_64_M54_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_64
x_PM_TMRDFFSNRNQNX1\%noxref_65 ( N_noxref_65_c_12455_n N_noxref_65_c_12438_n \
 N_noxref_65_c_12441_n N_noxref_65_c_12444_n N_noxref_65_c_12445_n \
 N_noxref_65_c_12447_n N_noxref_65_M56_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_65
x_PM_TMRDFFSNRNQNX1\%noxref_66 ( N_noxref_66_c_12509_n N_noxref_66_c_12493_n \
 N_noxref_66_c_12496_n N_noxref_66_c_12499_n N_noxref_66_c_12500_n \
 N_noxref_66_c_12502_n N_noxref_66_M58_noxref_s )  PM_TMRDFFSNRNQNX1\%noxref_66
cc_1 ( N_GND_c_1_p N_VDD_c_1063_n ) capacitor c=0.00989031f //x=0.74 //y=0 \
 //x2=0.74 //y2=7.4
cc_2 ( N_GND_c_2_p N_VDD_c_1064_n ) capacitor c=0.00989031f //x=95.83 //y=0 \
 //x2=95.83 //y2=7.4
cc_3 ( N_GND_c_3_p N_VDD_c_1065_n ) capacitor c=0.00576465f //x=4.81 //y=0 \
 //x2=4.81 //y2=7.4
cc_4 ( N_GND_c_4_p N_VDD_c_1066_n ) capacitor c=0.0057235f //x=9.62 //y=0 \
 //x2=9.62 //y2=7.4
cc_5 ( N_GND_c_5_p N_VDD_c_1067_n ) capacitor c=0.0057235f //x=14.43 //y=0 \
 //x2=14.43 //y2=7.4
cc_6 ( N_GND_c_6_p N_VDD_c_1068_n ) capacitor c=0.00474727f //x=19.24 //y=0 \
 //x2=19.24 //y2=7.4
cc_7 ( N_GND_c_7_p N_VDD_c_1069_n ) capacitor c=0.0057235f //x=24.05 //y=0 \
 //x2=24.05 //y2=7.4
cc_8 ( N_GND_c_8_p N_VDD_c_1070_n ) capacitor c=0.00482014f //x=28.86 //y=0 \
 //x2=28.86 //y2=7.4
cc_9 ( N_GND_c_9_p N_VDD_c_1071_n ) capacitor c=0.00576465f //x=33.67 //y=0 \
 //x2=33.67 //y2=7.4
cc_10 ( N_GND_c_10_p N_VDD_c_1072_n ) capacitor c=0.0057235f //x=38.48 //y=0 \
 //x2=38.48 //y2=7.4
cc_11 ( N_GND_c_11_p N_VDD_c_1073_n ) capacitor c=0.0057235f //x=43.29 //y=0 \
 //x2=43.29 //y2=7.4
cc_12 ( N_GND_c_12_p N_VDD_c_1074_n ) capacitor c=0.00474727f //x=48.1 //y=0 \
 //x2=48.1 //y2=7.4
cc_13 ( N_GND_c_13_p N_VDD_c_1075_n ) capacitor c=0.0057235f //x=52.91 //y=0 \
 //x2=52.91 //y2=7.4
cc_14 ( N_GND_c_14_p N_VDD_c_1076_n ) capacitor c=0.00474727f //x=57.72 //y=0 \
 //x2=57.72 //y2=7.4
cc_15 ( N_GND_c_15_p N_VDD_c_1077_n ) capacitor c=0.00989031f //x=62.53 //y=0 \
 //x2=62.53 //y2=7.4
cc_16 ( N_GND_c_16_p N_VDD_c_1078_n ) capacitor c=0.0057235f //x=67.34 //y=0 \
 //x2=67.34 //y2=7.4
cc_17 ( N_GND_c_17_p N_VDD_c_1079_n ) capacitor c=0.0057235f //x=72.15 //y=0 \
 //x2=72.15 //y2=7.4
cc_18 ( N_GND_c_18_p N_VDD_c_1080_n ) capacitor c=0.00474727f //x=76.96 //y=0 \
 //x2=76.96 //y2=7.4
cc_19 ( N_GND_c_19_p N_VDD_c_1081_n ) capacitor c=0.0057235f //x=81.77 //y=0 \
 //x2=81.77 //y2=7.4
cc_20 ( N_GND_c_20_p N_VDD_c_1082_n ) capacitor c=0.00553002f //x=86.58 //y=0 \
 //x2=86.58 //y2=7.4
cc_21 ( N_GND_c_21_p N_VDD_c_1083_n ) capacitor c=0.00553002f //x=89.91 //y=0 \
 //x2=89.91 //y2=7.4
cc_22 ( N_GND_c_22_p N_VDD_c_1084_n ) capacitor c=0.00553669f //x=93.24 //y=0 \
 //x2=93.24 //y2=7.4
cc_23 ( N_GND_c_3_p N_noxref_3_c_2221_n ) capacitor c=0.0238274f //x=4.81 \
 //y=0 //x2=5.805 //y2=2.59
cc_24 ( N_GND_c_3_p N_noxref_3_c_2222_n ) capacitor c=0.00102529f //x=4.81 \
 //y=0 //x2=4.185 //y2=2.59
cc_25 ( N_GND_c_4_p N_noxref_3_c_2223_n ) capacitor c=0.0253329f //x=9.62 \
 //y=0 //x2=10.615 //y2=2.59
cc_26 ( N_GND_c_3_p N_noxref_3_c_2224_n ) capacitor c=7.16565e-19 //x=4.81 \
 //y=0 //x2=6.035 //y2=2.59
cc_27 ( N_GND_c_3_p N_noxref_3_c_2225_n ) capacitor c=0.04008f //x=4.81 //y=0 \
 //x2=3.985 //y2=1.665
cc_28 ( N_GND_c_3_p N_noxref_3_c_2226_n ) capacitor c=5.56859e-19 //x=4.81 \
 //y=0 //x2=4.07 //y2=2.59
cc_29 ( N_GND_c_3_p N_noxref_3_c_2227_n ) capacitor c=0.0128021f //x=4.81 \
 //y=0 //x2=5.92 //y2=2.08
cc_30 ( N_GND_c_4_p N_noxref_3_c_2228_n ) capacitor c=0.0126655f //x=9.62 \
 //y=0 //x2=10.73 //y2=2.08
cc_31 ( N_GND_c_31_p N_noxref_3_c_2229_n ) capacitor c=0.00132755f //x=5.8 \
 //y=0 //x2=5.62 //y2=0.875
cc_32 ( N_GND_M3_noxref_d N_noxref_3_c_2229_n ) capacitor c=0.00211996f \
 //x=5.695 //y=0.875 //x2=5.62 //y2=0.875
cc_33 ( N_GND_M3_noxref_d N_noxref_3_c_2231_n ) capacitor c=0.00255985f \
 //x=5.695 //y=0.875 //x2=5.62 //y2=1.22
cc_34 ( N_GND_c_3_p N_noxref_3_c_2232_n ) capacitor c=0.00204716f //x=4.81 \
 //y=0 //x2=5.62 //y2=1.53
cc_35 ( N_GND_c_3_p N_noxref_3_c_2233_n ) capacitor c=0.0110952f //x=4.81 \
 //y=0 //x2=5.62 //y2=1.915
cc_36 ( N_GND_M3_noxref_d N_noxref_3_c_2234_n ) capacitor c=0.0131341f \
 //x=5.695 //y=0.875 //x2=5.995 //y2=0.72
cc_37 ( N_GND_M3_noxref_d N_noxref_3_c_2235_n ) capacitor c=0.00193146f \
 //x=5.695 //y=0.875 //x2=5.995 //y2=1.375
cc_38 ( N_GND_c_38_p N_noxref_3_c_2236_n ) capacitor c=0.00129018f //x=9.45 \
 //y=0 //x2=6.15 //y2=0.875
cc_39 ( N_GND_M3_noxref_d N_noxref_3_c_2236_n ) capacitor c=0.00257848f \
 //x=5.695 //y=0.875 //x2=6.15 //y2=0.875
cc_40 ( N_GND_M3_noxref_d N_noxref_3_c_2238_n ) capacitor c=0.00255985f \
 //x=5.695 //y=0.875 //x2=6.15 //y2=1.22
cc_41 ( N_GND_c_41_p N_noxref_3_c_2239_n ) capacitor c=0.00132755f //x=10.61 \
 //y=0 //x2=10.43 //y2=0.875
cc_42 ( N_GND_M6_noxref_d N_noxref_3_c_2239_n ) capacitor c=0.00211996f \
 //x=10.505 //y=0.875 //x2=10.43 //y2=0.875
cc_43 ( N_GND_M6_noxref_d N_noxref_3_c_2241_n ) capacitor c=0.00255985f \
 //x=10.505 //y=0.875 //x2=10.43 //y2=1.22
cc_44 ( N_GND_c_4_p N_noxref_3_c_2242_n ) capacitor c=0.00204716f //x=9.62 \
 //y=0 //x2=10.43 //y2=1.53
cc_45 ( N_GND_c_4_p N_noxref_3_c_2243_n ) capacitor c=0.0112696f //x=9.62 \
 //y=0 //x2=10.43 //y2=1.915
cc_46 ( N_GND_M6_noxref_d N_noxref_3_c_2244_n ) capacitor c=0.0131341f \
 //x=10.505 //y=0.875 //x2=10.805 //y2=0.72
cc_47 ( N_GND_M6_noxref_d N_noxref_3_c_2245_n ) capacitor c=0.00193146f \
 //x=10.505 //y=0.875 //x2=10.805 //y2=1.375
cc_48 ( N_GND_c_48_p N_noxref_3_c_2246_n ) capacitor c=0.00129018f //x=14.26 \
 //y=0 //x2=10.96 //y2=0.875
cc_49 ( N_GND_M6_noxref_d N_noxref_3_c_2246_n ) capacitor c=0.00257848f \
 //x=10.505 //y=0.875 //x2=10.96 //y2=0.875
cc_50 ( N_GND_M6_noxref_d N_noxref_3_c_2248_n ) capacitor c=0.00255985f \
 //x=10.505 //y=0.875 //x2=10.96 //y2=1.22
cc_51 ( N_GND_c_3_p N_noxref_3_M2_noxref_d ) capacitor c=0.00591582f //x=4.81 \
 //y=0 //x2=3.395 //y2=0.915
cc_52 ( N_GND_c_5_p N_noxref_4_c_2461_n ) capacitor c=0.0222748f //x=14.43 \
 //y=0 //x2=15.425 //y2=2.59
cc_53 ( N_GND_c_5_p N_noxref_4_c_2462_n ) capacitor c=0.00102529f //x=14.43 \
 //y=0 //x2=13.805 //y2=2.59
cc_54 ( N_GND_c_5_p N_noxref_4_c_2463_n ) capacitor c=0.0401826f //x=14.43 \
 //y=0 //x2=13.605 //y2=1.665
cc_55 ( N_GND_c_5_p N_noxref_4_c_2464_n ) capacitor c=5.56859e-19 //x=14.43 \
 //y=0 //x2=13.69 //y2=2.59
cc_56 ( N_GND_c_5_p N_noxref_4_c_2465_n ) capacitor c=0.0127664f //x=14.43 \
 //y=0 //x2=15.54 //y2=2.08
cc_57 ( N_GND_c_57_p N_noxref_4_c_2466_n ) capacitor c=0.00132755f //x=15.42 \
 //y=0 //x2=15.24 //y2=0.875
cc_58 ( N_GND_M9_noxref_d N_noxref_4_c_2466_n ) capacitor c=0.00211996f \
 //x=15.315 //y=0.875 //x2=15.24 //y2=0.875
cc_59 ( N_GND_M9_noxref_d N_noxref_4_c_2468_n ) capacitor c=0.00255985f \
 //x=15.315 //y=0.875 //x2=15.24 //y2=1.22
cc_60 ( N_GND_c_5_p N_noxref_4_c_2469_n ) capacitor c=0.00204716f //x=14.43 \
 //y=0 //x2=15.24 //y2=1.53
cc_61 ( N_GND_c_5_p N_noxref_4_c_2470_n ) capacitor c=0.0110952f //x=14.43 \
 //y=0 //x2=15.24 //y2=1.915
cc_62 ( N_GND_M9_noxref_d N_noxref_4_c_2471_n ) capacitor c=0.0131341f \
 //x=15.315 //y=0.875 //x2=15.615 //y2=0.72
cc_63 ( N_GND_M9_noxref_d N_noxref_4_c_2472_n ) capacitor c=0.00193146f \
 //x=15.315 //y=0.875 //x2=15.615 //y2=1.375
cc_64 ( N_GND_c_64_p N_noxref_4_c_2473_n ) capacitor c=0.00129018f //x=19.07 \
 //y=0 //x2=15.77 //y2=0.875
cc_65 ( N_GND_M9_noxref_d N_noxref_4_c_2473_n ) capacitor c=0.00257848f \
 //x=15.315 //y=0.875 //x2=15.77 //y2=0.875
cc_66 ( N_GND_M9_noxref_d N_noxref_4_c_2475_n ) capacitor c=0.00255985f \
 //x=15.315 //y=0.875 //x2=15.77 //y2=1.22
cc_67 ( N_GND_c_5_p N_noxref_4_M8_noxref_d ) capacitor c=0.00591582f //x=14.43 \
 //y=0 //x2=13.015 //y2=0.915
cc_68 ( N_GND_c_3_p N_noxref_5_c_2626_n ) capacitor c=0.00505527f //x=4.81 \
 //y=0 //x2=8.765 //y2=3.33
cc_69 ( N_GND_c_4_p N_noxref_5_c_2627_n ) capacitor c=0.00505527f //x=9.62 \
 //y=0 //x2=20.235 //y2=3.33
cc_70 ( N_GND_c_3_p N_noxref_5_c_2628_n ) capacitor c=0.00101012f //x=4.81 \
 //y=0 //x2=3.33 //y2=2.08
cc_71 ( N_GND_c_4_p N_noxref_5_c_2629_n ) capacitor c=0.0405987f //x=9.62 \
 //y=0 //x2=8.795 //y2=1.665
cc_72 ( N_GND_c_6_p N_noxref_5_c_2630_n ) capacitor c=0.0155796f //x=19.24 \
 //y=0 //x2=20.35 //y2=2.08
cc_73 ( N_GND_c_73_p N_noxref_5_c_2631_n ) capacitor c=0.00132755f //x=20.23 \
 //y=0 //x2=20.05 //y2=0.875
cc_74 ( N_GND_M12_noxref_d N_noxref_5_c_2631_n ) capacitor c=0.00211996f \
 //x=20.125 //y=0.875 //x2=20.05 //y2=0.875
cc_75 ( N_GND_M12_noxref_d N_noxref_5_c_2633_n ) capacitor c=0.00255985f \
 //x=20.125 //y=0.875 //x2=20.05 //y2=1.22
cc_76 ( N_GND_c_6_p N_noxref_5_c_2634_n ) capacitor c=0.00204716f //x=19.24 \
 //y=0 //x2=20.05 //y2=1.53
cc_77 ( N_GND_c_6_p N_noxref_5_c_2635_n ) capacitor c=0.0110952f //x=19.24 \
 //y=0 //x2=20.05 //y2=1.915
cc_78 ( N_GND_M12_noxref_d N_noxref_5_c_2636_n ) capacitor c=0.0131341f \
 //x=20.125 //y=0.875 //x2=20.425 //y2=0.72
cc_79 ( N_GND_M12_noxref_d N_noxref_5_c_2637_n ) capacitor c=0.00193146f \
 //x=20.125 //y=0.875 //x2=20.425 //y2=1.375
cc_80 ( N_GND_c_80_p N_noxref_5_c_2638_n ) capacitor c=0.00129018f //x=23.88 \
 //y=0 //x2=20.58 //y2=0.875
cc_81 ( N_GND_M12_noxref_d N_noxref_5_c_2638_n ) capacitor c=0.00257848f \
 //x=20.125 //y=0.875 //x2=20.58 //y2=0.875
cc_82 ( N_GND_M12_noxref_d N_noxref_5_c_2640_n ) capacitor c=0.00255985f \
 //x=20.125 //y=0.875 //x2=20.58 //y2=1.22
cc_83 ( N_GND_c_4_p N_noxref_5_M5_noxref_d ) capacitor c=0.00591582f //x=9.62 \
 //y=0 //x2=8.205 //y2=0.915
cc_84 ( N_GND_c_7_p N_noxref_6_c_2893_n ) capacitor c=0.0222748f //x=24.05 \
 //y=0 //x2=25.045 //y2=2.59
cc_85 ( N_GND_c_7_p N_noxref_6_c_2894_n ) capacitor c=0.00102529f //x=24.05 \
 //y=0 //x2=23.425 //y2=2.59
cc_86 ( N_GND_c_7_p N_noxref_6_c_2895_n ) capacitor c=0.04008f //x=24.05 //y=0 \
 //x2=23.225 //y2=1.665
cc_87 ( N_GND_c_7_p N_noxref_6_c_2896_n ) capacitor c=5.56859e-19 //x=24.05 \
 //y=0 //x2=23.31 //y2=2.59
cc_88 ( N_GND_c_7_p N_noxref_6_c_2897_n ) capacitor c=0.0128021f //x=24.05 \
 //y=0 //x2=25.16 //y2=2.08
cc_89 ( N_GND_c_89_p N_noxref_6_c_2898_n ) capacitor c=2.87616e-19 //x=95.83 \
 //y=0 //x2=87.32 //y2=2.08
cc_90 ( N_GND_c_20_p N_noxref_6_c_2898_n ) capacitor c=0.0264258f //x=86.58 \
 //y=0 //x2=87.32 //y2=2.08
cc_91 ( N_GND_c_21_p N_noxref_6_c_2898_n ) capacitor c=2.56782e-19 //x=89.91 \
 //y=0 //x2=87.32 //y2=2.08
cc_92 ( N_GND_c_21_p N_noxref_6_c_2901_n ) capacitor c=0.0156614f //x=89.91 \
 //y=0 //x2=91.02 //y2=2.08
cc_93 ( N_GND_c_22_p N_noxref_6_c_2901_n ) capacitor c=8.26235e-19 //x=93.24 \
 //y=0 //x2=91.02 //y2=2.08
cc_94 ( N_GND_c_94_p N_noxref_6_c_2903_n ) capacitor c=0.00132755f //x=25.04 \
 //y=0 //x2=24.86 //y2=0.875
cc_95 ( N_GND_M15_noxref_d N_noxref_6_c_2903_n ) capacitor c=0.00211996f \
 //x=24.935 //y=0.875 //x2=24.86 //y2=0.875
cc_96 ( N_GND_M15_noxref_d N_noxref_6_c_2905_n ) capacitor c=0.00255985f \
 //x=24.935 //y=0.875 //x2=24.86 //y2=1.22
cc_97 ( N_GND_c_7_p N_noxref_6_c_2906_n ) capacitor c=0.00204716f //x=24.05 \
 //y=0 //x2=24.86 //y2=1.53
cc_98 ( N_GND_c_7_p N_noxref_6_c_2907_n ) capacitor c=0.0110952f //x=24.05 \
 //y=0 //x2=24.86 //y2=1.915
cc_99 ( N_GND_M15_noxref_d N_noxref_6_c_2908_n ) capacitor c=0.0131341f \
 //x=24.935 //y=0.875 //x2=25.235 //y2=0.72
cc_100 ( N_GND_M15_noxref_d N_noxref_6_c_2909_n ) capacitor c=0.00193146f \
 //x=24.935 //y=0.875 //x2=25.235 //y2=1.375
cc_101 ( N_GND_c_101_p N_noxref_6_c_2910_n ) capacitor c=0.00129018f //x=28.69 \
 //y=0 //x2=25.39 //y2=0.875
cc_102 ( N_GND_M15_noxref_d N_noxref_6_c_2910_n ) capacitor c=0.00257848f \
 //x=24.935 //y=0.875 //x2=25.39 //y2=0.875
cc_103 ( N_GND_M15_noxref_d N_noxref_6_c_2912_n ) capacitor c=0.00255985f \
 //x=24.935 //y=0.875 //x2=25.39 //y2=1.22
cc_104 ( N_GND_c_104_p N_noxref_6_c_2913_n ) capacitor c=0.0013864f //x=87.675 \
 //y=0 //x2=87.495 //y2=0.865
cc_105 ( N_GND_M54_noxref_d N_noxref_6_c_2913_n ) capacitor c=0.00220047f \
 //x=87.57 //y=0.865 //x2=87.495 //y2=0.865
cc_106 ( N_GND_M54_noxref_d N_noxref_6_c_2915_n ) capacitor c=0.00255985f \
 //x=87.57 //y=0.865 //x2=87.495 //y2=1.21
cc_107 ( N_GND_c_20_p N_noxref_6_c_2916_n ) capacitor c=0.00189421f //x=86.58 \
 //y=0 //x2=87.495 //y2=1.52
cc_108 ( N_GND_c_20_p N_noxref_6_c_2917_n ) capacitor c=0.00369987f //x=86.58 \
 //y=0 //x2=87.495 //y2=1.915
cc_109 ( N_GND_M54_noxref_d N_noxref_6_c_2918_n ) capacitor c=0.0131326f \
 //x=87.57 //y=0.865 //x2=87.87 //y2=0.71
cc_110 ( N_GND_M54_noxref_d N_noxref_6_c_2919_n ) capacitor c=0.00193127f \
 //x=87.57 //y=0.865 //x2=87.87 //y2=1.365
cc_111 ( N_GND_c_111_p N_noxref_6_c_2920_n ) capacitor c=0.00130622f //x=89.74 \
 //y=0 //x2=88.025 //y2=0.865
cc_112 ( N_GND_M54_noxref_d N_noxref_6_c_2920_n ) capacitor c=0.00257848f \
 //x=87.57 //y=0.865 //x2=88.025 //y2=0.865
cc_113 ( N_GND_M54_noxref_d N_noxref_6_c_2922_n ) capacitor c=0.00255985f \
 //x=87.57 //y=0.865 //x2=88.025 //y2=1.21
cc_114 ( N_GND_c_114_p N_noxref_6_c_2923_n ) capacitor c=0.00135046f \
 //x=91.005 //y=0 //x2=90.825 //y2=0.865
cc_115 ( N_GND_M56_noxref_d N_noxref_6_c_2923_n ) capacitor c=0.00220047f \
 //x=90.9 //y=0.865 //x2=90.825 //y2=0.865
cc_116 ( N_GND_M56_noxref_d N_noxref_6_c_2925_n ) capacitor c=0.00272336f \
 //x=90.9 //y=0.865 //x2=90.825 //y2=1.21
cc_117 ( N_GND_c_21_p N_noxref_6_c_2926_n ) capacitor c=0.00902164f //x=89.91 \
 //y=0 //x2=90.825 //y2=1.915
cc_118 ( N_GND_M56_noxref_d N_noxref_6_c_2927_n ) capacitor c=0.0131326f \
 //x=90.9 //y=0.865 //x2=91.2 //y2=0.71
cc_119 ( N_GND_M56_noxref_d N_noxref_6_c_2928_n ) capacitor c=0.00167494f \
 //x=90.9 //y=0.865 //x2=91.2 //y2=1.365
cc_120 ( N_GND_c_120_p N_noxref_6_c_2929_n ) capacitor c=0.00130622f //x=93.07 \
 //y=0 //x2=91.355 //y2=0.865
cc_121 ( N_GND_M56_noxref_d N_noxref_6_c_2929_n ) capacitor c=0.00257848f \
 //x=90.9 //y=0.865 //x2=91.355 //y2=0.865
cc_122 ( N_GND_M56_noxref_d N_noxref_6_c_2931_n ) capacitor c=0.00272336f \
 //x=90.9 //y=0.865 //x2=91.355 //y2=1.21
cc_123 ( N_GND_c_20_p N_noxref_6_c_2932_n ) capacitor c=0.00917003f //x=86.58 \
 //y=0 //x2=87.32 //y2=2.08
cc_124 ( N_GND_c_7_p N_noxref_6_M14_noxref_d ) capacitor c=0.00591582f \
 //x=24.05 //y=0 //x2=22.635 //y2=0.915
cc_125 ( N_GND_c_4_p N_noxref_7_c_3527_n ) capacitor c=6.0472e-19 //x=9.62 \
 //y=0 //x2=8.14 //y2=2.08
cc_126 ( N_GND_c_5_p N_noxref_7_c_3528_n ) capacitor c=9.24123e-19 //x=14.43 \
 //y=0 //x2=12.95 //y2=2.08
cc_127 ( N_GND_c_6_p N_noxref_7_c_3529_n ) capacitor c=0.0430857f //x=19.24 \
 //y=0 //x2=18.415 //y2=1.665
cc_128 ( N_GND_c_8_p N_noxref_7_c_3530_n ) capacitor c=7.76678e-19 //x=28.86 \
 //y=0 //x2=27.38 //y2=2.08
cc_129 ( N_GND_c_6_p N_noxref_7_M11_noxref_d ) capacitor c=0.00591582f \
 //x=19.24 //y=0 //x2=17.825 //y2=0.915
cc_130 ( N_GND_c_7_p N_noxref_8_c_3866_n ) capacitor c=0.00101012f //x=24.05 \
 //y=0 //x2=22.57 //y2=2.08
cc_131 ( N_GND_c_8_p N_noxref_8_c_3867_n ) capacitor c=0.0432429f //x=28.86 \
 //y=0 //x2=28.035 //y2=1.665
cc_132 ( N_GND_c_8_p N_noxref_8_M17_noxref_d ) capacitor c=0.00591582f \
 //x=28.86 //y=0 //x2=27.445 //y2=0.915
cc_133 ( N_GND_c_9_p N_noxref_9_c_4042_n ) capacitor c=0.0215583f //x=33.67 \
 //y=0 //x2=34.665 //y2=2.59
cc_134 ( N_GND_c_9_p N_noxref_9_c_4043_n ) capacitor c=0.00102529f //x=33.67 \
 //y=0 //x2=33.045 //y2=2.59
cc_135 ( N_GND_c_10_p N_noxref_9_c_4044_n ) capacitor c=0.0230638f //x=38.48 \
 //y=0 //x2=39.475 //y2=2.59
cc_136 ( N_GND_c_9_p N_noxref_9_c_4045_n ) capacitor c=7.16565e-19 //x=33.67 \
 //y=0 //x2=34.895 //y2=2.59
cc_137 ( N_GND_c_9_p N_noxref_9_c_4046_n ) capacitor c=0.04008f //x=33.67 \
 //y=0 //x2=32.845 //y2=1.665
cc_138 ( N_GND_c_9_p N_noxref_9_c_4047_n ) capacitor c=5.56859e-19 //x=33.67 \
 //y=0 //x2=32.93 //y2=2.59
cc_139 ( N_GND_c_9_p N_noxref_9_c_4048_n ) capacitor c=0.0128021f //x=33.67 \
 //y=0 //x2=34.78 //y2=2.08
cc_140 ( N_GND_c_10_p N_noxref_9_c_4049_n ) capacitor c=0.0126655f //x=38.48 \
 //y=0 //x2=39.59 //y2=2.08
cc_141 ( N_GND_c_141_p N_noxref_9_c_4050_n ) capacitor c=0.00132755f //x=34.66 \
 //y=0 //x2=34.48 //y2=0.875
cc_142 ( N_GND_M21_noxref_d N_noxref_9_c_4050_n ) capacitor c=0.00211996f \
 //x=34.555 //y=0.875 //x2=34.48 //y2=0.875
cc_143 ( N_GND_M21_noxref_d N_noxref_9_c_4052_n ) capacitor c=0.00255985f \
 //x=34.555 //y=0.875 //x2=34.48 //y2=1.22
cc_144 ( N_GND_c_9_p N_noxref_9_c_4053_n ) capacitor c=0.00204716f //x=33.67 \
 //y=0 //x2=34.48 //y2=1.53
cc_145 ( N_GND_c_9_p N_noxref_9_c_4054_n ) capacitor c=0.0110952f //x=33.67 \
 //y=0 //x2=34.48 //y2=1.915
cc_146 ( N_GND_M21_noxref_d N_noxref_9_c_4055_n ) capacitor c=0.0131341f \
 //x=34.555 //y=0.875 //x2=34.855 //y2=0.72
cc_147 ( N_GND_M21_noxref_d N_noxref_9_c_4056_n ) capacitor c=0.00193146f \
 //x=34.555 //y=0.875 //x2=34.855 //y2=1.375
cc_148 ( N_GND_c_148_p N_noxref_9_c_4057_n ) capacitor c=0.00129018f //x=38.31 \
 //y=0 //x2=35.01 //y2=0.875
cc_149 ( N_GND_M21_noxref_d N_noxref_9_c_4057_n ) capacitor c=0.00257848f \
 //x=34.555 //y=0.875 //x2=35.01 //y2=0.875
cc_150 ( N_GND_M21_noxref_d N_noxref_9_c_4059_n ) capacitor c=0.00255985f \
 //x=34.555 //y=0.875 //x2=35.01 //y2=1.22
cc_151 ( N_GND_c_151_p N_noxref_9_c_4060_n ) capacitor c=0.00132755f //x=39.47 \
 //y=0 //x2=39.29 //y2=0.875
cc_152 ( N_GND_M24_noxref_d N_noxref_9_c_4060_n ) capacitor c=0.00211996f \
 //x=39.365 //y=0.875 //x2=39.29 //y2=0.875
cc_153 ( N_GND_M24_noxref_d N_noxref_9_c_4062_n ) capacitor c=0.00255985f \
 //x=39.365 //y=0.875 //x2=39.29 //y2=1.22
cc_154 ( N_GND_c_10_p N_noxref_9_c_4063_n ) capacitor c=0.00204716f //x=38.48 \
 //y=0 //x2=39.29 //y2=1.53
cc_155 ( N_GND_c_10_p N_noxref_9_c_4064_n ) capacitor c=0.0112696f //x=38.48 \
 //y=0 //x2=39.29 //y2=1.915
cc_156 ( N_GND_M24_noxref_d N_noxref_9_c_4065_n ) capacitor c=0.0131341f \
 //x=39.365 //y=0.875 //x2=39.665 //y2=0.72
cc_157 ( N_GND_M24_noxref_d N_noxref_9_c_4066_n ) capacitor c=0.00193146f \
 //x=39.365 //y=0.875 //x2=39.665 //y2=1.375
cc_158 ( N_GND_c_158_p N_noxref_9_c_4067_n ) capacitor c=0.00129018f //x=43.12 \
 //y=0 //x2=39.82 //y2=0.875
cc_159 ( N_GND_M24_noxref_d N_noxref_9_c_4067_n ) capacitor c=0.00257848f \
 //x=39.365 //y=0.875 //x2=39.82 //y2=0.875
cc_160 ( N_GND_M24_noxref_d N_noxref_9_c_4069_n ) capacitor c=0.00255985f \
 //x=39.365 //y=0.875 //x2=39.82 //y2=1.22
cc_161 ( N_GND_c_9_p N_noxref_9_M20_noxref_d ) capacitor c=0.00591582f \
 //x=33.67 //y=0 //x2=32.255 //y2=0.915
cc_162 ( N_GND_c_11_p N_noxref_10_c_4295_n ) capacitor c=0.0222748f //x=43.29 \
 //y=0 //x2=44.285 //y2=2.59
cc_163 ( N_GND_c_11_p N_noxref_10_c_4296_n ) capacitor c=0.00102529f //x=43.29 \
 //y=0 //x2=42.665 //y2=2.59
cc_164 ( N_GND_c_11_p N_noxref_10_c_4297_n ) capacitor c=0.0401826f //x=43.29 \
 //y=0 //x2=42.465 //y2=1.665
cc_165 ( N_GND_c_11_p N_noxref_10_c_4298_n ) capacitor c=5.56859e-19 //x=43.29 \
 //y=0 //x2=42.55 //y2=2.59
cc_166 ( N_GND_c_11_p N_noxref_10_c_4299_n ) capacitor c=0.0127664f //x=43.29 \
 //y=0 //x2=44.4 //y2=2.08
cc_167 ( N_GND_c_167_p N_noxref_10_c_4300_n ) capacitor c=0.00132755f \
 //x=44.28 //y=0 //x2=44.1 //y2=0.875
cc_168 ( N_GND_M27_noxref_d N_noxref_10_c_4300_n ) capacitor c=0.00211996f \
 //x=44.175 //y=0.875 //x2=44.1 //y2=0.875
cc_169 ( N_GND_M27_noxref_d N_noxref_10_c_4302_n ) capacitor c=0.00255985f \
 //x=44.175 //y=0.875 //x2=44.1 //y2=1.22
cc_170 ( N_GND_c_11_p N_noxref_10_c_4303_n ) capacitor c=0.00204716f //x=43.29 \
 //y=0 //x2=44.1 //y2=1.53
cc_171 ( N_GND_c_11_p N_noxref_10_c_4304_n ) capacitor c=0.0110952f //x=43.29 \
 //y=0 //x2=44.1 //y2=1.915
cc_172 ( N_GND_M27_noxref_d N_noxref_10_c_4305_n ) capacitor c=0.0131341f \
 //x=44.175 //y=0.875 //x2=44.475 //y2=0.72
cc_173 ( N_GND_M27_noxref_d N_noxref_10_c_4306_n ) capacitor c=0.00193146f \
 //x=44.175 //y=0.875 //x2=44.475 //y2=1.375
cc_174 ( N_GND_c_174_p N_noxref_10_c_4307_n ) capacitor c=0.00129018f \
 //x=47.93 //y=0 //x2=44.63 //y2=0.875
cc_175 ( N_GND_M27_noxref_d N_noxref_10_c_4307_n ) capacitor c=0.00257848f \
 //x=44.175 //y=0.875 //x2=44.63 //y2=0.875
cc_176 ( N_GND_M27_noxref_d N_noxref_10_c_4309_n ) capacitor c=0.00255985f \
 //x=44.175 //y=0.875 //x2=44.63 //y2=1.22
cc_177 ( N_GND_c_11_p N_noxref_10_M26_noxref_d ) capacitor c=0.00591582f \
 //x=43.29 //y=0 //x2=41.875 //y2=0.915
cc_178 ( N_GND_c_9_p N_noxref_11_c_4464_n ) capacitor c=0.00101012f //x=33.67 \
 //y=0 //x2=32.19 //y2=2.08
cc_179 ( N_GND_c_10_p N_noxref_11_c_4465_n ) capacitor c=0.0405987f //x=38.48 \
 //y=0 //x2=37.655 //y2=1.665
cc_180 ( N_GND_c_12_p N_noxref_11_c_4466_n ) capacitor c=0.0153237f //x=48.1 \
 //y=0 //x2=49.21 //y2=2.08
cc_181 ( N_GND_c_181_p N_noxref_11_c_4467_n ) capacitor c=0.00132755f \
 //x=49.09 //y=0 //x2=48.91 //y2=0.875
cc_182 ( N_GND_M30_noxref_d N_noxref_11_c_4467_n ) capacitor c=0.00211996f \
 //x=48.985 //y=0.875 //x2=48.91 //y2=0.875
cc_183 ( N_GND_M30_noxref_d N_noxref_11_c_4469_n ) capacitor c=0.00255985f \
 //x=48.985 //y=0.875 //x2=48.91 //y2=1.22
cc_184 ( N_GND_c_12_p N_noxref_11_c_4470_n ) capacitor c=0.00204716f //x=48.1 \
 //y=0 //x2=48.91 //y2=1.53
cc_185 ( N_GND_c_12_p N_noxref_11_c_4471_n ) capacitor c=0.0110952f //x=48.1 \
 //y=0 //x2=48.91 //y2=1.915
cc_186 ( N_GND_M30_noxref_d N_noxref_11_c_4472_n ) capacitor c=0.0131341f \
 //x=48.985 //y=0.875 //x2=49.285 //y2=0.72
cc_187 ( N_GND_M30_noxref_d N_noxref_11_c_4473_n ) capacitor c=0.00193146f \
 //x=48.985 //y=0.875 //x2=49.285 //y2=1.375
cc_188 ( N_GND_c_188_p N_noxref_11_c_4474_n ) capacitor c=0.00129018f \
 //x=52.74 //y=0 //x2=49.44 //y2=0.875
cc_189 ( N_GND_M30_noxref_d N_noxref_11_c_4474_n ) capacitor c=0.00257848f \
 //x=48.985 //y=0.875 //x2=49.44 //y2=0.875
cc_190 ( N_GND_M30_noxref_d N_noxref_11_c_4476_n ) capacitor c=0.00255985f \
 //x=48.985 //y=0.875 //x2=49.44 //y2=1.22
cc_191 ( N_GND_c_10_p N_noxref_11_M23_noxref_d ) capacitor c=0.00591582f \
 //x=38.48 //y=0 //x2=37.065 //y2=0.915
cc_192 ( N_GND_c_10_p N_noxref_12_c_4745_n ) capacitor c=6.0472e-19 //x=38.48 \
 //y=0 //x2=37 //y2=2.08
cc_193 ( N_GND_c_11_p N_noxref_12_c_4746_n ) capacitor c=9.24123e-19 //x=43.29 \
 //y=0 //x2=41.81 //y2=2.08
cc_194 ( N_GND_c_12_p N_noxref_12_c_4747_n ) capacitor c=0.0430857f //x=48.1 \
 //y=0 //x2=47.275 //y2=1.665
cc_195 ( N_GND_c_14_p N_noxref_12_c_4748_n ) capacitor c=9.84397e-19 //x=57.72 \
 //y=0 //x2=56.24 //y2=2.08
cc_196 ( N_GND_c_12_p N_noxref_12_M29_noxref_d ) capacitor c=0.00591582f \
 //x=48.1 //y=0 //x2=46.685 //y2=0.915
cc_197 ( N_GND_c_13_p N_noxref_13_c_5099_n ) capacitor c=0.0215583f //x=52.91 \
 //y=0 //x2=56.865 //y2=2.59
cc_198 ( N_GND_c_14_p N_noxref_13_c_5099_n ) capacitor c=0.00916039f //x=57.72 \
 //y=0 //x2=56.865 //y2=2.59
cc_199 ( N_GND_c_13_p N_noxref_13_c_5101_n ) capacitor c=6.60802e-19 //x=52.91 \
 //y=0 //x2=51.43 //y2=2.08
cc_200 ( N_GND_c_14_p N_noxref_13_c_5102_n ) capacitor c=0.0404948f //x=57.72 \
 //y=0 //x2=56.895 //y2=1.665
cc_201 ( N_GND_c_14_p N_noxref_13_c_5103_n ) capacitor c=5.56859e-19 //x=57.72 \
 //y=0 //x2=56.98 //y2=2.59
cc_202 ( N_GND_c_14_p N_noxref_13_M35_noxref_d ) capacitor c=0.00591582f \
 //x=57.72 //y=0 //x2=56.305 //y2=0.915
cc_203 ( N_GND_c_89_p N_D_c_5277_n ) capacitor c=0.00600344f //x=95.83 //y=0 \
 //x2=29.855 //y2=4.07
cc_204 ( N_GND_c_89_p N_D_c_5278_n ) capacitor c=0.00234563f //x=95.83 //y=0 \
 //x2=1.225 //y2=4.07
cc_205 ( N_GND_c_1_p N_D_c_5279_n ) capacitor c=0.0178706f //x=0.74 //y=0 \
 //x2=1.11 //y2=2.08
cc_206 ( N_GND_c_8_p N_D_c_5280_n ) capacitor c=0.0156304f //x=28.86 //y=0 \
 //x2=29.97 //y2=2.08
cc_207 ( N_GND_c_14_p N_D_c_5281_n ) capacitor c=0.0152886f //x=57.72 //y=0 \
 //x2=58.83 //y2=2.08
cc_208 ( N_GND_c_208_p N_D_c_5282_n ) capacitor c=0.00132755f //x=0.99 //y=0 \
 //x2=0.81 //y2=0.875
cc_209 ( N_GND_M0_noxref_d N_D_c_5282_n ) capacitor c=0.00211996f //x=0.885 \
 //y=0.875 //x2=0.81 //y2=0.875
cc_210 ( N_GND_M0_noxref_d N_D_c_5284_n ) capacitor c=0.00255985f //x=0.885 \
 //y=0.875 //x2=0.81 //y2=1.22
cc_211 ( N_GND_c_1_p N_D_c_5285_n ) capacitor c=0.00295461f //x=0.74 //y=0 \
 //x2=0.81 //y2=1.53
cc_212 ( N_GND_c_1_p N_D_c_5286_n ) capacitor c=0.0126075f //x=0.74 //y=0 \
 //x2=0.81 //y2=1.915
cc_213 ( N_GND_M0_noxref_d N_D_c_5287_n ) capacitor c=0.0131341f //x=0.885 \
 //y=0.875 //x2=1.185 //y2=0.72
cc_214 ( N_GND_M0_noxref_d N_D_c_5288_n ) capacitor c=0.00193146f //x=0.885 \
 //y=0.875 //x2=1.185 //y2=1.375
cc_215 ( N_GND_c_215_p N_D_c_5289_n ) capacitor c=0.00129018f //x=4.64 //y=0 \
 //x2=1.34 //y2=0.875
cc_216 ( N_GND_M0_noxref_d N_D_c_5289_n ) capacitor c=0.00257848f //x=0.885 \
 //y=0.875 //x2=1.34 //y2=0.875
cc_217 ( N_GND_M0_noxref_d N_D_c_5291_n ) capacitor c=0.00255985f //x=0.885 \
 //y=0.875 //x2=1.34 //y2=1.22
cc_218 ( N_GND_c_218_p N_D_c_5292_n ) capacitor c=0.00132755f //x=29.85 //y=0 \
 //x2=29.67 //y2=0.875
cc_219 ( N_GND_M18_noxref_d N_D_c_5292_n ) capacitor c=0.00211996f //x=29.745 \
 //y=0.875 //x2=29.67 //y2=0.875
cc_220 ( N_GND_M18_noxref_d N_D_c_5294_n ) capacitor c=0.00255985f //x=29.745 \
 //y=0.875 //x2=29.67 //y2=1.22
cc_221 ( N_GND_c_8_p N_D_c_5295_n ) capacitor c=0.00204716f //x=28.86 //y=0 \
 //x2=29.67 //y2=1.53
cc_222 ( N_GND_c_8_p N_D_c_5296_n ) capacitor c=0.0110952f //x=28.86 //y=0 \
 //x2=29.67 //y2=1.915
cc_223 ( N_GND_M18_noxref_d N_D_c_5297_n ) capacitor c=0.0131341f //x=29.745 \
 //y=0.875 //x2=30.045 //y2=0.72
cc_224 ( N_GND_M18_noxref_d N_D_c_5298_n ) capacitor c=0.00193146f //x=29.745 \
 //y=0.875 //x2=30.045 //y2=1.375
cc_225 ( N_GND_c_225_p N_D_c_5299_n ) capacitor c=0.00129018f //x=33.5 //y=0 \
 //x2=30.2 //y2=0.875
cc_226 ( N_GND_M18_noxref_d N_D_c_5299_n ) capacitor c=0.00257848f //x=29.745 \
 //y=0.875 //x2=30.2 //y2=0.875
cc_227 ( N_GND_M18_noxref_d N_D_c_5301_n ) capacitor c=0.00255985f //x=29.745 \
 //y=0.875 //x2=30.2 //y2=1.22
cc_228 ( N_GND_c_228_p N_D_c_5302_n ) capacitor c=0.00132755f //x=58.71 //y=0 \
 //x2=58.53 //y2=0.875
cc_229 ( N_GND_M36_noxref_d N_D_c_5302_n ) capacitor c=0.00211996f //x=58.605 \
 //y=0.875 //x2=58.53 //y2=0.875
cc_230 ( N_GND_M36_noxref_d N_D_c_5304_n ) capacitor c=0.00255985f //x=58.605 \
 //y=0.875 //x2=58.53 //y2=1.22
cc_231 ( N_GND_c_14_p N_D_c_5305_n ) capacitor c=0.00204716f //x=57.72 //y=0 \
 //x2=58.53 //y2=1.53
cc_232 ( N_GND_c_14_p N_D_c_5306_n ) capacitor c=0.0110952f //x=57.72 //y=0 \
 //x2=58.53 //y2=1.915
cc_233 ( N_GND_M36_noxref_d N_D_c_5307_n ) capacitor c=0.0131341f //x=58.605 \
 //y=0.875 //x2=58.905 //y2=0.72
cc_234 ( N_GND_M36_noxref_d N_D_c_5308_n ) capacitor c=0.00193146f //x=58.605 \
 //y=0.875 //x2=58.905 //y2=1.375
cc_235 ( N_GND_c_235_p N_D_c_5309_n ) capacitor c=0.00129018f //x=62.36 //y=0 \
 //x2=59.06 //y2=0.875
cc_236 ( N_GND_M36_noxref_d N_D_c_5309_n ) capacitor c=0.00257848f //x=58.605 \
 //y=0.875 //x2=59.06 //y2=0.875
cc_237 ( N_GND_M36_noxref_d N_D_c_5311_n ) capacitor c=0.00255985f //x=58.605 \
 //y=0.875 //x2=59.06 //y2=1.22
cc_238 ( N_GND_c_15_p N_noxref_15_c_5619_n ) capacitor c=0.0215583f //x=62.53 \
 //y=0 //x2=63.525 //y2=2.59
cc_239 ( N_GND_c_15_p N_noxref_15_c_5620_n ) capacitor c=0.00102529f //x=62.53 \
 //y=0 //x2=61.905 //y2=2.59
cc_240 ( N_GND_c_16_p N_noxref_15_c_5621_n ) capacitor c=0.0230638f //x=67.34 \
 //y=0 //x2=68.335 //y2=2.59
cc_241 ( N_GND_c_15_p N_noxref_15_c_5622_n ) capacitor c=7.16565e-19 //x=62.53 \
 //y=0 //x2=63.755 //y2=2.59
cc_242 ( N_GND_c_15_p N_noxref_15_c_5623_n ) capacitor c=0.04008f //x=62.53 \
 //y=0 //x2=61.705 //y2=1.665
cc_243 ( N_GND_c_15_p N_noxref_15_c_5624_n ) capacitor c=5.56859e-19 //x=62.53 \
 //y=0 //x2=61.79 //y2=2.59
cc_244 ( N_GND_c_15_p N_noxref_15_c_5625_n ) capacitor c=0.0128021f //x=62.53 \
 //y=0 //x2=63.64 //y2=2.08
cc_245 ( N_GND_c_16_p N_noxref_15_c_5626_n ) capacitor c=0.0126655f //x=67.34 \
 //y=0 //x2=68.45 //y2=2.08
cc_246 ( N_GND_c_246_p N_noxref_15_c_5627_n ) capacitor c=0.00132755f \
 //x=63.52 //y=0 //x2=63.34 //y2=0.875
cc_247 ( N_GND_M39_noxref_d N_noxref_15_c_5627_n ) capacitor c=0.00211996f \
 //x=63.415 //y=0.875 //x2=63.34 //y2=0.875
cc_248 ( N_GND_M39_noxref_d N_noxref_15_c_5629_n ) capacitor c=0.00255985f \
 //x=63.415 //y=0.875 //x2=63.34 //y2=1.22
cc_249 ( N_GND_c_15_p N_noxref_15_c_5630_n ) capacitor c=0.00204716f //x=62.53 \
 //y=0 //x2=63.34 //y2=1.53
cc_250 ( N_GND_c_15_p N_noxref_15_c_5631_n ) capacitor c=0.0110952f //x=62.53 \
 //y=0 //x2=63.34 //y2=1.915
cc_251 ( N_GND_M39_noxref_d N_noxref_15_c_5632_n ) capacitor c=0.0131341f \
 //x=63.415 //y=0.875 //x2=63.715 //y2=0.72
cc_252 ( N_GND_M39_noxref_d N_noxref_15_c_5633_n ) capacitor c=0.00193146f \
 //x=63.415 //y=0.875 //x2=63.715 //y2=1.375
cc_253 ( N_GND_c_253_p N_noxref_15_c_5634_n ) capacitor c=0.00129018f \
 //x=67.17 //y=0 //x2=63.87 //y2=0.875
cc_254 ( N_GND_M39_noxref_d N_noxref_15_c_5634_n ) capacitor c=0.00257848f \
 //x=63.415 //y=0.875 //x2=63.87 //y2=0.875
cc_255 ( N_GND_M39_noxref_d N_noxref_15_c_5636_n ) capacitor c=0.00255985f \
 //x=63.415 //y=0.875 //x2=63.87 //y2=1.22
cc_256 ( N_GND_c_256_p N_noxref_15_c_5637_n ) capacitor c=0.00132755f \
 //x=68.33 //y=0 //x2=68.15 //y2=0.875
cc_257 ( N_GND_M42_noxref_d N_noxref_15_c_5637_n ) capacitor c=0.00211996f \
 //x=68.225 //y=0.875 //x2=68.15 //y2=0.875
cc_258 ( N_GND_M42_noxref_d N_noxref_15_c_5639_n ) capacitor c=0.00255985f \
 //x=68.225 //y=0.875 //x2=68.15 //y2=1.22
cc_259 ( N_GND_c_16_p N_noxref_15_c_5640_n ) capacitor c=0.00204716f //x=67.34 \
 //y=0 //x2=68.15 //y2=1.53
cc_260 ( N_GND_c_16_p N_noxref_15_c_5641_n ) capacitor c=0.0112696f //x=67.34 \
 //y=0 //x2=68.15 //y2=1.915
cc_261 ( N_GND_M42_noxref_d N_noxref_15_c_5642_n ) capacitor c=0.0131341f \
 //x=68.225 //y=0.875 //x2=68.525 //y2=0.72
cc_262 ( N_GND_M42_noxref_d N_noxref_15_c_5643_n ) capacitor c=0.00193146f \
 //x=68.225 //y=0.875 //x2=68.525 //y2=1.375
cc_263 ( N_GND_c_263_p N_noxref_15_c_5644_n ) capacitor c=0.00129018f \
 //x=71.98 //y=0 //x2=68.68 //y2=0.875
cc_264 ( N_GND_M42_noxref_d N_noxref_15_c_5644_n ) capacitor c=0.00257848f \
 //x=68.225 //y=0.875 //x2=68.68 //y2=0.875
cc_265 ( N_GND_M42_noxref_d N_noxref_15_c_5646_n ) capacitor c=0.00255985f \
 //x=68.225 //y=0.875 //x2=68.68 //y2=1.22
cc_266 ( N_GND_c_15_p N_noxref_15_M38_noxref_d ) capacitor c=0.00591582f \
 //x=62.53 //y=0 //x2=61.115 //y2=0.915
cc_267 ( N_GND_c_17_p N_noxref_16_c_5872_n ) capacitor c=0.0222748f //x=72.15 \
 //y=0 //x2=73.145 //y2=2.59
cc_268 ( N_GND_c_17_p N_noxref_16_c_5873_n ) capacitor c=0.00102529f //x=72.15 \
 //y=0 //x2=71.525 //y2=2.59
cc_269 ( N_GND_c_17_p N_noxref_16_c_5874_n ) capacitor c=0.0401826f //x=72.15 \
 //y=0 //x2=71.325 //y2=1.665
cc_270 ( N_GND_c_17_p N_noxref_16_c_5875_n ) capacitor c=5.56859e-19 //x=72.15 \
 //y=0 //x2=71.41 //y2=2.59
cc_271 ( N_GND_c_17_p N_noxref_16_c_5876_n ) capacitor c=0.0127664f //x=72.15 \
 //y=0 //x2=73.26 //y2=2.08
cc_272 ( N_GND_c_272_p N_noxref_16_c_5877_n ) capacitor c=0.00132755f \
 //x=73.14 //y=0 //x2=72.96 //y2=0.875
cc_273 ( N_GND_M45_noxref_d N_noxref_16_c_5877_n ) capacitor c=0.00211996f \
 //x=73.035 //y=0.875 //x2=72.96 //y2=0.875
cc_274 ( N_GND_M45_noxref_d N_noxref_16_c_5879_n ) capacitor c=0.00255985f \
 //x=73.035 //y=0.875 //x2=72.96 //y2=1.22
cc_275 ( N_GND_c_17_p N_noxref_16_c_5880_n ) capacitor c=0.00204716f //x=72.15 \
 //y=0 //x2=72.96 //y2=1.53
cc_276 ( N_GND_c_17_p N_noxref_16_c_5881_n ) capacitor c=0.0110952f //x=72.15 \
 //y=0 //x2=72.96 //y2=1.915
cc_277 ( N_GND_M45_noxref_d N_noxref_16_c_5882_n ) capacitor c=0.0131341f \
 //x=73.035 //y=0.875 //x2=73.335 //y2=0.72
cc_278 ( N_GND_M45_noxref_d N_noxref_16_c_5883_n ) capacitor c=0.00193146f \
 //x=73.035 //y=0.875 //x2=73.335 //y2=1.375
cc_279 ( N_GND_c_279_p N_noxref_16_c_5884_n ) capacitor c=0.00129018f \
 //x=76.79 //y=0 //x2=73.49 //y2=0.875
cc_280 ( N_GND_M45_noxref_d N_noxref_16_c_5884_n ) capacitor c=0.00257848f \
 //x=73.035 //y=0.875 //x2=73.49 //y2=0.875
cc_281 ( N_GND_M45_noxref_d N_noxref_16_c_5886_n ) capacitor c=0.00255985f \
 //x=73.035 //y=0.875 //x2=73.49 //y2=1.22
cc_282 ( N_GND_c_17_p N_noxref_16_M44_noxref_d ) capacitor c=0.00591582f \
 //x=72.15 //y=0 //x2=70.735 //y2=0.915
cc_283 ( N_GND_c_3_p N_CLK_c_6040_n ) capacitor c=5.58077e-19 //x=4.81 //y=0 \
 //x2=7.03 //y2=2.08
cc_284 ( N_GND_c_5_p N_CLK_c_6041_n ) capacitor c=7.67786e-19 //x=14.43 //y=0 \
 //x2=16.65 //y2=2.08
cc_285 ( N_GND_c_9_p N_CLK_c_6042_n ) capacitor c=5.58077e-19 //x=33.67 //y=0 \
 //x2=35.89 //y2=2.08
cc_286 ( N_GND_c_11_p N_CLK_c_6043_n ) capacitor c=7.67786e-19 //x=43.29 //y=0 \
 //x2=45.51 //y2=2.08
cc_287 ( N_GND_c_15_p N_CLK_c_6044_n ) capacitor c=5.58077e-19 //x=62.53 //y=0 \
 //x2=64.75 //y2=2.08
cc_288 ( N_GND_c_17_p N_CLK_c_6045_n ) capacitor c=7.67786e-19 //x=72.15 //y=0 \
 //x2=74.37 //y2=2.08
cc_289 ( N_GND_c_15_p N_noxref_18_c_6747_n ) capacitor c=0.00101012f //x=62.53 \
 //y=0 //x2=61.05 //y2=2.08
cc_290 ( N_GND_c_16_p N_noxref_18_c_6748_n ) capacitor c=0.0405987f //x=67.34 \
 //y=0 //x2=66.515 //y2=1.665
cc_291 ( N_GND_c_18_p N_noxref_18_c_6749_n ) capacitor c=0.0153237f //x=76.96 \
 //y=0 //x2=78.07 //y2=2.08
cc_292 ( N_GND_c_292_p N_noxref_18_c_6750_n ) capacitor c=0.00132755f \
 //x=77.95 //y=0 //x2=77.77 //y2=0.875
cc_293 ( N_GND_M48_noxref_d N_noxref_18_c_6750_n ) capacitor c=0.00211996f \
 //x=77.845 //y=0.875 //x2=77.77 //y2=0.875
cc_294 ( N_GND_M48_noxref_d N_noxref_18_c_6752_n ) capacitor c=0.00255985f \
 //x=77.845 //y=0.875 //x2=77.77 //y2=1.22
cc_295 ( N_GND_c_18_p N_noxref_18_c_6753_n ) capacitor c=0.00204716f //x=76.96 \
 //y=0 //x2=77.77 //y2=1.53
cc_296 ( N_GND_c_18_p N_noxref_18_c_6754_n ) capacitor c=0.0110952f //x=76.96 \
 //y=0 //x2=77.77 //y2=1.915
cc_297 ( N_GND_M48_noxref_d N_noxref_18_c_6755_n ) capacitor c=0.0131341f \
 //x=77.845 //y=0.875 //x2=78.145 //y2=0.72
cc_298 ( N_GND_M48_noxref_d N_noxref_18_c_6756_n ) capacitor c=0.00193146f \
 //x=77.845 //y=0.875 //x2=78.145 //y2=1.375
cc_299 ( N_GND_c_299_p N_noxref_18_c_6757_n ) capacitor c=0.00129018f //x=81.6 \
 //y=0 //x2=78.3 //y2=0.875
cc_300 ( N_GND_M48_noxref_d N_noxref_18_c_6757_n ) capacitor c=0.00257848f \
 //x=77.845 //y=0.875 //x2=78.3 //y2=0.875
cc_301 ( N_GND_M48_noxref_d N_noxref_18_c_6759_n ) capacitor c=0.00255985f \
 //x=77.845 //y=0.875 //x2=78.3 //y2=1.22
cc_302 ( N_GND_c_16_p N_noxref_18_M41_noxref_d ) capacitor c=0.00591582f \
 //x=67.34 //y=0 //x2=65.925 //y2=0.915
cc_303 ( N_GND_c_89_p N_RN_c_7021_n ) capacitor c=0.145588f //x=95.83 //y=0 \
 //x2=17.645 //y2=2.22
cc_304 ( N_GND_c_215_p N_RN_c_7021_n ) capacitor c=0.00447829f //x=4.64 //y=0 \
 //x2=17.645 //y2=2.22
cc_305 ( N_GND_c_31_p N_RN_c_7021_n ) capacitor c=0.00274252f //x=5.8 //y=0 \
 //x2=17.645 //y2=2.22
cc_306 ( N_GND_c_38_p N_RN_c_7021_n ) capacitor c=0.00450506f //x=9.45 //y=0 \
 //x2=17.645 //y2=2.22
cc_307 ( N_GND_c_41_p N_RN_c_7021_n ) capacitor c=0.00274252f //x=10.61 //y=0 \
 //x2=17.645 //y2=2.22
cc_308 ( N_GND_c_48_p N_RN_c_7021_n ) capacitor c=0.00450506f //x=14.26 //y=0 \
 //x2=17.645 //y2=2.22
cc_309 ( N_GND_c_57_p N_RN_c_7021_n ) capacitor c=0.00274252f //x=15.42 //y=0 \
 //x2=17.645 //y2=2.22
cc_310 ( N_GND_c_64_p N_RN_c_7021_n ) capacitor c=0.00111309f //x=19.07 //y=0 \
 //x2=17.645 //y2=2.22
cc_311 ( N_GND_c_3_p N_RN_c_7021_n ) capacitor c=0.0379964f //x=4.81 //y=0 \
 //x2=17.645 //y2=2.22
cc_312 ( N_GND_c_4_p N_RN_c_7021_n ) capacitor c=0.0379964f //x=9.62 //y=0 \
 //x2=17.645 //y2=2.22
cc_313 ( N_GND_c_5_p N_RN_c_7021_n ) capacitor c=0.0379964f //x=14.43 //y=0 \
 //x2=17.645 //y2=2.22
cc_314 ( N_GND_c_89_p N_RN_c_7032_n ) capacitor c=0.0019104f //x=95.83 //y=0 \
 //x2=2.335 //y2=2.22
cc_315 ( N_GND_c_89_p N_RN_c_7033_n ) capacitor c=0.0336613f //x=95.83 //y=0 \
 //x2=21.345 //y2=2.22
cc_316 ( N_GND_c_64_p N_RN_c_7033_n ) capacitor c=0.00318526f //x=19.07 //y=0 \
 //x2=21.345 //y2=2.22
cc_317 ( N_GND_c_73_p N_RN_c_7033_n ) capacitor c=0.00274252f //x=20.23 //y=0 \
 //x2=21.345 //y2=2.22
cc_318 ( N_GND_c_6_p N_RN_c_7033_n ) capacitor c=0.0401775f //x=19.24 //y=0 \
 //x2=21.345 //y2=2.22
cc_319 ( N_GND_c_89_p N_RN_c_7037_n ) capacitor c=0.00195247f //x=95.83 //y=0 \
 //x2=17.875 //y2=2.22
cc_320 ( N_GND_c_89_p N_RN_c_7038_n ) capacitor c=0.0897026f //x=95.83 //y=0 \
 //x2=30.965 //y2=2.22
cc_321 ( N_GND_c_80_p N_RN_c_7038_n ) capacitor c=0.00447829f //x=23.88 //y=0 \
 //x2=30.965 //y2=2.22
cc_322 ( N_GND_c_94_p N_RN_c_7038_n ) capacitor c=0.00274252f //x=25.04 //y=0 \
 //x2=30.965 //y2=2.22
cc_323 ( N_GND_c_101_p N_RN_c_7038_n ) capacitor c=0.00450506f //x=28.69 //y=0 \
 //x2=30.965 //y2=2.22
cc_324 ( N_GND_c_218_p N_RN_c_7038_n ) capacitor c=0.00274252f //x=29.85 //y=0 \
 //x2=30.965 //y2=2.22
cc_325 ( N_GND_c_7_p N_RN_c_7038_n ) capacitor c=0.0379964f //x=24.05 //y=0 \
 //x2=30.965 //y2=2.22
cc_326 ( N_GND_c_8_p N_RN_c_7038_n ) capacitor c=0.0401775f //x=28.86 //y=0 \
 //x2=30.965 //y2=2.22
cc_327 ( N_GND_c_89_p N_RN_c_7045_n ) capacitor c=0.00168059f //x=95.83 //y=0 \
 //x2=21.575 //y2=2.22
cc_328 ( N_GND_c_89_p N_RN_c_7046_n ) capacitor c=0.145588f //x=95.83 //y=0 \
 //x2=46.505 //y2=2.22
cc_329 ( N_GND_c_225_p N_RN_c_7046_n ) capacitor c=0.00447829f //x=33.5 //y=0 \
 //x2=46.505 //y2=2.22
cc_330 ( N_GND_c_141_p N_RN_c_7046_n ) capacitor c=0.00274252f //x=34.66 //y=0 \
 //x2=46.505 //y2=2.22
cc_331 ( N_GND_c_148_p N_RN_c_7046_n ) capacitor c=0.00450506f //x=38.31 //y=0 \
 //x2=46.505 //y2=2.22
cc_332 ( N_GND_c_151_p N_RN_c_7046_n ) capacitor c=0.00274252f //x=39.47 //y=0 \
 //x2=46.505 //y2=2.22
cc_333 ( N_GND_c_158_p N_RN_c_7046_n ) capacitor c=0.00450506f //x=43.12 //y=0 \
 //x2=46.505 //y2=2.22
cc_334 ( N_GND_c_167_p N_RN_c_7046_n ) capacitor c=0.00274252f //x=44.28 //y=0 \
 //x2=46.505 //y2=2.22
cc_335 ( N_GND_c_174_p N_RN_c_7046_n ) capacitor c=0.00111309f //x=47.93 //y=0 \
 //x2=46.505 //y2=2.22
cc_336 ( N_GND_c_9_p N_RN_c_7046_n ) capacitor c=0.0379964f //x=33.67 //y=0 \
 //x2=46.505 //y2=2.22
cc_337 ( N_GND_c_10_p N_RN_c_7046_n ) capacitor c=0.0379964f //x=38.48 //y=0 \
 //x2=46.505 //y2=2.22
cc_338 ( N_GND_c_11_p N_RN_c_7046_n ) capacitor c=0.0379964f //x=43.29 //y=0 \
 //x2=46.505 //y2=2.22
cc_339 ( N_GND_c_89_p N_RN_c_7057_n ) capacitor c=0.00168059f //x=95.83 //y=0 \
 //x2=31.195 //y2=2.22
cc_340 ( N_GND_c_89_p N_RN_c_7058_n ) capacitor c=0.0336613f //x=95.83 //y=0 \
 //x2=50.205 //y2=2.22
cc_341 ( N_GND_c_174_p N_RN_c_7058_n ) capacitor c=0.00318526f //x=47.93 //y=0 \
 //x2=50.205 //y2=2.22
cc_342 ( N_GND_c_181_p N_RN_c_7058_n ) capacitor c=0.00274252f //x=49.09 //y=0 \
 //x2=50.205 //y2=2.22
cc_343 ( N_GND_c_12_p N_RN_c_7058_n ) capacitor c=0.0401775f //x=48.1 //y=0 \
 //x2=50.205 //y2=2.22
cc_344 ( N_GND_c_89_p N_RN_c_7062_n ) capacitor c=0.00195247f //x=95.83 //y=0 \
 //x2=46.735 //y2=2.22
cc_345 ( N_GND_c_89_p N_RN_c_7063_n ) capacitor c=0.0897026f //x=95.83 //y=0 \
 //x2=59.825 //y2=2.22
cc_346 ( N_GND_c_188_p N_RN_c_7063_n ) capacitor c=0.00447829f //x=52.74 //y=0 \
 //x2=59.825 //y2=2.22
cc_347 ( N_GND_c_347_p N_RN_c_7063_n ) capacitor c=0.00274252f //x=53.9 //y=0 \
 //x2=59.825 //y2=2.22
cc_348 ( N_GND_c_348_p N_RN_c_7063_n ) capacitor c=0.00450506f //x=57.55 //y=0 \
 //x2=59.825 //y2=2.22
cc_349 ( N_GND_c_228_p N_RN_c_7063_n ) capacitor c=0.00274252f //x=58.71 //y=0 \
 //x2=59.825 //y2=2.22
cc_350 ( N_GND_c_13_p N_RN_c_7063_n ) capacitor c=0.0379964f //x=52.91 //y=0 \
 //x2=59.825 //y2=2.22
cc_351 ( N_GND_c_14_p N_RN_c_7063_n ) capacitor c=0.0401775f //x=57.72 //y=0 \
 //x2=59.825 //y2=2.22
cc_352 ( N_GND_c_89_p N_RN_c_7070_n ) capacitor c=0.00168059f //x=95.83 //y=0 \
 //x2=50.435 //y2=2.22
cc_353 ( N_GND_c_89_p N_RN_c_7071_n ) capacitor c=0.145588f //x=95.83 //y=0 \
 //x2=75.365 //y2=2.22
cc_354 ( N_GND_c_235_p N_RN_c_7071_n ) capacitor c=0.00447829f //x=62.36 //y=0 \
 //x2=75.365 //y2=2.22
cc_355 ( N_GND_c_246_p N_RN_c_7071_n ) capacitor c=0.00274252f //x=63.52 //y=0 \
 //x2=75.365 //y2=2.22
cc_356 ( N_GND_c_253_p N_RN_c_7071_n ) capacitor c=0.00450506f //x=67.17 //y=0 \
 //x2=75.365 //y2=2.22
cc_357 ( N_GND_c_256_p N_RN_c_7071_n ) capacitor c=0.00274252f //x=68.33 //y=0 \
 //x2=75.365 //y2=2.22
cc_358 ( N_GND_c_263_p N_RN_c_7071_n ) capacitor c=0.00450506f //x=71.98 //y=0 \
 //x2=75.365 //y2=2.22
cc_359 ( N_GND_c_272_p N_RN_c_7071_n ) capacitor c=0.00274252f //x=73.14 //y=0 \
 //x2=75.365 //y2=2.22
cc_360 ( N_GND_c_279_p N_RN_c_7071_n ) capacitor c=0.00111309f //x=76.79 //y=0 \
 //x2=75.365 //y2=2.22
cc_361 ( N_GND_c_15_p N_RN_c_7071_n ) capacitor c=0.0379964f //x=62.53 //y=0 \
 //x2=75.365 //y2=2.22
cc_362 ( N_GND_c_16_p N_RN_c_7071_n ) capacitor c=0.0379964f //x=67.34 //y=0 \
 //x2=75.365 //y2=2.22
cc_363 ( N_GND_c_17_p N_RN_c_7071_n ) capacitor c=0.0379964f //x=72.15 //y=0 \
 //x2=75.365 //y2=2.22
cc_364 ( N_GND_c_89_p N_RN_c_7082_n ) capacitor c=0.00168059f //x=95.83 //y=0 \
 //x2=60.055 //y2=2.22
cc_365 ( N_GND_c_89_p N_RN_c_7083_n ) capacitor c=0.0355717f //x=95.83 //y=0 \
 //x2=79.065 //y2=2.22
cc_366 ( N_GND_c_279_p N_RN_c_7083_n ) capacitor c=0.00318526f //x=76.79 //y=0 \
 //x2=79.065 //y2=2.22
cc_367 ( N_GND_c_292_p N_RN_c_7083_n ) capacitor c=0.00274252f //x=77.95 //y=0 \
 //x2=79.065 //y2=2.22
cc_368 ( N_GND_c_18_p N_RN_c_7083_n ) capacitor c=0.0401775f //x=76.96 //y=0 \
 //x2=79.065 //y2=2.22
cc_369 ( N_GND_c_89_p N_RN_c_7087_n ) capacitor c=0.00195247f //x=95.83 //y=0 \
 //x2=75.595 //y2=2.22
cc_370 ( N_GND_c_1_p N_RN_c_7088_n ) capacitor c=8.20622e-19 //x=0.74 //y=0 \
 //x2=2.22 //y2=2.08
cc_371 ( N_GND_c_6_p N_RN_c_7089_n ) capacitor c=8.37259e-19 //x=19.24 //y=0 \
 //x2=17.76 //y2=2.08
cc_372 ( N_GND_c_6_p N_RN_c_7090_n ) capacitor c=5.94159e-19 //x=19.24 //y=0 \
 //x2=21.46 //y2=2.08
cc_373 ( N_GND_c_8_p N_RN_c_7091_n ) capacitor c=5.94159e-19 //x=28.86 //y=0 \
 //x2=31.08 //y2=2.08
cc_374 ( N_GND_c_12_p N_RN_c_7092_n ) capacitor c=8.37259e-19 //x=48.1 //y=0 \
 //x2=46.62 //y2=2.08
cc_375 ( N_GND_c_12_p N_RN_c_7093_n ) capacitor c=8.27581e-19 //x=48.1 //y=0 \
 //x2=50.32 //y2=2.08
cc_376 ( N_GND_c_14_p N_RN_c_7094_n ) capacitor c=7.9303e-19 //x=57.72 //y=0 \
 //x2=59.94 //y2=2.08
cc_377 ( N_GND_c_18_p N_RN_c_7095_n ) capacitor c=8.37259e-19 //x=76.96 //y=0 \
 //x2=75.48 //y2=2.08
cc_378 ( N_GND_c_18_p N_RN_c_7096_n ) capacitor c=8.27581e-19 //x=76.96 //y=0 \
 //x2=79.18 //y2=2.08
cc_379 ( N_GND_c_5_p N_SN_c_8129_n ) capacitor c=0.00750857f //x=14.43 //y=0 \
 //x2=26.155 //y2=2.96
cc_380 ( N_GND_c_6_p N_SN_c_8129_n ) capacitor c=0.00949826f //x=19.24 //y=0 \
 //x2=26.155 //y2=2.96
cc_381 ( N_GND_c_7_p N_SN_c_8129_n ) capacitor c=0.00750857f //x=24.05 //y=0 \
 //x2=26.155 //y2=2.96
cc_382 ( N_GND_c_8_p N_SN_c_8132_n ) capacitor c=0.00949826f //x=28.86 //y=0 \
 //x2=40.585 //y2=2.96
cc_383 ( N_GND_c_9_p N_SN_c_8132_n ) capacitor c=0.00750857f //x=33.67 //y=0 \
 //x2=40.585 //y2=2.96
cc_384 ( N_GND_c_10_p N_SN_c_8132_n ) capacitor c=0.00750857f //x=38.48 //y=0 \
 //x2=40.585 //y2=2.96
cc_385 ( N_GND_c_11_p N_SN_c_8135_n ) capacitor c=0.00750857f //x=43.29 //y=0 \
 //x2=55.015 //y2=2.96
cc_386 ( N_GND_c_12_p N_SN_c_8135_n ) capacitor c=0.00949826f //x=48.1 //y=0 \
 //x2=55.015 //y2=2.96
cc_387 ( N_GND_c_13_p N_SN_c_8135_n ) capacitor c=0.00750857f //x=52.91 //y=0 \
 //x2=55.015 //y2=2.96
cc_388 ( N_GND_c_14_p N_SN_c_8138_n ) capacitor c=0.00949826f //x=57.72 //y=0 \
 //x2=69.445 //y2=2.96
cc_389 ( N_GND_c_15_p N_SN_c_8138_n ) capacitor c=0.00750857f //x=62.53 //y=0 \
 //x2=69.445 //y2=2.96
cc_390 ( N_GND_c_16_p N_SN_c_8138_n ) capacitor c=0.00750857f //x=67.34 //y=0 \
 //x2=69.445 //y2=2.96
cc_391 ( N_GND_c_89_p N_SN_c_8141_n ) capacitor c=0.025494f //x=95.83 //y=0 \
 //x2=83.875 //y2=2.96
cc_392 ( N_GND_c_17_p N_SN_c_8141_n ) capacitor c=0.00750857f //x=72.15 //y=0 \
 //x2=83.875 //y2=2.96
cc_393 ( N_GND_c_18_p N_SN_c_8141_n ) capacitor c=0.00949826f //x=76.96 //y=0 \
 //x2=83.875 //y2=2.96
cc_394 ( N_GND_c_19_p N_SN_c_8141_n ) capacitor c=0.00750857f //x=81.77 //y=0 \
 //x2=83.875 //y2=2.96
cc_395 ( N_GND_c_4_p N_SN_c_8145_n ) capacitor c=7.37634e-19 //x=9.62 //y=0 \
 //x2=11.84 //y2=2.08
cc_396 ( N_GND_c_7_p N_SN_c_8146_n ) capacitor c=7.37634e-19 //x=24.05 //y=0 \
 //x2=26.27 //y2=2.08
cc_397 ( N_GND_c_10_p N_SN_c_8147_n ) capacitor c=7.37634e-19 //x=38.48 //y=0 \
 //x2=40.7 //y2=2.08
cc_398 ( N_GND_c_13_p N_SN_c_8148_n ) capacitor c=4.59642e-19 //x=52.91 //y=0 \
 //x2=55.13 //y2=2.08
cc_399 ( N_GND_c_16_p N_SN_c_8149_n ) capacitor c=7.37634e-19 //x=67.34 //y=0 \
 //x2=69.56 //y2=2.08
cc_400 ( N_GND_c_19_p N_SN_c_8150_n ) capacitor c=5.04543e-19 //x=81.77 //y=0 \
 //x2=83.99 //y2=2.08
cc_401 ( N_GND_c_16_p N_noxref_21_c_8828_n ) capacitor c=6.0472e-19 //x=67.34 \
 //y=0 //x2=65.86 //y2=2.08
cc_402 ( N_GND_c_17_p N_noxref_21_c_8829_n ) capacitor c=9.24123e-19 //x=72.15 \
 //y=0 //x2=70.67 //y2=2.08
cc_403 ( N_GND_c_18_p N_noxref_21_c_8830_n ) capacitor c=0.0430857f //x=76.96 \
 //y=0 //x2=76.135 //y2=1.665
cc_404 ( N_GND_c_20_p N_noxref_21_c_8831_n ) capacitor c=9.84397e-19 //x=86.58 \
 //y=0 //x2=85.1 //y2=2.08
cc_405 ( N_GND_c_18_p N_noxref_21_M47_noxref_d ) capacitor c=0.00591582f \
 //x=76.96 //y=0 //x2=75.545 //y2=0.915
cc_406 ( N_GND_c_89_p N_noxref_22_c_9171_n ) capacitor c=0.0235457f //x=95.83 \
 //y=0 //x2=85.725 //y2=2.59
cc_407 ( N_GND_c_19_p N_noxref_22_c_9171_n ) capacitor c=0.0215583f //x=81.77 \
 //y=0 //x2=85.725 //y2=2.59
cc_408 ( N_GND_c_20_p N_noxref_22_c_9171_n ) capacitor c=0.00916039f //x=86.58 \
 //y=0 //x2=85.725 //y2=2.59
cc_409 ( N_GND_c_89_p N_noxref_22_c_9174_n ) capacitor c=0.00220767f //x=95.83 \
 //y=0 //x2=80.405 //y2=2.59
cc_410 ( N_GND_c_19_p N_noxref_22_c_9175_n ) capacitor c=7.6469e-19 //x=81.77 \
 //y=0 //x2=80.29 //y2=2.08
cc_411 ( N_GND_c_20_p N_noxref_22_c_9176_n ) capacitor c=0.0405953f //x=86.58 \
 //y=0 //x2=85.755 //y2=1.665
cc_412 ( N_GND_c_20_p N_noxref_22_c_9177_n ) capacitor c=5.56859e-19 //x=86.58 \
 //y=0 //x2=85.84 //y2=2.59
cc_413 ( N_GND_c_20_p N_noxref_22_M53_noxref_d ) capacitor c=0.00591203f \
 //x=86.58 //y=0 //x2=85.165 //y2=0.915
cc_414 ( N_GND_c_89_p N_noxref_24_c_9433_n ) capacitor c=0.016597f //x=95.83 \
 //y=0 //x2=82.765 //y2=2.22
cc_415 ( N_GND_c_299_p N_noxref_24_c_9433_n ) capacitor c=0.00296191f //x=81.6 \
 //y=0 //x2=82.765 //y2=2.22
cc_416 ( N_GND_c_416_p N_noxref_24_c_9433_n ) capacitor c=0.00274252f \
 //x=82.76 //y=0 //x2=82.765 //y2=2.22
cc_417 ( N_GND_c_19_p N_noxref_24_c_9433_n ) capacitor c=0.0379964f //x=81.77 \
 //y=0 //x2=82.765 //y2=2.22
cc_418 ( N_GND_c_89_p N_noxref_24_c_9437_n ) capacitor c=0.00266116f //x=95.83 \
 //y=0 //x2=81.145 //y2=2.22
cc_419 ( N_GND_c_299_p N_noxref_24_c_9437_n ) capacitor c=2.28037e-19 //x=81.6 \
 //y=0 //x2=81.145 //y2=2.22
cc_420 ( N_GND_c_19_p N_noxref_24_c_9437_n ) capacitor c=0.00102529f //x=81.77 \
 //y=0 //x2=81.145 //y2=2.22
cc_421 ( N_GND_c_89_p N_noxref_24_c_9440_n ) capacitor c=0.0578533f //x=95.83 \
 //y=0 //x2=92.355 //y2=2.22
cc_422 ( N_GND_c_422_p N_noxref_24_c_9440_n ) capacitor c=0.00450506f \
 //x=86.41 //y=0 //x2=92.355 //y2=2.22
cc_423 ( N_GND_c_104_p N_noxref_24_c_9440_n ) capacitor c=0.00291512f \
 //x=87.675 //y=0 //x2=92.355 //y2=2.22
cc_424 ( N_GND_c_111_p N_noxref_24_c_9440_n ) capacitor c=0.0010086f //x=89.74 \
 //y=0 //x2=92.355 //y2=2.22
cc_425 ( N_GND_c_20_p N_noxref_24_c_9440_n ) capacitor c=0.0426726f //x=86.58 \
 //y=0 //x2=92.355 //y2=2.22
cc_426 ( N_GND_c_21_p N_noxref_24_c_9440_n ) capacitor c=0.0413498f //x=89.91 \
 //y=0 //x2=92.355 //y2=2.22
cc_427 ( N_GND_c_89_p N_noxref_24_c_9446_n ) capacitor c=0.00184466f //x=95.83 \
 //y=0 //x2=82.995 //y2=2.22
cc_428 ( N_GND_c_19_p N_noxref_24_c_9446_n ) capacitor c=8.25398e-19 //x=81.77 \
 //y=0 //x2=82.995 //y2=2.22
cc_429 ( N_GND_c_22_p N_noxref_24_c_9448_n ) capacitor c=0.0396043f //x=93.24 \
 //y=0 //x2=93.865 //y2=2.08
cc_430 ( N_GND_c_22_p N_noxref_24_c_9449_n ) capacitor c=0.00542298f //x=93.24 \
 //y=0 //x2=92.5 //y2=2.08
cc_431 ( N_GND_c_19_p N_noxref_24_c_9450_n ) capacitor c=0.0400254f //x=81.77 \
 //y=0 //x2=80.945 //y2=1.665
cc_432 ( N_GND_c_19_p N_noxref_24_c_9451_n ) capacitor c=5.56859e-19 //x=81.77 \
 //y=0 //x2=81.03 //y2=2.22
cc_433 ( N_GND_c_19_p N_noxref_24_c_9452_n ) capacitor c=0.0127447f //x=81.77 \
 //y=0 //x2=82.88 //y2=2.08
cc_434 ( N_GND_c_21_p N_noxref_24_c_9453_n ) capacitor c=5.16477e-19 //x=89.91 \
 //y=0 //x2=92.5 //y2=2.08
cc_435 ( N_GND_c_22_p N_noxref_24_c_9453_n ) capacitor c=0.0255016f //x=93.24 \
 //y=0 //x2=92.5 //y2=2.08
cc_436 ( N_GND_c_22_p N_noxref_24_c_9455_n ) capacitor c=0.0264827f //x=93.24 \
 //y=0 //x2=93.98 //y2=2.08
cc_437 ( N_GND_c_416_p N_noxref_24_c_9456_n ) capacitor c=0.00132755f \
 //x=82.76 //y=0 //x2=82.58 //y2=0.875
cc_438 ( N_GND_M51_noxref_d N_noxref_24_c_9456_n ) capacitor c=0.00211996f \
 //x=82.655 //y=0.875 //x2=82.58 //y2=0.875
cc_439 ( N_GND_M51_noxref_d N_noxref_24_c_9458_n ) capacitor c=0.00255985f \
 //x=82.655 //y=0.875 //x2=82.58 //y2=1.22
cc_440 ( N_GND_c_19_p N_noxref_24_c_9459_n ) capacitor c=0.00204716f //x=81.77 \
 //y=0 //x2=82.58 //y2=1.53
cc_441 ( N_GND_c_19_p N_noxref_24_c_9460_n ) capacitor c=0.0110952f //x=81.77 \
 //y=0 //x2=82.58 //y2=1.915
cc_442 ( N_GND_M51_noxref_d N_noxref_24_c_9461_n ) capacitor c=0.0131341f \
 //x=82.655 //y=0.875 //x2=82.955 //y2=0.72
cc_443 ( N_GND_M51_noxref_d N_noxref_24_c_9462_n ) capacitor c=0.00193146f \
 //x=82.655 //y=0.875 //x2=82.955 //y2=1.375
cc_444 ( N_GND_c_422_p N_noxref_24_c_9463_n ) capacitor c=0.00129018f \
 //x=86.41 //y=0 //x2=83.11 //y2=0.875
cc_445 ( N_GND_M51_noxref_d N_noxref_24_c_9463_n ) capacitor c=0.00257848f \
 //x=82.655 //y=0.875 //x2=83.11 //y2=0.875
cc_446 ( N_GND_M51_noxref_d N_noxref_24_c_9465_n ) capacitor c=0.00255985f \
 //x=82.655 //y=0.875 //x2=83.11 //y2=1.22
cc_447 ( N_GND_c_22_p N_noxref_24_c_9466_n ) capacitor c=0.0103285f //x=93.24 \
 //y=0 //x2=92.325 //y2=1.915
cc_448 ( N_GND_c_448_p N_noxref_24_c_9467_n ) capacitor c=0.0013864f \
 //x=94.335 //y=0 //x2=94.155 //y2=0.865
cc_449 ( N_GND_M58_noxref_d N_noxref_24_c_9467_n ) capacitor c=0.00220047f \
 //x=94.23 //y=0.865 //x2=94.155 //y2=0.865
cc_450 ( N_GND_M58_noxref_d N_noxref_24_c_9469_n ) capacitor c=0.00272336f \
 //x=94.23 //y=0.865 //x2=94.155 //y2=1.21
cc_451 ( N_GND_c_22_p N_noxref_24_c_9470_n ) capacitor c=0.00369763f //x=93.24 \
 //y=0 //x2=94.155 //y2=1.915
cc_452 ( N_GND_M58_noxref_d N_noxref_24_c_9471_n ) capacitor c=0.0131326f \
 //x=94.23 //y=0.865 //x2=94.53 //y2=0.71
cc_453 ( N_GND_M58_noxref_d N_noxref_24_c_9472_n ) capacitor c=0.00167494f \
 //x=94.23 //y=0.865 //x2=94.53 //y2=1.365
cc_454 ( N_GND_c_2_p N_noxref_24_c_9473_n ) capacitor c=0.00130622f //x=95.83 \
 //y=0 //x2=94.685 //y2=0.865
cc_455 ( N_GND_M58_noxref_d N_noxref_24_c_9473_n ) capacitor c=0.00257848f \
 //x=94.23 //y=0.865 //x2=94.685 //y2=0.865
cc_456 ( N_GND_M58_noxref_d N_noxref_24_c_9475_n ) capacitor c=0.00272336f \
 //x=94.23 //y=0.865 //x2=94.685 //y2=1.21
cc_457 ( N_GND_c_22_p N_noxref_24_c_9476_n ) capacitor c=0.00662863f //x=93.24 \
 //y=0 //x2=93.98 //y2=2.08
cc_458 ( N_GND_c_19_p N_noxref_24_M50_noxref_d ) capacitor c=0.00591582f \
 //x=81.77 //y=0 //x2=80.355 //y2=0.915
cc_459 ( N_GND_c_20_p N_noxref_26_c_9912_n ) capacitor c=0.00273037f //x=86.58 \
 //y=0 //x2=88.315 //y2=4.07
cc_460 ( N_GND_c_21_p N_noxref_26_c_9913_n ) capacitor c=0.00273037f //x=89.91 \
 //y=0 //x2=94.975 //y2=4.07
cc_461 ( N_GND_c_22_p N_noxref_26_c_9913_n ) capacitor c=0.00281233f //x=93.24 \
 //y=0 //x2=94.975 //y2=4.07
cc_462 ( N_GND_c_13_p N_noxref_26_c_9915_n ) capacitor c=0.0404651f //x=52.91 \
 //y=0 //x2=52.085 //y2=1.665
cc_463 ( N_GND_c_13_p N_noxref_26_c_9916_n ) capacitor c=0.0130159f //x=52.91 \
 //y=0 //x2=54.02 //y2=2.08
cc_464 ( N_GND_c_20_p N_noxref_26_c_9917_n ) capacitor c=0.00112925f //x=86.58 \
 //y=0 //x2=88.43 //y2=2.08
cc_465 ( N_GND_c_21_p N_noxref_26_c_9917_n ) capacitor c=0.0105756f //x=89.91 \
 //y=0 //x2=88.43 //y2=2.08
cc_466 ( N_GND_c_2_p N_noxref_26_c_9919_n ) capacitor c=0.00128267f //x=95.83 \
 //y=0 //x2=95.09 //y2=2.08
cc_467 ( N_GND_c_22_p N_noxref_26_c_9919_n ) capacitor c=9.01984e-19 //x=93.24 \
 //y=0 //x2=95.09 //y2=2.08
cc_468 ( N_GND_c_347_p N_noxref_26_c_9921_n ) capacitor c=0.00132755f //x=53.9 \
 //y=0 //x2=53.72 //y2=0.875
cc_469 ( N_GND_M33_noxref_d N_noxref_26_c_9921_n ) capacitor c=0.00211996f \
 //x=53.795 //y=0.875 //x2=53.72 //y2=0.875
cc_470 ( N_GND_M33_noxref_d N_noxref_26_c_9923_n ) capacitor c=0.00255985f \
 //x=53.795 //y=0.875 //x2=53.72 //y2=1.22
cc_471 ( N_GND_c_13_p N_noxref_26_c_9924_n ) capacitor c=0.00204716f //x=52.91 \
 //y=0 //x2=53.72 //y2=1.53
cc_472 ( N_GND_c_13_p N_noxref_26_c_9925_n ) capacitor c=0.0110952f //x=52.91 \
 //y=0 //x2=53.72 //y2=1.915
cc_473 ( N_GND_M33_noxref_d N_noxref_26_c_9926_n ) capacitor c=0.0131341f \
 //x=53.795 //y=0.875 //x2=54.095 //y2=0.72
cc_474 ( N_GND_M33_noxref_d N_noxref_26_c_9927_n ) capacitor c=0.00193146f \
 //x=53.795 //y=0.875 //x2=54.095 //y2=1.375
cc_475 ( N_GND_c_348_p N_noxref_26_c_9928_n ) capacitor c=0.00129018f \
 //x=57.55 //y=0 //x2=54.25 //y2=0.875
cc_476 ( N_GND_M33_noxref_d N_noxref_26_c_9928_n ) capacitor c=0.00257848f \
 //x=53.795 //y=0.875 //x2=54.25 //y2=0.875
cc_477 ( N_GND_M33_noxref_d N_noxref_26_c_9930_n ) capacitor c=0.00255985f \
 //x=53.795 //y=0.875 //x2=54.25 //y2=1.22
cc_478 ( N_GND_c_21_p N_noxref_26_c_9931_n ) capacitor c=2.63786e-19 //x=89.91 \
 //y=0 //x2=88.43 //y2=2.08
cc_479 ( N_GND_c_13_p N_noxref_26_M32_noxref_d ) capacitor c=0.00591582f \
 //x=52.91 //y=0 //x2=51.495 //y2=0.915
cc_480 ( N_GND_c_89_p Q ) capacitor c=0.00233821f //x=95.83 //y=0 //x2=95.83 \
 //y2=4.07
cc_481 ( N_GND_c_89_p N_Q_c_10368_n ) capacitor c=0.0695894f //x=95.83 //y=0 \
 //x2=91.945 //y2=1.18
cc_482 ( N_GND_c_111_p N_Q_c_10368_n ) capacitor c=0.0081414f //x=89.74 //y=0 \
 //x2=91.945 //y2=1.18
cc_483 ( N_GND_c_114_p N_Q_c_10368_n ) capacitor c=0.0101988f //x=91.005 //y=0 \
 //x2=91.945 //y2=1.18
cc_484 ( N_GND_c_120_p N_Q_c_10368_n ) capacitor c=0.00469062f //x=93.07 //y=0 \
 //x2=91.945 //y2=1.18
cc_485 ( N_GND_c_2_p N_Q_c_10368_n ) capacitor c=0.00131115f //x=95.83 //y=0 \
 //x2=91.945 //y2=1.18
cc_486 ( N_GND_c_21_p N_Q_c_10368_n ) capacitor c=0.039515f //x=89.91 //y=0 \
 //x2=91.945 //y2=1.18
cc_487 ( N_GND_M56_noxref_d N_Q_c_10368_n ) capacitor c=0.00960943f //x=90.9 \
 //y=0.865 //x2=91.945 //y2=1.18
cc_488 ( N_GND_c_89_p N_Q_c_10375_n ) capacitor c=0.00715563f //x=95.83 //y=0 \
 //x2=88.845 //y2=1.18
cc_489 ( N_GND_c_89_p N_Q_c_10376_n ) capacitor c=0.0769193f //x=95.83 //y=0 \
 //x2=95.275 //y2=1.18
cc_490 ( N_GND_c_120_p N_Q_c_10376_n ) capacitor c=0.00788597f //x=93.07 //y=0 \
 //x2=95.275 //y2=1.18
cc_491 ( N_GND_c_448_p N_Q_c_10376_n ) capacitor c=0.00974891f //x=94.335 \
 //y=0 //x2=95.275 //y2=1.18
cc_492 ( N_GND_c_2_p N_Q_c_10376_n ) capacitor c=0.00577123f //x=95.83 //y=0 \
 //x2=95.275 //y2=1.18
cc_493 ( N_GND_c_22_p N_Q_c_10376_n ) capacitor c=0.0384312f //x=93.24 //y=0 \
 //x2=95.275 //y2=1.18
cc_494 ( N_GND_M58_noxref_d N_Q_c_10376_n ) capacitor c=0.00960943f //x=94.23 \
 //y=0.865 //x2=95.275 //y2=1.18
cc_495 ( N_GND_c_89_p N_Q_c_10382_n ) capacitor c=0.00664346f //x=95.83 //y=0 \
 //x2=92.175 //y2=1.18
cc_496 ( N_GND_c_2_p N_Q_c_10383_n ) capacitor c=0.04686f //x=95.83 //y=0 \
 //x2=95.745 //y2=1.645
cc_497 ( N_GND_c_22_p N_Q_c_10384_n ) capacitor c=0.00109945f //x=93.24 //y=0 \
 //x2=95.83 //y2=4.07
cc_498 ( N_GND_c_89_p N_Q_M55_noxref_d ) capacitor c=2.00936e-19 //x=95.83 \
 //y=0 //x2=88.54 //y2=0.905
cc_499 ( N_GND_c_21_p N_Q_M55_noxref_d ) capacitor c=0.00141366f //x=89.91 \
 //y=0 //x2=88.54 //y2=0.905
cc_500 ( N_GND_M54_noxref_d N_Q_M55_noxref_d ) capacitor c=0.00128667f \
 //x=87.57 //y=0.865 //x2=88.54 //y2=0.905
cc_501 ( N_GND_c_89_p N_Q_M57_noxref_d ) capacitor c=2.00936e-19 //x=95.83 \
 //y=0 //x2=91.87 //y2=0.905
cc_502 ( N_GND_c_22_p N_Q_M57_noxref_d ) capacitor c=0.0014176f //x=93.24 \
 //y=0 //x2=91.87 //y2=0.905
cc_503 ( N_GND_M56_noxref_d N_Q_M57_noxref_d ) capacitor c=0.0012247f //x=90.9 \
 //y=0.865 //x2=91.87 //y2=0.905
cc_504 ( N_GND_c_89_p N_Q_M59_noxref_d ) capacitor c=2.00936e-19 //x=95.83 \
 //y=0 //x2=95.2 //y2=0.905
cc_505 ( N_GND_c_2_p N_Q_M59_noxref_d ) capacitor c=0.00524992f //x=95.83 \
 //y=0 //x2=95.2 //y2=0.905
cc_506 ( N_GND_c_22_p N_Q_M59_noxref_d ) capacitor c=8.62423e-19 //x=93.24 \
 //y=0 //x2=95.2 //y2=0.905
cc_507 ( N_GND_M58_noxref_d N_Q_M59_noxref_d ) capacitor c=0.0012247f \
 //x=94.23 //y=0.865 //x2=95.2 //y2=0.905
cc_508 ( N_GND_c_89_p N_noxref_28_c_10542_n ) capacitor c=0.0059534f //x=95.83 \
 //y=0 //x2=1.475 //y2=1.59
cc_509 ( N_GND_c_208_p N_noxref_28_c_10542_n ) capacitor c=0.00110021f \
 //x=0.99 //y=0 //x2=1.475 //y2=1.59
cc_510 ( N_GND_c_215_p N_noxref_28_c_10542_n ) capacitor c=0.00179185f \
 //x=4.64 //y=0 //x2=1.475 //y2=1.59
cc_511 ( N_GND_M0_noxref_d N_noxref_28_c_10542_n ) capacitor c=0.00894788f \
 //x=0.885 //y=0.875 //x2=1.475 //y2=1.59
cc_512 ( N_GND_c_89_p N_noxref_28_c_10546_n ) capacitor c=0.00575184f \
 //x=95.83 //y=0 //x2=1.56 //y2=0.625
cc_513 ( N_GND_c_215_p N_noxref_28_c_10546_n ) capacitor c=0.0140218f //x=4.64 \
 //y=0 //x2=1.56 //y2=0.625
cc_514 ( N_GND_M0_noxref_d N_noxref_28_c_10546_n ) capacitor c=0.033954f \
 //x=0.885 //y=0.875 //x2=1.56 //y2=0.625
cc_515 ( N_GND_c_89_p N_noxref_28_c_10549_n ) capacitor c=0.0122695f //x=95.83 \
 //y=0 //x2=2.445 //y2=0.54
cc_516 ( N_GND_c_215_p N_noxref_28_c_10549_n ) capacitor c=0.0358309f //x=4.64 \
 //y=0 //x2=2.445 //y2=0.54
cc_517 ( N_GND_c_89_p N_noxref_28_M0_noxref_s ) capacitor c=0.00962687f \
 //x=95.83 //y=0 //x2=0.455 //y2=0.375
cc_518 ( N_GND_c_208_p N_noxref_28_M0_noxref_s ) capacitor c=0.0140218f \
 //x=0.99 //y=0 //x2=0.455 //y2=0.375
cc_519 ( N_GND_c_1_p N_noxref_28_M0_noxref_s ) capacitor c=0.0712607f //x=0.74 \
 //y=0 //x2=0.455 //y2=0.375
cc_520 ( N_GND_c_215_p N_noxref_28_M0_noxref_s ) capacitor c=0.0131437f \
 //x=4.64 //y=0 //x2=0.455 //y2=0.375
cc_521 ( N_GND_c_3_p N_noxref_28_M0_noxref_s ) capacitor c=3.31601e-19 \
 //x=4.81 //y=0 //x2=0.455 //y2=0.375
cc_522 ( N_GND_M0_noxref_d N_noxref_28_M0_noxref_s ) capacitor c=0.033718f \
 //x=0.885 //y=0.875 //x2=0.455 //y2=0.375
cc_523 ( N_GND_c_89_p N_noxref_29_c_10591_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=3.015 //y2=0.995
cc_524 ( N_GND_c_215_p N_noxref_29_c_10591_n ) capacitor c=0.00934524f \
 //x=4.64 //y=0 //x2=3.015 //y2=0.995
cc_525 ( N_GND_c_89_p N_noxref_29_c_10593_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=3.1 //y2=0.625
cc_526 ( N_GND_c_215_p N_noxref_29_c_10593_n ) capacitor c=0.0140928f //x=4.64 \
 //y=0 //x2=3.1 //y2=0.625
cc_527 ( N_GND_M0_noxref_d N_noxref_29_c_10593_n ) capacitor c=6.21394e-19 \
 //x=0.885 //y=0.875 //x2=3.1 //y2=0.625
cc_528 ( N_GND_c_89_p N_noxref_29_c_10596_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=3.985 //y2=0.54
cc_529 ( N_GND_c_215_p N_noxref_29_c_10596_n ) capacitor c=0.0363691f //x=4.64 \
 //y=0 //x2=3.985 //y2=0.54
cc_530 ( N_GND_c_89_p N_noxref_29_c_10598_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=4.07 //y2=0.625
cc_531 ( N_GND_c_215_p N_noxref_29_c_10598_n ) capacitor c=0.0140304f //x=4.64 \
 //y=0 //x2=4.07 //y2=0.625
cc_532 ( N_GND_c_3_p N_noxref_29_c_10598_n ) capacitor c=0.0404137f //x=4.81 \
 //y=0 //x2=4.07 //y2=0.625
cc_533 ( N_GND_M0_noxref_d N_noxref_29_M1_noxref_d ) capacitor c=0.00162435f \
 //x=0.885 //y=0.875 //x2=1.86 //y2=0.91
cc_534 ( N_GND_c_1_p N_noxref_29_M2_noxref_s ) capacitor c=8.16352e-19 \
 //x=0.74 //y=0 //x2=2.965 //y2=0.375
cc_535 ( N_GND_c_3_p N_noxref_29_M2_noxref_s ) capacitor c=0.00183204f \
 //x=4.81 //y=0 //x2=2.965 //y2=0.375
cc_536 ( N_GND_c_89_p N_noxref_30_c_10643_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=6.285 //y2=1.59
cc_537 ( N_GND_c_31_p N_noxref_30_c_10643_n ) capacitor c=0.00111448f //x=5.8 \
 //y=0 //x2=6.285 //y2=1.59
cc_538 ( N_GND_c_38_p N_noxref_30_c_10643_n ) capacitor c=0.00180612f //x=9.45 \
 //y=0 //x2=6.285 //y2=1.59
cc_539 ( N_GND_M3_noxref_d N_noxref_30_c_10643_n ) capacitor c=0.00853078f \
 //x=5.695 //y=0.875 //x2=6.285 //y2=1.59
cc_540 ( N_GND_c_89_p N_noxref_30_c_10647_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=6.37 //y2=0.625
cc_541 ( N_GND_c_38_p N_noxref_30_c_10647_n ) capacitor c=0.0140928f //x=9.45 \
 //y=0 //x2=6.37 //y2=0.625
cc_542 ( N_GND_M3_noxref_d N_noxref_30_c_10647_n ) capacitor c=0.033954f \
 //x=5.695 //y=0.875 //x2=6.37 //y2=0.625
cc_543 ( N_GND_c_89_p N_noxref_30_c_10650_n ) capacitor c=0.0104506f //x=95.83 \
 //y=0 //x2=7.255 //y2=0.54
cc_544 ( N_GND_c_38_p N_noxref_30_c_10650_n ) capacitor c=0.0360726f //x=9.45 \
 //y=0 //x2=7.255 //y2=0.54
cc_545 ( N_GND_c_89_p N_noxref_30_M3_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=5.265 //y2=0.375
cc_546 ( N_GND_c_31_p N_noxref_30_M3_noxref_s ) capacitor c=0.0140928f //x=5.8 \
 //y=0 //x2=5.265 //y2=0.375
cc_547 ( N_GND_c_38_p N_noxref_30_M3_noxref_s ) capacitor c=0.0136651f \
 //x=9.45 //y=0 //x2=5.265 //y2=0.375
cc_548 ( N_GND_c_3_p N_noxref_30_M3_noxref_s ) capacitor c=0.0696963f //x=4.81 \
 //y=0 //x2=5.265 //y2=0.375
cc_549 ( N_GND_c_4_p N_noxref_30_M3_noxref_s ) capacitor c=3.31601e-19 \
 //x=9.62 //y=0 //x2=5.265 //y2=0.375
cc_550 ( N_GND_M3_noxref_d N_noxref_30_M3_noxref_s ) capacitor c=0.033718f \
 //x=5.695 //y=0.875 //x2=5.265 //y2=0.375
cc_551 ( N_GND_c_89_p N_noxref_31_c_10692_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=7.825 //y2=0.995
cc_552 ( N_GND_c_38_p N_noxref_31_c_10692_n ) capacitor c=0.00934524f //x=9.45 \
 //y=0 //x2=7.825 //y2=0.995
cc_553 ( N_GND_c_89_p N_noxref_31_c_10694_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=7.91 //y2=0.625
cc_554 ( N_GND_c_38_p N_noxref_31_c_10694_n ) capacitor c=0.0140928f //x=9.45 \
 //y=0 //x2=7.91 //y2=0.625
cc_555 ( N_GND_M3_noxref_d N_noxref_31_c_10694_n ) capacitor c=6.21394e-19 \
 //x=5.695 //y=0.875 //x2=7.91 //y2=0.625
cc_556 ( N_GND_c_89_p N_noxref_31_c_10697_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=8.795 //y2=0.54
cc_557 ( N_GND_c_38_p N_noxref_31_c_10697_n ) capacitor c=0.0364215f //x=9.45 \
 //y=0 //x2=8.795 //y2=0.54
cc_558 ( N_GND_c_89_p N_noxref_31_c_10699_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=8.88 //y2=0.625
cc_559 ( N_GND_c_38_p N_noxref_31_c_10699_n ) capacitor c=0.0140304f //x=9.45 \
 //y=0 //x2=8.88 //y2=0.625
cc_560 ( N_GND_c_4_p N_noxref_31_c_10699_n ) capacitor c=0.0404137f //x=9.62 \
 //y=0 //x2=8.88 //y2=0.625
cc_561 ( N_GND_M3_noxref_d N_noxref_31_M4_noxref_d ) capacitor c=0.00162435f \
 //x=5.695 //y=0.875 //x2=6.67 //y2=0.91
cc_562 ( N_GND_c_3_p N_noxref_31_M5_noxref_s ) capacitor c=8.16352e-19 \
 //x=4.81 //y=0 //x2=7.775 //y2=0.375
cc_563 ( N_GND_c_4_p N_noxref_31_M5_noxref_s ) capacitor c=0.00183204f \
 //x=9.62 //y=0 //x2=7.775 //y2=0.375
cc_564 ( N_GND_c_89_p N_noxref_32_c_10744_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=11.095 //y2=1.59
cc_565 ( N_GND_c_41_p N_noxref_32_c_10744_n ) capacitor c=0.00111448f \
 //x=10.61 //y=0 //x2=11.095 //y2=1.59
cc_566 ( N_GND_c_48_p N_noxref_32_c_10744_n ) capacitor c=0.00180612f \
 //x=14.26 //y=0 //x2=11.095 //y2=1.59
cc_567 ( N_GND_M6_noxref_d N_noxref_32_c_10744_n ) capacitor c=0.00853078f \
 //x=10.505 //y=0.875 //x2=11.095 //y2=1.59
cc_568 ( N_GND_c_89_p N_noxref_32_c_10748_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=11.18 //y2=0.625
cc_569 ( N_GND_c_48_p N_noxref_32_c_10748_n ) capacitor c=0.0140928f //x=14.26 \
 //y=0 //x2=11.18 //y2=0.625
cc_570 ( N_GND_M6_noxref_d N_noxref_32_c_10748_n ) capacitor c=0.033954f \
 //x=10.505 //y=0.875 //x2=11.18 //y2=0.625
cc_571 ( N_GND_c_89_p N_noxref_32_c_10751_n ) capacitor c=0.0104506f //x=95.83 \
 //y=0 //x2=12.065 //y2=0.54
cc_572 ( N_GND_c_48_p N_noxref_32_c_10751_n ) capacitor c=0.0360726f //x=14.26 \
 //y=0 //x2=12.065 //y2=0.54
cc_573 ( N_GND_c_89_p N_noxref_32_M6_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=10.075 //y2=0.375
cc_574 ( N_GND_c_41_p N_noxref_32_M6_noxref_s ) capacitor c=0.0140928f \
 //x=10.61 //y=0 //x2=10.075 //y2=0.375
cc_575 ( N_GND_c_48_p N_noxref_32_M6_noxref_s ) capacitor c=0.0131437f \
 //x=14.26 //y=0 //x2=10.075 //y2=0.375
cc_576 ( N_GND_c_4_p N_noxref_32_M6_noxref_s ) capacitor c=0.0696963f //x=9.62 \
 //y=0 //x2=10.075 //y2=0.375
cc_577 ( N_GND_c_5_p N_noxref_32_M6_noxref_s ) capacitor c=3.31601e-19 \
 //x=14.43 //y=0 //x2=10.075 //y2=0.375
cc_578 ( N_GND_M6_noxref_d N_noxref_32_M6_noxref_s ) capacitor c=0.033718f \
 //x=10.505 //y=0.875 //x2=10.075 //y2=0.375
cc_579 ( N_GND_c_89_p N_noxref_33_c_10793_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=12.635 //y2=0.995
cc_580 ( N_GND_c_48_p N_noxref_33_c_10793_n ) capacitor c=0.00934524f \
 //x=14.26 //y=0 //x2=12.635 //y2=0.995
cc_581 ( N_GND_c_89_p N_noxref_33_c_10795_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=12.72 //y2=0.625
cc_582 ( N_GND_c_48_p N_noxref_33_c_10795_n ) capacitor c=0.0140928f //x=14.26 \
 //y=0 //x2=12.72 //y2=0.625
cc_583 ( N_GND_M6_noxref_d N_noxref_33_c_10795_n ) capacitor c=6.21394e-19 \
 //x=10.505 //y=0.875 //x2=12.72 //y2=0.625
cc_584 ( N_GND_c_89_p N_noxref_33_c_10798_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=13.605 //y2=0.54
cc_585 ( N_GND_c_48_p N_noxref_33_c_10798_n ) capacitor c=0.0364215f //x=14.26 \
 //y=0 //x2=13.605 //y2=0.54
cc_586 ( N_GND_c_89_p N_noxref_33_c_10800_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=13.69 //y2=0.625
cc_587 ( N_GND_c_48_p N_noxref_33_c_10800_n ) capacitor c=0.0140304f //x=14.26 \
 //y=0 //x2=13.69 //y2=0.625
cc_588 ( N_GND_c_5_p N_noxref_33_c_10800_n ) capacitor c=0.0404137f //x=14.43 \
 //y=0 //x2=13.69 //y2=0.625
cc_589 ( N_GND_M6_noxref_d N_noxref_33_M7_noxref_d ) capacitor c=0.00162435f \
 //x=10.505 //y=0.875 //x2=11.48 //y2=0.91
cc_590 ( N_GND_c_4_p N_noxref_33_M8_noxref_s ) capacitor c=8.16352e-19 \
 //x=9.62 //y=0 //x2=12.585 //y2=0.375
cc_591 ( N_GND_c_5_p N_noxref_33_M8_noxref_s ) capacitor c=0.00183204f \
 //x=14.43 //y=0 //x2=12.585 //y2=0.375
cc_592 ( N_GND_c_89_p N_noxref_34_c_10845_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=15.905 //y2=1.59
cc_593 ( N_GND_c_57_p N_noxref_34_c_10845_n ) capacitor c=0.00111448f \
 //x=15.42 //y=0 //x2=15.905 //y2=1.59
cc_594 ( N_GND_c_64_p N_noxref_34_c_10845_n ) capacitor c=0.00180612f \
 //x=19.07 //y=0 //x2=15.905 //y2=1.59
cc_595 ( N_GND_M9_noxref_d N_noxref_34_c_10845_n ) capacitor c=0.00853078f \
 //x=15.315 //y=0.875 //x2=15.905 //y2=1.59
cc_596 ( N_GND_c_89_p N_noxref_34_c_10849_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=15.99 //y2=0.625
cc_597 ( N_GND_c_64_p N_noxref_34_c_10849_n ) capacitor c=0.0140928f //x=19.07 \
 //y=0 //x2=15.99 //y2=0.625
cc_598 ( N_GND_M9_noxref_d N_noxref_34_c_10849_n ) capacitor c=0.033954f \
 //x=15.315 //y=0.875 //x2=15.99 //y2=0.625
cc_599 ( N_GND_c_89_p N_noxref_34_c_10852_n ) capacitor c=0.0104506f //x=95.83 \
 //y=0 //x2=16.875 //y2=0.54
cc_600 ( N_GND_c_64_p N_noxref_34_c_10852_n ) capacitor c=0.0360726f //x=19.07 \
 //y=0 //x2=16.875 //y2=0.54
cc_601 ( N_GND_c_89_p N_noxref_34_M9_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=14.885 //y2=0.375
cc_602 ( N_GND_c_57_p N_noxref_34_M9_noxref_s ) capacitor c=0.0140928f \
 //x=15.42 //y=0 //x2=14.885 //y2=0.375
cc_603 ( N_GND_c_64_p N_noxref_34_M9_noxref_s ) capacitor c=0.0131437f \
 //x=19.07 //y=0 //x2=14.885 //y2=0.375
cc_604 ( N_GND_c_5_p N_noxref_34_M9_noxref_s ) capacitor c=0.0696963f \
 //x=14.43 //y=0 //x2=14.885 //y2=0.375
cc_605 ( N_GND_c_6_p N_noxref_34_M9_noxref_s ) capacitor c=3.31601e-19 \
 //x=19.24 //y=0 //x2=14.885 //y2=0.375
cc_606 ( N_GND_M9_noxref_d N_noxref_34_M9_noxref_s ) capacitor c=0.033718f \
 //x=15.315 //y=0.875 //x2=14.885 //y2=0.375
cc_607 ( N_GND_c_89_p N_noxref_35_c_10894_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=17.445 //y2=0.995
cc_608 ( N_GND_c_64_p N_noxref_35_c_10894_n ) capacitor c=0.00934524f \
 //x=19.07 //y=0 //x2=17.445 //y2=0.995
cc_609 ( N_GND_c_89_p N_noxref_35_c_10896_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=17.53 //y2=0.625
cc_610 ( N_GND_c_64_p N_noxref_35_c_10896_n ) capacitor c=0.0140928f //x=19.07 \
 //y=0 //x2=17.53 //y2=0.625
cc_611 ( N_GND_M9_noxref_d N_noxref_35_c_10896_n ) capacitor c=6.21394e-19 \
 //x=15.315 //y=0.875 //x2=17.53 //y2=0.625
cc_612 ( N_GND_c_89_p N_noxref_35_c_10899_n ) capacitor c=0.0105197f //x=95.83 \
 //y=0 //x2=18.415 //y2=0.54
cc_613 ( N_GND_c_64_p N_noxref_35_c_10899_n ) capacitor c=0.0364139f //x=19.07 \
 //y=0 //x2=18.415 //y2=0.54
cc_614 ( N_GND_c_89_p N_noxref_35_c_10901_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=18.5 //y2=0.625
cc_615 ( N_GND_c_64_p N_noxref_35_c_10901_n ) capacitor c=0.0140304f //x=19.07 \
 //y=0 //x2=18.5 //y2=0.625
cc_616 ( N_GND_c_6_p N_noxref_35_c_10901_n ) capacitor c=0.0404137f //x=19.24 \
 //y=0 //x2=18.5 //y2=0.625
cc_617 ( N_GND_M9_noxref_d N_noxref_35_M10_noxref_d ) capacitor c=0.00162435f \
 //x=15.315 //y=0.875 //x2=16.29 //y2=0.91
cc_618 ( N_GND_c_5_p N_noxref_35_M11_noxref_s ) capacitor c=8.16352e-19 \
 //x=14.43 //y=0 //x2=17.395 //y2=0.375
cc_619 ( N_GND_c_6_p N_noxref_35_M11_noxref_s ) capacitor c=0.00183204f \
 //x=19.24 //y=0 //x2=17.395 //y2=0.375
cc_620 ( N_GND_c_89_p N_noxref_36_c_10947_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=20.715 //y2=1.59
cc_621 ( N_GND_c_73_p N_noxref_36_c_10947_n ) capacitor c=0.00111448f \
 //x=20.23 //y=0 //x2=20.715 //y2=1.59
cc_622 ( N_GND_c_80_p N_noxref_36_c_10947_n ) capacitor c=0.00180612f \
 //x=23.88 //y=0 //x2=20.715 //y2=1.59
cc_623 ( N_GND_M12_noxref_d N_noxref_36_c_10947_n ) capacitor c=0.00853078f \
 //x=20.125 //y=0.875 //x2=20.715 //y2=1.59
cc_624 ( N_GND_c_89_p N_noxref_36_c_10951_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=20.8 //y2=0.625
cc_625 ( N_GND_c_80_p N_noxref_36_c_10951_n ) capacitor c=0.0140928f //x=23.88 \
 //y=0 //x2=20.8 //y2=0.625
cc_626 ( N_GND_M12_noxref_d N_noxref_36_c_10951_n ) capacitor c=0.033954f \
 //x=20.125 //y=0.875 //x2=20.8 //y2=0.625
cc_627 ( N_GND_c_89_p N_noxref_36_c_10954_n ) capacitor c=0.0104386f //x=95.83 \
 //y=0 //x2=21.685 //y2=0.54
cc_628 ( N_GND_c_80_p N_noxref_36_c_10954_n ) capacitor c=0.0360726f //x=23.88 \
 //y=0 //x2=21.685 //y2=0.54
cc_629 ( N_GND_c_89_p N_noxref_36_M12_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=19.695 //y2=0.375
cc_630 ( N_GND_c_73_p N_noxref_36_M12_noxref_s ) capacitor c=0.0140928f \
 //x=20.23 //y=0 //x2=19.695 //y2=0.375
cc_631 ( N_GND_c_80_p N_noxref_36_M12_noxref_s ) capacitor c=0.0136651f \
 //x=23.88 //y=0 //x2=19.695 //y2=0.375
cc_632 ( N_GND_c_6_p N_noxref_36_M12_noxref_s ) capacitor c=0.0696963f \
 //x=19.24 //y=0 //x2=19.695 //y2=0.375
cc_633 ( N_GND_c_7_p N_noxref_36_M12_noxref_s ) capacitor c=3.31601e-19 \
 //x=24.05 //y=0 //x2=19.695 //y2=0.375
cc_634 ( N_GND_M12_noxref_d N_noxref_36_M12_noxref_s ) capacitor c=0.033718f \
 //x=20.125 //y=0.875 //x2=19.695 //y2=0.375
cc_635 ( N_GND_c_89_p N_noxref_37_c_10999_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=22.255 //y2=0.995
cc_636 ( N_GND_c_80_p N_noxref_37_c_10999_n ) capacitor c=0.00934524f \
 //x=23.88 //y=0 //x2=22.255 //y2=0.995
cc_637 ( N_GND_c_89_p N_noxref_37_c_11001_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=22.34 //y2=0.625
cc_638 ( N_GND_c_80_p N_noxref_37_c_11001_n ) capacitor c=0.0140928f //x=23.88 \
 //y=0 //x2=22.34 //y2=0.625
cc_639 ( N_GND_M12_noxref_d N_noxref_37_c_11001_n ) capacitor c=6.21394e-19 \
 //x=20.125 //y=0.875 //x2=22.34 //y2=0.625
cc_640 ( N_GND_c_89_p N_noxref_37_c_11004_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=23.225 //y2=0.54
cc_641 ( N_GND_c_80_p N_noxref_37_c_11004_n ) capacitor c=0.0363691f //x=23.88 \
 //y=0 //x2=23.225 //y2=0.54
cc_642 ( N_GND_c_89_p N_noxref_37_c_11006_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=23.31 //y2=0.625
cc_643 ( N_GND_c_80_p N_noxref_37_c_11006_n ) capacitor c=0.0140304f //x=23.88 \
 //y=0 //x2=23.31 //y2=0.625
cc_644 ( N_GND_c_7_p N_noxref_37_c_11006_n ) capacitor c=0.0404137f //x=24.05 \
 //y=0 //x2=23.31 //y2=0.625
cc_645 ( N_GND_M12_noxref_d N_noxref_37_M13_noxref_d ) capacitor c=0.00162435f \
 //x=20.125 //y=0.875 //x2=21.1 //y2=0.91
cc_646 ( N_GND_c_6_p N_noxref_37_M14_noxref_s ) capacitor c=8.16352e-19 \
 //x=19.24 //y=0 //x2=22.205 //y2=0.375
cc_647 ( N_GND_c_7_p N_noxref_37_M14_noxref_s ) capacitor c=0.00183204f \
 //x=24.05 //y=0 //x2=22.205 //y2=0.375
cc_648 ( N_GND_c_89_p N_noxref_38_c_11051_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=25.525 //y2=1.59
cc_649 ( N_GND_c_94_p N_noxref_38_c_11051_n ) capacitor c=0.00111448f \
 //x=25.04 //y=0 //x2=25.525 //y2=1.59
cc_650 ( N_GND_c_101_p N_noxref_38_c_11051_n ) capacitor c=0.00180612f \
 //x=28.69 //y=0 //x2=25.525 //y2=1.59
cc_651 ( N_GND_M15_noxref_d N_noxref_38_c_11051_n ) capacitor c=0.00853078f \
 //x=24.935 //y=0.875 //x2=25.525 //y2=1.59
cc_652 ( N_GND_c_89_p N_noxref_38_c_11055_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=25.61 //y2=0.625
cc_653 ( N_GND_c_101_p N_noxref_38_c_11055_n ) capacitor c=0.0140928f \
 //x=28.69 //y=0 //x2=25.61 //y2=0.625
cc_654 ( N_GND_M15_noxref_d N_noxref_38_c_11055_n ) capacitor c=0.033954f \
 //x=24.935 //y=0.875 //x2=25.61 //y2=0.625
cc_655 ( N_GND_c_89_p N_noxref_38_c_11058_n ) capacitor c=0.0104506f //x=95.83 \
 //y=0 //x2=26.495 //y2=0.54
cc_656 ( N_GND_c_101_p N_noxref_38_c_11058_n ) capacitor c=0.0360726f \
 //x=28.69 //y=0 //x2=26.495 //y2=0.54
cc_657 ( N_GND_c_89_p N_noxref_38_M15_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=24.505 //y2=0.375
cc_658 ( N_GND_c_94_p N_noxref_38_M15_noxref_s ) capacitor c=0.0140928f \
 //x=25.04 //y=0 //x2=24.505 //y2=0.375
cc_659 ( N_GND_c_101_p N_noxref_38_M15_noxref_s ) capacitor c=0.0131437f \
 //x=28.69 //y=0 //x2=24.505 //y2=0.375
cc_660 ( N_GND_c_7_p N_noxref_38_M15_noxref_s ) capacitor c=0.0696963f \
 //x=24.05 //y=0 //x2=24.505 //y2=0.375
cc_661 ( N_GND_c_8_p N_noxref_38_M15_noxref_s ) capacitor c=3.31601e-19 \
 //x=28.86 //y=0 //x2=24.505 //y2=0.375
cc_662 ( N_GND_M15_noxref_d N_noxref_38_M15_noxref_s ) capacitor c=0.033718f \
 //x=24.935 //y=0.875 //x2=24.505 //y2=0.375
cc_663 ( N_GND_c_89_p N_noxref_39_c_11100_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=27.065 //y2=0.995
cc_664 ( N_GND_c_101_p N_noxref_39_c_11100_n ) capacitor c=0.00934524f \
 //x=28.69 //y=0 //x2=27.065 //y2=0.995
cc_665 ( N_GND_c_89_p N_noxref_39_c_11102_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=27.15 //y2=0.625
cc_666 ( N_GND_c_101_p N_noxref_39_c_11102_n ) capacitor c=0.0140928f \
 //x=28.69 //y=0 //x2=27.15 //y2=0.625
cc_667 ( N_GND_M15_noxref_d N_noxref_39_c_11102_n ) capacitor c=6.21394e-19 \
 //x=24.935 //y=0.875 //x2=27.15 //y2=0.625
cc_668 ( N_GND_c_89_p N_noxref_39_c_11105_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=28.035 //y2=0.54
cc_669 ( N_GND_c_101_p N_noxref_39_c_11105_n ) capacitor c=0.0364215f \
 //x=28.69 //y=0 //x2=28.035 //y2=0.54
cc_670 ( N_GND_c_89_p N_noxref_39_c_11107_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=28.12 //y2=0.625
cc_671 ( N_GND_c_101_p N_noxref_39_c_11107_n ) capacitor c=0.0140304f \
 //x=28.69 //y=0 //x2=28.12 //y2=0.625
cc_672 ( N_GND_c_8_p N_noxref_39_c_11107_n ) capacitor c=0.0404137f //x=28.86 \
 //y=0 //x2=28.12 //y2=0.625
cc_673 ( N_GND_M15_noxref_d N_noxref_39_M16_noxref_d ) capacitor c=0.00162435f \
 //x=24.935 //y=0.875 //x2=25.91 //y2=0.91
cc_674 ( N_GND_c_7_p N_noxref_39_M17_noxref_s ) capacitor c=8.16352e-19 \
 //x=24.05 //y=0 //x2=27.015 //y2=0.375
cc_675 ( N_GND_c_8_p N_noxref_39_M17_noxref_s ) capacitor c=0.00183204f \
 //x=28.86 //y=0 //x2=27.015 //y2=0.375
cc_676 ( N_GND_c_89_p N_noxref_40_c_11152_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=30.335 //y2=1.59
cc_677 ( N_GND_c_218_p N_noxref_40_c_11152_n ) capacitor c=0.00111448f \
 //x=29.85 //y=0 //x2=30.335 //y2=1.59
cc_678 ( N_GND_c_225_p N_noxref_40_c_11152_n ) capacitor c=0.00180612f \
 //x=33.5 //y=0 //x2=30.335 //y2=1.59
cc_679 ( N_GND_M18_noxref_d N_noxref_40_c_11152_n ) capacitor c=0.00853078f \
 //x=29.745 //y=0.875 //x2=30.335 //y2=1.59
cc_680 ( N_GND_c_89_p N_noxref_40_c_11156_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=30.42 //y2=0.625
cc_681 ( N_GND_c_225_p N_noxref_40_c_11156_n ) capacitor c=0.0140928f //x=33.5 \
 //y=0 //x2=30.42 //y2=0.625
cc_682 ( N_GND_M18_noxref_d N_noxref_40_c_11156_n ) capacitor c=0.033954f \
 //x=29.745 //y=0.875 //x2=30.42 //y2=0.625
cc_683 ( N_GND_c_89_p N_noxref_40_c_11159_n ) capacitor c=0.0104386f //x=95.83 \
 //y=0 //x2=31.305 //y2=0.54
cc_684 ( N_GND_c_225_p N_noxref_40_c_11159_n ) capacitor c=0.0360726f //x=33.5 \
 //y=0 //x2=31.305 //y2=0.54
cc_685 ( N_GND_c_89_p N_noxref_40_M18_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=29.315 //y2=0.375
cc_686 ( N_GND_c_218_p N_noxref_40_M18_noxref_s ) capacitor c=0.0140928f \
 //x=29.85 //y=0 //x2=29.315 //y2=0.375
cc_687 ( N_GND_c_225_p N_noxref_40_M18_noxref_s ) capacitor c=0.0131437f \
 //x=33.5 //y=0 //x2=29.315 //y2=0.375
cc_688 ( N_GND_c_8_p N_noxref_40_M18_noxref_s ) capacitor c=0.0696963f \
 //x=28.86 //y=0 //x2=29.315 //y2=0.375
cc_689 ( N_GND_c_9_p N_noxref_40_M18_noxref_s ) capacitor c=3.31601e-19 \
 //x=33.67 //y=0 //x2=29.315 //y2=0.375
cc_690 ( N_GND_M18_noxref_d N_noxref_40_M18_noxref_s ) capacitor c=0.033718f \
 //x=29.745 //y=0.875 //x2=29.315 //y2=0.375
cc_691 ( N_GND_c_89_p N_noxref_41_c_11204_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=31.875 //y2=0.995
cc_692 ( N_GND_c_225_p N_noxref_41_c_11204_n ) capacitor c=0.00934524f \
 //x=33.5 //y=0 //x2=31.875 //y2=0.995
cc_693 ( N_GND_c_89_p N_noxref_41_c_11206_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=31.96 //y2=0.625
cc_694 ( N_GND_c_225_p N_noxref_41_c_11206_n ) capacitor c=0.0140928f //x=33.5 \
 //y=0 //x2=31.96 //y2=0.625
cc_695 ( N_GND_M18_noxref_d N_noxref_41_c_11206_n ) capacitor c=6.21394e-19 \
 //x=29.745 //y=0.875 //x2=31.96 //y2=0.625
cc_696 ( N_GND_c_89_p N_noxref_41_c_11209_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=32.845 //y2=0.54
cc_697 ( N_GND_c_225_p N_noxref_41_c_11209_n ) capacitor c=0.0363691f //x=33.5 \
 //y=0 //x2=32.845 //y2=0.54
cc_698 ( N_GND_c_89_p N_noxref_41_c_11211_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=32.93 //y2=0.625
cc_699 ( N_GND_c_225_p N_noxref_41_c_11211_n ) capacitor c=0.0140304f //x=33.5 \
 //y=0 //x2=32.93 //y2=0.625
cc_700 ( N_GND_c_9_p N_noxref_41_c_11211_n ) capacitor c=0.0404137f //x=33.67 \
 //y=0 //x2=32.93 //y2=0.625
cc_701 ( N_GND_M18_noxref_d N_noxref_41_M19_noxref_d ) capacitor c=0.00162435f \
 //x=29.745 //y=0.875 //x2=30.72 //y2=0.91
cc_702 ( N_GND_c_8_p N_noxref_41_M20_noxref_s ) capacitor c=8.16352e-19 \
 //x=28.86 //y=0 //x2=31.825 //y2=0.375
cc_703 ( N_GND_c_9_p N_noxref_41_M20_noxref_s ) capacitor c=0.00183204f \
 //x=33.67 //y=0 //x2=31.825 //y2=0.375
cc_704 ( N_GND_c_89_p N_noxref_42_c_11256_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=35.145 //y2=1.59
cc_705 ( N_GND_c_141_p N_noxref_42_c_11256_n ) capacitor c=0.00111448f \
 //x=34.66 //y=0 //x2=35.145 //y2=1.59
cc_706 ( N_GND_c_148_p N_noxref_42_c_11256_n ) capacitor c=0.00180612f \
 //x=38.31 //y=0 //x2=35.145 //y2=1.59
cc_707 ( N_GND_M21_noxref_d N_noxref_42_c_11256_n ) capacitor c=0.00853078f \
 //x=34.555 //y=0.875 //x2=35.145 //y2=1.59
cc_708 ( N_GND_c_89_p N_noxref_42_c_11260_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=35.23 //y2=0.625
cc_709 ( N_GND_c_148_p N_noxref_42_c_11260_n ) capacitor c=0.0140928f \
 //x=38.31 //y=0 //x2=35.23 //y2=0.625
cc_710 ( N_GND_M21_noxref_d N_noxref_42_c_11260_n ) capacitor c=0.033954f \
 //x=34.555 //y=0.875 //x2=35.23 //y2=0.625
cc_711 ( N_GND_c_89_p N_noxref_42_c_11263_n ) capacitor c=0.0104506f //x=95.83 \
 //y=0 //x2=36.115 //y2=0.54
cc_712 ( N_GND_c_148_p N_noxref_42_c_11263_n ) capacitor c=0.0360726f \
 //x=38.31 //y=0 //x2=36.115 //y2=0.54
cc_713 ( N_GND_c_89_p N_noxref_42_M21_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=34.125 //y2=0.375
cc_714 ( N_GND_c_141_p N_noxref_42_M21_noxref_s ) capacitor c=0.0140928f \
 //x=34.66 //y=0 //x2=34.125 //y2=0.375
cc_715 ( N_GND_c_148_p N_noxref_42_M21_noxref_s ) capacitor c=0.0131437f \
 //x=38.31 //y=0 //x2=34.125 //y2=0.375
cc_716 ( N_GND_c_9_p N_noxref_42_M21_noxref_s ) capacitor c=0.0696963f \
 //x=33.67 //y=0 //x2=34.125 //y2=0.375
cc_717 ( N_GND_c_10_p N_noxref_42_M21_noxref_s ) capacitor c=3.31601e-19 \
 //x=38.48 //y=0 //x2=34.125 //y2=0.375
cc_718 ( N_GND_M21_noxref_d N_noxref_42_M21_noxref_s ) capacitor c=0.033718f \
 //x=34.555 //y=0.875 //x2=34.125 //y2=0.375
cc_719 ( N_GND_c_89_p N_noxref_43_c_11305_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=36.685 //y2=0.995
cc_720 ( N_GND_c_148_p N_noxref_43_c_11305_n ) capacitor c=0.00934524f \
 //x=38.31 //y=0 //x2=36.685 //y2=0.995
cc_721 ( N_GND_c_89_p N_noxref_43_c_11307_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=36.77 //y2=0.625
cc_722 ( N_GND_c_148_p N_noxref_43_c_11307_n ) capacitor c=0.0140928f \
 //x=38.31 //y=0 //x2=36.77 //y2=0.625
cc_723 ( N_GND_M21_noxref_d N_noxref_43_c_11307_n ) capacitor c=6.21394e-19 \
 //x=34.555 //y=0.875 //x2=36.77 //y2=0.625
cc_724 ( N_GND_c_89_p N_noxref_43_c_11310_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=37.655 //y2=0.54
cc_725 ( N_GND_c_148_p N_noxref_43_c_11310_n ) capacitor c=0.0364215f \
 //x=38.31 //y=0 //x2=37.655 //y2=0.54
cc_726 ( N_GND_c_89_p N_noxref_43_c_11312_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=37.74 //y2=0.625
cc_727 ( N_GND_c_148_p N_noxref_43_c_11312_n ) capacitor c=0.0140304f \
 //x=38.31 //y=0 //x2=37.74 //y2=0.625
cc_728 ( N_GND_c_10_p N_noxref_43_c_11312_n ) capacitor c=0.0404137f //x=38.48 \
 //y=0 //x2=37.74 //y2=0.625
cc_729 ( N_GND_M21_noxref_d N_noxref_43_M22_noxref_d ) capacitor c=0.00162435f \
 //x=34.555 //y=0.875 //x2=35.53 //y2=0.91
cc_730 ( N_GND_c_9_p N_noxref_43_M23_noxref_s ) capacitor c=8.16352e-19 \
 //x=33.67 //y=0 //x2=36.635 //y2=0.375
cc_731 ( N_GND_c_10_p N_noxref_43_M23_noxref_s ) capacitor c=0.00183204f \
 //x=38.48 //y=0 //x2=36.635 //y2=0.375
cc_732 ( N_GND_c_89_p N_noxref_44_c_11357_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=39.955 //y2=1.59
cc_733 ( N_GND_c_151_p N_noxref_44_c_11357_n ) capacitor c=0.00111448f \
 //x=39.47 //y=0 //x2=39.955 //y2=1.59
cc_734 ( N_GND_c_158_p N_noxref_44_c_11357_n ) capacitor c=0.00180612f \
 //x=43.12 //y=0 //x2=39.955 //y2=1.59
cc_735 ( N_GND_M24_noxref_d N_noxref_44_c_11357_n ) capacitor c=0.00853078f \
 //x=39.365 //y=0.875 //x2=39.955 //y2=1.59
cc_736 ( N_GND_c_89_p N_noxref_44_c_11361_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=40.04 //y2=0.625
cc_737 ( N_GND_c_158_p N_noxref_44_c_11361_n ) capacitor c=0.0140928f \
 //x=43.12 //y=0 //x2=40.04 //y2=0.625
cc_738 ( N_GND_M24_noxref_d N_noxref_44_c_11361_n ) capacitor c=0.033954f \
 //x=39.365 //y=0.875 //x2=40.04 //y2=0.625
cc_739 ( N_GND_c_89_p N_noxref_44_c_11364_n ) capacitor c=0.0104506f //x=95.83 \
 //y=0 //x2=40.925 //y2=0.54
cc_740 ( N_GND_c_158_p N_noxref_44_c_11364_n ) capacitor c=0.0360726f \
 //x=43.12 //y=0 //x2=40.925 //y2=0.54
cc_741 ( N_GND_c_89_p N_noxref_44_M24_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=38.935 //y2=0.375
cc_742 ( N_GND_c_151_p N_noxref_44_M24_noxref_s ) capacitor c=0.0140928f \
 //x=39.47 //y=0 //x2=38.935 //y2=0.375
cc_743 ( N_GND_c_158_p N_noxref_44_M24_noxref_s ) capacitor c=0.0131437f \
 //x=43.12 //y=0 //x2=38.935 //y2=0.375
cc_744 ( N_GND_c_10_p N_noxref_44_M24_noxref_s ) capacitor c=0.0696963f \
 //x=38.48 //y=0 //x2=38.935 //y2=0.375
cc_745 ( N_GND_c_11_p N_noxref_44_M24_noxref_s ) capacitor c=3.31601e-19 \
 //x=43.29 //y=0 //x2=38.935 //y2=0.375
cc_746 ( N_GND_M24_noxref_d N_noxref_44_M24_noxref_s ) capacitor c=0.033718f \
 //x=39.365 //y=0.875 //x2=38.935 //y2=0.375
cc_747 ( N_GND_c_89_p N_noxref_45_c_11406_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=41.495 //y2=0.995
cc_748 ( N_GND_c_158_p N_noxref_45_c_11406_n ) capacitor c=0.00934524f \
 //x=43.12 //y=0 //x2=41.495 //y2=0.995
cc_749 ( N_GND_c_89_p N_noxref_45_c_11408_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=41.58 //y2=0.625
cc_750 ( N_GND_c_158_p N_noxref_45_c_11408_n ) capacitor c=0.0140928f \
 //x=43.12 //y=0 //x2=41.58 //y2=0.625
cc_751 ( N_GND_M24_noxref_d N_noxref_45_c_11408_n ) capacitor c=6.21394e-19 \
 //x=39.365 //y=0.875 //x2=41.58 //y2=0.625
cc_752 ( N_GND_c_89_p N_noxref_45_c_11411_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=42.465 //y2=0.54
cc_753 ( N_GND_c_158_p N_noxref_45_c_11411_n ) capacitor c=0.0364215f \
 //x=43.12 //y=0 //x2=42.465 //y2=0.54
cc_754 ( N_GND_c_89_p N_noxref_45_c_11413_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=42.55 //y2=0.625
cc_755 ( N_GND_c_158_p N_noxref_45_c_11413_n ) capacitor c=0.0140304f \
 //x=43.12 //y=0 //x2=42.55 //y2=0.625
cc_756 ( N_GND_c_11_p N_noxref_45_c_11413_n ) capacitor c=0.0404137f //x=43.29 \
 //y=0 //x2=42.55 //y2=0.625
cc_757 ( N_GND_M24_noxref_d N_noxref_45_M25_noxref_d ) capacitor c=0.00162435f \
 //x=39.365 //y=0.875 //x2=40.34 //y2=0.91
cc_758 ( N_GND_c_10_p N_noxref_45_M26_noxref_s ) capacitor c=8.16352e-19 \
 //x=38.48 //y=0 //x2=41.445 //y2=0.375
cc_759 ( N_GND_c_11_p N_noxref_45_M26_noxref_s ) capacitor c=0.00183204f \
 //x=43.29 //y=0 //x2=41.445 //y2=0.375
cc_760 ( N_GND_c_89_p N_noxref_46_c_11458_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=44.765 //y2=1.59
cc_761 ( N_GND_c_167_p N_noxref_46_c_11458_n ) capacitor c=0.00111448f \
 //x=44.28 //y=0 //x2=44.765 //y2=1.59
cc_762 ( N_GND_c_174_p N_noxref_46_c_11458_n ) capacitor c=0.00180612f \
 //x=47.93 //y=0 //x2=44.765 //y2=1.59
cc_763 ( N_GND_M27_noxref_d N_noxref_46_c_11458_n ) capacitor c=0.00853078f \
 //x=44.175 //y=0.875 //x2=44.765 //y2=1.59
cc_764 ( N_GND_c_89_p N_noxref_46_c_11462_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=44.85 //y2=0.625
cc_765 ( N_GND_c_174_p N_noxref_46_c_11462_n ) capacitor c=0.0140928f \
 //x=47.93 //y=0 //x2=44.85 //y2=0.625
cc_766 ( N_GND_M27_noxref_d N_noxref_46_c_11462_n ) capacitor c=0.033954f \
 //x=44.175 //y=0.875 //x2=44.85 //y2=0.625
cc_767 ( N_GND_c_89_p N_noxref_46_c_11465_n ) capacitor c=0.0104506f //x=95.83 \
 //y=0 //x2=45.735 //y2=0.54
cc_768 ( N_GND_c_174_p N_noxref_46_c_11465_n ) capacitor c=0.0360726f \
 //x=47.93 //y=0 //x2=45.735 //y2=0.54
cc_769 ( N_GND_c_89_p N_noxref_46_M27_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=43.745 //y2=0.375
cc_770 ( N_GND_c_167_p N_noxref_46_M27_noxref_s ) capacitor c=0.0140928f \
 //x=44.28 //y=0 //x2=43.745 //y2=0.375
cc_771 ( N_GND_c_174_p N_noxref_46_M27_noxref_s ) capacitor c=0.0131437f \
 //x=47.93 //y=0 //x2=43.745 //y2=0.375
cc_772 ( N_GND_c_11_p N_noxref_46_M27_noxref_s ) capacitor c=0.0696963f \
 //x=43.29 //y=0 //x2=43.745 //y2=0.375
cc_773 ( N_GND_c_12_p N_noxref_46_M27_noxref_s ) capacitor c=3.31601e-19 \
 //x=48.1 //y=0 //x2=43.745 //y2=0.375
cc_774 ( N_GND_M27_noxref_d N_noxref_46_M27_noxref_s ) capacitor c=0.033718f \
 //x=44.175 //y=0.875 //x2=43.745 //y2=0.375
cc_775 ( N_GND_c_89_p N_noxref_47_c_11507_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=46.305 //y2=0.995
cc_776 ( N_GND_c_174_p N_noxref_47_c_11507_n ) capacitor c=0.00934524f \
 //x=47.93 //y=0 //x2=46.305 //y2=0.995
cc_777 ( N_GND_c_89_p N_noxref_47_c_11509_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=46.39 //y2=0.625
cc_778 ( N_GND_c_174_p N_noxref_47_c_11509_n ) capacitor c=0.0140928f \
 //x=47.93 //y=0 //x2=46.39 //y2=0.625
cc_779 ( N_GND_M27_noxref_d N_noxref_47_c_11509_n ) capacitor c=6.21394e-19 \
 //x=44.175 //y=0.875 //x2=46.39 //y2=0.625
cc_780 ( N_GND_c_89_p N_noxref_47_c_11512_n ) capacitor c=0.0105197f //x=95.83 \
 //y=0 //x2=47.275 //y2=0.54
cc_781 ( N_GND_c_174_p N_noxref_47_c_11512_n ) capacitor c=0.0364139f \
 //x=47.93 //y=0 //x2=47.275 //y2=0.54
cc_782 ( N_GND_c_89_p N_noxref_47_c_11514_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=47.36 //y2=0.625
cc_783 ( N_GND_c_174_p N_noxref_47_c_11514_n ) capacitor c=0.0140304f \
 //x=47.93 //y=0 //x2=47.36 //y2=0.625
cc_784 ( N_GND_c_12_p N_noxref_47_c_11514_n ) capacitor c=0.0404137f //x=48.1 \
 //y=0 //x2=47.36 //y2=0.625
cc_785 ( N_GND_M27_noxref_d N_noxref_47_M28_noxref_d ) capacitor c=0.00162435f \
 //x=44.175 //y=0.875 //x2=45.15 //y2=0.91
cc_786 ( N_GND_c_11_p N_noxref_47_M29_noxref_s ) capacitor c=8.16352e-19 \
 //x=43.29 //y=0 //x2=46.255 //y2=0.375
cc_787 ( N_GND_c_12_p N_noxref_47_M29_noxref_s ) capacitor c=0.00183204f \
 //x=48.1 //y=0 //x2=46.255 //y2=0.375
cc_788 ( N_GND_c_89_p N_noxref_48_c_11560_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=49.575 //y2=1.59
cc_789 ( N_GND_c_181_p N_noxref_48_c_11560_n ) capacitor c=0.00111448f \
 //x=49.09 //y=0 //x2=49.575 //y2=1.59
cc_790 ( N_GND_c_188_p N_noxref_48_c_11560_n ) capacitor c=0.00180612f \
 //x=52.74 //y=0 //x2=49.575 //y2=1.59
cc_791 ( N_GND_M30_noxref_d N_noxref_48_c_11560_n ) capacitor c=0.00853078f \
 //x=48.985 //y=0.875 //x2=49.575 //y2=1.59
cc_792 ( N_GND_c_89_p N_noxref_48_c_11564_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=49.66 //y2=0.625
cc_793 ( N_GND_c_188_p N_noxref_48_c_11564_n ) capacitor c=0.0140928f \
 //x=52.74 //y=0 //x2=49.66 //y2=0.625
cc_794 ( N_GND_M30_noxref_d N_noxref_48_c_11564_n ) capacitor c=0.033954f \
 //x=48.985 //y=0.875 //x2=49.66 //y2=0.625
cc_795 ( N_GND_c_89_p N_noxref_48_c_11567_n ) capacitor c=0.0104386f //x=95.83 \
 //y=0 //x2=50.545 //y2=0.54
cc_796 ( N_GND_c_188_p N_noxref_48_c_11567_n ) capacitor c=0.0360726f \
 //x=52.74 //y=0 //x2=50.545 //y2=0.54
cc_797 ( N_GND_c_89_p N_noxref_48_M30_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=48.555 //y2=0.375
cc_798 ( N_GND_c_181_p N_noxref_48_M30_noxref_s ) capacitor c=0.0140928f \
 //x=49.09 //y=0 //x2=48.555 //y2=0.375
cc_799 ( N_GND_c_188_p N_noxref_48_M30_noxref_s ) capacitor c=0.0136651f \
 //x=52.74 //y=0 //x2=48.555 //y2=0.375
cc_800 ( N_GND_c_12_p N_noxref_48_M30_noxref_s ) capacitor c=0.0696963f \
 //x=48.1 //y=0 //x2=48.555 //y2=0.375
cc_801 ( N_GND_c_13_p N_noxref_48_M30_noxref_s ) capacitor c=3.31601e-19 \
 //x=52.91 //y=0 //x2=48.555 //y2=0.375
cc_802 ( N_GND_M30_noxref_d N_noxref_48_M30_noxref_s ) capacitor c=0.033718f \
 //x=48.985 //y=0.875 //x2=48.555 //y2=0.375
cc_803 ( N_GND_c_89_p N_noxref_49_c_11612_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=51.115 //y2=0.995
cc_804 ( N_GND_c_188_p N_noxref_49_c_11612_n ) capacitor c=0.00934524f \
 //x=52.74 //y=0 //x2=51.115 //y2=0.995
cc_805 ( N_GND_c_89_p N_noxref_49_c_11614_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=51.2 //y2=0.625
cc_806 ( N_GND_c_188_p N_noxref_49_c_11614_n ) capacitor c=0.0140928f \
 //x=52.74 //y=0 //x2=51.2 //y2=0.625
cc_807 ( N_GND_M30_noxref_d N_noxref_49_c_11614_n ) capacitor c=6.21394e-19 \
 //x=48.985 //y=0.875 //x2=51.2 //y2=0.625
cc_808 ( N_GND_c_89_p N_noxref_49_c_11617_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=52.085 //y2=0.54
cc_809 ( N_GND_c_188_p N_noxref_49_c_11617_n ) capacitor c=0.0363691f \
 //x=52.74 //y=0 //x2=52.085 //y2=0.54
cc_810 ( N_GND_c_89_p N_noxref_49_c_11619_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=52.17 //y2=0.625
cc_811 ( N_GND_c_188_p N_noxref_49_c_11619_n ) capacitor c=0.0140304f \
 //x=52.74 //y=0 //x2=52.17 //y2=0.625
cc_812 ( N_GND_c_13_p N_noxref_49_c_11619_n ) capacitor c=0.0404137f //x=52.91 \
 //y=0 //x2=52.17 //y2=0.625
cc_813 ( N_GND_M30_noxref_d N_noxref_49_M31_noxref_d ) capacitor c=0.00162435f \
 //x=48.985 //y=0.875 //x2=49.96 //y2=0.91
cc_814 ( N_GND_c_12_p N_noxref_49_M32_noxref_s ) capacitor c=8.16352e-19 \
 //x=48.1 //y=0 //x2=51.065 //y2=0.375
cc_815 ( N_GND_c_13_p N_noxref_49_M32_noxref_s ) capacitor c=0.00183204f \
 //x=52.91 //y=0 //x2=51.065 //y2=0.375
cc_816 ( N_GND_c_89_p N_noxref_50_c_11664_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=54.385 //y2=1.59
cc_817 ( N_GND_c_347_p N_noxref_50_c_11664_n ) capacitor c=0.00111448f \
 //x=53.9 //y=0 //x2=54.385 //y2=1.59
cc_818 ( N_GND_c_348_p N_noxref_50_c_11664_n ) capacitor c=0.00180612f \
 //x=57.55 //y=0 //x2=54.385 //y2=1.59
cc_819 ( N_GND_M33_noxref_d N_noxref_50_c_11664_n ) capacitor c=0.00853078f \
 //x=53.795 //y=0.875 //x2=54.385 //y2=1.59
cc_820 ( N_GND_c_89_p N_noxref_50_c_11668_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=54.47 //y2=0.625
cc_821 ( N_GND_c_348_p N_noxref_50_c_11668_n ) capacitor c=0.0140928f \
 //x=57.55 //y=0 //x2=54.47 //y2=0.625
cc_822 ( N_GND_M33_noxref_d N_noxref_50_c_11668_n ) capacitor c=0.033954f \
 //x=53.795 //y=0.875 //x2=54.47 //y2=0.625
cc_823 ( N_GND_c_89_p N_noxref_50_c_11671_n ) capacitor c=0.0104506f //x=95.83 \
 //y=0 //x2=55.355 //y2=0.54
cc_824 ( N_GND_c_348_p N_noxref_50_c_11671_n ) capacitor c=0.0360726f \
 //x=57.55 //y=0 //x2=55.355 //y2=0.54
cc_825 ( N_GND_c_89_p N_noxref_50_M33_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=53.365 //y2=0.375
cc_826 ( N_GND_c_347_p N_noxref_50_M33_noxref_s ) capacitor c=0.0140928f \
 //x=53.9 //y=0 //x2=53.365 //y2=0.375
cc_827 ( N_GND_c_348_p N_noxref_50_M33_noxref_s ) capacitor c=0.0136651f \
 //x=57.55 //y=0 //x2=53.365 //y2=0.375
cc_828 ( N_GND_c_13_p N_noxref_50_M33_noxref_s ) capacitor c=0.0696963f \
 //x=52.91 //y=0 //x2=53.365 //y2=0.375
cc_829 ( N_GND_c_14_p N_noxref_50_M33_noxref_s ) capacitor c=3.31601e-19 \
 //x=57.72 //y=0 //x2=53.365 //y2=0.375
cc_830 ( N_GND_M33_noxref_d N_noxref_50_M33_noxref_s ) capacitor c=0.033718f \
 //x=53.795 //y=0.875 //x2=53.365 //y2=0.375
cc_831 ( N_GND_c_89_p N_noxref_51_c_11713_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=55.925 //y2=0.995
cc_832 ( N_GND_c_348_p N_noxref_51_c_11713_n ) capacitor c=0.00934524f \
 //x=57.55 //y=0 //x2=55.925 //y2=0.995
cc_833 ( N_GND_c_89_p N_noxref_51_c_11715_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=56.01 //y2=0.625
cc_834 ( N_GND_c_348_p N_noxref_51_c_11715_n ) capacitor c=0.0140928f \
 //x=57.55 //y=0 //x2=56.01 //y2=0.625
cc_835 ( N_GND_M33_noxref_d N_noxref_51_c_11715_n ) capacitor c=6.21394e-19 \
 //x=53.795 //y=0.875 //x2=56.01 //y2=0.625
cc_836 ( N_GND_c_89_p N_noxref_51_c_11718_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=56.895 //y2=0.54
cc_837 ( N_GND_c_348_p N_noxref_51_c_11718_n ) capacitor c=0.0364215f \
 //x=57.55 //y=0 //x2=56.895 //y2=0.54
cc_838 ( N_GND_c_89_p N_noxref_51_c_11720_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=56.98 //y2=0.625
cc_839 ( N_GND_c_348_p N_noxref_51_c_11720_n ) capacitor c=0.0140304f \
 //x=57.55 //y=0 //x2=56.98 //y2=0.625
cc_840 ( N_GND_c_14_p N_noxref_51_c_11720_n ) capacitor c=0.0404137f //x=57.72 \
 //y=0 //x2=56.98 //y2=0.625
cc_841 ( N_GND_M33_noxref_d N_noxref_51_M34_noxref_d ) capacitor c=0.00162435f \
 //x=53.795 //y=0.875 //x2=54.77 //y2=0.91
cc_842 ( N_GND_c_13_p N_noxref_51_M35_noxref_s ) capacitor c=8.16352e-19 \
 //x=52.91 //y=0 //x2=55.875 //y2=0.375
cc_843 ( N_GND_c_14_p N_noxref_51_M35_noxref_s ) capacitor c=0.00183204f \
 //x=57.72 //y=0 //x2=55.875 //y2=0.375
cc_844 ( N_GND_c_89_p N_noxref_52_c_11765_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=59.195 //y2=1.59
cc_845 ( N_GND_c_228_p N_noxref_52_c_11765_n ) capacitor c=0.00111448f \
 //x=58.71 //y=0 //x2=59.195 //y2=1.59
cc_846 ( N_GND_c_235_p N_noxref_52_c_11765_n ) capacitor c=0.00180612f \
 //x=62.36 //y=0 //x2=59.195 //y2=1.59
cc_847 ( N_GND_M36_noxref_d N_noxref_52_c_11765_n ) capacitor c=0.00853078f \
 //x=58.605 //y=0.875 //x2=59.195 //y2=1.59
cc_848 ( N_GND_c_89_p N_noxref_52_c_11769_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=59.28 //y2=0.625
cc_849 ( N_GND_c_235_p N_noxref_52_c_11769_n ) capacitor c=0.0140928f \
 //x=62.36 //y=0 //x2=59.28 //y2=0.625
cc_850 ( N_GND_M36_noxref_d N_noxref_52_c_11769_n ) capacitor c=0.033954f \
 //x=58.605 //y=0.875 //x2=59.28 //y2=0.625
cc_851 ( N_GND_c_89_p N_noxref_52_c_11772_n ) capacitor c=0.0104386f //x=95.83 \
 //y=0 //x2=60.165 //y2=0.54
cc_852 ( N_GND_c_235_p N_noxref_52_c_11772_n ) capacitor c=0.0360726f \
 //x=62.36 //y=0 //x2=60.165 //y2=0.54
cc_853 ( N_GND_c_89_p N_noxref_52_M36_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=58.175 //y2=0.375
cc_854 ( N_GND_c_228_p N_noxref_52_M36_noxref_s ) capacitor c=0.0140928f \
 //x=58.71 //y=0 //x2=58.175 //y2=0.375
cc_855 ( N_GND_c_235_p N_noxref_52_M36_noxref_s ) capacitor c=0.0136651f \
 //x=62.36 //y=0 //x2=58.175 //y2=0.375
cc_856 ( N_GND_c_14_p N_noxref_52_M36_noxref_s ) capacitor c=0.0696963f \
 //x=57.72 //y=0 //x2=58.175 //y2=0.375
cc_857 ( N_GND_c_15_p N_noxref_52_M36_noxref_s ) capacitor c=3.31601e-19 \
 //x=62.53 //y=0 //x2=58.175 //y2=0.375
cc_858 ( N_GND_M36_noxref_d N_noxref_52_M36_noxref_s ) capacitor c=0.033718f \
 //x=58.605 //y=0.875 //x2=58.175 //y2=0.375
cc_859 ( N_GND_c_89_p N_noxref_53_c_11817_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=60.735 //y2=0.995
cc_860 ( N_GND_c_235_p N_noxref_53_c_11817_n ) capacitor c=0.00934524f \
 //x=62.36 //y=0 //x2=60.735 //y2=0.995
cc_861 ( N_GND_c_89_p N_noxref_53_c_11819_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=60.82 //y2=0.625
cc_862 ( N_GND_c_235_p N_noxref_53_c_11819_n ) capacitor c=0.0140928f \
 //x=62.36 //y=0 //x2=60.82 //y2=0.625
cc_863 ( N_GND_M36_noxref_d N_noxref_53_c_11819_n ) capacitor c=6.21394e-19 \
 //x=58.605 //y=0.875 //x2=60.82 //y2=0.625
cc_864 ( N_GND_c_89_p N_noxref_53_c_11822_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=61.705 //y2=0.54
cc_865 ( N_GND_c_235_p N_noxref_53_c_11822_n ) capacitor c=0.0363691f \
 //x=62.36 //y=0 //x2=61.705 //y2=0.54
cc_866 ( N_GND_c_89_p N_noxref_53_c_11824_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=61.79 //y2=0.625
cc_867 ( N_GND_c_235_p N_noxref_53_c_11824_n ) capacitor c=0.0140304f \
 //x=62.36 //y=0 //x2=61.79 //y2=0.625
cc_868 ( N_GND_c_15_p N_noxref_53_c_11824_n ) capacitor c=0.0404137f //x=62.53 \
 //y=0 //x2=61.79 //y2=0.625
cc_869 ( N_GND_M36_noxref_d N_noxref_53_M37_noxref_d ) capacitor c=0.00162435f \
 //x=58.605 //y=0.875 //x2=59.58 //y2=0.91
cc_870 ( N_GND_c_14_p N_noxref_53_M38_noxref_s ) capacitor c=8.16352e-19 \
 //x=57.72 //y=0 //x2=60.685 //y2=0.375
cc_871 ( N_GND_c_15_p N_noxref_53_M38_noxref_s ) capacitor c=0.00183204f \
 //x=62.53 //y=0 //x2=60.685 //y2=0.375
cc_872 ( N_GND_c_89_p N_noxref_54_c_11869_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=64.005 //y2=1.59
cc_873 ( N_GND_c_246_p N_noxref_54_c_11869_n ) capacitor c=0.00111448f \
 //x=63.52 //y=0 //x2=64.005 //y2=1.59
cc_874 ( N_GND_c_253_p N_noxref_54_c_11869_n ) capacitor c=0.00180612f \
 //x=67.17 //y=0 //x2=64.005 //y2=1.59
cc_875 ( N_GND_M39_noxref_d N_noxref_54_c_11869_n ) capacitor c=0.00853078f \
 //x=63.415 //y=0.875 //x2=64.005 //y2=1.59
cc_876 ( N_GND_c_89_p N_noxref_54_c_11873_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=64.09 //y2=0.625
cc_877 ( N_GND_c_253_p N_noxref_54_c_11873_n ) capacitor c=0.0140928f \
 //x=67.17 //y=0 //x2=64.09 //y2=0.625
cc_878 ( N_GND_M39_noxref_d N_noxref_54_c_11873_n ) capacitor c=0.033954f \
 //x=63.415 //y=0.875 //x2=64.09 //y2=0.625
cc_879 ( N_GND_c_89_p N_noxref_54_c_11876_n ) capacitor c=0.0104506f //x=95.83 \
 //y=0 //x2=64.975 //y2=0.54
cc_880 ( N_GND_c_253_p N_noxref_54_c_11876_n ) capacitor c=0.0360726f \
 //x=67.17 //y=0 //x2=64.975 //y2=0.54
cc_881 ( N_GND_c_89_p N_noxref_54_M39_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=62.985 //y2=0.375
cc_882 ( N_GND_c_246_p N_noxref_54_M39_noxref_s ) capacitor c=0.0140928f \
 //x=63.52 //y=0 //x2=62.985 //y2=0.375
cc_883 ( N_GND_c_253_p N_noxref_54_M39_noxref_s ) capacitor c=0.0136651f \
 //x=67.17 //y=0 //x2=62.985 //y2=0.375
cc_884 ( N_GND_c_15_p N_noxref_54_M39_noxref_s ) capacitor c=0.0696963f \
 //x=62.53 //y=0 //x2=62.985 //y2=0.375
cc_885 ( N_GND_c_16_p N_noxref_54_M39_noxref_s ) capacitor c=3.31601e-19 \
 //x=67.34 //y=0 //x2=62.985 //y2=0.375
cc_886 ( N_GND_M39_noxref_d N_noxref_54_M39_noxref_s ) capacitor c=0.033718f \
 //x=63.415 //y=0.875 //x2=62.985 //y2=0.375
cc_887 ( N_GND_c_89_p N_noxref_55_c_11918_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=65.545 //y2=0.995
cc_888 ( N_GND_c_253_p N_noxref_55_c_11918_n ) capacitor c=0.00934524f \
 //x=67.17 //y=0 //x2=65.545 //y2=0.995
cc_889 ( N_GND_c_89_p N_noxref_55_c_11920_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=65.63 //y2=0.625
cc_890 ( N_GND_c_253_p N_noxref_55_c_11920_n ) capacitor c=0.0140928f \
 //x=67.17 //y=0 //x2=65.63 //y2=0.625
cc_891 ( N_GND_M39_noxref_d N_noxref_55_c_11920_n ) capacitor c=6.21394e-19 \
 //x=63.415 //y=0.875 //x2=65.63 //y2=0.625
cc_892 ( N_GND_c_89_p N_noxref_55_c_11923_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=66.515 //y2=0.54
cc_893 ( N_GND_c_253_p N_noxref_55_c_11923_n ) capacitor c=0.0364215f \
 //x=67.17 //y=0 //x2=66.515 //y2=0.54
cc_894 ( N_GND_c_89_p N_noxref_55_c_11925_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=66.6 //y2=0.625
cc_895 ( N_GND_c_253_p N_noxref_55_c_11925_n ) capacitor c=0.0140304f \
 //x=67.17 //y=0 //x2=66.6 //y2=0.625
cc_896 ( N_GND_c_16_p N_noxref_55_c_11925_n ) capacitor c=0.0404137f //x=67.34 \
 //y=0 //x2=66.6 //y2=0.625
cc_897 ( N_GND_M39_noxref_d N_noxref_55_M40_noxref_d ) capacitor c=0.00162435f \
 //x=63.415 //y=0.875 //x2=64.39 //y2=0.91
cc_898 ( N_GND_c_15_p N_noxref_55_M41_noxref_s ) capacitor c=8.16352e-19 \
 //x=62.53 //y=0 //x2=65.495 //y2=0.375
cc_899 ( N_GND_c_16_p N_noxref_55_M41_noxref_s ) capacitor c=0.00183204f \
 //x=67.34 //y=0 //x2=65.495 //y2=0.375
cc_900 ( N_GND_c_89_p N_noxref_56_c_11970_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=68.815 //y2=1.59
cc_901 ( N_GND_c_256_p N_noxref_56_c_11970_n ) capacitor c=0.00111448f \
 //x=68.33 //y=0 //x2=68.815 //y2=1.59
cc_902 ( N_GND_c_263_p N_noxref_56_c_11970_n ) capacitor c=0.00180612f \
 //x=71.98 //y=0 //x2=68.815 //y2=1.59
cc_903 ( N_GND_M42_noxref_d N_noxref_56_c_11970_n ) capacitor c=0.00853078f \
 //x=68.225 //y=0.875 //x2=68.815 //y2=1.59
cc_904 ( N_GND_c_89_p N_noxref_56_c_11974_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=68.9 //y2=0.625
cc_905 ( N_GND_c_263_p N_noxref_56_c_11974_n ) capacitor c=0.0140928f \
 //x=71.98 //y=0 //x2=68.9 //y2=0.625
cc_906 ( N_GND_M42_noxref_d N_noxref_56_c_11974_n ) capacitor c=0.033954f \
 //x=68.225 //y=0.875 //x2=68.9 //y2=0.625
cc_907 ( N_GND_c_89_p N_noxref_56_c_11977_n ) capacitor c=0.0104506f //x=95.83 \
 //y=0 //x2=69.785 //y2=0.54
cc_908 ( N_GND_c_263_p N_noxref_56_c_11977_n ) capacitor c=0.0360726f \
 //x=71.98 //y=0 //x2=69.785 //y2=0.54
cc_909 ( N_GND_c_89_p N_noxref_56_M42_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=67.795 //y2=0.375
cc_910 ( N_GND_c_256_p N_noxref_56_M42_noxref_s ) capacitor c=0.0140928f \
 //x=68.33 //y=0 //x2=67.795 //y2=0.375
cc_911 ( N_GND_c_263_p N_noxref_56_M42_noxref_s ) capacitor c=0.0131437f \
 //x=71.98 //y=0 //x2=67.795 //y2=0.375
cc_912 ( N_GND_c_16_p N_noxref_56_M42_noxref_s ) capacitor c=0.0696963f \
 //x=67.34 //y=0 //x2=67.795 //y2=0.375
cc_913 ( N_GND_c_17_p N_noxref_56_M42_noxref_s ) capacitor c=3.31601e-19 \
 //x=72.15 //y=0 //x2=67.795 //y2=0.375
cc_914 ( N_GND_M42_noxref_d N_noxref_56_M42_noxref_s ) capacitor c=0.033718f \
 //x=68.225 //y=0.875 //x2=67.795 //y2=0.375
cc_915 ( N_GND_c_89_p N_noxref_57_c_12019_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=70.355 //y2=0.995
cc_916 ( N_GND_c_263_p N_noxref_57_c_12019_n ) capacitor c=0.00934524f \
 //x=71.98 //y=0 //x2=70.355 //y2=0.995
cc_917 ( N_GND_c_89_p N_noxref_57_c_12021_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=70.44 //y2=0.625
cc_918 ( N_GND_c_263_p N_noxref_57_c_12021_n ) capacitor c=0.0140928f \
 //x=71.98 //y=0 //x2=70.44 //y2=0.625
cc_919 ( N_GND_M42_noxref_d N_noxref_57_c_12021_n ) capacitor c=6.21394e-19 \
 //x=68.225 //y=0.875 //x2=70.44 //y2=0.625
cc_920 ( N_GND_c_89_p N_noxref_57_c_12024_n ) capacitor c=0.0105317f //x=95.83 \
 //y=0 //x2=71.325 //y2=0.54
cc_921 ( N_GND_c_263_p N_noxref_57_c_12024_n ) capacitor c=0.0364215f \
 //x=71.98 //y=0 //x2=71.325 //y2=0.54
cc_922 ( N_GND_c_89_p N_noxref_57_c_12026_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=71.41 //y2=0.625
cc_923 ( N_GND_c_263_p N_noxref_57_c_12026_n ) capacitor c=0.0140304f \
 //x=71.98 //y=0 //x2=71.41 //y2=0.625
cc_924 ( N_GND_c_17_p N_noxref_57_c_12026_n ) capacitor c=0.0404137f //x=72.15 \
 //y=0 //x2=71.41 //y2=0.625
cc_925 ( N_GND_M42_noxref_d N_noxref_57_M43_noxref_d ) capacitor c=0.00162435f \
 //x=68.225 //y=0.875 //x2=69.2 //y2=0.91
cc_926 ( N_GND_c_16_p N_noxref_57_M44_noxref_s ) capacitor c=8.16352e-19 \
 //x=67.34 //y=0 //x2=70.305 //y2=0.375
cc_927 ( N_GND_c_17_p N_noxref_57_M44_noxref_s ) capacitor c=0.00183204f \
 //x=72.15 //y=0 //x2=70.305 //y2=0.375
cc_928 ( N_GND_c_89_p N_noxref_58_c_12071_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=73.625 //y2=1.59
cc_929 ( N_GND_c_272_p N_noxref_58_c_12071_n ) capacitor c=0.00111448f \
 //x=73.14 //y=0 //x2=73.625 //y2=1.59
cc_930 ( N_GND_c_279_p N_noxref_58_c_12071_n ) capacitor c=0.00180612f \
 //x=76.79 //y=0 //x2=73.625 //y2=1.59
cc_931 ( N_GND_M45_noxref_d N_noxref_58_c_12071_n ) capacitor c=0.00853078f \
 //x=73.035 //y=0.875 //x2=73.625 //y2=1.59
cc_932 ( N_GND_c_89_p N_noxref_58_c_12075_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=73.71 //y2=0.625
cc_933 ( N_GND_c_279_p N_noxref_58_c_12075_n ) capacitor c=0.0140928f \
 //x=76.79 //y=0 //x2=73.71 //y2=0.625
cc_934 ( N_GND_M45_noxref_d N_noxref_58_c_12075_n ) capacitor c=0.033954f \
 //x=73.035 //y=0.875 //x2=73.71 //y2=0.625
cc_935 ( N_GND_c_89_p N_noxref_58_c_12078_n ) capacitor c=0.0104506f //x=95.83 \
 //y=0 //x2=74.595 //y2=0.54
cc_936 ( N_GND_c_279_p N_noxref_58_c_12078_n ) capacitor c=0.0360726f \
 //x=76.79 //y=0 //x2=74.595 //y2=0.54
cc_937 ( N_GND_c_89_p N_noxref_58_M45_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=72.605 //y2=0.375
cc_938 ( N_GND_c_272_p N_noxref_58_M45_noxref_s ) capacitor c=0.0140928f \
 //x=73.14 //y=0 //x2=72.605 //y2=0.375
cc_939 ( N_GND_c_279_p N_noxref_58_M45_noxref_s ) capacitor c=0.0131437f \
 //x=76.79 //y=0 //x2=72.605 //y2=0.375
cc_940 ( N_GND_c_17_p N_noxref_58_M45_noxref_s ) capacitor c=0.0696963f \
 //x=72.15 //y=0 //x2=72.605 //y2=0.375
cc_941 ( N_GND_c_18_p N_noxref_58_M45_noxref_s ) capacitor c=3.31601e-19 \
 //x=76.96 //y=0 //x2=72.605 //y2=0.375
cc_942 ( N_GND_M45_noxref_d N_noxref_58_M45_noxref_s ) capacitor c=0.033718f \
 //x=73.035 //y=0.875 //x2=72.605 //y2=0.375
cc_943 ( N_GND_c_89_p N_noxref_59_c_12120_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=75.165 //y2=0.995
cc_944 ( N_GND_c_279_p N_noxref_59_c_12120_n ) capacitor c=0.00934524f \
 //x=76.79 //y=0 //x2=75.165 //y2=0.995
cc_945 ( N_GND_c_89_p N_noxref_59_c_12122_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=75.25 //y2=0.625
cc_946 ( N_GND_c_279_p N_noxref_59_c_12122_n ) capacitor c=0.0140928f \
 //x=76.79 //y=0 //x2=75.25 //y2=0.625
cc_947 ( N_GND_M45_noxref_d N_noxref_59_c_12122_n ) capacitor c=6.21394e-19 \
 //x=73.035 //y=0.875 //x2=75.25 //y2=0.625
cc_948 ( N_GND_c_89_p N_noxref_59_c_12125_n ) capacitor c=0.0105197f //x=95.83 \
 //y=0 //x2=76.135 //y2=0.54
cc_949 ( N_GND_c_279_p N_noxref_59_c_12125_n ) capacitor c=0.0364139f \
 //x=76.79 //y=0 //x2=76.135 //y2=0.54
cc_950 ( N_GND_c_89_p N_noxref_59_c_12127_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=76.22 //y2=0.625
cc_951 ( N_GND_c_279_p N_noxref_59_c_12127_n ) capacitor c=0.0140304f \
 //x=76.79 //y=0 //x2=76.22 //y2=0.625
cc_952 ( N_GND_c_18_p N_noxref_59_c_12127_n ) capacitor c=0.0404137f //x=76.96 \
 //y=0 //x2=76.22 //y2=0.625
cc_953 ( N_GND_M45_noxref_d N_noxref_59_M46_noxref_d ) capacitor c=0.00162435f \
 //x=73.035 //y=0.875 //x2=74.01 //y2=0.91
cc_954 ( N_GND_c_17_p N_noxref_59_M47_noxref_s ) capacitor c=8.16352e-19 \
 //x=72.15 //y=0 //x2=75.115 //y2=0.375
cc_955 ( N_GND_c_18_p N_noxref_59_M47_noxref_s ) capacitor c=0.00183204f \
 //x=76.96 //y=0 //x2=75.115 //y2=0.375
cc_956 ( N_GND_c_89_p N_noxref_60_c_12173_n ) capacitor c=0.00517576f \
 //x=95.83 //y=0 //x2=78.435 //y2=1.59
cc_957 ( N_GND_c_292_p N_noxref_60_c_12173_n ) capacitor c=0.00111448f \
 //x=77.95 //y=0 //x2=78.435 //y2=1.59
cc_958 ( N_GND_c_299_p N_noxref_60_c_12173_n ) capacitor c=0.00180612f \
 //x=81.6 //y=0 //x2=78.435 //y2=1.59
cc_959 ( N_GND_M48_noxref_d N_noxref_60_c_12173_n ) capacitor c=0.00853078f \
 //x=77.845 //y=0.875 //x2=78.435 //y2=1.59
cc_960 ( N_GND_c_89_p N_noxref_60_c_12177_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=78.52 //y2=0.625
cc_961 ( N_GND_c_299_p N_noxref_60_c_12177_n ) capacitor c=0.0140928f //x=81.6 \
 //y=0 //x2=78.52 //y2=0.625
cc_962 ( N_GND_M48_noxref_d N_noxref_60_c_12177_n ) capacitor c=0.033954f \
 //x=77.845 //y=0.875 //x2=78.52 //y2=0.625
cc_963 ( N_GND_c_89_p N_noxref_60_c_12180_n ) capacitor c=0.0105304f //x=95.83 \
 //y=0 //x2=79.405 //y2=0.54
cc_964 ( N_GND_c_299_p N_noxref_60_c_12180_n ) capacitor c=0.0361183f //x=81.6 \
 //y=0 //x2=79.405 //y2=0.54
cc_965 ( N_GND_c_89_p N_noxref_60_M48_noxref_s ) capacitor c=0.00531539f \
 //x=95.83 //y=0 //x2=77.415 //y2=0.375
cc_966 ( N_GND_c_292_p N_noxref_60_M48_noxref_s ) capacitor c=0.0140928f \
 //x=77.95 //y=0 //x2=77.415 //y2=0.375
cc_967 ( N_GND_c_299_p N_noxref_60_M48_noxref_s ) capacitor c=0.0133155f \
 //x=81.6 //y=0 //x2=77.415 //y2=0.375
cc_968 ( N_GND_c_18_p N_noxref_60_M48_noxref_s ) capacitor c=0.0696963f \
 //x=76.96 //y=0 //x2=77.415 //y2=0.375
cc_969 ( N_GND_c_19_p N_noxref_60_M48_noxref_s ) capacitor c=3.31601e-19 \
 //x=81.77 //y=0 //x2=77.415 //y2=0.375
cc_970 ( N_GND_M48_noxref_d N_noxref_60_M48_noxref_s ) capacitor c=0.033718f \
 //x=77.845 //y=0.875 //x2=77.415 //y2=0.375
cc_971 ( N_GND_c_89_p N_noxref_61_c_12224_n ) capacitor c=0.00375441f \
 //x=95.83 //y=0 //x2=79.975 //y2=0.995
cc_972 ( N_GND_c_299_p N_noxref_61_c_12224_n ) capacitor c=0.00944862f \
 //x=81.6 //y=0 //x2=79.975 //y2=0.995
cc_973 ( N_GND_c_89_p N_noxref_61_c_12226_n ) capacitor c=0.00277579f \
 //x=95.83 //y=0 //x2=80.06 //y2=0.625
cc_974 ( N_GND_c_299_p N_noxref_61_c_12226_n ) capacitor c=0.0142586f //x=81.6 \
 //y=0 //x2=80.06 //y2=0.625
cc_975 ( N_GND_M48_noxref_d N_noxref_61_c_12226_n ) capacitor c=6.21394e-19 \
 //x=77.845 //y=0.875 //x2=80.06 //y2=0.625
cc_976 ( N_GND_c_89_p N_noxref_61_c_12229_n ) capacitor c=0.010965f //x=95.83 \
 //y=0 //x2=80.945 //y2=0.54
cc_977 ( N_GND_c_299_p N_noxref_61_c_12229_n ) capacitor c=0.0363907f //x=81.6 \
 //y=0 //x2=80.945 //y2=0.54
cc_978 ( N_GND_c_89_p N_noxref_61_c_12231_n ) capacitor c=0.00253183f \
 //x=95.83 //y=0 //x2=81.03 //y2=0.625
cc_979 ( N_GND_c_299_p N_noxref_61_c_12231_n ) capacitor c=0.0140226f //x=81.6 \
 //y=0 //x2=81.03 //y2=0.625
cc_980 ( N_GND_c_19_p N_noxref_61_c_12231_n ) capacitor c=0.0404137f //x=81.77 \
 //y=0 //x2=81.03 //y2=0.625
cc_981 ( N_GND_M48_noxref_d N_noxref_61_M49_noxref_d ) capacitor c=0.00162435f \
 //x=77.845 //y=0.875 //x2=78.82 //y2=0.91
cc_982 ( N_GND_c_18_p N_noxref_61_M50_noxref_s ) capacitor c=8.16352e-19 \
 //x=76.96 //y=0 //x2=79.925 //y2=0.375
cc_983 ( N_GND_c_19_p N_noxref_61_M50_noxref_s ) capacitor c=0.00183204f \
 //x=81.77 //y=0 //x2=79.925 //y2=0.375
cc_984 ( N_GND_c_89_p N_noxref_62_c_12278_n ) capacitor c=0.00517235f \
 //x=95.83 //y=0 //x2=83.245 //y2=1.59
cc_985 ( N_GND_c_416_p N_noxref_62_c_12278_n ) capacitor c=0.00111448f \
 //x=82.76 //y=0 //x2=83.245 //y2=1.59
cc_986 ( N_GND_c_422_p N_noxref_62_c_12278_n ) capacitor c=0.00180612f \
 //x=86.41 //y=0 //x2=83.245 //y2=1.59
cc_987 ( N_GND_M51_noxref_d N_noxref_62_c_12278_n ) capacitor c=0.00851489f \
 //x=82.655 //y=0.875 //x2=83.245 //y2=1.59
cc_988 ( N_GND_c_89_p N_noxref_62_c_12282_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=83.33 //y2=0.625
cc_989 ( N_GND_c_422_p N_noxref_62_c_12282_n ) capacitor c=0.0140928f \
 //x=86.41 //y=0 //x2=83.33 //y2=0.625
cc_990 ( N_GND_M51_noxref_d N_noxref_62_c_12282_n ) capacitor c=0.033954f \
 //x=82.655 //y=0.875 //x2=83.33 //y2=0.625
cc_991 ( N_GND_c_89_p N_noxref_62_c_12285_n ) capacitor c=0.0104506f //x=95.83 \
 //y=0 //x2=84.215 //y2=0.54
cc_992 ( N_GND_c_422_p N_noxref_62_c_12285_n ) capacitor c=0.0360726f \
 //x=86.41 //y=0 //x2=84.215 //y2=0.54
cc_993 ( N_GND_c_89_p N_noxref_62_M51_noxref_s ) capacitor c=0.00507657f \
 //x=95.83 //y=0 //x2=82.225 //y2=0.375
cc_994 ( N_GND_c_416_p N_noxref_62_M51_noxref_s ) capacitor c=0.0140928f \
 //x=82.76 //y=0 //x2=82.225 //y2=0.375
cc_995 ( N_GND_c_422_p N_noxref_62_M51_noxref_s ) capacitor c=0.0136651f \
 //x=86.41 //y=0 //x2=82.225 //y2=0.375
cc_996 ( N_GND_c_19_p N_noxref_62_M51_noxref_s ) capacitor c=0.0696963f \
 //x=81.77 //y=0 //x2=82.225 //y2=0.375
cc_997 ( N_GND_c_20_p N_noxref_62_M51_noxref_s ) capacitor c=3.31601e-19 \
 //x=86.58 //y=0 //x2=82.225 //y2=0.375
cc_998 ( N_GND_M51_noxref_d N_noxref_62_M51_noxref_s ) capacitor c=0.033718f \
 //x=82.655 //y=0.875 //x2=82.225 //y2=0.375
cc_999 ( N_GND_c_89_p N_noxref_63_c_12329_n ) capacitor c=0.00352952f \
 //x=95.83 //y=0 //x2=84.785 //y2=0.995
cc_1000 ( N_GND_c_422_p N_noxref_63_c_12329_n ) capacitor c=0.00934524f \
 //x=86.41 //y=0 //x2=84.785 //y2=0.995
cc_1001 ( N_GND_c_89_p N_noxref_63_c_12331_n ) capacitor c=0.00254475f \
 //x=95.83 //y=0 //x2=84.87 //y2=0.625
cc_1002 ( N_GND_c_422_p N_noxref_63_c_12331_n ) capacitor c=0.0140928f \
 //x=86.41 //y=0 //x2=84.87 //y2=0.625
cc_1003 ( N_GND_M51_noxref_d N_noxref_63_c_12331_n ) capacitor c=6.21394e-19 \
 //x=82.655 //y=0.875 //x2=84.87 //y2=0.625
cc_1004 ( N_GND_c_89_p N_noxref_63_c_12334_n ) capacitor c=0.0105317f \
 //x=95.83 //y=0 //x2=85.755 //y2=0.54
cc_1005 ( N_GND_c_422_p N_noxref_63_c_12334_n ) capacitor c=0.0364215f \
 //x=86.41 //y=0 //x2=85.755 //y2=0.54
cc_1006 ( N_GND_c_89_p N_noxref_63_c_12336_n ) capacitor c=0.00254232f \
 //x=95.83 //y=0 //x2=85.84 //y2=0.625
cc_1007 ( N_GND_c_422_p N_noxref_63_c_12336_n ) capacitor c=0.0140304f \
 //x=86.41 //y=0 //x2=85.84 //y2=0.625
cc_1008 ( N_GND_c_20_p N_noxref_63_c_12336_n ) capacitor c=0.0400472f \
 //x=86.58 //y=0 //x2=85.84 //y2=0.625
cc_1009 ( N_GND_M51_noxref_d N_noxref_63_M52_noxref_d ) capacitor \
 c=0.00162435f //x=82.655 //y=0.875 //x2=83.63 //y2=0.91
cc_1010 ( N_GND_c_19_p N_noxref_63_M53_noxref_s ) capacitor c=8.16352e-19 \
 //x=81.77 //y=0 //x2=84.735 //y2=0.375
cc_1011 ( N_GND_c_20_p N_noxref_63_M53_noxref_s ) capacitor c=0.00183576f \
 //x=86.58 //y=0 //x2=84.735 //y2=0.375
cc_1012 ( N_GND_c_89_p N_noxref_64_c_12381_n ) capacitor c=0.00521624f \
 //x=95.83 //y=0 //x2=88.16 //y2=1.58
cc_1013 ( N_GND_c_104_p N_noxref_64_c_12381_n ) capacitor c=0.00112872f \
 //x=87.675 //y=0 //x2=88.16 //y2=1.58
cc_1014 ( N_GND_c_111_p N_noxref_64_c_12381_n ) capacitor c=0.0018229f \
 //x=89.74 //y=0 //x2=88.16 //y2=1.58
cc_1015 ( N_GND_M54_noxref_d N_noxref_64_c_12381_n ) capacitor c=0.00892401f \
 //x=87.57 //y=0.865 //x2=88.16 //y2=1.58
cc_1016 ( N_GND_c_89_p N_noxref_64_c_12385_n ) capacitor c=0.00259029f \
 //x=95.83 //y=0 //x2=88.245 //y2=0.615
cc_1017 ( N_GND_c_111_p N_noxref_64_c_12385_n ) capacitor c=0.0146901f \
 //x=89.74 //y=0 //x2=88.245 //y2=0.615
cc_1018 ( N_GND_M54_noxref_d N_noxref_64_c_12385_n ) capacitor c=0.0336822f \
 //x=87.57 //y=0.865 //x2=88.245 //y2=0.615
cc_1019 ( N_GND_c_20_p N_noxref_64_c_12388_n ) capacitor c=2.91423e-19 \
 //x=86.58 //y=0 //x2=88.245 //y2=1.495
cc_1020 ( N_GND_c_89_p N_noxref_64_c_12389_n ) capacitor c=0.00942819f \
 //x=95.83 //y=0 //x2=89.13 //y2=0.53
cc_1021 ( N_GND_c_111_p N_noxref_64_c_12389_n ) capacitor c=0.0374778f \
 //x=89.74 //y=0 //x2=89.13 //y2=0.53
cc_1022 ( N_GND_c_89_p N_noxref_64_c_12391_n ) capacitor c=0.00212661f \
 //x=95.83 //y=0 //x2=89.215 //y2=0.615
cc_1023 ( N_GND_c_111_p N_noxref_64_c_12391_n ) capacitor c=0.0143168f \
 //x=89.74 //y=0 //x2=89.215 //y2=0.615
cc_1024 ( N_GND_c_21_p N_noxref_64_c_12391_n ) capacitor c=0.0554337f \
 //x=89.91 //y=0 //x2=89.215 //y2=0.615
cc_1025 ( N_GND_c_89_p N_noxref_64_M54_noxref_s ) capacitor c=0.00259029f \
 //x=95.83 //y=0 //x2=87.14 //y2=0.365
cc_1026 ( N_GND_c_104_p N_noxref_64_M54_noxref_s ) capacitor c=0.0146901f \
 //x=87.675 //y=0 //x2=87.14 //y2=0.365
cc_1027 ( N_GND_c_20_p N_noxref_64_M54_noxref_s ) capacitor c=0.058813f \
 //x=86.58 //y=0 //x2=87.14 //y2=0.365
cc_1028 ( N_GND_c_21_p N_noxref_64_M54_noxref_s ) capacitor c=0.00181744f \
 //x=89.91 //y=0 //x2=87.14 //y2=0.365
cc_1029 ( N_GND_M54_noxref_d N_noxref_64_M54_noxref_s ) capacitor c=0.0333456f \
 //x=87.57 //y=0.865 //x2=87.14 //y2=0.365
cc_1030 ( N_GND_c_114_p N_noxref_65_c_12438_n ) capacitor c=8.01905e-19 \
 //x=91.005 //y=0 //x2=91.49 //y2=1.58
cc_1031 ( N_GND_c_120_p N_noxref_65_c_12438_n ) capacitor c=0.00161527f \
 //x=93.07 //y=0 //x2=91.49 //y2=1.58
cc_1032 ( N_GND_M56_noxref_d N_noxref_65_c_12438_n ) capacitor c=0.0073276f \
 //x=90.9 //y=0.865 //x2=91.49 //y2=1.58
cc_1033 ( N_GND_c_89_p N_noxref_65_c_12441_n ) capacitor c=0.00212661f \
 //x=95.83 //y=0 //x2=91.575 //y2=0.615
cc_1034 ( N_GND_c_120_p N_noxref_65_c_12441_n ) capacitor c=0.0143168f \
 //x=93.07 //y=0 //x2=91.575 //y2=0.615
cc_1035 ( N_GND_M56_noxref_d N_noxref_65_c_12441_n ) capacitor c=0.0336587f \
 //x=90.9 //y=0.865 //x2=91.575 //y2=0.615
cc_1036 ( N_GND_c_21_p N_noxref_65_c_12444_n ) capacitor c=2.91423e-19 \
 //x=89.91 //y=0 //x2=91.575 //y2=1.495
cc_1037 ( N_GND_c_89_p N_noxref_65_c_12445_n ) capacitor c=0.00884129f \
 //x=95.83 //y=0 //x2=92.46 //y2=0.53
cc_1038 ( N_GND_c_120_p N_noxref_65_c_12445_n ) capacitor c=0.0373651f \
 //x=93.07 //y=0 //x2=92.46 //y2=0.53
cc_1039 ( N_GND_c_89_p N_noxref_65_c_12447_n ) capacitor c=0.00212661f \
 //x=95.83 //y=0 //x2=92.545 //y2=0.615
cc_1040 ( N_GND_c_120_p N_noxref_65_c_12447_n ) capacitor c=0.0143168f \
 //x=93.07 //y=0 //x2=92.545 //y2=0.615
cc_1041 ( N_GND_c_22_p N_noxref_65_c_12447_n ) capacitor c=0.0548042f \
 //x=93.24 //y=0 //x2=92.545 //y2=0.615
cc_1042 ( N_GND_c_89_p N_noxref_65_M56_noxref_s ) capacitor c=0.00212661f \
 //x=95.83 //y=0 //x2=90.47 //y2=0.365
cc_1043 ( N_GND_c_114_p N_noxref_65_M56_noxref_s ) capacitor c=0.0143168f \
 //x=91.005 //y=0 //x2=90.47 //y2=0.365
cc_1044 ( N_GND_c_21_p N_noxref_65_M56_noxref_s ) capacitor c=0.0561194f \
 //x=89.91 //y=0 //x2=90.47 //y2=0.365
cc_1045 ( N_GND_c_22_p N_noxref_65_M56_noxref_s ) capacitor c=0.0022128f \
 //x=93.24 //y=0 //x2=90.47 //y2=0.365
cc_1046 ( N_GND_M56_noxref_d N_noxref_65_M56_noxref_s ) capacitor c=0.0332904f \
 //x=90.9 //y=0.865 //x2=90.47 //y2=0.365
cc_1047 ( N_GND_c_448_p N_noxref_66_c_12493_n ) capacitor c=8.01912e-19 \
 //x=94.335 //y=0 //x2=94.82 //y2=1.58
cc_1048 ( N_GND_c_2_p N_noxref_66_c_12493_n ) capacitor c=0.00161527f \
 //x=95.83 //y=0 //x2=94.82 //y2=1.58
cc_1049 ( N_GND_M58_noxref_d N_noxref_66_c_12493_n ) capacitor c=0.0073482f \
 //x=94.23 //y=0.865 //x2=94.82 //y2=1.58
cc_1050 ( N_GND_c_89_p N_noxref_66_c_12496_n ) capacitor c=0.00212661f \
 //x=95.83 //y=0 //x2=94.905 //y2=0.615
cc_1051 ( N_GND_c_2_p N_noxref_66_c_12496_n ) capacitor c=0.0143168f //x=95.83 \
 //y=0 //x2=94.905 //y2=0.615
cc_1052 ( N_GND_M58_noxref_d N_noxref_66_c_12496_n ) capacitor c=0.0336587f \
 //x=94.23 //y=0.865 //x2=94.905 //y2=0.615
cc_1053 ( N_GND_c_22_p N_noxref_66_c_12499_n ) capacitor c=2.91423e-19 \
 //x=93.24 //y=0 //x2=94.905 //y2=1.495
cc_1054 ( N_GND_c_89_p N_noxref_66_c_12500_n ) capacitor c=0.0119802f \
 //x=95.83 //y=0 //x2=95.79 //y2=0.53
cc_1055 ( N_GND_c_2_p N_noxref_66_c_12500_n ) capacitor c=0.0371788f //x=95.83 \
 //y=0 //x2=95.79 //y2=0.53
cc_1056 ( N_GND_c_89_p N_noxref_66_c_12502_n ) capacitor c=0.00579412f \
 //x=95.83 //y=0 //x2=95.875 //y2=0.615
cc_1057 ( N_GND_c_2_p N_noxref_66_c_12502_n ) capacitor c=0.0581858f //x=95.83 \
 //y=0 //x2=95.875 //y2=0.615
cc_1058 ( N_GND_c_89_p N_noxref_66_M58_noxref_s ) capacitor c=0.00212661f \
 //x=95.83 //y=0 //x2=93.8 //y2=0.365
cc_1059 ( N_GND_c_448_p N_noxref_66_M58_noxref_s ) capacitor c=0.0143168f \
 //x=94.335 //y=0 //x2=93.8 //y2=0.365
cc_1060 ( N_GND_c_2_p N_noxref_66_M58_noxref_s ) capacitor c=0.00202267f \
 //x=95.83 //y=0 //x2=93.8 //y2=0.365
cc_1061 ( N_GND_c_22_p N_noxref_66_M58_noxref_s ) capacitor c=0.0555228f \
 //x=93.24 //y=0 //x2=93.8 //y2=0.365
cc_1062 ( N_GND_M58_noxref_d N_noxref_66_M58_noxref_s ) capacitor c=0.0332904f \
 //x=94.23 //y=0.865 //x2=93.8 //y2=0.365
cc_1063 ( N_VDD_c_1085_p N_noxref_3_c_2250_n ) capacitor c=0.004515f //x=95.83 \
 //y=7.4 //x2=2.325 //y2=5.155
cc_1064 ( N_VDD_c_1086_p N_noxref_3_c_2250_n ) capacitor c=4.32228e-19 \
 //x=1.885 //y=7.4 //x2=2.325 //y2=5.155
cc_1065 ( N_VDD_c_1087_p N_noxref_3_c_2250_n ) capacitor c=4.32228e-19 \
 //x=2.765 //y=7.4 //x2=2.325 //y2=5.155
cc_1066 ( N_VDD_M61_noxref_d N_noxref_3_c_2250_n ) capacitor c=0.0115147f \
 //x=1.825 //y=5.02 //x2=2.325 //y2=5.155
cc_1067 ( N_VDD_c_1063_n N_noxref_3_c_2254_n ) capacitor c=0.00880189f \
 //x=0.74 //y=7.4 //x2=1.615 //y2=5.155
cc_1068 ( N_VDD_M60_noxref_s N_noxref_3_c_2254_n ) capacitor c=0.0831083f \
 //x=0.955 //y=5.02 //x2=1.615 //y2=5.155
cc_1069 ( N_VDD_c_1085_p N_noxref_3_c_2256_n ) capacitor c=0.00448996f \
 //x=95.83 //y=7.4 //x2=3.205 //y2=5.155
cc_1070 ( N_VDD_c_1087_p N_noxref_3_c_2256_n ) capacitor c=4.32228e-19 \
 //x=2.765 //y=7.4 //x2=3.205 //y2=5.155
cc_1071 ( N_VDD_c_1093_p N_noxref_3_c_2256_n ) capacitor c=4.32228e-19 \
 //x=3.645 //y=7.4 //x2=3.205 //y2=5.155
cc_1072 ( N_VDD_M63_noxref_d N_noxref_3_c_2256_n ) capacitor c=0.0115147f \
 //x=2.705 //y=5.02 //x2=3.205 //y2=5.155
cc_1073 ( N_VDD_c_1085_p N_noxref_3_c_2260_n ) capacitor c=0.00442621f \
 //x=95.83 //y=7.4 //x2=3.985 //y2=5.155
cc_1074 ( N_VDD_c_1093_p N_noxref_3_c_2260_n ) capacitor c=7.47666e-19 \
 //x=3.645 //y=7.4 //x2=3.985 //y2=5.155
cc_1075 ( N_VDD_c_1097_p N_noxref_3_c_2260_n ) capacitor c=0.00198981f \
 //x=4.64 //y=7.4 //x2=3.985 //y2=5.155
cc_1076 ( N_VDD_M65_noxref_d N_noxref_3_c_2260_n ) capacitor c=0.0115147f \
 //x=3.585 //y=5.02 //x2=3.985 //y2=5.155
cc_1077 ( N_VDD_c_1065_n N_noxref_3_c_2226_n ) capacitor c=0.0450638f //x=4.81 \
 //y=7.4 //x2=4.07 //y2=2.59
cc_1078 ( N_VDD_c_1085_p N_noxref_3_c_2227_n ) capacitor c=9.23542e-19 \
 //x=95.83 //y=7.4 //x2=5.92 //y2=2.08
cc_1079 ( N_VDD_c_1065_n N_noxref_3_c_2227_n ) capacitor c=0.015772f //x=4.81 \
 //y=7.4 //x2=5.92 //y2=2.08
cc_1080 ( N_VDD_M66_noxref_s N_noxref_3_c_2227_n ) capacitor c=0.0123142f \
 //x=5.765 //y=5.02 //x2=5.92 //y2=2.08
cc_1081 ( N_VDD_c_1085_p N_noxref_3_c_2228_n ) capacitor c=9.10347e-19 \
 //x=95.83 //y=7.4 //x2=10.73 //y2=2.08
cc_1082 ( N_VDD_c_1066_n N_noxref_3_c_2228_n ) capacitor c=0.0134711f //x=9.62 \
 //y=7.4 //x2=10.73 //y2=2.08
cc_1083 ( N_VDD_M72_noxref_s N_noxref_3_c_2228_n ) capacitor c=0.0125322f \
 //x=10.575 //y=5.02 //x2=10.73 //y2=2.08
cc_1084 ( N_VDD_c_1106_p N_noxref_3_M66_noxref_g ) capacitor c=0.00749687f \
 //x=6.695 //y=7.4 //x2=6.12 //y2=6.02
cc_1085 ( N_VDD_M66_noxref_s N_noxref_3_M66_noxref_g ) capacitor c=0.0477201f \
 //x=5.765 //y=5.02 //x2=6.12 //y2=6.02
cc_1086 ( N_VDD_c_1106_p N_noxref_3_M67_noxref_g ) capacitor c=0.00675175f \
 //x=6.695 //y=7.4 //x2=6.56 //y2=6.02
cc_1087 ( N_VDD_M67_noxref_d N_noxref_3_M67_noxref_g ) capacitor c=0.015318f \
 //x=6.635 //y=5.02 //x2=6.56 //y2=6.02
cc_1088 ( N_VDD_c_1110_p N_noxref_3_M72_noxref_g ) capacitor c=0.00749687f \
 //x=11.505 //y=7.4 //x2=10.93 //y2=6.02
cc_1089 ( N_VDD_M72_noxref_s N_noxref_3_M72_noxref_g ) capacitor c=0.0477201f \
 //x=10.575 //y=5.02 //x2=10.93 //y2=6.02
cc_1090 ( N_VDD_c_1110_p N_noxref_3_M73_noxref_g ) capacitor c=0.00675175f \
 //x=11.505 //y=7.4 //x2=11.37 //y2=6.02
cc_1091 ( N_VDD_M73_noxref_d N_noxref_3_M73_noxref_g ) capacitor c=0.015318f \
 //x=11.445 //y=5.02 //x2=11.37 //y2=6.02
cc_1092 ( N_VDD_c_1065_n N_noxref_3_c_2279_n ) capacitor c=0.00757682f \
 //x=4.81 //y=7.4 //x2=6.195 //y2=4.79
cc_1093 ( N_VDD_M66_noxref_s N_noxref_3_c_2279_n ) capacitor c=0.00445134f \
 //x=5.765 //y=5.02 //x2=6.195 //y2=4.79
cc_1094 ( N_VDD_c_1066_n N_noxref_3_c_2281_n ) capacitor c=0.00757682f \
 //x=9.62 //y=7.4 //x2=11.005 //y2=4.79
cc_1095 ( N_VDD_M72_noxref_s N_noxref_3_c_2281_n ) capacitor c=0.00444914f \
 //x=10.575 //y=5.02 //x2=11.005 //y2=4.79
cc_1096 ( N_VDD_c_1085_p N_noxref_3_M60_noxref_d ) capacitor c=0.00285091f \
 //x=95.83 //y=7.4 //x2=1.385 //y2=5.02
cc_1097 ( N_VDD_c_1086_p N_noxref_3_M60_noxref_d ) capacitor c=0.0141016f \
 //x=1.885 //y=7.4 //x2=1.385 //y2=5.02
cc_1098 ( N_VDD_M61_noxref_d N_noxref_3_M60_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=1.385 //y2=5.02
cc_1099 ( N_VDD_c_1085_p N_noxref_3_M62_noxref_d ) capacitor c=0.00285091f \
 //x=95.83 //y=7.4 //x2=2.265 //y2=5.02
cc_1100 ( N_VDD_c_1087_p N_noxref_3_M62_noxref_d ) capacitor c=0.0141016f \
 //x=2.765 //y=7.4 //x2=2.265 //y2=5.02
cc_1101 ( N_VDD_c_1065_n N_noxref_3_M62_noxref_d ) capacitor c=4.9285e-19 \
 //x=4.81 //y=7.4 //x2=2.265 //y2=5.02
cc_1102 ( N_VDD_M60_noxref_s N_noxref_3_M62_noxref_d ) capacitor c=0.00130656f \
 //x=0.955 //y=5.02 //x2=2.265 //y2=5.02
cc_1103 ( N_VDD_M61_noxref_d N_noxref_3_M62_noxref_d ) capacitor c=0.0664752f \
 //x=1.825 //y=5.02 //x2=2.265 //y2=5.02
cc_1104 ( N_VDD_M63_noxref_d N_noxref_3_M62_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=2.265 //y2=5.02
cc_1105 ( N_VDD_c_1085_p N_noxref_3_M64_noxref_d ) capacitor c=0.00285091f \
 //x=95.83 //y=7.4 //x2=3.145 //y2=5.02
cc_1106 ( N_VDD_c_1093_p N_noxref_3_M64_noxref_d ) capacitor c=0.0141016f \
 //x=3.645 //y=7.4 //x2=3.145 //y2=5.02
cc_1107 ( N_VDD_c_1065_n N_noxref_3_M64_noxref_d ) capacitor c=0.00939849f \
 //x=4.81 //y=7.4 //x2=3.145 //y2=5.02
cc_1108 ( N_VDD_M63_noxref_d N_noxref_3_M64_noxref_d ) capacitor c=0.0664752f \
 //x=2.705 //y=5.02 //x2=3.145 //y2=5.02
cc_1109 ( N_VDD_M65_noxref_d N_noxref_3_M64_noxref_d ) capacitor c=0.0664752f \
 //x=3.585 //y=5.02 //x2=3.145 //y2=5.02
cc_1110 ( N_VDD_M66_noxref_s N_noxref_3_M64_noxref_d ) capacitor c=3.57641e-19 \
 //x=5.765 //y=5.02 //x2=3.145 //y2=5.02
cc_1111 ( N_VDD_c_1085_p N_noxref_4_c_2477_n ) capacitor c=0.00444892f \
 //x=95.83 //y=7.4 //x2=11.945 //y2=5.155
cc_1112 ( N_VDD_c_1110_p N_noxref_4_c_2477_n ) capacitor c=4.31931e-19 \
 //x=11.505 //y=7.4 //x2=11.945 //y2=5.155
cc_1113 ( N_VDD_c_1135_p N_noxref_4_c_2477_n ) capacitor c=4.31931e-19 \
 //x=12.385 //y=7.4 //x2=11.945 //y2=5.155
cc_1114 ( N_VDD_M73_noxref_d N_noxref_4_c_2477_n ) capacitor c=0.0112985f \
 //x=11.445 //y=5.02 //x2=11.945 //y2=5.155
cc_1115 ( N_VDD_c_1066_n N_noxref_4_c_2481_n ) capacitor c=0.00863585f \
 //x=9.62 //y=7.4 //x2=11.235 //y2=5.155
cc_1116 ( N_VDD_M72_noxref_s N_noxref_4_c_2481_n ) capacitor c=0.0831083f \
 //x=10.575 //y=5.02 //x2=11.235 //y2=5.155
cc_1117 ( N_VDD_c_1085_p N_noxref_4_c_2483_n ) capacitor c=0.0044221f \
 //x=95.83 //y=7.4 //x2=12.825 //y2=5.155
cc_1118 ( N_VDD_c_1135_p N_noxref_4_c_2483_n ) capacitor c=4.31931e-19 \
 //x=12.385 //y=7.4 //x2=12.825 //y2=5.155
cc_1119 ( N_VDD_c_1141_p N_noxref_4_c_2483_n ) capacitor c=4.31931e-19 \
 //x=13.265 //y=7.4 //x2=12.825 //y2=5.155
cc_1120 ( N_VDD_M75_noxref_d N_noxref_4_c_2483_n ) capacitor c=0.0112985f \
 //x=12.325 //y=5.02 //x2=12.825 //y2=5.155
cc_1121 ( N_VDD_c_1085_p N_noxref_4_c_2487_n ) capacitor c=0.00434174f \
 //x=95.83 //y=7.4 //x2=13.605 //y2=5.155
cc_1122 ( N_VDD_c_1141_p N_noxref_4_c_2487_n ) capacitor c=7.46626e-19 \
 //x=13.265 //y=7.4 //x2=13.605 //y2=5.155
cc_1123 ( N_VDD_c_1145_p N_noxref_4_c_2487_n ) capacitor c=0.00198565f \
 //x=14.26 //y=7.4 //x2=13.605 //y2=5.155
cc_1124 ( N_VDD_M77_noxref_d N_noxref_4_c_2487_n ) capacitor c=0.0112985f \
 //x=13.205 //y=5.02 //x2=13.605 //y2=5.155
cc_1125 ( N_VDD_c_1067_n N_noxref_4_c_2464_n ) capacitor c=0.0427199f \
 //x=14.43 //y=7.4 //x2=13.69 //y2=2.59
cc_1126 ( N_VDD_c_1085_p N_noxref_4_c_2465_n ) capacitor c=9.10347e-19 \
 //x=95.83 //y=7.4 //x2=15.54 //y2=2.08
cc_1127 ( N_VDD_c_1067_n N_noxref_4_c_2465_n ) capacitor c=0.0134112f \
 //x=14.43 //y=7.4 //x2=15.54 //y2=2.08
cc_1128 ( N_VDD_M78_noxref_s N_noxref_4_c_2465_n ) capacitor c=0.0126798f \
 //x=15.385 //y=5.02 //x2=15.54 //y2=2.08
cc_1129 ( N_VDD_c_1151_p N_noxref_4_M78_noxref_g ) capacitor c=0.00749687f \
 //x=16.315 //y=7.4 //x2=15.74 //y2=6.02
cc_1130 ( N_VDD_M78_noxref_s N_noxref_4_M78_noxref_g ) capacitor c=0.0477201f \
 //x=15.385 //y=5.02 //x2=15.74 //y2=6.02
cc_1131 ( N_VDD_c_1151_p N_noxref_4_M79_noxref_g ) capacitor c=0.00675175f \
 //x=16.315 //y=7.4 //x2=16.18 //y2=6.02
cc_1132 ( N_VDD_M79_noxref_d N_noxref_4_M79_noxref_g ) capacitor c=0.015318f \
 //x=16.255 //y=5.02 //x2=16.18 //y2=6.02
cc_1133 ( N_VDD_c_1067_n N_noxref_4_c_2499_n ) capacitor c=0.00757682f \
 //x=14.43 //y=7.4 //x2=15.815 //y2=4.79
cc_1134 ( N_VDD_M78_noxref_s N_noxref_4_c_2499_n ) capacitor c=0.00444914f \
 //x=15.385 //y=5.02 //x2=15.815 //y2=4.79
cc_1135 ( N_VDD_c_1085_p N_noxref_4_M72_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=11.005 //y2=5.02
cc_1136 ( N_VDD_c_1110_p N_noxref_4_M72_noxref_d ) capacitor c=0.014035f \
 //x=11.505 //y=7.4 //x2=11.005 //y2=5.02
cc_1137 ( N_VDD_M73_noxref_d N_noxref_4_M72_noxref_d ) capacitor c=0.0664752f \
 //x=11.445 //y=5.02 //x2=11.005 //y2=5.02
cc_1138 ( N_VDD_c_1085_p N_noxref_4_M74_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=11.885 //y2=5.02
cc_1139 ( N_VDD_c_1135_p N_noxref_4_M74_noxref_d ) capacitor c=0.014035f \
 //x=12.385 //y=7.4 //x2=11.885 //y2=5.02
cc_1140 ( N_VDD_c_1067_n N_noxref_4_M74_noxref_d ) capacitor c=4.9285e-19 \
 //x=14.43 //y=7.4 //x2=11.885 //y2=5.02
cc_1141 ( N_VDD_M72_noxref_s N_noxref_4_M74_noxref_d ) capacitor c=0.00130656f \
 //x=10.575 //y=5.02 //x2=11.885 //y2=5.02
cc_1142 ( N_VDD_M73_noxref_d N_noxref_4_M74_noxref_d ) capacitor c=0.0664752f \
 //x=11.445 //y=5.02 //x2=11.885 //y2=5.02
cc_1143 ( N_VDD_M75_noxref_d N_noxref_4_M74_noxref_d ) capacitor c=0.0664752f \
 //x=12.325 //y=5.02 //x2=11.885 //y2=5.02
cc_1144 ( N_VDD_c_1085_p N_noxref_4_M76_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=12.765 //y2=5.02
cc_1145 ( N_VDD_c_1141_p N_noxref_4_M76_noxref_d ) capacitor c=0.014035f \
 //x=13.265 //y=7.4 //x2=12.765 //y2=5.02
cc_1146 ( N_VDD_c_1067_n N_noxref_4_M76_noxref_d ) capacitor c=0.00939849f \
 //x=14.43 //y=7.4 //x2=12.765 //y2=5.02
cc_1147 ( N_VDD_M75_noxref_d N_noxref_4_M76_noxref_d ) capacitor c=0.0664752f \
 //x=12.325 //y=5.02 //x2=12.765 //y2=5.02
cc_1148 ( N_VDD_M77_noxref_d N_noxref_4_M76_noxref_d ) capacitor c=0.0664752f \
 //x=13.205 //y=5.02 //x2=12.765 //y2=5.02
cc_1149 ( N_VDD_M78_noxref_s N_noxref_4_M76_noxref_d ) capacitor c=3.57641e-19 \
 //x=15.385 //y=5.02 //x2=12.765 //y2=5.02
cc_1150 ( N_VDD_c_1065_n N_noxref_5_c_2628_n ) capacitor c=8.16879e-19 \
 //x=4.81 //y=7.4 //x2=3.33 //y2=2.08
cc_1151 ( N_VDD_c_1085_p N_noxref_5_c_2643_n ) capacitor c=0.00449316f \
 //x=95.83 //y=7.4 //x2=7.135 //y2=5.155
cc_1152 ( N_VDD_c_1106_p N_noxref_5_c_2643_n ) capacitor c=4.32228e-19 \
 //x=6.695 //y=7.4 //x2=7.135 //y2=5.155
cc_1153 ( N_VDD_c_1175_p N_noxref_5_c_2643_n ) capacitor c=4.31906e-19 \
 //x=7.575 //y=7.4 //x2=7.135 //y2=5.155
cc_1154 ( N_VDD_M67_noxref_d N_noxref_5_c_2643_n ) capacitor c=0.0115147f \
 //x=6.635 //y=5.02 //x2=7.135 //y2=5.155
cc_1155 ( N_VDD_c_1065_n N_noxref_5_c_2647_n ) capacitor c=0.00863585f \
 //x=4.81 //y=7.4 //x2=6.425 //y2=5.155
cc_1156 ( N_VDD_M66_noxref_s N_noxref_5_c_2647_n ) capacitor c=0.0831083f \
 //x=5.765 //y=5.02 //x2=6.425 //y2=5.155
cc_1157 ( N_VDD_c_1085_p N_noxref_5_c_2649_n ) capacitor c=0.0044221f \
 //x=95.83 //y=7.4 //x2=8.015 //y2=5.155
cc_1158 ( N_VDD_c_1175_p N_noxref_5_c_2649_n ) capacitor c=4.31931e-19 \
 //x=7.575 //y=7.4 //x2=8.015 //y2=5.155
cc_1159 ( N_VDD_c_1181_p N_noxref_5_c_2649_n ) capacitor c=4.31931e-19 \
 //x=8.455 //y=7.4 //x2=8.015 //y2=5.155
cc_1160 ( N_VDD_M69_noxref_d N_noxref_5_c_2649_n ) capacitor c=0.0112985f \
 //x=7.515 //y=5.02 //x2=8.015 //y2=5.155
cc_1161 ( N_VDD_c_1085_p N_noxref_5_c_2653_n ) capacitor c=0.00434174f \
 //x=95.83 //y=7.4 //x2=8.795 //y2=5.155
cc_1162 ( N_VDD_c_1181_p N_noxref_5_c_2653_n ) capacitor c=7.46626e-19 \
 //x=8.455 //y=7.4 //x2=8.795 //y2=5.155
cc_1163 ( N_VDD_c_1185_p N_noxref_5_c_2653_n ) capacitor c=0.00198565f \
 //x=9.45 //y=7.4 //x2=8.795 //y2=5.155
cc_1164 ( N_VDD_M71_noxref_d N_noxref_5_c_2653_n ) capacitor c=0.0112985f \
 //x=8.395 //y=5.02 //x2=8.795 //y2=5.155
cc_1165 ( N_VDD_c_1066_n N_noxref_5_c_2657_n ) capacitor c=0.0427116f //x=9.62 \
 //y=7.4 //x2=8.88 //y2=3.33
cc_1166 ( N_VDD_c_1085_p N_noxref_5_c_2630_n ) capacitor c=9.10347e-19 \
 //x=95.83 //y=7.4 //x2=20.35 //y2=2.08
cc_1167 ( N_VDD_c_1068_n N_noxref_5_c_2630_n ) capacitor c=0.0134711f \
 //x=19.24 //y=7.4 //x2=20.35 //y2=2.08
cc_1168 ( N_VDD_M84_noxref_s N_noxref_5_c_2630_n ) capacitor c=0.0125322f \
 //x=20.195 //y=5.02 //x2=20.35 //y2=2.08
cc_1169 ( N_VDD_c_1093_p N_noxref_5_M64_noxref_g ) capacitor c=0.00675175f \
 //x=3.645 //y=7.4 //x2=3.07 //y2=6.02
cc_1170 ( N_VDD_M63_noxref_d N_noxref_5_M64_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=3.07 //y2=6.02
cc_1171 ( N_VDD_c_1093_p N_noxref_5_M65_noxref_g ) capacitor c=0.00675379f \
 //x=3.645 //y=7.4 //x2=3.51 //y2=6.02
cc_1172 ( N_VDD_M65_noxref_d N_noxref_5_M65_noxref_g ) capacitor c=0.0394719f \
 //x=3.585 //y=5.02 //x2=3.51 //y2=6.02
cc_1173 ( N_VDD_c_1195_p N_noxref_5_M84_noxref_g ) capacitor c=0.00749687f \
 //x=21.125 //y=7.4 //x2=20.55 //y2=6.02
cc_1174 ( N_VDD_M84_noxref_s N_noxref_5_M84_noxref_g ) capacitor c=0.0477201f \
 //x=20.195 //y=5.02 //x2=20.55 //y2=6.02
cc_1175 ( N_VDD_c_1195_p N_noxref_5_M85_noxref_g ) capacitor c=0.00675175f \
 //x=21.125 //y=7.4 //x2=20.99 //y2=6.02
cc_1176 ( N_VDD_M85_noxref_d N_noxref_5_M85_noxref_g ) capacitor c=0.015318f \
 //x=21.065 //y=5.02 //x2=20.99 //y2=6.02
cc_1177 ( N_VDD_c_1068_n N_noxref_5_c_2669_n ) capacitor c=0.00757682f \
 //x=19.24 //y=7.4 //x2=20.625 //y2=4.79
cc_1178 ( N_VDD_M84_noxref_s N_noxref_5_c_2669_n ) capacitor c=0.00444914f \
 //x=20.195 //y=5.02 //x2=20.625 //y2=4.79
cc_1179 ( N_VDD_c_1085_p N_noxref_5_M66_noxref_d ) capacitor c=0.00285091f \
 //x=95.83 //y=7.4 //x2=6.195 //y2=5.02
cc_1180 ( N_VDD_c_1106_p N_noxref_5_M66_noxref_d ) capacitor c=0.0141016f \
 //x=6.695 //y=7.4 //x2=6.195 //y2=5.02
cc_1181 ( N_VDD_M67_noxref_d N_noxref_5_M66_noxref_d ) capacitor c=0.0664752f \
 //x=6.635 //y=5.02 //x2=6.195 //y2=5.02
cc_1182 ( N_VDD_c_1085_p N_noxref_5_M68_noxref_d ) capacitor c=0.00275186f \
 //x=95.83 //y=7.4 //x2=7.075 //y2=5.02
cc_1183 ( N_VDD_c_1175_p N_noxref_5_M68_noxref_d ) capacitor c=0.0140346f \
 //x=7.575 //y=7.4 //x2=7.075 //y2=5.02
cc_1184 ( N_VDD_c_1066_n N_noxref_5_M68_noxref_d ) capacitor c=4.9285e-19 \
 //x=9.62 //y=7.4 //x2=7.075 //y2=5.02
cc_1185 ( N_VDD_M66_noxref_s N_noxref_5_M68_noxref_d ) capacitor c=0.00130656f \
 //x=5.765 //y=5.02 //x2=7.075 //y2=5.02
cc_1186 ( N_VDD_M67_noxref_d N_noxref_5_M68_noxref_d ) capacitor c=0.0664752f \
 //x=6.635 //y=5.02 //x2=7.075 //y2=5.02
cc_1187 ( N_VDD_M69_noxref_d N_noxref_5_M68_noxref_d ) capacitor c=0.0664752f \
 //x=7.515 //y=5.02 //x2=7.075 //y2=5.02
cc_1188 ( N_VDD_c_1085_p N_noxref_5_M70_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=7.955 //y2=5.02
cc_1189 ( N_VDD_c_1181_p N_noxref_5_M70_noxref_d ) capacitor c=0.014035f \
 //x=8.455 //y=7.4 //x2=7.955 //y2=5.02
cc_1190 ( N_VDD_c_1066_n N_noxref_5_M70_noxref_d ) capacitor c=0.00939849f \
 //x=9.62 //y=7.4 //x2=7.955 //y2=5.02
cc_1191 ( N_VDD_M69_noxref_d N_noxref_5_M70_noxref_d ) capacitor c=0.0664752f \
 //x=7.515 //y=5.02 //x2=7.955 //y2=5.02
cc_1192 ( N_VDD_M71_noxref_d N_noxref_5_M70_noxref_d ) capacitor c=0.0664752f \
 //x=8.395 //y=5.02 //x2=7.955 //y2=5.02
cc_1193 ( N_VDD_M72_noxref_s N_noxref_5_M70_noxref_d ) capacitor c=3.57641e-19 \
 //x=10.575 //y=5.02 //x2=7.955 //y2=5.02
cc_1194 ( N_VDD_c_1085_p N_noxref_6_c_2934_n ) capacitor c=0.42938f //x=95.83 \
 //y=7.4 //x2=75.025 //y2=4.81
cc_1195 ( N_VDD_c_1217_p N_noxref_6_c_2934_n ) capacitor c=0.00238461f \
 //x=23.88 //y=7.4 //x2=75.025 //y2=4.81
cc_1196 ( N_VDD_c_1218_p N_noxref_6_c_2934_n ) capacitor c=0.00393349f \
 //x=25.055 //y=7.4 //x2=75.025 //y2=4.81
cc_1197 ( N_VDD_c_1219_p N_noxref_6_c_2934_n ) capacitor c=0.00257486f \
 //x=25.935 //y=7.4 //x2=75.025 //y2=4.81
cc_1198 ( N_VDD_c_1220_p N_noxref_6_c_2934_n ) capacitor c=0.00309625f \
 //x=28.69 //y=7.4 //x2=75.025 //y2=4.81
cc_1199 ( N_VDD_c_1221_p N_noxref_6_c_2934_n ) capacitor c=0.00393349f \
 //x=29.865 //y=7.4 //x2=75.025 //y2=4.81
cc_1200 ( N_VDD_c_1222_p N_noxref_6_c_2934_n ) capacitor c=0.00257486f \
 //x=30.745 //y=7.4 //x2=75.025 //y2=4.81
cc_1201 ( N_VDD_c_1223_p N_noxref_6_c_2934_n ) capacitor c=0.00309625f \
 //x=33.5 //y=7.4 //x2=75.025 //y2=4.81
cc_1202 ( N_VDD_c_1224_p N_noxref_6_c_2934_n ) capacitor c=0.00393349f \
 //x=34.675 //y=7.4 //x2=75.025 //y2=4.81
cc_1203 ( N_VDD_c_1225_p N_noxref_6_c_2934_n ) capacitor c=0.00257486f \
 //x=35.555 //y=7.4 //x2=75.025 //y2=4.81
cc_1204 ( N_VDD_c_1226_p N_noxref_6_c_2934_n ) capacitor c=0.00309625f \
 //x=38.31 //y=7.4 //x2=75.025 //y2=4.81
cc_1205 ( N_VDD_c_1227_p N_noxref_6_c_2934_n ) capacitor c=0.00393349f \
 //x=39.485 //y=7.4 //x2=75.025 //y2=4.81
cc_1206 ( N_VDD_c_1228_p N_noxref_6_c_2934_n ) capacitor c=0.00257486f \
 //x=40.365 //y=7.4 //x2=75.025 //y2=4.81
cc_1207 ( N_VDD_c_1229_p N_noxref_6_c_2934_n ) capacitor c=0.00309625f \
 //x=43.12 //y=7.4 //x2=75.025 //y2=4.81
cc_1208 ( N_VDD_c_1230_p N_noxref_6_c_2934_n ) capacitor c=0.00393349f \
 //x=44.295 //y=7.4 //x2=75.025 //y2=4.81
cc_1209 ( N_VDD_c_1231_p N_noxref_6_c_2934_n ) capacitor c=0.00257486f \
 //x=45.175 //y=7.4 //x2=75.025 //y2=4.81
cc_1210 ( N_VDD_c_1232_p N_noxref_6_c_2934_n ) capacitor c=0.00309625f \
 //x=47.93 //y=7.4 //x2=75.025 //y2=4.81
cc_1211 ( N_VDD_c_1233_p N_noxref_6_c_2934_n ) capacitor c=0.00393349f \
 //x=49.105 //y=7.4 //x2=75.025 //y2=4.81
cc_1212 ( N_VDD_c_1234_p N_noxref_6_c_2934_n ) capacitor c=0.00257486f \
 //x=49.985 //y=7.4 //x2=75.025 //y2=4.81
cc_1213 ( N_VDD_c_1235_p N_noxref_6_c_2934_n ) capacitor c=0.00309625f \
 //x=52.74 //y=7.4 //x2=75.025 //y2=4.81
cc_1214 ( N_VDD_c_1236_p N_noxref_6_c_2934_n ) capacitor c=0.00393349f \
 //x=53.915 //y=7.4 //x2=75.025 //y2=4.81
cc_1215 ( N_VDD_c_1237_p N_noxref_6_c_2934_n ) capacitor c=0.00257486f \
 //x=54.795 //y=7.4 //x2=75.025 //y2=4.81
cc_1216 ( N_VDD_c_1238_p N_noxref_6_c_2934_n ) capacitor c=0.00309625f \
 //x=57.55 //y=7.4 //x2=75.025 //y2=4.81
cc_1217 ( N_VDD_c_1239_p N_noxref_6_c_2934_n ) capacitor c=0.00393349f \
 //x=58.725 //y=7.4 //x2=75.025 //y2=4.81
cc_1218 ( N_VDD_c_1240_p N_noxref_6_c_2934_n ) capacitor c=0.00257486f \
 //x=59.605 //y=7.4 //x2=75.025 //y2=4.81
cc_1219 ( N_VDD_c_1241_p N_noxref_6_c_2934_n ) capacitor c=0.00309625f \
 //x=62.36 //y=7.4 //x2=75.025 //y2=4.81
cc_1220 ( N_VDD_c_1242_p N_noxref_6_c_2934_n ) capacitor c=0.00393349f \
 //x=63.535 //y=7.4 //x2=75.025 //y2=4.81
cc_1221 ( N_VDD_c_1243_p N_noxref_6_c_2934_n ) capacitor c=0.00257486f \
 //x=64.415 //y=7.4 //x2=75.025 //y2=4.81
cc_1222 ( N_VDD_c_1244_p N_noxref_6_c_2934_n ) capacitor c=0.00309625f \
 //x=67.17 //y=7.4 //x2=75.025 //y2=4.81
cc_1223 ( N_VDD_c_1245_p N_noxref_6_c_2934_n ) capacitor c=0.00393349f \
 //x=68.345 //y=7.4 //x2=75.025 //y2=4.81
cc_1224 ( N_VDD_c_1246_p N_noxref_6_c_2934_n ) capacitor c=0.00257486f \
 //x=69.225 //y=7.4 //x2=75.025 //y2=4.81
cc_1225 ( N_VDD_c_1247_p N_noxref_6_c_2934_n ) capacitor c=0.00309625f \
 //x=71.98 //y=7.4 //x2=75.025 //y2=4.81
cc_1226 ( N_VDD_c_1248_p N_noxref_6_c_2934_n ) capacitor c=0.00393349f \
 //x=73.155 //y=7.4 //x2=75.025 //y2=4.81
cc_1227 ( N_VDD_c_1249_p N_noxref_6_c_2934_n ) capacitor c=0.00257486f \
 //x=74.035 //y=7.4 //x2=75.025 //y2=4.81
cc_1228 ( N_VDD_c_1069_n N_noxref_6_c_2934_n ) capacitor c=0.0387886f \
 //x=24.05 //y=7.4 //x2=75.025 //y2=4.81
cc_1229 ( N_VDD_c_1070_n N_noxref_6_c_2934_n ) capacitor c=0.0387886f \
 //x=28.86 //y=7.4 //x2=75.025 //y2=4.81
cc_1230 ( N_VDD_c_1071_n N_noxref_6_c_2934_n ) capacitor c=0.0387886f \
 //x=33.67 //y=7.4 //x2=75.025 //y2=4.81
cc_1231 ( N_VDD_c_1072_n N_noxref_6_c_2934_n ) capacitor c=0.0387886f \
 //x=38.48 //y=7.4 //x2=75.025 //y2=4.81
cc_1232 ( N_VDD_c_1073_n N_noxref_6_c_2934_n ) capacitor c=0.0387886f \
 //x=43.29 //y=7.4 //x2=75.025 //y2=4.81
cc_1233 ( N_VDD_c_1074_n N_noxref_6_c_2934_n ) capacitor c=0.0387886f //x=48.1 \
 //y=7.4 //x2=75.025 //y2=4.81
cc_1234 ( N_VDD_c_1075_n N_noxref_6_c_2934_n ) capacitor c=0.0387886f \
 //x=52.91 //y=7.4 //x2=75.025 //y2=4.81
cc_1235 ( N_VDD_c_1076_n N_noxref_6_c_2934_n ) capacitor c=0.0387886f \
 //x=57.72 //y=7.4 //x2=75.025 //y2=4.81
cc_1236 ( N_VDD_c_1077_n N_noxref_6_c_2934_n ) capacitor c=0.0387886f \
 //x=62.53 //y=7.4 //x2=75.025 //y2=4.81
cc_1237 ( N_VDD_c_1078_n N_noxref_6_c_2934_n ) capacitor c=0.0387886f \
 //x=67.34 //y=7.4 //x2=75.025 //y2=4.81
cc_1238 ( N_VDD_c_1079_n N_noxref_6_c_2934_n ) capacitor c=0.0387869f \
 //x=72.15 //y=7.4 //x2=75.025 //y2=4.81
cc_1239 ( N_VDD_M90_noxref_s N_noxref_6_c_2934_n ) capacitor c=0.00433388f \
 //x=25.005 //y=5.02 //x2=75.025 //y2=4.81
cc_1240 ( N_VDD_M96_noxref_s N_noxref_6_c_2934_n ) capacitor c=0.00433388f \
 //x=29.815 //y=5.02 //x2=75.025 //y2=4.81
cc_1241 ( N_VDD_M102_noxref_s N_noxref_6_c_2934_n ) capacitor c=0.00433388f \
 //x=34.625 //y=5.02 //x2=75.025 //y2=4.81
cc_1242 ( N_VDD_M108_noxref_s N_noxref_6_c_2934_n ) capacitor c=0.00433388f \
 //x=39.435 //y=5.02 //x2=75.025 //y2=4.81
cc_1243 ( N_VDD_M114_noxref_s N_noxref_6_c_2934_n ) capacitor c=0.00433388f \
 //x=44.245 //y=5.02 //x2=75.025 //y2=4.81
cc_1244 ( N_VDD_M120_noxref_s N_noxref_6_c_2934_n ) capacitor c=0.00433388f \
 //x=49.055 //y=5.02 //x2=75.025 //y2=4.81
cc_1245 ( N_VDD_M126_noxref_s N_noxref_6_c_2934_n ) capacitor c=0.00433388f \
 //x=53.865 //y=5.02 //x2=75.025 //y2=4.81
cc_1246 ( N_VDD_M132_noxref_s N_noxref_6_c_2934_n ) capacitor c=0.00433388f \
 //x=58.675 //y=5.02 //x2=75.025 //y2=4.81
cc_1247 ( N_VDD_M138_noxref_s N_noxref_6_c_2934_n ) capacitor c=0.00433388f \
 //x=63.485 //y=5.02 //x2=75.025 //y2=4.81
cc_1248 ( N_VDD_M144_noxref_s N_noxref_6_c_2934_n ) capacitor c=0.00433388f \
 //x=68.295 //y=5.02 //x2=75.025 //y2=4.81
cc_1249 ( N_VDD_M150_noxref_s N_noxref_6_c_2934_n ) capacitor c=0.00433388f \
 //x=73.105 //y=5.02 //x2=75.025 //y2=4.81
cc_1250 ( N_VDD_c_1085_p N_noxref_6_c_2990_n ) capacitor c=0.00247397f \
 //x=95.83 //y=7.4 //x2=23.425 //y2=4.81
cc_1251 ( N_VDD_c_1217_p N_noxref_6_c_2990_n ) capacitor c=7.12616e-19 \
 //x=23.88 //y=7.4 //x2=23.425 //y2=4.81
cc_1252 ( N_VDD_c_1069_n N_noxref_6_c_2990_n ) capacitor c=0.00190934f \
 //x=24.05 //y=7.4 //x2=23.425 //y2=4.81
cc_1253 ( N_VDD_c_1085_p N_noxref_6_c_2993_n ) capacitor c=0.0898237f \
 //x=95.83 //y=7.4 //x2=87.205 //y2=4.44
cc_1254 ( N_VDD_c_1276_p N_noxref_6_c_2993_n ) capacitor c=0.00258496f \
 //x=76.79 //y=7.4 //x2=87.205 //y2=4.44
cc_1255 ( N_VDD_c_1277_p N_noxref_6_c_2993_n ) capacitor c=0.00328994f \
 //x=77.965 //y=7.4 //x2=87.205 //y2=4.44
cc_1256 ( N_VDD_c_1278_p N_noxref_6_c_2993_n ) capacitor c=0.00135925f \
 //x=78.845 //y=7.4 //x2=87.205 //y2=4.44
cc_1257 ( N_VDD_c_1279_p N_noxref_6_c_2993_n ) capacitor c=0.00258496f \
 //x=81.6 //y=7.4 //x2=87.205 //y2=4.44
cc_1258 ( N_VDD_c_1280_p N_noxref_6_c_2993_n ) capacitor c=0.00328994f \
 //x=82.775 //y=7.4 //x2=87.205 //y2=4.44
cc_1259 ( N_VDD_c_1281_p N_noxref_6_c_2993_n ) capacitor c=0.00135925f \
 //x=83.655 //y=7.4 //x2=87.205 //y2=4.44
cc_1260 ( N_VDD_c_1282_p N_noxref_6_c_2993_n ) capacitor c=0.00258496f \
 //x=86.41 //y=7.4 //x2=87.205 //y2=4.44
cc_1261 ( N_VDD_c_1283_p N_noxref_6_c_2993_n ) capacitor c=0.00196539f \
 //x=87.285 //y=7.4 //x2=87.205 //y2=4.44
cc_1262 ( N_VDD_c_1080_n N_noxref_6_c_2993_n ) capacitor c=0.0389825f \
 //x=76.96 //y=7.4 //x2=87.205 //y2=4.44
cc_1263 ( N_VDD_c_1081_n N_noxref_6_c_2993_n ) capacitor c=0.0389825f \
 //x=81.77 //y=7.4 //x2=87.205 //y2=4.44
cc_1264 ( N_VDD_c_1082_n N_noxref_6_c_2993_n ) capacitor c=0.0377357f \
 //x=86.58 //y=7.4 //x2=87.205 //y2=4.44
cc_1265 ( N_VDD_M156_noxref_s N_noxref_6_c_2993_n ) capacitor c=0.00179496f \
 //x=77.915 //y=5.02 //x2=87.205 //y2=4.44
cc_1266 ( N_VDD_M162_noxref_s N_noxref_6_c_2993_n ) capacitor c=0.00179496f \
 //x=82.725 //y=5.02 //x2=87.205 //y2=4.44
cc_1267 ( N_VDD_c_1085_p N_noxref_6_c_3007_n ) capacitor c=0.014626f //x=95.83 \
 //y=7.4 //x2=90.905 //y2=4.44
cc_1268 ( N_VDD_c_1290_p N_noxref_6_c_3007_n ) capacitor c=0.00134165f \
 //x=88.165 //y=7.4 //x2=90.905 //y2=4.44
cc_1269 ( N_VDD_c_1083_n N_noxref_6_c_3007_n ) capacitor c=0.03415f //x=89.91 \
 //y=7.4 //x2=90.905 //y2=4.44
cc_1270 ( N_VDD_M168_noxref_s N_noxref_6_c_3007_n ) capacitor c=6.29527e-19 \
 //x=87.235 //y=5.025 //x2=90.905 //y2=4.44
cc_1271 ( N_VDD_M171_noxref_d N_noxref_6_c_3007_n ) capacitor c=0.0033086f \
 //x=88.985 //y=5.025 //x2=90.905 //y2=4.44
cc_1272 ( N_VDD_c_1085_p N_noxref_6_c_3012_n ) capacitor c=0.00140297f \
 //x=95.83 //y=7.4 //x2=87.435 //y2=4.44
cc_1273 ( N_VDD_c_1283_p N_noxref_6_c_3012_n ) capacitor c=3.1987e-19 \
 //x=87.285 //y=7.4 //x2=87.435 //y2=4.44
cc_1274 ( N_VDD_c_1082_n N_noxref_6_c_3012_n ) capacitor c=0.00205902f \
 //x=86.58 //y=7.4 //x2=87.435 //y2=4.44
cc_1275 ( N_VDD_M168_noxref_s N_noxref_6_c_3012_n ) capacitor c=0.00225389f \
 //x=87.235 //y=5.025 //x2=87.435 //y2=4.44
cc_1276 ( N_VDD_c_1085_p N_noxref_6_c_3016_n ) capacitor c=0.00444892f \
 //x=95.83 //y=7.4 //x2=21.565 //y2=5.155
cc_1277 ( N_VDD_c_1195_p N_noxref_6_c_3016_n ) capacitor c=4.31931e-19 \
 //x=21.125 //y=7.4 //x2=21.565 //y2=5.155
cc_1278 ( N_VDD_c_1300_p N_noxref_6_c_3016_n ) capacitor c=4.31931e-19 \
 //x=22.005 //y=7.4 //x2=21.565 //y2=5.155
cc_1279 ( N_VDD_M85_noxref_d N_noxref_6_c_3016_n ) capacitor c=0.0112985f \
 //x=21.065 //y=5.02 //x2=21.565 //y2=5.155
cc_1280 ( N_VDD_c_1068_n N_noxref_6_c_3020_n ) capacitor c=0.00863585f \
 //x=19.24 //y=7.4 //x2=20.855 //y2=5.155
cc_1281 ( N_VDD_M84_noxref_s N_noxref_6_c_3020_n ) capacitor c=0.0831083f \
 //x=20.195 //y=5.02 //x2=20.855 //y2=5.155
cc_1282 ( N_VDD_c_1085_p N_noxref_6_c_3022_n ) capacitor c=0.0044221f \
 //x=95.83 //y=7.4 //x2=22.445 //y2=5.155
cc_1283 ( N_VDD_c_1300_p N_noxref_6_c_3022_n ) capacitor c=4.31931e-19 \
 //x=22.005 //y=7.4 //x2=22.445 //y2=5.155
cc_1284 ( N_VDD_c_1306_p N_noxref_6_c_3022_n ) capacitor c=4.31931e-19 \
 //x=22.885 //y=7.4 //x2=22.445 //y2=5.155
cc_1285 ( N_VDD_M87_noxref_d N_noxref_6_c_3022_n ) capacitor c=0.0112985f \
 //x=21.945 //y=5.02 //x2=22.445 //y2=5.155
cc_1286 ( N_VDD_c_1085_p N_noxref_6_c_3026_n ) capacitor c=0.00431542f \
 //x=95.83 //y=7.4 //x2=23.225 //y2=5.155
cc_1287 ( N_VDD_c_1306_p N_noxref_6_c_3026_n ) capacitor c=7.46626e-19 \
 //x=22.885 //y=7.4 //x2=23.225 //y2=5.155
cc_1288 ( N_VDD_c_1217_p N_noxref_6_c_3026_n ) capacitor c=0.0019817f \
 //x=23.88 //y=7.4 //x2=23.225 //y2=5.155
cc_1289 ( N_VDD_M89_noxref_d N_noxref_6_c_3026_n ) capacitor c=0.0112985f \
 //x=22.825 //y=5.02 //x2=23.225 //y2=5.155
cc_1290 ( N_VDD_c_1069_n N_noxref_6_c_2896_n ) capacitor c=0.0400289f \
 //x=24.05 //y=7.4 //x2=23.31 //y2=2.59
cc_1291 ( N_VDD_c_1085_p N_noxref_6_c_2897_n ) capacitor c=6.51035e-19 \
 //x=95.83 //y=7.4 //x2=25.16 //y2=2.08
cc_1292 ( N_VDD_c_1069_n N_noxref_6_c_2897_n ) capacitor c=0.011472f //x=24.05 \
 //y=7.4 //x2=25.16 //y2=2.08
cc_1293 ( N_VDD_M90_noxref_s N_noxref_6_c_2897_n ) capacitor c=0.00923513f \
 //x=25.005 //y=5.02 //x2=25.16 //y2=2.08
cc_1294 ( N_VDD_c_1085_p N_noxref_6_c_2898_n ) capacitor c=0.00142825f \
 //x=95.83 //y=7.4 //x2=87.32 //y2=2.08
cc_1295 ( N_VDD_c_1082_n N_noxref_6_c_2898_n ) capacitor c=0.0239954f \
 //x=86.58 //y=7.4 //x2=87.32 //y2=2.08
cc_1296 ( N_VDD_c_1083_n N_noxref_6_c_2898_n ) capacitor c=3.70458e-19 \
 //x=89.91 //y=7.4 //x2=87.32 //y2=2.08
cc_1297 ( N_VDD_M168_noxref_s N_noxref_6_c_2898_n ) capacitor c=0.0119799f \
 //x=87.235 //y=5.025 //x2=87.32 //y2=2.08
cc_1298 ( N_VDD_c_1083_n N_noxref_6_c_2901_n ) capacitor c=0.0131686f \
 //x=89.91 //y=7.4 //x2=91.02 //y2=2.08
cc_1299 ( N_VDD_c_1084_n N_noxref_6_c_2901_n ) capacitor c=0.00133861f \
 //x=93.24 //y=7.4 //x2=91.02 //y2=2.08
cc_1300 ( N_VDD_c_1219_p N_noxref_6_M90_noxref_g ) capacitor c=0.00749687f \
 //x=25.935 //y=7.4 //x2=25.36 //y2=6.02
cc_1301 ( N_VDD_M90_noxref_s N_noxref_6_M90_noxref_g ) capacitor c=0.0477201f \
 //x=25.005 //y=5.02 //x2=25.36 //y2=6.02
cc_1302 ( N_VDD_c_1219_p N_noxref_6_M91_noxref_g ) capacitor c=0.00675175f \
 //x=25.935 //y=7.4 //x2=25.8 //y2=6.02
cc_1303 ( N_VDD_M91_noxref_d N_noxref_6_M91_noxref_g ) capacitor c=0.015318f \
 //x=25.875 //y=5.02 //x2=25.8 //y2=6.02
cc_1304 ( N_VDD_c_1290_p N_noxref_6_M168_noxref_g ) capacitor c=0.00754867f \
 //x=88.165 //y=7.4 //x2=87.59 //y2=6.025
cc_1305 ( N_VDD_c_1082_n N_noxref_6_M168_noxref_g ) capacitor c=0.00694765f \
 //x=86.58 //y=7.4 //x2=87.59 //y2=6.025
cc_1306 ( N_VDD_M168_noxref_s N_noxref_6_M168_noxref_g ) capacitor \
 c=0.0547553f //x=87.235 //y=5.025 //x2=87.59 //y2=6.025
cc_1307 ( N_VDD_c_1290_p N_noxref_6_M169_noxref_g ) capacitor c=0.00678153f \
 //x=88.165 //y=7.4 //x2=88.03 //y2=6.025
cc_1308 ( N_VDD_M169_noxref_d N_noxref_6_M169_noxref_g ) capacitor c=0.015501f \
 //x=88.105 //y=5.025 //x2=88.03 //y2=6.025
cc_1309 ( N_VDD_c_1331_p N_noxref_6_M172_noxref_g ) capacitor c=0.00513227f \
 //x=93.07 //y=7.4 //x2=90.91 //y2=6.025
cc_1310 ( N_VDD_c_1083_n N_noxref_6_M172_noxref_g ) capacitor c=0.00316281f \
 //x=89.91 //y=7.4 //x2=90.91 //y2=6.025
cc_1311 ( N_VDD_c_1331_p N_noxref_6_M173_noxref_g ) capacitor c=0.00512552f \
 //x=93.07 //y=7.4 //x2=91.35 //y2=6.025
cc_1312 ( N_VDD_c_1069_n N_noxref_6_c_3052_n ) capacitor c=0.00522674f \
 //x=24.05 //y=7.4 //x2=25.435 //y2=4.79
cc_1313 ( N_VDD_M90_noxref_s N_noxref_6_c_3052_n ) capacitor c=0.00433385f \
 //x=25.005 //y=5.02 //x2=25.435 //y2=4.79
cc_1314 ( N_VDD_c_1082_n N_noxref_6_c_3054_n ) capacitor c=0.0110236f \
 //x=86.58 //y=7.4 //x2=87.665 //y2=4.795
cc_1315 ( N_VDD_M168_noxref_s N_noxref_6_c_3054_n ) capacitor c=0.00628155f \
 //x=87.235 //y=5.025 //x2=87.665 //y2=4.795
cc_1316 ( N_VDD_c_1083_n N_noxref_6_c_3056_n ) capacitor c=0.0115029f \
 //x=89.91 //y=7.4 //x2=91.02 //y2=4.705
cc_1317 ( N_VDD_c_1085_p N_noxref_6_M84_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=20.625 //y2=5.02
cc_1318 ( N_VDD_c_1195_p N_noxref_6_M84_noxref_d ) capacitor c=0.014035f \
 //x=21.125 //y=7.4 //x2=20.625 //y2=5.02
cc_1319 ( N_VDD_M85_noxref_d N_noxref_6_M84_noxref_d ) capacitor c=0.0664752f \
 //x=21.065 //y=5.02 //x2=20.625 //y2=5.02
cc_1320 ( N_VDD_c_1085_p N_noxref_6_M86_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=21.505 //y2=5.02
cc_1321 ( N_VDD_c_1300_p N_noxref_6_M86_noxref_d ) capacitor c=0.014035f \
 //x=22.005 //y=7.4 //x2=21.505 //y2=5.02
cc_1322 ( N_VDD_c_1069_n N_noxref_6_M86_noxref_d ) capacitor c=4.9285e-19 \
 //x=24.05 //y=7.4 //x2=21.505 //y2=5.02
cc_1323 ( N_VDD_M84_noxref_s N_noxref_6_M86_noxref_d ) capacitor c=0.00130656f \
 //x=20.195 //y=5.02 //x2=21.505 //y2=5.02
cc_1324 ( N_VDD_M85_noxref_d N_noxref_6_M86_noxref_d ) capacitor c=0.0664752f \
 //x=21.065 //y=5.02 //x2=21.505 //y2=5.02
cc_1325 ( N_VDD_M87_noxref_d N_noxref_6_M86_noxref_d ) capacitor c=0.0664752f \
 //x=21.945 //y=5.02 //x2=21.505 //y2=5.02
cc_1326 ( N_VDD_c_1085_p N_noxref_6_M88_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=22.385 //y2=5.02
cc_1327 ( N_VDD_c_1306_p N_noxref_6_M88_noxref_d ) capacitor c=0.014035f \
 //x=22.885 //y=7.4 //x2=22.385 //y2=5.02
cc_1328 ( N_VDD_c_1069_n N_noxref_6_M88_noxref_d ) capacitor c=0.00939849f \
 //x=24.05 //y=7.4 //x2=22.385 //y2=5.02
cc_1329 ( N_VDD_M87_noxref_d N_noxref_6_M88_noxref_d ) capacitor c=0.0664752f \
 //x=21.945 //y=5.02 //x2=22.385 //y2=5.02
cc_1330 ( N_VDD_M89_noxref_d N_noxref_6_M88_noxref_d ) capacitor c=0.0664752f \
 //x=22.825 //y=5.02 //x2=22.385 //y2=5.02
cc_1331 ( N_VDD_M90_noxref_s N_noxref_6_M88_noxref_d ) capacitor c=3.57641e-19 \
 //x=25.005 //y=5.02 //x2=22.385 //y2=5.02
cc_1332 ( N_VDD_c_1066_n N_noxref_7_c_3527_n ) capacitor c=6.58823e-19 \
 //x=9.62 //y=7.4 //x2=8.14 //y2=2.08
cc_1333 ( N_VDD_c_1067_n N_noxref_7_c_3528_n ) capacitor c=5.72823e-19 \
 //x=14.43 //y=7.4 //x2=12.95 //y2=2.08
cc_1334 ( N_VDD_c_1085_p N_noxref_7_c_3534_n ) capacitor c=0.00444751f \
 //x=95.83 //y=7.4 //x2=16.755 //y2=5.155
cc_1335 ( N_VDD_c_1151_p N_noxref_7_c_3534_n ) capacitor c=4.31931e-19 \
 //x=16.315 //y=7.4 //x2=16.755 //y2=5.155
cc_1336 ( N_VDD_c_1358_p N_noxref_7_c_3534_n ) capacitor c=4.31906e-19 \
 //x=17.195 //y=7.4 //x2=16.755 //y2=5.155
cc_1337 ( N_VDD_M79_noxref_d N_noxref_7_c_3534_n ) capacitor c=0.0112985f \
 //x=16.255 //y=5.02 //x2=16.755 //y2=5.155
cc_1338 ( N_VDD_c_1067_n N_noxref_7_c_3538_n ) capacitor c=0.00863585f \
 //x=14.43 //y=7.4 //x2=16.045 //y2=5.155
cc_1339 ( N_VDD_M78_noxref_s N_noxref_7_c_3538_n ) capacitor c=0.0831083f \
 //x=15.385 //y=5.02 //x2=16.045 //y2=5.155
cc_1340 ( N_VDD_c_1085_p N_noxref_7_c_3540_n ) capacitor c=0.0044221f \
 //x=95.83 //y=7.4 //x2=17.635 //y2=5.155
cc_1341 ( N_VDD_c_1358_p N_noxref_7_c_3540_n ) capacitor c=4.31931e-19 \
 //x=17.195 //y=7.4 //x2=17.635 //y2=5.155
cc_1342 ( N_VDD_c_1364_p N_noxref_7_c_3540_n ) capacitor c=4.31931e-19 \
 //x=18.075 //y=7.4 //x2=17.635 //y2=5.155
cc_1343 ( N_VDD_M81_noxref_d N_noxref_7_c_3540_n ) capacitor c=0.0112985f \
 //x=17.135 //y=5.02 //x2=17.635 //y2=5.155
cc_1344 ( N_VDD_c_1085_p N_noxref_7_c_3544_n ) capacitor c=0.00434174f \
 //x=95.83 //y=7.4 //x2=18.415 //y2=5.155
cc_1345 ( N_VDD_c_1364_p N_noxref_7_c_3544_n ) capacitor c=7.46626e-19 \
 //x=18.075 //y=7.4 //x2=18.415 //y2=5.155
cc_1346 ( N_VDD_c_1368_p N_noxref_7_c_3544_n ) capacitor c=0.00198565f \
 //x=19.07 //y=7.4 //x2=18.415 //y2=5.155
cc_1347 ( N_VDD_M83_noxref_d N_noxref_7_c_3544_n ) capacitor c=0.0112985f \
 //x=18.015 //y=5.02 //x2=18.415 //y2=5.155
cc_1348 ( N_VDD_c_1068_n N_noxref_7_c_3548_n ) capacitor c=0.0427116f \
 //x=19.24 //y=7.4 //x2=18.5 //y2=3.7
cc_1349 ( N_VDD_c_1070_n N_noxref_7_c_3530_n ) capacitor c=4.93757e-19 \
 //x=28.86 //y=7.4 //x2=27.38 //y2=2.08
cc_1350 ( N_VDD_c_1181_p N_noxref_7_M70_noxref_g ) capacitor c=0.00675175f \
 //x=8.455 //y=7.4 //x2=7.88 //y2=6.02
cc_1351 ( N_VDD_M69_noxref_d N_noxref_7_M70_noxref_g ) capacitor c=0.015318f \
 //x=7.515 //y=5.02 //x2=7.88 //y2=6.02
cc_1352 ( N_VDD_c_1181_p N_noxref_7_M71_noxref_g ) capacitor c=0.00675379f \
 //x=8.455 //y=7.4 //x2=8.32 //y2=6.02
cc_1353 ( N_VDD_M71_noxref_d N_noxref_7_M71_noxref_g ) capacitor c=0.0394719f \
 //x=8.395 //y=5.02 //x2=8.32 //y2=6.02
cc_1354 ( N_VDD_c_1141_p N_noxref_7_M76_noxref_g ) capacitor c=0.00675175f \
 //x=13.265 //y=7.4 //x2=12.69 //y2=6.02
cc_1355 ( N_VDD_M75_noxref_d N_noxref_7_M76_noxref_g ) capacitor c=0.015318f \
 //x=12.325 //y=5.02 //x2=12.69 //y2=6.02
cc_1356 ( N_VDD_c_1141_p N_noxref_7_M77_noxref_g ) capacitor c=0.00675379f \
 //x=13.265 //y=7.4 //x2=13.13 //y2=6.02
cc_1357 ( N_VDD_M77_noxref_d N_noxref_7_M77_noxref_g ) capacitor c=0.0394719f \
 //x=13.205 //y=5.02 //x2=13.13 //y2=6.02
cc_1358 ( N_VDD_c_1380_p N_noxref_7_M94_noxref_g ) capacitor c=0.00675175f \
 //x=27.695 //y=7.4 //x2=27.12 //y2=6.02
cc_1359 ( N_VDD_M93_noxref_d N_noxref_7_M94_noxref_g ) capacitor c=0.015318f \
 //x=26.755 //y=5.02 //x2=27.12 //y2=6.02
cc_1360 ( N_VDD_c_1380_p N_noxref_7_M95_noxref_g ) capacitor c=0.00675379f \
 //x=27.695 //y=7.4 //x2=27.56 //y2=6.02
cc_1361 ( N_VDD_M95_noxref_d N_noxref_7_M95_noxref_g ) capacitor c=0.0394719f \
 //x=27.635 //y=5.02 //x2=27.56 //y2=6.02
cc_1362 ( N_VDD_c_1085_p N_noxref_7_M78_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=15.815 //y2=5.02
cc_1363 ( N_VDD_c_1151_p N_noxref_7_M78_noxref_d ) capacitor c=0.014035f \
 //x=16.315 //y=7.4 //x2=15.815 //y2=5.02
cc_1364 ( N_VDD_M79_noxref_d N_noxref_7_M78_noxref_d ) capacitor c=0.0664752f \
 //x=16.255 //y=5.02 //x2=15.815 //y2=5.02
cc_1365 ( N_VDD_c_1085_p N_noxref_7_M80_noxref_d ) capacitor c=0.00275186f \
 //x=95.83 //y=7.4 //x2=16.695 //y2=5.02
cc_1366 ( N_VDD_c_1358_p N_noxref_7_M80_noxref_d ) capacitor c=0.0140346f \
 //x=17.195 //y=7.4 //x2=16.695 //y2=5.02
cc_1367 ( N_VDD_c_1068_n N_noxref_7_M80_noxref_d ) capacitor c=4.9285e-19 \
 //x=19.24 //y=7.4 //x2=16.695 //y2=5.02
cc_1368 ( N_VDD_M78_noxref_s N_noxref_7_M80_noxref_d ) capacitor c=0.00130656f \
 //x=15.385 //y=5.02 //x2=16.695 //y2=5.02
cc_1369 ( N_VDD_M79_noxref_d N_noxref_7_M80_noxref_d ) capacitor c=0.0664752f \
 //x=16.255 //y=5.02 //x2=16.695 //y2=5.02
cc_1370 ( N_VDD_M81_noxref_d N_noxref_7_M80_noxref_d ) capacitor c=0.0664752f \
 //x=17.135 //y=5.02 //x2=16.695 //y2=5.02
cc_1371 ( N_VDD_c_1085_p N_noxref_7_M82_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=17.575 //y2=5.02
cc_1372 ( N_VDD_c_1364_p N_noxref_7_M82_noxref_d ) capacitor c=0.014035f \
 //x=18.075 //y=7.4 //x2=17.575 //y2=5.02
cc_1373 ( N_VDD_c_1068_n N_noxref_7_M82_noxref_d ) capacitor c=0.00939849f \
 //x=19.24 //y=7.4 //x2=17.575 //y2=5.02
cc_1374 ( N_VDD_M81_noxref_d N_noxref_7_M82_noxref_d ) capacitor c=0.0664752f \
 //x=17.135 //y=5.02 //x2=17.575 //y2=5.02
cc_1375 ( N_VDD_M83_noxref_d N_noxref_7_M82_noxref_d ) capacitor c=0.0664752f \
 //x=18.015 //y=5.02 //x2=17.575 //y2=5.02
cc_1376 ( N_VDD_M84_noxref_s N_noxref_7_M82_noxref_d ) capacitor c=3.57641e-19 \
 //x=20.195 //y=5.02 //x2=17.575 //y2=5.02
cc_1377 ( N_VDD_c_1069_n N_noxref_8_c_3866_n ) capacitor c=4.9109e-19 \
 //x=24.05 //y=7.4 //x2=22.57 //y2=2.08
cc_1378 ( N_VDD_c_1085_p N_noxref_8_c_3870_n ) capacitor c=0.00437246f \
 //x=95.83 //y=7.4 //x2=26.375 //y2=5.155
cc_1379 ( N_VDD_c_1219_p N_noxref_8_c_3870_n ) capacitor c=4.31596e-19 \
 //x=25.935 //y=7.4 //x2=26.375 //y2=5.155
cc_1380 ( N_VDD_c_1402_p N_noxref_8_c_3870_n ) capacitor c=4.31596e-19 \
 //x=26.815 //y=7.4 //x2=26.375 //y2=5.155
cc_1381 ( N_VDD_M91_noxref_d N_noxref_8_c_3870_n ) capacitor c=0.0109802f \
 //x=25.875 //y=5.02 //x2=26.375 //y2=5.155
cc_1382 ( N_VDD_c_1069_n N_noxref_8_c_3874_n ) capacitor c=0.00863585f \
 //x=24.05 //y=7.4 //x2=25.665 //y2=5.155
cc_1383 ( N_VDD_M90_noxref_s N_noxref_8_c_3874_n ) capacitor c=0.0831083f \
 //x=25.005 //y=5.02 //x2=25.665 //y2=5.155
cc_1384 ( N_VDD_c_1085_p N_noxref_8_c_3876_n ) capacitor c=0.00434259f \
 //x=95.83 //y=7.4 //x2=27.255 //y2=5.155
cc_1385 ( N_VDD_c_1402_p N_noxref_8_c_3876_n ) capacitor c=4.31596e-19 \
 //x=26.815 //y=7.4 //x2=27.255 //y2=5.155
cc_1386 ( N_VDD_c_1380_p N_noxref_8_c_3876_n ) capacitor c=4.31596e-19 \
 //x=27.695 //y=7.4 //x2=27.255 //y2=5.155
cc_1387 ( N_VDD_M93_noxref_d N_noxref_8_c_3876_n ) capacitor c=0.0109802f \
 //x=26.755 //y=5.02 //x2=27.255 //y2=5.155
cc_1388 ( N_VDD_c_1085_p N_noxref_8_c_3880_n ) capacitor c=0.00424413f \
 //x=95.83 //y=7.4 //x2=28.035 //y2=5.155
cc_1389 ( N_VDD_c_1380_p N_noxref_8_c_3880_n ) capacitor c=7.45454e-19 \
 //x=27.695 //y=7.4 //x2=28.035 //y2=5.155
cc_1390 ( N_VDD_c_1220_p N_noxref_8_c_3880_n ) capacitor c=0.00198097f \
 //x=28.69 //y=7.4 //x2=28.035 //y2=5.155
cc_1391 ( N_VDD_M95_noxref_d N_noxref_8_c_3880_n ) capacitor c=0.0109802f \
 //x=27.635 //y=5.02 //x2=28.035 //y2=5.155
cc_1392 ( N_VDD_c_1070_n N_noxref_8_c_3884_n ) capacitor c=0.0401063f \
 //x=28.86 //y=7.4 //x2=28.12 //y2=3.33
cc_1393 ( N_VDD_c_1306_p N_noxref_8_M88_noxref_g ) capacitor c=0.00675175f \
 //x=22.885 //y=7.4 //x2=22.31 //y2=6.02
cc_1394 ( N_VDD_M87_noxref_d N_noxref_8_M88_noxref_g ) capacitor c=0.015318f \
 //x=21.945 //y=5.02 //x2=22.31 //y2=6.02
cc_1395 ( N_VDD_c_1306_p N_noxref_8_M89_noxref_g ) capacitor c=0.00675379f \
 //x=22.885 //y=7.4 //x2=22.75 //y2=6.02
cc_1396 ( N_VDD_M89_noxref_d N_noxref_8_M89_noxref_g ) capacitor c=0.0394719f \
 //x=22.825 //y=5.02 //x2=22.75 //y2=6.02
cc_1397 ( N_VDD_c_1085_p N_noxref_8_M90_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=25.435 //y2=5.02
cc_1398 ( N_VDD_c_1219_p N_noxref_8_M90_noxref_d ) capacitor c=0.0139598f \
 //x=25.935 //y=7.4 //x2=25.435 //y2=5.02
cc_1399 ( N_VDD_M91_noxref_d N_noxref_8_M90_noxref_d ) capacitor c=0.0664752f \
 //x=25.875 //y=5.02 //x2=25.435 //y2=5.02
cc_1400 ( N_VDD_c_1085_p N_noxref_8_M92_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=26.315 //y2=5.02
cc_1401 ( N_VDD_c_1402_p N_noxref_8_M92_noxref_d ) capacitor c=0.0139598f \
 //x=26.815 //y=7.4 //x2=26.315 //y2=5.02
cc_1402 ( N_VDD_c_1070_n N_noxref_8_M92_noxref_d ) capacitor c=4.9285e-19 \
 //x=28.86 //y=7.4 //x2=26.315 //y2=5.02
cc_1403 ( N_VDD_M90_noxref_s N_noxref_8_M92_noxref_d ) capacitor c=0.00130656f \
 //x=25.005 //y=5.02 //x2=26.315 //y2=5.02
cc_1404 ( N_VDD_M91_noxref_d N_noxref_8_M92_noxref_d ) capacitor c=0.0664752f \
 //x=25.875 //y=5.02 //x2=26.315 //y2=5.02
cc_1405 ( N_VDD_M93_noxref_d N_noxref_8_M92_noxref_d ) capacitor c=0.0664752f \
 //x=26.755 //y=5.02 //x2=26.315 //y2=5.02
cc_1406 ( N_VDD_c_1085_p N_noxref_8_M94_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=27.195 //y2=5.02
cc_1407 ( N_VDD_c_1380_p N_noxref_8_M94_noxref_d ) capacitor c=0.0139598f \
 //x=27.695 //y=7.4 //x2=27.195 //y2=5.02
cc_1408 ( N_VDD_c_1070_n N_noxref_8_M94_noxref_d ) capacitor c=0.00939849f \
 //x=28.86 //y=7.4 //x2=27.195 //y2=5.02
cc_1409 ( N_VDD_M93_noxref_d N_noxref_8_M94_noxref_d ) capacitor c=0.0664752f \
 //x=26.755 //y=5.02 //x2=27.195 //y2=5.02
cc_1410 ( N_VDD_M95_noxref_d N_noxref_8_M94_noxref_d ) capacitor c=0.0664752f \
 //x=27.635 //y=5.02 //x2=27.195 //y2=5.02
cc_1411 ( N_VDD_M96_noxref_s N_noxref_8_M94_noxref_d ) capacitor c=3.57641e-19 \
 //x=29.815 //y=5.02 //x2=27.195 //y2=5.02
cc_1412 ( N_VDD_c_1085_p N_noxref_9_c_4071_n ) capacitor c=0.00437246f \
 //x=95.83 //y=7.4 //x2=31.185 //y2=5.155
cc_1413 ( N_VDD_c_1222_p N_noxref_9_c_4071_n ) capacitor c=4.31596e-19 \
 //x=30.745 //y=7.4 //x2=31.185 //y2=5.155
cc_1414 ( N_VDD_c_1436_p N_noxref_9_c_4071_n ) capacitor c=4.31596e-19 \
 //x=31.625 //y=7.4 //x2=31.185 //y2=5.155
cc_1415 ( N_VDD_M97_noxref_d N_noxref_9_c_4071_n ) capacitor c=0.0109802f \
 //x=30.685 //y=5.02 //x2=31.185 //y2=5.155
cc_1416 ( N_VDD_c_1070_n N_noxref_9_c_4075_n ) capacitor c=0.00863585f \
 //x=28.86 //y=7.4 //x2=30.475 //y2=5.155
cc_1417 ( N_VDD_M96_noxref_s N_noxref_9_c_4075_n ) capacitor c=0.0831083f \
 //x=29.815 //y=5.02 //x2=30.475 //y2=5.155
cc_1418 ( N_VDD_c_1085_p N_noxref_9_c_4077_n ) capacitor c=0.00434259f \
 //x=95.83 //y=7.4 //x2=32.065 //y2=5.155
cc_1419 ( N_VDD_c_1436_p N_noxref_9_c_4077_n ) capacitor c=4.31596e-19 \
 //x=31.625 //y=7.4 //x2=32.065 //y2=5.155
cc_1420 ( N_VDD_c_1442_p N_noxref_9_c_4077_n ) capacitor c=4.31596e-19 \
 //x=32.505 //y=7.4 //x2=32.065 //y2=5.155
cc_1421 ( N_VDD_M99_noxref_d N_noxref_9_c_4077_n ) capacitor c=0.0109802f \
 //x=31.565 //y=5.02 //x2=32.065 //y2=5.155
cc_1422 ( N_VDD_c_1085_p N_noxref_9_c_4081_n ) capacitor c=0.00424413f \
 //x=95.83 //y=7.4 //x2=32.845 //y2=5.155
cc_1423 ( N_VDD_c_1442_p N_noxref_9_c_4081_n ) capacitor c=7.45454e-19 \
 //x=32.505 //y=7.4 //x2=32.845 //y2=5.155
cc_1424 ( N_VDD_c_1223_p N_noxref_9_c_4081_n ) capacitor c=0.00198097f \
 //x=33.5 //y=7.4 //x2=32.845 //y2=5.155
cc_1425 ( N_VDD_M101_noxref_d N_noxref_9_c_4081_n ) capacitor c=0.0109802f \
 //x=32.445 //y=5.02 //x2=32.845 //y2=5.155
cc_1426 ( N_VDD_c_1071_n N_noxref_9_c_4047_n ) capacitor c=0.0400751f \
 //x=33.67 //y=7.4 //x2=32.93 //y2=2.59
cc_1427 ( N_VDD_c_1085_p N_noxref_9_c_4048_n ) capacitor c=6.51035e-19 \
 //x=95.83 //y=7.4 //x2=34.78 //y2=2.08
cc_1428 ( N_VDD_c_1071_n N_noxref_9_c_4048_n ) capacitor c=0.0114465f \
 //x=33.67 //y=7.4 //x2=34.78 //y2=2.08
cc_1429 ( N_VDD_M102_noxref_s N_noxref_9_c_4048_n ) capacitor c=0.00909681f \
 //x=34.625 //y=5.02 //x2=34.78 //y2=2.08
cc_1430 ( N_VDD_c_1085_p N_noxref_9_c_4049_n ) capacitor c=6.51035e-19 \
 //x=95.83 //y=7.4 //x2=39.59 //y2=2.08
cc_1431 ( N_VDD_c_1072_n N_noxref_9_c_4049_n ) capacitor c=0.0115064f \
 //x=38.48 //y=7.4 //x2=39.59 //y2=2.08
cc_1432 ( N_VDD_M108_noxref_s N_noxref_9_c_4049_n ) capacitor c=0.00923513f \
 //x=39.435 //y=5.02 //x2=39.59 //y2=2.08
cc_1433 ( N_VDD_c_1225_p N_noxref_9_M102_noxref_g ) capacitor c=0.00749687f \
 //x=35.555 //y=7.4 //x2=34.98 //y2=6.02
cc_1434 ( N_VDD_M102_noxref_s N_noxref_9_M102_noxref_g ) capacitor \
 c=0.0477201f //x=34.625 //y=5.02 //x2=34.98 //y2=6.02
cc_1435 ( N_VDD_c_1225_p N_noxref_9_M103_noxref_g ) capacitor c=0.00675175f \
 //x=35.555 //y=7.4 //x2=35.42 //y2=6.02
cc_1436 ( N_VDD_M103_noxref_d N_noxref_9_M103_noxref_g ) capacitor c=0.015318f \
 //x=35.495 //y=5.02 //x2=35.42 //y2=6.02
cc_1437 ( N_VDD_c_1228_p N_noxref_9_M108_noxref_g ) capacitor c=0.00749687f \
 //x=40.365 //y=7.4 //x2=39.79 //y2=6.02
cc_1438 ( N_VDD_M108_noxref_s N_noxref_9_M108_noxref_g ) capacitor \
 c=0.0477201f //x=39.435 //y=5.02 //x2=39.79 //y2=6.02
cc_1439 ( N_VDD_c_1228_p N_noxref_9_M109_noxref_g ) capacitor c=0.00675175f \
 //x=40.365 //y=7.4 //x2=40.23 //y2=6.02
cc_1440 ( N_VDD_M109_noxref_d N_noxref_9_M109_noxref_g ) capacitor c=0.015318f \
 //x=40.305 //y=5.02 //x2=40.23 //y2=6.02
cc_1441 ( N_VDD_c_1071_n N_noxref_9_c_4100_n ) capacitor c=0.00528488f \
 //x=33.67 //y=7.4 //x2=35.055 //y2=4.79
cc_1442 ( N_VDD_M102_noxref_s N_noxref_9_c_4100_n ) capacitor c=0.00433385f \
 //x=34.625 //y=5.02 //x2=35.055 //y2=4.79
cc_1443 ( N_VDD_c_1072_n N_noxref_9_c_4102_n ) capacitor c=0.00528488f \
 //x=38.48 //y=7.4 //x2=39.865 //y2=4.79
cc_1444 ( N_VDD_M108_noxref_s N_noxref_9_c_4102_n ) capacitor c=0.00433385f \
 //x=39.435 //y=5.02 //x2=39.865 //y2=4.79
cc_1445 ( N_VDD_c_1085_p N_noxref_9_M96_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=30.245 //y2=5.02
cc_1446 ( N_VDD_c_1222_p N_noxref_9_M96_noxref_d ) capacitor c=0.0139598f \
 //x=30.745 //y=7.4 //x2=30.245 //y2=5.02
cc_1447 ( N_VDD_M97_noxref_d N_noxref_9_M96_noxref_d ) capacitor c=0.0664752f \
 //x=30.685 //y=5.02 //x2=30.245 //y2=5.02
cc_1448 ( N_VDD_c_1085_p N_noxref_9_M98_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=31.125 //y2=5.02
cc_1449 ( N_VDD_c_1436_p N_noxref_9_M98_noxref_d ) capacitor c=0.0139598f \
 //x=31.625 //y=7.4 //x2=31.125 //y2=5.02
cc_1450 ( N_VDD_c_1071_n N_noxref_9_M98_noxref_d ) capacitor c=4.9285e-19 \
 //x=33.67 //y=7.4 //x2=31.125 //y2=5.02
cc_1451 ( N_VDD_M96_noxref_s N_noxref_9_M98_noxref_d ) capacitor c=0.00130656f \
 //x=29.815 //y=5.02 //x2=31.125 //y2=5.02
cc_1452 ( N_VDD_M97_noxref_d N_noxref_9_M98_noxref_d ) capacitor c=0.0664752f \
 //x=30.685 //y=5.02 //x2=31.125 //y2=5.02
cc_1453 ( N_VDD_M99_noxref_d N_noxref_9_M98_noxref_d ) capacitor c=0.0664752f \
 //x=31.565 //y=5.02 //x2=31.125 //y2=5.02
cc_1454 ( N_VDD_c_1085_p N_noxref_9_M100_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=32.005 //y2=5.02
cc_1455 ( N_VDD_c_1442_p N_noxref_9_M100_noxref_d ) capacitor c=0.0139598f \
 //x=32.505 //y=7.4 //x2=32.005 //y2=5.02
cc_1456 ( N_VDD_c_1071_n N_noxref_9_M100_noxref_d ) capacitor c=0.00939849f \
 //x=33.67 //y=7.4 //x2=32.005 //y2=5.02
cc_1457 ( N_VDD_M99_noxref_d N_noxref_9_M100_noxref_d ) capacitor c=0.0664752f \
 //x=31.565 //y=5.02 //x2=32.005 //y2=5.02
cc_1458 ( N_VDD_M101_noxref_d N_noxref_9_M100_noxref_d ) capacitor \
 c=0.0664752f //x=32.445 //y=5.02 //x2=32.005 //y2=5.02
cc_1459 ( N_VDD_M102_noxref_s N_noxref_9_M100_noxref_d ) capacitor \
 c=3.57641e-19 //x=34.625 //y=5.02 //x2=32.005 //y2=5.02
cc_1460 ( N_VDD_c_1085_p N_noxref_10_c_4311_n ) capacitor c=0.00437246f \
 //x=95.83 //y=7.4 //x2=40.805 //y2=5.155
cc_1461 ( N_VDD_c_1228_p N_noxref_10_c_4311_n ) capacitor c=4.31596e-19 \
 //x=40.365 //y=7.4 //x2=40.805 //y2=5.155
cc_1462 ( N_VDD_c_1484_p N_noxref_10_c_4311_n ) capacitor c=4.31596e-19 \
 //x=41.245 //y=7.4 //x2=40.805 //y2=5.155
cc_1463 ( N_VDD_M109_noxref_d N_noxref_10_c_4311_n ) capacitor c=0.0109802f \
 //x=40.305 //y=5.02 //x2=40.805 //y2=5.155
cc_1464 ( N_VDD_c_1072_n N_noxref_10_c_4315_n ) capacitor c=0.00863585f \
 //x=38.48 //y=7.4 //x2=40.095 //y2=5.155
cc_1465 ( N_VDD_M108_noxref_s N_noxref_10_c_4315_n ) capacitor c=0.0831083f \
 //x=39.435 //y=5.02 //x2=40.095 //y2=5.155
cc_1466 ( N_VDD_c_1085_p N_noxref_10_c_4317_n ) capacitor c=0.00434259f \
 //x=95.83 //y=7.4 //x2=41.685 //y2=5.155
cc_1467 ( N_VDD_c_1484_p N_noxref_10_c_4317_n ) capacitor c=4.31596e-19 \
 //x=41.245 //y=7.4 //x2=41.685 //y2=5.155
cc_1468 ( N_VDD_c_1490_p N_noxref_10_c_4317_n ) capacitor c=4.31596e-19 \
 //x=42.125 //y=7.4 //x2=41.685 //y2=5.155
cc_1469 ( N_VDD_M111_noxref_d N_noxref_10_c_4317_n ) capacitor c=0.0109802f \
 //x=41.185 //y=5.02 //x2=41.685 //y2=5.155
cc_1470 ( N_VDD_c_1085_p N_noxref_10_c_4321_n ) capacitor c=0.00424413f \
 //x=95.83 //y=7.4 //x2=42.465 //y2=5.155
cc_1471 ( N_VDD_c_1490_p N_noxref_10_c_4321_n ) capacitor c=7.45454e-19 \
 //x=42.125 //y=7.4 //x2=42.465 //y2=5.155
cc_1472 ( N_VDD_c_1229_p N_noxref_10_c_4321_n ) capacitor c=0.00198097f \
 //x=43.12 //y=7.4 //x2=42.465 //y2=5.155
cc_1473 ( N_VDD_M113_noxref_d N_noxref_10_c_4321_n ) capacitor c=0.0109802f \
 //x=42.065 //y=5.02 //x2=42.465 //y2=5.155
cc_1474 ( N_VDD_c_1073_n N_noxref_10_c_4298_n ) capacitor c=0.0400751f \
 //x=43.29 //y=7.4 //x2=42.55 //y2=2.59
cc_1475 ( N_VDD_c_1085_p N_noxref_10_c_4299_n ) capacitor c=6.51035e-19 \
 //x=95.83 //y=7.4 //x2=44.4 //y2=2.08
cc_1476 ( N_VDD_c_1073_n N_noxref_10_c_4299_n ) capacitor c=0.0114465f \
 //x=43.29 //y=7.4 //x2=44.4 //y2=2.08
cc_1477 ( N_VDD_M114_noxref_s N_noxref_10_c_4299_n ) capacitor c=0.00923513f \
 //x=44.245 //y=5.02 //x2=44.4 //y2=2.08
cc_1478 ( N_VDD_c_1231_p N_noxref_10_M114_noxref_g ) capacitor c=0.00749687f \
 //x=45.175 //y=7.4 //x2=44.6 //y2=6.02
cc_1479 ( N_VDD_M114_noxref_s N_noxref_10_M114_noxref_g ) capacitor \
 c=0.0477201f //x=44.245 //y=5.02 //x2=44.6 //y2=6.02
cc_1480 ( N_VDD_c_1231_p N_noxref_10_M115_noxref_g ) capacitor c=0.00675175f \
 //x=45.175 //y=7.4 //x2=45.04 //y2=6.02
cc_1481 ( N_VDD_M115_noxref_d N_noxref_10_M115_noxref_g ) capacitor \
 c=0.015318f //x=45.115 //y=5.02 //x2=45.04 //y2=6.02
cc_1482 ( N_VDD_c_1073_n N_noxref_10_c_4333_n ) capacitor c=0.00528488f \
 //x=43.29 //y=7.4 //x2=44.675 //y2=4.79
cc_1483 ( N_VDD_M114_noxref_s N_noxref_10_c_4333_n ) capacitor c=0.00433385f \
 //x=44.245 //y=5.02 //x2=44.675 //y2=4.79
cc_1484 ( N_VDD_c_1085_p N_noxref_10_M108_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=39.865 //y2=5.02
cc_1485 ( N_VDD_c_1228_p N_noxref_10_M108_noxref_d ) capacitor c=0.0139598f \
 //x=40.365 //y=7.4 //x2=39.865 //y2=5.02
cc_1486 ( N_VDD_M109_noxref_d N_noxref_10_M108_noxref_d ) capacitor \
 c=0.0664752f //x=40.305 //y=5.02 //x2=39.865 //y2=5.02
cc_1487 ( N_VDD_c_1085_p N_noxref_10_M110_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=40.745 //y2=5.02
cc_1488 ( N_VDD_c_1484_p N_noxref_10_M110_noxref_d ) capacitor c=0.0139598f \
 //x=41.245 //y=7.4 //x2=40.745 //y2=5.02
cc_1489 ( N_VDD_c_1073_n N_noxref_10_M110_noxref_d ) capacitor c=4.9285e-19 \
 //x=43.29 //y=7.4 //x2=40.745 //y2=5.02
cc_1490 ( N_VDD_M108_noxref_s N_noxref_10_M110_noxref_d ) capacitor \
 c=0.00130656f //x=39.435 //y=5.02 //x2=40.745 //y2=5.02
cc_1491 ( N_VDD_M109_noxref_d N_noxref_10_M110_noxref_d ) capacitor \
 c=0.0664752f //x=40.305 //y=5.02 //x2=40.745 //y2=5.02
cc_1492 ( N_VDD_M111_noxref_d N_noxref_10_M110_noxref_d ) capacitor \
 c=0.0664752f //x=41.185 //y=5.02 //x2=40.745 //y2=5.02
cc_1493 ( N_VDD_c_1085_p N_noxref_10_M112_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=41.625 //y2=5.02
cc_1494 ( N_VDD_c_1490_p N_noxref_10_M112_noxref_d ) capacitor c=0.0139598f \
 //x=42.125 //y=7.4 //x2=41.625 //y2=5.02
cc_1495 ( N_VDD_c_1073_n N_noxref_10_M112_noxref_d ) capacitor c=0.00939849f \
 //x=43.29 //y=7.4 //x2=41.625 //y2=5.02
cc_1496 ( N_VDD_M111_noxref_d N_noxref_10_M112_noxref_d ) capacitor \
 c=0.0664752f //x=41.185 //y=5.02 //x2=41.625 //y2=5.02
cc_1497 ( N_VDD_M113_noxref_d N_noxref_10_M112_noxref_d ) capacitor \
 c=0.0664752f //x=42.065 //y=5.02 //x2=41.625 //y2=5.02
cc_1498 ( N_VDD_M114_noxref_s N_noxref_10_M112_noxref_d ) capacitor \
 c=3.57641e-19 //x=44.245 //y=5.02 //x2=41.625 //y2=5.02
cc_1499 ( N_VDD_c_1071_n N_noxref_11_c_4464_n ) capacitor c=4.57708e-19 \
 //x=33.67 //y=7.4 //x2=32.19 //y2=2.08
cc_1500 ( N_VDD_c_1085_p N_noxref_11_c_4479_n ) capacitor c=0.00437246f \
 //x=95.83 //y=7.4 //x2=35.995 //y2=5.155
cc_1501 ( N_VDD_c_1225_p N_noxref_11_c_4479_n ) capacitor c=4.31596e-19 \
 //x=35.555 //y=7.4 //x2=35.995 //y2=5.155
cc_1502 ( N_VDD_c_1524_p N_noxref_11_c_4479_n ) capacitor c=4.31596e-19 \
 //x=36.435 //y=7.4 //x2=35.995 //y2=5.155
cc_1503 ( N_VDD_M103_noxref_d N_noxref_11_c_4479_n ) capacitor c=0.0109802f \
 //x=35.495 //y=5.02 //x2=35.995 //y2=5.155
cc_1504 ( N_VDD_c_1071_n N_noxref_11_c_4483_n ) capacitor c=0.00863585f \
 //x=33.67 //y=7.4 //x2=35.285 //y2=5.155
cc_1505 ( N_VDD_M102_noxref_s N_noxref_11_c_4483_n ) capacitor c=0.0831083f \
 //x=34.625 //y=5.02 //x2=35.285 //y2=5.155
cc_1506 ( N_VDD_c_1085_p N_noxref_11_c_4485_n ) capacitor c=0.00434259f \
 //x=95.83 //y=7.4 //x2=36.875 //y2=5.155
cc_1507 ( N_VDD_c_1524_p N_noxref_11_c_4485_n ) capacitor c=4.31596e-19 \
 //x=36.435 //y=7.4 //x2=36.875 //y2=5.155
cc_1508 ( N_VDD_c_1530_p N_noxref_11_c_4485_n ) capacitor c=4.31596e-19 \
 //x=37.315 //y=7.4 //x2=36.875 //y2=5.155
cc_1509 ( N_VDD_M105_noxref_d N_noxref_11_c_4485_n ) capacitor c=0.0109802f \
 //x=36.375 //y=5.02 //x2=36.875 //y2=5.155
cc_1510 ( N_VDD_c_1085_p N_noxref_11_c_4489_n ) capacitor c=0.00424413f \
 //x=95.83 //y=7.4 //x2=37.655 //y2=5.155
cc_1511 ( N_VDD_c_1530_p N_noxref_11_c_4489_n ) capacitor c=7.45454e-19 \
 //x=37.315 //y=7.4 //x2=37.655 //y2=5.155
cc_1512 ( N_VDD_c_1226_p N_noxref_11_c_4489_n ) capacitor c=0.00198097f \
 //x=38.31 //y=7.4 //x2=37.655 //y2=5.155
cc_1513 ( N_VDD_M107_noxref_d N_noxref_11_c_4489_n ) capacitor c=0.0109802f \
 //x=37.255 //y=5.02 //x2=37.655 //y2=5.155
cc_1514 ( N_VDD_c_1072_n N_noxref_11_c_4493_n ) capacitor c=0.0400668f \
 //x=38.48 //y=7.4 //x2=37.74 //y2=3.33
cc_1515 ( N_VDD_c_1085_p N_noxref_11_c_4466_n ) capacitor c=6.51035e-19 \
 //x=95.83 //y=7.4 //x2=49.21 //y2=2.08
cc_1516 ( N_VDD_c_1074_n N_noxref_11_c_4466_n ) capacitor c=0.0115064f \
 //x=48.1 //y=7.4 //x2=49.21 //y2=2.08
cc_1517 ( N_VDD_M120_noxref_s N_noxref_11_c_4466_n ) capacitor c=0.00909681f \
 //x=49.055 //y=5.02 //x2=49.21 //y2=2.08
cc_1518 ( N_VDD_c_1442_p N_noxref_11_M100_noxref_g ) capacitor c=0.00675175f \
 //x=32.505 //y=7.4 //x2=31.93 //y2=6.02
cc_1519 ( N_VDD_M99_noxref_d N_noxref_11_M100_noxref_g ) capacitor c=0.015318f \
 //x=31.565 //y=5.02 //x2=31.93 //y2=6.02
cc_1520 ( N_VDD_c_1442_p N_noxref_11_M101_noxref_g ) capacitor c=0.00675379f \
 //x=32.505 //y=7.4 //x2=32.37 //y2=6.02
cc_1521 ( N_VDD_M101_noxref_d N_noxref_11_M101_noxref_g ) capacitor \
 c=0.0394719f //x=32.445 //y=5.02 //x2=32.37 //y2=6.02
cc_1522 ( N_VDD_c_1234_p N_noxref_11_M120_noxref_g ) capacitor c=0.00749687f \
 //x=49.985 //y=7.4 //x2=49.41 //y2=6.02
cc_1523 ( N_VDD_M120_noxref_s N_noxref_11_M120_noxref_g ) capacitor \
 c=0.0477201f //x=49.055 //y=5.02 //x2=49.41 //y2=6.02
cc_1524 ( N_VDD_c_1234_p N_noxref_11_M121_noxref_g ) capacitor c=0.00675175f \
 //x=49.985 //y=7.4 //x2=49.85 //y2=6.02
cc_1525 ( N_VDD_M121_noxref_d N_noxref_11_M121_noxref_g ) capacitor \
 c=0.015318f //x=49.925 //y=5.02 //x2=49.85 //y2=6.02
cc_1526 ( N_VDD_c_1074_n N_noxref_11_c_4505_n ) capacitor c=0.00528488f \
 //x=48.1 //y=7.4 //x2=49.485 //y2=4.79
cc_1527 ( N_VDD_M120_noxref_s N_noxref_11_c_4505_n ) capacitor c=0.00433385f \
 //x=49.055 //y=5.02 //x2=49.485 //y2=4.79
cc_1528 ( N_VDD_c_1085_p N_noxref_11_M102_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=35.055 //y2=5.02
cc_1529 ( N_VDD_c_1225_p N_noxref_11_M102_noxref_d ) capacitor c=0.0139598f \
 //x=35.555 //y=7.4 //x2=35.055 //y2=5.02
cc_1530 ( N_VDD_M103_noxref_d N_noxref_11_M102_noxref_d ) capacitor \
 c=0.0664752f //x=35.495 //y=5.02 //x2=35.055 //y2=5.02
cc_1531 ( N_VDD_c_1085_p N_noxref_11_M104_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=35.935 //y2=5.02
cc_1532 ( N_VDD_c_1524_p N_noxref_11_M104_noxref_d ) capacitor c=0.0139598f \
 //x=36.435 //y=7.4 //x2=35.935 //y2=5.02
cc_1533 ( N_VDD_c_1072_n N_noxref_11_M104_noxref_d ) capacitor c=4.9285e-19 \
 //x=38.48 //y=7.4 //x2=35.935 //y2=5.02
cc_1534 ( N_VDD_M102_noxref_s N_noxref_11_M104_noxref_d ) capacitor \
 c=0.00130656f //x=34.625 //y=5.02 //x2=35.935 //y2=5.02
cc_1535 ( N_VDD_M103_noxref_d N_noxref_11_M104_noxref_d ) capacitor \
 c=0.0664752f //x=35.495 //y=5.02 //x2=35.935 //y2=5.02
cc_1536 ( N_VDD_M105_noxref_d N_noxref_11_M104_noxref_d ) capacitor \
 c=0.0664752f //x=36.375 //y=5.02 //x2=35.935 //y2=5.02
cc_1537 ( N_VDD_c_1085_p N_noxref_11_M106_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=36.815 //y2=5.02
cc_1538 ( N_VDD_c_1530_p N_noxref_11_M106_noxref_d ) capacitor c=0.0139598f \
 //x=37.315 //y=7.4 //x2=36.815 //y2=5.02
cc_1539 ( N_VDD_c_1072_n N_noxref_11_M106_noxref_d ) capacitor c=0.00939849f \
 //x=38.48 //y=7.4 //x2=36.815 //y2=5.02
cc_1540 ( N_VDD_M105_noxref_d N_noxref_11_M106_noxref_d ) capacitor \
 c=0.0664752f //x=36.375 //y=5.02 //x2=36.815 //y2=5.02
cc_1541 ( N_VDD_M107_noxref_d N_noxref_11_M106_noxref_d ) capacitor \
 c=0.0664752f //x=37.255 //y=5.02 //x2=36.815 //y2=5.02
cc_1542 ( N_VDD_M108_noxref_s N_noxref_11_M106_noxref_d ) capacitor \
 c=3.57641e-19 //x=39.435 //y=5.02 //x2=36.815 //y2=5.02
cc_1543 ( N_VDD_c_1072_n N_noxref_12_c_4745_n ) capacitor c=5.43708e-19 \
 //x=38.48 //y=7.4 //x2=37 //y2=2.08
cc_1544 ( N_VDD_c_1073_n N_noxref_12_c_4746_n ) capacitor c=4.57708e-19 \
 //x=43.29 //y=7.4 //x2=41.81 //y2=2.08
cc_1545 ( N_VDD_c_1085_p N_noxref_12_c_4752_n ) capacitor c=0.00437246f \
 //x=95.83 //y=7.4 //x2=45.615 //y2=5.155
cc_1546 ( N_VDD_c_1231_p N_noxref_12_c_4752_n ) capacitor c=4.31596e-19 \
 //x=45.175 //y=7.4 //x2=45.615 //y2=5.155
cc_1547 ( N_VDD_c_1569_p N_noxref_12_c_4752_n ) capacitor c=4.31596e-19 \
 //x=46.055 //y=7.4 //x2=45.615 //y2=5.155
cc_1548 ( N_VDD_M115_noxref_d N_noxref_12_c_4752_n ) capacitor c=0.0109802f \
 //x=45.115 //y=5.02 //x2=45.615 //y2=5.155
cc_1549 ( N_VDD_c_1073_n N_noxref_12_c_4756_n ) capacitor c=0.00863585f \
 //x=43.29 //y=7.4 //x2=44.905 //y2=5.155
cc_1550 ( N_VDD_M114_noxref_s N_noxref_12_c_4756_n ) capacitor c=0.0831083f \
 //x=44.245 //y=5.02 //x2=44.905 //y2=5.155
cc_1551 ( N_VDD_c_1085_p N_noxref_12_c_4758_n ) capacitor c=0.00434259f \
 //x=95.83 //y=7.4 //x2=46.495 //y2=5.155
cc_1552 ( N_VDD_c_1569_p N_noxref_12_c_4758_n ) capacitor c=4.31596e-19 \
 //x=46.055 //y=7.4 //x2=46.495 //y2=5.155
cc_1553 ( N_VDD_c_1575_p N_noxref_12_c_4758_n ) capacitor c=4.31596e-19 \
 //x=46.935 //y=7.4 //x2=46.495 //y2=5.155
cc_1554 ( N_VDD_M117_noxref_d N_noxref_12_c_4758_n ) capacitor c=0.0109802f \
 //x=45.995 //y=5.02 //x2=46.495 //y2=5.155
cc_1555 ( N_VDD_c_1085_p N_noxref_12_c_4762_n ) capacitor c=0.00424413f \
 //x=95.83 //y=7.4 //x2=47.275 //y2=5.155
cc_1556 ( N_VDD_c_1575_p N_noxref_12_c_4762_n ) capacitor c=7.45454e-19 \
 //x=46.935 //y=7.4 //x2=47.275 //y2=5.155
cc_1557 ( N_VDD_c_1232_p N_noxref_12_c_4762_n ) capacitor c=0.00198097f \
 //x=47.93 //y=7.4 //x2=47.275 //y2=5.155
cc_1558 ( N_VDD_M119_noxref_d N_noxref_12_c_4762_n ) capacitor c=0.0109802f \
 //x=46.875 //y=5.02 //x2=47.275 //y2=5.155
cc_1559 ( N_VDD_c_1074_n N_noxref_12_c_4766_n ) capacitor c=0.0400668f \
 //x=48.1 //y=7.4 //x2=47.36 //y2=3.7
cc_1560 ( N_VDD_c_1076_n N_noxref_12_c_4748_n ) capacitor c=4.93757e-19 \
 //x=57.72 //y=7.4 //x2=56.24 //y2=2.08
cc_1561 ( N_VDD_c_1530_p N_noxref_12_M106_noxref_g ) capacitor c=0.00675175f \
 //x=37.315 //y=7.4 //x2=36.74 //y2=6.02
cc_1562 ( N_VDD_M105_noxref_d N_noxref_12_M106_noxref_g ) capacitor \
 c=0.015318f //x=36.375 //y=5.02 //x2=36.74 //y2=6.02
cc_1563 ( N_VDD_c_1530_p N_noxref_12_M107_noxref_g ) capacitor c=0.00675379f \
 //x=37.315 //y=7.4 //x2=37.18 //y2=6.02
cc_1564 ( N_VDD_M107_noxref_d N_noxref_12_M107_noxref_g ) capacitor \
 c=0.0394719f //x=37.255 //y=5.02 //x2=37.18 //y2=6.02
cc_1565 ( N_VDD_c_1490_p N_noxref_12_M112_noxref_g ) capacitor c=0.00675175f \
 //x=42.125 //y=7.4 //x2=41.55 //y2=6.02
cc_1566 ( N_VDD_M111_noxref_d N_noxref_12_M112_noxref_g ) capacitor \
 c=0.015318f //x=41.185 //y=5.02 //x2=41.55 //y2=6.02
cc_1567 ( N_VDD_c_1490_p N_noxref_12_M113_noxref_g ) capacitor c=0.00675379f \
 //x=42.125 //y=7.4 //x2=41.99 //y2=6.02
cc_1568 ( N_VDD_M113_noxref_d N_noxref_12_M113_noxref_g ) capacitor \
 c=0.0394719f //x=42.065 //y=5.02 //x2=41.99 //y2=6.02
cc_1569 ( N_VDD_c_1591_p N_noxref_12_M130_noxref_g ) capacitor c=0.00675175f \
 //x=56.555 //y=7.4 //x2=55.98 //y2=6.02
cc_1570 ( N_VDD_M129_noxref_d N_noxref_12_M130_noxref_g ) capacitor \
 c=0.015318f //x=55.615 //y=5.02 //x2=55.98 //y2=6.02
cc_1571 ( N_VDD_c_1591_p N_noxref_12_M131_noxref_g ) capacitor c=0.00675379f \
 //x=56.555 //y=7.4 //x2=56.42 //y2=6.02
cc_1572 ( N_VDD_M131_noxref_d N_noxref_12_M131_noxref_g ) capacitor \
 c=0.0394719f //x=56.495 //y=5.02 //x2=56.42 //y2=6.02
cc_1573 ( N_VDD_c_1085_p N_noxref_12_M114_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=44.675 //y2=5.02
cc_1574 ( N_VDD_c_1231_p N_noxref_12_M114_noxref_d ) capacitor c=0.0139598f \
 //x=45.175 //y=7.4 //x2=44.675 //y2=5.02
cc_1575 ( N_VDD_M115_noxref_d N_noxref_12_M114_noxref_d ) capacitor \
 c=0.0664752f //x=45.115 //y=5.02 //x2=44.675 //y2=5.02
cc_1576 ( N_VDD_c_1085_p N_noxref_12_M116_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=45.555 //y2=5.02
cc_1577 ( N_VDD_c_1569_p N_noxref_12_M116_noxref_d ) capacitor c=0.0139598f \
 //x=46.055 //y=7.4 //x2=45.555 //y2=5.02
cc_1578 ( N_VDD_c_1074_n N_noxref_12_M116_noxref_d ) capacitor c=4.9285e-19 \
 //x=48.1 //y=7.4 //x2=45.555 //y2=5.02
cc_1579 ( N_VDD_M114_noxref_s N_noxref_12_M116_noxref_d ) capacitor \
 c=0.00130656f //x=44.245 //y=5.02 //x2=45.555 //y2=5.02
cc_1580 ( N_VDD_M115_noxref_d N_noxref_12_M116_noxref_d ) capacitor \
 c=0.0664752f //x=45.115 //y=5.02 //x2=45.555 //y2=5.02
cc_1581 ( N_VDD_M117_noxref_d N_noxref_12_M116_noxref_d ) capacitor \
 c=0.0664752f //x=45.995 //y=5.02 //x2=45.555 //y2=5.02
cc_1582 ( N_VDD_c_1085_p N_noxref_12_M118_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=46.435 //y2=5.02
cc_1583 ( N_VDD_c_1575_p N_noxref_12_M118_noxref_d ) capacitor c=0.0139598f \
 //x=46.935 //y=7.4 //x2=46.435 //y2=5.02
cc_1584 ( N_VDD_c_1074_n N_noxref_12_M118_noxref_d ) capacitor c=0.00939849f \
 //x=48.1 //y=7.4 //x2=46.435 //y2=5.02
cc_1585 ( N_VDD_M117_noxref_d N_noxref_12_M118_noxref_d ) capacitor \
 c=0.0664752f //x=45.995 //y=5.02 //x2=46.435 //y2=5.02
cc_1586 ( N_VDD_M119_noxref_d N_noxref_12_M118_noxref_d ) capacitor \
 c=0.0664752f //x=46.875 //y=5.02 //x2=46.435 //y2=5.02
cc_1587 ( N_VDD_M120_noxref_s N_noxref_12_M118_noxref_d ) capacitor \
 c=3.57641e-19 //x=49.055 //y=5.02 //x2=46.435 //y2=5.02
cc_1588 ( N_VDD_c_1075_n N_noxref_13_c_5101_n ) capacitor c=4.57708e-19 \
 //x=52.91 //y=7.4 //x2=51.43 //y2=2.08
cc_1589 ( N_VDD_c_1085_p N_noxref_13_c_5106_n ) capacitor c=0.00437246f \
 //x=95.83 //y=7.4 //x2=55.235 //y2=5.155
cc_1590 ( N_VDD_c_1237_p N_noxref_13_c_5106_n ) capacitor c=4.31596e-19 \
 //x=54.795 //y=7.4 //x2=55.235 //y2=5.155
cc_1591 ( N_VDD_c_1613_p N_noxref_13_c_5106_n ) capacitor c=4.31596e-19 \
 //x=55.675 //y=7.4 //x2=55.235 //y2=5.155
cc_1592 ( N_VDD_M127_noxref_d N_noxref_13_c_5106_n ) capacitor c=0.0109802f \
 //x=54.735 //y=5.02 //x2=55.235 //y2=5.155
cc_1593 ( N_VDD_c_1075_n N_noxref_13_c_5110_n ) capacitor c=0.00863585f \
 //x=52.91 //y=7.4 //x2=54.525 //y2=5.155
cc_1594 ( N_VDD_M126_noxref_s N_noxref_13_c_5110_n ) capacitor c=0.0831083f \
 //x=53.865 //y=5.02 //x2=54.525 //y2=5.155
cc_1595 ( N_VDD_c_1085_p N_noxref_13_c_5112_n ) capacitor c=0.00434259f \
 //x=95.83 //y=7.4 //x2=56.115 //y2=5.155
cc_1596 ( N_VDD_c_1613_p N_noxref_13_c_5112_n ) capacitor c=4.31596e-19 \
 //x=55.675 //y=7.4 //x2=56.115 //y2=5.155
cc_1597 ( N_VDD_c_1591_p N_noxref_13_c_5112_n ) capacitor c=4.31596e-19 \
 //x=56.555 //y=7.4 //x2=56.115 //y2=5.155
cc_1598 ( N_VDD_M129_noxref_d N_noxref_13_c_5112_n ) capacitor c=0.0109802f \
 //x=55.615 //y=5.02 //x2=56.115 //y2=5.155
cc_1599 ( N_VDD_c_1085_p N_noxref_13_c_5116_n ) capacitor c=0.0042353f \
 //x=95.83 //y=7.4 //x2=56.895 //y2=5.155
cc_1600 ( N_VDD_c_1591_p N_noxref_13_c_5116_n ) capacitor c=7.45454e-19 \
 //x=56.555 //y=7.4 //x2=56.895 //y2=5.155
cc_1601 ( N_VDD_c_1238_p N_noxref_13_c_5116_n ) capacitor c=0.00198097f \
 //x=57.55 //y=7.4 //x2=56.895 //y2=5.155
cc_1602 ( N_VDD_M131_noxref_d N_noxref_13_c_5116_n ) capacitor c=0.0109802f \
 //x=56.495 //y=5.02 //x2=56.895 //y2=5.155
cc_1603 ( N_VDD_c_1076_n N_noxref_13_c_5103_n ) capacitor c=0.0401063f \
 //x=57.72 //y=7.4 //x2=56.98 //y2=2.59
cc_1604 ( N_VDD_c_1626_p N_noxref_13_M124_noxref_g ) capacitor c=0.00675175f \
 //x=51.745 //y=7.4 //x2=51.17 //y2=6.02
cc_1605 ( N_VDD_M123_noxref_d N_noxref_13_M124_noxref_g ) capacitor \
 c=0.015318f //x=50.805 //y=5.02 //x2=51.17 //y2=6.02
cc_1606 ( N_VDD_c_1626_p N_noxref_13_M125_noxref_g ) capacitor c=0.00675379f \
 //x=51.745 //y=7.4 //x2=51.61 //y2=6.02
cc_1607 ( N_VDD_M125_noxref_d N_noxref_13_M125_noxref_g ) capacitor \
 c=0.0394719f //x=51.685 //y=5.02 //x2=51.61 //y2=6.02
cc_1608 ( N_VDD_c_1085_p N_noxref_13_M126_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=54.295 //y2=5.02
cc_1609 ( N_VDD_c_1237_p N_noxref_13_M126_noxref_d ) capacitor c=0.0139598f \
 //x=54.795 //y=7.4 //x2=54.295 //y2=5.02
cc_1610 ( N_VDD_M127_noxref_d N_noxref_13_M126_noxref_d ) capacitor \
 c=0.0664752f //x=54.735 //y=5.02 //x2=54.295 //y2=5.02
cc_1611 ( N_VDD_c_1085_p N_noxref_13_M128_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=55.175 //y2=5.02
cc_1612 ( N_VDD_c_1613_p N_noxref_13_M128_noxref_d ) capacitor c=0.0139598f \
 //x=55.675 //y=7.4 //x2=55.175 //y2=5.02
cc_1613 ( N_VDD_c_1076_n N_noxref_13_M128_noxref_d ) capacitor c=4.9285e-19 \
 //x=57.72 //y=7.4 //x2=55.175 //y2=5.02
cc_1614 ( N_VDD_M126_noxref_s N_noxref_13_M128_noxref_d ) capacitor \
 c=0.00130656f //x=53.865 //y=5.02 //x2=55.175 //y2=5.02
cc_1615 ( N_VDD_M127_noxref_d N_noxref_13_M128_noxref_d ) capacitor \
 c=0.0664752f //x=54.735 //y=5.02 //x2=55.175 //y2=5.02
cc_1616 ( N_VDD_M129_noxref_d N_noxref_13_M128_noxref_d ) capacitor \
 c=0.0664752f //x=55.615 //y=5.02 //x2=55.175 //y2=5.02
cc_1617 ( N_VDD_c_1085_p N_noxref_13_M130_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=56.055 //y2=5.02
cc_1618 ( N_VDD_c_1591_p N_noxref_13_M130_noxref_d ) capacitor c=0.0139598f \
 //x=56.555 //y=7.4 //x2=56.055 //y2=5.02
cc_1619 ( N_VDD_c_1076_n N_noxref_13_M130_noxref_d ) capacitor c=0.00939849f \
 //x=57.72 //y=7.4 //x2=56.055 //y2=5.02
cc_1620 ( N_VDD_M129_noxref_d N_noxref_13_M130_noxref_d ) capacitor \
 c=0.0664752f //x=55.615 //y=5.02 //x2=56.055 //y2=5.02
cc_1621 ( N_VDD_M131_noxref_d N_noxref_13_M130_noxref_d ) capacitor \
 c=0.0664752f //x=56.495 //y=5.02 //x2=56.055 //y2=5.02
cc_1622 ( N_VDD_M132_noxref_s N_noxref_13_M130_noxref_d ) capacitor \
 c=3.57641e-19 //x=58.675 //y=5.02 //x2=56.055 //y2=5.02
cc_1623 ( N_VDD_c_1085_p N_D_c_5277_n ) capacitor c=0.104182f //x=95.83 \
 //y=7.4 //x2=29.855 //y2=4.07
cc_1624 ( N_VDD_c_1086_p N_D_c_5277_n ) capacitor c=0.00113322f //x=1.885 \
 //y=7.4 //x2=29.855 //y2=4.07
cc_1625 ( N_VDD_c_1097_p N_D_c_5277_n ) capacitor c=0.00214241f //x=4.64 \
 //y=7.4 //x2=29.855 //y2=4.07
cc_1626 ( N_VDD_c_1648_p N_D_c_5277_n ) capacitor c=0.0027159f //x=5.815 \
 //y=7.4 //x2=29.855 //y2=4.07
cc_1627 ( N_VDD_c_1106_p N_D_c_5277_n ) capacitor c=0.00113459f //x=6.695 \
 //y=7.4 //x2=29.855 //y2=4.07
cc_1628 ( N_VDD_c_1065_n N_D_c_5277_n ) capacitor c=0.0272312f //x=4.81 \
 //y=7.4 //x2=29.855 //y2=4.07
cc_1629 ( N_VDD_c_1066_n N_D_c_5277_n ) capacitor c=0.0140578f //x=9.62 \
 //y=7.4 //x2=29.855 //y2=4.07
cc_1630 ( N_VDD_c_1067_n N_D_c_5277_n ) capacitor c=0.0140578f //x=14.43 \
 //y=7.4 //x2=29.855 //y2=4.07
cc_1631 ( N_VDD_c_1068_n N_D_c_5277_n ) capacitor c=0.0140578f //x=19.24 \
 //y=7.4 //x2=29.855 //y2=4.07
cc_1632 ( N_VDD_c_1069_n N_D_c_5277_n ) capacitor c=0.0140578f //x=24.05 \
 //y=7.4 //x2=29.855 //y2=4.07
cc_1633 ( N_VDD_c_1070_n N_D_c_5277_n ) capacitor c=0.0145592f //x=28.86 \
 //y=7.4 //x2=29.855 //y2=4.07
cc_1634 ( N_VDD_M66_noxref_s N_D_c_5277_n ) capacitor c=0.00122826f //x=5.765 \
 //y=5.02 //x2=29.855 //y2=4.07
cc_1635 ( N_VDD_c_1085_p N_D_c_5278_n ) capacitor c=0.00284951f //x=95.83 \
 //y=7.4 //x2=1.225 //y2=4.07
cc_1636 ( N_VDD_c_1658_p N_D_c_5278_n ) capacitor c=3.84396e-19 //x=1.005 \
 //y=7.4 //x2=1.225 //y2=4.07
cc_1637 ( N_VDD_c_1063_n N_D_c_5278_n ) capacitor c=0.0019001f //x=0.74 \
 //y=7.4 //x2=1.225 //y2=4.07
cc_1638 ( N_VDD_M60_noxref_s N_D_c_5278_n ) capacitor c=0.00128242f //x=0.955 \
 //y=5.02 //x2=1.225 //y2=4.07
cc_1639 ( N_VDD_c_1071_n N_D_c_5328_n ) capacitor c=0.0143396f //x=33.67 \
 //y=7.4 //x2=58.715 //y2=4.07
cc_1640 ( N_VDD_c_1072_n N_D_c_5328_n ) capacitor c=0.0140578f //x=38.48 \
 //y=7.4 //x2=58.715 //y2=4.07
cc_1641 ( N_VDD_c_1073_n N_D_c_5328_n ) capacitor c=0.0140578f //x=43.29 \
 //y=7.4 //x2=58.715 //y2=4.07
cc_1642 ( N_VDD_c_1074_n N_D_c_5328_n ) capacitor c=0.0140578f //x=48.1 \
 //y=7.4 //x2=58.715 //y2=4.07
cc_1643 ( N_VDD_c_1075_n N_D_c_5328_n ) capacitor c=0.0140578f //x=52.91 \
 //y=7.4 //x2=58.715 //y2=4.07
cc_1644 ( N_VDD_c_1076_n N_D_c_5328_n ) capacitor c=0.0148105f //x=57.72 \
 //y=7.4 //x2=58.715 //y2=4.07
cc_1645 ( N_VDD_c_1070_n N_D_c_5334_n ) capacitor c=7.52739e-19 //x=28.86 \
 //y=7.4 //x2=30.085 //y2=4.07
cc_1646 ( N_VDD_c_1085_p N_D_c_5279_n ) capacitor c=9.2251e-19 //x=95.83 \
 //y=7.4 //x2=1.11 //y2=2.08
cc_1647 ( N_VDD_c_1063_n N_D_c_5279_n ) capacitor c=0.016255f //x=0.74 //y=7.4 \
 //x2=1.11 //y2=2.08
cc_1648 ( N_VDD_M60_noxref_s N_D_c_5279_n ) capacitor c=0.0122951f //x=0.955 \
 //y=5.02 //x2=1.11 //y2=2.08
cc_1649 ( N_VDD_c_1085_p N_D_c_5280_n ) capacitor c=6.51035e-19 //x=95.83 \
 //y=7.4 //x2=29.97 //y2=2.08
cc_1650 ( N_VDD_c_1070_n N_D_c_5280_n ) capacitor c=0.0113781f //x=28.86 \
 //y=7.4 //x2=29.97 //y2=2.08
cc_1651 ( N_VDD_M96_noxref_s N_D_c_5280_n ) capacitor c=0.00862885f //x=29.815 \
 //y=5.02 //x2=29.97 //y2=2.08
cc_1652 ( N_VDD_c_1085_p N_D_c_5281_n ) capacitor c=6.51035e-19 //x=95.83 \
 //y=7.4 //x2=58.83 //y2=2.08
cc_1653 ( N_VDD_c_1076_n N_D_c_5281_n ) capacitor c=0.0113781f //x=57.72 \
 //y=7.4 //x2=58.83 //y2=2.08
cc_1654 ( N_VDD_M132_noxref_s N_D_c_5281_n ) capacitor c=0.00862885f \
 //x=58.675 //y=5.02 //x2=58.83 //y2=2.08
cc_1655 ( N_VDD_c_1086_p N_D_M60_noxref_g ) capacitor c=0.00749687f //x=1.885 \
 //y=7.4 //x2=1.31 //y2=6.02
cc_1656 ( N_VDD_M60_noxref_s N_D_M60_noxref_g ) capacitor c=0.0477201f \
 //x=0.955 //y=5.02 //x2=1.31 //y2=6.02
cc_1657 ( N_VDD_c_1086_p N_D_M61_noxref_g ) capacitor c=0.00675175f //x=1.885 \
 //y=7.4 //x2=1.75 //y2=6.02
cc_1658 ( N_VDD_M61_noxref_d N_D_M61_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=1.75 //y2=6.02
cc_1659 ( N_VDD_c_1222_p N_D_M96_noxref_g ) capacitor c=0.00749687f //x=30.745 \
 //y=7.4 //x2=30.17 //y2=6.02
cc_1660 ( N_VDD_M96_noxref_s N_D_M96_noxref_g ) capacitor c=0.0477201f \
 //x=29.815 //y=5.02 //x2=30.17 //y2=6.02
cc_1661 ( N_VDD_c_1222_p N_D_M97_noxref_g ) capacitor c=0.00675175f //x=30.745 \
 //y=7.4 //x2=30.61 //y2=6.02
cc_1662 ( N_VDD_M97_noxref_d N_D_M97_noxref_g ) capacitor c=0.015318f \
 //x=30.685 //y=5.02 //x2=30.61 //y2=6.02
cc_1663 ( N_VDD_c_1240_p N_D_M132_noxref_g ) capacitor c=0.00749687f \
 //x=59.605 //y=7.4 //x2=59.03 //y2=6.02
cc_1664 ( N_VDD_M132_noxref_s N_D_M132_noxref_g ) capacitor c=0.0477201f \
 //x=58.675 //y=5.02 //x2=59.03 //y2=6.02
cc_1665 ( N_VDD_c_1240_p N_D_M133_noxref_g ) capacitor c=0.00675175f \
 //x=59.605 //y=7.4 //x2=59.47 //y2=6.02
cc_1666 ( N_VDD_M133_noxref_d N_D_M133_noxref_g ) capacitor c=0.015318f \
 //x=59.545 //y=5.02 //x2=59.47 //y2=6.02
cc_1667 ( N_VDD_c_1063_n N_D_c_5356_n ) capacitor c=0.0076931f //x=0.74 \
 //y=7.4 //x2=1.385 //y2=4.79
cc_1668 ( N_VDD_M60_noxref_s N_D_c_5356_n ) capacitor c=0.00445117f //x=0.955 \
 //y=5.02 //x2=1.385 //y2=4.79
cc_1669 ( N_VDD_c_1070_n N_D_c_5358_n ) capacitor c=0.00540116f //x=28.86 \
 //y=7.4 //x2=30.245 //y2=4.79
cc_1670 ( N_VDD_M96_noxref_s N_D_c_5358_n ) capacitor c=0.00433385f //x=29.815 \
 //y=5.02 //x2=30.245 //y2=4.79
cc_1671 ( N_VDD_c_1076_n N_D_c_5360_n ) capacitor c=0.00540116f //x=57.72 \
 //y=7.4 //x2=59.105 //y2=4.79
cc_1672 ( N_VDD_M132_noxref_s N_D_c_5360_n ) capacitor c=0.00433385f \
 //x=58.675 //y=5.02 //x2=59.105 //y2=4.79
cc_1673 ( N_VDD_c_1085_p N_noxref_15_c_5648_n ) capacitor c=0.00437246f \
 //x=95.83 //y=7.4 //x2=60.045 //y2=5.155
cc_1674 ( N_VDD_c_1240_p N_noxref_15_c_5648_n ) capacitor c=4.31596e-19 \
 //x=59.605 //y=7.4 //x2=60.045 //y2=5.155
cc_1675 ( N_VDD_c_1697_p N_noxref_15_c_5648_n ) capacitor c=4.31596e-19 \
 //x=60.485 //y=7.4 //x2=60.045 //y2=5.155
cc_1676 ( N_VDD_M133_noxref_d N_noxref_15_c_5648_n ) capacitor c=0.0109802f \
 //x=59.545 //y=5.02 //x2=60.045 //y2=5.155
cc_1677 ( N_VDD_c_1076_n N_noxref_15_c_5652_n ) capacitor c=0.00863585f \
 //x=57.72 //y=7.4 //x2=59.335 //y2=5.155
cc_1678 ( N_VDD_M132_noxref_s N_noxref_15_c_5652_n ) capacitor c=0.0831083f \
 //x=58.675 //y=5.02 //x2=59.335 //y2=5.155
cc_1679 ( N_VDD_c_1085_p N_noxref_15_c_5654_n ) capacitor c=0.00434259f \
 //x=95.83 //y=7.4 //x2=60.925 //y2=5.155
cc_1680 ( N_VDD_c_1697_p N_noxref_15_c_5654_n ) capacitor c=4.31596e-19 \
 //x=60.485 //y=7.4 //x2=60.925 //y2=5.155
cc_1681 ( N_VDD_c_1703_p N_noxref_15_c_5654_n ) capacitor c=4.31596e-19 \
 //x=61.365 //y=7.4 //x2=60.925 //y2=5.155
cc_1682 ( N_VDD_M135_noxref_d N_noxref_15_c_5654_n ) capacitor c=0.0109802f \
 //x=60.425 //y=5.02 //x2=60.925 //y2=5.155
cc_1683 ( N_VDD_c_1085_p N_noxref_15_c_5658_n ) capacitor c=0.00424413f \
 //x=95.83 //y=7.4 //x2=61.705 //y2=5.155
cc_1684 ( N_VDD_c_1703_p N_noxref_15_c_5658_n ) capacitor c=7.45454e-19 \
 //x=61.365 //y=7.4 //x2=61.705 //y2=5.155
cc_1685 ( N_VDD_c_1241_p N_noxref_15_c_5658_n ) capacitor c=0.00198097f \
 //x=62.36 //y=7.4 //x2=61.705 //y2=5.155
cc_1686 ( N_VDD_M137_noxref_d N_noxref_15_c_5658_n ) capacitor c=0.0109802f \
 //x=61.305 //y=5.02 //x2=61.705 //y2=5.155
cc_1687 ( N_VDD_c_1077_n N_noxref_15_c_5624_n ) capacitor c=0.0406991f \
 //x=62.53 //y=7.4 //x2=61.79 //y2=2.59
cc_1688 ( N_VDD_c_1085_p N_noxref_15_c_5625_n ) capacitor c=6.51035e-19 \
 //x=95.83 //y=7.4 //x2=63.64 //y2=2.08
cc_1689 ( N_VDD_c_1077_n N_noxref_15_c_5625_n ) capacitor c=0.0120774f \
 //x=62.53 //y=7.4 //x2=63.64 //y2=2.08
cc_1690 ( N_VDD_M138_noxref_s N_noxref_15_c_5625_n ) capacitor c=0.00909681f \
 //x=63.485 //y=5.02 //x2=63.64 //y2=2.08
cc_1691 ( N_VDD_c_1085_p N_noxref_15_c_5626_n ) capacitor c=6.51035e-19 \
 //x=95.83 //y=7.4 //x2=68.45 //y2=2.08
cc_1692 ( N_VDD_c_1078_n N_noxref_15_c_5626_n ) capacitor c=0.0115064f \
 //x=67.34 //y=7.4 //x2=68.45 //y2=2.08
cc_1693 ( N_VDD_M144_noxref_s N_noxref_15_c_5626_n ) capacitor c=0.00923513f \
 //x=68.295 //y=5.02 //x2=68.45 //y2=2.08
cc_1694 ( N_VDD_c_1243_p N_noxref_15_M138_noxref_g ) capacitor c=0.00749687f \
 //x=64.415 //y=7.4 //x2=63.84 //y2=6.02
cc_1695 ( N_VDD_M138_noxref_s N_noxref_15_M138_noxref_g ) capacitor \
 c=0.0477201f //x=63.485 //y=5.02 //x2=63.84 //y2=6.02
cc_1696 ( N_VDD_c_1243_p N_noxref_15_M139_noxref_g ) capacitor c=0.00675175f \
 //x=64.415 //y=7.4 //x2=64.28 //y2=6.02
cc_1697 ( N_VDD_M139_noxref_d N_noxref_15_M139_noxref_g ) capacitor \
 c=0.015318f //x=64.355 //y=5.02 //x2=64.28 //y2=6.02
cc_1698 ( N_VDD_c_1246_p N_noxref_15_M144_noxref_g ) capacitor c=0.00749687f \
 //x=69.225 //y=7.4 //x2=68.65 //y2=6.02
cc_1699 ( N_VDD_M144_noxref_s N_noxref_15_M144_noxref_g ) capacitor \
 c=0.0477201f //x=68.295 //y=5.02 //x2=68.65 //y2=6.02
cc_1700 ( N_VDD_c_1246_p N_noxref_15_M145_noxref_g ) capacitor c=0.00675175f \
 //x=69.225 //y=7.4 //x2=69.09 //y2=6.02
cc_1701 ( N_VDD_M145_noxref_d N_noxref_15_M145_noxref_g ) capacitor \
 c=0.015318f //x=69.165 //y=5.02 //x2=69.09 //y2=6.02
cc_1702 ( N_VDD_c_1077_n N_noxref_15_c_5677_n ) capacitor c=0.00528488f \
 //x=62.53 //y=7.4 //x2=63.915 //y2=4.79
cc_1703 ( N_VDD_M138_noxref_s N_noxref_15_c_5677_n ) capacitor c=0.00433385f \
 //x=63.485 //y=5.02 //x2=63.915 //y2=4.79
cc_1704 ( N_VDD_c_1078_n N_noxref_15_c_5679_n ) capacitor c=0.00528488f \
 //x=67.34 //y=7.4 //x2=68.725 //y2=4.79
cc_1705 ( N_VDD_M144_noxref_s N_noxref_15_c_5679_n ) capacitor c=0.00433385f \
 //x=68.295 //y=5.02 //x2=68.725 //y2=4.79
cc_1706 ( N_VDD_c_1085_p N_noxref_15_M132_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=59.105 //y2=5.02
cc_1707 ( N_VDD_c_1240_p N_noxref_15_M132_noxref_d ) capacitor c=0.0139598f \
 //x=59.605 //y=7.4 //x2=59.105 //y2=5.02
cc_1708 ( N_VDD_M133_noxref_d N_noxref_15_M132_noxref_d ) capacitor \
 c=0.0664752f //x=59.545 //y=5.02 //x2=59.105 //y2=5.02
cc_1709 ( N_VDD_c_1085_p N_noxref_15_M134_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=59.985 //y2=5.02
cc_1710 ( N_VDD_c_1697_p N_noxref_15_M134_noxref_d ) capacitor c=0.0139598f \
 //x=60.485 //y=7.4 //x2=59.985 //y2=5.02
cc_1711 ( N_VDD_c_1077_n N_noxref_15_M134_noxref_d ) capacitor c=4.9285e-19 \
 //x=62.53 //y=7.4 //x2=59.985 //y2=5.02
cc_1712 ( N_VDD_M132_noxref_s N_noxref_15_M134_noxref_d ) capacitor \
 c=0.00130656f //x=58.675 //y=5.02 //x2=59.985 //y2=5.02
cc_1713 ( N_VDD_M133_noxref_d N_noxref_15_M134_noxref_d ) capacitor \
 c=0.0664752f //x=59.545 //y=5.02 //x2=59.985 //y2=5.02
cc_1714 ( N_VDD_M135_noxref_d N_noxref_15_M134_noxref_d ) capacitor \
 c=0.0664752f //x=60.425 //y=5.02 //x2=59.985 //y2=5.02
cc_1715 ( N_VDD_c_1085_p N_noxref_15_M136_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=60.865 //y2=5.02
cc_1716 ( N_VDD_c_1703_p N_noxref_15_M136_noxref_d ) capacitor c=0.0139598f \
 //x=61.365 //y=7.4 //x2=60.865 //y2=5.02
cc_1717 ( N_VDD_c_1077_n N_noxref_15_M136_noxref_d ) capacitor c=0.00939849f \
 //x=62.53 //y=7.4 //x2=60.865 //y2=5.02
cc_1718 ( N_VDD_M135_noxref_d N_noxref_15_M136_noxref_d ) capacitor \
 c=0.0664752f //x=60.425 //y=5.02 //x2=60.865 //y2=5.02
cc_1719 ( N_VDD_M137_noxref_d N_noxref_15_M136_noxref_d ) capacitor \
 c=0.0664752f //x=61.305 //y=5.02 //x2=60.865 //y2=5.02
cc_1720 ( N_VDD_M138_noxref_s N_noxref_15_M136_noxref_d ) capacitor \
 c=3.57641e-19 //x=63.485 //y=5.02 //x2=60.865 //y2=5.02
cc_1721 ( N_VDD_c_1085_p N_noxref_16_c_5888_n ) capacitor c=0.00437246f \
 //x=95.83 //y=7.4 //x2=69.665 //y2=5.155
cc_1722 ( N_VDD_c_1246_p N_noxref_16_c_5888_n ) capacitor c=4.31596e-19 \
 //x=69.225 //y=7.4 //x2=69.665 //y2=5.155
cc_1723 ( N_VDD_c_1745_p N_noxref_16_c_5888_n ) capacitor c=4.31596e-19 \
 //x=70.105 //y=7.4 //x2=69.665 //y2=5.155
cc_1724 ( N_VDD_M145_noxref_d N_noxref_16_c_5888_n ) capacitor c=0.0109802f \
 //x=69.165 //y=5.02 //x2=69.665 //y2=5.155
cc_1725 ( N_VDD_c_1078_n N_noxref_16_c_5892_n ) capacitor c=0.00863585f \
 //x=67.34 //y=7.4 //x2=68.955 //y2=5.155
cc_1726 ( N_VDD_M144_noxref_s N_noxref_16_c_5892_n ) capacitor c=0.0831083f \
 //x=68.295 //y=5.02 //x2=68.955 //y2=5.155
cc_1727 ( N_VDD_c_1085_p N_noxref_16_c_5894_n ) capacitor c=0.00434259f \
 //x=95.83 //y=7.4 //x2=70.545 //y2=5.155
cc_1728 ( N_VDD_c_1745_p N_noxref_16_c_5894_n ) capacitor c=4.31596e-19 \
 //x=70.105 //y=7.4 //x2=70.545 //y2=5.155
cc_1729 ( N_VDD_c_1751_p N_noxref_16_c_5894_n ) capacitor c=4.31596e-19 \
 //x=70.985 //y=7.4 //x2=70.545 //y2=5.155
cc_1730 ( N_VDD_M147_noxref_d N_noxref_16_c_5894_n ) capacitor c=0.0109802f \
 //x=70.045 //y=5.02 //x2=70.545 //y2=5.155
cc_1731 ( N_VDD_c_1085_p N_noxref_16_c_5898_n ) capacitor c=0.00424413f \
 //x=95.83 //y=7.4 //x2=71.325 //y2=5.155
cc_1732 ( N_VDD_c_1751_p N_noxref_16_c_5898_n ) capacitor c=7.45454e-19 \
 //x=70.985 //y=7.4 //x2=71.325 //y2=5.155
cc_1733 ( N_VDD_c_1247_p N_noxref_16_c_5898_n ) capacitor c=0.00198097f \
 //x=71.98 //y=7.4 //x2=71.325 //y2=5.155
cc_1734 ( N_VDD_M149_noxref_d N_noxref_16_c_5898_n ) capacitor c=0.0109802f \
 //x=70.925 //y=5.02 //x2=71.325 //y2=5.155
cc_1735 ( N_VDD_c_1079_n N_noxref_16_c_5875_n ) capacitor c=0.0400751f \
 //x=72.15 //y=7.4 //x2=71.41 //y2=2.59
cc_1736 ( N_VDD_c_1085_p N_noxref_16_c_5876_n ) capacitor c=6.51035e-19 \
 //x=95.83 //y=7.4 //x2=73.26 //y2=2.08
cc_1737 ( N_VDD_c_1079_n N_noxref_16_c_5876_n ) capacitor c=0.0114261f \
 //x=72.15 //y=7.4 //x2=73.26 //y2=2.08
cc_1738 ( N_VDD_M150_noxref_s N_noxref_16_c_5876_n ) capacitor c=0.00923513f \
 //x=73.105 //y=5.02 //x2=73.26 //y2=2.08
cc_1739 ( N_VDD_c_1249_p N_noxref_16_M150_noxref_g ) capacitor c=0.00749687f \
 //x=74.035 //y=7.4 //x2=73.46 //y2=6.02
cc_1740 ( N_VDD_M150_noxref_s N_noxref_16_M150_noxref_g ) capacitor \
 c=0.0477201f //x=73.105 //y=5.02 //x2=73.46 //y2=6.02
cc_1741 ( N_VDD_c_1249_p N_noxref_16_M151_noxref_g ) capacitor c=0.00675175f \
 //x=74.035 //y=7.4 //x2=73.9 //y2=6.02
cc_1742 ( N_VDD_M151_noxref_d N_noxref_16_M151_noxref_g ) capacitor \
 c=0.015318f //x=73.975 //y=5.02 //x2=73.9 //y2=6.02
cc_1743 ( N_VDD_c_1079_n N_noxref_16_c_5910_n ) capacitor c=0.00429651f \
 //x=72.15 //y=7.4 //x2=73.535 //y2=4.79
cc_1744 ( N_VDD_M150_noxref_s N_noxref_16_c_5910_n ) capacitor c=0.00433385f \
 //x=73.105 //y=5.02 //x2=73.535 //y2=4.79
cc_1745 ( N_VDD_c_1085_p N_noxref_16_M144_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=68.725 //y2=5.02
cc_1746 ( N_VDD_c_1246_p N_noxref_16_M144_noxref_d ) capacitor c=0.0139598f \
 //x=69.225 //y=7.4 //x2=68.725 //y2=5.02
cc_1747 ( N_VDD_M145_noxref_d N_noxref_16_M144_noxref_d ) capacitor \
 c=0.0664752f //x=69.165 //y=5.02 //x2=68.725 //y2=5.02
cc_1748 ( N_VDD_c_1085_p N_noxref_16_M146_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=69.605 //y2=5.02
cc_1749 ( N_VDD_c_1745_p N_noxref_16_M146_noxref_d ) capacitor c=0.0139598f \
 //x=70.105 //y=7.4 //x2=69.605 //y2=5.02
cc_1750 ( N_VDD_c_1079_n N_noxref_16_M146_noxref_d ) capacitor c=4.9285e-19 \
 //x=72.15 //y=7.4 //x2=69.605 //y2=5.02
cc_1751 ( N_VDD_M144_noxref_s N_noxref_16_M146_noxref_d ) capacitor \
 c=0.00130656f //x=68.295 //y=5.02 //x2=69.605 //y2=5.02
cc_1752 ( N_VDD_M145_noxref_d N_noxref_16_M146_noxref_d ) capacitor \
 c=0.0664752f //x=69.165 //y=5.02 //x2=69.605 //y2=5.02
cc_1753 ( N_VDD_M147_noxref_d N_noxref_16_M146_noxref_d ) capacitor \
 c=0.0664752f //x=70.045 //y=5.02 //x2=69.605 //y2=5.02
cc_1754 ( N_VDD_c_1085_p N_noxref_16_M148_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=70.485 //y2=5.02
cc_1755 ( N_VDD_c_1751_p N_noxref_16_M148_noxref_d ) capacitor c=0.0139598f \
 //x=70.985 //y=7.4 //x2=70.485 //y2=5.02
cc_1756 ( N_VDD_c_1079_n N_noxref_16_M148_noxref_d ) capacitor c=0.00939849f \
 //x=72.15 //y=7.4 //x2=70.485 //y2=5.02
cc_1757 ( N_VDD_M147_noxref_d N_noxref_16_M148_noxref_d ) capacitor \
 c=0.0664752f //x=70.045 //y=5.02 //x2=70.485 //y2=5.02
cc_1758 ( N_VDD_M149_noxref_d N_noxref_16_M148_noxref_d ) capacitor \
 c=0.0664752f //x=70.925 //y=5.02 //x2=70.485 //y2=5.02
cc_1759 ( N_VDD_M150_noxref_s N_noxref_16_M148_noxref_d ) capacitor \
 c=3.57641e-19 //x=73.105 //y=5.02 //x2=70.485 //y2=5.02
cc_1760 ( N_VDD_c_1085_p N_CLK_c_6046_n ) capacitor c=0.071114f //x=95.83 \
 //y=7.4 //x2=16.535 //y2=4.44
cc_1761 ( N_VDD_c_1185_p N_CLK_c_6046_n ) capacitor c=0.00258496f //x=9.45 \
 //y=7.4 //x2=16.535 //y2=4.44
cc_1762 ( N_VDD_c_1784_p N_CLK_c_6046_n ) capacitor c=0.00328994f //x=10.625 \
 //y=7.4 //x2=16.535 //y2=4.44
cc_1763 ( N_VDD_c_1110_p N_CLK_c_6046_n ) capacitor c=0.00135925f //x=11.505 \
 //y=7.4 //x2=16.535 //y2=4.44
cc_1764 ( N_VDD_c_1145_p N_CLK_c_6046_n ) capacitor c=0.00258496f //x=14.26 \
 //y=7.4 //x2=16.535 //y2=4.44
cc_1765 ( N_VDD_c_1787_p N_CLK_c_6046_n ) capacitor c=0.00328994f //x=15.435 \
 //y=7.4 //x2=16.535 //y2=4.44
cc_1766 ( N_VDD_c_1151_p N_CLK_c_6046_n ) capacitor c=0.00135925f //x=16.315 \
 //y=7.4 //x2=16.535 //y2=4.44
cc_1767 ( N_VDD_c_1066_n N_CLK_c_6046_n ) capacitor c=0.0389825f //x=9.62 \
 //y=7.4 //x2=16.535 //y2=4.44
cc_1768 ( N_VDD_c_1067_n N_CLK_c_6046_n ) capacitor c=0.0389825f //x=14.43 \
 //y=7.4 //x2=16.535 //y2=4.44
cc_1769 ( N_VDD_M72_noxref_s N_CLK_c_6046_n ) capacitor c=0.00179496f \
 //x=10.575 //y=5.02 //x2=16.535 //y2=4.44
cc_1770 ( N_VDD_M78_noxref_s N_CLK_c_6046_n ) capacitor c=0.00179496f \
 //x=15.385 //y=5.02 //x2=16.535 //y2=4.44
cc_1771 ( N_VDD_c_1085_p N_CLK_c_6057_n ) capacitor c=0.00146064f //x=95.83 \
 //y=7.4 //x2=7.145 //y2=4.44
cc_1772 ( N_VDD_c_1085_p N_CLK_c_6058_n ) capacitor c=0.0974885f //x=95.83 \
 //y=7.4 //x2=35.775 //y2=4.44
cc_1773 ( N_VDD_c_1368_p N_CLK_c_6058_n ) capacitor c=0.00258496f //x=19.07 \
 //y=7.4 //x2=35.775 //y2=4.44
cc_1774 ( N_VDD_c_1796_p N_CLK_c_6058_n ) capacitor c=0.00328994f //x=20.245 \
 //y=7.4 //x2=35.775 //y2=4.44
cc_1775 ( N_VDD_c_1195_p N_CLK_c_6058_n ) capacitor c=0.00135925f //x=21.125 \
 //y=7.4 //x2=35.775 //y2=4.44
cc_1776 ( N_VDD_c_1068_n N_CLK_c_6058_n ) capacitor c=0.0389825f //x=19.24 \
 //y=7.4 //x2=35.775 //y2=4.44
cc_1777 ( N_VDD_c_1069_n N_CLK_c_6058_n ) capacitor c=0.0263454f //x=24.05 \
 //y=7.4 //x2=35.775 //y2=4.44
cc_1778 ( N_VDD_c_1070_n N_CLK_c_6058_n ) capacitor c=0.0263454f //x=28.86 \
 //y=7.4 //x2=35.775 //y2=4.44
cc_1779 ( N_VDD_c_1071_n N_CLK_c_6058_n ) capacitor c=0.0263454f //x=33.67 \
 //y=7.4 //x2=35.775 //y2=4.44
cc_1780 ( N_VDD_M84_noxref_s N_CLK_c_6058_n ) capacitor c=0.00179496f \
 //x=20.195 //y=5.02 //x2=35.775 //y2=4.44
cc_1781 ( N_VDD_c_1085_p N_CLK_c_6067_n ) capacitor c=0.00120845f //x=95.83 \
 //y=7.4 //x2=16.765 //y2=4.44
cc_1782 ( N_VDD_c_1072_n N_CLK_c_6068_n ) capacitor c=0.0263454f //x=38.48 \
 //y=7.4 //x2=45.395 //y2=4.44
cc_1783 ( N_VDD_c_1073_n N_CLK_c_6068_n ) capacitor c=0.0263454f //x=43.29 \
 //y=7.4 //x2=45.395 //y2=4.44
cc_1784 ( N_VDD_c_1074_n N_CLK_c_6070_n ) capacitor c=0.0263454f //x=48.1 \
 //y=7.4 //x2=64.635 //y2=4.44
cc_1785 ( N_VDD_c_1075_n N_CLK_c_6070_n ) capacitor c=0.0263454f //x=52.91 \
 //y=7.4 //x2=64.635 //y2=4.44
cc_1786 ( N_VDD_c_1076_n N_CLK_c_6070_n ) capacitor c=0.0263454f //x=57.72 \
 //y=7.4 //x2=64.635 //y2=4.44
cc_1787 ( N_VDD_c_1077_n N_CLK_c_6070_n ) capacitor c=0.0249242f //x=62.53 \
 //y=7.4 //x2=64.635 //y2=4.44
cc_1788 ( N_VDD_c_1078_n N_CLK_c_6074_n ) capacitor c=0.0263454f //x=67.34 \
 //y=7.4 //x2=74.255 //y2=4.44
cc_1789 ( N_VDD_c_1079_n N_CLK_c_6074_n ) capacitor c=0.0263454f //x=72.15 \
 //y=7.4 //x2=74.255 //y2=4.44
cc_1790 ( N_VDD_c_1085_p N_CLK_c_6040_n ) capacitor c=2.03287e-19 //x=95.83 \
 //y=7.4 //x2=7.03 //y2=2.08
cc_1791 ( N_VDD_c_1065_n N_CLK_c_6040_n ) capacitor c=8.47879e-19 //x=4.81 \
 //y=7.4 //x2=7.03 //y2=2.08
cc_1792 ( N_VDD_c_1085_p N_CLK_c_6041_n ) capacitor c=2.03287e-19 //x=95.83 \
 //y=7.4 //x2=16.65 //y2=2.08
cc_1793 ( N_VDD_c_1067_n N_CLK_c_6041_n ) capacitor c=6.15921e-19 //x=14.43 \
 //y=7.4 //x2=16.65 //y2=2.08
cc_1794 ( N_VDD_c_1071_n N_CLK_c_6042_n ) capacitor c=4.26258e-19 //x=33.67 \
 //y=7.4 //x2=35.89 //y2=2.08
cc_1795 ( N_VDD_c_1073_n N_CLK_c_6043_n ) capacitor c=4.26258e-19 //x=43.29 \
 //y=7.4 //x2=45.51 //y2=2.08
cc_1796 ( N_VDD_c_1077_n N_CLK_c_6044_n ) capacitor c=5.01735e-19 //x=62.53 \
 //y=7.4 //x2=64.75 //y2=2.08
cc_1797 ( N_VDD_c_1079_n N_CLK_c_6045_n ) capacitor c=4.23657e-19 //x=72.15 \
 //y=7.4 //x2=74.37 //y2=2.08
cc_1798 ( N_VDD_c_1175_p N_CLK_M68_noxref_g ) capacitor c=0.00676195f \
 //x=7.575 //y=7.4 //x2=7 //y2=6.02
cc_1799 ( N_VDD_M67_noxref_d N_CLK_M68_noxref_g ) capacitor c=0.015318f \
 //x=6.635 //y=5.02 //x2=7 //y2=6.02
cc_1800 ( N_VDD_c_1175_p N_CLK_M69_noxref_g ) capacitor c=0.00675175f \
 //x=7.575 //y=7.4 //x2=7.44 //y2=6.02
cc_1801 ( N_VDD_M69_noxref_d N_CLK_M69_noxref_g ) capacitor c=0.015318f \
 //x=7.515 //y=5.02 //x2=7.44 //y2=6.02
cc_1802 ( N_VDD_c_1358_p N_CLK_M80_noxref_g ) capacitor c=0.00676195f \
 //x=17.195 //y=7.4 //x2=16.62 //y2=6.02
cc_1803 ( N_VDD_M79_noxref_d N_CLK_M80_noxref_g ) capacitor c=0.015318f \
 //x=16.255 //y=5.02 //x2=16.62 //y2=6.02
cc_1804 ( N_VDD_c_1358_p N_CLK_M81_noxref_g ) capacitor c=0.00675175f \
 //x=17.195 //y=7.4 //x2=17.06 //y2=6.02
cc_1805 ( N_VDD_M81_noxref_d N_CLK_M81_noxref_g ) capacitor c=0.015318f \
 //x=17.135 //y=5.02 //x2=17.06 //y2=6.02
cc_1806 ( N_VDD_c_1524_p N_CLK_M104_noxref_g ) capacitor c=0.00676195f \
 //x=36.435 //y=7.4 //x2=35.86 //y2=6.02
cc_1807 ( N_VDD_M103_noxref_d N_CLK_M104_noxref_g ) capacitor c=0.015318f \
 //x=35.495 //y=5.02 //x2=35.86 //y2=6.02
cc_1808 ( N_VDD_c_1524_p N_CLK_M105_noxref_g ) capacitor c=0.00675175f \
 //x=36.435 //y=7.4 //x2=36.3 //y2=6.02
cc_1809 ( N_VDD_M105_noxref_d N_CLK_M105_noxref_g ) capacitor c=0.015318f \
 //x=36.375 //y=5.02 //x2=36.3 //y2=6.02
cc_1810 ( N_VDD_c_1569_p N_CLK_M116_noxref_g ) capacitor c=0.00676195f \
 //x=46.055 //y=7.4 //x2=45.48 //y2=6.02
cc_1811 ( N_VDD_M115_noxref_d N_CLK_M116_noxref_g ) capacitor c=0.015318f \
 //x=45.115 //y=5.02 //x2=45.48 //y2=6.02
cc_1812 ( N_VDD_c_1569_p N_CLK_M117_noxref_g ) capacitor c=0.00675175f \
 //x=46.055 //y=7.4 //x2=45.92 //y2=6.02
cc_1813 ( N_VDD_M117_noxref_d N_CLK_M117_noxref_g ) capacitor c=0.015318f \
 //x=45.995 //y=5.02 //x2=45.92 //y2=6.02
cc_1814 ( N_VDD_c_1836_p N_CLK_M140_noxref_g ) capacitor c=0.00676195f \
 //x=65.295 //y=7.4 //x2=64.72 //y2=6.02
cc_1815 ( N_VDD_M139_noxref_d N_CLK_M140_noxref_g ) capacitor c=0.015318f \
 //x=64.355 //y=5.02 //x2=64.72 //y2=6.02
cc_1816 ( N_VDD_c_1836_p N_CLK_M141_noxref_g ) capacitor c=0.00675175f \
 //x=65.295 //y=7.4 //x2=65.16 //y2=6.02
cc_1817 ( N_VDD_M141_noxref_d N_CLK_M141_noxref_g ) capacitor c=0.015318f \
 //x=65.235 //y=5.02 //x2=65.16 //y2=6.02
cc_1818 ( N_VDD_c_1840_p N_CLK_M152_noxref_g ) capacitor c=0.00676195f \
 //x=74.915 //y=7.4 //x2=74.34 //y2=6.02
cc_1819 ( N_VDD_M151_noxref_d N_CLK_M152_noxref_g ) capacitor c=0.015318f \
 //x=73.975 //y=5.02 //x2=74.34 //y2=6.02
cc_1820 ( N_VDD_c_1840_p N_CLK_M153_noxref_g ) capacitor c=0.00675175f \
 //x=74.915 //y=7.4 //x2=74.78 //y2=6.02
cc_1821 ( N_VDD_M153_noxref_d N_CLK_M153_noxref_g ) capacitor c=0.015318f \
 //x=74.855 //y=5.02 //x2=74.78 //y2=6.02
cc_1822 ( N_VDD_c_1077_n N_noxref_18_c_6747_n ) capacitor c=5.22311e-19 \
 //x=62.53 //y=7.4 //x2=61.05 //y2=2.08
cc_1823 ( N_VDD_c_1085_p N_noxref_18_c_6762_n ) capacitor c=0.00437246f \
 //x=95.83 //y=7.4 //x2=64.855 //y2=5.155
cc_1824 ( N_VDD_c_1243_p N_noxref_18_c_6762_n ) capacitor c=4.31596e-19 \
 //x=64.415 //y=7.4 //x2=64.855 //y2=5.155
cc_1825 ( N_VDD_c_1836_p N_noxref_18_c_6762_n ) capacitor c=4.31596e-19 \
 //x=65.295 //y=7.4 //x2=64.855 //y2=5.155
cc_1826 ( N_VDD_M139_noxref_d N_noxref_18_c_6762_n ) capacitor c=0.0109802f \
 //x=64.355 //y=5.02 //x2=64.855 //y2=5.155
cc_1827 ( N_VDD_c_1077_n N_noxref_18_c_6766_n ) capacitor c=0.00863585f \
 //x=62.53 //y=7.4 //x2=64.145 //y2=5.155
cc_1828 ( N_VDD_M138_noxref_s N_noxref_18_c_6766_n ) capacitor c=0.0831083f \
 //x=63.485 //y=5.02 //x2=64.145 //y2=5.155
cc_1829 ( N_VDD_c_1085_p N_noxref_18_c_6768_n ) capacitor c=0.00434259f \
 //x=95.83 //y=7.4 //x2=65.735 //y2=5.155
cc_1830 ( N_VDD_c_1836_p N_noxref_18_c_6768_n ) capacitor c=4.31596e-19 \
 //x=65.295 //y=7.4 //x2=65.735 //y2=5.155
cc_1831 ( N_VDD_c_1853_p N_noxref_18_c_6768_n ) capacitor c=4.31596e-19 \
 //x=66.175 //y=7.4 //x2=65.735 //y2=5.155
cc_1832 ( N_VDD_M141_noxref_d N_noxref_18_c_6768_n ) capacitor c=0.0109802f \
 //x=65.235 //y=5.02 //x2=65.735 //y2=5.155
cc_1833 ( N_VDD_c_1085_p N_noxref_18_c_6772_n ) capacitor c=0.00424413f \
 //x=95.83 //y=7.4 //x2=66.515 //y2=5.155
cc_1834 ( N_VDD_c_1853_p N_noxref_18_c_6772_n ) capacitor c=7.45454e-19 \
 //x=66.175 //y=7.4 //x2=66.515 //y2=5.155
cc_1835 ( N_VDD_c_1244_p N_noxref_18_c_6772_n ) capacitor c=0.00198097f \
 //x=67.17 //y=7.4 //x2=66.515 //y2=5.155
cc_1836 ( N_VDD_M143_noxref_d N_noxref_18_c_6772_n ) capacitor c=0.0109802f \
 //x=66.115 //y=5.02 //x2=66.515 //y2=5.155
cc_1837 ( N_VDD_c_1078_n N_noxref_18_c_6776_n ) capacitor c=0.0400668f \
 //x=67.34 //y=7.4 //x2=66.6 //y2=3.33
cc_1838 ( N_VDD_c_1085_p N_noxref_18_c_6749_n ) capacitor c=9.10347e-19 \
 //x=95.83 //y=7.4 //x2=78.07 //y2=2.08
cc_1839 ( N_VDD_c_1080_n N_noxref_18_c_6749_n ) capacitor c=0.0133494f \
 //x=76.96 //y=7.4 //x2=78.07 //y2=2.08
cc_1840 ( N_VDD_M156_noxref_s N_noxref_18_c_6749_n ) capacitor c=0.0125322f \
 //x=77.915 //y=5.02 //x2=78.07 //y2=2.08
cc_1841 ( N_VDD_c_1703_p N_noxref_18_M136_noxref_g ) capacitor c=0.00675175f \
 //x=61.365 //y=7.4 //x2=60.79 //y2=6.02
cc_1842 ( N_VDD_M135_noxref_d N_noxref_18_M136_noxref_g ) capacitor \
 c=0.015318f //x=60.425 //y=5.02 //x2=60.79 //y2=6.02
cc_1843 ( N_VDD_c_1703_p N_noxref_18_M137_noxref_g ) capacitor c=0.00675379f \
 //x=61.365 //y=7.4 //x2=61.23 //y2=6.02
cc_1844 ( N_VDD_M137_noxref_d N_noxref_18_M137_noxref_g ) capacitor \
 c=0.0394719f //x=61.305 //y=5.02 //x2=61.23 //y2=6.02
cc_1845 ( N_VDD_c_1278_p N_noxref_18_M156_noxref_g ) capacitor c=0.00749687f \
 //x=78.845 //y=7.4 //x2=78.27 //y2=6.02
cc_1846 ( N_VDD_M156_noxref_s N_noxref_18_M156_noxref_g ) capacitor \
 c=0.0477201f //x=77.915 //y=5.02 //x2=78.27 //y2=6.02
cc_1847 ( N_VDD_c_1278_p N_noxref_18_M157_noxref_g ) capacitor c=0.00675175f \
 //x=78.845 //y=7.4 //x2=78.71 //y2=6.02
cc_1848 ( N_VDD_M157_noxref_d N_noxref_18_M157_noxref_g ) capacitor \
 c=0.015318f //x=78.785 //y=5.02 //x2=78.71 //y2=6.02
cc_1849 ( N_VDD_c_1080_n N_noxref_18_c_6788_n ) capacitor c=0.0057745f \
 //x=76.96 //y=7.4 //x2=78.345 //y2=4.79
cc_1850 ( N_VDD_M156_noxref_s N_noxref_18_c_6788_n ) capacitor c=0.00444914f \
 //x=77.915 //y=5.02 //x2=78.345 //y2=4.79
cc_1851 ( N_VDD_c_1085_p N_noxref_18_M138_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=63.915 //y2=5.02
cc_1852 ( N_VDD_c_1243_p N_noxref_18_M138_noxref_d ) capacitor c=0.0139598f \
 //x=64.415 //y=7.4 //x2=63.915 //y2=5.02
cc_1853 ( N_VDD_M139_noxref_d N_noxref_18_M138_noxref_d ) capacitor \
 c=0.0664752f //x=64.355 //y=5.02 //x2=63.915 //y2=5.02
cc_1854 ( N_VDD_c_1085_p N_noxref_18_M140_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=64.795 //y2=5.02
cc_1855 ( N_VDD_c_1836_p N_noxref_18_M140_noxref_d ) capacitor c=0.0139598f \
 //x=65.295 //y=7.4 //x2=64.795 //y2=5.02
cc_1856 ( N_VDD_c_1078_n N_noxref_18_M140_noxref_d ) capacitor c=4.9285e-19 \
 //x=67.34 //y=7.4 //x2=64.795 //y2=5.02
cc_1857 ( N_VDD_M138_noxref_s N_noxref_18_M140_noxref_d ) capacitor \
 c=0.00130656f //x=63.485 //y=5.02 //x2=64.795 //y2=5.02
cc_1858 ( N_VDD_M139_noxref_d N_noxref_18_M140_noxref_d ) capacitor \
 c=0.0664752f //x=64.355 //y=5.02 //x2=64.795 //y2=5.02
cc_1859 ( N_VDD_M141_noxref_d N_noxref_18_M140_noxref_d ) capacitor \
 c=0.0664752f //x=65.235 //y=5.02 //x2=64.795 //y2=5.02
cc_1860 ( N_VDD_c_1085_p N_noxref_18_M142_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=65.675 //y2=5.02
cc_1861 ( N_VDD_c_1853_p N_noxref_18_M142_noxref_d ) capacitor c=0.0139598f \
 //x=66.175 //y=7.4 //x2=65.675 //y2=5.02
cc_1862 ( N_VDD_c_1078_n N_noxref_18_M142_noxref_d ) capacitor c=0.00939849f \
 //x=67.34 //y=7.4 //x2=65.675 //y2=5.02
cc_1863 ( N_VDD_M141_noxref_d N_noxref_18_M142_noxref_d ) capacitor \
 c=0.0664752f //x=65.235 //y=5.02 //x2=65.675 //y2=5.02
cc_1864 ( N_VDD_M143_noxref_d N_noxref_18_M142_noxref_d ) capacitor \
 c=0.0664752f //x=66.115 //y=5.02 //x2=65.675 //y2=5.02
cc_1865 ( N_VDD_M144_noxref_s N_noxref_18_M142_noxref_d ) capacitor \
 c=3.57641e-19 //x=68.295 //y=5.02 //x2=65.675 //y2=5.02
cc_1866 ( N_VDD_c_1085_p N_RN_c_7088_n ) capacitor c=2.05828e-19 //x=95.83 \
 //y=7.4 //x2=2.22 //y2=2.08
cc_1867 ( N_VDD_c_1063_n N_RN_c_7088_n ) capacitor c=8.08669e-19 //x=0.74 \
 //y=7.4 //x2=2.22 //y2=2.08
cc_1868 ( N_VDD_c_1068_n N_RN_c_7089_n ) capacitor c=6.58823e-19 //x=19.24 \
 //y=7.4 //x2=17.76 //y2=2.08
cc_1869 ( N_VDD_c_1085_p N_RN_c_7090_n ) capacitor c=2.03486e-19 //x=95.83 \
 //y=7.4 //x2=21.46 //y2=2.08
cc_1870 ( N_VDD_c_1068_n N_RN_c_7090_n ) capacitor c=5.89117e-19 //x=19.24 \
 //y=7.4 //x2=21.46 //y2=2.08
cc_1871 ( N_VDD_c_1070_n N_RN_c_7091_n ) capacitor c=4.48671e-19 //x=28.86 \
 //y=7.4 //x2=31.08 //y2=2.08
cc_1872 ( N_VDD_c_1074_n N_RN_c_7092_n ) capacitor c=5.43708e-19 //x=48.1 \
 //y=7.4 //x2=46.62 //y2=2.08
cc_1873 ( N_VDD_c_1074_n N_RN_c_7093_n ) capacitor c=3.99454e-19 //x=48.1 \
 //y=7.4 //x2=50.32 //y2=2.08
cc_1874 ( N_VDD_c_1076_n N_RN_c_7094_n ) capacitor c=4.96201e-19 //x=57.72 \
 //y=7.4 //x2=59.94 //y2=2.08
cc_1875 ( N_VDD_c_1080_n N_RN_c_7095_n ) capacitor c=0.00108383f //x=76.96 \
 //y=7.4 //x2=75.48 //y2=2.08
cc_1876 ( N_VDD_c_1085_p N_RN_c_7096_n ) capacitor c=2.03486e-19 //x=95.83 \
 //y=7.4 //x2=79.18 //y2=2.08
cc_1877 ( N_VDD_c_1080_n N_RN_c_7096_n ) capacitor c=5.89117e-19 //x=76.96 \
 //y=7.4 //x2=79.18 //y2=2.08
cc_1878 ( N_VDD_c_1087_p N_RN_M62_noxref_g ) capacitor c=0.00676195f //x=2.765 \
 //y=7.4 //x2=2.19 //y2=6.02
cc_1879 ( N_VDD_M61_noxref_d N_RN_M62_noxref_g ) capacitor c=0.015318f \
 //x=1.825 //y=5.02 //x2=2.19 //y2=6.02
cc_1880 ( N_VDD_c_1087_p N_RN_M63_noxref_g ) capacitor c=0.00675175f //x=2.765 \
 //y=7.4 //x2=2.63 //y2=6.02
cc_1881 ( N_VDD_M63_noxref_d N_RN_M63_noxref_g ) capacitor c=0.015318f \
 //x=2.705 //y=5.02 //x2=2.63 //y2=6.02
cc_1882 ( N_VDD_c_1364_p N_RN_M82_noxref_g ) capacitor c=0.00675175f \
 //x=18.075 //y=7.4 //x2=17.5 //y2=6.02
cc_1883 ( N_VDD_M81_noxref_d N_RN_M82_noxref_g ) capacitor c=0.015318f \
 //x=17.135 //y=5.02 //x2=17.5 //y2=6.02
cc_1884 ( N_VDD_c_1364_p N_RN_M83_noxref_g ) capacitor c=0.00675379f \
 //x=18.075 //y=7.4 //x2=17.94 //y2=6.02
cc_1885 ( N_VDD_M83_noxref_d N_RN_M83_noxref_g ) capacitor c=0.0394719f \
 //x=18.015 //y=5.02 //x2=17.94 //y2=6.02
cc_1886 ( N_VDD_c_1300_p N_RN_M86_noxref_g ) capacitor c=0.00676195f \
 //x=22.005 //y=7.4 //x2=21.43 //y2=6.02
cc_1887 ( N_VDD_M85_noxref_d N_RN_M86_noxref_g ) capacitor c=0.015318f \
 //x=21.065 //y=5.02 //x2=21.43 //y2=6.02
cc_1888 ( N_VDD_c_1300_p N_RN_M87_noxref_g ) capacitor c=0.00675175f \
 //x=22.005 //y=7.4 //x2=21.87 //y2=6.02
cc_1889 ( N_VDD_M87_noxref_d N_RN_M87_noxref_g ) capacitor c=0.015318f \
 //x=21.945 //y=5.02 //x2=21.87 //y2=6.02
cc_1890 ( N_VDD_c_1436_p N_RN_M98_noxref_g ) capacitor c=0.00676195f \
 //x=31.625 //y=7.4 //x2=31.05 //y2=6.02
cc_1891 ( N_VDD_M97_noxref_d N_RN_M98_noxref_g ) capacitor c=0.015318f \
 //x=30.685 //y=5.02 //x2=31.05 //y2=6.02
cc_1892 ( N_VDD_c_1436_p N_RN_M99_noxref_g ) capacitor c=0.00675175f \
 //x=31.625 //y=7.4 //x2=31.49 //y2=6.02
cc_1893 ( N_VDD_M99_noxref_d N_RN_M99_noxref_g ) capacitor c=0.015318f \
 //x=31.565 //y=5.02 //x2=31.49 //y2=6.02
cc_1894 ( N_VDD_c_1575_p N_RN_M118_noxref_g ) capacitor c=0.00675175f \
 //x=46.935 //y=7.4 //x2=46.36 //y2=6.02
cc_1895 ( N_VDD_M117_noxref_d N_RN_M118_noxref_g ) capacitor c=0.015318f \
 //x=45.995 //y=5.02 //x2=46.36 //y2=6.02
cc_1896 ( N_VDD_c_1575_p N_RN_M119_noxref_g ) capacitor c=0.00675379f \
 //x=46.935 //y=7.4 //x2=46.8 //y2=6.02
cc_1897 ( N_VDD_M119_noxref_d N_RN_M119_noxref_g ) capacitor c=0.0394719f \
 //x=46.875 //y=5.02 //x2=46.8 //y2=6.02
cc_1898 ( N_VDD_c_1920_p N_RN_M122_noxref_g ) capacitor c=0.00676195f \
 //x=50.865 //y=7.4 //x2=50.29 //y2=6.02
cc_1899 ( N_VDD_M121_noxref_d N_RN_M122_noxref_g ) capacitor c=0.015318f \
 //x=49.925 //y=5.02 //x2=50.29 //y2=6.02
cc_1900 ( N_VDD_c_1920_p N_RN_M123_noxref_g ) capacitor c=0.00675175f \
 //x=50.865 //y=7.4 //x2=50.73 //y2=6.02
cc_1901 ( N_VDD_M123_noxref_d N_RN_M123_noxref_g ) capacitor c=0.015318f \
 //x=50.805 //y=5.02 //x2=50.73 //y2=6.02
cc_1902 ( N_VDD_c_1697_p N_RN_M134_noxref_g ) capacitor c=0.00676195f \
 //x=60.485 //y=7.4 //x2=59.91 //y2=6.02
cc_1903 ( N_VDD_M133_noxref_d N_RN_M134_noxref_g ) capacitor c=0.015318f \
 //x=59.545 //y=5.02 //x2=59.91 //y2=6.02
cc_1904 ( N_VDD_c_1697_p N_RN_M135_noxref_g ) capacitor c=0.00675175f \
 //x=60.485 //y=7.4 //x2=60.35 //y2=6.02
cc_1905 ( N_VDD_M135_noxref_d N_RN_M135_noxref_g ) capacitor c=0.015318f \
 //x=60.425 //y=5.02 //x2=60.35 //y2=6.02
cc_1906 ( N_VDD_c_1928_p N_RN_M154_noxref_g ) capacitor c=0.00675175f \
 //x=75.795 //y=7.4 //x2=75.22 //y2=6.02
cc_1907 ( N_VDD_M153_noxref_d N_RN_M154_noxref_g ) capacitor c=0.015318f \
 //x=74.855 //y=5.02 //x2=75.22 //y2=6.02
cc_1908 ( N_VDD_c_1928_p N_RN_M155_noxref_g ) capacitor c=0.00675379f \
 //x=75.795 //y=7.4 //x2=75.66 //y2=6.02
cc_1909 ( N_VDD_M155_noxref_d N_RN_M155_noxref_g ) capacitor c=0.0394719f \
 //x=75.735 //y=5.02 //x2=75.66 //y2=6.02
cc_1910 ( N_VDD_c_1932_p N_RN_M158_noxref_g ) capacitor c=0.00676195f \
 //x=79.725 //y=7.4 //x2=79.15 //y2=6.02
cc_1911 ( N_VDD_M157_noxref_d N_RN_M158_noxref_g ) capacitor c=0.015318f \
 //x=78.785 //y=5.02 //x2=79.15 //y2=6.02
cc_1912 ( N_VDD_c_1932_p N_RN_M159_noxref_g ) capacitor c=0.00675175f \
 //x=79.725 //y=7.4 //x2=79.59 //y2=6.02
cc_1913 ( N_VDD_M159_noxref_d N_RN_M159_noxref_g ) capacitor c=0.015318f \
 //x=79.665 //y=5.02 //x2=79.59 //y2=6.02
cc_1914 ( N_VDD_c_1085_p N_SN_c_8145_n ) capacitor c=2.03486e-19 //x=95.83 \
 //y=7.4 //x2=11.84 //y2=2.08
cc_1915 ( N_VDD_c_1066_n N_SN_c_8145_n ) capacitor c=5.89117e-19 //x=9.62 \
 //y=7.4 //x2=11.84 //y2=2.08
cc_1916 ( N_VDD_c_1069_n N_SN_c_8146_n ) capacitor c=3.99454e-19 //x=24.05 \
 //y=7.4 //x2=26.27 //y2=2.08
cc_1917 ( N_VDD_c_1072_n N_SN_c_8147_n ) capacitor c=3.99454e-19 //x=38.48 \
 //y=7.4 //x2=40.7 //y2=2.08
cc_1918 ( N_VDD_c_1075_n N_SN_c_8148_n ) capacitor c=3.99454e-19 //x=52.91 \
 //y=7.4 //x2=55.13 //y2=2.08
cc_1919 ( N_VDD_c_1078_n N_SN_c_8149_n ) capacitor c=3.99454e-19 //x=67.34 \
 //y=7.4 //x2=69.56 //y2=2.08
cc_1920 ( N_VDD_c_1085_p N_SN_c_8150_n ) capacitor c=2.03486e-19 //x=95.83 \
 //y=7.4 //x2=83.99 //y2=2.08
cc_1921 ( N_VDD_c_1081_n N_SN_c_8150_n ) capacitor c=5.89117e-19 //x=81.77 \
 //y=7.4 //x2=83.99 //y2=2.08
cc_1922 ( N_VDD_c_1135_p N_SN_M74_noxref_g ) capacitor c=0.00676195f \
 //x=12.385 //y=7.4 //x2=11.81 //y2=6.02
cc_1923 ( N_VDD_M73_noxref_d N_SN_M74_noxref_g ) capacitor c=0.015318f \
 //x=11.445 //y=5.02 //x2=11.81 //y2=6.02
cc_1924 ( N_VDD_c_1135_p N_SN_M75_noxref_g ) capacitor c=0.00675175f \
 //x=12.385 //y=7.4 //x2=12.25 //y2=6.02
cc_1925 ( N_VDD_M75_noxref_d N_SN_M75_noxref_g ) capacitor c=0.015318f \
 //x=12.325 //y=5.02 //x2=12.25 //y2=6.02
cc_1926 ( N_VDD_c_1402_p N_SN_M92_noxref_g ) capacitor c=0.00676195f \
 //x=26.815 //y=7.4 //x2=26.24 //y2=6.02
cc_1927 ( N_VDD_M91_noxref_d N_SN_M92_noxref_g ) capacitor c=0.015318f \
 //x=25.875 //y=5.02 //x2=26.24 //y2=6.02
cc_1928 ( N_VDD_c_1402_p N_SN_M93_noxref_g ) capacitor c=0.00675175f \
 //x=26.815 //y=7.4 //x2=26.68 //y2=6.02
cc_1929 ( N_VDD_M93_noxref_d N_SN_M93_noxref_g ) capacitor c=0.015318f \
 //x=26.755 //y=5.02 //x2=26.68 //y2=6.02
cc_1930 ( N_VDD_c_1484_p N_SN_M110_noxref_g ) capacitor c=0.00676195f \
 //x=41.245 //y=7.4 //x2=40.67 //y2=6.02
cc_1931 ( N_VDD_M109_noxref_d N_SN_M110_noxref_g ) capacitor c=0.015318f \
 //x=40.305 //y=5.02 //x2=40.67 //y2=6.02
cc_1932 ( N_VDD_c_1484_p N_SN_M111_noxref_g ) capacitor c=0.00675175f \
 //x=41.245 //y=7.4 //x2=41.11 //y2=6.02
cc_1933 ( N_VDD_M111_noxref_d N_SN_M111_noxref_g ) capacitor c=0.015318f \
 //x=41.185 //y=5.02 //x2=41.11 //y2=6.02
cc_1934 ( N_VDD_c_1613_p N_SN_M128_noxref_g ) capacitor c=0.00676195f \
 //x=55.675 //y=7.4 //x2=55.1 //y2=6.02
cc_1935 ( N_VDD_M127_noxref_d N_SN_M128_noxref_g ) capacitor c=0.015318f \
 //x=54.735 //y=5.02 //x2=55.1 //y2=6.02
cc_1936 ( N_VDD_c_1613_p N_SN_M129_noxref_g ) capacitor c=0.00675175f \
 //x=55.675 //y=7.4 //x2=55.54 //y2=6.02
cc_1937 ( N_VDD_M129_noxref_d N_SN_M129_noxref_g ) capacitor c=0.015318f \
 //x=55.615 //y=5.02 //x2=55.54 //y2=6.02
cc_1938 ( N_VDD_c_1745_p N_SN_M146_noxref_g ) capacitor c=0.00676195f \
 //x=70.105 //y=7.4 //x2=69.53 //y2=6.02
cc_1939 ( N_VDD_M145_noxref_d N_SN_M146_noxref_g ) capacitor c=0.015318f \
 //x=69.165 //y=5.02 //x2=69.53 //y2=6.02
cc_1940 ( N_VDD_c_1745_p N_SN_M147_noxref_g ) capacitor c=0.00675175f \
 //x=70.105 //y=7.4 //x2=69.97 //y2=6.02
cc_1941 ( N_VDD_M147_noxref_d N_SN_M147_noxref_g ) capacitor c=0.015318f \
 //x=70.045 //y=5.02 //x2=69.97 //y2=6.02
cc_1942 ( N_VDD_c_1964_p N_SN_M164_noxref_g ) capacitor c=0.00676195f \
 //x=84.535 //y=7.4 //x2=83.96 //y2=6.02
cc_1943 ( N_VDD_M163_noxref_d N_SN_M164_noxref_g ) capacitor c=0.015318f \
 //x=83.595 //y=5.02 //x2=83.96 //y2=6.02
cc_1944 ( N_VDD_c_1964_p N_SN_M165_noxref_g ) capacitor c=0.00675175f \
 //x=84.535 //y=7.4 //x2=84.4 //y2=6.02
cc_1945 ( N_VDD_M165_noxref_d N_SN_M165_noxref_g ) capacitor c=0.015318f \
 //x=84.475 //y=5.02 //x2=84.4 //y2=6.02
cc_1946 ( N_VDD_c_1078_n N_noxref_21_c_8828_n ) capacitor c=5.43708e-19 \
 //x=67.34 //y=7.4 //x2=65.86 //y2=2.08
cc_1947 ( N_VDD_c_1079_n N_noxref_21_c_8829_n ) capacitor c=4.57708e-19 \
 //x=72.15 //y=7.4 //x2=70.67 //y2=2.08
cc_1948 ( N_VDD_c_1085_p N_noxref_21_c_8835_n ) capacitor c=0.00437246f \
 //x=95.83 //y=7.4 //x2=74.475 //y2=5.155
cc_1949 ( N_VDD_c_1249_p N_noxref_21_c_8835_n ) capacitor c=4.31596e-19 \
 //x=74.035 //y=7.4 //x2=74.475 //y2=5.155
cc_1950 ( N_VDD_c_1840_p N_noxref_21_c_8835_n ) capacitor c=4.31596e-19 \
 //x=74.915 //y=7.4 //x2=74.475 //y2=5.155
cc_1951 ( N_VDD_M151_noxref_d N_noxref_21_c_8835_n ) capacitor c=0.0109802f \
 //x=73.975 //y=5.02 //x2=74.475 //y2=5.155
cc_1952 ( N_VDD_c_1079_n N_noxref_21_c_8839_n ) capacitor c=0.00863585f \
 //x=72.15 //y=7.4 //x2=73.765 //y2=5.155
cc_1953 ( N_VDD_M150_noxref_s N_noxref_21_c_8839_n ) capacitor c=0.0831083f \
 //x=73.105 //y=5.02 //x2=73.765 //y2=5.155
cc_1954 ( N_VDD_c_1085_p N_noxref_21_c_8841_n ) capacitor c=0.00435431f \
 //x=95.83 //y=7.4 //x2=75.355 //y2=5.155
cc_1955 ( N_VDD_c_1840_p N_noxref_21_c_8841_n ) capacitor c=4.31596e-19 \
 //x=74.915 //y=7.4 //x2=75.355 //y2=5.155
cc_1956 ( N_VDD_c_1928_p N_noxref_21_c_8841_n ) capacitor c=4.31764e-19 \
 //x=75.795 //y=7.4 //x2=75.355 //y2=5.155
cc_1957 ( N_VDD_M153_noxref_d N_noxref_21_c_8841_n ) capacitor c=0.0109802f \
 //x=74.855 //y=5.02 //x2=75.355 //y2=5.155
cc_1958 ( N_VDD_c_1085_p N_noxref_21_c_8845_n ) capacitor c=0.00434174f \
 //x=95.83 //y=7.4 //x2=76.135 //y2=5.155
cc_1959 ( N_VDD_c_1928_p N_noxref_21_c_8845_n ) capacitor c=7.46626e-19 \
 //x=75.795 //y=7.4 //x2=76.135 //y2=5.155
cc_1960 ( N_VDD_c_1276_p N_noxref_21_c_8845_n ) capacitor c=0.00198565f \
 //x=76.79 //y=7.4 //x2=76.135 //y2=5.155
cc_1961 ( N_VDD_M155_noxref_d N_noxref_21_c_8845_n ) capacitor c=0.0112985f \
 //x=75.735 //y=5.02 //x2=76.135 //y2=5.155
cc_1962 ( N_VDD_c_1080_n N_noxref_21_c_8849_n ) capacitor c=0.0420055f \
 //x=76.96 //y=7.4 //x2=76.22 //y2=3.7
cc_1963 ( N_VDD_c_1082_n N_noxref_21_c_8831_n ) capacitor c=6.56791e-19 \
 //x=86.58 //y=7.4 //x2=85.1 //y2=2.08
cc_1964 ( N_VDD_c_1853_p N_noxref_21_M142_noxref_g ) capacitor c=0.00675175f \
 //x=66.175 //y=7.4 //x2=65.6 //y2=6.02
cc_1965 ( N_VDD_M141_noxref_d N_noxref_21_M142_noxref_g ) capacitor \
 c=0.015318f //x=65.235 //y=5.02 //x2=65.6 //y2=6.02
cc_1966 ( N_VDD_c_1853_p N_noxref_21_M143_noxref_g ) capacitor c=0.00675379f \
 //x=66.175 //y=7.4 //x2=66.04 //y2=6.02
cc_1967 ( N_VDD_M143_noxref_d N_noxref_21_M143_noxref_g ) capacitor \
 c=0.0394719f //x=66.115 //y=5.02 //x2=66.04 //y2=6.02
cc_1968 ( N_VDD_c_1751_p N_noxref_21_M148_noxref_g ) capacitor c=0.00675175f \
 //x=70.985 //y=7.4 //x2=70.41 //y2=6.02
cc_1969 ( N_VDD_M147_noxref_d N_noxref_21_M148_noxref_g ) capacitor \
 c=0.015318f //x=70.045 //y=5.02 //x2=70.41 //y2=6.02
cc_1970 ( N_VDD_c_1751_p N_noxref_21_M149_noxref_g ) capacitor c=0.00675379f \
 //x=70.985 //y=7.4 //x2=70.85 //y2=6.02
cc_1971 ( N_VDD_M149_noxref_d N_noxref_21_M149_noxref_g ) capacitor \
 c=0.0394719f //x=70.925 //y=5.02 //x2=70.85 //y2=6.02
cc_1972 ( N_VDD_c_1994_p N_noxref_21_M166_noxref_g ) capacitor c=0.00675175f \
 //x=85.415 //y=7.4 //x2=84.84 //y2=6.02
cc_1973 ( N_VDD_M165_noxref_d N_noxref_21_M166_noxref_g ) capacitor \
 c=0.015318f //x=84.475 //y=5.02 //x2=84.84 //y2=6.02
cc_1974 ( N_VDD_c_1994_p N_noxref_21_M167_noxref_g ) capacitor c=0.00675379f \
 //x=85.415 //y=7.4 //x2=85.28 //y2=6.02
cc_1975 ( N_VDD_M167_noxref_d N_noxref_21_M167_noxref_g ) capacitor \
 c=0.0394719f //x=85.355 //y=5.02 //x2=85.28 //y2=6.02
cc_1976 ( N_VDD_c_1085_p N_noxref_21_M150_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=73.535 //y2=5.02
cc_1977 ( N_VDD_c_1249_p N_noxref_21_M150_noxref_d ) capacitor c=0.0139598f \
 //x=74.035 //y=7.4 //x2=73.535 //y2=5.02
cc_1978 ( N_VDD_M151_noxref_d N_noxref_21_M150_noxref_d ) capacitor \
 c=0.0664752f //x=73.975 //y=5.02 //x2=73.535 //y2=5.02
cc_1979 ( N_VDD_c_1085_p N_noxref_21_M152_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=74.415 //y2=5.02
cc_1980 ( N_VDD_c_1840_p N_noxref_21_M152_noxref_d ) capacitor c=0.0139598f \
 //x=74.915 //y=7.4 //x2=74.415 //y2=5.02
cc_1981 ( N_VDD_c_1080_n N_noxref_21_M152_noxref_d ) capacitor c=4.9285e-19 \
 //x=76.96 //y=7.4 //x2=74.415 //y2=5.02
cc_1982 ( N_VDD_M150_noxref_s N_noxref_21_M152_noxref_d ) capacitor \
 c=0.00130656f //x=73.105 //y=5.02 //x2=74.415 //y2=5.02
cc_1983 ( N_VDD_M151_noxref_d N_noxref_21_M152_noxref_d ) capacitor \
 c=0.0664752f //x=73.975 //y=5.02 //x2=74.415 //y2=5.02
cc_1984 ( N_VDD_M153_noxref_d N_noxref_21_M152_noxref_d ) capacitor \
 c=0.0664752f //x=74.855 //y=5.02 //x2=74.415 //y2=5.02
cc_1985 ( N_VDD_c_1085_p N_noxref_21_M154_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=75.295 //y2=5.02
cc_1986 ( N_VDD_c_1928_p N_noxref_21_M154_noxref_d ) capacitor c=0.014035f \
 //x=75.795 //y=7.4 //x2=75.295 //y2=5.02
cc_1987 ( N_VDD_c_1080_n N_noxref_21_M154_noxref_d ) capacitor c=0.00939849f \
 //x=76.96 //y=7.4 //x2=75.295 //y2=5.02
cc_1988 ( N_VDD_M153_noxref_d N_noxref_21_M154_noxref_d ) capacitor \
 c=0.0664752f //x=74.855 //y=5.02 //x2=75.295 //y2=5.02
cc_1989 ( N_VDD_M155_noxref_d N_noxref_21_M154_noxref_d ) capacitor \
 c=0.0664752f //x=75.735 //y=5.02 //x2=75.295 //y2=5.02
cc_1990 ( N_VDD_M156_noxref_s N_noxref_21_M154_noxref_d ) capacitor \
 c=3.57641e-19 //x=77.915 //y=5.02 //x2=75.295 //y2=5.02
cc_1991 ( N_VDD_c_1081_n N_noxref_22_c_9175_n ) capacitor c=5.72823e-19 \
 //x=81.77 //y=7.4 //x2=80.29 //y2=2.08
cc_1992 ( N_VDD_c_1085_p N_noxref_22_c_9180_n ) capacitor c=0.00444892f \
 //x=95.83 //y=7.4 //x2=84.095 //y2=5.155
cc_1993 ( N_VDD_c_1281_p N_noxref_22_c_9180_n ) capacitor c=4.31931e-19 \
 //x=83.655 //y=7.4 //x2=84.095 //y2=5.155
cc_1994 ( N_VDD_c_1964_p N_noxref_22_c_9180_n ) capacitor c=4.31931e-19 \
 //x=84.535 //y=7.4 //x2=84.095 //y2=5.155
cc_1995 ( N_VDD_M163_noxref_d N_noxref_22_c_9180_n ) capacitor c=0.0112985f \
 //x=83.595 //y=5.02 //x2=84.095 //y2=5.155
cc_1996 ( N_VDD_c_1081_n N_noxref_22_c_9184_n ) capacitor c=0.00863585f \
 //x=81.77 //y=7.4 //x2=83.385 //y2=5.155
cc_1997 ( N_VDD_M162_noxref_s N_noxref_22_c_9184_n ) capacitor c=0.0831083f \
 //x=82.725 //y=5.02 //x2=83.385 //y2=5.155
cc_1998 ( N_VDD_c_1085_p N_noxref_22_c_9186_n ) capacitor c=0.0044221f \
 //x=95.83 //y=7.4 //x2=84.975 //y2=5.155
cc_1999 ( N_VDD_c_1964_p N_noxref_22_c_9186_n ) capacitor c=4.31931e-19 \
 //x=84.535 //y=7.4 //x2=84.975 //y2=5.155
cc_2000 ( N_VDD_c_1994_p N_noxref_22_c_9186_n ) capacitor c=4.31931e-19 \
 //x=85.415 //y=7.4 //x2=84.975 //y2=5.155
cc_2001 ( N_VDD_M165_noxref_d N_noxref_22_c_9186_n ) capacitor c=0.0112985f \
 //x=84.475 //y=5.02 //x2=84.975 //y2=5.155
cc_2002 ( N_VDD_c_1085_p N_noxref_22_c_9190_n ) capacitor c=0.00434174f \
 //x=95.83 //y=7.4 //x2=85.755 //y2=5.155
cc_2003 ( N_VDD_c_1994_p N_noxref_22_c_9190_n ) capacitor c=7.46626e-19 \
 //x=85.415 //y=7.4 //x2=85.755 //y2=5.155
cc_2004 ( N_VDD_c_1282_p N_noxref_22_c_9190_n ) capacitor c=0.00198565f \
 //x=86.41 //y=7.4 //x2=85.755 //y2=5.155
cc_2005 ( N_VDD_M167_noxref_d N_noxref_22_c_9190_n ) capacitor c=0.0112985f \
 //x=85.355 //y=5.02 //x2=85.755 //y2=5.155
cc_2006 ( N_VDD_M168_noxref_s N_noxref_22_c_9190_n ) capacitor c=4.06494e-19 \
 //x=87.235 //y=5.025 //x2=85.755 //y2=5.155
cc_2007 ( N_VDD_c_1082_n N_noxref_22_c_9177_n ) capacitor c=0.0423183f \
 //x=86.58 //y=7.4 //x2=85.84 //y2=2.59
cc_2008 ( N_VDD_c_2030_p N_noxref_22_M160_noxref_g ) capacitor c=0.00675175f \
 //x=80.605 //y=7.4 //x2=80.03 //y2=6.02
cc_2009 ( N_VDD_M159_noxref_d N_noxref_22_M160_noxref_g ) capacitor \
 c=0.015318f //x=79.665 //y=5.02 //x2=80.03 //y2=6.02
cc_2010 ( N_VDD_c_2030_p N_noxref_22_M161_noxref_g ) capacitor c=0.00675379f \
 //x=80.605 //y=7.4 //x2=80.47 //y2=6.02
cc_2011 ( N_VDD_M161_noxref_d N_noxref_22_M161_noxref_g ) capacitor \
 c=0.0394719f //x=80.545 //y=5.02 //x2=80.47 //y2=6.02
cc_2012 ( N_VDD_c_1085_p N_noxref_22_M162_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=83.155 //y2=5.02
cc_2013 ( N_VDD_c_1281_p N_noxref_22_M162_noxref_d ) capacitor c=0.014035f \
 //x=83.655 //y=7.4 //x2=83.155 //y2=5.02
cc_2014 ( N_VDD_M163_noxref_d N_noxref_22_M162_noxref_d ) capacitor \
 c=0.0664752f //x=83.595 //y=5.02 //x2=83.155 //y2=5.02
cc_2015 ( N_VDD_c_1085_p N_noxref_22_M164_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=84.035 //y2=5.02
cc_2016 ( N_VDD_c_1964_p N_noxref_22_M164_noxref_d ) capacitor c=0.014035f \
 //x=84.535 //y=7.4 //x2=84.035 //y2=5.02
cc_2017 ( N_VDD_c_1082_n N_noxref_22_M164_noxref_d ) capacitor c=4.9285e-19 \
 //x=86.58 //y=7.4 //x2=84.035 //y2=5.02
cc_2018 ( N_VDD_M162_noxref_s N_noxref_22_M164_noxref_d ) capacitor \
 c=0.00130656f //x=82.725 //y=5.02 //x2=84.035 //y2=5.02
cc_2019 ( N_VDD_M163_noxref_d N_noxref_22_M164_noxref_d ) capacitor \
 c=0.0664752f //x=83.595 //y=5.02 //x2=84.035 //y2=5.02
cc_2020 ( N_VDD_M165_noxref_d N_noxref_22_M164_noxref_d ) capacitor \
 c=0.0664752f //x=84.475 //y=5.02 //x2=84.035 //y2=5.02
cc_2021 ( N_VDD_c_1085_p N_noxref_22_M166_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=84.915 //y2=5.02
cc_2022 ( N_VDD_c_1994_p N_noxref_22_M166_noxref_d ) capacitor c=0.014035f \
 //x=85.415 //y=7.4 //x2=84.915 //y2=5.02
cc_2023 ( N_VDD_c_1082_n N_noxref_22_M166_noxref_d ) capacitor c=0.00939849f \
 //x=86.58 //y=7.4 //x2=84.915 //y2=5.02
cc_2024 ( N_VDD_M165_noxref_d N_noxref_22_M166_noxref_d ) capacitor \
 c=0.0664752f //x=84.475 //y=5.02 //x2=84.915 //y2=5.02
cc_2025 ( N_VDD_M167_noxref_d N_noxref_22_M166_noxref_d ) capacitor \
 c=0.0664752f //x=85.355 //y=5.02 //x2=84.915 //y2=5.02
cc_2026 ( N_VDD_M168_noxref_s N_noxref_22_M166_noxref_d ) capacitor \
 c=4.52683e-19 //x=87.235 //y=5.025 //x2=84.915 //y2=5.02
cc_2027 ( N_VDD_c_1085_p N_noxref_23_c_9342_n ) capacitor c=0.0206457f \
 //x=95.83 //y=7.4 //x2=90.575 //y2=5.21
cc_2028 ( N_VDD_c_2050_p N_noxref_23_c_9342_n ) capacitor c=0.00213763f \
 //x=89.045 //y=7.4 //x2=90.575 //y2=5.21
cc_2029 ( N_VDD_c_2051_p N_noxref_23_c_9342_n ) capacitor c=0.003172f \
 //x=89.74 //y=7.4 //x2=90.575 //y2=5.21
cc_2030 ( N_VDD_c_1331_p N_noxref_23_c_9342_n ) capacitor c=0.00424633f \
 //x=93.07 //y=7.4 //x2=90.575 //y2=5.21
cc_2031 ( N_VDD_c_1083_n N_noxref_23_c_9342_n ) capacitor c=0.0430305f \
 //x=89.91 //y=7.4 //x2=90.575 //y2=5.21
cc_2032 ( N_VDD_M171_noxref_d N_noxref_23_c_9342_n ) capacitor c=0.0197937f \
 //x=88.985 //y=5.025 //x2=90.575 //y2=5.21
cc_2033 ( N_VDD_c_1085_p N_noxref_23_c_9348_n ) capacitor c=0.00274812f \
 //x=95.83 //y=7.4 //x2=88.805 //y2=5.21
cc_2034 ( N_VDD_c_2050_p N_noxref_23_c_9348_n ) capacitor c=0.00107267f \
 //x=89.045 //y=7.4 //x2=88.805 //y2=5.21
cc_2035 ( N_VDD_c_1082_n N_noxref_23_c_9348_n ) capacitor c=2.89592e-19 \
 //x=86.58 //y=7.4 //x2=88.805 //y2=5.21
cc_2036 ( N_VDD_c_1083_n N_noxref_23_c_9348_n ) capacitor c=3.35418e-19 \
 //x=89.91 //y=7.4 //x2=88.805 //y2=5.21
cc_2037 ( N_VDD_M171_noxref_d N_noxref_23_c_9348_n ) capacitor c=6.02701e-19 \
 //x=88.985 //y=5.025 //x2=88.805 //y2=5.21
cc_2038 ( N_VDD_c_1085_p N_noxref_23_c_9353_n ) capacitor c=0.00453889f \
 //x=95.83 //y=7.4 //x2=88.605 //y2=5.21
cc_2039 ( N_VDD_c_1290_p N_noxref_23_c_9353_n ) capacitor c=4.52207e-19 \
 //x=88.165 //y=7.4 //x2=88.605 //y2=5.21
cc_2040 ( N_VDD_c_2050_p N_noxref_23_c_9353_n ) capacitor c=4.11408e-19 \
 //x=89.045 //y=7.4 //x2=88.605 //y2=5.21
cc_2041 ( N_VDD_M169_noxref_d N_noxref_23_c_9353_n ) capacitor c=0.0127968f \
 //x=88.105 //y=5.025 //x2=88.605 //y2=5.21
cc_2042 ( N_VDD_c_1082_n N_noxref_23_c_9357_n ) capacitor c=0.00914165f \
 //x=86.58 //y=7.4 //x2=87.895 //y2=5.21
cc_2043 ( N_VDD_M168_noxref_s N_noxref_23_c_9357_n ) capacitor c=0.0872987f \
 //x=87.235 //y=5.025 //x2=87.895 //y2=5.21
cc_2044 ( N_VDD_c_1082_n N_noxref_23_c_9359_n ) capacitor c=6.3991e-19 \
 //x=86.58 //y=7.4 //x2=88.69 //y2=5.295
cc_2045 ( N_VDD_c_1083_n N_noxref_23_c_9359_n ) capacitor c=0.00985441f \
 //x=89.91 //y=7.4 //x2=88.69 //y2=5.295
cc_2046 ( N_VDD_M171_noxref_d N_noxref_23_c_9359_n ) capacitor c=0.0873334f \
 //x=88.985 //y=5.025 //x2=88.69 //y2=5.295
cc_2047 ( N_VDD_c_1083_n N_noxref_23_c_9362_n ) capacitor c=0.0674112f \
 //x=89.91 //y=7.4 //x2=90.69 //y2=5.21
cc_2048 ( N_VDD_M171_noxref_d N_noxref_23_c_9362_n ) capacitor c=0.00235009f \
 //x=88.985 //y=5.025 //x2=90.69 //y2=5.21
cc_2049 ( N_VDD_c_1085_p N_noxref_23_c_9364_n ) capacitor c=0.0296361f \
 //x=95.83 //y=7.4 //x2=90.775 //y2=6.91
cc_2050 ( N_VDD_c_1331_p N_noxref_23_c_9364_n ) capacitor c=0.109938f \
 //x=93.07 //y=7.4 //x2=90.775 //y2=6.91
cc_2051 ( N_VDD_c_1085_p N_noxref_23_M168_noxref_d ) capacitor c=0.00291898f \
 //x=95.83 //y=7.4 //x2=87.665 //y2=5.025
cc_2052 ( N_VDD_c_1290_p N_noxref_23_M168_noxref_d ) capacitor c=0.0137097f \
 //x=88.165 //y=7.4 //x2=87.665 //y2=5.025
cc_2053 ( N_VDD_M169_noxref_d N_noxref_23_M168_noxref_d ) capacitor \
 c=0.067695f //x=88.105 //y=5.025 //x2=87.665 //y2=5.025
cc_2054 ( N_VDD_M171_noxref_d N_noxref_23_M168_noxref_d ) capacitor \
 c=0.00105738f //x=88.985 //y=5.025 //x2=87.665 //y2=5.025
cc_2055 ( N_VDD_c_1085_p N_noxref_23_M170_noxref_d ) capacitor c=0.00241371f \
 //x=95.83 //y=7.4 //x2=88.545 //y2=5.025
cc_2056 ( N_VDD_c_2050_p N_noxref_23_M170_noxref_d ) capacitor c=0.01268f \
 //x=89.045 //y=7.4 //x2=88.545 //y2=5.025
cc_2057 ( N_VDD_M168_noxref_s N_noxref_23_M170_noxref_d ) capacitor \
 c=0.00103189f //x=87.235 //y=5.025 //x2=88.545 //y2=5.025
cc_2058 ( N_VDD_M169_noxref_d N_noxref_23_M170_noxref_d ) capacitor \
 c=0.0653408f //x=88.105 //y=5.025 //x2=88.545 //y2=5.025
cc_2059 ( N_VDD_c_1083_n N_noxref_23_M173_noxref_d ) capacitor c=8.96067e-19 \
 //x=89.91 //y=7.4 //x2=91.425 //y2=5.025
cc_2060 ( N_VDD_c_1084_n N_noxref_23_M173_noxref_d ) capacitor c=8.88629e-19 \
 //x=93.24 //y=7.4 //x2=91.425 //y2=5.025
cc_2061 ( N_VDD_c_1084_n N_noxref_23_M175_noxref_d ) capacitor c=0.0575594f \
 //x=93.24 //y=7.4 //x2=92.305 //y2=5.025
cc_2062 ( N_VDD_c_1085_p N_noxref_24_c_9478_n ) capacitor c=0.00444892f \
 //x=95.83 //y=7.4 //x2=79.285 //y2=5.155
cc_2063 ( N_VDD_c_1278_p N_noxref_24_c_9478_n ) capacitor c=4.31931e-19 \
 //x=78.845 //y=7.4 //x2=79.285 //y2=5.155
cc_2064 ( N_VDD_c_1932_p N_noxref_24_c_9478_n ) capacitor c=4.31931e-19 \
 //x=79.725 //y=7.4 //x2=79.285 //y2=5.155
cc_2065 ( N_VDD_M157_noxref_d N_noxref_24_c_9478_n ) capacitor c=0.0112985f \
 //x=78.785 //y=5.02 //x2=79.285 //y2=5.155
cc_2066 ( N_VDD_c_1080_n N_noxref_24_c_9482_n ) capacitor c=0.00863585f \
 //x=76.96 //y=7.4 //x2=78.575 //y2=5.155
cc_2067 ( N_VDD_M156_noxref_s N_noxref_24_c_9482_n ) capacitor c=0.0831083f \
 //x=77.915 //y=5.02 //x2=78.575 //y2=5.155
cc_2068 ( N_VDD_c_1085_p N_noxref_24_c_9484_n ) capacitor c=0.0044221f \
 //x=95.83 //y=7.4 //x2=80.165 //y2=5.155
cc_2069 ( N_VDD_c_1932_p N_noxref_24_c_9484_n ) capacitor c=4.31931e-19 \
 //x=79.725 //y=7.4 //x2=80.165 //y2=5.155
cc_2070 ( N_VDD_c_2030_p N_noxref_24_c_9484_n ) capacitor c=4.31931e-19 \
 //x=80.605 //y=7.4 //x2=80.165 //y2=5.155
cc_2071 ( N_VDD_M159_noxref_d N_noxref_24_c_9484_n ) capacitor c=0.0112985f \
 //x=79.665 //y=5.02 //x2=80.165 //y2=5.155
cc_2072 ( N_VDD_c_1085_p N_noxref_24_c_9488_n ) capacitor c=0.00434174f \
 //x=95.83 //y=7.4 //x2=80.945 //y2=5.155
cc_2073 ( N_VDD_c_2030_p N_noxref_24_c_9488_n ) capacitor c=7.46626e-19 \
 //x=80.605 //y=7.4 //x2=80.945 //y2=5.155
cc_2074 ( N_VDD_c_1279_p N_noxref_24_c_9488_n ) capacitor c=0.00198565f \
 //x=81.6 //y=7.4 //x2=80.945 //y2=5.155
cc_2075 ( N_VDD_M161_noxref_d N_noxref_24_c_9488_n ) capacitor c=0.0112985f \
 //x=80.545 //y=5.02 //x2=80.945 //y2=5.155
cc_2076 ( N_VDD_c_1081_n N_noxref_24_c_9451_n ) capacitor c=0.0428142f \
 //x=81.77 //y=7.4 //x2=81.03 //y2=2.22
cc_2077 ( N_VDD_c_1085_p N_noxref_24_c_9452_n ) capacitor c=9.10347e-19 \
 //x=95.83 //y=7.4 //x2=82.88 //y2=2.08
cc_2078 ( N_VDD_c_1081_n N_noxref_24_c_9452_n ) capacitor c=0.0134711f \
 //x=81.77 //y=7.4 //x2=82.88 //y2=2.08
cc_2079 ( N_VDD_M162_noxref_s N_noxref_24_c_9452_n ) capacitor c=0.0125322f \
 //x=82.725 //y=5.02 //x2=82.88 //y2=2.08
cc_2080 ( N_VDD_c_1083_n N_noxref_24_c_9453_n ) capacitor c=7.57423e-19 \
 //x=89.91 //y=7.4 //x2=92.5 //y2=2.08
cc_2081 ( N_VDD_c_1084_n N_noxref_24_c_9453_n ) capacitor c=0.0263215f \
 //x=93.24 //y=7.4 //x2=92.5 //y2=2.08
cc_2082 ( N_VDD_c_1084_n N_noxref_24_c_9455_n ) capacitor c=0.0263871f \
 //x=93.24 //y=7.4 //x2=93.98 //y2=2.08
cc_2083 ( N_VDD_c_1281_p N_noxref_24_M162_noxref_g ) capacitor c=0.00749687f \
 //x=83.655 //y=7.4 //x2=83.08 //y2=6.02
cc_2084 ( N_VDD_M162_noxref_s N_noxref_24_M162_noxref_g ) capacitor \
 c=0.0477201f //x=82.725 //y=5.02 //x2=83.08 //y2=6.02
cc_2085 ( N_VDD_c_1281_p N_noxref_24_M163_noxref_g ) capacitor c=0.00675175f \
 //x=83.655 //y=7.4 //x2=83.52 //y2=6.02
cc_2086 ( N_VDD_M163_noxref_d N_noxref_24_M163_noxref_g ) capacitor \
 c=0.015318f //x=83.595 //y=5.02 //x2=83.52 //y2=6.02
cc_2087 ( N_VDD_c_1331_p N_noxref_24_M174_noxref_g ) capacitor c=0.00512552f \
 //x=93.07 //y=7.4 //x2=91.79 //y2=6.025
cc_2088 ( N_VDD_c_1331_p N_noxref_24_M175_noxref_g ) capacitor c=0.00512552f \
 //x=93.07 //y=7.4 //x2=92.23 //y2=6.025
cc_2089 ( N_VDD_c_1084_n N_noxref_24_M175_noxref_g ) capacitor c=0.010355f \
 //x=93.24 //y=7.4 //x2=92.23 //y2=6.025
cc_2090 ( N_VDD_c_1064_n N_noxref_24_M176_noxref_g ) capacitor c=0.00512552f \
 //x=95.83 //y=7.4 //x2=94.25 //y2=6.025
cc_2091 ( N_VDD_c_1084_n N_noxref_24_M176_noxref_g ) capacitor c=0.00767856f \
 //x=93.24 //y=7.4 //x2=94.25 //y2=6.025
cc_2092 ( N_VDD_c_1064_n N_noxref_24_M177_noxref_g ) capacitor c=0.00512552f \
 //x=95.83 //y=7.4 //x2=94.69 //y2=6.025
cc_2093 ( N_VDD_c_1081_n N_noxref_24_c_9509_n ) capacitor c=0.0076931f \
 //x=81.77 //y=7.4 //x2=83.155 //y2=4.79
cc_2094 ( N_VDD_M162_noxref_s N_noxref_24_c_9509_n ) capacitor c=0.00444914f \
 //x=82.725 //y=5.02 //x2=83.155 //y2=4.79
cc_2095 ( N_VDD_c_1084_n N_noxref_24_c_9511_n ) capacitor c=0.00803198f \
 //x=93.24 //y=7.4 //x2=92.23 //y2=4.87
cc_2096 ( N_VDD_c_1084_n N_noxref_24_c_9512_n ) capacitor c=0.00803198f \
 //x=93.24 //y=7.4 //x2=94.325 //y2=4.795
cc_2097 ( N_VDD_c_1085_p N_noxref_24_M156_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=78.345 //y2=5.02
cc_2098 ( N_VDD_c_1278_p N_noxref_24_M156_noxref_d ) capacitor c=0.014035f \
 //x=78.845 //y=7.4 //x2=78.345 //y2=5.02
cc_2099 ( N_VDD_M157_noxref_d N_noxref_24_M156_noxref_d ) capacitor \
 c=0.0664752f //x=78.785 //y=5.02 //x2=78.345 //y2=5.02
cc_2100 ( N_VDD_c_1085_p N_noxref_24_M158_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=79.225 //y2=5.02
cc_2101 ( N_VDD_c_1932_p N_noxref_24_M158_noxref_d ) capacitor c=0.014035f \
 //x=79.725 //y=7.4 //x2=79.225 //y2=5.02
cc_2102 ( N_VDD_c_1081_n N_noxref_24_M158_noxref_d ) capacitor c=4.9285e-19 \
 //x=81.77 //y=7.4 //x2=79.225 //y2=5.02
cc_2103 ( N_VDD_M156_noxref_s N_noxref_24_M158_noxref_d ) capacitor \
 c=0.00130656f //x=77.915 //y=5.02 //x2=79.225 //y2=5.02
cc_2104 ( N_VDD_M157_noxref_d N_noxref_24_M158_noxref_d ) capacitor \
 c=0.0664752f //x=78.785 //y=5.02 //x2=79.225 //y2=5.02
cc_2105 ( N_VDD_M159_noxref_d N_noxref_24_M158_noxref_d ) capacitor \
 c=0.0664752f //x=79.665 //y=5.02 //x2=79.225 //y2=5.02
cc_2106 ( N_VDD_c_1085_p N_noxref_24_M160_noxref_d ) capacitor c=0.00275235f \
 //x=95.83 //y=7.4 //x2=80.105 //y2=5.02
cc_2107 ( N_VDD_c_2030_p N_noxref_24_M160_noxref_d ) capacitor c=0.014035f \
 //x=80.605 //y=7.4 //x2=80.105 //y2=5.02
cc_2108 ( N_VDD_c_1081_n N_noxref_24_M160_noxref_d ) capacitor c=0.00939849f \
 //x=81.77 //y=7.4 //x2=80.105 //y2=5.02
cc_2109 ( N_VDD_M159_noxref_d N_noxref_24_M160_noxref_d ) capacitor \
 c=0.0664752f //x=79.665 //y=5.02 //x2=80.105 //y2=5.02
cc_2110 ( N_VDD_M161_noxref_d N_noxref_24_M160_noxref_d ) capacitor \
 c=0.0664752f //x=80.545 //y=5.02 //x2=80.105 //y2=5.02
cc_2111 ( N_VDD_M162_noxref_s N_noxref_24_M160_noxref_d ) capacitor \
 c=3.57641e-19 //x=82.725 //y=5.02 //x2=80.105 //y2=5.02
cc_2112 ( N_VDD_c_1085_p N_noxref_25_c_9823_n ) capacitor c=0.0212729f \
 //x=95.83 //y=7.4 //x2=93.915 //y2=5.21
cc_2113 ( N_VDD_c_1331_p N_noxref_25_c_9823_n ) capacitor c=0.00386143f \
 //x=93.07 //y=7.4 //x2=93.915 //y2=5.21
cc_2114 ( N_VDD_c_1064_n N_noxref_25_c_9823_n ) capacitor c=0.00403412f \
 //x=95.83 //y=7.4 //x2=93.915 //y2=5.21
cc_2115 ( N_VDD_c_1084_n N_noxref_25_c_9823_n ) capacitor c=0.0473381f \
 //x=93.24 //y=7.4 //x2=93.915 //y2=5.21
cc_2116 ( N_VDD_c_1085_p N_noxref_25_c_9827_n ) capacitor c=0.00264311f \
 //x=95.83 //y=7.4 //x2=92.125 //y2=5.21
cc_2117 ( N_VDD_c_1084_n N_noxref_25_c_9827_n ) capacitor c=6.67754e-19 \
 //x=93.24 //y=7.4 //x2=92.125 //y2=5.21
cc_2118 ( N_VDD_c_1083_n N_noxref_25_c_9829_n ) capacitor c=0.00662411f \
 //x=89.91 //y=7.4 //x2=91.215 //y2=5.21
cc_2119 ( N_VDD_c_1084_n N_noxref_25_c_9830_n ) capacitor c=0.00999961f \
 //x=93.24 //y=7.4 //x2=92.01 //y2=5.295
cc_2120 ( N_VDD_c_1064_n N_noxref_25_c_9831_n ) capacitor c=6.48751e-19 \
 //x=95.83 //y=7.4 //x2=94.03 //y2=5.21
cc_2121 ( N_VDD_c_1084_n N_noxref_25_c_9831_n ) capacitor c=0.0664301f \
 //x=93.24 //y=7.4 //x2=94.03 //y2=5.21
cc_2122 ( N_VDD_c_1085_p N_noxref_25_c_9833_n ) capacitor c=0.0387208f \
 //x=95.83 //y=7.4 //x2=94.115 //y2=6.91
cc_2123 ( N_VDD_c_1064_n N_noxref_25_c_9833_n ) capacitor c=0.108798f \
 //x=95.83 //y=7.4 //x2=94.115 //y2=6.91
cc_2124 ( N_VDD_c_1064_n N_noxref_25_M177_noxref_d ) capacitor c=8.96067e-19 \
 //x=95.83 //y=7.4 //x2=94.765 //y2=5.025
cc_2125 ( N_VDD_c_1084_n N_noxref_25_M177_noxref_d ) capacitor c=8.88629e-19 \
 //x=93.24 //y=7.4 //x2=94.765 //y2=5.025
cc_2126 ( N_VDD_c_1064_n N_noxref_25_M179_noxref_d ) capacitor c=0.0529764f \
 //x=95.83 //y=7.4 //x2=95.645 //y2=5.025
cc_2127 ( N_VDD_c_1077_n N_noxref_26_c_9933_n ) capacitor c=0.00686843f \
 //x=62.53 //y=7.4 //x2=65.035 //y2=3.7
cc_2128 ( N_VDD_c_1078_n N_noxref_26_c_9912_n ) capacitor c=0.0140578f \
 //x=67.34 //y=7.4 //x2=88.315 //y2=4.07
cc_2129 ( N_VDD_c_1079_n N_noxref_26_c_9912_n ) capacitor c=0.0140578f \
 //x=72.15 //y=7.4 //x2=88.315 //y2=4.07
cc_2130 ( N_VDD_c_1080_n N_noxref_26_c_9912_n ) capacitor c=0.0140578f \
 //x=76.96 //y=7.4 //x2=88.315 //y2=4.07
cc_2131 ( N_VDD_c_1081_n N_noxref_26_c_9912_n ) capacitor c=0.0140578f \
 //x=81.77 //y=7.4 //x2=88.315 //y2=4.07
cc_2132 ( N_VDD_c_1082_n N_noxref_26_c_9912_n ) capacitor c=0.0145414f \
 //x=86.58 //y=7.4 //x2=88.315 //y2=4.07
cc_2133 ( N_VDD_c_1085_p N_noxref_26_c_9913_n ) capacitor c=0.0151699f \
 //x=95.83 //y=7.4 //x2=94.975 //y2=4.07
cc_2134 ( N_VDD_c_1064_n N_noxref_26_c_9913_n ) capacitor c=4.075e-19 \
 //x=95.83 //y=7.4 //x2=94.975 //y2=4.07
cc_2135 ( N_VDD_c_1083_n N_noxref_26_c_9913_n ) capacitor c=0.0153579f \
 //x=89.91 //y=7.4 //x2=94.975 //y2=4.07
cc_2136 ( N_VDD_c_1084_n N_noxref_26_c_9913_n ) capacitor c=0.0225025f \
 //x=93.24 //y=7.4 //x2=94.975 //y2=4.07
cc_2137 ( N_VDD_c_1083_n N_noxref_26_c_9943_n ) capacitor c=5.4458e-19 \
 //x=89.91 //y=7.4 //x2=88.545 //y2=4.07
cc_2138 ( N_VDD_c_1085_p N_noxref_26_c_9944_n ) capacitor c=0.00437246f \
 //x=95.83 //y=7.4 //x2=50.425 //y2=5.155
cc_2139 ( N_VDD_c_1234_p N_noxref_26_c_9944_n ) capacitor c=4.31596e-19 \
 //x=49.985 //y=7.4 //x2=50.425 //y2=5.155
cc_2140 ( N_VDD_c_1920_p N_noxref_26_c_9944_n ) capacitor c=4.31596e-19 \
 //x=50.865 //y=7.4 //x2=50.425 //y2=5.155
cc_2141 ( N_VDD_M121_noxref_d N_noxref_26_c_9944_n ) capacitor c=0.0109802f \
 //x=49.925 //y=5.02 //x2=50.425 //y2=5.155
cc_2142 ( N_VDD_c_1074_n N_noxref_26_c_9948_n ) capacitor c=0.00863585f \
 //x=48.1 //y=7.4 //x2=49.715 //y2=5.155
cc_2143 ( N_VDD_M120_noxref_s N_noxref_26_c_9948_n ) capacitor c=0.0831083f \
 //x=49.055 //y=5.02 //x2=49.715 //y2=5.155
cc_2144 ( N_VDD_c_1085_p N_noxref_26_c_9950_n ) capacitor c=0.00434259f \
 //x=95.83 //y=7.4 //x2=51.305 //y2=5.155
cc_2145 ( N_VDD_c_1920_p N_noxref_26_c_9950_n ) capacitor c=4.31596e-19 \
 //x=50.865 //y=7.4 //x2=51.305 //y2=5.155
cc_2146 ( N_VDD_c_1626_p N_noxref_26_c_9950_n ) capacitor c=4.31596e-19 \
 //x=51.745 //y=7.4 //x2=51.305 //y2=5.155
cc_2147 ( N_VDD_M123_noxref_d N_noxref_26_c_9950_n ) capacitor c=0.0109802f \
 //x=50.805 //y=5.02 //x2=51.305 //y2=5.155
cc_2148 ( N_VDD_c_1085_p N_noxref_26_c_9954_n ) capacitor c=0.00424413f \
 //x=95.83 //y=7.4 //x2=52.085 //y2=5.155
cc_2149 ( N_VDD_c_1626_p N_noxref_26_c_9954_n ) capacitor c=7.45454e-19 \
 //x=51.745 //y=7.4 //x2=52.085 //y2=5.155
cc_2150 ( N_VDD_c_1235_p N_noxref_26_c_9954_n ) capacitor c=0.00198097f \
 //x=52.74 //y=7.4 //x2=52.085 //y2=5.155
cc_2151 ( N_VDD_M125_noxref_d N_noxref_26_c_9954_n ) capacitor c=0.0109802f \
 //x=51.685 //y=5.02 //x2=52.085 //y2=5.155
cc_2152 ( N_VDD_c_1075_n N_noxref_26_c_9958_n ) capacitor c=0.0401694f \
 //x=52.91 //y=7.4 //x2=52.17 //y2=3.33
cc_2153 ( N_VDD_c_1085_p N_noxref_26_c_9916_n ) capacitor c=6.51035e-19 \
 //x=95.83 //y=7.4 //x2=54.02 //y2=2.08
cc_2154 ( N_VDD_c_1075_n N_noxref_26_c_9916_n ) capacitor c=0.0115064f \
 //x=52.91 //y=7.4 //x2=54.02 //y2=2.08
cc_2155 ( N_VDD_M126_noxref_s N_noxref_26_c_9916_n ) capacitor c=0.00923513f \
 //x=53.865 //y=5.02 //x2=54.02 //y2=2.08
cc_2156 ( N_VDD_c_1083_n N_noxref_26_c_9962_n ) capacitor c=0.00491684f \
 //x=89.91 //y=7.4 //x2=88.43 //y2=4.54
cc_2157 ( N_VDD_c_1082_n N_noxref_26_c_9917_n ) capacitor c=7.12079e-19 \
 //x=86.58 //y=7.4 //x2=88.43 //y2=2.08
cc_2158 ( N_VDD_c_1083_n N_noxref_26_c_9917_n ) capacitor c=0.0042566f \
 //x=89.91 //y=7.4 //x2=88.43 //y2=2.08
cc_2159 ( N_VDD_c_1064_n N_noxref_26_c_9919_n ) capacitor c=6.51778e-19 \
 //x=95.83 //y=7.4 //x2=95.09 //y2=2.08
cc_2160 ( N_VDD_c_1084_n N_noxref_26_c_9919_n ) capacitor c=0.00116377f \
 //x=93.24 //y=7.4 //x2=95.09 //y2=2.08
cc_2161 ( N_VDD_c_1237_p N_noxref_26_M126_noxref_g ) capacitor c=0.00749687f \
 //x=54.795 //y=7.4 //x2=54.22 //y2=6.02
cc_2162 ( N_VDD_M126_noxref_s N_noxref_26_M126_noxref_g ) capacitor \
 c=0.0477201f //x=53.865 //y=5.02 //x2=54.22 //y2=6.02
cc_2163 ( N_VDD_c_1237_p N_noxref_26_M127_noxref_g ) capacitor c=0.00675175f \
 //x=54.795 //y=7.4 //x2=54.66 //y2=6.02
cc_2164 ( N_VDD_M127_noxref_d N_noxref_26_M127_noxref_g ) capacitor \
 c=0.015318f //x=54.735 //y=5.02 //x2=54.66 //y2=6.02
cc_2165 ( N_VDD_c_2050_p N_noxref_26_M170_noxref_g ) capacitor c=0.0067918f \
 //x=89.045 //y=7.4 //x2=88.47 //y2=6.025
cc_2166 ( N_VDD_M169_noxref_d N_noxref_26_M170_noxref_g ) capacitor \
 c=0.015526f //x=88.105 //y=5.025 //x2=88.47 //y2=6.025
cc_2167 ( N_VDD_c_2050_p N_noxref_26_M171_noxref_g ) capacitor c=0.00754867f \
 //x=89.045 //y=7.4 //x2=88.91 //y2=6.025
cc_2168 ( N_VDD_M171_noxref_d N_noxref_26_M171_noxref_g ) capacitor \
 c=0.0537676f //x=88.985 //y=5.025 //x2=88.91 //y2=6.025
cc_2169 ( N_VDD_c_1064_n N_noxref_26_M178_noxref_g ) capacitor c=0.00513565f \
 //x=95.83 //y=7.4 //x2=95.13 //y2=6.025
cc_2170 ( N_VDD_c_1064_n N_noxref_26_M179_noxref_g ) capacitor c=0.0309137f \
 //x=95.83 //y=7.4 //x2=95.57 //y2=6.025
cc_2171 ( N_VDD_c_1075_n N_noxref_26_c_9977_n ) capacitor c=0.00540116f \
 //x=52.91 //y=7.4 //x2=54.295 //y2=4.79
cc_2172 ( N_VDD_M126_noxref_s N_noxref_26_c_9977_n ) capacitor c=0.00433385f \
 //x=53.865 //y=5.02 //x2=54.295 //y2=4.79
cc_2173 ( N_VDD_c_1083_n N_noxref_26_c_9979_n ) capacitor c=0.00985898f \
 //x=89.91 //y=7.4 //x2=88.835 //y2=4.795
cc_2174 ( N_VDD_c_1083_n N_noxref_26_c_9980_n ) capacitor c=2.76772e-19 \
 //x=89.91 //y=7.4 //x2=88.47 //y2=4.705
cc_2175 ( N_VDD_c_1085_p N_noxref_26_M120_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=49.485 //y2=5.02
cc_2176 ( N_VDD_c_1234_p N_noxref_26_M120_noxref_d ) capacitor c=0.0139598f \
 //x=49.985 //y=7.4 //x2=49.485 //y2=5.02
cc_2177 ( N_VDD_M121_noxref_d N_noxref_26_M120_noxref_d ) capacitor \
 c=0.0664752f //x=49.925 //y=5.02 //x2=49.485 //y2=5.02
cc_2178 ( N_VDD_c_1085_p N_noxref_26_M122_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=50.365 //y2=5.02
cc_2179 ( N_VDD_c_1920_p N_noxref_26_M122_noxref_d ) capacitor c=0.0139598f \
 //x=50.865 //y=7.4 //x2=50.365 //y2=5.02
cc_2180 ( N_VDD_c_1075_n N_noxref_26_M122_noxref_d ) capacitor c=4.9285e-19 \
 //x=52.91 //y=7.4 //x2=50.365 //y2=5.02
cc_2181 ( N_VDD_M120_noxref_s N_noxref_26_M122_noxref_d ) capacitor \
 c=0.00130656f //x=49.055 //y=5.02 //x2=50.365 //y2=5.02
cc_2182 ( N_VDD_M121_noxref_d N_noxref_26_M122_noxref_d ) capacitor \
 c=0.0664752f //x=49.925 //y=5.02 //x2=50.365 //y2=5.02
cc_2183 ( N_VDD_M123_noxref_d N_noxref_26_M122_noxref_d ) capacitor \
 c=0.0664752f //x=50.805 //y=5.02 //x2=50.365 //y2=5.02
cc_2184 ( N_VDD_c_1085_p N_noxref_26_M124_noxref_d ) capacitor c=0.00264488f \
 //x=95.83 //y=7.4 //x2=51.245 //y2=5.02
cc_2185 ( N_VDD_c_1626_p N_noxref_26_M124_noxref_d ) capacitor c=0.0139598f \
 //x=51.745 //y=7.4 //x2=51.245 //y2=5.02
cc_2186 ( N_VDD_c_1075_n N_noxref_26_M124_noxref_d ) capacitor c=0.00939849f \
 //x=52.91 //y=7.4 //x2=51.245 //y2=5.02
cc_2187 ( N_VDD_M123_noxref_d N_noxref_26_M124_noxref_d ) capacitor \
 c=0.0664752f //x=50.805 //y=5.02 //x2=51.245 //y2=5.02
cc_2188 ( N_VDD_M125_noxref_d N_noxref_26_M124_noxref_d ) capacitor \
 c=0.0664752f //x=51.685 //y=5.02 //x2=51.245 //y2=5.02
cc_2189 ( N_VDD_M126_noxref_s N_noxref_26_M124_noxref_d ) capacitor \
 c=3.57641e-19 //x=53.865 //y=5.02 //x2=51.245 //y2=5.02
cc_2190 ( N_VDD_c_1085_p Q ) capacitor c=0.00298795f //x=95.83 //y=7.4 \
 //x2=95.83 //y2=4.07
cc_2191 ( N_VDD_c_1064_n Q ) capacitor c=0.00255307f //x=95.83 //y=7.4 \
 //x2=95.83 //y2=4.07
cc_2192 ( N_VDD_c_1084_n N_Q_c_10397_n ) capacitor c=0.00660621f //x=93.24 \
 //y=7.4 //x2=94.555 //y2=5.21
cc_2193 ( N_VDD_c_1085_p N_Q_c_10398_n ) capacitor c=0.0017748f //x=95.83 \
 //y=7.4 //x2=95.745 //y2=5.21
cc_2194 ( N_VDD_c_1064_n N_Q_c_10398_n ) capacitor c=0.00139502f //x=95.83 \
 //y=7.4 //x2=95.745 //y2=5.21
cc_2195 ( N_VDD_c_1064_n N_Q_c_10384_n ) capacitor c=0.0468676f //x=95.83 \
 //y=7.4 //x2=95.83 //y2=4.07
cc_2196 ( N_VDD_c_1084_n N_Q_c_10384_n ) capacitor c=0.00147633f //x=93.24 \
 //y=7.4 //x2=95.83 //y2=4.07
cc_2197 ( N_VDD_c_1064_n N_Q_M176_noxref_d ) capacitor c=6.67979e-19 //x=95.83 \
 //y=7.4 //x2=94.325 //y2=5.025
cc_2198 ( N_VDD_c_1064_n N_Q_M178_noxref_d ) capacitor c=0.0099096f //x=95.83 \
 //y=7.4 //x2=95.205 //y2=5.025
cc_2199 ( N_noxref_3_c_2223_n N_noxref_4_c_2462_n ) capacitor c=0.00564994f \
 //x=10.615 //y=2.59 //x2=13.805 //y2=2.59
cc_2200 ( N_noxref_3_M73_noxref_g N_noxref_4_c_2477_n ) capacitor c=0.0168349f \
 //x=11.37 //y=6.02 //x2=11.945 //y2=5.155
cc_2201 ( N_noxref_3_M72_noxref_g N_noxref_4_c_2481_n ) capacitor c=0.0213876f \
 //x=10.93 //y=6.02 //x2=11.235 //y2=5.155
cc_2202 ( N_noxref_3_c_2301_p N_noxref_4_c_2481_n ) capacitor c=0.00428486f \
 //x=11.295 //y=4.79 //x2=11.235 //y2=5.155
cc_2203 ( N_noxref_3_M73_noxref_g N_noxref_4_M72_noxref_d ) capacitor \
 c=0.0180032f //x=11.37 //y=6.02 //x2=11.005 //y2=5.02
cc_2204 ( N_noxref_3_c_2221_n N_noxref_5_c_2626_n ) capacitor c=0.0709582f \
 //x=5.805 //y=2.59 //x2=8.765 //y2=3.33
cc_2205 ( N_noxref_3_c_2222_n N_noxref_5_c_2626_n ) capacitor c=0.0134806f \
 //x=4.185 //y=2.59 //x2=8.765 //y2=3.33
cc_2206 ( N_noxref_3_c_2223_n N_noxref_5_c_2626_n ) capacitor c=0.114019f \
 //x=10.615 //y=2.59 //x2=8.765 //y2=3.33
cc_2207 ( N_noxref_3_c_2224_n N_noxref_5_c_2626_n ) capacitor c=0.0123232f \
 //x=6.035 //y=2.59 //x2=8.765 //y2=3.33
cc_2208 ( N_noxref_3_c_2226_n N_noxref_5_c_2626_n ) capacitor c=0.0237657f \
 //x=4.07 //y=2.59 //x2=8.765 //y2=3.33
cc_2209 ( N_noxref_3_c_2227_n N_noxref_5_c_2626_n ) capacitor c=0.0247707f \
 //x=5.92 //y=2.08 //x2=8.765 //y2=3.33
cc_2210 ( N_noxref_3_c_2226_n N_noxref_5_c_2692_n ) capacitor c=0.00179385f \
 //x=4.07 //y=2.59 //x2=3.445 //y2=3.33
cc_2211 ( N_noxref_3_c_2223_n N_noxref_5_c_2627_n ) capacitor c=0.0846302f \
 //x=10.615 //y=2.59 //x2=20.235 //y2=3.33
cc_2212 ( N_noxref_3_c_2228_n N_noxref_5_c_2627_n ) capacitor c=0.0224325f \
 //x=10.73 //y=2.08 //x2=20.235 //y2=3.33
cc_2213 ( N_noxref_3_c_2223_n N_noxref_5_c_2695_n ) capacitor c=0.0120889f \
 //x=10.615 //y=2.59 //x2=8.995 //y2=3.33
cc_2214 ( N_noxref_3_c_2228_n N_noxref_5_c_2695_n ) capacitor c=7.01366e-19 \
 //x=10.73 //y=2.08 //x2=8.995 //y2=3.33
cc_2215 ( N_noxref_3_c_2222_n N_noxref_5_c_2628_n ) capacitor c=0.00687545f \
 //x=4.185 //y=2.59 //x2=3.33 //y2=2.08
cc_2216 ( N_noxref_3_c_2226_n N_noxref_5_c_2628_n ) capacitor c=0.0835358f \
 //x=4.07 //y=2.59 //x2=3.33 //y2=2.08
cc_2217 ( N_noxref_3_c_2227_n N_noxref_5_c_2628_n ) capacitor c=7.74334e-19 \
 //x=5.92 //y=2.08 //x2=3.33 //y2=2.08
cc_2218 ( N_noxref_3_c_2317_p N_noxref_5_c_2628_n ) capacitor c=0.0174995f \
 //x=3.29 //y=5.155 //x2=3.33 //y2=2.08
cc_2219 ( N_noxref_3_M67_noxref_g N_noxref_5_c_2643_n ) capacitor c=0.0178794f \
 //x=6.56 //y=6.02 //x2=7.135 //y2=5.155
cc_2220 ( N_noxref_3_c_2260_n N_noxref_5_c_2647_n ) capacitor c=3.10026e-19 \
 //x=3.985 //y=5.155 //x2=6.425 //y2=5.155
cc_2221 ( N_noxref_3_M66_noxref_g N_noxref_5_c_2647_n ) capacitor c=0.0213876f \
 //x=6.12 //y=6.02 //x2=6.425 //y2=5.155
cc_2222 ( N_noxref_3_c_2321_p N_noxref_5_c_2647_n ) capacitor c=0.00429591f \
 //x=6.485 //y=4.79 //x2=6.425 //y2=5.155
cc_2223 ( N_noxref_3_c_2223_n N_noxref_5_c_2657_n ) capacitor c=0.0192483f \
 //x=10.615 //y=2.59 //x2=8.88 //y2=3.33
cc_2224 ( N_noxref_3_c_2228_n N_noxref_5_c_2657_n ) capacitor c=0.0122828f \
 //x=10.73 //y=2.08 //x2=8.88 //y2=3.33
cc_2225 ( N_noxref_3_c_2256_n N_noxref_5_M64_noxref_g ) capacitor c=0.0184045f \
 //x=3.205 //y=5.155 //x2=3.07 //y2=6.02
cc_2226 ( N_noxref_3_M64_noxref_d N_noxref_5_M64_noxref_g ) capacitor \
 c=0.0180032f //x=3.145 //y=5.02 //x2=3.07 //y2=6.02
cc_2227 ( N_noxref_3_c_2260_n N_noxref_5_M65_noxref_g ) capacitor c=0.0205426f \
 //x=3.985 //y=5.155 //x2=3.51 //y2=6.02
cc_2228 ( N_noxref_3_M64_noxref_d N_noxref_5_M65_noxref_g ) capacitor \
 c=0.0194246f //x=3.145 //y=5.02 //x2=3.51 //y2=6.02
cc_2229 ( N_noxref_3_M2_noxref_d N_noxref_5_c_2711_n ) capacitor c=0.00217566f \
 //x=3.395 //y=0.915 //x2=3.32 //y2=0.915
cc_2230 ( N_noxref_3_M2_noxref_d N_noxref_5_c_2712_n ) capacitor c=0.0034598f \
 //x=3.395 //y=0.915 //x2=3.32 //y2=1.26
cc_2231 ( N_noxref_3_M2_noxref_d N_noxref_5_c_2713_n ) capacitor c=0.00546784f \
 //x=3.395 //y=0.915 //x2=3.32 //y2=1.57
cc_2232 ( N_noxref_3_M2_noxref_d N_noxref_5_c_2714_n ) capacitor c=0.00241102f \
 //x=3.395 //y=0.915 //x2=3.695 //y2=0.76
cc_2233 ( N_noxref_3_c_2225_n N_noxref_5_c_2715_n ) capacitor c=0.00371277f \
 //x=3.985 //y=1.665 //x2=3.695 //y2=1.415
cc_2234 ( N_noxref_3_M2_noxref_d N_noxref_5_c_2715_n ) capacitor c=0.0138621f \
 //x=3.395 //y=0.915 //x2=3.695 //y2=1.415
cc_2235 ( N_noxref_3_M2_noxref_d N_noxref_5_c_2717_n ) capacitor c=0.00219619f \
 //x=3.395 //y=0.915 //x2=3.85 //y2=0.915
cc_2236 ( N_noxref_3_c_2225_n N_noxref_5_c_2718_n ) capacitor c=0.00457401f \
 //x=3.985 //y=1.665 //x2=3.85 //y2=1.26
cc_2237 ( N_noxref_3_M2_noxref_d N_noxref_5_c_2718_n ) capacitor c=0.00603828f \
 //x=3.395 //y=0.915 //x2=3.85 //y2=1.26
cc_2238 ( N_noxref_3_c_2226_n N_noxref_5_c_2720_n ) capacitor c=0.00709342f \
 //x=4.07 //y=2.59 //x2=3.33 //y2=2.08
cc_2239 ( N_noxref_3_c_2226_n N_noxref_5_c_2721_n ) capacitor c=0.00283672f \
 //x=4.07 //y=2.59 //x2=3.33 //y2=1.915
cc_2240 ( N_noxref_3_M2_noxref_d N_noxref_5_c_2721_n ) capacitor c=0.00661782f \
 //x=3.395 //y=0.915 //x2=3.33 //y2=1.915
cc_2241 ( N_noxref_3_c_2260_n N_noxref_5_c_2723_n ) capacitor c=0.00201851f \
 //x=3.985 //y=5.155 //x2=3.33 //y2=4.7
cc_2242 ( N_noxref_3_c_2226_n N_noxref_5_c_2723_n ) capacitor c=0.013693f \
 //x=4.07 //y=2.59 //x2=3.33 //y2=4.7
cc_2243 ( N_noxref_3_c_2317_p N_noxref_5_c_2723_n ) capacitor c=0.00475729f \
 //x=3.29 //y=5.155 //x2=3.33 //y2=4.7
cc_2244 ( N_noxref_3_M67_noxref_g N_noxref_5_M66_noxref_d ) capacitor \
 c=0.0180032f //x=6.56 //y=6.02 //x2=6.195 //y2=5.02
cc_2245 ( N_noxref_3_c_2223_n N_noxref_7_c_3577_n ) capacitor c=0.0121818f \
 //x=10.615 //y=2.59 //x2=12.835 //y2=3.7
cc_2246 ( N_noxref_3_c_2228_n N_noxref_7_c_3577_n ) capacitor c=0.0197627f \
 //x=10.73 //y=2.08 //x2=12.835 //y2=3.7
cc_2247 ( N_noxref_3_c_2223_n N_noxref_7_c_3579_n ) capacitor c=5.84956e-19 \
 //x=10.615 //y=2.59 //x2=8.255 //y2=3.7
cc_2248 ( N_noxref_3_c_2223_n N_noxref_7_c_3527_n ) capacitor c=0.0203032f \
 //x=10.615 //y=2.59 //x2=8.14 //y2=2.08
cc_2249 ( N_noxref_3_c_2227_n N_noxref_7_c_3527_n ) capacitor c=0.00136793f \
 //x=5.92 //y=2.08 //x2=8.14 //y2=2.08
cc_2250 ( N_noxref_3_c_2228_n N_noxref_7_c_3527_n ) capacitor c=7.41683e-19 \
 //x=10.73 //y=2.08 //x2=8.14 //y2=2.08
cc_2251 ( N_noxref_3_c_2228_n N_noxref_7_c_3528_n ) capacitor c=0.00124614f \
 //x=10.73 //y=2.08 //x2=12.95 //y2=2.08
cc_2252 ( N_noxref_3_c_2221_n N_D_c_5277_n ) capacitor c=0.00327657f //x=5.805 \
 //y=2.59 //x2=29.855 //y2=4.07
cc_2253 ( N_noxref_3_c_2222_n N_D_c_5277_n ) capacitor c=3.66073e-19 //x=4.185 \
 //y=2.59 //x2=29.855 //y2=4.07
cc_2254 ( N_noxref_3_c_2223_n N_D_c_5277_n ) capacitor c=0.00875976f \
 //x=10.615 //y=2.59 //x2=29.855 //y2=4.07
cc_2255 ( N_noxref_3_c_2224_n N_D_c_5277_n ) capacitor c=2.46147e-19 //x=6.035 \
 //y=2.59 //x2=29.855 //y2=4.07
cc_2256 ( N_noxref_3_c_2250_n N_D_c_5277_n ) capacitor c=0.0244187f //x=2.325 \
 //y=5.155 //x2=29.855 //y2=4.07
cc_2257 ( N_noxref_3_c_2254_n N_D_c_5277_n ) capacitor c=0.0169078f //x=1.615 \
 //y=5.155 //x2=29.855 //y2=4.07
cc_2258 ( N_noxref_3_c_2260_n N_D_c_5277_n ) capacitor c=0.0138556f //x=3.985 \
 //y=5.155 //x2=29.855 //y2=4.07
cc_2259 ( N_noxref_3_c_2226_n N_D_c_5277_n ) capacitor c=0.0256324f //x=4.07 \
 //y=2.59 //x2=29.855 //y2=4.07
cc_2260 ( N_noxref_3_c_2227_n N_D_c_5277_n ) capacitor c=0.0257995f //x=5.92 \
 //y=2.08 //x2=29.855 //y2=4.07
cc_2261 ( N_noxref_3_c_2228_n N_D_c_5277_n ) capacitor c=0.0194977f //x=10.73 \
 //y=2.08 //x2=29.855 //y2=4.07
cc_2262 ( N_noxref_3_c_2279_n N_D_c_5277_n ) capacitor c=0.0116469f //x=6.195 \
 //y=4.79 //x2=29.855 //y2=4.07
cc_2263 ( N_noxref_3_c_2254_n N_D_M60_noxref_g ) capacitor c=0.0213876f \
 //x=1.615 //y=5.155 //x2=1.31 //y2=6.02
cc_2264 ( N_noxref_3_c_2250_n N_D_M61_noxref_g ) capacitor c=0.0178794f \
 //x=2.325 //y=5.155 //x2=1.75 //y2=6.02
cc_2265 ( N_noxref_3_M60_noxref_d N_D_M61_noxref_g ) capacitor c=0.0180032f \
 //x=1.385 //y=5.02 //x2=1.75 //y2=6.02
cc_2266 ( N_noxref_3_c_2254_n N_D_c_5376_n ) capacitor c=0.00429591f //x=1.615 \
 //y=5.155 //x2=1.675 //y2=4.79
cc_2267 ( N_noxref_3_c_2228_n N_CLK_c_6046_n ) capacitor c=0.0208709f \
 //x=10.73 //y=2.08 //x2=16.535 //y2=4.44
cc_2268 ( N_noxref_3_c_2281_n N_CLK_c_6046_n ) capacitor c=0.0166984f \
 //x=11.005 //y=4.79 //x2=16.535 //y2=4.44
cc_2269 ( N_noxref_3_c_2227_n N_CLK_c_6057_n ) capacitor c=0.00551083f \
 //x=5.92 //y=2.08 //x2=7.145 //y2=4.44
cc_2270 ( N_noxref_3_c_2223_n N_CLK_c_6040_n ) capacitor c=0.0213409f \
 //x=10.615 //y=2.59 //x2=7.03 //y2=2.08
cc_2271 ( N_noxref_3_c_2224_n N_CLK_c_6040_n ) capacitor c=9.95819e-19 \
 //x=6.035 //y=2.59 //x2=7.03 //y2=2.08
cc_2272 ( N_noxref_3_c_2226_n N_CLK_c_6040_n ) capacitor c=4.30656e-19 \
 //x=4.07 //y=2.59 //x2=7.03 //y2=2.08
cc_2273 ( N_noxref_3_c_2227_n N_CLK_c_6040_n ) capacitor c=0.0467743f //x=5.92 \
 //y=2.08 //x2=7.03 //y2=2.08
cc_2274 ( N_noxref_3_c_2233_n N_CLK_c_6040_n ) capacitor c=0.00210802f \
 //x=5.62 //y=1.915 //x2=7.03 //y2=2.08
cc_2275 ( N_noxref_3_c_2321_p N_CLK_c_6040_n ) capacitor c=0.00147352f \
 //x=6.485 //y=4.79 //x2=7.03 //y2=2.08
cc_2276 ( N_noxref_3_c_2279_n N_CLK_c_6040_n ) capacitor c=0.00141297f \
 //x=6.195 //y=4.79 //x2=7.03 //y2=2.08
cc_2277 ( N_noxref_3_M66_noxref_g N_CLK_M68_noxref_g ) capacitor c=0.0105869f \
 //x=6.12 //y=6.02 //x2=7 //y2=6.02
cc_2278 ( N_noxref_3_M67_noxref_g N_CLK_M68_noxref_g ) capacitor c=0.10632f \
 //x=6.56 //y=6.02 //x2=7 //y2=6.02
cc_2279 ( N_noxref_3_M67_noxref_g N_CLK_M69_noxref_g ) capacitor c=0.0101598f \
 //x=6.56 //y=6.02 //x2=7.44 //y2=6.02
cc_2280 ( N_noxref_3_c_2229_n N_CLK_c_6121_n ) capacitor c=5.72482e-19 \
 //x=5.62 //y=0.875 //x2=6.595 //y2=0.91
cc_2281 ( N_noxref_3_c_2231_n N_CLK_c_6121_n ) capacitor c=0.00149976f \
 //x=5.62 //y=1.22 //x2=6.595 //y2=0.91
cc_2282 ( N_noxref_3_c_2236_n N_CLK_c_6121_n ) capacitor c=0.0160123f //x=6.15 \
 //y=0.875 //x2=6.595 //y2=0.91
cc_2283 ( N_noxref_3_c_2232_n N_CLK_c_6124_n ) capacitor c=0.00111227f \
 //x=5.62 //y=1.53 //x2=6.595 //y2=1.22
cc_2284 ( N_noxref_3_c_2238_n N_CLK_c_6124_n ) capacitor c=0.0124075f //x=6.15 \
 //y=1.22 //x2=6.595 //y2=1.22
cc_2285 ( N_noxref_3_c_2236_n N_CLK_c_6126_n ) capacitor c=0.00103227f \
 //x=6.15 //y=0.875 //x2=7.12 //y2=0.91
cc_2286 ( N_noxref_3_c_2238_n N_CLK_c_6127_n ) capacitor c=0.0010154f //x=6.15 \
 //y=1.22 //x2=7.12 //y2=1.22
cc_2287 ( N_noxref_3_c_2238_n N_CLK_c_6128_n ) capacitor c=9.23422e-19 \
 //x=6.15 //y=1.22 //x2=7.12 //y2=1.45
cc_2288 ( N_noxref_3_c_2227_n N_CLK_c_6129_n ) capacitor c=0.00203769f \
 //x=5.92 //y=2.08 //x2=7.12 //y2=1.915
cc_2289 ( N_noxref_3_c_2233_n N_CLK_c_6129_n ) capacitor c=0.00834532f \
 //x=5.62 //y=1.915 //x2=7.12 //y2=1.915
cc_2290 ( N_noxref_3_c_2227_n N_CLK_c_6131_n ) capacitor c=0.00183762f \
 //x=5.92 //y=2.08 //x2=7.03 //y2=4.7
cc_2291 ( N_noxref_3_c_2321_p N_CLK_c_6131_n ) capacitor c=0.0168581f \
 //x=6.485 //y=4.79 //x2=7.03 //y2=4.7
cc_2292 ( N_noxref_3_c_2279_n N_CLK_c_6131_n ) capacitor c=0.00484466f \
 //x=6.195 //y=4.79 //x2=7.03 //y2=4.7
cc_2293 ( N_noxref_3_c_2221_n N_RN_c_7021_n ) capacitor c=0.143487f //x=5.805 \
 //y=2.59 //x2=17.645 //y2=2.22
cc_2294 ( N_noxref_3_c_2222_n N_RN_c_7021_n ) capacitor c=0.0291301f //x=4.185 \
 //y=2.59 //x2=17.645 //y2=2.22
cc_2295 ( N_noxref_3_c_2223_n N_RN_c_7021_n ) capacitor c=0.42762f //x=10.615 \
 //y=2.59 //x2=17.645 //y2=2.22
cc_2296 ( N_noxref_3_c_2224_n N_RN_c_7021_n ) capacitor c=0.0264401f //x=6.035 \
 //y=2.59 //x2=17.645 //y2=2.22
cc_2297 ( N_noxref_3_c_2396_p N_RN_c_7021_n ) capacitor c=0.016327f //x=3.67 \
 //y=1.665 //x2=17.645 //y2=2.22
cc_2298 ( N_noxref_3_c_2226_n N_RN_c_7021_n ) capacitor c=0.0215653f //x=4.07 \
 //y=2.59 //x2=17.645 //y2=2.22
cc_2299 ( N_noxref_3_c_2227_n N_RN_c_7021_n ) capacitor c=0.021104f //x=5.92 \
 //y=2.08 //x2=17.645 //y2=2.22
cc_2300 ( N_noxref_3_c_2228_n N_RN_c_7021_n ) capacitor c=0.021104f //x=10.73 \
 //y=2.08 //x2=17.645 //y2=2.22
cc_2301 ( N_noxref_3_c_2233_n N_RN_c_7021_n ) capacitor c=0.011987f //x=5.62 \
 //y=1.915 //x2=17.645 //y2=2.22
cc_2302 ( N_noxref_3_c_2243_n N_RN_c_7021_n ) capacitor c=0.011987f //x=10.43 \
 //y=1.915 //x2=17.645 //y2=2.22
cc_2303 ( N_noxref_3_c_2250_n N_RN_c_7088_n ) capacitor c=0.0148665f //x=2.325 \
 //y=5.155 //x2=2.22 //y2=2.08
cc_2304 ( N_noxref_3_c_2226_n N_RN_c_7088_n ) capacitor c=0.00309416f //x=4.07 \
 //y=2.59 //x2=2.22 //y2=2.08
cc_2305 ( N_noxref_3_c_2250_n N_RN_M62_noxref_g ) capacitor c=0.0166659f \
 //x=2.325 //y=5.155 //x2=2.19 //y2=6.02
cc_2306 ( N_noxref_3_M62_noxref_d N_RN_M62_noxref_g ) capacitor c=0.0180032f \
 //x=2.265 //y=5.02 //x2=2.19 //y2=6.02
cc_2307 ( N_noxref_3_c_2256_n N_RN_M63_noxref_g ) capacitor c=0.0184045f \
 //x=3.205 //y=5.155 //x2=2.63 //y2=6.02
cc_2308 ( N_noxref_3_M62_noxref_d N_RN_M63_noxref_g ) capacitor c=0.0180032f \
 //x=2.265 //y=5.02 //x2=2.63 //y2=6.02
cc_2309 ( N_noxref_3_c_2408_p N_RN_c_7161_n ) capacitor c=0.00427862f //x=2.41 \
 //y=5.155 //x2=2.555 //y2=4.79
cc_2310 ( N_noxref_3_c_2250_n N_RN_c_7162_n ) capacitor c=0.00322396f \
 //x=2.325 //y=5.155 //x2=2.22 //y2=4.7
cc_2311 ( N_noxref_3_c_2228_n N_SN_c_8183_n ) capacitor c=0.00526349f \
 //x=10.73 //y=2.08 //x2=11.955 //y2=2.96
cc_2312 ( N_noxref_3_c_2223_n N_SN_c_8145_n ) capacitor c=0.00311593f \
 //x=10.615 //y=2.59 //x2=11.84 //y2=2.08
cc_2313 ( N_noxref_3_c_2228_n N_SN_c_8145_n ) capacitor c=0.0436559f //x=10.73 \
 //y=2.08 //x2=11.84 //y2=2.08
cc_2314 ( N_noxref_3_c_2243_n N_SN_c_8145_n ) capacitor c=0.00210802f \
 //x=10.43 //y=1.915 //x2=11.84 //y2=2.08
cc_2315 ( N_noxref_3_c_2301_p N_SN_c_8145_n ) capacitor c=0.00147352f \
 //x=11.295 //y=4.79 //x2=11.84 //y2=2.08
cc_2316 ( N_noxref_3_c_2281_n N_SN_c_8145_n ) capacitor c=0.00142741f \
 //x=11.005 //y=4.79 //x2=11.84 //y2=2.08
cc_2317 ( N_noxref_3_M72_noxref_g N_SN_M74_noxref_g ) capacitor c=0.0105869f \
 //x=10.93 //y=6.02 //x2=11.81 //y2=6.02
cc_2318 ( N_noxref_3_M73_noxref_g N_SN_M74_noxref_g ) capacitor c=0.10632f \
 //x=11.37 //y=6.02 //x2=11.81 //y2=6.02
cc_2319 ( N_noxref_3_M73_noxref_g N_SN_M75_noxref_g ) capacitor c=0.0101598f \
 //x=11.37 //y=6.02 //x2=12.25 //y2=6.02
cc_2320 ( N_noxref_3_c_2239_n N_SN_c_8192_n ) capacitor c=5.72482e-19 \
 //x=10.43 //y=0.875 //x2=11.405 //y2=0.91
cc_2321 ( N_noxref_3_c_2241_n N_SN_c_8192_n ) capacitor c=0.00149976f \
 //x=10.43 //y=1.22 //x2=11.405 //y2=0.91
cc_2322 ( N_noxref_3_c_2246_n N_SN_c_8192_n ) capacitor c=0.0160123f //x=10.96 \
 //y=0.875 //x2=11.405 //y2=0.91
cc_2323 ( N_noxref_3_c_2242_n N_SN_c_8195_n ) capacitor c=0.00111227f \
 //x=10.43 //y=1.53 //x2=11.405 //y2=1.22
cc_2324 ( N_noxref_3_c_2248_n N_SN_c_8195_n ) capacitor c=0.0124075f //x=10.96 \
 //y=1.22 //x2=11.405 //y2=1.22
cc_2325 ( N_noxref_3_c_2246_n N_SN_c_8197_n ) capacitor c=0.00103227f \
 //x=10.96 //y=0.875 //x2=11.93 //y2=0.91
cc_2326 ( N_noxref_3_c_2248_n N_SN_c_8198_n ) capacitor c=0.0010154f //x=10.96 \
 //y=1.22 //x2=11.93 //y2=1.22
cc_2327 ( N_noxref_3_c_2248_n N_SN_c_8199_n ) capacitor c=9.23422e-19 \
 //x=10.96 //y=1.22 //x2=11.93 //y2=1.45
cc_2328 ( N_noxref_3_c_2228_n N_SN_c_8200_n ) capacitor c=0.00203769f \
 //x=10.73 //y=2.08 //x2=11.93 //y2=1.915
cc_2329 ( N_noxref_3_c_2243_n N_SN_c_8200_n ) capacitor c=0.00834532f \
 //x=10.43 //y=1.915 //x2=11.93 //y2=1.915
cc_2330 ( N_noxref_3_c_2228_n N_SN_c_8202_n ) capacitor c=0.00183762f \
 //x=10.73 //y=2.08 //x2=11.84 //y2=4.7
cc_2331 ( N_noxref_3_c_2301_p N_SN_c_8202_n ) capacitor c=0.0168581f \
 //x=11.295 //y=4.79 //x2=11.84 //y2=4.7
cc_2332 ( N_noxref_3_c_2281_n N_SN_c_8202_n ) capacitor c=0.00484466f \
 //x=11.005 //y=4.79 //x2=11.84 //y2=4.7
cc_2333 ( N_noxref_3_M2_noxref_d N_noxref_28_M0_noxref_s ) capacitor \
 c=0.00309936f //x=3.395 //y=0.915 //x2=0.455 //y2=0.375
cc_2334 ( N_noxref_3_c_2225_n N_noxref_29_c_10596_n ) capacitor c=0.00457167f \
 //x=3.985 //y=1.665 //x2=3.985 //y2=0.54
cc_2335 ( N_noxref_3_M2_noxref_d N_noxref_29_c_10596_n ) capacitor \
 c=0.0115903f //x=3.395 //y=0.915 //x2=3.985 //y2=0.54
cc_2336 ( N_noxref_3_c_2396_p N_noxref_29_c_10606_n ) capacitor c=0.0200405f \
 //x=3.67 //y=1.665 //x2=3.1 //y2=0.995
cc_2337 ( N_noxref_3_M2_noxref_d N_noxref_29_M1_noxref_d ) capacitor \
 c=5.27807e-19 //x=3.395 //y=0.915 //x2=1.86 //y2=0.91
cc_2338 ( N_noxref_3_c_2225_n N_noxref_29_M2_noxref_s ) capacitor c=0.0184051f \
 //x=3.985 //y=1.665 //x2=2.965 //y2=0.375
cc_2339 ( N_noxref_3_M2_noxref_d N_noxref_29_M2_noxref_s ) capacitor \
 c=0.0426368f //x=3.395 //y=0.915 //x2=2.965 //y2=0.375
cc_2340 ( N_noxref_3_c_2225_n N_noxref_30_c_10658_n ) capacitor c=3.84569e-19 \
 //x=3.985 //y=1.665 //x2=5.4 //y2=1.505
cc_2341 ( N_noxref_3_c_2233_n N_noxref_30_c_10658_n ) capacitor c=0.0034165f \
 //x=5.62 //y=1.915 //x2=5.4 //y2=1.505
cc_2342 ( N_noxref_3_c_2227_n N_noxref_30_c_10643_n ) capacitor c=0.0119952f \
 //x=5.92 //y=2.08 //x2=6.285 //y2=1.59
cc_2343 ( N_noxref_3_c_2232_n N_noxref_30_c_10643_n ) capacitor c=0.00697148f \
 //x=5.62 //y=1.53 //x2=6.285 //y2=1.59
cc_2344 ( N_noxref_3_c_2233_n N_noxref_30_c_10643_n ) capacitor c=0.0204849f \
 //x=5.62 //y=1.915 //x2=6.285 //y2=1.59
cc_2345 ( N_noxref_3_c_2235_n N_noxref_30_c_10643_n ) capacitor c=0.00610316f \
 //x=5.995 //y=1.375 //x2=6.285 //y2=1.59
cc_2346 ( N_noxref_3_c_2238_n N_noxref_30_c_10643_n ) capacitor c=0.00698822f \
 //x=6.15 //y=1.22 //x2=6.285 //y2=1.59
cc_2347 ( N_noxref_3_c_2229_n N_noxref_30_M3_noxref_s ) capacitor c=0.0327271f \
 //x=5.62 //y=0.875 //x2=5.265 //y2=0.375
cc_2348 ( N_noxref_3_c_2232_n N_noxref_30_M3_noxref_s ) capacitor \
 c=7.99997e-19 //x=5.62 //y=1.53 //x2=5.265 //y2=0.375
cc_2349 ( N_noxref_3_c_2233_n N_noxref_30_M3_noxref_s ) capacitor \
 c=0.00122123f //x=5.62 //y=1.915 //x2=5.265 //y2=0.375
cc_2350 ( N_noxref_3_c_2236_n N_noxref_30_M3_noxref_s ) capacitor c=0.0121427f \
 //x=6.15 //y=0.875 //x2=5.265 //y2=0.375
cc_2351 ( N_noxref_3_M2_noxref_d N_noxref_30_M3_noxref_s ) capacitor \
 c=2.55333e-19 //x=3.395 //y=0.915 //x2=5.265 //y2=0.375
cc_2352 ( N_noxref_3_c_2243_n N_noxref_32_c_10759_n ) capacitor c=0.0034165f \
 //x=10.43 //y=1.915 //x2=10.21 //y2=1.505
cc_2353 ( N_noxref_3_c_2228_n N_noxref_32_c_10744_n ) capacitor c=0.0115578f \
 //x=10.73 //y=2.08 //x2=11.095 //y2=1.59
cc_2354 ( N_noxref_3_c_2242_n N_noxref_32_c_10744_n ) capacitor c=0.00697148f \
 //x=10.43 //y=1.53 //x2=11.095 //y2=1.59
cc_2355 ( N_noxref_3_c_2243_n N_noxref_32_c_10744_n ) capacitor c=0.0204849f \
 //x=10.43 //y=1.915 //x2=11.095 //y2=1.59
cc_2356 ( N_noxref_3_c_2245_n N_noxref_32_c_10744_n ) capacitor c=0.00610316f \
 //x=10.805 //y=1.375 //x2=11.095 //y2=1.59
cc_2357 ( N_noxref_3_c_2248_n N_noxref_32_c_10744_n ) capacitor c=0.00698822f \
 //x=10.96 //y=1.22 //x2=11.095 //y2=1.59
cc_2358 ( N_noxref_3_c_2239_n N_noxref_32_M6_noxref_s ) capacitor c=0.0327271f \
 //x=10.43 //y=0.875 //x2=10.075 //y2=0.375
cc_2359 ( N_noxref_3_c_2242_n N_noxref_32_M6_noxref_s ) capacitor \
 c=7.99997e-19 //x=10.43 //y=1.53 //x2=10.075 //y2=0.375
cc_2360 ( N_noxref_3_c_2243_n N_noxref_32_M6_noxref_s ) capacitor \
 c=0.00122123f //x=10.43 //y=1.915 //x2=10.075 //y2=0.375
cc_2361 ( N_noxref_3_c_2246_n N_noxref_32_M6_noxref_s ) capacitor c=0.0121427f \
 //x=10.96 //y=0.875 //x2=10.075 //y2=0.375
cc_2362 ( N_noxref_4_c_2461_n N_noxref_5_c_2627_n ) capacitor c=0.0119023f \
 //x=15.425 //y=2.59 //x2=20.235 //y2=3.33
cc_2363 ( N_noxref_4_c_2462_n N_noxref_5_c_2627_n ) capacitor c=8.87672e-19 \
 //x=13.805 //y=2.59 //x2=20.235 //y2=3.33
cc_2364 ( N_noxref_4_c_2464_n N_noxref_5_c_2627_n ) capacitor c=0.018769f \
 //x=13.69 //y=2.59 //x2=20.235 //y2=3.33
cc_2365 ( N_noxref_4_c_2465_n N_noxref_5_c_2627_n ) capacitor c=0.0198064f \
 //x=15.54 //y=2.08 //x2=20.235 //y2=3.33
cc_2366 ( N_noxref_4_c_2481_n N_noxref_5_c_2653_n ) capacitor c=3.10026e-19 \
 //x=11.235 //y=5.155 //x2=8.795 //y2=5.155
cc_2367 ( N_noxref_4_c_2464_n N_noxref_7_c_3584_n ) capacitor c=0.0187698f \
 //x=13.69 //y=2.59 //x2=18.385 //y2=3.7
cc_2368 ( N_noxref_4_c_2465_n N_noxref_7_c_3584_n ) capacitor c=0.0197889f \
 //x=15.54 //y=2.08 //x2=18.385 //y2=3.7
cc_2369 ( N_noxref_4_c_2464_n N_noxref_7_c_3586_n ) capacitor c=0.00179385f \
 //x=13.69 //y=2.59 //x2=13.065 //y2=3.7
cc_2370 ( N_noxref_4_c_2462_n N_noxref_7_c_3528_n ) capacitor c=0.00456439f \
 //x=13.805 //y=2.59 //x2=12.95 //y2=2.08
cc_2371 ( N_noxref_4_c_2464_n N_noxref_7_c_3528_n ) capacitor c=0.0769512f \
 //x=13.69 //y=2.59 //x2=12.95 //y2=2.08
cc_2372 ( N_noxref_4_c_2465_n N_noxref_7_c_3528_n ) capacitor c=5.32619e-19 \
 //x=15.54 //y=2.08 //x2=12.95 //y2=2.08
cc_2373 ( N_noxref_4_c_2532_p N_noxref_7_c_3528_n ) capacitor c=0.016476f \
 //x=12.91 //y=5.155 //x2=12.95 //y2=2.08
cc_2374 ( N_noxref_4_M79_noxref_g N_noxref_7_c_3534_n ) capacitor c=0.0168349f \
 //x=16.18 //y=6.02 //x2=16.755 //y2=5.155
cc_2375 ( N_noxref_4_c_2487_n N_noxref_7_c_3538_n ) capacitor c=3.10026e-19 \
 //x=13.605 //y=5.155 //x2=16.045 //y2=5.155
cc_2376 ( N_noxref_4_M78_noxref_g N_noxref_7_c_3538_n ) capacitor c=0.0213876f \
 //x=15.74 //y=6.02 //x2=16.045 //y2=5.155
cc_2377 ( N_noxref_4_c_2536_p N_noxref_7_c_3538_n ) capacitor c=0.00428486f \
 //x=16.105 //y=4.79 //x2=16.045 //y2=5.155
cc_2378 ( N_noxref_4_c_2483_n N_noxref_7_M76_noxref_g ) capacitor c=0.01736f \
 //x=12.825 //y=5.155 //x2=12.69 //y2=6.02
cc_2379 ( N_noxref_4_M76_noxref_d N_noxref_7_M76_noxref_g ) capacitor \
 c=0.0180032f //x=12.765 //y=5.02 //x2=12.69 //y2=6.02
cc_2380 ( N_noxref_4_c_2487_n N_noxref_7_M77_noxref_g ) capacitor c=0.0194981f \
 //x=13.605 //y=5.155 //x2=13.13 //y2=6.02
cc_2381 ( N_noxref_4_M76_noxref_d N_noxref_7_M77_noxref_g ) capacitor \
 c=0.0194246f //x=12.765 //y=5.02 //x2=13.13 //y2=6.02
cc_2382 ( N_noxref_4_M8_noxref_d N_noxref_7_c_3599_n ) capacitor c=0.00217566f \
 //x=13.015 //y=0.915 //x2=12.94 //y2=0.915
cc_2383 ( N_noxref_4_M8_noxref_d N_noxref_7_c_3600_n ) capacitor c=0.0034598f \
 //x=13.015 //y=0.915 //x2=12.94 //y2=1.26
cc_2384 ( N_noxref_4_M8_noxref_d N_noxref_7_c_3601_n ) capacitor c=0.00546784f \
 //x=13.015 //y=0.915 //x2=12.94 //y2=1.57
cc_2385 ( N_noxref_4_M8_noxref_d N_noxref_7_c_3602_n ) capacitor c=0.00241102f \
 //x=13.015 //y=0.915 //x2=13.315 //y2=0.76
cc_2386 ( N_noxref_4_c_2463_n N_noxref_7_c_3603_n ) capacitor c=0.00371277f \
 //x=13.605 //y=1.665 //x2=13.315 //y2=1.415
cc_2387 ( N_noxref_4_M8_noxref_d N_noxref_7_c_3603_n ) capacitor c=0.0138621f \
 //x=13.015 //y=0.915 //x2=13.315 //y2=1.415
cc_2388 ( N_noxref_4_M8_noxref_d N_noxref_7_c_3605_n ) capacitor c=0.00219619f \
 //x=13.015 //y=0.915 //x2=13.47 //y2=0.915
cc_2389 ( N_noxref_4_c_2463_n N_noxref_7_c_3606_n ) capacitor c=0.00457401f \
 //x=13.605 //y=1.665 //x2=13.47 //y2=1.26
cc_2390 ( N_noxref_4_M8_noxref_d N_noxref_7_c_3606_n ) capacitor c=0.00603828f \
 //x=13.015 //y=0.915 //x2=13.47 //y2=1.26
cc_2391 ( N_noxref_4_c_2464_n N_noxref_7_c_3608_n ) capacitor c=0.00731987f \
 //x=13.69 //y=2.59 //x2=12.95 //y2=2.08
cc_2392 ( N_noxref_4_c_2464_n N_noxref_7_c_3609_n ) capacitor c=0.00283672f \
 //x=13.69 //y=2.59 //x2=12.95 //y2=1.915
cc_2393 ( N_noxref_4_M8_noxref_d N_noxref_7_c_3609_n ) capacitor c=0.00661782f \
 //x=13.015 //y=0.915 //x2=12.95 //y2=1.915
cc_2394 ( N_noxref_4_c_2487_n N_noxref_7_c_3611_n ) capacitor c=0.00201851f \
 //x=13.605 //y=5.155 //x2=12.95 //y2=4.7
cc_2395 ( N_noxref_4_c_2464_n N_noxref_7_c_3611_n ) capacitor c=0.013693f \
 //x=13.69 //y=2.59 //x2=12.95 //y2=4.7
cc_2396 ( N_noxref_4_c_2532_p N_noxref_7_c_3611_n ) capacitor c=0.00475601f \
 //x=12.91 //y=5.155 //x2=12.95 //y2=4.7
cc_2397 ( N_noxref_4_M79_noxref_g N_noxref_7_M78_noxref_d ) capacitor \
 c=0.0180032f //x=16.18 //y=6.02 //x2=15.815 //y2=5.02
cc_2398 ( N_noxref_4_c_2464_n N_D_c_5277_n ) capacitor c=0.0181982f //x=13.69 \
 //y=2.59 //x2=29.855 //y2=4.07
cc_2399 ( N_noxref_4_c_2465_n N_D_c_5277_n ) capacitor c=0.019517f //x=15.54 \
 //y=2.08 //x2=29.855 //y2=4.07
cc_2400 ( N_noxref_4_c_2477_n N_CLK_c_6046_n ) capacitor c=0.032141f \
 //x=11.945 //y=5.155 //x2=16.535 //y2=4.44
cc_2401 ( N_noxref_4_c_2481_n N_CLK_c_6046_n ) capacitor c=0.0230136f \
 //x=11.235 //y=5.155 //x2=16.535 //y2=4.44
cc_2402 ( N_noxref_4_c_2487_n N_CLK_c_6046_n ) capacitor c=0.0183122f \
 //x=13.605 //y=5.155 //x2=16.535 //y2=4.44
cc_2403 ( N_noxref_4_c_2464_n N_CLK_c_6046_n ) capacitor c=0.0210274f \
 //x=13.69 //y=2.59 //x2=16.535 //y2=4.44
cc_2404 ( N_noxref_4_c_2465_n N_CLK_c_6046_n ) capacitor c=0.0208709f \
 //x=15.54 //y=2.08 //x2=16.535 //y2=4.44
cc_2405 ( N_noxref_4_c_2499_n N_CLK_c_6046_n ) capacitor c=0.0166984f \
 //x=15.815 //y=4.79 //x2=16.535 //y2=4.44
cc_2406 ( N_noxref_4_c_2465_n N_CLK_c_6067_n ) capacitor c=0.00153281f \
 //x=15.54 //y=2.08 //x2=16.765 //y2=4.44
cc_2407 ( N_noxref_4_c_2461_n N_CLK_c_6041_n ) capacitor c=0.00520283f \
 //x=15.425 //y=2.59 //x2=16.65 //y2=2.08
cc_2408 ( N_noxref_4_c_2464_n N_CLK_c_6041_n ) capacitor c=2.96936e-19 \
 //x=13.69 //y=2.59 //x2=16.65 //y2=2.08
cc_2409 ( N_noxref_4_c_2465_n N_CLK_c_6041_n ) capacitor c=0.0422272f \
 //x=15.54 //y=2.08 //x2=16.65 //y2=2.08
cc_2410 ( N_noxref_4_c_2470_n N_CLK_c_6041_n ) capacitor c=0.00210802f \
 //x=15.24 //y=1.915 //x2=16.65 //y2=2.08
cc_2411 ( N_noxref_4_c_2536_p N_CLK_c_6041_n ) capacitor c=0.00147352f \
 //x=16.105 //y=4.79 //x2=16.65 //y2=2.08
cc_2412 ( N_noxref_4_c_2499_n N_CLK_c_6041_n ) capacitor c=0.00141297f \
 //x=15.815 //y=4.79 //x2=16.65 //y2=2.08
cc_2413 ( N_noxref_4_M78_noxref_g N_CLK_M80_noxref_g ) capacitor c=0.0105869f \
 //x=15.74 //y=6.02 //x2=16.62 //y2=6.02
cc_2414 ( N_noxref_4_M79_noxref_g N_CLK_M80_noxref_g ) capacitor c=0.10632f \
 //x=16.18 //y=6.02 //x2=16.62 //y2=6.02
cc_2415 ( N_noxref_4_M79_noxref_g N_CLK_M81_noxref_g ) capacitor c=0.0101598f \
 //x=16.18 //y=6.02 //x2=17.06 //y2=6.02
cc_2416 ( N_noxref_4_c_2466_n N_CLK_c_6150_n ) capacitor c=5.72482e-19 \
 //x=15.24 //y=0.875 //x2=16.215 //y2=0.91
cc_2417 ( N_noxref_4_c_2468_n N_CLK_c_6150_n ) capacitor c=0.00149976f \
 //x=15.24 //y=1.22 //x2=16.215 //y2=0.91
cc_2418 ( N_noxref_4_c_2473_n N_CLK_c_6150_n ) capacitor c=0.0160123f \
 //x=15.77 //y=0.875 //x2=16.215 //y2=0.91
cc_2419 ( N_noxref_4_c_2469_n N_CLK_c_6153_n ) capacitor c=0.00111227f \
 //x=15.24 //y=1.53 //x2=16.215 //y2=1.22
cc_2420 ( N_noxref_4_c_2475_n N_CLK_c_6153_n ) capacitor c=0.0124075f \
 //x=15.77 //y=1.22 //x2=16.215 //y2=1.22
cc_2421 ( N_noxref_4_c_2473_n N_CLK_c_6155_n ) capacitor c=0.00103227f \
 //x=15.77 //y=0.875 //x2=16.74 //y2=0.91
cc_2422 ( N_noxref_4_c_2475_n N_CLK_c_6156_n ) capacitor c=0.0010154f \
 //x=15.77 //y=1.22 //x2=16.74 //y2=1.22
cc_2423 ( N_noxref_4_c_2475_n N_CLK_c_6157_n ) capacitor c=9.23422e-19 \
 //x=15.77 //y=1.22 //x2=16.74 //y2=1.45
cc_2424 ( N_noxref_4_c_2465_n N_CLK_c_6158_n ) capacitor c=0.00203769f \
 //x=15.54 //y=2.08 //x2=16.74 //y2=1.915
cc_2425 ( N_noxref_4_c_2470_n N_CLK_c_6158_n ) capacitor c=0.00834532f \
 //x=15.24 //y=1.915 //x2=16.74 //y2=1.915
cc_2426 ( N_noxref_4_c_2465_n N_CLK_c_6160_n ) capacitor c=0.00183762f \
 //x=15.54 //y=2.08 //x2=16.65 //y2=4.7
cc_2427 ( N_noxref_4_c_2536_p N_CLK_c_6160_n ) capacitor c=0.0168581f \
 //x=16.105 //y=4.79 //x2=16.65 //y2=4.7
cc_2428 ( N_noxref_4_c_2499_n N_CLK_c_6160_n ) capacitor c=0.00484466f \
 //x=15.815 //y=4.79 //x2=16.65 //y2=4.7
cc_2429 ( N_noxref_4_c_2461_n N_RN_c_7021_n ) capacitor c=0.172592f //x=15.425 \
 //y=2.59 //x2=17.645 //y2=2.22
cc_2430 ( N_noxref_4_c_2462_n N_RN_c_7021_n ) capacitor c=0.0291301f \
 //x=13.805 //y=2.59 //x2=17.645 //y2=2.22
cc_2431 ( N_noxref_4_c_2590_p N_RN_c_7021_n ) capacitor c=0.016327f //x=13.29 \
 //y=1.665 //x2=17.645 //y2=2.22
cc_2432 ( N_noxref_4_c_2464_n N_RN_c_7021_n ) capacitor c=0.0215653f //x=13.69 \
 //y=2.59 //x2=17.645 //y2=2.22
cc_2433 ( N_noxref_4_c_2465_n N_RN_c_7021_n ) capacitor c=0.021104f //x=15.54 \
 //y=2.08 //x2=17.645 //y2=2.22
cc_2434 ( N_noxref_4_c_2470_n N_RN_c_7021_n ) capacitor c=0.011987f //x=15.24 \
 //y=1.915 //x2=17.645 //y2=2.22
cc_2435 ( N_noxref_4_c_2465_n N_RN_c_7089_n ) capacitor c=0.00107158f \
 //x=15.54 //y=2.08 //x2=17.76 //y2=2.08
cc_2436 ( N_noxref_4_c_2461_n N_SN_c_8129_n ) capacitor c=0.172781f //x=15.425 \
 //y=2.59 //x2=26.155 //y2=2.96
cc_2437 ( N_noxref_4_c_2462_n N_SN_c_8129_n ) capacitor c=0.0293832f \
 //x=13.805 //y=2.59 //x2=26.155 //y2=2.96
cc_2438 ( N_noxref_4_c_2464_n N_SN_c_8129_n ) capacitor c=0.0206007f //x=13.69 \
 //y=2.59 //x2=26.155 //y2=2.96
cc_2439 ( N_noxref_4_c_2465_n N_SN_c_8129_n ) capacitor c=0.0216195f //x=15.54 \
 //y=2.08 //x2=26.155 //y2=2.96
cc_2440 ( N_noxref_4_c_2477_n N_SN_c_8145_n ) capacitor c=0.0146f //x=11.945 \
 //y=5.155 //x2=11.84 //y2=2.08
cc_2441 ( N_noxref_4_c_2464_n N_SN_c_8145_n ) capacitor c=0.00240615f \
 //x=13.69 //y=2.59 //x2=11.84 //y2=2.08
cc_2442 ( N_noxref_4_c_2477_n N_SN_M74_noxref_g ) capacitor c=0.0165266f \
 //x=11.945 //y=5.155 //x2=11.81 //y2=6.02
cc_2443 ( N_noxref_4_M74_noxref_d N_SN_M74_noxref_g ) capacitor c=0.0180032f \
 //x=11.885 //y=5.02 //x2=11.81 //y2=6.02
cc_2444 ( N_noxref_4_c_2483_n N_SN_M75_noxref_g ) capacitor c=0.01736f \
 //x=12.825 //y=5.155 //x2=12.25 //y2=6.02
cc_2445 ( N_noxref_4_M74_noxref_d N_SN_M75_noxref_g ) capacitor c=0.0180032f \
 //x=11.885 //y=5.02 //x2=12.25 //y2=6.02
cc_2446 ( N_noxref_4_c_2605_p N_SN_c_8215_n ) capacitor c=0.00426767f \
 //x=12.03 //y=5.155 //x2=12.175 //y2=4.79
cc_2447 ( N_noxref_4_c_2477_n N_SN_c_8202_n ) capacitor c=0.00322054f \
 //x=11.945 //y=5.155 //x2=11.84 //y2=4.7
cc_2448 ( N_noxref_4_M8_noxref_d N_noxref_32_M6_noxref_s ) capacitor \
 c=0.00309936f //x=13.015 //y=0.915 //x2=10.075 //y2=0.375
cc_2449 ( N_noxref_4_c_2463_n N_noxref_33_c_10798_n ) capacitor c=0.00457167f \
 //x=13.605 //y=1.665 //x2=13.605 //y2=0.54
cc_2450 ( N_noxref_4_M8_noxref_d N_noxref_33_c_10798_n ) capacitor \
 c=0.0115903f //x=13.015 //y=0.915 //x2=13.605 //y2=0.54
cc_2451 ( N_noxref_4_c_2590_p N_noxref_33_c_10808_n ) capacitor c=0.0200405f \
 //x=13.29 //y=1.665 //x2=12.72 //y2=0.995
cc_2452 ( N_noxref_4_M8_noxref_d N_noxref_33_M7_noxref_d ) capacitor \
 c=5.27807e-19 //x=13.015 //y=0.915 //x2=11.48 //y2=0.91
cc_2453 ( N_noxref_4_c_2463_n N_noxref_33_M8_noxref_s ) capacitor c=0.0184051f \
 //x=13.605 //y=1.665 //x2=12.585 //y2=0.375
cc_2454 ( N_noxref_4_M8_noxref_d N_noxref_33_M8_noxref_s ) capacitor \
 c=0.0426368f //x=13.015 //y=0.915 //x2=12.585 //y2=0.375
cc_2455 ( N_noxref_4_c_2463_n N_noxref_34_c_10860_n ) capacitor c=3.84569e-19 \
 //x=13.605 //y=1.665 //x2=15.02 //y2=1.505
cc_2456 ( N_noxref_4_c_2470_n N_noxref_34_c_10860_n ) capacitor c=0.0034165f \
 //x=15.24 //y=1.915 //x2=15.02 //y2=1.505
cc_2457 ( N_noxref_4_c_2465_n N_noxref_34_c_10845_n ) capacitor c=0.0115578f \
 //x=15.54 //y=2.08 //x2=15.905 //y2=1.59
cc_2458 ( N_noxref_4_c_2469_n N_noxref_34_c_10845_n ) capacitor c=0.00697148f \
 //x=15.24 //y=1.53 //x2=15.905 //y2=1.59
cc_2459 ( N_noxref_4_c_2470_n N_noxref_34_c_10845_n ) capacitor c=0.0204849f \
 //x=15.24 //y=1.915 //x2=15.905 //y2=1.59
cc_2460 ( N_noxref_4_c_2472_n N_noxref_34_c_10845_n ) capacitor c=0.00610316f \
 //x=15.615 //y=1.375 //x2=15.905 //y2=1.59
cc_2461 ( N_noxref_4_c_2475_n N_noxref_34_c_10845_n ) capacitor c=0.00698822f \
 //x=15.77 //y=1.22 //x2=15.905 //y2=1.59
cc_2462 ( N_noxref_4_c_2466_n N_noxref_34_M9_noxref_s ) capacitor c=0.0327271f \
 //x=15.24 //y=0.875 //x2=14.885 //y2=0.375
cc_2463 ( N_noxref_4_c_2469_n N_noxref_34_M9_noxref_s ) capacitor \
 c=7.99997e-19 //x=15.24 //y=1.53 //x2=14.885 //y2=0.375
cc_2464 ( N_noxref_4_c_2470_n N_noxref_34_M9_noxref_s ) capacitor \
 c=0.00122123f //x=15.24 //y=1.915 //x2=14.885 //y2=0.375
cc_2465 ( N_noxref_4_c_2473_n N_noxref_34_M9_noxref_s ) capacitor c=0.0121427f \
 //x=15.77 //y=0.875 //x2=14.885 //y2=0.375
cc_2466 ( N_noxref_4_M8_noxref_d N_noxref_34_M9_noxref_s ) capacitor \
 c=2.55333e-19 //x=13.015 //y=0.915 //x2=14.885 //y2=0.375
cc_2467 ( N_noxref_5_M85_noxref_g N_noxref_6_c_3016_n ) capacitor c=0.0168349f \
 //x=20.99 //y=6.02 //x2=21.565 //y2=5.155
cc_2468 ( N_noxref_5_M84_noxref_g N_noxref_6_c_3020_n ) capacitor c=0.0213876f \
 //x=20.55 //y=6.02 //x2=20.855 //y2=5.155
cc_2469 ( N_noxref_5_c_2734_p N_noxref_6_c_3020_n ) capacitor c=0.00428486f \
 //x=20.915 //y=4.79 //x2=20.855 //y2=5.155
cc_2470 ( N_noxref_5_M85_noxref_g N_noxref_6_M84_noxref_d ) capacitor \
 c=0.0180032f //x=20.99 //y=6.02 //x2=20.625 //y2=5.02
cc_2471 ( N_noxref_5_c_2626_n N_noxref_7_c_3577_n ) capacitor c=0.0446157f \
 //x=8.765 //y=3.33 //x2=12.835 //y2=3.7
cc_2472 ( N_noxref_5_c_2627_n N_noxref_7_c_3577_n ) capacitor c=0.340407f \
 //x=20.235 //y=3.33 //x2=12.835 //y2=3.7
cc_2473 ( N_noxref_5_c_2695_n N_noxref_7_c_3577_n ) capacitor c=0.0268386f \
 //x=8.995 //y=3.33 //x2=12.835 //y2=3.7
cc_2474 ( N_noxref_5_c_2657_n N_noxref_7_c_3577_n ) capacitor c=0.0205782f \
 //x=8.88 //y=3.33 //x2=12.835 //y2=3.7
cc_2475 ( N_noxref_5_c_2626_n N_noxref_7_c_3579_n ) capacitor c=0.029444f \
 //x=8.765 //y=3.33 //x2=8.255 //y2=3.7
cc_2476 ( N_noxref_5_c_2657_n N_noxref_7_c_3579_n ) capacitor c=0.00179385f \
 //x=8.88 //y=3.33 //x2=8.255 //y2=3.7
cc_2477 ( N_noxref_5_c_2627_n N_noxref_7_c_3584_n ) capacitor c=0.468734f \
 //x=20.235 //y=3.33 //x2=18.385 //y2=3.7
cc_2478 ( N_noxref_5_c_2627_n N_noxref_7_c_3586_n ) capacitor c=0.026734f \
 //x=20.235 //y=3.33 //x2=13.065 //y2=3.7
cc_2479 ( N_noxref_5_c_2627_n N_noxref_7_c_3623_n ) capacitor c=0.176086f \
 //x=20.235 //y=3.33 //x2=27.265 //y2=3.7
cc_2480 ( N_noxref_5_c_2630_n N_noxref_7_c_3623_n ) capacitor c=0.0215974f \
 //x=20.35 //y=2.08 //x2=27.265 //y2=3.7
cc_2481 ( N_noxref_5_c_2627_n N_noxref_7_c_3625_n ) capacitor c=0.0268461f \
 //x=20.235 //y=3.33 //x2=18.615 //y2=3.7
cc_2482 ( N_noxref_5_c_2630_n N_noxref_7_c_3625_n ) capacitor c=7.01366e-19 \
 //x=20.35 //y=2.08 //x2=18.615 //y2=3.7
cc_2483 ( N_noxref_5_c_2626_n N_noxref_7_c_3527_n ) capacitor c=0.0221941f \
 //x=8.765 //y=3.33 //x2=8.14 //y2=2.08
cc_2484 ( N_noxref_5_c_2695_n N_noxref_7_c_3527_n ) capacitor c=0.00179385f \
 //x=8.995 //y=3.33 //x2=8.14 //y2=2.08
cc_2485 ( N_noxref_5_c_2657_n N_noxref_7_c_3527_n ) capacitor c=0.0777866f \
 //x=8.88 //y=3.33 //x2=8.14 //y2=2.08
cc_2486 ( N_noxref_5_c_2751_p N_noxref_7_c_3527_n ) capacitor c=0.016476f \
 //x=8.1 //y=5.155 //x2=8.14 //y2=2.08
cc_2487 ( N_noxref_5_c_2627_n N_noxref_7_c_3528_n ) capacitor c=0.0198536f \
 //x=20.235 //y=3.33 //x2=12.95 //y2=2.08
cc_2488 ( N_noxref_5_c_2627_n N_noxref_7_c_3548_n ) capacitor c=0.0212788f \
 //x=20.235 //y=3.33 //x2=18.5 //y2=3.7
cc_2489 ( N_noxref_5_c_2630_n N_noxref_7_c_3548_n ) capacitor c=0.0105909f \
 //x=20.35 //y=2.08 //x2=18.5 //y2=3.7
cc_2490 ( N_noxref_5_c_2649_n N_noxref_7_M70_noxref_g ) capacitor c=0.01736f \
 //x=8.015 //y=5.155 //x2=7.88 //y2=6.02
cc_2491 ( N_noxref_5_M70_noxref_d N_noxref_7_M70_noxref_g ) capacitor \
 c=0.0180032f //x=7.955 //y=5.02 //x2=7.88 //y2=6.02
cc_2492 ( N_noxref_5_c_2653_n N_noxref_7_M71_noxref_g ) capacitor c=0.0194981f \
 //x=8.795 //y=5.155 //x2=8.32 //y2=6.02
cc_2493 ( N_noxref_5_M70_noxref_d N_noxref_7_M71_noxref_g ) capacitor \
 c=0.0194246f //x=7.955 //y=5.02 //x2=8.32 //y2=6.02
cc_2494 ( N_noxref_5_M5_noxref_d N_noxref_7_c_3638_n ) capacitor c=0.00217566f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=0.915
cc_2495 ( N_noxref_5_M5_noxref_d N_noxref_7_c_3639_n ) capacitor c=0.0034598f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=1.26
cc_2496 ( N_noxref_5_M5_noxref_d N_noxref_7_c_3640_n ) capacitor c=0.00546784f \
 //x=8.205 //y=0.915 //x2=8.13 //y2=1.57
cc_2497 ( N_noxref_5_M5_noxref_d N_noxref_7_c_3641_n ) capacitor c=0.00241102f \
 //x=8.205 //y=0.915 //x2=8.505 //y2=0.76
cc_2498 ( N_noxref_5_c_2629_n N_noxref_7_c_3642_n ) capacitor c=0.00371277f \
 //x=8.795 //y=1.665 //x2=8.505 //y2=1.415
cc_2499 ( N_noxref_5_M5_noxref_d N_noxref_7_c_3642_n ) capacitor c=0.0138621f \
 //x=8.205 //y=0.915 //x2=8.505 //y2=1.415
cc_2500 ( N_noxref_5_M5_noxref_d N_noxref_7_c_3644_n ) capacitor c=0.00219619f \
 //x=8.205 //y=0.915 //x2=8.66 //y2=0.915
cc_2501 ( N_noxref_5_c_2629_n N_noxref_7_c_3645_n ) capacitor c=0.00457401f \
 //x=8.795 //y=1.665 //x2=8.66 //y2=1.26
cc_2502 ( N_noxref_5_M5_noxref_d N_noxref_7_c_3645_n ) capacitor c=0.00603828f \
 //x=8.205 //y=0.915 //x2=8.66 //y2=1.26
cc_2503 ( N_noxref_5_c_2657_n N_noxref_7_c_3647_n ) capacitor c=0.00731987f \
 //x=8.88 //y=3.33 //x2=8.14 //y2=2.08
cc_2504 ( N_noxref_5_c_2657_n N_noxref_7_c_3648_n ) capacitor c=0.00283672f \
 //x=8.88 //y=3.33 //x2=8.14 //y2=1.915
cc_2505 ( N_noxref_5_M5_noxref_d N_noxref_7_c_3648_n ) capacitor c=0.00661782f \
 //x=8.205 //y=0.915 //x2=8.14 //y2=1.915
cc_2506 ( N_noxref_5_c_2653_n N_noxref_7_c_3650_n ) capacitor c=0.00201851f \
 //x=8.795 //y=5.155 //x2=8.14 //y2=4.7
cc_2507 ( N_noxref_5_c_2657_n N_noxref_7_c_3650_n ) capacitor c=0.013693f \
 //x=8.88 //y=3.33 //x2=8.14 //y2=4.7
cc_2508 ( N_noxref_5_c_2751_p N_noxref_7_c_3650_n ) capacitor c=0.00475601f \
 //x=8.1 //y=5.155 //x2=8.14 //y2=4.7
cc_2509 ( N_noxref_5_c_2627_n N_noxref_8_c_3904_n ) capacitor c=0.00740361f \
 //x=20.235 //y=3.33 //x2=22.685 //y2=3.33
cc_2510 ( N_noxref_5_c_2630_n N_noxref_8_c_3866_n ) capacitor c=0.0010247f \
 //x=20.35 //y=2.08 //x2=22.57 //y2=2.08
cc_2511 ( N_noxref_5_c_2626_n N_D_c_5277_n ) capacitor c=0.202839f //x=8.765 \
 //y=3.33 //x2=29.855 //y2=4.07
cc_2512 ( N_noxref_5_c_2692_n N_D_c_5277_n ) capacitor c=0.0135672f //x=3.445 \
 //y=3.33 //x2=29.855 //y2=4.07
cc_2513 ( N_noxref_5_c_2627_n N_D_c_5277_n ) capacitor c=0.0809428f //x=20.235 \
 //y=3.33 //x2=29.855 //y2=4.07
cc_2514 ( N_noxref_5_c_2695_n N_D_c_5277_n ) capacitor c=4.80262e-19 //x=8.995 \
 //y=3.33 //x2=29.855 //y2=4.07
cc_2515 ( N_noxref_5_c_2628_n N_D_c_5277_n ) capacitor c=0.0245725f //x=3.33 \
 //y=2.08 //x2=29.855 //y2=4.07
cc_2516 ( N_noxref_5_c_2647_n N_D_c_5277_n ) capacitor c=0.0157836f //x=6.425 \
 //y=5.155 //x2=29.855 //y2=4.07
cc_2517 ( N_noxref_5_c_2657_n N_D_c_5277_n ) capacitor c=0.0181789f //x=8.88 \
 //y=3.33 //x2=29.855 //y2=4.07
cc_2518 ( N_noxref_5_c_2630_n N_D_c_5277_n ) capacitor c=0.0194977f //x=20.35 \
 //y=2.08 //x2=29.855 //y2=4.07
cc_2519 ( N_noxref_5_c_2723_n N_D_c_5277_n ) capacitor c=0.00652255f //x=3.33 \
 //y=4.7 //x2=29.855 //y2=4.07
cc_2520 ( N_noxref_5_c_2628_n N_D_c_5279_n ) capacitor c=0.00168488f //x=3.33 \
 //y=2.08 //x2=1.11 //y2=2.08
cc_2521 ( N_noxref_5_c_2626_n N_CLK_c_6046_n ) capacitor c=0.00667512f \
 //x=8.765 //y=3.33 //x2=16.535 //y2=4.44
cc_2522 ( N_noxref_5_c_2653_n N_CLK_c_6046_n ) capacitor c=0.0183122f \
 //x=8.795 //y=5.155 //x2=16.535 //y2=4.44
cc_2523 ( N_noxref_5_c_2657_n N_CLK_c_6046_n ) capacitor c=0.0210274f //x=8.88 \
 //y=3.33 //x2=16.535 //y2=4.44
cc_2524 ( N_noxref_5_c_2789_p N_CLK_c_6046_n ) capacitor c=0.0311227f //x=7.22 \
 //y=5.155 //x2=16.535 //y2=4.44
cc_2525 ( N_noxref_5_c_2626_n N_CLK_c_6057_n ) capacitor c=7.37203e-19 \
 //x=8.765 //y=3.33 //x2=7.145 //y2=4.44
cc_2526 ( N_noxref_5_c_2643_n N_CLK_c_6057_n ) capacitor c=0.00330099f \
 //x=7.135 //y=5.155 //x2=7.145 //y2=4.44
cc_2527 ( N_noxref_5_c_2630_n N_CLK_c_6058_n ) capacitor c=0.0208709f \
 //x=20.35 //y=2.08 //x2=35.775 //y2=4.44
cc_2528 ( N_noxref_5_c_2669_n N_CLK_c_6058_n ) capacitor c=0.0166984f \
 //x=20.625 //y=4.79 //x2=35.775 //y2=4.44
cc_2529 ( N_noxref_5_c_2626_n N_CLK_c_6040_n ) capacitor c=0.0237264f \
 //x=8.765 //y=3.33 //x2=7.03 //y2=2.08
cc_2530 ( N_noxref_5_c_2643_n N_CLK_c_6040_n ) capacitor c=0.0143918f \
 //x=7.135 //y=5.155 //x2=7.03 //y2=2.08
cc_2531 ( N_noxref_5_c_2657_n N_CLK_c_6040_n ) capacitor c=0.00260293f \
 //x=8.88 //y=3.33 //x2=7.03 //y2=2.08
cc_2532 ( N_noxref_5_c_2627_n N_CLK_c_6041_n ) capacitor c=0.0190562f \
 //x=20.235 //y=3.33 //x2=16.65 //y2=2.08
cc_2533 ( N_noxref_5_c_2643_n N_CLK_M68_noxref_g ) capacitor c=0.016514f \
 //x=7.135 //y=5.155 //x2=7 //y2=6.02
cc_2534 ( N_noxref_5_M68_noxref_d N_CLK_M68_noxref_g ) capacitor c=0.0180032f \
 //x=7.075 //y=5.02 //x2=7 //y2=6.02
cc_2535 ( N_noxref_5_c_2649_n N_CLK_M69_noxref_g ) capacitor c=0.01736f \
 //x=8.015 //y=5.155 //x2=7.44 //y2=6.02
cc_2536 ( N_noxref_5_M68_noxref_d N_CLK_M69_noxref_g ) capacitor c=0.0180032f \
 //x=7.075 //y=5.02 //x2=7.44 //y2=6.02
cc_2537 ( N_noxref_5_c_2789_p N_CLK_c_6179_n ) capacitor c=0.00426767f \
 //x=7.22 //y=5.155 //x2=7.365 //y2=4.79
cc_2538 ( N_noxref_5_c_2643_n N_CLK_c_6131_n ) capacitor c=0.00322046f \
 //x=7.135 //y=5.155 //x2=7.03 //y2=4.7
cc_2539 ( N_noxref_5_c_2626_n N_RN_c_7021_n ) capacitor c=0.0392678f //x=8.765 \
 //y=3.33 //x2=17.645 //y2=2.22
cc_2540 ( N_noxref_5_c_2692_n N_RN_c_7021_n ) capacitor c=0.00751886f \
 //x=3.445 //y=3.33 //x2=17.645 //y2=2.22
cc_2541 ( N_noxref_5_c_2627_n N_RN_c_7021_n ) capacitor c=0.0561264f \
 //x=20.235 //y=3.33 //x2=17.645 //y2=2.22
cc_2542 ( N_noxref_5_c_2695_n N_RN_c_7021_n ) capacitor c=3.9466e-19 //x=8.995 \
 //y=3.33 //x2=17.645 //y2=2.22
cc_2543 ( N_noxref_5_c_2628_n N_RN_c_7021_n ) capacitor c=0.0225728f //x=3.33 \
 //y=2.08 //x2=17.645 //y2=2.22
cc_2544 ( N_noxref_5_c_2809_p N_RN_c_7021_n ) capacitor c=0.016327f //x=8.48 \
 //y=1.665 //x2=17.645 //y2=2.22
cc_2545 ( N_noxref_5_c_2657_n N_RN_c_7021_n ) capacitor c=0.0197307f //x=8.88 \
 //y=3.33 //x2=17.645 //y2=2.22
cc_2546 ( N_noxref_5_c_2715_n N_RN_c_7021_n ) capacitor c=3.13485e-19 \
 //x=3.695 //y=1.415 //x2=17.645 //y2=2.22
cc_2547 ( N_noxref_5_c_2720_n N_RN_c_7021_n ) capacitor c=0.00583286f //x=3.33 \
 //y=2.08 //x2=17.645 //y2=2.22
cc_2548 ( N_noxref_5_c_2628_n N_RN_c_7032_n ) capacitor c=0.00165648f //x=3.33 \
 //y=2.08 //x2=2.335 //y2=2.22
cc_2549 ( N_noxref_5_c_2720_n N_RN_c_7032_n ) capacitor c=2.3323e-19 //x=3.33 \
 //y=2.08 //x2=2.335 //y2=2.22
cc_2550 ( N_noxref_5_c_2627_n N_RN_c_7033_n ) capacitor c=0.014255f //x=20.235 \
 //y=3.33 //x2=21.345 //y2=2.22
cc_2551 ( N_noxref_5_c_2630_n N_RN_c_7033_n ) capacitor c=0.0216101f //x=20.35 \
 //y=2.08 //x2=21.345 //y2=2.22
cc_2552 ( N_noxref_5_c_2635_n N_RN_c_7033_n ) capacitor c=0.011987f //x=20.05 \
 //y=1.915 //x2=21.345 //y2=2.22
cc_2553 ( N_noxref_5_c_2627_n N_RN_c_7037_n ) capacitor c=4.86139e-19 \
 //x=20.235 //y=3.33 //x2=17.875 //y2=2.22
cc_2554 ( N_noxref_5_c_2630_n N_RN_c_7045_n ) capacitor c=0.00100368f \
 //x=20.35 //y=2.08 //x2=21.575 //y2=2.22
cc_2555 ( N_noxref_5_c_2635_n N_RN_c_7045_n ) capacitor c=2.11894e-19 \
 //x=20.05 //y=1.915 //x2=21.575 //y2=2.22
cc_2556 ( N_noxref_5_c_2692_n N_RN_c_7088_n ) capacitor c=0.00526349f \
 //x=3.445 //y=3.33 //x2=2.22 //y2=2.08
cc_2557 ( N_noxref_5_c_2628_n N_RN_c_7088_n ) capacitor c=0.0515337f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_2558 ( N_noxref_5_c_2720_n N_RN_c_7088_n ) capacitor c=0.0019893f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_2559 ( N_noxref_5_c_2723_n N_RN_c_7088_n ) capacitor c=0.00219458f //x=3.33 \
 //y=4.7 //x2=2.22 //y2=2.08
cc_2560 ( N_noxref_5_c_2627_n N_RN_c_7089_n ) capacitor c=0.0180187f \
 //x=20.235 //y=3.33 //x2=17.76 //y2=2.08
cc_2561 ( N_noxref_5_c_2630_n N_RN_c_7089_n ) capacitor c=6.89573e-19 \
 //x=20.35 //y=2.08 //x2=17.76 //y2=2.08
cc_2562 ( N_noxref_5_c_2627_n N_RN_c_7090_n ) capacitor c=0.0027353f \
 //x=20.235 //y=3.33 //x2=21.46 //y2=2.08
cc_2563 ( N_noxref_5_c_2630_n N_RN_c_7090_n ) capacitor c=0.0449054f //x=20.35 \
 //y=2.08 //x2=21.46 //y2=2.08
cc_2564 ( N_noxref_5_c_2635_n N_RN_c_7090_n ) capacitor c=0.00208635f \
 //x=20.05 //y=1.915 //x2=21.46 //y2=2.08
cc_2565 ( N_noxref_5_c_2734_p N_RN_c_7090_n ) capacitor c=0.00147352f \
 //x=20.915 //y=4.79 //x2=21.46 //y2=2.08
cc_2566 ( N_noxref_5_c_2669_n N_RN_c_7090_n ) capacitor c=0.00142741f \
 //x=20.625 //y=4.79 //x2=21.46 //y2=2.08
cc_2567 ( N_noxref_5_M64_noxref_g N_RN_M62_noxref_g ) capacitor c=0.0101598f \
 //x=3.07 //y=6.02 //x2=2.19 //y2=6.02
cc_2568 ( N_noxref_5_M64_noxref_g N_RN_M63_noxref_g ) capacitor c=0.0602553f \
 //x=3.07 //y=6.02 //x2=2.63 //y2=6.02
cc_2569 ( N_noxref_5_M65_noxref_g N_RN_M63_noxref_g ) capacitor c=0.0101598f \
 //x=3.51 //y=6.02 //x2=2.63 //y2=6.02
cc_2570 ( N_noxref_5_M84_noxref_g N_RN_M86_noxref_g ) capacitor c=0.0105869f \
 //x=20.55 //y=6.02 //x2=21.43 //y2=6.02
cc_2571 ( N_noxref_5_M85_noxref_g N_RN_M86_noxref_g ) capacitor c=0.10632f \
 //x=20.99 //y=6.02 //x2=21.43 //y2=6.02
cc_2572 ( N_noxref_5_M85_noxref_g N_RN_M87_noxref_g ) capacitor c=0.0101598f \
 //x=20.99 //y=6.02 //x2=21.87 //y2=6.02
cc_2573 ( N_noxref_5_c_2711_n N_RN_c_7204_n ) capacitor c=0.00456962f //x=3.32 \
 //y=0.915 //x2=2.31 //y2=0.91
cc_2574 ( N_noxref_5_c_2712_n N_RN_c_7205_n ) capacitor c=0.00438372f //x=3.32 \
 //y=1.26 //x2=2.31 //y2=1.22
cc_2575 ( N_noxref_5_c_2713_n N_RN_c_7206_n ) capacitor c=0.00438372f //x=3.32 \
 //y=1.57 //x2=2.31 //y2=1.45
cc_2576 ( N_noxref_5_c_2628_n N_RN_c_7207_n ) capacitor c=0.00205895f //x=3.33 \
 //y=2.08 //x2=2.31 //y2=1.915
cc_2577 ( N_noxref_5_c_2720_n N_RN_c_7207_n ) capacitor c=0.00828003f //x=3.33 \
 //y=2.08 //x2=2.31 //y2=1.915
cc_2578 ( N_noxref_5_c_2721_n N_RN_c_7207_n ) capacitor c=0.00438372f //x=3.33 \
 //y=1.915 //x2=2.31 //y2=1.915
cc_2579 ( N_noxref_5_c_2723_n N_RN_c_7161_n ) capacitor c=0.0611812f //x=3.33 \
 //y=4.7 //x2=2.555 //y2=4.79
cc_2580 ( N_noxref_5_c_2631_n N_RN_c_7211_n ) capacitor c=5.72482e-19 \
 //x=20.05 //y=0.875 //x2=21.025 //y2=0.91
cc_2581 ( N_noxref_5_c_2633_n N_RN_c_7211_n ) capacitor c=0.00149976f \
 //x=20.05 //y=1.22 //x2=21.025 //y2=0.91
cc_2582 ( N_noxref_5_c_2638_n N_RN_c_7211_n ) capacitor c=0.0160123f //x=20.58 \
 //y=0.875 //x2=21.025 //y2=0.91
cc_2583 ( N_noxref_5_c_2634_n N_RN_c_7214_n ) capacitor c=0.00111227f \
 //x=20.05 //y=1.53 //x2=21.025 //y2=1.22
cc_2584 ( N_noxref_5_c_2640_n N_RN_c_7214_n ) capacitor c=0.0124075f //x=20.58 \
 //y=1.22 //x2=21.025 //y2=1.22
cc_2585 ( N_noxref_5_c_2638_n N_RN_c_7216_n ) capacitor c=0.00103227f \
 //x=20.58 //y=0.875 //x2=21.55 //y2=0.91
cc_2586 ( N_noxref_5_c_2640_n N_RN_c_7217_n ) capacitor c=0.0010154f //x=20.58 \
 //y=1.22 //x2=21.55 //y2=1.22
cc_2587 ( N_noxref_5_c_2640_n N_RN_c_7218_n ) capacitor c=9.23422e-19 \
 //x=20.58 //y=1.22 //x2=21.55 //y2=1.45
cc_2588 ( N_noxref_5_c_2630_n N_RN_c_7219_n ) capacitor c=0.00203769f \
 //x=20.35 //y=2.08 //x2=21.55 //y2=1.915
cc_2589 ( N_noxref_5_c_2635_n N_RN_c_7219_n ) capacitor c=0.00834532f \
 //x=20.05 //y=1.915 //x2=21.55 //y2=1.915
cc_2590 ( N_noxref_5_c_2628_n N_RN_c_7162_n ) capacitor c=0.00142741f //x=3.33 \
 //y=2.08 //x2=2.22 //y2=4.7
cc_2591 ( N_noxref_5_c_2723_n N_RN_c_7162_n ) capacitor c=0.00487508f //x=3.33 \
 //y=4.7 //x2=2.22 //y2=4.7
cc_2592 ( N_noxref_5_c_2630_n N_RN_c_7223_n ) capacitor c=0.00183762f \
 //x=20.35 //y=2.08 //x2=21.46 //y2=4.7
cc_2593 ( N_noxref_5_c_2734_p N_RN_c_7223_n ) capacitor c=0.0168581f \
 //x=20.915 //y=4.79 //x2=21.46 //y2=4.7
cc_2594 ( N_noxref_5_c_2669_n N_RN_c_7223_n ) capacitor c=0.00484466f \
 //x=20.625 //y=4.79 //x2=21.46 //y2=4.7
cc_2595 ( N_noxref_5_c_2627_n N_SN_c_8129_n ) capacitor c=0.756732f //x=20.235 \
 //y=3.33 //x2=26.155 //y2=2.96
cc_2596 ( N_noxref_5_c_2630_n N_SN_c_8129_n ) capacitor c=0.0238838f //x=20.35 \
 //y=2.08 //x2=26.155 //y2=2.96
cc_2597 ( N_noxref_5_c_2627_n N_SN_c_8183_n ) capacitor c=0.0292094f \
 //x=20.235 //y=3.33 //x2=11.955 //y2=2.96
cc_2598 ( N_noxref_5_c_2627_n N_SN_c_8145_n ) capacitor c=0.0208912f \
 //x=20.235 //y=3.33 //x2=11.84 //y2=2.08
cc_2599 ( N_noxref_5_c_2657_n N_SN_c_8145_n ) capacitor c=4.63641e-19 //x=8.88 \
 //y=3.33 //x2=11.84 //y2=2.08
cc_2600 ( N_noxref_5_c_2628_n N_noxref_29_c_10596_n ) capacitor c=0.00204385f \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_2601 ( N_noxref_5_c_2711_n N_noxref_29_c_10596_n ) capacitor c=0.0194423f \
 //x=3.32 //y=0.915 //x2=3.985 //y2=0.54
cc_2602 ( N_noxref_5_c_2717_n N_noxref_29_c_10596_n ) capacitor c=0.00656458f \
 //x=3.85 //y=0.915 //x2=3.985 //y2=0.54
cc_2603 ( N_noxref_5_c_2720_n N_noxref_29_c_10596_n ) capacitor c=2.20712e-19 \
 //x=3.33 //y=2.08 //x2=3.985 //y2=0.54
cc_2604 ( N_noxref_5_c_2712_n N_noxref_29_c_10606_n ) capacitor c=0.00538829f \
 //x=3.32 //y=1.26 //x2=3.1 //y2=0.995
cc_2605 ( N_noxref_5_c_2711_n N_noxref_29_M2_noxref_s ) capacitor \
 c=0.00538829f //x=3.32 //y=0.915 //x2=2.965 //y2=0.375
cc_2606 ( N_noxref_5_c_2713_n N_noxref_29_M2_noxref_s ) capacitor \
 c=0.00538829f //x=3.32 //y=1.57 //x2=2.965 //y2=0.375
cc_2607 ( N_noxref_5_c_2717_n N_noxref_29_M2_noxref_s ) capacitor c=0.0143002f \
 //x=3.85 //y=0.915 //x2=2.965 //y2=0.375
cc_2608 ( N_noxref_5_c_2718_n N_noxref_29_M2_noxref_s ) capacitor \
 c=0.00290153f //x=3.85 //y=1.26 //x2=2.965 //y2=0.375
cc_2609 ( N_noxref_5_M5_noxref_d N_noxref_30_M3_noxref_s ) capacitor \
 c=0.00309936f //x=8.205 //y=0.915 //x2=5.265 //y2=0.375
cc_2610 ( N_noxref_5_c_2629_n N_noxref_31_c_10697_n ) capacitor c=0.00457167f \
 //x=8.795 //y=1.665 //x2=8.795 //y2=0.54
cc_2611 ( N_noxref_5_M5_noxref_d N_noxref_31_c_10697_n ) capacitor \
 c=0.0115903f //x=8.205 //y=0.915 //x2=8.795 //y2=0.54
cc_2612 ( N_noxref_5_c_2809_p N_noxref_31_c_10707_n ) capacitor c=0.0200405f \
 //x=8.48 //y=1.665 //x2=7.91 //y2=0.995
cc_2613 ( N_noxref_5_M5_noxref_d N_noxref_31_M4_noxref_d ) capacitor \
 c=5.27807e-19 //x=8.205 //y=0.915 //x2=6.67 //y2=0.91
cc_2614 ( N_noxref_5_c_2629_n N_noxref_31_M5_noxref_s ) capacitor c=0.0196084f \
 //x=8.795 //y=1.665 //x2=7.775 //y2=0.375
cc_2615 ( N_noxref_5_M5_noxref_d N_noxref_31_M5_noxref_s ) capacitor \
 c=0.0426368f //x=8.205 //y=0.915 //x2=7.775 //y2=0.375
cc_2616 ( N_noxref_5_c_2629_n N_noxref_32_c_10759_n ) capacitor c=3.84569e-19 \
 //x=8.795 //y=1.665 //x2=10.21 //y2=1.505
cc_2617 ( N_noxref_5_M5_noxref_d N_noxref_32_M6_noxref_s ) capacitor \
 c=2.55333e-19 //x=8.205 //y=0.915 //x2=10.075 //y2=0.375
cc_2618 ( N_noxref_5_c_2635_n N_noxref_36_c_10962_n ) capacitor c=0.0034165f \
 //x=20.05 //y=1.915 //x2=19.83 //y2=1.505
cc_2619 ( N_noxref_5_c_2630_n N_noxref_36_c_10947_n ) capacitor c=0.0115578f \
 //x=20.35 //y=2.08 //x2=20.715 //y2=1.59
cc_2620 ( N_noxref_5_c_2634_n N_noxref_36_c_10947_n ) capacitor c=0.00697148f \
 //x=20.05 //y=1.53 //x2=20.715 //y2=1.59
cc_2621 ( N_noxref_5_c_2635_n N_noxref_36_c_10947_n ) capacitor c=0.0204849f \
 //x=20.05 //y=1.915 //x2=20.715 //y2=1.59
cc_2622 ( N_noxref_5_c_2637_n N_noxref_36_c_10947_n ) capacitor c=0.00610316f \
 //x=20.425 //y=1.375 //x2=20.715 //y2=1.59
cc_2623 ( N_noxref_5_c_2640_n N_noxref_36_c_10947_n ) capacitor c=0.00698822f \
 //x=20.58 //y=1.22 //x2=20.715 //y2=1.59
cc_2624 ( N_noxref_5_c_2631_n N_noxref_36_M12_noxref_s ) capacitor \
 c=0.0327271f //x=20.05 //y=0.875 //x2=19.695 //y2=0.375
cc_2625 ( N_noxref_5_c_2634_n N_noxref_36_M12_noxref_s ) capacitor \
 c=7.99997e-19 //x=20.05 //y=1.53 //x2=19.695 //y2=0.375
cc_2626 ( N_noxref_5_c_2635_n N_noxref_36_M12_noxref_s ) capacitor \
 c=0.00122123f //x=20.05 //y=1.915 //x2=19.695 //y2=0.375
cc_2627 ( N_noxref_5_c_2638_n N_noxref_36_M12_noxref_s ) capacitor \
 c=0.0121427f //x=20.58 //y=0.875 //x2=19.695 //y2=0.375
cc_2628 ( N_noxref_6_c_2896_n N_noxref_7_c_3623_n ) capacitor c=0.0187698f \
 //x=23.31 //y=2.59 //x2=27.265 //y2=3.7
cc_2629 ( N_noxref_6_c_2897_n N_noxref_7_c_3623_n ) capacitor c=0.0197889f \
 //x=25.16 //y=2.08 //x2=27.265 //y2=3.7
cc_2630 ( N_noxref_6_c_3020_n N_noxref_7_c_3544_n ) capacitor c=3.10026e-19 \
 //x=20.855 //y=5.155 //x2=18.415 //y2=5.155
cc_2631 ( N_noxref_6_c_2934_n N_noxref_7_c_3530_n ) capacitor c=0.012757f \
 //x=75.025 //y=4.81 //x2=27.38 //y2=2.08
cc_2632 ( N_noxref_6_c_2897_n N_noxref_7_c_3530_n ) capacitor c=0.00111863f \
 //x=25.16 //y=2.08 //x2=27.38 //y2=2.08
cc_2633 ( N_noxref_6_c_2934_n N_noxref_7_M94_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=27.12 //y2=6.02
cc_2634 ( N_noxref_6_c_2934_n N_noxref_7_M95_noxref_g ) capacitor \
 c=0.00288422f //x=75.025 //y=4.81 //x2=27.56 //y2=6.02
cc_2635 ( N_noxref_6_c_2934_n N_noxref_7_c_3660_n ) capacitor c=0.00205991f \
 //x=75.025 //y=4.81 //x2=27.38 //y2=4.7
cc_2636 ( N_noxref_6_c_2893_n N_noxref_8_c_3906_n ) capacitor c=0.0119023f \
 //x=25.045 //y=2.59 //x2=28.005 //y2=3.33
cc_2637 ( N_noxref_6_c_2894_n N_noxref_8_c_3906_n ) capacitor c=8.87672e-19 \
 //x=23.425 //y=2.59 //x2=28.005 //y2=3.33
cc_2638 ( N_noxref_6_c_2896_n N_noxref_8_c_3906_n ) capacitor c=0.018769f \
 //x=23.31 //y=2.59 //x2=28.005 //y2=3.33
cc_2639 ( N_noxref_6_c_2897_n N_noxref_8_c_3906_n ) capacitor c=0.0197803f \
 //x=25.16 //y=2.08 //x2=28.005 //y2=3.33
cc_2640 ( N_noxref_6_c_2896_n N_noxref_8_c_3904_n ) capacitor c=0.00131333f \
 //x=23.31 //y=2.59 //x2=22.685 //y2=3.33
cc_2641 ( N_noxref_6_c_2894_n N_noxref_8_c_3866_n ) capacitor c=0.00720056f \
 //x=23.425 //y=2.59 //x2=22.57 //y2=2.08
cc_2642 ( N_noxref_6_c_2990_n N_noxref_8_c_3866_n ) capacitor c=0.0045659f \
 //x=23.425 //y=4.81 //x2=22.57 //y2=2.08
cc_2643 ( N_noxref_6_c_2896_n N_noxref_8_c_3866_n ) capacitor c=0.0747906f \
 //x=23.31 //y=2.59 //x2=22.57 //y2=2.08
cc_2644 ( N_noxref_6_c_2897_n N_noxref_8_c_3866_n ) capacitor c=5.32619e-19 \
 //x=25.16 //y=2.08 //x2=22.57 //y2=2.08
cc_2645 ( N_noxref_6_c_3093_p N_noxref_8_c_3866_n ) capacitor c=0.0166016f \
 //x=22.53 //y=5.155 //x2=22.57 //y2=2.08
cc_2646 ( N_noxref_6_M91_noxref_g N_noxref_8_c_3870_n ) capacitor c=0.0157304f \
 //x=25.8 //y=6.02 //x2=26.375 //y2=5.155
cc_2647 ( N_noxref_6_c_2934_n N_noxref_8_c_3874_n ) capacitor c=0.112727f \
 //x=75.025 //y=4.81 //x2=25.665 //y2=5.155
cc_2648 ( N_noxref_6_c_3026_n N_noxref_8_c_3874_n ) capacitor c=3.10026e-19 \
 //x=23.225 //y=5.155 //x2=25.665 //y2=5.155
cc_2649 ( N_noxref_6_M90_noxref_g N_noxref_8_c_3874_n ) capacitor c=0.0213876f \
 //x=25.36 //y=6.02 //x2=25.665 //y2=5.155
cc_2650 ( N_noxref_6_c_3098_p N_noxref_8_c_3874_n ) capacitor c=0.00393496f \
 //x=25.725 //y=4.79 //x2=25.665 //y2=5.155
cc_2651 ( N_noxref_6_c_2934_n N_noxref_8_c_3884_n ) capacitor c=0.0187537f \
 //x=75.025 //y=4.81 //x2=28.12 //y2=3.33
cc_2652 ( N_noxref_6_c_3022_n N_noxref_8_M88_noxref_g ) capacitor c=0.01736f \
 //x=22.445 //y=5.155 //x2=22.31 //y2=6.02
cc_2653 ( N_noxref_6_M88_noxref_d N_noxref_8_M88_noxref_g ) capacitor \
 c=0.0180032f //x=22.385 //y=5.02 //x2=22.31 //y2=6.02
cc_2654 ( N_noxref_6_c_2990_n N_noxref_8_M89_noxref_g ) capacitor \
 c=5.47828e-19 //x=23.425 //y=4.81 //x2=22.75 //y2=6.02
cc_2655 ( N_noxref_6_c_3026_n N_noxref_8_M89_noxref_g ) capacitor c=0.0194981f \
 //x=23.225 //y=5.155 //x2=22.75 //y2=6.02
cc_2656 ( N_noxref_6_M88_noxref_d N_noxref_8_M89_noxref_g ) capacitor \
 c=0.0194246f //x=22.385 //y=5.02 //x2=22.75 //y2=6.02
cc_2657 ( N_noxref_6_M14_noxref_d N_noxref_8_c_3927_n ) capacitor \
 c=0.00217566f //x=22.635 //y=0.915 //x2=22.56 //y2=0.915
cc_2658 ( N_noxref_6_M14_noxref_d N_noxref_8_c_3928_n ) capacitor c=0.0034598f \
 //x=22.635 //y=0.915 //x2=22.56 //y2=1.26
cc_2659 ( N_noxref_6_M14_noxref_d N_noxref_8_c_3929_n ) capacitor \
 c=0.00546784f //x=22.635 //y=0.915 //x2=22.56 //y2=1.57
cc_2660 ( N_noxref_6_M14_noxref_d N_noxref_8_c_3930_n ) capacitor \
 c=0.00241102f //x=22.635 //y=0.915 //x2=22.935 //y2=0.76
cc_2661 ( N_noxref_6_c_2895_n N_noxref_8_c_3931_n ) capacitor c=0.00371277f \
 //x=23.225 //y=1.665 //x2=22.935 //y2=1.415
cc_2662 ( N_noxref_6_M14_noxref_d N_noxref_8_c_3931_n ) capacitor c=0.0138621f \
 //x=22.635 //y=0.915 //x2=22.935 //y2=1.415
cc_2663 ( N_noxref_6_M14_noxref_d N_noxref_8_c_3933_n ) capacitor \
 c=0.00219619f //x=22.635 //y=0.915 //x2=23.09 //y2=0.915
cc_2664 ( N_noxref_6_c_2895_n N_noxref_8_c_3934_n ) capacitor c=0.00457401f \
 //x=23.225 //y=1.665 //x2=23.09 //y2=1.26
cc_2665 ( N_noxref_6_M14_noxref_d N_noxref_8_c_3934_n ) capacitor \
 c=0.00603828f //x=22.635 //y=0.915 //x2=23.09 //y2=1.26
cc_2666 ( N_noxref_6_c_2896_n N_noxref_8_c_3936_n ) capacitor c=0.00709342f \
 //x=23.31 //y=2.59 //x2=22.57 //y2=2.08
cc_2667 ( N_noxref_6_c_2896_n N_noxref_8_c_3937_n ) capacitor c=0.00283672f \
 //x=23.31 //y=2.59 //x2=22.57 //y2=1.915
cc_2668 ( N_noxref_6_M14_noxref_d N_noxref_8_c_3937_n ) capacitor \
 c=0.00661782f //x=22.635 //y=0.915 //x2=22.57 //y2=1.915
cc_2669 ( N_noxref_6_c_2990_n N_noxref_8_c_3939_n ) capacitor c=0.00660462f \
 //x=23.425 //y=4.81 //x2=22.57 //y2=4.7
cc_2670 ( N_noxref_6_c_3026_n N_noxref_8_c_3939_n ) capacitor c=0.00201851f \
 //x=23.225 //y=5.155 //x2=22.57 //y2=4.7
cc_2671 ( N_noxref_6_c_2896_n N_noxref_8_c_3939_n ) capacitor c=0.0121399f \
 //x=23.31 //y=2.59 //x2=22.57 //y2=4.7
cc_2672 ( N_noxref_6_c_3093_p N_noxref_8_c_3939_n ) capacitor c=0.00475601f \
 //x=22.53 //y=5.155 //x2=22.57 //y2=4.7
cc_2673 ( N_noxref_6_M91_noxref_g N_noxref_8_M90_noxref_d ) capacitor \
 c=0.0180032f //x=25.8 //y=6.02 //x2=25.435 //y2=5.02
cc_2674 ( N_noxref_6_c_2934_n N_noxref_9_c_4075_n ) capacitor c=0.112727f \
 //x=75.025 //y=4.81 //x2=30.475 //y2=5.155
cc_2675 ( N_noxref_6_c_2934_n N_noxref_9_c_4047_n ) capacitor c=0.0187537f \
 //x=75.025 //y=4.81 //x2=32.93 //y2=2.59
cc_2676 ( N_noxref_6_c_2934_n N_noxref_9_c_4048_n ) capacitor c=0.0139535f \
 //x=75.025 //y=4.81 //x2=34.78 //y2=2.08
cc_2677 ( N_noxref_6_c_2934_n N_noxref_9_c_4049_n ) capacitor c=0.0139535f \
 //x=75.025 //y=4.81 //x2=39.59 //y2=2.08
cc_2678 ( N_noxref_6_c_2934_n N_noxref_9_M102_noxref_g ) capacitor \
 c=0.00558442f //x=75.025 //y=4.81 //x2=34.98 //y2=6.02
cc_2679 ( N_noxref_6_c_2934_n N_noxref_9_M103_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=35.42 //y2=6.02
cc_2680 ( N_noxref_6_c_2934_n N_noxref_9_M108_noxref_g ) capacitor \
 c=0.00558442f //x=75.025 //y=4.81 //x2=39.79 //y2=6.02
cc_2681 ( N_noxref_6_c_2934_n N_noxref_9_M109_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=40.23 //y2=6.02
cc_2682 ( N_noxref_6_c_2934_n N_noxref_9_c_4127_n ) capacitor c=0.00458471f \
 //x=75.025 //y=4.81 //x2=35.345 //y2=4.79
cc_2683 ( N_noxref_6_c_2934_n N_noxref_9_c_4100_n ) capacitor c=0.00184926f \
 //x=75.025 //y=4.81 //x2=35.055 //y2=4.79
cc_2684 ( N_noxref_6_c_2934_n N_noxref_9_c_4129_n ) capacitor c=0.00458471f \
 //x=75.025 //y=4.81 //x2=40.155 //y2=4.79
cc_2685 ( N_noxref_6_c_2934_n N_noxref_9_c_4102_n ) capacitor c=0.00184926f \
 //x=75.025 //y=4.81 //x2=39.865 //y2=4.79
cc_2686 ( N_noxref_6_c_2934_n N_noxref_10_c_4315_n ) capacitor c=0.112727f \
 //x=75.025 //y=4.81 //x2=40.095 //y2=5.155
cc_2687 ( N_noxref_6_c_2934_n N_noxref_10_c_4298_n ) capacitor c=0.0187537f \
 //x=75.025 //y=4.81 //x2=42.55 //y2=2.59
cc_2688 ( N_noxref_6_c_2934_n N_noxref_10_c_4299_n ) capacitor c=0.0139535f \
 //x=75.025 //y=4.81 //x2=44.4 //y2=2.08
cc_2689 ( N_noxref_6_c_2934_n N_noxref_10_M114_noxref_g ) capacitor \
 c=0.00558442f //x=75.025 //y=4.81 //x2=44.6 //y2=6.02
cc_2690 ( N_noxref_6_c_2934_n N_noxref_10_M115_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=45.04 //y2=6.02
cc_2691 ( N_noxref_6_c_2934_n N_noxref_10_c_4355_n ) capacitor c=0.00458471f \
 //x=75.025 //y=4.81 //x2=44.965 //y2=4.79
cc_2692 ( N_noxref_6_c_2934_n N_noxref_10_c_4333_n ) capacitor c=0.00184926f \
 //x=75.025 //y=4.81 //x2=44.675 //y2=4.79
cc_2693 ( N_noxref_6_c_2934_n N_noxref_11_c_4464_n ) capacitor c=0.012757f \
 //x=75.025 //y=4.81 //x2=32.19 //y2=2.08
cc_2694 ( N_noxref_6_c_2934_n N_noxref_11_c_4483_n ) capacitor c=0.112727f \
 //x=75.025 //y=4.81 //x2=35.285 //y2=5.155
cc_2695 ( N_noxref_6_c_2934_n N_noxref_11_c_4493_n ) capacitor c=0.0187537f \
 //x=75.025 //y=4.81 //x2=37.74 //y2=3.33
cc_2696 ( N_noxref_6_c_2934_n N_noxref_11_c_4466_n ) capacitor c=0.0139535f \
 //x=75.025 //y=4.81 //x2=49.21 //y2=2.08
cc_2697 ( N_noxref_6_c_2934_n N_noxref_11_M100_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=31.93 //y2=6.02
cc_2698 ( N_noxref_6_c_2934_n N_noxref_11_M101_noxref_g ) capacitor \
 c=0.00288422f //x=75.025 //y=4.81 //x2=32.37 //y2=6.02
cc_2699 ( N_noxref_6_c_2934_n N_noxref_11_M120_noxref_g ) capacitor \
 c=0.00558442f //x=75.025 //y=4.81 //x2=49.41 //y2=6.02
cc_2700 ( N_noxref_6_c_2934_n N_noxref_11_M121_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=49.85 //y2=6.02
cc_2701 ( N_noxref_6_c_2934_n N_noxref_11_c_4530_n ) capacitor c=0.00458471f \
 //x=75.025 //y=4.81 //x2=49.775 //y2=4.79
cc_2702 ( N_noxref_6_c_2934_n N_noxref_11_c_4505_n ) capacitor c=0.00184926f \
 //x=75.025 //y=4.81 //x2=49.485 //y2=4.79
cc_2703 ( N_noxref_6_c_2934_n N_noxref_11_c_4532_n ) capacitor c=0.00205991f \
 //x=75.025 //y=4.81 //x2=32.19 //y2=4.7
cc_2704 ( N_noxref_6_c_2934_n N_noxref_12_c_4745_n ) capacitor c=0.012757f \
 //x=75.025 //y=4.81 //x2=37 //y2=2.08
cc_2705 ( N_noxref_6_c_2934_n N_noxref_12_c_4746_n ) capacitor c=0.012757f \
 //x=75.025 //y=4.81 //x2=41.81 //y2=2.08
cc_2706 ( N_noxref_6_c_2934_n N_noxref_12_c_4756_n ) capacitor c=0.112727f \
 //x=75.025 //y=4.81 //x2=44.905 //y2=5.155
cc_2707 ( N_noxref_6_c_2934_n N_noxref_12_c_4766_n ) capacitor c=0.0187537f \
 //x=75.025 //y=4.81 //x2=47.36 //y2=3.7
cc_2708 ( N_noxref_6_c_2934_n N_noxref_12_c_4748_n ) capacitor c=0.012757f \
 //x=75.025 //y=4.81 //x2=56.24 //y2=2.08
cc_2709 ( N_noxref_6_c_2934_n N_noxref_12_M106_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=36.74 //y2=6.02
cc_2710 ( N_noxref_6_c_2934_n N_noxref_12_M107_noxref_g ) capacitor \
 c=0.00288422f //x=75.025 //y=4.81 //x2=37.18 //y2=6.02
cc_2711 ( N_noxref_6_c_2934_n N_noxref_12_M112_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=41.55 //y2=6.02
cc_2712 ( N_noxref_6_c_2934_n N_noxref_12_M113_noxref_g ) capacitor \
 c=0.00288422f //x=75.025 //y=4.81 //x2=41.99 //y2=6.02
cc_2713 ( N_noxref_6_c_2934_n N_noxref_12_M130_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=55.98 //y2=6.02
cc_2714 ( N_noxref_6_c_2934_n N_noxref_12_M131_noxref_g ) capacitor \
 c=0.00288422f //x=75.025 //y=4.81 //x2=56.42 //y2=6.02
cc_2715 ( N_noxref_6_c_2934_n N_noxref_12_c_4806_n ) capacitor c=0.00205991f \
 //x=75.025 //y=4.81 //x2=37 //y2=4.7
cc_2716 ( N_noxref_6_c_2934_n N_noxref_12_c_4807_n ) capacitor c=0.00205991f \
 //x=75.025 //y=4.81 //x2=41.81 //y2=4.7
cc_2717 ( N_noxref_6_c_2934_n N_noxref_12_c_4808_n ) capacitor c=0.00205991f \
 //x=75.025 //y=4.81 //x2=56.24 //y2=4.7
cc_2718 ( N_noxref_6_c_2934_n N_noxref_13_c_5101_n ) capacitor c=0.012757f \
 //x=75.025 //y=4.81 //x2=51.43 //y2=2.08
cc_2719 ( N_noxref_6_c_2934_n N_noxref_13_c_5110_n ) capacitor c=0.112727f \
 //x=75.025 //y=4.81 //x2=54.525 //y2=5.155
cc_2720 ( N_noxref_6_c_2934_n N_noxref_13_c_5103_n ) capacitor c=0.0187537f \
 //x=75.025 //y=4.81 //x2=56.98 //y2=2.59
cc_2721 ( N_noxref_6_c_2934_n N_noxref_13_M124_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=51.17 //y2=6.02
cc_2722 ( N_noxref_6_c_2934_n N_noxref_13_M125_noxref_g ) capacitor \
 c=0.00288422f //x=75.025 //y=4.81 //x2=51.61 //y2=6.02
cc_2723 ( N_noxref_6_c_2934_n N_noxref_13_c_5145_n ) capacitor c=0.00205991f \
 //x=75.025 //y=4.81 //x2=51.43 //y2=4.7
cc_2724 ( N_noxref_6_c_2934_n N_D_c_5277_n ) capacitor c=0.0387198f //x=75.025 \
 //y=4.81 //x2=29.855 //y2=4.07
cc_2725 ( N_noxref_6_c_2990_n N_D_c_5277_n ) capacitor c=8.80731e-19 \
 //x=23.425 //y=4.81 //x2=29.855 //y2=4.07
cc_2726 ( N_noxref_6_c_2896_n N_D_c_5277_n ) capacitor c=0.0181982f //x=23.31 \
 //y=2.59 //x2=29.855 //y2=4.07
cc_2727 ( N_noxref_6_c_2897_n N_D_c_5277_n ) capacitor c=0.019517f //x=25.16 \
 //y=2.08 //x2=29.855 //y2=4.07
cc_2728 ( N_noxref_6_c_2934_n N_D_c_5328_n ) capacitor c=0.167266f //x=75.025 \
 //y=4.81 //x2=58.715 //y2=4.07
cc_2729 ( N_noxref_6_c_2934_n N_D_c_5280_n ) capacitor c=0.0139535f //x=75.025 \
 //y=4.81 //x2=29.97 //y2=2.08
cc_2730 ( N_noxref_6_c_2934_n N_D_c_5281_n ) capacitor c=0.0139535f //x=75.025 \
 //y=4.81 //x2=58.83 //y2=2.08
cc_2731 ( N_noxref_6_c_2934_n N_D_M96_noxref_g ) capacitor c=0.00558442f \
 //x=75.025 //y=4.81 //x2=30.17 //y2=6.02
cc_2732 ( N_noxref_6_c_2934_n N_D_M97_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=30.61 //y2=6.02
cc_2733 ( N_noxref_6_c_2934_n N_D_M132_noxref_g ) capacitor c=0.00558442f \
 //x=75.025 //y=4.81 //x2=59.03 //y2=6.02
cc_2734 ( N_noxref_6_c_2934_n N_D_M133_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=59.47 //y2=6.02
cc_2735 ( N_noxref_6_c_2934_n N_D_c_5400_n ) capacitor c=0.00458471f \
 //x=75.025 //y=4.81 //x2=30.535 //y2=4.79
cc_2736 ( N_noxref_6_c_2934_n N_D_c_5358_n ) capacitor c=0.00184926f \
 //x=75.025 //y=4.81 //x2=30.245 //y2=4.79
cc_2737 ( N_noxref_6_c_2934_n N_D_c_5402_n ) capacitor c=0.00458471f \
 //x=75.025 //y=4.81 //x2=59.395 //y2=4.79
cc_2738 ( N_noxref_6_c_2934_n N_D_c_5360_n ) capacitor c=0.00184926f \
 //x=75.025 //y=4.81 //x2=59.105 //y2=4.79
cc_2739 ( N_noxref_6_c_2934_n N_noxref_15_c_5652_n ) capacitor c=0.112727f \
 //x=75.025 //y=4.81 //x2=59.335 //y2=5.155
cc_2740 ( N_noxref_6_c_2934_n N_noxref_15_c_5624_n ) capacitor c=0.0187537f \
 //x=75.025 //y=4.81 //x2=61.79 //y2=2.59
cc_2741 ( N_noxref_6_c_2934_n N_noxref_15_c_5625_n ) capacitor c=0.0139535f \
 //x=75.025 //y=4.81 //x2=63.64 //y2=2.08
cc_2742 ( N_noxref_6_c_2934_n N_noxref_15_c_5626_n ) capacitor c=0.0139535f \
 //x=75.025 //y=4.81 //x2=68.45 //y2=2.08
cc_2743 ( N_noxref_6_c_2934_n N_noxref_15_M138_noxref_g ) capacitor \
 c=0.00558442f //x=75.025 //y=4.81 //x2=63.84 //y2=6.02
cc_2744 ( N_noxref_6_c_2934_n N_noxref_15_M139_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=64.28 //y2=6.02
cc_2745 ( N_noxref_6_c_2934_n N_noxref_15_M144_noxref_g ) capacitor \
 c=0.00558442f //x=75.025 //y=4.81 //x2=68.65 //y2=6.02
cc_2746 ( N_noxref_6_c_2934_n N_noxref_15_M145_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=69.09 //y2=6.02
cc_2747 ( N_noxref_6_c_2934_n N_noxref_15_c_5704_n ) capacitor c=0.00458471f \
 //x=75.025 //y=4.81 //x2=64.205 //y2=4.79
cc_2748 ( N_noxref_6_c_2934_n N_noxref_15_c_5677_n ) capacitor c=0.00184926f \
 //x=75.025 //y=4.81 //x2=63.915 //y2=4.79
cc_2749 ( N_noxref_6_c_2934_n N_noxref_15_c_5706_n ) capacitor c=0.00458471f \
 //x=75.025 //y=4.81 //x2=69.015 //y2=4.79
cc_2750 ( N_noxref_6_c_2934_n N_noxref_15_c_5679_n ) capacitor c=0.00184926f \
 //x=75.025 //y=4.81 //x2=68.725 //y2=4.79
cc_2751 ( N_noxref_6_c_2934_n N_noxref_16_c_5892_n ) capacitor c=0.112727f \
 //x=75.025 //y=4.81 //x2=68.955 //y2=5.155
cc_2752 ( N_noxref_6_c_2934_n N_noxref_16_c_5875_n ) capacitor c=0.0187537f \
 //x=75.025 //y=4.81 //x2=71.41 //y2=2.59
cc_2753 ( N_noxref_6_c_2934_n N_noxref_16_c_5876_n ) capacitor c=0.0139535f \
 //x=75.025 //y=4.81 //x2=73.26 //y2=2.08
cc_2754 ( N_noxref_6_c_2934_n N_noxref_16_M150_noxref_g ) capacitor \
 c=0.00558442f //x=75.025 //y=4.81 //x2=73.46 //y2=6.02
cc_2755 ( N_noxref_6_c_2934_n N_noxref_16_M151_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=73.9 //y2=6.02
cc_2756 ( N_noxref_6_c_2934_n N_noxref_16_c_5932_n ) capacitor c=0.00458471f \
 //x=75.025 //y=4.81 //x2=73.825 //y2=4.79
cc_2757 ( N_noxref_6_c_2934_n N_noxref_16_c_5910_n ) capacitor c=0.00184926f \
 //x=75.025 //y=4.81 //x2=73.535 //y2=4.79
cc_2758 ( N_noxref_6_c_2934_n N_CLK_c_6058_n ) capacitor c=1.07152f //x=75.025 \
 //y=4.81 //x2=35.775 //y2=4.44
cc_2759 ( N_noxref_6_c_2990_n N_CLK_c_6058_n ) capacitor c=0.0292847f \
 //x=23.425 //y=4.81 //x2=35.775 //y2=4.44
cc_2760 ( N_noxref_6_c_3016_n N_CLK_c_6058_n ) capacitor c=0.032141f \
 //x=21.565 //y=5.155 //x2=35.775 //y2=4.44
cc_2761 ( N_noxref_6_c_3020_n N_CLK_c_6058_n ) capacitor c=0.0230136f \
 //x=20.855 //y=5.155 //x2=35.775 //y2=4.44
cc_2762 ( N_noxref_6_c_3026_n N_CLK_c_6058_n ) capacitor c=0.0165623f \
 //x=23.225 //y=5.155 //x2=35.775 //y2=4.44
cc_2763 ( N_noxref_6_c_2896_n N_CLK_c_6058_n ) capacitor c=0.0184447f \
 //x=23.31 //y=2.59 //x2=35.775 //y2=4.44
cc_2764 ( N_noxref_6_c_2897_n N_CLK_c_6058_n ) capacitor c=0.018786f //x=25.16 \
 //y=2.08 //x2=35.775 //y2=4.44
cc_2765 ( N_noxref_6_c_3052_n N_CLK_c_6058_n ) capacitor c=0.0112124f \
 //x=25.435 //y=4.79 //x2=35.775 //y2=4.44
cc_2766 ( N_noxref_6_c_2934_n N_CLK_c_6068_n ) capacitor c=0.813498f \
 //x=75.025 //y=4.81 //x2=45.395 //y2=4.44
cc_2767 ( N_noxref_6_c_2934_n N_CLK_c_6190_n ) capacitor c=0.0274297f \
 //x=75.025 //y=4.81 //x2=36.005 //y2=4.44
cc_2768 ( N_noxref_6_c_2934_n N_CLK_c_6070_n ) capacitor c=1.64653f //x=75.025 \
 //y=4.81 //x2=64.635 //y2=4.44
cc_2769 ( N_noxref_6_c_2934_n N_CLK_c_6192_n ) capacitor c=0.0274297f \
 //x=75.025 //y=4.81 //x2=45.625 //y2=4.44
cc_2770 ( N_noxref_6_c_2934_n N_CLK_c_6074_n ) capacitor c=0.843459f \
 //x=75.025 //y=4.81 //x2=74.255 //y2=4.44
cc_2771 ( N_noxref_6_c_3219_p N_CLK_c_6074_n ) capacitor c=0.00143832f \
 //x=75.11 //y=4.725 //x2=74.255 //y2=4.44
cc_2772 ( N_noxref_6_c_3220_p N_CLK_c_6074_n ) capacitor c=0.015699f \
 //x=75.195 //y=4.44 //x2=74.255 //y2=4.44
cc_2773 ( N_noxref_6_c_2934_n N_CLK_c_6196_n ) capacitor c=0.0274297f \
 //x=75.025 //y=4.81 //x2=64.865 //y2=4.44
cc_2774 ( N_noxref_6_c_2934_n N_CLK_c_6042_n ) capacitor c=0.015102f \
 //x=75.025 //y=4.81 //x2=35.89 //y2=2.08
cc_2775 ( N_noxref_6_c_2934_n N_CLK_c_6043_n ) capacitor c=0.015102f \
 //x=75.025 //y=4.81 //x2=45.51 //y2=2.08
cc_2776 ( N_noxref_6_c_2934_n N_CLK_c_6044_n ) capacitor c=0.015102f \
 //x=75.025 //y=4.81 //x2=64.75 //y2=2.08
cc_2777 ( N_noxref_6_c_2934_n N_CLK_c_6045_n ) capacitor c=0.015097f \
 //x=75.025 //y=4.81 //x2=74.37 //y2=2.08
cc_2778 ( N_noxref_6_c_3219_p N_CLK_c_6045_n ) capacitor c=0.00452835f \
 //x=75.11 //y=4.725 //x2=74.37 //y2=2.08
cc_2779 ( N_noxref_6_c_3220_p N_CLK_c_6045_n ) capacitor c=0.00267376f \
 //x=75.195 //y=4.44 //x2=74.37 //y2=2.08
cc_2780 ( N_noxref_6_c_2934_n N_CLK_M104_noxref_g ) capacitor c=0.00246676f \
 //x=75.025 //y=4.81 //x2=35.86 //y2=6.02
cc_2781 ( N_noxref_6_c_2934_n N_CLK_M105_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=36.3 //y2=6.02
cc_2782 ( N_noxref_6_c_2934_n N_CLK_M116_noxref_g ) capacitor c=0.00246676f \
 //x=75.025 //y=4.81 //x2=45.48 //y2=6.02
cc_2783 ( N_noxref_6_c_2934_n N_CLK_M117_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=45.92 //y2=6.02
cc_2784 ( N_noxref_6_c_2934_n N_CLK_M140_noxref_g ) capacitor c=0.00246676f \
 //x=75.025 //y=4.81 //x2=64.72 //y2=6.02
cc_2785 ( N_noxref_6_c_2934_n N_CLK_M141_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=65.16 //y2=6.02
cc_2786 ( N_noxref_6_c_2934_n N_CLK_M152_noxref_g ) capacitor c=0.00246676f \
 //x=75.025 //y=4.81 //x2=74.34 //y2=6.02
cc_2787 ( N_noxref_6_c_2934_n N_CLK_M153_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=74.78 //y2=6.02
cc_2788 ( N_noxref_6_c_2934_n N_CLK_c_6211_n ) capacitor c=0.00356032f \
 //x=75.025 //y=4.81 //x2=36.225 //y2=4.79
cc_2789 ( N_noxref_6_c_2934_n N_CLK_c_6212_n ) capacitor c=0.00356032f \
 //x=75.025 //y=4.81 //x2=45.845 //y2=4.79
cc_2790 ( N_noxref_6_c_2934_n N_CLK_c_6213_n ) capacitor c=0.00356032f \
 //x=75.025 //y=4.81 //x2=65.085 //y2=4.79
cc_2791 ( N_noxref_6_c_2934_n N_CLK_c_6214_n ) capacitor c=0.00458005f \
 //x=75.025 //y=4.81 //x2=74.705 //y2=4.79
cc_2792 ( N_noxref_6_c_2934_n N_CLK_c_6215_n ) capacitor c=9.51445e-19 \
 //x=75.025 //y=4.81 //x2=35.89 //y2=4.7
cc_2793 ( N_noxref_6_c_2934_n N_CLK_c_6216_n ) capacitor c=9.51445e-19 \
 //x=75.025 //y=4.81 //x2=45.51 //y2=4.7
cc_2794 ( N_noxref_6_c_2934_n N_CLK_c_6217_n ) capacitor c=9.51445e-19 \
 //x=75.025 //y=4.81 //x2=64.75 //y2=4.7
cc_2795 ( N_noxref_6_c_2934_n N_CLK_c_6218_n ) capacitor c=9.51445e-19 \
 //x=75.025 //y=4.81 //x2=74.37 //y2=4.7
cc_2796 ( N_noxref_6_c_3219_p N_CLK_c_6218_n ) capacitor c=0.00252294f \
 //x=75.11 //y=4.725 //x2=74.37 //y2=4.7
cc_2797 ( N_noxref_6_c_2934_n N_noxref_18_c_6747_n ) capacitor c=0.012757f \
 //x=75.025 //y=4.81 //x2=61.05 //y2=2.08
cc_2798 ( N_noxref_6_c_2934_n N_noxref_18_c_6766_n ) capacitor c=0.112846f \
 //x=75.025 //y=4.81 //x2=64.145 //y2=5.155
cc_2799 ( N_noxref_6_c_2934_n N_noxref_18_c_6776_n ) capacitor c=0.0187537f \
 //x=75.025 //y=4.81 //x2=66.6 //y2=3.33
cc_2800 ( N_noxref_6_c_2993_n N_noxref_18_c_6749_n ) capacitor c=0.0208709f \
 //x=87.205 //y=4.44 //x2=78.07 //y2=2.08
cc_2801 ( N_noxref_6_c_2934_n N_noxref_18_M136_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=60.79 //y2=6.02
cc_2802 ( N_noxref_6_c_2934_n N_noxref_18_M137_noxref_g ) capacitor \
 c=0.00288422f //x=75.025 //y=4.81 //x2=61.23 //y2=6.02
cc_2803 ( N_noxref_6_c_2993_n N_noxref_18_c_6788_n ) capacitor c=0.0166984f \
 //x=87.205 //y=4.44 //x2=78.345 //y2=4.79
cc_2804 ( N_noxref_6_c_2934_n N_noxref_18_c_6812_n ) capacitor c=0.00205991f \
 //x=75.025 //y=4.81 //x2=61.05 //y2=4.7
cc_2805 ( N_noxref_6_c_2893_n N_RN_c_7038_n ) capacitor c=0.172592f //x=25.045 \
 //y=2.59 //x2=30.965 //y2=2.22
cc_2806 ( N_noxref_6_c_2894_n N_RN_c_7038_n ) capacitor c=0.0291301f \
 //x=23.425 //y=2.59 //x2=30.965 //y2=2.22
cc_2807 ( N_noxref_6_c_3255_p N_RN_c_7038_n ) capacitor c=0.016327f //x=22.91 \
 //y=1.665 //x2=30.965 //y2=2.22
cc_2808 ( N_noxref_6_c_2896_n N_RN_c_7038_n ) capacitor c=0.0215653f //x=23.31 \
 //y=2.59 //x2=30.965 //y2=2.22
cc_2809 ( N_noxref_6_c_2897_n N_RN_c_7038_n ) capacitor c=0.021104f //x=25.16 \
 //y=2.08 //x2=30.965 //y2=2.22
cc_2810 ( N_noxref_6_c_2907_n N_RN_c_7038_n ) capacitor c=0.011987f //x=24.86 \
 //y=1.915 //x2=30.965 //y2=2.22
cc_2811 ( N_noxref_6_c_3016_n N_RN_c_7090_n ) capacitor c=0.0144268f \
 //x=21.565 //y=5.155 //x2=21.46 //y2=2.08
cc_2812 ( N_noxref_6_c_2896_n N_RN_c_7090_n ) capacitor c=0.00226806f \
 //x=23.31 //y=2.59 //x2=21.46 //y2=2.08
cc_2813 ( N_noxref_6_c_2934_n N_RN_c_7091_n ) capacitor c=0.0132674f \
 //x=75.025 //y=4.81 //x2=31.08 //y2=2.08
cc_2814 ( N_noxref_6_c_2934_n N_RN_c_7092_n ) capacitor c=0.012757f //x=75.025 \
 //y=4.81 //x2=46.62 //y2=2.08
cc_2815 ( N_noxref_6_c_2934_n N_RN_c_7093_n ) capacitor c=0.0132674f \
 //x=75.025 //y=4.81 //x2=50.32 //y2=2.08
cc_2816 ( N_noxref_6_c_2934_n N_RN_c_7094_n ) capacitor c=0.0132674f \
 //x=75.025 //y=4.81 //x2=59.94 //y2=2.08
cc_2817 ( N_noxref_6_c_3219_p N_RN_c_7095_n ) capacitor c=0.0133429f //x=75.11 \
 //y=4.725 //x2=75.48 //y2=2.08
cc_2818 ( N_noxref_6_c_2993_n N_RN_c_7095_n ) capacitor c=0.0191507f \
 //x=87.205 //y=4.44 //x2=75.48 //y2=2.08
cc_2819 ( N_noxref_6_c_2993_n N_RN_c_7096_n ) capacitor c=0.0210462f \
 //x=87.205 //y=4.44 //x2=79.18 //y2=2.08
cc_2820 ( N_noxref_6_c_3016_n N_RN_M86_noxref_g ) capacitor c=0.0165266f \
 //x=21.565 //y=5.155 //x2=21.43 //y2=6.02
cc_2821 ( N_noxref_6_M86_noxref_d N_RN_M86_noxref_g ) capacitor c=0.0180032f \
 //x=21.505 //y=5.02 //x2=21.43 //y2=6.02
cc_2822 ( N_noxref_6_c_3022_n N_RN_M87_noxref_g ) capacitor c=0.01736f \
 //x=22.445 //y=5.155 //x2=21.87 //y2=6.02
cc_2823 ( N_noxref_6_M86_noxref_d N_RN_M87_noxref_g ) capacitor c=0.0180032f \
 //x=21.505 //y=5.02 //x2=21.87 //y2=6.02
cc_2824 ( N_noxref_6_c_2934_n N_RN_M98_noxref_g ) capacitor c=0.00246676f \
 //x=75.025 //y=4.81 //x2=31.05 //y2=6.02
cc_2825 ( N_noxref_6_c_2934_n N_RN_M99_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=31.49 //y2=6.02
cc_2826 ( N_noxref_6_c_2934_n N_RN_M118_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=46.36 //y2=6.02
cc_2827 ( N_noxref_6_c_2934_n N_RN_M119_noxref_g ) capacitor c=0.00288422f \
 //x=75.025 //y=4.81 //x2=46.8 //y2=6.02
cc_2828 ( N_noxref_6_c_2934_n N_RN_M122_noxref_g ) capacitor c=0.00246676f \
 //x=75.025 //y=4.81 //x2=50.29 //y2=6.02
cc_2829 ( N_noxref_6_c_2934_n N_RN_M123_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=50.73 //y2=6.02
cc_2830 ( N_noxref_6_c_2934_n N_RN_M134_noxref_g ) capacitor c=0.00246676f \
 //x=75.025 //y=4.81 //x2=59.91 //y2=6.02
cc_2831 ( N_noxref_6_c_2934_n N_RN_M135_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=60.35 //y2=6.02
cc_2832 ( N_noxref_6_c_2934_n N_RN_M154_noxref_g ) capacitor c=0.00178866f \
 //x=75.025 //y=4.81 //x2=75.22 //y2=6.02
cc_2833 ( N_noxref_6_c_2934_n N_RN_M155_noxref_g ) capacitor c=3.26891e-19 \
 //x=75.025 //y=4.81 //x2=75.66 //y2=6.02
cc_2834 ( N_noxref_6_c_3282_p N_RN_c_7255_n ) capacitor c=0.00426767f \
 //x=21.65 //y=5.155 //x2=21.795 //y2=4.79
cc_2835 ( N_noxref_6_c_2934_n N_RN_c_7256_n ) capacitor c=0.00356032f \
 //x=75.025 //y=4.81 //x2=31.415 //y2=4.79
cc_2836 ( N_noxref_6_c_2934_n N_RN_c_7257_n ) capacitor c=0.00356032f \
 //x=75.025 //y=4.81 //x2=50.655 //y2=4.79
cc_2837 ( N_noxref_6_c_2934_n N_RN_c_7258_n ) capacitor c=0.00356032f \
 //x=75.025 //y=4.81 //x2=60.275 //y2=4.79
cc_2838 ( N_noxref_6_c_2993_n N_RN_c_7259_n ) capacitor c=0.0085986f \
 //x=87.205 //y=4.44 //x2=79.515 //y2=4.79
cc_2839 ( N_noxref_6_c_3016_n N_RN_c_7223_n ) capacitor c=0.00322054f \
 //x=21.565 //y=5.155 //x2=21.46 //y2=4.7
cc_2840 ( N_noxref_6_c_2934_n N_RN_c_7261_n ) capacitor c=5.37461e-19 \
 //x=75.025 //y=4.81 //x2=31.08 //y2=4.7
cc_2841 ( N_noxref_6_c_2934_n N_RN_c_7262_n ) capacitor c=0.00205991f \
 //x=75.025 //y=4.81 //x2=46.62 //y2=4.7
cc_2842 ( N_noxref_6_c_2934_n N_RN_c_7263_n ) capacitor c=5.37461e-19 \
 //x=75.025 //y=4.81 //x2=50.32 //y2=4.7
cc_2843 ( N_noxref_6_c_2934_n N_RN_c_7264_n ) capacitor c=5.37461e-19 \
 //x=75.025 //y=4.81 //x2=59.94 //y2=4.7
cc_2844 ( N_noxref_6_c_2934_n N_RN_c_7265_n ) capacitor c=0.00244717f \
 //x=75.025 //y=4.81 //x2=75.48 //y2=4.7
cc_2845 ( N_noxref_6_c_3219_p N_RN_c_7265_n ) capacitor c=0.00370337f \
 //x=75.11 //y=4.725 //x2=75.48 //y2=4.7
cc_2846 ( N_noxref_6_c_2993_n N_RN_c_7265_n ) capacitor c=0.00989126f \
 //x=87.205 //y=4.44 //x2=75.48 //y2=4.7
cc_2847 ( N_noxref_6_c_2993_n N_RN_c_7268_n ) capacitor c=0.00293313f \
 //x=87.205 //y=4.44 //x2=79.18 //y2=4.7
cc_2848 ( N_noxref_6_c_2893_n N_SN_c_8129_n ) capacitor c=0.172781f //x=25.045 \
 //y=2.59 //x2=26.155 //y2=2.96
cc_2849 ( N_noxref_6_c_2894_n N_SN_c_8129_n ) capacitor c=0.0293832f \
 //x=23.425 //y=2.59 //x2=26.155 //y2=2.96
cc_2850 ( N_noxref_6_c_2896_n N_SN_c_8129_n ) capacitor c=0.0206007f //x=23.31 \
 //y=2.59 //x2=26.155 //y2=2.96
cc_2851 ( N_noxref_6_c_2897_n N_SN_c_8129_n ) capacitor c=0.0216195f //x=25.16 \
 //y=2.08 //x2=26.155 //y2=2.96
cc_2852 ( N_noxref_6_c_2897_n N_SN_c_8226_n ) capacitor c=0.00128547f \
 //x=25.16 //y=2.08 //x2=26.385 //y2=2.96
cc_2853 ( N_noxref_6_c_2893_n N_SN_c_8146_n ) capacitor c=0.00520283f \
 //x=25.045 //y=2.59 //x2=26.27 //y2=2.08
cc_2854 ( N_noxref_6_c_2934_n N_SN_c_8146_n ) capacitor c=0.0132674f \
 //x=75.025 //y=4.81 //x2=26.27 //y2=2.08
cc_2855 ( N_noxref_6_c_2896_n N_SN_c_8146_n ) capacitor c=3.11441e-19 \
 //x=23.31 //y=2.59 //x2=26.27 //y2=2.08
cc_2856 ( N_noxref_6_c_2897_n N_SN_c_8146_n ) capacitor c=0.0402779f //x=25.16 \
 //y=2.08 //x2=26.27 //y2=2.08
cc_2857 ( N_noxref_6_c_2907_n N_SN_c_8146_n ) capacitor c=0.00210802f \
 //x=24.86 //y=1.915 //x2=26.27 //y2=2.08
cc_2858 ( N_noxref_6_c_3098_p N_SN_c_8146_n ) capacitor c=0.00120758f \
 //x=25.725 //y=4.79 //x2=26.27 //y2=2.08
cc_2859 ( N_noxref_6_c_3052_n N_SN_c_8146_n ) capacitor c=0.00142741f \
 //x=25.435 //y=4.79 //x2=26.27 //y2=2.08
cc_2860 ( N_noxref_6_c_2934_n N_SN_c_8147_n ) capacitor c=0.0132674f \
 //x=75.025 //y=4.81 //x2=40.7 //y2=2.08
cc_2861 ( N_noxref_6_c_2934_n N_SN_c_8148_n ) capacitor c=0.0132674f \
 //x=75.025 //y=4.81 //x2=55.13 //y2=2.08
cc_2862 ( N_noxref_6_c_2934_n N_SN_c_8149_n ) capacitor c=0.0132674f \
 //x=75.025 //y=4.81 //x2=69.56 //y2=2.08
cc_2863 ( N_noxref_6_c_2993_n N_SN_c_8150_n ) capacitor c=0.0210462f \
 //x=87.205 //y=4.44 //x2=83.99 //y2=2.08
cc_2864 ( N_noxref_6_c_2934_n N_SN_M92_noxref_g ) capacitor c=0.00246676f \
 //x=75.025 //y=4.81 //x2=26.24 //y2=6.02
cc_2865 ( N_noxref_6_M90_noxref_g N_SN_M92_noxref_g ) capacitor c=0.0105174f \
 //x=25.36 //y=6.02 //x2=26.24 //y2=6.02
cc_2866 ( N_noxref_6_M91_noxref_g N_SN_M92_noxref_g ) capacitor c=0.10624f \
 //x=25.8 //y=6.02 //x2=26.24 //y2=6.02
cc_2867 ( N_noxref_6_c_2934_n N_SN_M93_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=26.68 //y2=6.02
cc_2868 ( N_noxref_6_M91_noxref_g N_SN_M93_noxref_g ) capacitor c=0.0100903f \
 //x=25.8 //y=6.02 //x2=26.68 //y2=6.02
cc_2869 ( N_noxref_6_c_2934_n N_SN_M110_noxref_g ) capacitor c=0.00246676f \
 //x=75.025 //y=4.81 //x2=40.67 //y2=6.02
cc_2870 ( N_noxref_6_c_2934_n N_SN_M111_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=41.11 //y2=6.02
cc_2871 ( N_noxref_6_c_2934_n N_SN_M128_noxref_g ) capacitor c=0.00246676f \
 //x=75.025 //y=4.81 //x2=55.1 //y2=6.02
cc_2872 ( N_noxref_6_c_2934_n N_SN_M129_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=55.54 //y2=6.02
cc_2873 ( N_noxref_6_c_2934_n N_SN_M146_noxref_g ) capacitor c=0.00246676f \
 //x=75.025 //y=4.81 //x2=69.53 //y2=6.02
cc_2874 ( N_noxref_6_c_2934_n N_SN_M147_noxref_g ) capacitor c=0.00267973f \
 //x=75.025 //y=4.81 //x2=69.97 //y2=6.02
cc_2875 ( N_noxref_6_c_2903_n N_SN_c_8249_n ) capacitor c=5.72482e-19 \
 //x=24.86 //y=0.875 //x2=25.835 //y2=0.91
cc_2876 ( N_noxref_6_c_2905_n N_SN_c_8249_n ) capacitor c=0.00149976f \
 //x=24.86 //y=1.22 //x2=25.835 //y2=0.91
cc_2877 ( N_noxref_6_c_2910_n N_SN_c_8249_n ) capacitor c=0.0160123f //x=25.39 \
 //y=0.875 //x2=25.835 //y2=0.91
cc_2878 ( N_noxref_6_c_2906_n N_SN_c_8252_n ) capacitor c=0.00111227f \
 //x=24.86 //y=1.53 //x2=25.835 //y2=1.22
cc_2879 ( N_noxref_6_c_2912_n N_SN_c_8252_n ) capacitor c=0.0124075f //x=25.39 \
 //y=1.22 //x2=25.835 //y2=1.22
cc_2880 ( N_noxref_6_c_2910_n N_SN_c_8254_n ) capacitor c=0.00103227f \
 //x=25.39 //y=0.875 //x2=26.36 //y2=0.91
cc_2881 ( N_noxref_6_c_2912_n N_SN_c_8255_n ) capacitor c=0.0010154f //x=25.39 \
 //y=1.22 //x2=26.36 //y2=1.22
cc_2882 ( N_noxref_6_c_2912_n N_SN_c_8256_n ) capacitor c=9.23422e-19 \
 //x=25.39 //y=1.22 //x2=26.36 //y2=1.45
cc_2883 ( N_noxref_6_c_2897_n N_SN_c_8257_n ) capacitor c=0.00203769f \
 //x=25.16 //y=2.08 //x2=26.36 //y2=1.915
cc_2884 ( N_noxref_6_c_2907_n N_SN_c_8257_n ) capacitor c=0.00834532f \
 //x=24.86 //y=1.915 //x2=26.36 //y2=1.915
cc_2885 ( N_noxref_6_c_2934_n N_SN_c_8259_n ) capacitor c=0.00356032f \
 //x=75.025 //y=4.81 //x2=26.605 //y2=4.79
cc_2886 ( N_noxref_6_c_2934_n N_SN_c_8260_n ) capacitor c=0.00356032f \
 //x=75.025 //y=4.81 //x2=41.035 //y2=4.79
cc_2887 ( N_noxref_6_c_2934_n N_SN_c_8261_n ) capacitor c=0.00356032f \
 //x=75.025 //y=4.81 //x2=55.465 //y2=4.79
cc_2888 ( N_noxref_6_c_2934_n N_SN_c_8262_n ) capacitor c=0.00356032f \
 //x=75.025 //y=4.81 //x2=69.895 //y2=4.79
cc_2889 ( N_noxref_6_c_2993_n N_SN_c_8263_n ) capacitor c=0.0085986f \
 //x=87.205 //y=4.44 //x2=84.325 //y2=4.79
cc_2890 ( N_noxref_6_c_2934_n N_SN_c_8264_n ) capacitor c=5.37461e-19 \
 //x=75.025 //y=4.81 //x2=26.27 //y2=4.7
cc_2891 ( N_noxref_6_c_2897_n N_SN_c_8264_n ) capacitor c=0.0017365f //x=25.16 \
 //y=2.08 //x2=26.27 //y2=4.7
cc_2892 ( N_noxref_6_c_3098_p N_SN_c_8264_n ) capacitor c=0.0170104f \
 //x=25.725 //y=4.79 //x2=26.27 //y2=4.7
cc_2893 ( N_noxref_6_c_3052_n N_SN_c_8264_n ) capacitor c=0.00484466f \
 //x=25.435 //y=4.79 //x2=26.27 //y2=4.7
cc_2894 ( N_noxref_6_c_2934_n N_SN_c_8268_n ) capacitor c=5.37461e-19 \
 //x=75.025 //y=4.81 //x2=40.7 //y2=4.7
cc_2895 ( N_noxref_6_c_2934_n N_SN_c_8269_n ) capacitor c=5.37461e-19 \
 //x=75.025 //y=4.81 //x2=55.13 //y2=4.7
cc_2896 ( N_noxref_6_c_2934_n N_SN_c_8270_n ) capacitor c=5.37461e-19 \
 //x=75.025 //y=4.81 //x2=69.56 //y2=4.7
cc_2897 ( N_noxref_6_c_2993_n N_SN_c_8271_n ) capacitor c=0.00293313f \
 //x=87.205 //y=4.44 //x2=83.99 //y2=4.7
cc_2898 ( N_noxref_6_c_2934_n N_noxref_21_c_8878_n ) capacitor c=0.00279672f \
 //x=75.025 //y=4.81 //x2=76.105 //y2=3.7
cc_2899 ( N_noxref_6_c_3220_p N_noxref_21_c_8878_n ) capacitor c=0.00925922f \
 //x=75.195 //y=4.44 //x2=76.105 //y2=3.7
cc_2900 ( N_noxref_6_c_2993_n N_noxref_21_c_8880_n ) capacitor c=0.0644712f \
 //x=87.205 //y=4.44 //x2=84.985 //y2=3.7
cc_2901 ( N_noxref_6_c_2993_n N_noxref_21_c_8881_n ) capacitor c=4.78746e-19 \
 //x=87.205 //y=4.44 //x2=76.335 //y2=3.7
cc_2902 ( N_noxref_6_c_2934_n N_noxref_21_c_8828_n ) capacitor c=0.012757f \
 //x=75.025 //y=4.81 //x2=65.86 //y2=2.08
cc_2903 ( N_noxref_6_c_2934_n N_noxref_21_c_8829_n ) capacitor c=0.012757f \
 //x=75.025 //y=4.81 //x2=70.67 //y2=2.08
cc_2904 ( N_noxref_6_c_2934_n N_noxref_21_c_8839_n ) capacitor c=0.0728972f \
 //x=75.025 //y=4.81 //x2=73.765 //y2=5.155
cc_2905 ( N_noxref_6_c_2993_n N_noxref_21_c_8841_n ) capacitor c=0.0072467f \
 //x=87.205 //y=4.44 //x2=75.355 //y2=5.155
cc_2906 ( N_noxref_6_c_2993_n N_noxref_21_c_8845_n ) capacitor c=0.0183122f \
 //x=87.205 //y=4.44 //x2=76.135 //y2=5.155
cc_2907 ( N_noxref_6_c_2934_n N_noxref_21_c_8849_n ) capacitor c=0.00105091f \
 //x=75.025 //y=4.81 //x2=76.22 //y2=3.7
cc_2908 ( N_noxref_6_c_2993_n N_noxref_21_c_8849_n ) capacitor c=0.0210274f \
 //x=87.205 //y=4.44 //x2=76.22 //y2=3.7
cc_2909 ( N_noxref_6_c_2993_n N_noxref_21_c_8831_n ) capacitor c=0.0200057f \
 //x=87.205 //y=4.44 //x2=85.1 //y2=2.08
cc_2910 ( N_noxref_6_c_2898_n N_noxref_21_c_8831_n ) capacitor c=0.00118902f \
 //x=87.32 //y=2.08 //x2=85.1 //y2=2.08
cc_2911 ( N_noxref_6_c_2934_n N_noxref_21_M142_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=65.6 //y2=6.02
cc_2912 ( N_noxref_6_c_2934_n N_noxref_21_M143_noxref_g ) capacitor \
 c=0.00288422f //x=75.025 //y=4.81 //x2=66.04 //y2=6.02
cc_2913 ( N_noxref_6_c_2934_n N_noxref_21_M148_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=70.41 //y2=6.02
cc_2914 ( N_noxref_6_c_2934_n N_noxref_21_M149_noxref_g ) capacitor \
 c=0.00288422f //x=75.025 //y=4.81 //x2=70.85 //y2=6.02
cc_2915 ( N_noxref_6_c_2934_n N_noxref_21_c_8895_n ) capacitor c=0.00205991f \
 //x=75.025 //y=4.81 //x2=65.86 //y2=4.7
cc_2916 ( N_noxref_6_c_2934_n N_noxref_21_c_8896_n ) capacitor c=0.00205991f \
 //x=75.025 //y=4.81 //x2=70.67 //y2=4.7
cc_2917 ( N_noxref_6_c_2993_n N_noxref_21_c_8897_n ) capacitor c=0.0111881f \
 //x=87.205 //y=4.44 //x2=85.1 //y2=4.7
cc_2918 ( N_noxref_6_c_2993_n N_noxref_22_c_9171_n ) capacitor c=0.00343796f \
 //x=87.205 //y=4.44 //x2=85.725 //y2=2.59
cc_2919 ( N_noxref_6_c_2993_n N_noxref_22_c_9175_n ) capacitor c=0.0200057f \
 //x=87.205 //y=4.44 //x2=80.29 //y2=2.08
cc_2920 ( N_noxref_6_c_2993_n N_noxref_22_c_9180_n ) capacitor c=0.032141f \
 //x=87.205 //y=4.44 //x2=84.095 //y2=5.155
cc_2921 ( N_noxref_6_c_2993_n N_noxref_22_c_9184_n ) capacitor c=0.0230136f \
 //x=87.205 //y=4.44 //x2=83.385 //y2=5.155
cc_2922 ( N_noxref_6_c_2993_n N_noxref_22_c_9190_n ) capacitor c=0.0183122f \
 //x=87.205 //y=4.44 //x2=85.755 //y2=5.155
cc_2923 ( N_noxref_6_c_2993_n N_noxref_22_c_9177_n ) capacitor c=0.0210274f \
 //x=87.205 //y=4.44 //x2=85.84 //y2=2.59
cc_2924 ( N_noxref_6_c_2898_n N_noxref_22_c_9177_n ) capacitor c=0.0209332f \
 //x=87.32 //y=2.08 //x2=85.84 //y2=2.59
cc_2925 ( N_noxref_6_c_2993_n N_noxref_22_c_9222_n ) capacitor c=0.0111881f \
 //x=87.205 //y=4.44 //x2=80.29 //y2=4.7
cc_2926 ( N_noxref_6_c_3007_n N_noxref_23_c_9342_n ) capacitor c=0.0856654f \
 //x=90.905 //y=4.44 //x2=90.575 //y2=5.21
cc_2927 ( N_noxref_6_M172_noxref_g N_noxref_23_c_9342_n ) capacitor \
 c=0.00503498f //x=90.91 //y=6.025 //x2=90.575 //y2=5.21
cc_2928 ( N_noxref_6_c_3007_n N_noxref_23_c_9348_n ) capacitor c=0.0130311f \
 //x=90.905 //y=4.44 //x2=88.805 //y2=5.21
cc_2929 ( N_noxref_6_c_3007_n N_noxref_23_c_9353_n ) capacitor c=0.00145992f \
 //x=90.905 //y=4.44 //x2=88.605 //y2=5.21
cc_2930 ( N_noxref_6_M169_noxref_g N_noxref_23_c_9353_n ) capacitor \
 c=0.0169795f //x=88.03 //y=6.025 //x2=88.605 //y2=5.21
cc_2931 ( N_noxref_6_c_3007_n N_noxref_23_c_9357_n ) capacitor c=0.0197096f \
 //x=90.905 //y=4.44 //x2=87.895 //y2=5.21
cc_2932 ( N_noxref_6_M168_noxref_g N_noxref_23_c_9357_n ) capacitor \
 c=0.0172236f //x=87.59 //y=6.025 //x2=87.895 //y2=5.21
cc_2933 ( N_noxref_6_c_3381_p N_noxref_23_c_9357_n ) capacitor c=0.00405363f \
 //x=87.955 //y=4.795 //x2=87.895 //y2=5.21
cc_2934 ( N_noxref_6_c_3007_n N_noxref_23_c_9359_n ) capacitor c=0.00467548f \
 //x=90.905 //y=4.44 //x2=88.69 //y2=5.295
cc_2935 ( N_noxref_6_c_3007_n N_noxref_23_c_9362_n ) capacitor c=0.00439121f \
 //x=90.905 //y=4.44 //x2=90.69 //y2=5.21
cc_2936 ( N_noxref_6_M172_noxref_g N_noxref_23_c_9362_n ) capacitor \
 c=0.0481665f //x=90.91 //y=6.025 //x2=90.69 //y2=5.21
cc_2937 ( N_noxref_6_c_3007_n N_noxref_23_c_9388_n ) capacitor c=0.00249667f \
 //x=90.905 //y=4.44 //x2=91.485 //y2=6.91
cc_2938 ( N_noxref_6_c_2901_n N_noxref_23_c_9388_n ) capacitor c=8.81369e-19 \
 //x=91.02 //y=2.08 //x2=91.485 //y2=6.91
cc_2939 ( N_noxref_6_M172_noxref_g N_noxref_23_c_9388_n ) capacitor \
 c=0.0163949f //x=90.91 //y=6.025 //x2=91.485 //y2=6.91
cc_2940 ( N_noxref_6_M173_noxref_g N_noxref_23_c_9388_n ) capacitor \
 c=0.0150104f //x=91.35 //y=6.025 //x2=91.485 //y2=6.91
cc_2941 ( N_noxref_6_M169_noxref_g N_noxref_23_M168_noxref_d ) capacitor \
 c=0.0169879f //x=88.03 //y=6.025 //x2=87.665 //y2=5.025
cc_2942 ( N_noxref_6_M173_noxref_g N_noxref_23_M173_noxref_d ) capacitor \
 c=0.0130327f //x=91.35 //y=6.025 //x2=91.425 //y2=5.025
cc_2943 ( N_noxref_6_c_2993_n N_noxref_24_c_9440_n ) capacitor c=0.00223593f \
 //x=87.205 //y=4.44 //x2=92.355 //y2=2.22
cc_2944 ( N_noxref_6_c_3007_n N_noxref_24_c_9440_n ) capacitor c=0.0138862f \
 //x=90.905 //y=4.44 //x2=92.355 //y2=2.22
cc_2945 ( N_noxref_6_c_3012_n N_noxref_24_c_9440_n ) capacitor c=3.84749e-19 \
 //x=87.435 //y=4.44 //x2=92.355 //y2=2.22
cc_2946 ( N_noxref_6_c_2898_n N_noxref_24_c_9440_n ) capacitor c=0.0238027f \
 //x=87.32 //y=2.08 //x2=92.355 //y2=2.22
cc_2947 ( N_noxref_6_c_2901_n N_noxref_24_c_9440_n ) capacitor c=0.0236386f \
 //x=91.02 //y=2.08 //x2=92.355 //y2=2.22
cc_2948 ( N_noxref_6_c_2926_n N_noxref_24_c_9440_n ) capacitor c=0.00813982f \
 //x=90.825 //y=1.915 //x2=92.355 //y2=2.22
cc_2949 ( N_noxref_6_c_2932_n N_noxref_24_c_9440_n ) capacitor c=0.00825063f \
 //x=87.32 //y=2.08 //x2=92.355 //y2=2.22
cc_2950 ( N_noxref_6_c_2901_n N_noxref_24_c_9449_n ) capacitor c=0.00466111f \
 //x=91.02 //y=2.08 //x2=92.5 //y2=2.08
cc_2951 ( N_noxref_6_c_2993_n N_noxref_24_c_9478_n ) capacitor c=0.032141f \
 //x=87.205 //y=4.44 //x2=79.285 //y2=5.155
cc_2952 ( N_noxref_6_c_2993_n N_noxref_24_c_9482_n ) capacitor c=0.0230136f \
 //x=87.205 //y=4.44 //x2=78.575 //y2=5.155
cc_2953 ( N_noxref_6_c_2993_n N_noxref_24_c_9488_n ) capacitor c=0.0183122f \
 //x=87.205 //y=4.44 //x2=80.945 //y2=5.155
cc_2954 ( N_noxref_6_c_2993_n N_noxref_24_c_9451_n ) capacitor c=0.0210274f \
 //x=87.205 //y=4.44 //x2=81.03 //y2=2.22
cc_2955 ( N_noxref_6_c_2993_n N_noxref_24_c_9452_n ) capacitor c=0.0208709f \
 //x=87.205 //y=4.44 //x2=82.88 //y2=2.08
cc_2956 ( N_noxref_6_c_3007_n N_noxref_24_c_9453_n ) capacitor c=0.00408423f \
 //x=90.905 //y=4.44 //x2=92.5 //y2=2.08
cc_2957 ( N_noxref_6_c_2901_n N_noxref_24_c_9453_n ) capacitor c=0.0355675f \
 //x=91.02 //y=2.08 //x2=92.5 //y2=2.08
cc_2958 ( N_noxref_6_c_2926_n N_noxref_24_c_9453_n ) capacitor c=2.35599e-19 \
 //x=90.825 //y=1.915 //x2=92.5 //y2=2.08
cc_2959 ( N_noxref_6_c_3056_n N_noxref_24_c_9453_n ) capacitor c=2.35599e-19 \
 //x=91.02 //y=4.705 //x2=92.5 //y2=2.08
cc_2960 ( N_noxref_6_c_2901_n N_noxref_24_c_9455_n ) capacitor c=4.31424e-19 \
 //x=91.02 //y=2.08 //x2=93.98 //y2=2.08
cc_2961 ( N_noxref_6_M172_noxref_g N_noxref_24_M174_noxref_g ) capacitor \
 c=0.009459f //x=90.91 //y=6.025 //x2=91.79 //y2=6.025
cc_2962 ( N_noxref_6_M173_noxref_g N_noxref_24_M174_noxref_g ) capacitor \
 c=0.0626756f //x=91.35 //y=6.025 //x2=91.79 //y2=6.025
cc_2963 ( N_noxref_6_M173_noxref_g N_noxref_24_M175_noxref_g ) capacitor \
 c=0.00899012f //x=91.35 //y=6.025 //x2=92.23 //y2=6.025
cc_2964 ( N_noxref_6_c_2993_n N_noxref_24_c_9509_n ) capacitor c=0.0166984f \
 //x=87.205 //y=4.44 //x2=83.155 //y2=4.79
cc_2965 ( N_noxref_6_c_2923_n N_noxref_24_c_9550_n ) capacitor c=4.86506e-19 \
 //x=90.825 //y=0.865 //x2=91.795 //y2=0.905
cc_2966 ( N_noxref_6_c_2925_n N_noxref_24_c_9550_n ) capacitor c=0.00101233f \
 //x=90.825 //y=1.21 //x2=91.795 //y2=0.905
cc_2967 ( N_noxref_6_c_2929_n N_noxref_24_c_9550_n ) capacitor c=0.0168844f \
 //x=91.355 //y=0.865 //x2=91.795 //y2=0.905
cc_2968 ( N_noxref_6_c_3416_p N_noxref_24_c_9553_n ) capacitor c=7.88071e-19 \
 //x=90.825 //y=1.52 //x2=91.795 //y2=1.25
cc_2969 ( N_noxref_6_c_2931_n N_noxref_24_c_9553_n ) capacitor c=0.0168218f \
 //x=91.355 //y=1.21 //x2=91.795 //y2=1.25
cc_2970 ( N_noxref_6_c_2901_n N_noxref_24_c_9555_n ) capacitor c=9.39431e-19 \
 //x=91.02 //y=2.08 //x2=91.865 //y2=4.795
cc_2971 ( N_noxref_6_c_3056_n N_noxref_24_c_9555_n ) capacitor c=0.0634092f \
 //x=91.02 //y=4.705 //x2=91.865 //y2=4.795
cc_2972 ( N_noxref_6_c_2901_n N_noxref_24_c_9511_n ) capacitor c=2.35599e-19 \
 //x=91.02 //y=2.08 //x2=92.23 //y2=4.87
cc_2973 ( N_noxref_6_c_3056_n N_noxref_24_c_9511_n ) capacitor c=5.35364e-19 \
 //x=91.02 //y=4.705 //x2=92.23 //y2=4.87
cc_2974 ( N_noxref_6_c_2929_n N_noxref_24_c_9559_n ) capacitor c=0.00124821f \
 //x=91.355 //y=0.865 //x2=92.325 //y2=0.905
cc_2975 ( N_noxref_6_c_2931_n N_noxref_24_c_9560_n ) capacitor c=8.19575e-19 \
 //x=91.355 //y=1.21 //x2=92.325 //y2=1.25
cc_2976 ( N_noxref_6_c_2931_n N_noxref_24_c_9561_n ) capacitor c=3.60397e-19 \
 //x=91.355 //y=1.21 //x2=92.325 //y2=1.56
cc_2977 ( N_noxref_6_c_2901_n N_noxref_24_c_9466_n ) capacitor c=2.35599e-19 \
 //x=91.02 //y=2.08 //x2=92.325 //y2=1.915
cc_2978 ( N_noxref_6_c_2926_n N_noxref_24_c_9466_n ) capacitor c=4.61972e-19 \
 //x=90.825 //y=1.915 //x2=92.325 //y2=1.915
cc_2979 ( N_noxref_6_M173_noxref_g N_noxref_25_c_9838_n ) capacitor \
 c=0.0179287f //x=91.35 //y=6.025 //x2=91.925 //y2=5.21
cc_2980 ( N_noxref_6_c_3007_n N_noxref_25_c_9829_n ) capacitor c=0.0021588f \
 //x=90.905 //y=4.44 //x2=91.215 //y2=5.21
cc_2981 ( N_noxref_6_c_2901_n N_noxref_25_c_9829_n ) capacitor c=0.0056513f \
 //x=91.02 //y=2.08 //x2=91.215 //y2=5.21
cc_2982 ( N_noxref_6_M172_noxref_g N_noxref_25_c_9829_n ) capacitor \
 c=0.0132827f //x=90.91 //y=6.025 //x2=91.215 //y2=5.21
cc_2983 ( N_noxref_6_c_3056_n N_noxref_25_c_9829_n ) capacitor c=0.00554802f \
 //x=91.02 //y=4.705 //x2=91.215 //y2=5.21
cc_2984 ( N_noxref_6_M173_noxref_g N_noxref_25_M172_noxref_d ) capacitor \
 c=0.0130327f //x=91.35 //y=6.025 //x2=90.985 //y2=5.025
cc_2985 ( N_noxref_6_c_2934_n N_noxref_26_c_9933_n ) capacitor c=0.0208109f \
 //x=75.025 //y=4.81 //x2=65.035 //y2=3.7
cc_2986 ( N_noxref_6_c_3220_p N_noxref_26_c_9912_n ) capacitor c=1.06014f \
 //x=75.195 //y=4.44 //x2=88.315 //y2=4.07
cc_2987 ( N_noxref_6_c_3007_n N_noxref_26_c_9912_n ) capacitor c=0.0763193f \
 //x=90.905 //y=4.44 //x2=88.315 //y2=4.07
cc_2988 ( N_noxref_6_c_3012_n N_noxref_26_c_9912_n ) capacitor c=0.0265335f \
 //x=87.435 //y=4.44 //x2=88.315 //y2=4.07
cc_2989 ( N_noxref_6_c_2898_n N_noxref_26_c_9912_n ) capacitor c=0.0263238f \
 //x=87.32 //y=2.08 //x2=88.315 //y2=4.07
cc_2990 ( N_noxref_6_c_2934_n N_noxref_26_c_10001_n ) capacitor c=0.0774037f \
 //x=75.025 //y=4.81 //x2=65.205 //y2=4.07
cc_2991 ( N_noxref_6_c_3007_n N_noxref_26_c_9913_n ) capacitor c=0.23799f \
 //x=90.905 //y=4.44 //x2=94.975 //y2=4.07
cc_2992 ( N_noxref_6_c_2901_n N_noxref_26_c_9913_n ) capacitor c=0.0274281f \
 //x=91.02 //y=2.08 //x2=94.975 //y2=4.07
cc_2993 ( N_noxref_6_c_3056_n N_noxref_26_c_9913_n ) capacitor c=0.00381677f \
 //x=91.02 //y=4.705 //x2=94.975 //y2=4.07
cc_2994 ( N_noxref_6_c_3007_n N_noxref_26_c_9943_n ) capacitor c=0.0263445f \
 //x=90.905 //y=4.44 //x2=88.545 //y2=4.07
cc_2995 ( N_noxref_6_c_2898_n N_noxref_26_c_9943_n ) capacitor c=0.00128547f \
 //x=87.32 //y=2.08 //x2=88.545 //y2=4.07
cc_2996 ( N_noxref_6_c_2934_n N_noxref_26_c_9948_n ) capacitor c=0.112727f \
 //x=75.025 //y=4.81 //x2=49.715 //y2=5.155
cc_2997 ( N_noxref_6_c_2934_n N_noxref_26_c_9958_n ) capacitor c=0.0187537f \
 //x=75.025 //y=4.81 //x2=52.17 //y2=3.33
cc_2998 ( N_noxref_6_c_2934_n N_noxref_26_c_9916_n ) capacitor c=0.0139535f \
 //x=75.025 //y=4.81 //x2=54.02 //y2=2.08
cc_2999 ( N_noxref_6_c_3007_n N_noxref_26_c_9962_n ) capacitor c=0.00210648f \
 //x=90.905 //y=4.44 //x2=88.43 //y2=4.54
cc_3000 ( N_noxref_6_c_2898_n N_noxref_26_c_9962_n ) capacitor c=0.00227044f \
 //x=87.32 //y=2.08 //x2=88.43 //y2=4.54
cc_3001 ( N_noxref_6_c_3381_p N_noxref_26_c_9962_n ) capacitor c=0.00155256f \
 //x=87.955 //y=4.795 //x2=88.43 //y2=4.54
cc_3002 ( N_noxref_6_c_3054_n N_noxref_26_c_9962_n ) capacitor c=0.00180548f \
 //x=87.665 //y=4.795 //x2=88.43 //y2=4.54
cc_3003 ( N_noxref_6_c_3007_n N_noxref_26_c_9917_n ) capacitor c=0.0232321f \
 //x=90.905 //y=4.44 //x2=88.43 //y2=2.08
cc_3004 ( N_noxref_6_c_3012_n N_noxref_26_c_9917_n ) capacitor c=9.10428e-19 \
 //x=87.435 //y=4.44 //x2=88.43 //y2=2.08
cc_3005 ( N_noxref_6_c_2898_n N_noxref_26_c_9917_n ) capacitor c=0.0484612f \
 //x=87.32 //y=2.08 //x2=88.43 //y2=2.08
cc_3006 ( N_noxref_6_c_2901_n N_noxref_26_c_9917_n ) capacitor c=0.0109059f \
 //x=91.02 //y=2.08 //x2=88.43 //y2=2.08
cc_3007 ( N_noxref_6_c_2932_n N_noxref_26_c_9917_n ) capacitor c=0.00209193f \
 //x=87.32 //y=2.08 //x2=88.43 //y2=2.08
cc_3008 ( N_noxref_6_c_2934_n N_noxref_26_M126_noxref_g ) capacitor \
 c=0.00558442f //x=75.025 //y=4.81 //x2=54.22 //y2=6.02
cc_3009 ( N_noxref_6_c_2934_n N_noxref_26_M127_noxref_g ) capacitor \
 c=0.00267973f //x=75.025 //y=4.81 //x2=54.66 //y2=6.02
cc_3010 ( N_noxref_6_M168_noxref_g N_noxref_26_M170_noxref_g ) capacitor \
 c=0.010584f //x=87.59 //y=6.025 //x2=88.47 //y2=6.025
cc_3011 ( N_noxref_6_M169_noxref_g N_noxref_26_M170_noxref_g ) capacitor \
 c=0.106414f //x=88.03 //y=6.025 //x2=88.47 //y2=6.025
cc_3012 ( N_noxref_6_M169_noxref_g N_noxref_26_M171_noxref_g ) capacitor \
 c=0.0102479f //x=88.03 //y=6.025 //x2=88.91 //y2=6.025
cc_3013 ( N_noxref_6_c_2934_n N_noxref_26_c_10024_n ) capacitor c=0.00458471f \
 //x=75.025 //y=4.81 //x2=54.585 //y2=4.79
cc_3014 ( N_noxref_6_c_2934_n N_noxref_26_c_9977_n ) capacitor c=0.00184926f \
 //x=75.025 //y=4.81 //x2=54.295 //y2=4.79
cc_3015 ( N_noxref_6_c_2913_n N_noxref_26_c_10026_n ) capacitor c=4.86506e-19 \
 //x=87.495 //y=0.865 //x2=88.465 //y2=0.905
cc_3016 ( N_noxref_6_c_2915_n N_noxref_26_c_10026_n ) capacitor c=0.00152104f \
 //x=87.495 //y=1.21 //x2=88.465 //y2=0.905
cc_3017 ( N_noxref_6_c_2920_n N_noxref_26_c_10026_n ) capacitor c=0.0151475f \
 //x=88.025 //y=0.865 //x2=88.465 //y2=0.905
cc_3018 ( N_noxref_6_c_2916_n N_noxref_26_c_10029_n ) capacitor c=0.00109982f \
 //x=87.495 //y=1.52 //x2=88.465 //y2=1.25
cc_3019 ( N_noxref_6_c_2922_n N_noxref_26_c_10029_n ) capacitor c=0.0111064f \
 //x=88.025 //y=1.21 //x2=88.465 //y2=1.25
cc_3020 ( N_noxref_6_c_2916_n N_noxref_26_c_10031_n ) capacitor c=0.00182948f \
 //x=87.495 //y=1.52 //x2=88.465 //y2=1.56
cc_3021 ( N_noxref_6_c_2917_n N_noxref_26_c_10031_n ) capacitor c=0.00662747f \
 //x=87.495 //y=1.915 //x2=88.465 //y2=1.56
cc_3022 ( N_noxref_6_c_2922_n N_noxref_26_c_10031_n ) capacitor c=0.00862358f \
 //x=88.025 //y=1.21 //x2=88.465 //y2=1.56
cc_3023 ( N_noxref_6_c_3007_n N_noxref_26_c_9979_n ) capacitor c=0.0069773f \
 //x=90.905 //y=4.44 //x2=88.835 //y2=4.795
cc_3024 ( N_noxref_6_c_2920_n N_noxref_26_c_10035_n ) capacitor c=0.00124846f \
 //x=88.025 //y=0.865 //x2=88.995 //y2=0.905
cc_3025 ( N_noxref_6_c_2922_n N_noxref_26_c_10036_n ) capacitor c=0.00168739f \
 //x=88.025 //y=1.21 //x2=88.995 //y2=1.25
cc_3026 ( N_noxref_6_c_2898_n N_noxref_26_c_9931_n ) capacitor c=0.00197072f \
 //x=87.32 //y=2.08 //x2=88.43 //y2=2.08
cc_3027 ( N_noxref_6_c_2932_n N_noxref_26_c_9931_n ) capacitor c=0.00836805f \
 //x=87.32 //y=2.08 //x2=88.43 //y2=2.08
cc_3028 ( N_noxref_6_c_3007_n N_noxref_26_c_9980_n ) capacitor c=0.0014023f \
 //x=90.905 //y=4.44 //x2=88.47 //y2=4.705
cc_3029 ( N_noxref_6_c_2898_n N_noxref_26_c_9980_n ) capacitor c=0.00228787f \
 //x=87.32 //y=2.08 //x2=88.47 //y2=4.705
cc_3030 ( N_noxref_6_c_3381_p N_noxref_26_c_9980_n ) capacitor c=0.0201611f \
 //x=87.955 //y=4.795 //x2=88.47 //y2=4.705
cc_3031 ( N_noxref_6_c_3054_n N_noxref_26_c_9980_n ) capacitor c=0.00447195f \
 //x=87.665 //y=4.795 //x2=88.47 //y2=4.705
cc_3032 ( N_noxref_6_c_2925_n N_Q_c_10368_n ) capacitor c=0.00500281f \
 //x=90.825 //y=1.21 //x2=91.945 //y2=1.18
cc_3033 ( N_noxref_6_c_3416_p N_Q_c_10368_n ) capacitor c=0.00306895f \
 //x=90.825 //y=1.52 //x2=91.945 //y2=1.18
cc_3034 ( N_noxref_6_c_2927_n N_Q_c_10368_n ) capacitor c=4.02408e-19 //x=91.2 \
 //y=0.71 //x2=91.945 //y2=1.18
cc_3035 ( N_noxref_6_c_2928_n N_Q_c_10368_n ) capacitor c=0.00256926f //x=91.2 \
 //y=1.365 //x2=91.945 //y2=1.18
cc_3036 ( N_noxref_6_c_2931_n N_Q_c_10368_n ) capacitor c=0.00674619f \
 //x=91.355 //y=1.21 //x2=91.945 //y2=1.18
cc_3037 ( N_noxref_6_M14_noxref_d N_noxref_36_M12_noxref_s ) capacitor \
 c=0.00309936f //x=22.635 //y=0.915 //x2=19.695 //y2=0.375
cc_3038 ( N_noxref_6_c_2895_n N_noxref_37_c_11004_n ) capacitor c=0.00457167f \
 //x=23.225 //y=1.665 //x2=23.225 //y2=0.54
cc_3039 ( N_noxref_6_M14_noxref_d N_noxref_37_c_11004_n ) capacitor \
 c=0.0115903f //x=22.635 //y=0.915 //x2=23.225 //y2=0.54
cc_3040 ( N_noxref_6_c_3255_p N_noxref_37_c_11014_n ) capacitor c=0.0200405f \
 //x=22.91 //y=1.665 //x2=22.34 //y2=0.995
cc_3041 ( N_noxref_6_M14_noxref_d N_noxref_37_M13_noxref_d ) capacitor \
 c=5.27807e-19 //x=22.635 //y=0.915 //x2=21.1 //y2=0.91
cc_3042 ( N_noxref_6_c_2895_n N_noxref_37_M14_noxref_s ) capacitor \
 c=0.0184051f //x=23.225 //y=1.665 //x2=22.205 //y2=0.375
cc_3043 ( N_noxref_6_M14_noxref_d N_noxref_37_M14_noxref_s ) capacitor \
 c=0.0426368f //x=22.635 //y=0.915 //x2=22.205 //y2=0.375
cc_3044 ( N_noxref_6_c_2895_n N_noxref_38_c_11066_n ) capacitor c=3.84569e-19 \
 //x=23.225 //y=1.665 //x2=24.64 //y2=1.505
cc_3045 ( N_noxref_6_c_2907_n N_noxref_38_c_11066_n ) capacitor c=0.0034165f \
 //x=24.86 //y=1.915 //x2=24.64 //y2=1.505
cc_3046 ( N_noxref_6_c_2897_n N_noxref_38_c_11051_n ) capacitor c=0.0115578f \
 //x=25.16 //y=2.08 //x2=25.525 //y2=1.59
cc_3047 ( N_noxref_6_c_2906_n N_noxref_38_c_11051_n ) capacitor c=0.00697148f \
 //x=24.86 //y=1.53 //x2=25.525 //y2=1.59
cc_3048 ( N_noxref_6_c_2907_n N_noxref_38_c_11051_n ) capacitor c=0.0204849f \
 //x=24.86 //y=1.915 //x2=25.525 //y2=1.59
cc_3049 ( N_noxref_6_c_2909_n N_noxref_38_c_11051_n ) capacitor c=0.00610316f \
 //x=25.235 //y=1.375 //x2=25.525 //y2=1.59
cc_3050 ( N_noxref_6_c_2912_n N_noxref_38_c_11051_n ) capacitor c=0.00698822f \
 //x=25.39 //y=1.22 //x2=25.525 //y2=1.59
cc_3051 ( N_noxref_6_c_2903_n N_noxref_38_M15_noxref_s ) capacitor \
 c=0.0327271f //x=24.86 //y=0.875 //x2=24.505 //y2=0.375
cc_3052 ( N_noxref_6_c_2906_n N_noxref_38_M15_noxref_s ) capacitor \
 c=7.99997e-19 //x=24.86 //y=1.53 //x2=24.505 //y2=0.375
cc_3053 ( N_noxref_6_c_2907_n N_noxref_38_M15_noxref_s ) capacitor \
 c=0.00122123f //x=24.86 //y=1.915 //x2=24.505 //y2=0.375
cc_3054 ( N_noxref_6_c_2910_n N_noxref_38_M15_noxref_s ) capacitor \
 c=0.0121427f //x=25.39 //y=0.875 //x2=24.505 //y2=0.375
cc_3055 ( N_noxref_6_M14_noxref_d N_noxref_38_M15_noxref_s ) capacitor \
 c=2.55333e-19 //x=22.635 //y=0.915 //x2=24.505 //y2=0.375
cc_3056 ( N_noxref_6_c_2898_n N_noxref_64_c_12399_n ) capacitor c=0.015296f \
 //x=87.32 //y=2.08 //x2=87.275 //y2=1.495
cc_3057 ( N_noxref_6_c_2917_n N_noxref_64_c_12399_n ) capacitor c=0.0034165f \
 //x=87.495 //y=1.915 //x2=87.275 //y2=1.495
cc_3058 ( N_noxref_6_c_2932_n N_noxref_64_c_12399_n ) capacitor c=0.00780881f \
 //x=87.32 //y=2.08 //x2=87.275 //y2=1.495
cc_3059 ( N_noxref_6_c_2898_n N_noxref_64_c_12381_n ) capacitor c=0.00497226f \
 //x=87.32 //y=2.08 //x2=88.16 //y2=1.58
cc_3060 ( N_noxref_6_c_2916_n N_noxref_64_c_12381_n ) capacitor c=0.00700766f \
 //x=87.495 //y=1.52 //x2=88.16 //y2=1.58
cc_3061 ( N_noxref_6_c_2917_n N_noxref_64_c_12381_n ) capacitor c=0.0121133f \
 //x=87.495 //y=1.915 //x2=88.16 //y2=1.58
cc_3062 ( N_noxref_6_c_2919_n N_noxref_64_c_12381_n ) capacitor c=0.0103505f \
 //x=87.87 //y=1.365 //x2=88.16 //y2=1.58
cc_3063 ( N_noxref_6_c_2922_n N_noxref_64_c_12381_n ) capacitor c=0.00339872f \
 //x=88.025 //y=1.21 //x2=88.16 //y2=1.58
cc_3064 ( N_noxref_6_c_2932_n N_noxref_64_c_12381_n ) capacitor c=0.00324269f \
 //x=87.32 //y=2.08 //x2=88.16 //y2=1.58
cc_3065 ( N_noxref_6_c_2917_n N_noxref_64_c_12388_n ) capacitor c=6.71402e-19 \
 //x=87.495 //y=1.915 //x2=88.245 //y2=1.495
cc_3066 ( N_noxref_6_c_2913_n N_noxref_64_M54_noxref_s ) capacitor \
 c=0.0326926f //x=87.495 //y=0.865 //x2=87.14 //y2=0.365
cc_3067 ( N_noxref_6_c_2916_n N_noxref_64_M54_noxref_s ) capacitor \
 c=0.00110192f //x=87.495 //y=1.52 //x2=87.14 //y2=0.365
cc_3068 ( N_noxref_6_c_2920_n N_noxref_64_M54_noxref_s ) capacitor \
 c=0.0120759f //x=88.025 //y=0.865 //x2=87.14 //y2=0.365
cc_3069 ( N_noxref_6_c_2926_n N_noxref_65_c_12455_n ) capacitor c=0.0034165f \
 //x=90.825 //y=1.915 //x2=90.605 //y2=1.495
cc_3070 ( N_noxref_6_c_2901_n N_noxref_65_c_12438_n ) capacitor c=0.0107612f \
 //x=91.02 //y=2.08 //x2=91.49 //y2=1.58
cc_3071 ( N_noxref_6_c_3416_p N_noxref_65_c_12438_n ) capacitor c=0.0059182f \
 //x=90.825 //y=1.52 //x2=91.49 //y2=1.58
cc_3072 ( N_noxref_6_c_2926_n N_noxref_65_c_12438_n ) capacitor c=0.0178746f \
 //x=90.825 //y=1.915 //x2=91.49 //y2=1.58
cc_3073 ( N_noxref_6_c_2928_n N_noxref_65_c_12438_n ) capacitor c=0.00784927f \
 //x=91.2 //y=1.365 //x2=91.49 //y2=1.58
cc_3074 ( N_noxref_6_c_2931_n N_noxref_65_c_12438_n ) capacitor c=0.0059368f \
 //x=91.355 //y=1.21 //x2=91.49 //y2=1.58
cc_3075 ( N_noxref_6_c_2926_n N_noxref_65_c_12444_n ) capacitor c=0.00122123f \
 //x=90.825 //y=1.915 //x2=91.575 //y2=1.495
cc_3076 ( N_noxref_6_c_2923_n N_noxref_65_M56_noxref_s ) capacitor \
 c=0.0312776f //x=90.825 //y=0.865 //x2=90.47 //y2=0.365
cc_3077 ( N_noxref_6_c_3416_p N_noxref_65_M56_noxref_s ) capacitor \
 c=3.48408e-19 //x=90.825 //y=1.52 //x2=90.47 //y2=0.365
cc_3078 ( N_noxref_6_c_2929_n N_noxref_65_M56_noxref_s ) capacitor \
 c=0.0132463f //x=91.355 //y=0.865 //x2=90.47 //y2=0.365
cc_3079 ( N_noxref_7_c_3623_n N_noxref_8_c_3906_n ) capacitor c=0.433994f \
 //x=27.265 //y=3.7 //x2=28.005 //y2=3.33
cc_3080 ( N_noxref_7_c_3530_n N_noxref_8_c_3906_n ) capacitor c=0.0216474f \
 //x=27.38 //y=2.08 //x2=28.005 //y2=3.33
cc_3081 ( N_noxref_7_c_3623_n N_noxref_8_c_3904_n ) capacitor c=0.0293356f \
 //x=27.265 //y=3.7 //x2=22.685 //y2=3.33
cc_3082 ( N_noxref_7_c_3623_n N_noxref_8_c_3866_n ) capacitor c=0.0198345f \
 //x=27.265 //y=3.7 //x2=22.57 //y2=2.08
cc_3083 ( N_noxref_7_M94_noxref_g N_noxref_8_c_3876_n ) capacitor c=0.0162556f \
 //x=27.12 //y=6.02 //x2=27.255 //y2=5.155
cc_3084 ( N_noxref_7_M95_noxref_g N_noxref_8_c_3880_n ) capacitor c=0.0183937f \
 //x=27.56 //y=6.02 //x2=28.035 //y2=5.155
cc_3085 ( N_noxref_7_c_3660_n N_noxref_8_c_3880_n ) capacitor c=0.00201851f \
 //x=27.38 //y=4.7 //x2=28.035 //y2=5.155
cc_3086 ( N_noxref_7_c_3668_p N_noxref_8_c_3867_n ) capacitor c=0.00371277f \
 //x=27.745 //y=1.415 //x2=28.035 //y2=1.665
cc_3087 ( N_noxref_7_c_3669_p N_noxref_8_c_3867_n ) capacitor c=0.00457401f \
 //x=27.9 //y=1.26 //x2=28.035 //y2=1.665
cc_3088 ( N_noxref_7_c_3623_n N_noxref_8_c_3884_n ) capacitor c=0.00735597f \
 //x=27.265 //y=3.7 //x2=28.12 //y2=3.33
cc_3089 ( N_noxref_7_c_3530_n N_noxref_8_c_3884_n ) capacitor c=0.0763171f \
 //x=27.38 //y=2.08 //x2=28.12 //y2=3.33
cc_3090 ( N_noxref_7_c_3672_p N_noxref_8_c_3884_n ) capacitor c=0.00709342f \
 //x=27.38 //y=2.08 //x2=28.12 //y2=3.33
cc_3091 ( N_noxref_7_c_3673_p N_noxref_8_c_3884_n ) capacitor c=0.00283672f \
 //x=27.38 //y=1.915 //x2=28.12 //y2=3.33
cc_3092 ( N_noxref_7_c_3660_n N_noxref_8_c_3884_n ) capacitor c=0.0116291f \
 //x=27.38 //y=4.7 //x2=28.12 //y2=3.33
cc_3093 ( N_noxref_7_c_3530_n N_noxref_8_c_3958_n ) capacitor c=0.0126839f \
 //x=27.38 //y=2.08 //x2=27.34 //y2=5.155
cc_3094 ( N_noxref_7_c_3660_n N_noxref_8_c_3958_n ) capacitor c=0.00470675f \
 //x=27.38 //y=4.7 //x2=27.34 //y2=5.155
cc_3095 ( N_noxref_7_c_3677_p N_noxref_8_M17_noxref_d ) capacitor \
 c=0.00217566f //x=27.37 //y=0.915 //x2=27.445 //y2=0.915
cc_3096 ( N_noxref_7_c_3678_p N_noxref_8_M17_noxref_d ) capacitor c=0.0034598f \
 //x=27.37 //y=1.26 //x2=27.445 //y2=0.915
cc_3097 ( N_noxref_7_c_3679_p N_noxref_8_M17_noxref_d ) capacitor \
 c=0.00546784f //x=27.37 //y=1.57 //x2=27.445 //y2=0.915
cc_3098 ( N_noxref_7_c_3680_p N_noxref_8_M17_noxref_d ) capacitor \
 c=0.00241102f //x=27.745 //y=0.76 //x2=27.445 //y2=0.915
cc_3099 ( N_noxref_7_c_3668_p N_noxref_8_M17_noxref_d ) capacitor c=0.0138621f \
 //x=27.745 //y=1.415 //x2=27.445 //y2=0.915
cc_3100 ( N_noxref_7_c_3682_p N_noxref_8_M17_noxref_d ) capacitor \
 c=0.00219619f //x=27.9 //y=0.915 //x2=27.445 //y2=0.915
cc_3101 ( N_noxref_7_c_3669_p N_noxref_8_M17_noxref_d ) capacitor \
 c=0.00603828f //x=27.9 //y=1.26 //x2=27.445 //y2=0.915
cc_3102 ( N_noxref_7_c_3673_p N_noxref_8_M17_noxref_d ) capacitor \
 c=0.00661782f //x=27.38 //y=1.915 //x2=27.445 //y2=0.915
cc_3103 ( N_noxref_7_M94_noxref_g N_noxref_8_M94_noxref_d ) capacitor \
 c=0.0180032f //x=27.12 //y=6.02 //x2=27.195 //y2=5.02
cc_3104 ( N_noxref_7_M95_noxref_g N_noxref_8_M94_noxref_d ) capacitor \
 c=0.0194246f //x=27.56 //y=6.02 //x2=27.195 //y2=5.02
cc_3105 ( N_noxref_7_c_3577_n N_D_c_5277_n ) capacitor c=0.403974f //x=12.835 \
 //y=3.7 //x2=29.855 //y2=4.07
cc_3106 ( N_noxref_7_c_3579_n N_D_c_5277_n ) capacitor c=0.0292842f //x=8.255 \
 //y=3.7 //x2=29.855 //y2=4.07
cc_3107 ( N_noxref_7_c_3584_n N_D_c_5277_n ) capacitor c=0.468094f //x=18.385 \
 //y=3.7 //x2=29.855 //y2=4.07
cc_3108 ( N_noxref_7_c_3586_n N_D_c_5277_n ) capacitor c=0.026596f //x=13.065 \
 //y=3.7 //x2=29.855 //y2=4.07
cc_3109 ( N_noxref_7_c_3623_n N_D_c_5277_n ) capacitor c=0.792602f //x=27.265 \
 //y=3.7 //x2=29.855 //y2=4.07
cc_3110 ( N_noxref_7_c_3625_n N_D_c_5277_n ) capacitor c=0.026809f //x=18.615 \
 //y=3.7 //x2=29.855 //y2=4.07
cc_3111 ( N_noxref_7_c_3527_n N_D_c_5277_n ) capacitor c=0.0198068f //x=8.14 \
 //y=2.08 //x2=29.855 //y2=4.07
cc_3112 ( N_noxref_7_c_3528_n N_D_c_5277_n ) capacitor c=0.0198068f //x=12.95 \
 //y=2.08 //x2=29.855 //y2=4.07
cc_3113 ( N_noxref_7_c_3548_n N_D_c_5277_n ) capacitor c=0.0200135f //x=18.5 \
 //y=3.7 //x2=29.855 //y2=4.07
cc_3114 ( N_noxref_7_c_3530_n N_D_c_5277_n ) capacitor c=0.0198068f //x=27.38 \
 //y=2.08 //x2=29.855 //y2=4.07
cc_3115 ( N_noxref_7_c_3530_n N_D_c_5280_n ) capacitor c=8.68563e-19 //x=27.38 \
 //y=2.08 //x2=29.97 //y2=2.08
cc_3116 ( N_noxref_7_c_3577_n N_CLK_c_6046_n ) capacitor c=0.0344845f \
 //x=12.835 //y=3.7 //x2=16.535 //y2=4.44
cc_3117 ( N_noxref_7_c_3579_n N_CLK_c_6046_n ) capacitor c=7.0371e-19 \
 //x=8.255 //y=3.7 //x2=16.535 //y2=4.44
cc_3118 ( N_noxref_7_c_3584_n N_CLK_c_6046_n ) capacitor c=0.0246711f \
 //x=18.385 //y=3.7 //x2=16.535 //y2=4.44
cc_3119 ( N_noxref_7_c_3586_n N_CLK_c_6046_n ) capacitor c=4.78625e-19 \
 //x=13.065 //y=3.7 //x2=16.535 //y2=4.44
cc_3120 ( N_noxref_7_c_3527_n N_CLK_c_6046_n ) capacitor c=0.0200057f //x=8.14 \
 //y=2.08 //x2=16.535 //y2=4.44
cc_3121 ( N_noxref_7_c_3528_n N_CLK_c_6046_n ) capacitor c=0.0200057f \
 //x=12.95 //y=2.08 //x2=16.535 //y2=4.44
cc_3122 ( N_noxref_7_c_3538_n N_CLK_c_6046_n ) capacitor c=0.0219114f \
 //x=16.045 //y=5.155 //x2=16.535 //y2=4.44
cc_3123 ( N_noxref_7_c_3650_n N_CLK_c_6046_n ) capacitor c=0.0111881f //x=8.14 \
 //y=4.7 //x2=16.535 //y2=4.44
cc_3124 ( N_noxref_7_c_3611_n N_CLK_c_6046_n ) capacitor c=0.0111881f \
 //x=12.95 //y=4.7 //x2=16.535 //y2=4.44
cc_3125 ( N_noxref_7_c_3527_n N_CLK_c_6057_n ) capacitor c=0.00153281f \
 //x=8.14 //y=2.08 //x2=7.145 //y2=4.44
cc_3126 ( N_noxref_7_c_3584_n N_CLK_c_6058_n ) capacitor c=0.014831f \
 //x=18.385 //y=3.7 //x2=35.775 //y2=4.44
cc_3127 ( N_noxref_7_c_3623_n N_CLK_c_6058_n ) capacitor c=0.0644712f \
 //x=27.265 //y=3.7 //x2=35.775 //y2=4.44
cc_3128 ( N_noxref_7_c_3625_n N_CLK_c_6058_n ) capacitor c=4.78746e-19 \
 //x=18.615 //y=3.7 //x2=35.775 //y2=4.44
cc_3129 ( N_noxref_7_c_3544_n N_CLK_c_6058_n ) capacitor c=0.0183122f \
 //x=18.415 //y=5.155 //x2=35.775 //y2=4.44
cc_3130 ( N_noxref_7_c_3548_n N_CLK_c_6058_n ) capacitor c=0.0210274f //x=18.5 \
 //y=3.7 //x2=35.775 //y2=4.44
cc_3131 ( N_noxref_7_c_3530_n N_CLK_c_6058_n ) capacitor c=0.0178424f \
 //x=27.38 //y=2.08 //x2=35.775 //y2=4.44
cc_3132 ( N_noxref_7_c_3714_p N_CLK_c_6058_n ) capacitor c=0.0311227f \
 //x=16.84 //y=5.155 //x2=35.775 //y2=4.44
cc_3133 ( N_noxref_7_c_3660_n N_CLK_c_6058_n ) capacitor c=0.00731624f \
 //x=27.38 //y=4.7 //x2=35.775 //y2=4.44
cc_3134 ( N_noxref_7_c_3584_n N_CLK_c_6067_n ) capacitor c=6.6036e-19 \
 //x=18.385 //y=3.7 //x2=16.765 //y2=4.44
cc_3135 ( N_noxref_7_c_3534_n N_CLK_c_6067_n ) capacitor c=0.00241768f \
 //x=16.755 //y=5.155 //x2=16.765 //y2=4.44
cc_3136 ( N_noxref_7_c_3579_n N_CLK_c_6040_n ) capacitor c=0.00526349f \
 //x=8.255 //y=3.7 //x2=7.03 //y2=2.08
cc_3137 ( N_noxref_7_c_3527_n N_CLK_c_6040_n ) capacitor c=0.0446102f //x=8.14 \
 //y=2.08 //x2=7.03 //y2=2.08
cc_3138 ( N_noxref_7_c_3647_n N_CLK_c_6040_n ) capacitor c=0.00201097f \
 //x=8.14 //y=2.08 //x2=7.03 //y2=2.08
cc_3139 ( N_noxref_7_c_3650_n N_CLK_c_6040_n ) capacitor c=0.00218014f \
 //x=8.14 //y=4.7 //x2=7.03 //y2=2.08
cc_3140 ( N_noxref_7_c_3584_n N_CLK_c_6041_n ) capacitor c=0.0190398f \
 //x=18.385 //y=3.7 //x2=16.65 //y2=2.08
cc_3141 ( N_noxref_7_c_3534_n N_CLK_c_6041_n ) capacitor c=0.014564f \
 //x=16.755 //y=5.155 //x2=16.65 //y2=2.08
cc_3142 ( N_noxref_7_c_3548_n N_CLK_c_6041_n ) capacitor c=0.00256882f \
 //x=18.5 //y=3.7 //x2=16.65 //y2=2.08
cc_3143 ( N_noxref_7_M70_noxref_g N_CLK_M68_noxref_g ) capacitor c=0.0101598f \
 //x=7.88 //y=6.02 //x2=7 //y2=6.02
cc_3144 ( N_noxref_7_M70_noxref_g N_CLK_M69_noxref_g ) capacitor c=0.0602553f \
 //x=7.88 //y=6.02 //x2=7.44 //y2=6.02
cc_3145 ( N_noxref_7_M71_noxref_g N_CLK_M69_noxref_g ) capacitor c=0.0101598f \
 //x=8.32 //y=6.02 //x2=7.44 //y2=6.02
cc_3146 ( N_noxref_7_c_3534_n N_CLK_M80_noxref_g ) capacitor c=0.016514f \
 //x=16.755 //y=5.155 //x2=16.62 //y2=6.02
cc_3147 ( N_noxref_7_M80_noxref_d N_CLK_M80_noxref_g ) capacitor c=0.0180032f \
 //x=16.695 //y=5.02 //x2=16.62 //y2=6.02
cc_3148 ( N_noxref_7_c_3540_n N_CLK_M81_noxref_g ) capacitor c=0.01736f \
 //x=17.635 //y=5.155 //x2=17.06 //y2=6.02
cc_3149 ( N_noxref_7_M80_noxref_d N_CLK_M81_noxref_g ) capacitor c=0.0180032f \
 //x=16.695 //y=5.02 //x2=17.06 //y2=6.02
cc_3150 ( N_noxref_7_c_3638_n N_CLK_c_6126_n ) capacitor c=0.00456962f \
 //x=8.13 //y=0.915 //x2=7.12 //y2=0.91
cc_3151 ( N_noxref_7_c_3639_n N_CLK_c_6127_n ) capacitor c=0.00438372f \
 //x=8.13 //y=1.26 //x2=7.12 //y2=1.22
cc_3152 ( N_noxref_7_c_3640_n N_CLK_c_6128_n ) capacitor c=0.00438372f \
 //x=8.13 //y=1.57 //x2=7.12 //y2=1.45
cc_3153 ( N_noxref_7_c_3527_n N_CLK_c_6129_n ) capacitor c=0.00205895f \
 //x=8.14 //y=2.08 //x2=7.12 //y2=1.915
cc_3154 ( N_noxref_7_c_3647_n N_CLK_c_6129_n ) capacitor c=0.00828003f \
 //x=8.14 //y=2.08 //x2=7.12 //y2=1.915
cc_3155 ( N_noxref_7_c_3648_n N_CLK_c_6129_n ) capacitor c=0.00438372f \
 //x=8.14 //y=1.915 //x2=7.12 //y2=1.915
cc_3156 ( N_noxref_7_c_3650_n N_CLK_c_6179_n ) capacitor c=0.0611812f //x=8.14 \
 //y=4.7 //x2=7.365 //y2=4.79
cc_3157 ( N_noxref_7_c_3714_p N_CLK_c_6261_n ) capacitor c=0.00426767f \
 //x=16.84 //y=5.155 //x2=16.985 //y2=4.79
cc_3158 ( N_noxref_7_c_3527_n N_CLK_c_6131_n ) capacitor c=0.00142741f \
 //x=8.14 //y=2.08 //x2=7.03 //y2=4.7
cc_3159 ( N_noxref_7_c_3650_n N_CLK_c_6131_n ) capacitor c=0.00487508f \
 //x=8.14 //y=4.7 //x2=7.03 //y2=4.7
cc_3160 ( N_noxref_7_c_3534_n N_CLK_c_6160_n ) capacitor c=0.00322046f \
 //x=16.755 //y=5.155 //x2=16.65 //y2=4.7
cc_3161 ( N_noxref_7_c_3577_n N_RN_c_7021_n ) capacitor c=0.00548028f \
 //x=12.835 //y=3.7 //x2=17.645 //y2=2.22
cc_3162 ( N_noxref_7_c_3527_n N_RN_c_7021_n ) capacitor c=0.0186201f //x=8.14 \
 //y=2.08 //x2=17.645 //y2=2.22
cc_3163 ( N_noxref_7_c_3528_n N_RN_c_7021_n ) capacitor c=0.0209607f //x=12.95 \
 //y=2.08 //x2=17.645 //y2=2.22
cc_3164 ( N_noxref_7_c_3642_n N_RN_c_7021_n ) capacitor c=3.13485e-19 \
 //x=8.505 //y=1.415 //x2=17.645 //y2=2.22
cc_3165 ( N_noxref_7_c_3603_n N_RN_c_7021_n ) capacitor c=3.13485e-19 \
 //x=13.315 //y=1.415 //x2=17.645 //y2=2.22
cc_3166 ( N_noxref_7_c_3647_n N_RN_c_7021_n ) capacitor c=0.00584491f //x=8.14 \
 //y=2.08 //x2=17.645 //y2=2.22
cc_3167 ( N_noxref_7_c_3608_n N_RN_c_7021_n ) capacitor c=0.00584491f \
 //x=12.95 //y=2.08 //x2=17.645 //y2=2.22
cc_3168 ( N_noxref_7_c_3623_n N_RN_c_7033_n ) capacitor c=0.00400452f \
 //x=27.265 //y=3.7 //x2=21.345 //y2=2.22
cc_3169 ( N_noxref_7_c_3751_p N_RN_c_7033_n ) capacitor c=0.016327f //x=18.1 \
 //y=1.665 //x2=21.345 //y2=2.22
cc_3170 ( N_noxref_7_c_3548_n N_RN_c_7033_n ) capacitor c=0.0220713f //x=18.5 \
 //y=3.7 //x2=21.345 //y2=2.22
cc_3171 ( N_noxref_7_c_3548_n N_RN_c_7037_n ) capacitor c=0.0012045f //x=18.5 \
 //y=3.7 //x2=17.875 //y2=2.22
cc_3172 ( N_noxref_7_c_3623_n N_RN_c_7038_n ) capacitor c=0.00433536f \
 //x=27.265 //y=3.7 //x2=30.965 //y2=2.22
cc_3173 ( N_noxref_7_c_3530_n N_RN_c_7038_n ) capacitor c=0.0209607f //x=27.38 \
 //y=2.08 //x2=30.965 //y2=2.22
cc_3174 ( N_noxref_7_c_3668_p N_RN_c_7038_n ) capacitor c=3.13485e-19 \
 //x=27.745 //y=1.415 //x2=30.965 //y2=2.22
cc_3175 ( N_noxref_7_c_3672_p N_RN_c_7038_n ) capacitor c=0.00584491f \
 //x=27.38 //y=2.08 //x2=30.965 //y2=2.22
cc_3176 ( N_noxref_7_c_3623_n N_RN_c_7045_n ) capacitor c=3.18831e-19 \
 //x=27.265 //y=3.7 //x2=21.575 //y2=2.22
cc_3177 ( N_noxref_7_c_3584_n N_RN_c_7089_n ) capacitor c=0.0179999f \
 //x=18.385 //y=3.7 //x2=17.76 //y2=2.08
cc_3178 ( N_noxref_7_c_3625_n N_RN_c_7089_n ) capacitor c=0.00179385f \
 //x=18.615 //y=3.7 //x2=17.76 //y2=2.08
cc_3179 ( N_noxref_7_c_3548_n N_RN_c_7089_n ) capacitor c=0.0776213f //x=18.5 \
 //y=3.7 //x2=17.76 //y2=2.08
cc_3180 ( N_noxref_7_c_3762_p N_RN_c_7089_n ) capacitor c=0.0171303f //x=17.72 \
 //y=5.155 //x2=17.76 //y2=2.08
cc_3181 ( N_noxref_7_c_3623_n N_RN_c_7090_n ) capacitor c=0.0213788f \
 //x=27.265 //y=3.7 //x2=21.46 //y2=2.08
cc_3182 ( N_noxref_7_c_3548_n N_RN_c_7090_n ) capacitor c=5.91559e-19 //x=18.5 \
 //y=3.7 //x2=21.46 //y2=2.08
cc_3183 ( N_noxref_7_c_3540_n N_RN_M82_noxref_g ) capacitor c=0.01736f \
 //x=17.635 //y=5.155 //x2=17.5 //y2=6.02
cc_3184 ( N_noxref_7_M82_noxref_d N_RN_M82_noxref_g ) capacitor c=0.0180032f \
 //x=17.575 //y=5.02 //x2=17.5 //y2=6.02
cc_3185 ( N_noxref_7_c_3544_n N_RN_M83_noxref_g ) capacitor c=0.0194981f \
 //x=18.415 //y=5.155 //x2=17.94 //y2=6.02
cc_3186 ( N_noxref_7_M82_noxref_d N_RN_M83_noxref_g ) capacitor c=0.0194246f \
 //x=17.575 //y=5.02 //x2=17.94 //y2=6.02
cc_3187 ( N_noxref_7_M11_noxref_d N_RN_c_7295_n ) capacitor c=0.00217566f \
 //x=17.825 //y=0.915 //x2=17.75 //y2=0.915
cc_3188 ( N_noxref_7_M11_noxref_d N_RN_c_7296_n ) capacitor c=0.0034598f \
 //x=17.825 //y=0.915 //x2=17.75 //y2=1.26
cc_3189 ( N_noxref_7_M11_noxref_d N_RN_c_7297_n ) capacitor c=0.00546784f \
 //x=17.825 //y=0.915 //x2=17.75 //y2=1.57
cc_3190 ( N_noxref_7_M11_noxref_d N_RN_c_7298_n ) capacitor c=0.00241102f \
 //x=17.825 //y=0.915 //x2=18.125 //y2=0.76
cc_3191 ( N_noxref_7_c_3529_n N_RN_c_7299_n ) capacitor c=0.00371277f \
 //x=18.415 //y=1.665 //x2=18.125 //y2=1.415
cc_3192 ( N_noxref_7_M11_noxref_d N_RN_c_7299_n ) capacitor c=0.0138621f \
 //x=17.825 //y=0.915 //x2=18.125 //y2=1.415
cc_3193 ( N_noxref_7_M11_noxref_d N_RN_c_7301_n ) capacitor c=0.00219619f \
 //x=17.825 //y=0.915 //x2=18.28 //y2=0.915
cc_3194 ( N_noxref_7_c_3529_n N_RN_c_7302_n ) capacitor c=0.00457401f \
 //x=18.415 //y=1.665 //x2=18.28 //y2=1.26
cc_3195 ( N_noxref_7_M11_noxref_d N_RN_c_7302_n ) capacitor c=0.00603828f \
 //x=17.825 //y=0.915 //x2=18.28 //y2=1.26
cc_3196 ( N_noxref_7_c_3548_n N_RN_c_7304_n ) capacitor c=0.00709342f //x=18.5 \
 //y=3.7 //x2=17.76 //y2=2.08
cc_3197 ( N_noxref_7_c_3548_n N_RN_c_7305_n ) capacitor c=0.00283672f //x=18.5 \
 //y=3.7 //x2=17.76 //y2=1.915
cc_3198 ( N_noxref_7_M11_noxref_d N_RN_c_7305_n ) capacitor c=0.00661782f \
 //x=17.825 //y=0.915 //x2=17.76 //y2=1.915
cc_3199 ( N_noxref_7_c_3544_n N_RN_c_7307_n ) capacitor c=0.00201851f \
 //x=18.415 //y=5.155 //x2=17.76 //y2=4.7
cc_3200 ( N_noxref_7_c_3548_n N_RN_c_7307_n ) capacitor c=0.013693f //x=18.5 \
 //y=3.7 //x2=17.76 //y2=4.7
cc_3201 ( N_noxref_7_c_3762_p N_RN_c_7307_n ) capacitor c=0.00475601f \
 //x=17.72 //y=5.155 //x2=17.76 //y2=4.7
cc_3202 ( N_noxref_7_c_3577_n N_SN_c_8129_n ) capacitor c=0.0092394f \
 //x=12.835 //y=3.7 //x2=26.155 //y2=2.96
cc_3203 ( N_noxref_7_c_3584_n N_SN_c_8129_n ) capacitor c=0.041794f //x=18.385 \
 //y=3.7 //x2=26.155 //y2=2.96
cc_3204 ( N_noxref_7_c_3586_n N_SN_c_8129_n ) capacitor c=6.03896e-19 \
 //x=13.065 //y=3.7 //x2=26.155 //y2=2.96
cc_3205 ( N_noxref_7_c_3623_n N_SN_c_8129_n ) capacitor c=0.119625f //x=27.265 \
 //y=3.7 //x2=26.155 //y2=2.96
cc_3206 ( N_noxref_7_c_3625_n N_SN_c_8129_n ) capacitor c=4.80612e-19 \
 //x=18.615 //y=3.7 //x2=26.155 //y2=2.96
cc_3207 ( N_noxref_7_c_3528_n N_SN_c_8129_n ) capacitor c=0.0202855f //x=12.95 \
 //y=2.08 //x2=26.155 //y2=2.96
cc_3208 ( N_noxref_7_c_3548_n N_SN_c_8129_n ) capacitor c=0.0210712f //x=18.5 \
 //y=3.7 //x2=26.155 //y2=2.96
cc_3209 ( N_noxref_7_c_3577_n N_SN_c_8183_n ) capacitor c=9.83937e-19 \
 //x=12.835 //y=3.7 //x2=11.955 //y2=2.96
cc_3210 ( N_noxref_7_c_3528_n N_SN_c_8183_n ) capacitor c=0.00128547f \
 //x=12.95 //y=2.08 //x2=11.955 //y2=2.96
cc_3211 ( N_noxref_7_c_3623_n N_SN_c_8132_n ) capacitor c=0.0101624f \
 //x=27.265 //y=3.7 //x2=40.585 //y2=2.96
cc_3212 ( N_noxref_7_c_3530_n N_SN_c_8132_n ) capacitor c=0.0202855f //x=27.38 \
 //y=2.08 //x2=40.585 //y2=2.96
cc_3213 ( N_noxref_7_c_3623_n N_SN_c_8226_n ) capacitor c=6.65965e-19 \
 //x=27.265 //y=3.7 //x2=26.385 //y2=2.96
cc_3214 ( N_noxref_7_c_3530_n N_SN_c_8226_n ) capacitor c=0.00128547f \
 //x=27.38 //y=2.08 //x2=26.385 //y2=2.96
cc_3215 ( N_noxref_7_c_3577_n N_SN_c_8145_n ) capacitor c=0.0190398f \
 //x=12.835 //y=3.7 //x2=11.84 //y2=2.08
cc_3216 ( N_noxref_7_c_3586_n N_SN_c_8145_n ) capacitor c=0.00128547f \
 //x=13.065 //y=3.7 //x2=11.84 //y2=2.08
cc_3217 ( N_noxref_7_c_3528_n N_SN_c_8145_n ) capacitor c=0.0432923f //x=12.95 \
 //y=2.08 //x2=11.84 //y2=2.08
cc_3218 ( N_noxref_7_c_3608_n N_SN_c_8145_n ) capacitor c=0.00201097f \
 //x=12.95 //y=2.08 //x2=11.84 //y2=2.08
cc_3219 ( N_noxref_7_c_3611_n N_SN_c_8145_n ) capacitor c=0.00219458f \
 //x=12.95 //y=4.7 //x2=11.84 //y2=2.08
cc_3220 ( N_noxref_7_c_3623_n N_SN_c_8146_n ) capacitor c=0.0203253f \
 //x=27.265 //y=3.7 //x2=26.27 //y2=2.08
cc_3221 ( N_noxref_7_c_3530_n N_SN_c_8146_n ) capacitor c=0.0415826f //x=27.38 \
 //y=2.08 //x2=26.27 //y2=2.08
cc_3222 ( N_noxref_7_c_3672_p N_SN_c_8146_n ) capacitor c=0.00201097f \
 //x=27.38 //y=2.08 //x2=26.27 //y2=2.08
cc_3223 ( N_noxref_7_c_3660_n N_SN_c_8146_n ) capacitor c=0.00197875f \
 //x=27.38 //y=4.7 //x2=26.27 //y2=2.08
cc_3224 ( N_noxref_7_M76_noxref_g N_SN_M74_noxref_g ) capacitor c=0.0101598f \
 //x=12.69 //y=6.02 //x2=11.81 //y2=6.02
cc_3225 ( N_noxref_7_M76_noxref_g N_SN_M75_noxref_g ) capacitor c=0.0602553f \
 //x=12.69 //y=6.02 //x2=12.25 //y2=6.02
cc_3226 ( N_noxref_7_M77_noxref_g N_SN_M75_noxref_g ) capacitor c=0.0101598f \
 //x=13.13 //y=6.02 //x2=12.25 //y2=6.02
cc_3227 ( N_noxref_7_M94_noxref_g N_SN_M92_noxref_g ) capacitor c=0.0100903f \
 //x=27.12 //y=6.02 //x2=26.24 //y2=6.02
cc_3228 ( N_noxref_7_M94_noxref_g N_SN_M93_noxref_g ) capacitor c=0.0600064f \
 //x=27.12 //y=6.02 //x2=26.68 //y2=6.02
cc_3229 ( N_noxref_7_M95_noxref_g N_SN_M93_noxref_g ) capacitor c=0.0100903f \
 //x=27.56 //y=6.02 //x2=26.68 //y2=6.02
cc_3230 ( N_noxref_7_c_3599_n N_SN_c_8197_n ) capacitor c=0.00456962f \
 //x=12.94 //y=0.915 //x2=11.93 //y2=0.91
cc_3231 ( N_noxref_7_c_3600_n N_SN_c_8198_n ) capacitor c=0.00438372f \
 //x=12.94 //y=1.26 //x2=11.93 //y2=1.22
cc_3232 ( N_noxref_7_c_3601_n N_SN_c_8199_n ) capacitor c=0.00438372f \
 //x=12.94 //y=1.57 //x2=11.93 //y2=1.45
cc_3233 ( N_noxref_7_c_3528_n N_SN_c_8200_n ) capacitor c=0.00205895f \
 //x=12.95 //y=2.08 //x2=11.93 //y2=1.915
cc_3234 ( N_noxref_7_c_3608_n N_SN_c_8200_n ) capacitor c=0.00828003f \
 //x=12.95 //y=2.08 //x2=11.93 //y2=1.915
cc_3235 ( N_noxref_7_c_3609_n N_SN_c_8200_n ) capacitor c=0.00438372f \
 //x=12.95 //y=1.915 //x2=11.93 //y2=1.915
cc_3236 ( N_noxref_7_c_3611_n N_SN_c_8215_n ) capacitor c=0.0611812f //x=12.95 \
 //y=4.7 //x2=12.175 //y2=4.79
cc_3237 ( N_noxref_7_c_3677_p N_SN_c_8254_n ) capacitor c=0.00456962f \
 //x=27.37 //y=0.915 //x2=26.36 //y2=0.91
cc_3238 ( N_noxref_7_c_3678_p N_SN_c_8255_n ) capacitor c=0.00438372f \
 //x=27.37 //y=1.26 //x2=26.36 //y2=1.22
cc_3239 ( N_noxref_7_c_3679_p N_SN_c_8256_n ) capacitor c=0.00438372f \
 //x=27.37 //y=1.57 //x2=26.36 //y2=1.45
cc_3240 ( N_noxref_7_c_3530_n N_SN_c_8257_n ) capacitor c=0.00205895f \
 //x=27.38 //y=2.08 //x2=26.36 //y2=1.915
cc_3241 ( N_noxref_7_c_3672_p N_SN_c_8257_n ) capacitor c=0.00828003f \
 //x=27.38 //y=2.08 //x2=26.36 //y2=1.915
cc_3242 ( N_noxref_7_c_3673_p N_SN_c_8257_n ) capacitor c=0.00438372f \
 //x=27.38 //y=1.915 //x2=26.36 //y2=1.915
cc_3243 ( N_noxref_7_c_3660_n N_SN_c_8259_n ) capacitor c=0.0609323f //x=27.38 \
 //y=4.7 //x2=26.605 //y2=4.79
cc_3244 ( N_noxref_7_c_3528_n N_SN_c_8202_n ) capacitor c=0.00142741f \
 //x=12.95 //y=2.08 //x2=11.84 //y2=4.7
cc_3245 ( N_noxref_7_c_3611_n N_SN_c_8202_n ) capacitor c=0.00487508f \
 //x=12.95 //y=4.7 //x2=11.84 //y2=4.7
cc_3246 ( N_noxref_7_c_3530_n N_SN_c_8264_n ) capacitor c=0.00142741f \
 //x=27.38 //y=2.08 //x2=26.27 //y2=4.7
cc_3247 ( N_noxref_7_c_3660_n N_SN_c_8264_n ) capacitor c=0.00487508f \
 //x=27.38 //y=4.7 //x2=26.27 //y2=4.7
cc_3248 ( N_noxref_7_c_3527_n N_noxref_31_c_10697_n ) capacitor c=0.00204385f \
 //x=8.14 //y=2.08 //x2=8.795 //y2=0.54
cc_3249 ( N_noxref_7_c_3638_n N_noxref_31_c_10697_n ) capacitor c=0.0194423f \
 //x=8.13 //y=0.915 //x2=8.795 //y2=0.54
cc_3250 ( N_noxref_7_c_3644_n N_noxref_31_c_10697_n ) capacitor c=0.00656458f \
 //x=8.66 //y=0.915 //x2=8.795 //y2=0.54
cc_3251 ( N_noxref_7_c_3647_n N_noxref_31_c_10697_n ) capacitor c=2.20712e-19 \
 //x=8.14 //y=2.08 //x2=8.795 //y2=0.54
cc_3252 ( N_noxref_7_c_3639_n N_noxref_31_c_10707_n ) capacitor c=0.00538829f \
 //x=8.13 //y=1.26 //x2=7.91 //y2=0.995
cc_3253 ( N_noxref_7_c_3638_n N_noxref_31_M5_noxref_s ) capacitor \
 c=0.00538829f //x=8.13 //y=0.915 //x2=7.775 //y2=0.375
cc_3254 ( N_noxref_7_c_3640_n N_noxref_31_M5_noxref_s ) capacitor \
 c=0.00538829f //x=8.13 //y=1.57 //x2=7.775 //y2=0.375
cc_3255 ( N_noxref_7_c_3644_n N_noxref_31_M5_noxref_s ) capacitor c=0.0143002f \
 //x=8.66 //y=0.915 //x2=7.775 //y2=0.375
cc_3256 ( N_noxref_7_c_3645_n N_noxref_31_M5_noxref_s ) capacitor \
 c=0.00290153f //x=8.66 //y=1.26 //x2=7.775 //y2=0.375
cc_3257 ( N_noxref_7_c_3528_n N_noxref_33_c_10798_n ) capacitor c=0.00204385f \
 //x=12.95 //y=2.08 //x2=13.605 //y2=0.54
cc_3258 ( N_noxref_7_c_3599_n N_noxref_33_c_10798_n ) capacitor c=0.0194423f \
 //x=12.94 //y=0.915 //x2=13.605 //y2=0.54
cc_3259 ( N_noxref_7_c_3605_n N_noxref_33_c_10798_n ) capacitor c=0.00656458f \
 //x=13.47 //y=0.915 //x2=13.605 //y2=0.54
cc_3260 ( N_noxref_7_c_3608_n N_noxref_33_c_10798_n ) capacitor c=2.20712e-19 \
 //x=12.95 //y=2.08 //x2=13.605 //y2=0.54
cc_3261 ( N_noxref_7_c_3600_n N_noxref_33_c_10808_n ) capacitor c=0.00538829f \
 //x=12.94 //y=1.26 //x2=12.72 //y2=0.995
cc_3262 ( N_noxref_7_c_3599_n N_noxref_33_M8_noxref_s ) capacitor \
 c=0.00538829f //x=12.94 //y=0.915 //x2=12.585 //y2=0.375
cc_3263 ( N_noxref_7_c_3601_n N_noxref_33_M8_noxref_s ) capacitor \
 c=0.00538829f //x=12.94 //y=1.57 //x2=12.585 //y2=0.375
cc_3264 ( N_noxref_7_c_3605_n N_noxref_33_M8_noxref_s ) capacitor c=0.0143002f \
 //x=13.47 //y=0.915 //x2=12.585 //y2=0.375
cc_3265 ( N_noxref_7_c_3606_n N_noxref_33_M8_noxref_s ) capacitor \
 c=0.00290153f //x=13.47 //y=1.26 //x2=12.585 //y2=0.375
cc_3266 ( N_noxref_7_M11_noxref_d N_noxref_34_M9_noxref_s ) capacitor \
 c=0.00309936f //x=17.825 //y=0.915 //x2=14.885 //y2=0.375
cc_3267 ( N_noxref_7_c_3529_n N_noxref_35_c_10899_n ) capacitor c=0.00457167f \
 //x=18.415 //y=1.665 //x2=18.415 //y2=0.54
cc_3268 ( N_noxref_7_M11_noxref_d N_noxref_35_c_10899_n ) capacitor \
 c=0.0115903f //x=17.825 //y=0.915 //x2=18.415 //y2=0.54
cc_3269 ( N_noxref_7_c_3751_p N_noxref_35_c_10909_n ) capacitor c=0.0200405f \
 //x=18.1 //y=1.665 //x2=17.53 //y2=0.995
cc_3270 ( N_noxref_7_M11_noxref_d N_noxref_35_M10_noxref_d ) capacitor \
 c=5.27807e-19 //x=17.825 //y=0.915 //x2=16.29 //y2=0.91
cc_3271 ( N_noxref_7_c_3529_n N_noxref_35_M11_noxref_s ) capacitor \
 c=0.0196084f //x=18.415 //y=1.665 //x2=17.395 //y2=0.375
cc_3272 ( N_noxref_7_M11_noxref_d N_noxref_35_M11_noxref_s ) capacitor \
 c=0.0426368f //x=17.825 //y=0.915 //x2=17.395 //y2=0.375
cc_3273 ( N_noxref_7_c_3529_n N_noxref_36_c_10962_n ) capacitor c=3.84569e-19 \
 //x=18.415 //y=1.665 //x2=19.83 //y2=1.505
cc_3274 ( N_noxref_7_M11_noxref_d N_noxref_36_M12_noxref_s ) capacitor \
 c=2.55333e-19 //x=17.825 //y=0.915 //x2=19.695 //y2=0.375
cc_3275 ( N_noxref_7_c_3530_n N_noxref_39_c_11105_n ) capacitor c=0.00204385f \
 //x=27.38 //y=2.08 //x2=28.035 //y2=0.54
cc_3276 ( N_noxref_7_c_3677_p N_noxref_39_c_11105_n ) capacitor c=0.0194423f \
 //x=27.37 //y=0.915 //x2=28.035 //y2=0.54
cc_3277 ( N_noxref_7_c_3682_p N_noxref_39_c_11105_n ) capacitor c=0.00656458f \
 //x=27.9 //y=0.915 //x2=28.035 //y2=0.54
cc_3278 ( N_noxref_7_c_3672_p N_noxref_39_c_11105_n ) capacitor c=2.20712e-19 \
 //x=27.38 //y=2.08 //x2=28.035 //y2=0.54
cc_3279 ( N_noxref_7_c_3678_p N_noxref_39_c_11117_n ) capacitor c=0.00538829f \
 //x=27.37 //y=1.26 //x2=27.15 //y2=0.995
cc_3280 ( N_noxref_7_c_3677_p N_noxref_39_M17_noxref_s ) capacitor \
 c=0.00538829f //x=27.37 //y=0.915 //x2=27.015 //y2=0.375
cc_3281 ( N_noxref_7_c_3679_p N_noxref_39_M17_noxref_s ) capacitor \
 c=0.00538829f //x=27.37 //y=1.57 //x2=27.015 //y2=0.375
cc_3282 ( N_noxref_7_c_3682_p N_noxref_39_M17_noxref_s ) capacitor \
 c=0.0143002f //x=27.9 //y=0.915 //x2=27.015 //y2=0.375
cc_3283 ( N_noxref_7_c_3669_p N_noxref_39_M17_noxref_s ) capacitor \
 c=0.00290153f //x=27.9 //y=1.26 //x2=27.015 //y2=0.375
cc_3284 ( N_noxref_8_c_3880_n N_noxref_9_c_4075_n ) capacitor c=3.10026e-19 \
 //x=28.035 //y=5.155 //x2=30.475 //y2=5.155
cc_3285 ( N_noxref_8_c_3906_n N_noxref_11_c_4533_n ) capacitor c=0.00359266f \
 //x=28.005 //y=3.33 //x2=32.305 //y2=3.33
cc_3286 ( N_noxref_8_c_3906_n N_D_c_5277_n ) capacitor c=0.0693839f //x=28.005 \
 //y=3.33 //x2=29.855 //y2=4.07
cc_3287 ( N_noxref_8_c_3904_n N_D_c_5277_n ) capacitor c=7.1286e-19 //x=22.685 \
 //y=3.33 //x2=29.855 //y2=4.07
cc_3288 ( N_noxref_8_c_3866_n N_D_c_5277_n ) capacitor c=0.0179722f //x=22.57 \
 //y=2.08 //x2=29.855 //y2=4.07
cc_3289 ( N_noxref_8_c_3884_n N_D_c_5277_n ) capacitor c=0.0208368f //x=28.12 \
 //y=3.33 //x2=29.855 //y2=4.07
cc_3290 ( N_noxref_8_c_3884_n N_D_c_5334_n ) capacitor c=3.50683e-19 //x=28.12 \
 //y=3.33 //x2=30.085 //y2=4.07
cc_3291 ( N_noxref_8_c_3906_n N_D_c_5280_n ) capacitor c=0.00186218f \
 //x=28.005 //y=3.33 //x2=29.97 //y2=2.08
cc_3292 ( N_noxref_8_c_3884_n N_D_c_5280_n ) capacitor c=0.0130123f //x=28.12 \
 //y=3.33 //x2=29.97 //y2=2.08
cc_3293 ( N_noxref_8_c_3906_n N_CLK_c_6058_n ) capacitor c=0.00412696f \
 //x=28.005 //y=3.33 //x2=35.775 //y2=4.44
cc_3294 ( N_noxref_8_c_3866_n N_CLK_c_6058_n ) capacitor c=0.0200057f \
 //x=22.57 //y=2.08 //x2=35.775 //y2=4.44
cc_3295 ( N_noxref_8_c_3884_n N_CLK_c_6058_n ) capacitor c=0.0166101f \
 //x=28.12 //y=3.33 //x2=35.775 //y2=4.44
cc_3296 ( N_noxref_8_c_3939_n N_CLK_c_6058_n ) capacitor c=0.0111881f \
 //x=22.57 //y=4.7 //x2=35.775 //y2=4.44
cc_3297 ( N_noxref_8_c_3906_n N_RN_c_7038_n ) capacitor c=0.0225411f \
 //x=28.005 //y=3.33 //x2=30.965 //y2=2.22
cc_3298 ( N_noxref_8_c_3904_n N_RN_c_7038_n ) capacitor c=7.32243e-19 \
 //x=22.685 //y=3.33 //x2=30.965 //y2=2.22
cc_3299 ( N_noxref_8_c_3866_n N_RN_c_7038_n ) capacitor c=0.0209607f //x=22.57 \
 //y=2.08 //x2=30.965 //y2=2.22
cc_3300 ( N_noxref_8_c_3986_p N_RN_c_7038_n ) capacitor c=0.016327f //x=27.72 \
 //y=1.665 //x2=30.965 //y2=2.22
cc_3301 ( N_noxref_8_c_3884_n N_RN_c_7038_n ) capacitor c=0.0220713f //x=28.12 \
 //y=3.33 //x2=30.965 //y2=2.22
cc_3302 ( N_noxref_8_c_3931_n N_RN_c_7038_n ) capacitor c=3.13485e-19 \
 //x=22.935 //y=1.415 //x2=30.965 //y2=2.22
cc_3303 ( N_noxref_8_c_3936_n N_RN_c_7038_n ) capacitor c=0.00584491f \
 //x=22.57 //y=2.08 //x2=30.965 //y2=2.22
cc_3304 ( N_noxref_8_c_3866_n N_RN_c_7045_n ) capacitor c=0.00165648f \
 //x=22.57 //y=2.08 //x2=21.575 //y2=2.22
cc_3305 ( N_noxref_8_c_3936_n N_RN_c_7045_n ) capacitor c=2.3323e-19 //x=22.57 \
 //y=2.08 //x2=21.575 //y2=2.22
cc_3306 ( N_noxref_8_c_3904_n N_RN_c_7090_n ) capacitor c=0.0027353f \
 //x=22.685 //y=3.33 //x2=21.46 //y2=2.08
cc_3307 ( N_noxref_8_c_3866_n N_RN_c_7090_n ) capacitor c=0.044753f //x=22.57 \
 //y=2.08 //x2=21.46 //y2=2.08
cc_3308 ( N_noxref_8_c_3936_n N_RN_c_7090_n ) capacitor c=0.0019893f //x=22.57 \
 //y=2.08 //x2=21.46 //y2=2.08
cc_3309 ( N_noxref_8_c_3939_n N_RN_c_7090_n ) capacitor c=0.00219458f \
 //x=22.57 //y=4.7 //x2=21.46 //y2=2.08
cc_3310 ( N_noxref_8_c_3884_n N_RN_c_7091_n ) capacitor c=6.3801e-19 //x=28.12 \
 //y=3.33 //x2=31.08 //y2=2.08
cc_3311 ( N_noxref_8_M88_noxref_g N_RN_M86_noxref_g ) capacitor c=0.0101598f \
 //x=22.31 //y=6.02 //x2=21.43 //y2=6.02
cc_3312 ( N_noxref_8_M88_noxref_g N_RN_M87_noxref_g ) capacitor c=0.0602553f \
 //x=22.31 //y=6.02 //x2=21.87 //y2=6.02
cc_3313 ( N_noxref_8_M89_noxref_g N_RN_M87_noxref_g ) capacitor c=0.0101598f \
 //x=22.75 //y=6.02 //x2=21.87 //y2=6.02
cc_3314 ( N_noxref_8_c_3927_n N_RN_c_7216_n ) capacitor c=0.00456962f \
 //x=22.56 //y=0.915 //x2=21.55 //y2=0.91
cc_3315 ( N_noxref_8_c_3928_n N_RN_c_7217_n ) capacitor c=0.00438372f \
 //x=22.56 //y=1.26 //x2=21.55 //y2=1.22
cc_3316 ( N_noxref_8_c_3929_n N_RN_c_7218_n ) capacitor c=0.00438372f \
 //x=22.56 //y=1.57 //x2=21.55 //y2=1.45
cc_3317 ( N_noxref_8_c_3866_n N_RN_c_7219_n ) capacitor c=0.00205895f \
 //x=22.57 //y=2.08 //x2=21.55 //y2=1.915
cc_3318 ( N_noxref_8_c_3936_n N_RN_c_7219_n ) capacitor c=0.00828003f \
 //x=22.57 //y=2.08 //x2=21.55 //y2=1.915
cc_3319 ( N_noxref_8_c_3937_n N_RN_c_7219_n ) capacitor c=0.00438372f \
 //x=22.57 //y=1.915 //x2=21.55 //y2=1.915
cc_3320 ( N_noxref_8_c_3939_n N_RN_c_7255_n ) capacitor c=0.0611812f //x=22.57 \
 //y=4.7 //x2=21.795 //y2=4.79
cc_3321 ( N_noxref_8_c_3866_n N_RN_c_7223_n ) capacitor c=0.00142741f \
 //x=22.57 //y=2.08 //x2=21.46 //y2=4.7
cc_3322 ( N_noxref_8_c_3939_n N_RN_c_7223_n ) capacitor c=0.00487508f \
 //x=22.57 //y=4.7 //x2=21.46 //y2=4.7
cc_3323 ( N_noxref_8_c_3906_n N_SN_c_8129_n ) capacitor c=0.30592f //x=28.005 \
 //y=3.33 //x2=26.155 //y2=2.96
cc_3324 ( N_noxref_8_c_3904_n N_SN_c_8129_n ) capacitor c=0.0291389f \
 //x=22.685 //y=3.33 //x2=26.155 //y2=2.96
cc_3325 ( N_noxref_8_c_3866_n N_SN_c_8129_n ) capacitor c=0.0221202f //x=22.57 \
 //y=2.08 //x2=26.155 //y2=2.96
cc_3326 ( N_noxref_8_c_3906_n N_SN_c_8132_n ) capacitor c=0.170628f //x=28.005 \
 //y=3.33 //x2=40.585 //y2=2.96
cc_3327 ( N_noxref_8_c_3884_n N_SN_c_8132_n ) capacitor c=0.0229057f //x=28.12 \
 //y=3.33 //x2=40.585 //y2=2.96
cc_3328 ( N_noxref_8_c_3906_n N_SN_c_8226_n ) capacitor c=0.0265806f \
 //x=28.005 //y=3.33 //x2=26.385 //y2=2.96
cc_3329 ( N_noxref_8_c_3906_n N_SN_c_8146_n ) capacitor c=0.0208912f \
 //x=28.005 //y=3.33 //x2=26.27 //y2=2.08
cc_3330 ( N_noxref_8_c_3870_n N_SN_c_8146_n ) capacitor c=0.0121898f \
 //x=26.375 //y=5.155 //x2=26.27 //y2=2.08
cc_3331 ( N_noxref_8_c_3884_n N_SN_c_8146_n ) capacitor c=0.00267392f \
 //x=28.12 //y=3.33 //x2=26.27 //y2=2.08
cc_3332 ( N_noxref_8_c_3870_n N_SN_M92_noxref_g ) capacitor c=0.0163793f \
 //x=26.375 //y=5.155 //x2=26.24 //y2=6.02
cc_3333 ( N_noxref_8_M92_noxref_d N_SN_M92_noxref_g ) capacitor c=0.0180032f \
 //x=26.315 //y=5.02 //x2=26.24 //y2=6.02
cc_3334 ( N_noxref_8_c_3876_n N_SN_M93_noxref_g ) capacitor c=0.0162556f \
 //x=27.255 //y=5.155 //x2=26.68 //y2=6.02
cc_3335 ( N_noxref_8_M92_noxref_d N_SN_M93_noxref_g ) capacitor c=0.0180032f \
 //x=26.315 //y=5.02 //x2=26.68 //y2=6.02
cc_3336 ( N_noxref_8_c_4022_p N_SN_c_8259_n ) capacitor c=0.00392095f \
 //x=26.46 //y=5.155 //x2=26.605 //y2=4.79
cc_3337 ( N_noxref_8_c_3870_n N_SN_c_8264_n ) capacitor c=0.00309994f \
 //x=26.375 //y=5.155 //x2=26.27 //y2=4.7
cc_3338 ( N_noxref_8_c_3866_n N_noxref_37_c_11004_n ) capacitor c=0.00204385f \
 //x=22.57 //y=2.08 //x2=23.225 //y2=0.54
cc_3339 ( N_noxref_8_c_3927_n N_noxref_37_c_11004_n ) capacitor c=0.0194423f \
 //x=22.56 //y=0.915 //x2=23.225 //y2=0.54
cc_3340 ( N_noxref_8_c_3933_n N_noxref_37_c_11004_n ) capacitor c=0.00656458f \
 //x=23.09 //y=0.915 //x2=23.225 //y2=0.54
cc_3341 ( N_noxref_8_c_3936_n N_noxref_37_c_11004_n ) capacitor c=2.20712e-19 \
 //x=22.57 //y=2.08 //x2=23.225 //y2=0.54
cc_3342 ( N_noxref_8_c_3928_n N_noxref_37_c_11014_n ) capacitor c=0.00538829f \
 //x=22.56 //y=1.26 //x2=22.34 //y2=0.995
cc_3343 ( N_noxref_8_c_3927_n N_noxref_37_M14_noxref_s ) capacitor \
 c=0.00538829f //x=22.56 //y=0.915 //x2=22.205 //y2=0.375
cc_3344 ( N_noxref_8_c_3929_n N_noxref_37_M14_noxref_s ) capacitor \
 c=0.00538829f //x=22.56 //y=1.57 //x2=22.205 //y2=0.375
cc_3345 ( N_noxref_8_c_3933_n N_noxref_37_M14_noxref_s ) capacitor \
 c=0.0143002f //x=23.09 //y=0.915 //x2=22.205 //y2=0.375
cc_3346 ( N_noxref_8_c_3934_n N_noxref_37_M14_noxref_s ) capacitor \
 c=0.00290153f //x=23.09 //y=1.26 //x2=22.205 //y2=0.375
cc_3347 ( N_noxref_8_M17_noxref_d N_noxref_38_M15_noxref_s ) capacitor \
 c=0.00309936f //x=27.445 //y=0.915 //x2=24.505 //y2=0.375
cc_3348 ( N_noxref_8_c_3867_n N_noxref_39_c_11105_n ) capacitor c=0.00457167f \
 //x=28.035 //y=1.665 //x2=28.035 //y2=0.54
cc_3349 ( N_noxref_8_M17_noxref_d N_noxref_39_c_11105_n ) capacitor \
 c=0.0115903f //x=27.445 //y=0.915 //x2=28.035 //y2=0.54
cc_3350 ( N_noxref_8_c_3986_p N_noxref_39_c_11117_n ) capacitor c=0.0200405f \
 //x=27.72 //y=1.665 //x2=27.15 //y2=0.995
cc_3351 ( N_noxref_8_M17_noxref_d N_noxref_39_M16_noxref_d ) capacitor \
 c=5.27807e-19 //x=27.445 //y=0.915 //x2=25.91 //y2=0.91
cc_3352 ( N_noxref_8_c_3867_n N_noxref_39_M17_noxref_s ) capacitor \
 c=0.0196084f //x=28.035 //y=1.665 //x2=27.015 //y2=0.375
cc_3353 ( N_noxref_8_M17_noxref_d N_noxref_39_M17_noxref_s ) capacitor \
 c=0.0426368f //x=27.445 //y=0.915 //x2=27.015 //y2=0.375
cc_3354 ( N_noxref_8_c_3867_n N_noxref_40_c_11167_n ) capacitor c=3.84569e-19 \
 //x=28.035 //y=1.665 //x2=29.45 //y2=1.505
cc_3355 ( N_noxref_8_M17_noxref_d N_noxref_40_M18_noxref_s ) capacitor \
 c=2.55333e-19 //x=27.445 //y=0.915 //x2=29.315 //y2=0.375
cc_3356 ( N_noxref_9_c_4044_n N_noxref_10_c_4296_n ) capacitor c=0.00564994f \
 //x=39.475 //y=2.59 //x2=42.665 //y2=2.59
cc_3357 ( N_noxref_9_M109_noxref_g N_noxref_10_c_4311_n ) capacitor \
 c=0.0157304f //x=40.23 //y=6.02 //x2=40.805 //y2=5.155
cc_3358 ( N_noxref_9_M108_noxref_g N_noxref_10_c_4315_n ) capacitor \
 c=0.0213876f //x=39.79 //y=6.02 //x2=40.095 //y2=5.155
cc_3359 ( N_noxref_9_c_4129_n N_noxref_10_c_4315_n ) capacitor c=0.00393496f \
 //x=40.155 //y=4.79 //x2=40.095 //y2=5.155
cc_3360 ( N_noxref_9_M109_noxref_g N_noxref_10_M108_noxref_d ) capacitor \
 c=0.0180032f //x=40.23 //y=6.02 //x2=39.865 //y2=5.02
cc_3361 ( N_noxref_9_c_4042_n N_noxref_11_c_4534_n ) capacitor c=0.0111384f \
 //x=34.665 //y=2.59 //x2=37.625 //y2=3.33
cc_3362 ( N_noxref_9_c_4043_n N_noxref_11_c_4534_n ) capacitor c=8.87672e-19 \
 //x=33.045 //y=2.59 //x2=37.625 //y2=3.33
cc_3363 ( N_noxref_9_c_4044_n N_noxref_11_c_4534_n ) capacitor c=0.0246405f \
 //x=39.475 //y=2.59 //x2=37.625 //y2=3.33
cc_3364 ( N_noxref_9_c_4045_n N_noxref_11_c_4534_n ) capacitor c=5.36573e-19 \
 //x=34.895 //y=2.59 //x2=37.625 //y2=3.33
cc_3365 ( N_noxref_9_c_4047_n N_noxref_11_c_4534_n ) capacitor c=0.0211097f \
 //x=32.93 //y=2.59 //x2=37.625 //y2=3.33
cc_3366 ( N_noxref_9_c_4048_n N_noxref_11_c_4534_n ) capacitor c=0.0221185f \
 //x=34.78 //y=2.08 //x2=37.625 //y2=3.33
cc_3367 ( N_noxref_9_c_4047_n N_noxref_11_c_4533_n ) capacitor c=0.00179385f \
 //x=32.93 //y=2.59 //x2=32.305 //y2=3.33
cc_3368 ( N_noxref_9_c_4044_n N_noxref_11_c_4541_n ) capacitor c=0.0118993f \
 //x=39.475 //y=2.59 //x2=49.095 //y2=3.33
cc_3369 ( N_noxref_9_c_4049_n N_noxref_11_c_4541_n ) capacitor c=0.0197803f \
 //x=39.59 //y=2.08 //x2=49.095 //y2=3.33
cc_3370 ( N_noxref_9_c_4044_n N_noxref_11_c_4543_n ) capacitor c=5.76706e-19 \
 //x=39.475 //y=2.59 //x2=37.855 //y2=3.33
cc_3371 ( N_noxref_9_c_4049_n N_noxref_11_c_4543_n ) capacitor c=7.01366e-19 \
 //x=39.59 //y=2.08 //x2=37.855 //y2=3.33
cc_3372 ( N_noxref_9_c_4043_n N_noxref_11_c_4464_n ) capacitor c=0.00687545f \
 //x=33.045 //y=2.59 //x2=32.19 //y2=2.08
cc_3373 ( N_noxref_9_c_4047_n N_noxref_11_c_4464_n ) capacitor c=0.0766861f \
 //x=32.93 //y=2.59 //x2=32.19 //y2=2.08
cc_3374 ( N_noxref_9_c_4048_n N_noxref_11_c_4464_n ) capacitor c=6.53477e-19 \
 //x=34.78 //y=2.08 //x2=32.19 //y2=2.08
cc_3375 ( N_noxref_9_c_4151_p N_noxref_11_c_4464_n ) capacitor c=0.013297f \
 //x=32.15 //y=5.155 //x2=32.19 //y2=2.08
cc_3376 ( N_noxref_9_M103_noxref_g N_noxref_11_c_4479_n ) capacitor \
 c=0.0157304f //x=35.42 //y=6.02 //x2=35.995 //y2=5.155
cc_3377 ( N_noxref_9_c_4081_n N_noxref_11_c_4483_n ) capacitor c=3.10026e-19 \
 //x=32.845 //y=5.155 //x2=35.285 //y2=5.155
cc_3378 ( N_noxref_9_M102_noxref_g N_noxref_11_c_4483_n ) capacitor \
 c=0.0213876f //x=34.98 //y=6.02 //x2=35.285 //y2=5.155
cc_3379 ( N_noxref_9_c_4127_n N_noxref_11_c_4483_n ) capacitor c=0.00393496f \
 //x=35.345 //y=4.79 //x2=35.285 //y2=5.155
cc_3380 ( N_noxref_9_c_4044_n N_noxref_11_c_4493_n ) capacitor c=0.0165903f \
 //x=39.475 //y=2.59 //x2=37.74 //y2=3.33
cc_3381 ( N_noxref_9_c_4049_n N_noxref_11_c_4493_n ) capacitor c=0.0105286f \
 //x=39.59 //y=2.08 //x2=37.74 //y2=3.33
cc_3382 ( N_noxref_9_c_4077_n N_noxref_11_M100_noxref_g ) capacitor \
 c=0.0162556f //x=32.065 //y=5.155 //x2=31.93 //y2=6.02
cc_3383 ( N_noxref_9_M100_noxref_d N_noxref_11_M100_noxref_g ) capacitor \
 c=0.0180032f //x=32.005 //y=5.02 //x2=31.93 //y2=6.02
cc_3384 ( N_noxref_9_c_4081_n N_noxref_11_M101_noxref_g ) capacitor \
 c=0.0183937f //x=32.845 //y=5.155 //x2=32.37 //y2=6.02
cc_3385 ( N_noxref_9_M100_noxref_d N_noxref_11_M101_noxref_g ) capacitor \
 c=0.0194246f //x=32.005 //y=5.02 //x2=32.37 //y2=6.02
cc_3386 ( N_noxref_9_M20_noxref_d N_noxref_11_c_4559_n ) capacitor \
 c=0.00217566f //x=32.255 //y=0.915 //x2=32.18 //y2=0.915
cc_3387 ( N_noxref_9_M20_noxref_d N_noxref_11_c_4560_n ) capacitor \
 c=0.0034598f //x=32.255 //y=0.915 //x2=32.18 //y2=1.26
cc_3388 ( N_noxref_9_M20_noxref_d N_noxref_11_c_4561_n ) capacitor \
 c=0.00546784f //x=32.255 //y=0.915 //x2=32.18 //y2=1.57
cc_3389 ( N_noxref_9_M20_noxref_d N_noxref_11_c_4562_n ) capacitor \
 c=0.00241102f //x=32.255 //y=0.915 //x2=32.555 //y2=0.76
cc_3390 ( N_noxref_9_c_4046_n N_noxref_11_c_4563_n ) capacitor c=0.00371277f \
 //x=32.845 //y=1.665 //x2=32.555 //y2=1.415
cc_3391 ( N_noxref_9_M20_noxref_d N_noxref_11_c_4563_n ) capacitor \
 c=0.0138621f //x=32.255 //y=0.915 //x2=32.555 //y2=1.415
cc_3392 ( N_noxref_9_M20_noxref_d N_noxref_11_c_4565_n ) capacitor \
 c=0.00219619f //x=32.255 //y=0.915 //x2=32.71 //y2=0.915
cc_3393 ( N_noxref_9_c_4046_n N_noxref_11_c_4566_n ) capacitor c=0.00457401f \
 //x=32.845 //y=1.665 //x2=32.71 //y2=1.26
cc_3394 ( N_noxref_9_M20_noxref_d N_noxref_11_c_4566_n ) capacitor \
 c=0.00603828f //x=32.255 //y=0.915 //x2=32.71 //y2=1.26
cc_3395 ( N_noxref_9_c_4047_n N_noxref_11_c_4568_n ) capacitor c=0.00709342f \
 //x=32.93 //y=2.59 //x2=32.19 //y2=2.08
cc_3396 ( N_noxref_9_c_4047_n N_noxref_11_c_4569_n ) capacitor c=0.00283672f \
 //x=32.93 //y=2.59 //x2=32.19 //y2=1.915
cc_3397 ( N_noxref_9_M20_noxref_d N_noxref_11_c_4569_n ) capacitor \
 c=0.00661782f //x=32.255 //y=0.915 //x2=32.19 //y2=1.915
cc_3398 ( N_noxref_9_c_4081_n N_noxref_11_c_4532_n ) capacitor c=0.00201851f \
 //x=32.845 //y=5.155 //x2=32.19 //y2=4.7
cc_3399 ( N_noxref_9_c_4047_n N_noxref_11_c_4532_n ) capacitor c=0.0114782f \
 //x=32.93 //y=2.59 //x2=32.19 //y2=4.7
cc_3400 ( N_noxref_9_c_4151_p N_noxref_11_c_4532_n ) capacitor c=0.00470675f \
 //x=32.15 //y=5.155 //x2=32.19 //y2=4.7
cc_3401 ( N_noxref_9_M103_noxref_g N_noxref_11_M102_noxref_d ) capacitor \
 c=0.0180032f //x=35.42 //y=6.02 //x2=35.055 //y2=5.02
cc_3402 ( N_noxref_9_c_4049_n N_noxref_12_c_4809_n ) capacitor c=0.0197627f \
 //x=39.59 //y=2.08 //x2=41.695 //y2=3.7
cc_3403 ( N_noxref_9_c_4044_n N_noxref_12_c_4745_n ) capacitor c=0.0179628f \
 //x=39.475 //y=2.59 //x2=37 //y2=2.08
cc_3404 ( N_noxref_9_c_4048_n N_noxref_12_c_4745_n ) capacitor c=0.00108809f \
 //x=34.78 //y=2.08 //x2=37 //y2=2.08
cc_3405 ( N_noxref_9_c_4049_n N_noxref_12_c_4745_n ) capacitor c=6.20825e-19 \
 //x=39.59 //y=2.08 //x2=37 //y2=2.08
cc_3406 ( N_noxref_9_c_4049_n N_noxref_12_c_4746_n ) capacitor c=0.00106679f \
 //x=39.59 //y=2.08 //x2=41.81 //y2=2.08
cc_3407 ( N_noxref_9_c_4047_n N_D_c_5328_n ) capacitor c=0.0205387f //x=32.93 \
 //y=2.59 //x2=58.715 //y2=4.07
cc_3408 ( N_noxref_9_c_4048_n N_D_c_5328_n ) capacitor c=0.0218572f //x=34.78 \
 //y=2.08 //x2=58.715 //y2=4.07
cc_3409 ( N_noxref_9_c_4049_n N_D_c_5328_n ) capacitor c=0.0194977f //x=39.59 \
 //y=2.08 //x2=58.715 //y2=4.07
cc_3410 ( N_noxref_9_c_4075_n N_D_M96_noxref_g ) capacitor c=0.0213876f \
 //x=30.475 //y=5.155 //x2=30.17 //y2=6.02
cc_3411 ( N_noxref_9_c_4071_n N_D_M97_noxref_g ) capacitor c=0.0157304f \
 //x=31.185 //y=5.155 //x2=30.61 //y2=6.02
cc_3412 ( N_noxref_9_M96_noxref_d N_D_M97_noxref_g ) capacitor c=0.0180032f \
 //x=30.245 //y=5.02 //x2=30.61 //y2=6.02
cc_3413 ( N_noxref_9_c_4075_n N_D_c_5400_n ) capacitor c=0.00393496f \
 //x=30.475 //y=5.155 //x2=30.535 //y2=4.79
cc_3414 ( N_noxref_9_c_4047_n N_CLK_c_6058_n ) capacitor c=0.0166101f \
 //x=32.93 //y=2.59 //x2=35.775 //y2=4.44
cc_3415 ( N_noxref_9_c_4048_n N_CLK_c_6058_n ) capacitor c=0.018786f //x=34.78 \
 //y=2.08 //x2=35.775 //y2=4.44
cc_3416 ( N_noxref_9_c_4100_n N_CLK_c_6058_n ) capacitor c=0.0112124f \
 //x=35.055 //y=4.79 //x2=35.775 //y2=4.44
cc_3417 ( N_noxref_9_c_4049_n N_CLK_c_6068_n ) capacitor c=0.018786f //x=39.59 \
 //y=2.08 //x2=45.395 //y2=4.44
cc_3418 ( N_noxref_9_c_4102_n N_CLK_c_6068_n ) capacitor c=0.0112124f \
 //x=39.865 //y=4.79 //x2=45.395 //y2=4.44
cc_3419 ( N_noxref_9_c_4048_n N_CLK_c_6190_n ) capacitor c=0.00153281f \
 //x=34.78 //y=2.08 //x2=36.005 //y2=4.44
cc_3420 ( N_noxref_9_c_4044_n N_CLK_c_6042_n ) capacitor c=0.0190006f \
 //x=39.475 //y=2.59 //x2=35.89 //y2=2.08
cc_3421 ( N_noxref_9_c_4045_n N_CLK_c_6042_n ) capacitor c=9.95819e-19 \
 //x=34.895 //y=2.59 //x2=35.89 //y2=2.08
cc_3422 ( N_noxref_9_c_4047_n N_CLK_c_6042_n ) capacitor c=3.63796e-19 \
 //x=32.93 //y=2.59 //x2=35.89 //y2=2.08
cc_3423 ( N_noxref_9_c_4048_n N_CLK_c_6042_n ) capacitor c=0.0416208f \
 //x=34.78 //y=2.08 //x2=35.89 //y2=2.08
cc_3424 ( N_noxref_9_c_4054_n N_CLK_c_6042_n ) capacitor c=0.00210802f \
 //x=34.48 //y=1.915 //x2=35.89 //y2=2.08
cc_3425 ( N_noxref_9_c_4127_n N_CLK_c_6042_n ) capacitor c=0.00120758f \
 //x=35.345 //y=4.79 //x2=35.89 //y2=2.08
cc_3426 ( N_noxref_9_c_4100_n N_CLK_c_6042_n ) capacitor c=0.00141297f \
 //x=35.055 //y=4.79 //x2=35.89 //y2=2.08
cc_3427 ( N_noxref_9_M102_noxref_g N_CLK_M104_noxref_g ) capacitor \
 c=0.0105174f //x=34.98 //y=6.02 //x2=35.86 //y2=6.02
cc_3428 ( N_noxref_9_M103_noxref_g N_CLK_M104_noxref_g ) capacitor c=0.10624f \
 //x=35.42 //y=6.02 //x2=35.86 //y2=6.02
cc_3429 ( N_noxref_9_M103_noxref_g N_CLK_M105_noxref_g ) capacitor \
 c=0.0100903f //x=35.42 //y=6.02 //x2=36.3 //y2=6.02
cc_3430 ( N_noxref_9_c_4050_n N_CLK_c_6285_n ) capacitor c=5.72482e-19 \
 //x=34.48 //y=0.875 //x2=35.455 //y2=0.91
cc_3431 ( N_noxref_9_c_4052_n N_CLK_c_6285_n ) capacitor c=0.00149976f \
 //x=34.48 //y=1.22 //x2=35.455 //y2=0.91
cc_3432 ( N_noxref_9_c_4057_n N_CLK_c_6285_n ) capacitor c=0.0160123f \
 //x=35.01 //y=0.875 //x2=35.455 //y2=0.91
cc_3433 ( N_noxref_9_c_4053_n N_CLK_c_6288_n ) capacitor c=0.00111227f \
 //x=34.48 //y=1.53 //x2=35.455 //y2=1.22
cc_3434 ( N_noxref_9_c_4059_n N_CLK_c_6288_n ) capacitor c=0.0124075f \
 //x=35.01 //y=1.22 //x2=35.455 //y2=1.22
cc_3435 ( N_noxref_9_c_4057_n N_CLK_c_6290_n ) capacitor c=0.00103227f \
 //x=35.01 //y=0.875 //x2=35.98 //y2=0.91
cc_3436 ( N_noxref_9_c_4059_n N_CLK_c_6291_n ) capacitor c=0.0010154f \
 //x=35.01 //y=1.22 //x2=35.98 //y2=1.22
cc_3437 ( N_noxref_9_c_4059_n N_CLK_c_6292_n ) capacitor c=9.23422e-19 \
 //x=35.01 //y=1.22 //x2=35.98 //y2=1.45
cc_3438 ( N_noxref_9_c_4048_n N_CLK_c_6293_n ) capacitor c=0.00203769f \
 //x=34.78 //y=2.08 //x2=35.98 //y2=1.915
cc_3439 ( N_noxref_9_c_4054_n N_CLK_c_6293_n ) capacitor c=0.00834532f \
 //x=34.48 //y=1.915 //x2=35.98 //y2=1.915
cc_3440 ( N_noxref_9_c_4048_n N_CLK_c_6215_n ) capacitor c=0.0017365f \
 //x=34.78 //y=2.08 //x2=35.89 //y2=4.7
cc_3441 ( N_noxref_9_c_4127_n N_CLK_c_6215_n ) capacitor c=0.0170104f \
 //x=35.345 //y=4.79 //x2=35.89 //y2=4.7
cc_3442 ( N_noxref_9_c_4100_n N_CLK_c_6215_n ) capacitor c=0.00484466f \
 //x=35.055 //y=4.79 //x2=35.89 //y2=4.7
cc_3443 ( N_noxref_9_c_4042_n N_RN_c_7046_n ) capacitor c=0.143487f //x=34.665 \
 //y=2.59 //x2=46.505 //y2=2.22
cc_3444 ( N_noxref_9_c_4043_n N_RN_c_7046_n ) capacitor c=0.0291301f \
 //x=33.045 //y=2.59 //x2=46.505 //y2=2.22
cc_3445 ( N_noxref_9_c_4044_n N_RN_c_7046_n ) capacitor c=0.42762f //x=39.475 \
 //y=2.59 //x2=46.505 //y2=2.22
cc_3446 ( N_noxref_9_c_4045_n N_RN_c_7046_n ) capacitor c=0.0264401f \
 //x=34.895 //y=2.59 //x2=46.505 //y2=2.22
cc_3447 ( N_noxref_9_c_4223_p N_RN_c_7046_n ) capacitor c=0.016327f //x=32.53 \
 //y=1.665 //x2=46.505 //y2=2.22
cc_3448 ( N_noxref_9_c_4047_n N_RN_c_7046_n ) capacitor c=0.0215653f //x=32.93 \
 //y=2.59 //x2=46.505 //y2=2.22
cc_3449 ( N_noxref_9_c_4048_n N_RN_c_7046_n ) capacitor c=0.021104f //x=34.78 \
 //y=2.08 //x2=46.505 //y2=2.22
cc_3450 ( N_noxref_9_c_4049_n N_RN_c_7046_n ) capacitor c=0.021104f //x=39.59 \
 //y=2.08 //x2=46.505 //y2=2.22
cc_3451 ( N_noxref_9_c_4054_n N_RN_c_7046_n ) capacitor c=0.011987f //x=34.48 \
 //y=1.915 //x2=46.505 //y2=2.22
cc_3452 ( N_noxref_9_c_4064_n N_RN_c_7046_n ) capacitor c=0.011987f //x=39.29 \
 //y=1.915 //x2=46.505 //y2=2.22
cc_3453 ( N_noxref_9_c_4071_n N_RN_c_7091_n ) capacitor c=0.0120276f \
 //x=31.185 //y=5.155 //x2=31.08 //y2=2.08
cc_3454 ( N_noxref_9_c_4047_n N_RN_c_7091_n ) capacitor c=0.00254659f \
 //x=32.93 //y=2.59 //x2=31.08 //y2=2.08
cc_3455 ( N_noxref_9_c_4071_n N_RN_M98_noxref_g ) capacitor c=0.0163793f \
 //x=31.185 //y=5.155 //x2=31.05 //y2=6.02
cc_3456 ( N_noxref_9_M98_noxref_d N_RN_M98_noxref_g ) capacitor c=0.0180032f \
 //x=31.125 //y=5.02 //x2=31.05 //y2=6.02
cc_3457 ( N_noxref_9_c_4077_n N_RN_M99_noxref_g ) capacitor c=0.0162556f \
 //x=32.065 //y=5.155 //x2=31.49 //y2=6.02
cc_3458 ( N_noxref_9_M98_noxref_d N_RN_M99_noxref_g ) capacitor c=0.0180032f \
 //x=31.125 //y=5.02 //x2=31.49 //y2=6.02
cc_3459 ( N_noxref_9_c_4235_p N_RN_c_7256_n ) capacitor c=0.00392095f \
 //x=31.27 //y=5.155 //x2=31.415 //y2=4.79
cc_3460 ( N_noxref_9_c_4071_n N_RN_c_7261_n ) capacitor c=0.00309994f \
 //x=31.185 //y=5.155 //x2=31.08 //y2=4.7
cc_3461 ( N_noxref_9_c_4042_n N_SN_c_8132_n ) capacitor c=0.143324f //x=34.665 \
 //y=2.59 //x2=40.585 //y2=2.96
cc_3462 ( N_noxref_9_c_4043_n N_SN_c_8132_n ) capacitor c=0.0293832f \
 //x=33.045 //y=2.59 //x2=40.585 //y2=2.96
cc_3463 ( N_noxref_9_c_4044_n N_SN_c_8132_n ) capacitor c=0.429547f //x=39.475 \
 //y=2.59 //x2=40.585 //y2=2.96
cc_3464 ( N_noxref_9_c_4045_n N_SN_c_8132_n ) capacitor c=0.0267736f \
 //x=34.895 //y=2.59 //x2=40.585 //y2=2.96
cc_3465 ( N_noxref_9_c_4047_n N_SN_c_8132_n ) capacitor c=0.0206007f //x=32.93 \
 //y=2.59 //x2=40.585 //y2=2.96
cc_3466 ( N_noxref_9_c_4048_n N_SN_c_8132_n ) capacitor c=0.0216195f //x=34.78 \
 //y=2.08 //x2=40.585 //y2=2.96
cc_3467 ( N_noxref_9_c_4049_n N_SN_c_8132_n ) capacitor c=0.0215933f //x=39.59 \
 //y=2.08 //x2=40.585 //y2=2.96
cc_3468 ( N_noxref_9_c_4049_n N_SN_c_8340_n ) capacitor c=0.00128547f \
 //x=39.59 //y=2.08 //x2=40.815 //y2=2.96
cc_3469 ( N_noxref_9_c_4044_n N_SN_c_8147_n ) capacitor c=0.00311593f \
 //x=39.475 //y=2.59 //x2=40.7 //y2=2.08
cc_3470 ( N_noxref_9_c_4049_n N_SN_c_8147_n ) capacitor c=0.0408822f //x=39.59 \
 //y=2.08 //x2=40.7 //y2=2.08
cc_3471 ( N_noxref_9_c_4064_n N_SN_c_8147_n ) capacitor c=0.00210802f \
 //x=39.29 //y=1.915 //x2=40.7 //y2=2.08
cc_3472 ( N_noxref_9_c_4129_n N_SN_c_8147_n ) capacitor c=0.00120758f \
 //x=40.155 //y=4.79 //x2=40.7 //y2=2.08
cc_3473 ( N_noxref_9_c_4102_n N_SN_c_8147_n ) capacitor c=0.00142741f \
 //x=39.865 //y=4.79 //x2=40.7 //y2=2.08
cc_3474 ( N_noxref_9_M108_noxref_g N_SN_M110_noxref_g ) capacitor c=0.0105174f \
 //x=39.79 //y=6.02 //x2=40.67 //y2=6.02
cc_3475 ( N_noxref_9_M109_noxref_g N_SN_M110_noxref_g ) capacitor c=0.10624f \
 //x=40.23 //y=6.02 //x2=40.67 //y2=6.02
cc_3476 ( N_noxref_9_M109_noxref_g N_SN_M111_noxref_g ) capacitor c=0.0100903f \
 //x=40.23 //y=6.02 //x2=41.11 //y2=6.02
cc_3477 ( N_noxref_9_c_4060_n N_SN_c_8349_n ) capacitor c=5.72482e-19 \
 //x=39.29 //y=0.875 //x2=40.265 //y2=0.91
cc_3478 ( N_noxref_9_c_4062_n N_SN_c_8349_n ) capacitor c=0.00149976f \
 //x=39.29 //y=1.22 //x2=40.265 //y2=0.91
cc_3479 ( N_noxref_9_c_4067_n N_SN_c_8349_n ) capacitor c=0.0160123f //x=39.82 \
 //y=0.875 //x2=40.265 //y2=0.91
cc_3480 ( N_noxref_9_c_4063_n N_SN_c_8352_n ) capacitor c=0.00111227f \
 //x=39.29 //y=1.53 //x2=40.265 //y2=1.22
cc_3481 ( N_noxref_9_c_4069_n N_SN_c_8352_n ) capacitor c=0.0124075f //x=39.82 \
 //y=1.22 //x2=40.265 //y2=1.22
cc_3482 ( N_noxref_9_c_4067_n N_SN_c_8354_n ) capacitor c=0.00103227f \
 //x=39.82 //y=0.875 //x2=40.79 //y2=0.91
cc_3483 ( N_noxref_9_c_4069_n N_SN_c_8355_n ) capacitor c=0.0010154f //x=39.82 \
 //y=1.22 //x2=40.79 //y2=1.22
cc_3484 ( N_noxref_9_c_4069_n N_SN_c_8356_n ) capacitor c=9.23422e-19 \
 //x=39.82 //y=1.22 //x2=40.79 //y2=1.45
cc_3485 ( N_noxref_9_c_4049_n N_SN_c_8357_n ) capacitor c=0.00203769f \
 //x=39.59 //y=2.08 //x2=40.79 //y2=1.915
cc_3486 ( N_noxref_9_c_4064_n N_SN_c_8357_n ) capacitor c=0.00834532f \
 //x=39.29 //y=1.915 //x2=40.79 //y2=1.915
cc_3487 ( N_noxref_9_c_4049_n N_SN_c_8268_n ) capacitor c=0.0017365f //x=39.59 \
 //y=2.08 //x2=40.7 //y2=4.7
cc_3488 ( N_noxref_9_c_4129_n N_SN_c_8268_n ) capacitor c=0.0170104f \
 //x=40.155 //y=4.79 //x2=40.7 //y2=4.7
cc_3489 ( N_noxref_9_c_4102_n N_SN_c_8268_n ) capacitor c=0.00484466f \
 //x=39.865 //y=4.79 //x2=40.7 //y2=4.7
cc_3490 ( N_noxref_9_M20_noxref_d N_noxref_40_M18_noxref_s ) capacitor \
 c=0.00309936f //x=32.255 //y=0.915 //x2=29.315 //y2=0.375
cc_3491 ( N_noxref_9_c_4046_n N_noxref_41_c_11209_n ) capacitor c=0.00457167f \
 //x=32.845 //y=1.665 //x2=32.845 //y2=0.54
cc_3492 ( N_noxref_9_M20_noxref_d N_noxref_41_c_11209_n ) capacitor \
 c=0.0115903f //x=32.255 //y=0.915 //x2=32.845 //y2=0.54
cc_3493 ( N_noxref_9_c_4223_p N_noxref_41_c_11219_n ) capacitor c=0.0200405f \
 //x=32.53 //y=1.665 //x2=31.96 //y2=0.995
cc_3494 ( N_noxref_9_M20_noxref_d N_noxref_41_M19_noxref_d ) capacitor \
 c=5.27807e-19 //x=32.255 //y=0.915 //x2=30.72 //y2=0.91
cc_3495 ( N_noxref_9_c_4046_n N_noxref_41_M20_noxref_s ) capacitor \
 c=0.0184051f //x=32.845 //y=1.665 //x2=31.825 //y2=0.375
cc_3496 ( N_noxref_9_M20_noxref_d N_noxref_41_M20_noxref_s ) capacitor \
 c=0.0426368f //x=32.255 //y=0.915 //x2=31.825 //y2=0.375
cc_3497 ( N_noxref_9_c_4046_n N_noxref_42_c_11271_n ) capacitor c=3.84569e-19 \
 //x=32.845 //y=1.665 //x2=34.26 //y2=1.505
cc_3498 ( N_noxref_9_c_4054_n N_noxref_42_c_11271_n ) capacitor c=0.0034165f \
 //x=34.48 //y=1.915 //x2=34.26 //y2=1.505
cc_3499 ( N_noxref_9_c_4048_n N_noxref_42_c_11256_n ) capacitor c=0.0115578f \
 //x=34.78 //y=2.08 //x2=35.145 //y2=1.59
cc_3500 ( N_noxref_9_c_4053_n N_noxref_42_c_11256_n ) capacitor c=0.00697148f \
 //x=34.48 //y=1.53 //x2=35.145 //y2=1.59
cc_3501 ( N_noxref_9_c_4054_n N_noxref_42_c_11256_n ) capacitor c=0.0204849f \
 //x=34.48 //y=1.915 //x2=35.145 //y2=1.59
cc_3502 ( N_noxref_9_c_4056_n N_noxref_42_c_11256_n ) capacitor c=0.00610316f \
 //x=34.855 //y=1.375 //x2=35.145 //y2=1.59
cc_3503 ( N_noxref_9_c_4059_n N_noxref_42_c_11256_n ) capacitor c=0.00698822f \
 //x=35.01 //y=1.22 //x2=35.145 //y2=1.59
cc_3504 ( N_noxref_9_c_4050_n N_noxref_42_M21_noxref_s ) capacitor \
 c=0.0327271f //x=34.48 //y=0.875 //x2=34.125 //y2=0.375
cc_3505 ( N_noxref_9_c_4053_n N_noxref_42_M21_noxref_s ) capacitor \
 c=7.99997e-19 //x=34.48 //y=1.53 //x2=34.125 //y2=0.375
cc_3506 ( N_noxref_9_c_4054_n N_noxref_42_M21_noxref_s ) capacitor \
 c=0.00122123f //x=34.48 //y=1.915 //x2=34.125 //y2=0.375
cc_3507 ( N_noxref_9_c_4057_n N_noxref_42_M21_noxref_s ) capacitor \
 c=0.0121427f //x=35.01 //y=0.875 //x2=34.125 //y2=0.375
cc_3508 ( N_noxref_9_M20_noxref_d N_noxref_42_M21_noxref_s ) capacitor \
 c=2.55333e-19 //x=32.255 //y=0.915 //x2=34.125 //y2=0.375
cc_3509 ( N_noxref_9_c_4064_n N_noxref_44_c_11372_n ) capacitor c=0.0034165f \
 //x=39.29 //y=1.915 //x2=39.07 //y2=1.505
cc_3510 ( N_noxref_9_c_4049_n N_noxref_44_c_11357_n ) capacitor c=0.0115578f \
 //x=39.59 //y=2.08 //x2=39.955 //y2=1.59
cc_3511 ( N_noxref_9_c_4063_n N_noxref_44_c_11357_n ) capacitor c=0.00697148f \
 //x=39.29 //y=1.53 //x2=39.955 //y2=1.59
cc_3512 ( N_noxref_9_c_4064_n N_noxref_44_c_11357_n ) capacitor c=0.0204849f \
 //x=39.29 //y=1.915 //x2=39.955 //y2=1.59
cc_3513 ( N_noxref_9_c_4066_n N_noxref_44_c_11357_n ) capacitor c=0.00610316f \
 //x=39.665 //y=1.375 //x2=39.955 //y2=1.59
cc_3514 ( N_noxref_9_c_4069_n N_noxref_44_c_11357_n ) capacitor c=0.00698822f \
 //x=39.82 //y=1.22 //x2=39.955 //y2=1.59
cc_3515 ( N_noxref_9_c_4060_n N_noxref_44_M24_noxref_s ) capacitor \
 c=0.0327271f //x=39.29 //y=0.875 //x2=38.935 //y2=0.375
cc_3516 ( N_noxref_9_c_4063_n N_noxref_44_M24_noxref_s ) capacitor \
 c=7.99997e-19 //x=39.29 //y=1.53 //x2=38.935 //y2=0.375
cc_3517 ( N_noxref_9_c_4064_n N_noxref_44_M24_noxref_s ) capacitor \
 c=0.00122123f //x=39.29 //y=1.915 //x2=38.935 //y2=0.375
cc_3518 ( N_noxref_9_c_4067_n N_noxref_44_M24_noxref_s ) capacitor \
 c=0.0121427f //x=39.82 //y=0.875 //x2=38.935 //y2=0.375
cc_3519 ( N_noxref_10_c_4295_n N_noxref_11_c_4541_n ) capacitor c=0.0119023f \
 //x=44.285 //y=2.59 //x2=49.095 //y2=3.33
cc_3520 ( N_noxref_10_c_4296_n N_noxref_11_c_4541_n ) capacitor c=8.87672e-19 \
 //x=42.665 //y=2.59 //x2=49.095 //y2=3.33
cc_3521 ( N_noxref_10_c_4298_n N_noxref_11_c_4541_n ) capacitor c=0.018769f \
 //x=42.55 //y=2.59 //x2=49.095 //y2=3.33
cc_3522 ( N_noxref_10_c_4299_n N_noxref_11_c_4541_n ) capacitor c=0.0198064f \
 //x=44.4 //y=2.08 //x2=49.095 //y2=3.33
cc_3523 ( N_noxref_10_c_4315_n N_noxref_11_c_4489_n ) capacitor c=3.10026e-19 \
 //x=40.095 //y=5.155 //x2=37.655 //y2=5.155
cc_3524 ( N_noxref_10_c_4298_n N_noxref_12_c_4814_n ) capacitor c=0.0187698f \
 //x=42.55 //y=2.59 //x2=47.245 //y2=3.7
cc_3525 ( N_noxref_10_c_4299_n N_noxref_12_c_4814_n ) capacitor c=0.0197889f \
 //x=44.4 //y=2.08 //x2=47.245 //y2=3.7
cc_3526 ( N_noxref_10_c_4298_n N_noxref_12_c_4816_n ) capacitor c=0.00179385f \
 //x=42.55 //y=2.59 //x2=41.925 //y2=3.7
cc_3527 ( N_noxref_10_c_4296_n N_noxref_12_c_4746_n ) capacitor c=0.00456439f \
 //x=42.665 //y=2.59 //x2=41.81 //y2=2.08
cc_3528 ( N_noxref_10_c_4298_n N_noxref_12_c_4746_n ) capacitor c=0.0750956f \
 //x=42.55 //y=2.59 //x2=41.81 //y2=2.08
cc_3529 ( N_noxref_10_c_4299_n N_noxref_12_c_4746_n ) capacitor c=5.32619e-19 \
 //x=44.4 //y=2.08 //x2=41.81 //y2=2.08
cc_3530 ( N_noxref_10_c_4373_p N_noxref_12_c_4746_n ) capacitor c=0.0126839f \
 //x=41.77 //y=5.155 //x2=41.81 //y2=2.08
cc_3531 ( N_noxref_10_M115_noxref_g N_noxref_12_c_4752_n ) capacitor \
 c=0.0157304f //x=45.04 //y=6.02 //x2=45.615 //y2=5.155
cc_3532 ( N_noxref_10_c_4321_n N_noxref_12_c_4756_n ) capacitor c=3.10026e-19 \
 //x=42.465 //y=5.155 //x2=44.905 //y2=5.155
cc_3533 ( N_noxref_10_M114_noxref_g N_noxref_12_c_4756_n ) capacitor \
 c=0.0213876f //x=44.6 //y=6.02 //x2=44.905 //y2=5.155
cc_3534 ( N_noxref_10_c_4355_n N_noxref_12_c_4756_n ) capacitor c=0.00393496f \
 //x=44.965 //y=4.79 //x2=44.905 //y2=5.155
cc_3535 ( N_noxref_10_c_4317_n N_noxref_12_M112_noxref_g ) capacitor \
 c=0.0162556f //x=41.685 //y=5.155 //x2=41.55 //y2=6.02
cc_3536 ( N_noxref_10_M112_noxref_d N_noxref_12_M112_noxref_g ) capacitor \
 c=0.0180032f //x=41.625 //y=5.02 //x2=41.55 //y2=6.02
cc_3537 ( N_noxref_10_c_4321_n N_noxref_12_M113_noxref_g ) capacitor \
 c=0.0183937f //x=42.465 //y=5.155 //x2=41.99 //y2=6.02
cc_3538 ( N_noxref_10_M112_noxref_d N_noxref_12_M113_noxref_g ) capacitor \
 c=0.0194246f //x=41.625 //y=5.02 //x2=41.99 //y2=6.02
cc_3539 ( N_noxref_10_M26_noxref_d N_noxref_12_c_4829_n ) capacitor \
 c=0.00217566f //x=41.875 //y=0.915 //x2=41.8 //y2=0.915
cc_3540 ( N_noxref_10_M26_noxref_d N_noxref_12_c_4830_n ) capacitor \
 c=0.0034598f //x=41.875 //y=0.915 //x2=41.8 //y2=1.26
cc_3541 ( N_noxref_10_M26_noxref_d N_noxref_12_c_4831_n ) capacitor \
 c=0.00546784f //x=41.875 //y=0.915 //x2=41.8 //y2=1.57
cc_3542 ( N_noxref_10_M26_noxref_d N_noxref_12_c_4832_n ) capacitor \
 c=0.00241102f //x=41.875 //y=0.915 //x2=42.175 //y2=0.76
cc_3543 ( N_noxref_10_c_4297_n N_noxref_12_c_4833_n ) capacitor c=0.00371277f \
 //x=42.465 //y=1.665 //x2=42.175 //y2=1.415
cc_3544 ( N_noxref_10_M26_noxref_d N_noxref_12_c_4833_n ) capacitor \
 c=0.0138621f //x=41.875 //y=0.915 //x2=42.175 //y2=1.415
cc_3545 ( N_noxref_10_M26_noxref_d N_noxref_12_c_4835_n ) capacitor \
 c=0.00219619f //x=41.875 //y=0.915 //x2=42.33 //y2=0.915
cc_3546 ( N_noxref_10_c_4297_n N_noxref_12_c_4836_n ) capacitor c=0.00457401f \
 //x=42.465 //y=1.665 //x2=42.33 //y2=1.26
cc_3547 ( N_noxref_10_M26_noxref_d N_noxref_12_c_4836_n ) capacitor \
 c=0.00603828f //x=41.875 //y=0.915 //x2=42.33 //y2=1.26
cc_3548 ( N_noxref_10_c_4298_n N_noxref_12_c_4838_n ) capacitor c=0.00731987f \
 //x=42.55 //y=2.59 //x2=41.81 //y2=2.08
cc_3549 ( N_noxref_10_c_4298_n N_noxref_12_c_4839_n ) capacitor c=0.00283672f \
 //x=42.55 //y=2.59 //x2=41.81 //y2=1.915
cc_3550 ( N_noxref_10_M26_noxref_d N_noxref_12_c_4839_n ) capacitor \
 c=0.00661782f //x=41.875 //y=0.915 //x2=41.81 //y2=1.915
cc_3551 ( N_noxref_10_c_4321_n N_noxref_12_c_4807_n ) capacitor c=0.00201851f \
 //x=42.465 //y=5.155 //x2=41.81 //y2=4.7
cc_3552 ( N_noxref_10_c_4298_n N_noxref_12_c_4807_n ) capacitor c=0.0114782f \
 //x=42.55 //y=2.59 //x2=41.81 //y2=4.7
cc_3553 ( N_noxref_10_c_4373_p N_noxref_12_c_4807_n ) capacitor c=0.00470675f \
 //x=41.77 //y=5.155 //x2=41.81 //y2=4.7
cc_3554 ( N_noxref_10_M115_noxref_g N_noxref_12_M114_noxref_d ) capacitor \
 c=0.0180032f //x=45.04 //y=6.02 //x2=44.675 //y2=5.02
cc_3555 ( N_noxref_10_c_4298_n N_D_c_5328_n ) capacitor c=0.0181982f //x=42.55 \
 //y=2.59 //x2=58.715 //y2=4.07
cc_3556 ( N_noxref_10_c_4299_n N_D_c_5328_n ) capacitor c=0.019517f //x=44.4 \
 //y=2.08 //x2=58.715 //y2=4.07
cc_3557 ( N_noxref_10_c_4298_n N_CLK_c_6068_n ) capacitor c=0.0166101f \
 //x=42.55 //y=2.59 //x2=45.395 //y2=4.44
cc_3558 ( N_noxref_10_c_4299_n N_CLK_c_6068_n ) capacitor c=0.018786f //x=44.4 \
 //y=2.08 //x2=45.395 //y2=4.44
cc_3559 ( N_noxref_10_c_4333_n N_CLK_c_6068_n ) capacitor c=0.0112124f \
 //x=44.675 //y=4.79 //x2=45.395 //y2=4.44
cc_3560 ( N_noxref_10_c_4299_n N_CLK_c_6192_n ) capacitor c=0.00153281f \
 //x=44.4 //y=2.08 //x2=45.625 //y2=4.44
cc_3561 ( N_noxref_10_c_4295_n N_CLK_c_6043_n ) capacitor c=0.00520283f \
 //x=44.285 //y=2.59 //x2=45.51 //y2=2.08
cc_3562 ( N_noxref_10_c_4298_n N_CLK_c_6043_n ) capacitor c=2.96936e-19 \
 //x=42.55 //y=2.59 //x2=45.51 //y2=2.08
cc_3563 ( N_noxref_10_c_4299_n N_CLK_c_6043_n ) capacitor c=0.0403217f \
 //x=44.4 //y=2.08 //x2=45.51 //y2=2.08
cc_3564 ( N_noxref_10_c_4304_n N_CLK_c_6043_n ) capacitor c=0.00210802f \
 //x=44.1 //y=1.915 //x2=45.51 //y2=2.08
cc_3565 ( N_noxref_10_c_4355_n N_CLK_c_6043_n ) capacitor c=0.00120758f \
 //x=44.965 //y=4.79 //x2=45.51 //y2=2.08
cc_3566 ( N_noxref_10_c_4333_n N_CLK_c_6043_n ) capacitor c=0.00141297f \
 //x=44.675 //y=4.79 //x2=45.51 //y2=2.08
cc_3567 ( N_noxref_10_M114_noxref_g N_CLK_M116_noxref_g ) capacitor \
 c=0.0105174f //x=44.6 //y=6.02 //x2=45.48 //y2=6.02
cc_3568 ( N_noxref_10_M115_noxref_g N_CLK_M116_noxref_g ) capacitor c=0.10624f \
 //x=45.04 //y=6.02 //x2=45.48 //y2=6.02
cc_3569 ( N_noxref_10_M115_noxref_g N_CLK_M117_noxref_g ) capacitor \
 c=0.0100903f //x=45.04 //y=6.02 //x2=45.92 //y2=6.02
cc_3570 ( N_noxref_10_c_4300_n N_CLK_c_6311_n ) capacitor c=5.72482e-19 \
 //x=44.1 //y=0.875 //x2=45.075 //y2=0.91
cc_3571 ( N_noxref_10_c_4302_n N_CLK_c_6311_n ) capacitor c=0.00149976f \
 //x=44.1 //y=1.22 //x2=45.075 //y2=0.91
cc_3572 ( N_noxref_10_c_4307_n N_CLK_c_6311_n ) capacitor c=0.0160123f \
 //x=44.63 //y=0.875 //x2=45.075 //y2=0.91
cc_3573 ( N_noxref_10_c_4303_n N_CLK_c_6314_n ) capacitor c=0.00111227f \
 //x=44.1 //y=1.53 //x2=45.075 //y2=1.22
cc_3574 ( N_noxref_10_c_4309_n N_CLK_c_6314_n ) capacitor c=0.0124075f \
 //x=44.63 //y=1.22 //x2=45.075 //y2=1.22
cc_3575 ( N_noxref_10_c_4307_n N_CLK_c_6316_n ) capacitor c=0.00103227f \
 //x=44.63 //y=0.875 //x2=45.6 //y2=0.91
cc_3576 ( N_noxref_10_c_4309_n N_CLK_c_6317_n ) capacitor c=0.0010154f \
 //x=44.63 //y=1.22 //x2=45.6 //y2=1.22
cc_3577 ( N_noxref_10_c_4309_n N_CLK_c_6318_n ) capacitor c=9.23422e-19 \
 //x=44.63 //y=1.22 //x2=45.6 //y2=1.45
cc_3578 ( N_noxref_10_c_4299_n N_CLK_c_6319_n ) capacitor c=0.00203769f \
 //x=44.4 //y=2.08 //x2=45.6 //y2=1.915
cc_3579 ( N_noxref_10_c_4304_n N_CLK_c_6319_n ) capacitor c=0.00834532f \
 //x=44.1 //y=1.915 //x2=45.6 //y2=1.915
cc_3580 ( N_noxref_10_c_4299_n N_CLK_c_6216_n ) capacitor c=0.0017365f \
 //x=44.4 //y=2.08 //x2=45.51 //y2=4.7
cc_3581 ( N_noxref_10_c_4355_n N_CLK_c_6216_n ) capacitor c=0.0170104f \
 //x=44.965 //y=4.79 //x2=45.51 //y2=4.7
cc_3582 ( N_noxref_10_c_4333_n N_CLK_c_6216_n ) capacitor c=0.00484466f \
 //x=44.675 //y=4.79 //x2=45.51 //y2=4.7
cc_3583 ( N_noxref_10_c_4295_n N_RN_c_7046_n ) capacitor c=0.172592f \
 //x=44.285 //y=2.59 //x2=46.505 //y2=2.22
cc_3584 ( N_noxref_10_c_4296_n N_RN_c_7046_n ) capacitor c=0.0291301f \
 //x=42.665 //y=2.59 //x2=46.505 //y2=2.22
cc_3585 ( N_noxref_10_c_4428_p N_RN_c_7046_n ) capacitor c=0.016327f //x=42.15 \
 //y=1.665 //x2=46.505 //y2=2.22
cc_3586 ( N_noxref_10_c_4298_n N_RN_c_7046_n ) capacitor c=0.0215653f \
 //x=42.55 //y=2.59 //x2=46.505 //y2=2.22
cc_3587 ( N_noxref_10_c_4299_n N_RN_c_7046_n ) capacitor c=0.021104f //x=44.4 \
 //y=2.08 //x2=46.505 //y2=2.22
cc_3588 ( N_noxref_10_c_4304_n N_RN_c_7046_n ) capacitor c=0.011987f //x=44.1 \
 //y=1.915 //x2=46.505 //y2=2.22
cc_3589 ( N_noxref_10_c_4299_n N_RN_c_7092_n ) capacitor c=0.00107158f \
 //x=44.4 //y=2.08 //x2=46.62 //y2=2.08
cc_3590 ( N_noxref_10_c_4295_n N_SN_c_8135_n ) capacitor c=0.172781f \
 //x=44.285 //y=2.59 //x2=55.015 //y2=2.96
cc_3591 ( N_noxref_10_c_4296_n N_SN_c_8135_n ) capacitor c=0.0293832f \
 //x=42.665 //y=2.59 //x2=55.015 //y2=2.96
cc_3592 ( N_noxref_10_c_4298_n N_SN_c_8135_n ) capacitor c=0.0206007f \
 //x=42.55 //y=2.59 //x2=55.015 //y2=2.96
cc_3593 ( N_noxref_10_c_4299_n N_SN_c_8135_n ) capacitor c=0.0216195f //x=44.4 \
 //y=2.08 //x2=55.015 //y2=2.96
cc_3594 ( N_noxref_10_c_4311_n N_SN_c_8147_n ) capacitor c=0.0121898f \
 //x=40.805 //y=5.155 //x2=40.7 //y2=2.08
cc_3595 ( N_noxref_10_c_4298_n N_SN_c_8147_n ) capacitor c=0.00216737f \
 //x=42.55 //y=2.59 //x2=40.7 //y2=2.08
cc_3596 ( N_noxref_10_c_4311_n N_SN_M110_noxref_g ) capacitor c=0.0163793f \
 //x=40.805 //y=5.155 //x2=40.67 //y2=6.02
cc_3597 ( N_noxref_10_M110_noxref_d N_SN_M110_noxref_g ) capacitor \
 c=0.0180032f //x=40.745 //y=5.02 //x2=40.67 //y2=6.02
cc_3598 ( N_noxref_10_c_4317_n N_SN_M111_noxref_g ) capacitor c=0.0162556f \
 //x=41.685 //y=5.155 //x2=41.11 //y2=6.02
cc_3599 ( N_noxref_10_M110_noxref_d N_SN_M111_noxref_g ) capacitor \
 c=0.0180032f //x=40.745 //y=5.02 //x2=41.11 //y2=6.02
cc_3600 ( N_noxref_10_c_4443_p N_SN_c_8260_n ) capacitor c=0.00392095f \
 //x=40.89 //y=5.155 //x2=41.035 //y2=4.79
cc_3601 ( N_noxref_10_c_4311_n N_SN_c_8268_n ) capacitor c=0.00309994f \
 //x=40.805 //y=5.155 //x2=40.7 //y2=4.7
cc_3602 ( N_noxref_10_M26_noxref_d N_noxref_44_M24_noxref_s ) capacitor \
 c=0.00309936f //x=41.875 //y=0.915 //x2=38.935 //y2=0.375
cc_3603 ( N_noxref_10_c_4297_n N_noxref_45_c_11411_n ) capacitor c=0.00457167f \
 //x=42.465 //y=1.665 //x2=42.465 //y2=0.54
cc_3604 ( N_noxref_10_M26_noxref_d N_noxref_45_c_11411_n ) capacitor \
 c=0.0115903f //x=41.875 //y=0.915 //x2=42.465 //y2=0.54
cc_3605 ( N_noxref_10_c_4428_p N_noxref_45_c_11421_n ) capacitor c=0.0200405f \
 //x=42.15 //y=1.665 //x2=41.58 //y2=0.995
cc_3606 ( N_noxref_10_M26_noxref_d N_noxref_45_M25_noxref_d ) capacitor \
 c=5.27807e-19 //x=41.875 //y=0.915 //x2=40.34 //y2=0.91
cc_3607 ( N_noxref_10_c_4297_n N_noxref_45_M26_noxref_s ) capacitor \
 c=0.0184051f //x=42.465 //y=1.665 //x2=41.445 //y2=0.375
cc_3608 ( N_noxref_10_M26_noxref_d N_noxref_45_M26_noxref_s ) capacitor \
 c=0.0426368f //x=41.875 //y=0.915 //x2=41.445 //y2=0.375
cc_3609 ( N_noxref_10_c_4297_n N_noxref_46_c_11473_n ) capacitor c=3.84569e-19 \
 //x=42.465 //y=1.665 //x2=43.88 //y2=1.505
cc_3610 ( N_noxref_10_c_4304_n N_noxref_46_c_11473_n ) capacitor c=0.0034165f \
 //x=44.1 //y=1.915 //x2=43.88 //y2=1.505
cc_3611 ( N_noxref_10_c_4299_n N_noxref_46_c_11458_n ) capacitor c=0.0115578f \
 //x=44.4 //y=2.08 //x2=44.765 //y2=1.59
cc_3612 ( N_noxref_10_c_4303_n N_noxref_46_c_11458_n ) capacitor c=0.00697148f \
 //x=44.1 //y=1.53 //x2=44.765 //y2=1.59
cc_3613 ( N_noxref_10_c_4304_n N_noxref_46_c_11458_n ) capacitor c=0.0204849f \
 //x=44.1 //y=1.915 //x2=44.765 //y2=1.59
cc_3614 ( N_noxref_10_c_4306_n N_noxref_46_c_11458_n ) capacitor c=0.00610316f \
 //x=44.475 //y=1.375 //x2=44.765 //y2=1.59
cc_3615 ( N_noxref_10_c_4309_n N_noxref_46_c_11458_n ) capacitor c=0.00698822f \
 //x=44.63 //y=1.22 //x2=44.765 //y2=1.59
cc_3616 ( N_noxref_10_c_4300_n N_noxref_46_M27_noxref_s ) capacitor \
 c=0.0327271f //x=44.1 //y=0.875 //x2=43.745 //y2=0.375
cc_3617 ( N_noxref_10_c_4303_n N_noxref_46_M27_noxref_s ) capacitor \
 c=7.99997e-19 //x=44.1 //y=1.53 //x2=43.745 //y2=0.375
cc_3618 ( N_noxref_10_c_4304_n N_noxref_46_M27_noxref_s ) capacitor \
 c=0.00122123f //x=44.1 //y=1.915 //x2=43.745 //y2=0.375
cc_3619 ( N_noxref_10_c_4307_n N_noxref_46_M27_noxref_s ) capacitor \
 c=0.0121427f //x=44.63 //y=0.875 //x2=43.745 //y2=0.375
cc_3620 ( N_noxref_10_M26_noxref_d N_noxref_46_M27_noxref_s ) capacitor \
 c=2.55333e-19 //x=41.875 //y=0.915 //x2=43.745 //y2=0.375
cc_3621 ( N_noxref_11_c_4534_n N_noxref_12_c_4809_n ) capacitor c=0.0446157f \
 //x=37.625 //y=3.33 //x2=41.695 //y2=3.7
cc_3622 ( N_noxref_11_c_4541_n N_noxref_12_c_4809_n ) capacitor c=0.340407f \
 //x=49.095 //y=3.33 //x2=41.695 //y2=3.7
cc_3623 ( N_noxref_11_c_4543_n N_noxref_12_c_4809_n ) capacitor c=0.0268386f \
 //x=37.855 //y=3.33 //x2=41.695 //y2=3.7
cc_3624 ( N_noxref_11_c_4493_n N_noxref_12_c_4809_n ) capacitor c=0.0205782f \
 //x=37.74 //y=3.33 //x2=41.695 //y2=3.7
cc_3625 ( N_noxref_11_c_4534_n N_noxref_12_c_4849_n ) capacitor c=0.029444f \
 //x=37.625 //y=3.33 //x2=37.115 //y2=3.7
cc_3626 ( N_noxref_11_c_4493_n N_noxref_12_c_4849_n ) capacitor c=0.00179385f \
 //x=37.74 //y=3.33 //x2=37.115 //y2=3.7
cc_3627 ( N_noxref_11_c_4541_n N_noxref_12_c_4814_n ) capacitor c=0.468734f \
 //x=49.095 //y=3.33 //x2=47.245 //y2=3.7
cc_3628 ( N_noxref_11_c_4541_n N_noxref_12_c_4816_n ) capacitor c=0.026734f \
 //x=49.095 //y=3.33 //x2=41.925 //y2=3.7
cc_3629 ( N_noxref_11_c_4541_n N_noxref_12_c_4853_n ) capacitor c=0.176086f \
 //x=49.095 //y=3.33 //x2=56.125 //y2=3.7
cc_3630 ( N_noxref_11_c_4466_n N_noxref_12_c_4853_n ) capacitor c=0.0215974f \
 //x=49.21 //y=2.08 //x2=56.125 //y2=3.7
cc_3631 ( N_noxref_11_c_4541_n N_noxref_12_c_4855_n ) capacitor c=0.0268461f \
 //x=49.095 //y=3.33 //x2=47.475 //y2=3.7
cc_3632 ( N_noxref_11_c_4466_n N_noxref_12_c_4855_n ) capacitor c=7.01366e-19 \
 //x=49.21 //y=2.08 //x2=47.475 //y2=3.7
cc_3633 ( N_noxref_11_c_4534_n N_noxref_12_c_4745_n ) capacitor c=0.0198536f \
 //x=37.625 //y=3.33 //x2=37 //y2=2.08
cc_3634 ( N_noxref_11_c_4543_n N_noxref_12_c_4745_n ) capacitor c=0.00179385f \
 //x=37.855 //y=3.33 //x2=37 //y2=2.08
cc_3635 ( N_noxref_11_c_4493_n N_noxref_12_c_4745_n ) capacitor c=0.073434f \
 //x=37.74 //y=3.33 //x2=37 //y2=2.08
cc_3636 ( N_noxref_11_c_4595_p N_noxref_12_c_4745_n ) capacitor c=0.0126839f \
 //x=36.96 //y=5.155 //x2=37 //y2=2.08
cc_3637 ( N_noxref_11_c_4541_n N_noxref_12_c_4746_n ) capacitor c=0.0198536f \
 //x=49.095 //y=3.33 //x2=41.81 //y2=2.08
cc_3638 ( N_noxref_11_c_4541_n N_noxref_12_c_4766_n ) capacitor c=0.0212788f \
 //x=49.095 //y=3.33 //x2=47.36 //y2=3.7
cc_3639 ( N_noxref_11_c_4466_n N_noxref_12_c_4766_n ) capacitor c=0.0104866f \
 //x=49.21 //y=2.08 //x2=47.36 //y2=3.7
cc_3640 ( N_noxref_11_c_4485_n N_noxref_12_M106_noxref_g ) capacitor \
 c=0.0162556f //x=36.875 //y=5.155 //x2=36.74 //y2=6.02
cc_3641 ( N_noxref_11_M106_noxref_d N_noxref_12_M106_noxref_g ) capacitor \
 c=0.0180032f //x=36.815 //y=5.02 //x2=36.74 //y2=6.02
cc_3642 ( N_noxref_11_c_4489_n N_noxref_12_M107_noxref_g ) capacitor \
 c=0.0183937f //x=37.655 //y=5.155 //x2=37.18 //y2=6.02
cc_3643 ( N_noxref_11_M106_noxref_d N_noxref_12_M107_noxref_g ) capacitor \
 c=0.0194246f //x=36.815 //y=5.02 //x2=37.18 //y2=6.02
cc_3644 ( N_noxref_11_M23_noxref_d N_noxref_12_c_4868_n ) capacitor \
 c=0.00217566f //x=37.065 //y=0.915 //x2=36.99 //y2=0.915
cc_3645 ( N_noxref_11_M23_noxref_d N_noxref_12_c_4869_n ) capacitor \
 c=0.0034598f //x=37.065 //y=0.915 //x2=36.99 //y2=1.26
cc_3646 ( N_noxref_11_M23_noxref_d N_noxref_12_c_4870_n ) capacitor \
 c=0.00546784f //x=37.065 //y=0.915 //x2=36.99 //y2=1.57
cc_3647 ( N_noxref_11_M23_noxref_d N_noxref_12_c_4871_n ) capacitor \
 c=0.00241102f //x=37.065 //y=0.915 //x2=37.365 //y2=0.76
cc_3648 ( N_noxref_11_c_4465_n N_noxref_12_c_4872_n ) capacitor c=0.00371277f \
 //x=37.655 //y=1.665 //x2=37.365 //y2=1.415
cc_3649 ( N_noxref_11_M23_noxref_d N_noxref_12_c_4872_n ) capacitor \
 c=0.0138621f //x=37.065 //y=0.915 //x2=37.365 //y2=1.415
cc_3650 ( N_noxref_11_M23_noxref_d N_noxref_12_c_4874_n ) capacitor \
 c=0.00219619f //x=37.065 //y=0.915 //x2=37.52 //y2=0.915
cc_3651 ( N_noxref_11_c_4465_n N_noxref_12_c_4875_n ) capacitor c=0.00457401f \
 //x=37.655 //y=1.665 //x2=37.52 //y2=1.26
cc_3652 ( N_noxref_11_M23_noxref_d N_noxref_12_c_4875_n ) capacitor \
 c=0.00603828f //x=37.065 //y=0.915 //x2=37.52 //y2=1.26
cc_3653 ( N_noxref_11_c_4493_n N_noxref_12_c_4877_n ) capacitor c=0.00731987f \
 //x=37.74 //y=3.33 //x2=37 //y2=2.08
cc_3654 ( N_noxref_11_c_4493_n N_noxref_12_c_4878_n ) capacitor c=0.00283672f \
 //x=37.74 //y=3.33 //x2=37 //y2=1.915
cc_3655 ( N_noxref_11_M23_noxref_d N_noxref_12_c_4878_n ) capacitor \
 c=0.00661782f //x=37.065 //y=0.915 //x2=37 //y2=1.915
cc_3656 ( N_noxref_11_c_4489_n N_noxref_12_c_4806_n ) capacitor c=0.00201851f \
 //x=37.655 //y=5.155 //x2=37 //y2=4.7
cc_3657 ( N_noxref_11_c_4493_n N_noxref_12_c_4806_n ) capacitor c=0.0114782f \
 //x=37.74 //y=3.33 //x2=37 //y2=4.7
cc_3658 ( N_noxref_11_c_4595_p N_noxref_12_c_4806_n ) capacitor c=0.00470675f \
 //x=36.96 //y=5.155 //x2=37 //y2=4.7
cc_3659 ( N_noxref_11_c_4466_n N_noxref_13_c_5101_n ) capacitor c=0.00121487f \
 //x=49.21 //y=2.08 //x2=51.43 //y2=2.08
cc_3660 ( N_noxref_11_c_4534_n N_D_c_5328_n ) capacitor c=0.202839f //x=37.625 \
 //y=3.33 //x2=58.715 //y2=4.07
cc_3661 ( N_noxref_11_c_4533_n N_D_c_5328_n ) capacitor c=0.0135672f \
 //x=32.305 //y=3.33 //x2=58.715 //y2=4.07
cc_3662 ( N_noxref_11_c_4541_n N_D_c_5328_n ) capacitor c=0.0809428f \
 //x=49.095 //y=3.33 //x2=58.715 //y2=4.07
cc_3663 ( N_noxref_11_c_4543_n N_D_c_5328_n ) capacitor c=4.80262e-19 \
 //x=37.855 //y=3.33 //x2=58.715 //y2=4.07
cc_3664 ( N_noxref_11_c_4464_n N_D_c_5328_n ) capacitor c=0.0206302f //x=32.19 \
 //y=2.08 //x2=58.715 //y2=4.07
cc_3665 ( N_noxref_11_c_4493_n N_D_c_5328_n ) capacitor c=0.0181789f //x=37.74 \
 //y=3.33 //x2=58.715 //y2=4.07
cc_3666 ( N_noxref_11_c_4466_n N_D_c_5328_n ) capacitor c=0.0194977f //x=49.21 \
 //y=2.08 //x2=58.715 //y2=4.07
cc_3667 ( N_noxref_11_c_4464_n N_D_c_5280_n ) capacitor c=0.0014206f //x=32.19 \
 //y=2.08 //x2=29.97 //y2=2.08
cc_3668 ( N_noxref_11_c_4534_n N_CLK_c_6058_n ) capacitor c=0.0174494f \
 //x=37.625 //y=3.33 //x2=35.775 //y2=4.44
cc_3669 ( N_noxref_11_c_4533_n N_CLK_c_6058_n ) capacitor c=4.49102e-19 \
 //x=32.305 //y=3.33 //x2=35.775 //y2=4.44
cc_3670 ( N_noxref_11_c_4464_n N_CLK_c_6058_n ) capacitor c=0.0178424f \
 //x=32.19 //y=2.08 //x2=35.775 //y2=4.44
cc_3671 ( N_noxref_11_c_4532_n N_CLK_c_6058_n ) capacitor c=0.00731624f \
 //x=32.19 //y=4.7 //x2=35.775 //y2=4.44
cc_3672 ( N_noxref_11_c_4534_n N_CLK_c_6068_n ) capacitor c=0.00667512f \
 //x=37.625 //y=3.33 //x2=45.395 //y2=4.44
cc_3673 ( N_noxref_11_c_4493_n N_CLK_c_6068_n ) capacitor c=0.0166101f \
 //x=37.74 //y=3.33 //x2=45.395 //y2=4.44
cc_3674 ( N_noxref_11_c_4534_n N_CLK_c_6190_n ) capacitor c=5.01525e-19 \
 //x=37.625 //y=3.33 //x2=36.005 //y2=4.44
cc_3675 ( N_noxref_11_c_4466_n N_CLK_c_6070_n ) capacitor c=0.018786f \
 //x=49.21 //y=2.08 //x2=64.635 //y2=4.44
cc_3676 ( N_noxref_11_c_4505_n N_CLK_c_6070_n ) capacitor c=0.0112124f \
 //x=49.485 //y=4.79 //x2=64.635 //y2=4.44
cc_3677 ( N_noxref_11_c_4534_n N_CLK_c_6042_n ) capacitor c=0.0213922f \
 //x=37.625 //y=3.33 //x2=35.89 //y2=2.08
cc_3678 ( N_noxref_11_c_4479_n N_CLK_c_6042_n ) capacitor c=0.0121898f \
 //x=35.995 //y=5.155 //x2=35.89 //y2=2.08
cc_3679 ( N_noxref_11_c_4493_n N_CLK_c_6042_n ) capacitor c=0.00220975f \
 //x=37.74 //y=3.33 //x2=35.89 //y2=2.08
cc_3680 ( N_noxref_11_c_4541_n N_CLK_c_6043_n ) capacitor c=0.0190562f \
 //x=49.095 //y=3.33 //x2=45.51 //y2=2.08
cc_3681 ( N_noxref_11_c_4479_n N_CLK_M104_noxref_g ) capacitor c=0.0163793f \
 //x=35.995 //y=5.155 //x2=35.86 //y2=6.02
cc_3682 ( N_noxref_11_M104_noxref_d N_CLK_M104_noxref_g ) capacitor \
 c=0.0180032f //x=35.935 //y=5.02 //x2=35.86 //y2=6.02
cc_3683 ( N_noxref_11_c_4485_n N_CLK_M105_noxref_g ) capacitor c=0.0162556f \
 //x=36.875 //y=5.155 //x2=36.3 //y2=6.02
cc_3684 ( N_noxref_11_M104_noxref_d N_CLK_M105_noxref_g ) capacitor \
 c=0.0180032f //x=35.935 //y=5.02 //x2=36.3 //y2=6.02
cc_3685 ( N_noxref_11_c_4644_p N_CLK_c_6211_n ) capacitor c=0.00392095f \
 //x=36.08 //y=5.155 //x2=36.225 //y2=4.79
cc_3686 ( N_noxref_11_c_4479_n N_CLK_c_6215_n ) capacitor c=0.00309994f \
 //x=35.995 //y=5.155 //x2=35.89 //y2=4.7
cc_3687 ( N_noxref_11_c_4534_n N_RN_c_7046_n ) capacitor c=0.00374603f \
 //x=37.625 //y=3.33 //x2=46.505 //y2=2.22
cc_3688 ( N_noxref_11_c_4533_n N_RN_c_7046_n ) capacitor c=7.32243e-19 \
 //x=32.305 //y=3.33 //x2=46.505 //y2=2.22
cc_3689 ( N_noxref_11_c_4541_n N_RN_c_7046_n ) capacitor c=0.0316113f \
 //x=49.095 //y=3.33 //x2=46.505 //y2=2.22
cc_3690 ( N_noxref_11_c_4464_n N_RN_c_7046_n ) capacitor c=0.0209607f \
 //x=32.19 //y=2.08 //x2=46.505 //y2=2.22
cc_3691 ( N_noxref_11_c_4650_p N_RN_c_7046_n ) capacitor c=0.016327f //x=37.34 \
 //y=1.665 //x2=46.505 //y2=2.22
cc_3692 ( N_noxref_11_c_4493_n N_RN_c_7046_n ) capacitor c=0.0197307f \
 //x=37.74 //y=3.33 //x2=46.505 //y2=2.22
cc_3693 ( N_noxref_11_c_4563_n N_RN_c_7046_n ) capacitor c=3.13485e-19 \
 //x=32.555 //y=1.415 //x2=46.505 //y2=2.22
cc_3694 ( N_noxref_11_c_4568_n N_RN_c_7046_n ) capacitor c=0.00584491f \
 //x=32.19 //y=2.08 //x2=46.505 //y2=2.22
cc_3695 ( N_noxref_11_c_4464_n N_RN_c_7057_n ) capacitor c=0.00165648f \
 //x=32.19 //y=2.08 //x2=31.195 //y2=2.22
cc_3696 ( N_noxref_11_c_4568_n N_RN_c_7057_n ) capacitor c=2.3323e-19 \
 //x=32.19 //y=2.08 //x2=31.195 //y2=2.22
cc_3697 ( N_noxref_11_c_4541_n N_RN_c_7058_n ) capacitor c=0.014255f \
 //x=49.095 //y=3.33 //x2=50.205 //y2=2.22
cc_3698 ( N_noxref_11_c_4466_n N_RN_c_7058_n ) capacitor c=0.0216101f \
 //x=49.21 //y=2.08 //x2=50.205 //y2=2.22
cc_3699 ( N_noxref_11_c_4471_n N_RN_c_7058_n ) capacitor c=0.011987f //x=48.91 \
 //y=1.915 //x2=50.205 //y2=2.22
cc_3700 ( N_noxref_11_c_4541_n N_RN_c_7062_n ) capacitor c=4.86139e-19 \
 //x=49.095 //y=3.33 //x2=46.735 //y2=2.22
cc_3701 ( N_noxref_11_c_4466_n N_RN_c_7070_n ) capacitor c=0.00100368f \
 //x=49.21 //y=2.08 //x2=50.435 //y2=2.22
cc_3702 ( N_noxref_11_c_4471_n N_RN_c_7070_n ) capacitor c=2.11894e-19 \
 //x=48.91 //y=1.915 //x2=50.435 //y2=2.22
cc_3703 ( N_noxref_11_c_4533_n N_RN_c_7091_n ) capacitor c=0.00350495f \
 //x=32.305 //y=3.33 //x2=31.08 //y2=2.08
cc_3704 ( N_noxref_11_c_4464_n N_RN_c_7091_n ) capacitor c=0.0448384f \
 //x=32.19 //y=2.08 //x2=31.08 //y2=2.08
cc_3705 ( N_noxref_11_c_4568_n N_RN_c_7091_n ) capacitor c=0.0019893f \
 //x=32.19 //y=2.08 //x2=31.08 //y2=2.08
cc_3706 ( N_noxref_11_c_4532_n N_RN_c_7091_n ) capacitor c=0.00197875f \
 //x=32.19 //y=4.7 //x2=31.08 //y2=2.08
cc_3707 ( N_noxref_11_c_4541_n N_RN_c_7092_n ) capacitor c=0.0180187f \
 //x=49.095 //y=3.33 //x2=46.62 //y2=2.08
cc_3708 ( N_noxref_11_c_4466_n N_RN_c_7092_n ) capacitor c=6.89573e-19 \
 //x=49.21 //y=2.08 //x2=46.62 //y2=2.08
cc_3709 ( N_noxref_11_c_4541_n N_RN_c_7093_n ) capacitor c=0.00311593f \
 //x=49.095 //y=3.33 //x2=50.32 //y2=2.08
cc_3710 ( N_noxref_11_c_4466_n N_RN_c_7093_n ) capacitor c=0.0430926f \
 //x=49.21 //y=2.08 //x2=50.32 //y2=2.08
cc_3711 ( N_noxref_11_c_4471_n N_RN_c_7093_n ) capacitor c=0.00208635f \
 //x=48.91 //y=1.915 //x2=50.32 //y2=2.08
cc_3712 ( N_noxref_11_c_4530_n N_RN_c_7093_n ) capacitor c=0.00120758f \
 //x=49.775 //y=4.79 //x2=50.32 //y2=2.08
cc_3713 ( N_noxref_11_c_4505_n N_RN_c_7093_n ) capacitor c=0.00142741f \
 //x=49.485 //y=4.79 //x2=50.32 //y2=2.08
cc_3714 ( N_noxref_11_M100_noxref_g N_RN_M98_noxref_g ) capacitor c=0.0100903f \
 //x=31.93 //y=6.02 //x2=31.05 //y2=6.02
cc_3715 ( N_noxref_11_M100_noxref_g N_RN_M99_noxref_g ) capacitor c=0.0600064f \
 //x=31.93 //y=6.02 //x2=31.49 //y2=6.02
cc_3716 ( N_noxref_11_M101_noxref_g N_RN_M99_noxref_g ) capacitor c=0.0100903f \
 //x=32.37 //y=6.02 //x2=31.49 //y2=6.02
cc_3717 ( N_noxref_11_M120_noxref_g N_RN_M122_noxref_g ) capacitor \
 c=0.0105174f //x=49.41 //y=6.02 //x2=50.29 //y2=6.02
cc_3718 ( N_noxref_11_M121_noxref_g N_RN_M122_noxref_g ) capacitor c=0.10624f \
 //x=49.85 //y=6.02 //x2=50.29 //y2=6.02
cc_3719 ( N_noxref_11_M121_noxref_g N_RN_M123_noxref_g ) capacitor \
 c=0.0100903f //x=49.85 //y=6.02 //x2=50.73 //y2=6.02
cc_3720 ( N_noxref_11_c_4559_n N_RN_c_7394_n ) capacitor c=0.00456962f \
 //x=32.18 //y=0.915 //x2=31.17 //y2=0.91
cc_3721 ( N_noxref_11_c_4560_n N_RN_c_7395_n ) capacitor c=0.00438372f \
 //x=32.18 //y=1.26 //x2=31.17 //y2=1.22
cc_3722 ( N_noxref_11_c_4561_n N_RN_c_7396_n ) capacitor c=0.00438372f \
 //x=32.18 //y=1.57 //x2=31.17 //y2=1.45
cc_3723 ( N_noxref_11_c_4464_n N_RN_c_7397_n ) capacitor c=0.00205895f \
 //x=32.19 //y=2.08 //x2=31.17 //y2=1.915
cc_3724 ( N_noxref_11_c_4568_n N_RN_c_7397_n ) capacitor c=0.00828003f \
 //x=32.19 //y=2.08 //x2=31.17 //y2=1.915
cc_3725 ( N_noxref_11_c_4569_n N_RN_c_7397_n ) capacitor c=0.00438372f \
 //x=32.19 //y=1.915 //x2=31.17 //y2=1.915
cc_3726 ( N_noxref_11_c_4532_n N_RN_c_7256_n ) capacitor c=0.0609323f \
 //x=32.19 //y=4.7 //x2=31.415 //y2=4.79
cc_3727 ( N_noxref_11_c_4467_n N_RN_c_7401_n ) capacitor c=5.72482e-19 \
 //x=48.91 //y=0.875 //x2=49.885 //y2=0.91
cc_3728 ( N_noxref_11_c_4469_n N_RN_c_7401_n ) capacitor c=0.00149976f \
 //x=48.91 //y=1.22 //x2=49.885 //y2=0.91
cc_3729 ( N_noxref_11_c_4474_n N_RN_c_7401_n ) capacitor c=0.0160123f \
 //x=49.44 //y=0.875 //x2=49.885 //y2=0.91
cc_3730 ( N_noxref_11_c_4470_n N_RN_c_7404_n ) capacitor c=0.00111227f \
 //x=48.91 //y=1.53 //x2=49.885 //y2=1.22
cc_3731 ( N_noxref_11_c_4476_n N_RN_c_7404_n ) capacitor c=0.0124075f \
 //x=49.44 //y=1.22 //x2=49.885 //y2=1.22
cc_3732 ( N_noxref_11_c_4474_n N_RN_c_7406_n ) capacitor c=0.00103227f \
 //x=49.44 //y=0.875 //x2=50.41 //y2=0.91
cc_3733 ( N_noxref_11_c_4476_n N_RN_c_7407_n ) capacitor c=0.0010154f \
 //x=49.44 //y=1.22 //x2=50.41 //y2=1.22
cc_3734 ( N_noxref_11_c_4476_n N_RN_c_7408_n ) capacitor c=9.23422e-19 \
 //x=49.44 //y=1.22 //x2=50.41 //y2=1.45
cc_3735 ( N_noxref_11_c_4466_n N_RN_c_7409_n ) capacitor c=0.00203769f \
 //x=49.21 //y=2.08 //x2=50.41 //y2=1.915
cc_3736 ( N_noxref_11_c_4471_n N_RN_c_7409_n ) capacitor c=0.00834532f \
 //x=48.91 //y=1.915 //x2=50.41 //y2=1.915
cc_3737 ( N_noxref_11_c_4464_n N_RN_c_7261_n ) capacitor c=0.00142741f \
 //x=32.19 //y=2.08 //x2=31.08 //y2=4.7
cc_3738 ( N_noxref_11_c_4532_n N_RN_c_7261_n ) capacitor c=0.00487508f \
 //x=32.19 //y=4.7 //x2=31.08 //y2=4.7
cc_3739 ( N_noxref_11_c_4466_n N_RN_c_7263_n ) capacitor c=0.0017365f \
 //x=49.21 //y=2.08 //x2=50.32 //y2=4.7
cc_3740 ( N_noxref_11_c_4530_n N_RN_c_7263_n ) capacitor c=0.0170104f \
 //x=49.775 //y=4.79 //x2=50.32 //y2=4.7
cc_3741 ( N_noxref_11_c_4505_n N_RN_c_7263_n ) capacitor c=0.00484466f \
 //x=49.485 //y=4.79 //x2=50.32 //y2=4.7
cc_3742 ( N_noxref_11_c_4534_n N_SN_c_8132_n ) capacitor c=0.466581f \
 //x=37.625 //y=3.33 //x2=40.585 //y2=2.96
cc_3743 ( N_noxref_11_c_4533_n N_SN_c_8132_n ) capacitor c=0.0291389f \
 //x=32.305 //y=3.33 //x2=40.585 //y2=2.96
cc_3744 ( N_noxref_11_c_4541_n N_SN_c_8132_n ) capacitor c=0.241804f \
 //x=49.095 //y=3.33 //x2=40.585 //y2=2.96
cc_3745 ( N_noxref_11_c_4543_n N_SN_c_8132_n ) capacitor c=0.0266688f \
 //x=37.855 //y=3.33 //x2=40.585 //y2=2.96
cc_3746 ( N_noxref_11_c_4464_n N_SN_c_8132_n ) capacitor c=0.0221202f \
 //x=32.19 //y=2.08 //x2=40.585 //y2=2.96
cc_3747 ( N_noxref_11_c_4493_n N_SN_c_8132_n ) capacitor c=0.020574f //x=37.74 \
 //y=3.33 //x2=40.585 //y2=2.96
cc_3748 ( N_noxref_11_c_4541_n N_SN_c_8135_n ) capacitor c=0.756732f \
 //x=49.095 //y=3.33 //x2=55.015 //y2=2.96
cc_3749 ( N_noxref_11_c_4466_n N_SN_c_8135_n ) capacitor c=0.0238838f \
 //x=49.21 //y=2.08 //x2=55.015 //y2=2.96
cc_3750 ( N_noxref_11_c_4541_n N_SN_c_8340_n ) capacitor c=0.0265806f \
 //x=49.095 //y=3.33 //x2=40.815 //y2=2.96
cc_3751 ( N_noxref_11_c_4541_n N_SN_c_8147_n ) capacitor c=0.0208912f \
 //x=49.095 //y=3.33 //x2=40.7 //y2=2.08
cc_3752 ( N_noxref_11_c_4493_n N_SN_c_8147_n ) capacitor c=3.55725e-19 \
 //x=37.74 //y=3.33 //x2=40.7 //y2=2.08
cc_3753 ( N_noxref_11_c_4541_n N_noxref_26_c_10043_n ) capacitor c=0.00564994f \
 //x=49.095 //y=3.33 //x2=52.285 //y2=3.33
cc_3754 ( N_noxref_11_M121_noxref_g N_noxref_26_c_9944_n ) capacitor \
 c=0.0157304f //x=49.85 //y=6.02 //x2=50.425 //y2=5.155
cc_3755 ( N_noxref_11_M120_noxref_g N_noxref_26_c_9948_n ) capacitor \
 c=0.0213876f //x=49.41 //y=6.02 //x2=49.715 //y2=5.155
cc_3756 ( N_noxref_11_c_4530_n N_noxref_26_c_9948_n ) capacitor c=0.00393496f \
 //x=49.775 //y=4.79 //x2=49.715 //y2=5.155
cc_3757 ( N_noxref_11_M121_noxref_g N_noxref_26_M120_noxref_d ) capacitor \
 c=0.0180032f //x=49.85 //y=6.02 //x2=49.485 //y2=5.02
cc_3758 ( N_noxref_11_c_4464_n N_noxref_41_c_11209_n ) capacitor c=0.00204385f \
 //x=32.19 //y=2.08 //x2=32.845 //y2=0.54
cc_3759 ( N_noxref_11_c_4559_n N_noxref_41_c_11209_n ) capacitor c=0.0194423f \
 //x=32.18 //y=0.915 //x2=32.845 //y2=0.54
cc_3760 ( N_noxref_11_c_4565_n N_noxref_41_c_11209_n ) capacitor c=0.00656458f \
 //x=32.71 //y=0.915 //x2=32.845 //y2=0.54
cc_3761 ( N_noxref_11_c_4568_n N_noxref_41_c_11209_n ) capacitor c=2.20712e-19 \
 //x=32.19 //y=2.08 //x2=32.845 //y2=0.54
cc_3762 ( N_noxref_11_c_4560_n N_noxref_41_c_11219_n ) capacitor c=0.00538829f \
 //x=32.18 //y=1.26 //x2=31.96 //y2=0.995
cc_3763 ( N_noxref_11_c_4559_n N_noxref_41_M20_noxref_s ) capacitor \
 c=0.00538829f //x=32.18 //y=0.915 //x2=31.825 //y2=0.375
cc_3764 ( N_noxref_11_c_4561_n N_noxref_41_M20_noxref_s ) capacitor \
 c=0.00538829f //x=32.18 //y=1.57 //x2=31.825 //y2=0.375
cc_3765 ( N_noxref_11_c_4565_n N_noxref_41_M20_noxref_s ) capacitor \
 c=0.0143002f //x=32.71 //y=0.915 //x2=31.825 //y2=0.375
cc_3766 ( N_noxref_11_c_4566_n N_noxref_41_M20_noxref_s ) capacitor \
 c=0.00290153f //x=32.71 //y=1.26 //x2=31.825 //y2=0.375
cc_3767 ( N_noxref_11_M23_noxref_d N_noxref_42_M21_noxref_s ) capacitor \
 c=0.00309936f //x=37.065 //y=0.915 //x2=34.125 //y2=0.375
cc_3768 ( N_noxref_11_c_4465_n N_noxref_43_c_11310_n ) capacitor c=0.00457167f \
 //x=37.655 //y=1.665 //x2=37.655 //y2=0.54
cc_3769 ( N_noxref_11_M23_noxref_d N_noxref_43_c_11310_n ) capacitor \
 c=0.0115903f //x=37.065 //y=0.915 //x2=37.655 //y2=0.54
cc_3770 ( N_noxref_11_c_4650_p N_noxref_43_c_11320_n ) capacitor c=0.0200405f \
 //x=37.34 //y=1.665 //x2=36.77 //y2=0.995
cc_3771 ( N_noxref_11_M23_noxref_d N_noxref_43_M22_noxref_d ) capacitor \
 c=5.27807e-19 //x=37.065 //y=0.915 //x2=35.53 //y2=0.91
cc_3772 ( N_noxref_11_c_4465_n N_noxref_43_M23_noxref_s ) capacitor \
 c=0.0196084f //x=37.655 //y=1.665 //x2=36.635 //y2=0.375
cc_3773 ( N_noxref_11_M23_noxref_d N_noxref_43_M23_noxref_s ) capacitor \
 c=0.0426368f //x=37.065 //y=0.915 //x2=36.635 //y2=0.375
cc_3774 ( N_noxref_11_c_4465_n N_noxref_44_c_11372_n ) capacitor c=3.84569e-19 \
 //x=37.655 //y=1.665 //x2=39.07 //y2=1.505
cc_3775 ( N_noxref_11_M23_noxref_d N_noxref_44_M24_noxref_s ) capacitor \
 c=2.55333e-19 //x=37.065 //y=0.915 //x2=38.935 //y2=0.375
cc_3776 ( N_noxref_11_c_4471_n N_noxref_48_c_11575_n ) capacitor c=0.0034165f \
 //x=48.91 //y=1.915 //x2=48.69 //y2=1.505
cc_3777 ( N_noxref_11_c_4466_n N_noxref_48_c_11560_n ) capacitor c=0.0115578f \
 //x=49.21 //y=2.08 //x2=49.575 //y2=1.59
cc_3778 ( N_noxref_11_c_4470_n N_noxref_48_c_11560_n ) capacitor c=0.00697148f \
 //x=48.91 //y=1.53 //x2=49.575 //y2=1.59
cc_3779 ( N_noxref_11_c_4471_n N_noxref_48_c_11560_n ) capacitor c=0.0204849f \
 //x=48.91 //y=1.915 //x2=49.575 //y2=1.59
cc_3780 ( N_noxref_11_c_4473_n N_noxref_48_c_11560_n ) capacitor c=0.00610316f \
 //x=49.285 //y=1.375 //x2=49.575 //y2=1.59
cc_3781 ( N_noxref_11_c_4476_n N_noxref_48_c_11560_n ) capacitor c=0.00698822f \
 //x=49.44 //y=1.22 //x2=49.575 //y2=1.59
cc_3782 ( N_noxref_11_c_4467_n N_noxref_48_M30_noxref_s ) capacitor \
 c=0.0327271f //x=48.91 //y=0.875 //x2=48.555 //y2=0.375
cc_3783 ( N_noxref_11_c_4470_n N_noxref_48_M30_noxref_s ) capacitor \
 c=7.99997e-19 //x=48.91 //y=1.53 //x2=48.555 //y2=0.375
cc_3784 ( N_noxref_11_c_4471_n N_noxref_48_M30_noxref_s ) capacitor \
 c=0.00122123f //x=48.91 //y=1.915 //x2=48.555 //y2=0.375
cc_3785 ( N_noxref_11_c_4474_n N_noxref_48_M30_noxref_s ) capacitor \
 c=0.0121427f //x=49.44 //y=0.875 //x2=48.555 //y2=0.375
cc_3786 ( N_noxref_12_c_4853_n N_noxref_13_c_5099_n ) capacitor c=0.00376735f \
 //x=56.125 //y=3.7 //x2=56.865 //y2=2.59
cc_3787 ( N_noxref_12_c_4748_n N_noxref_13_c_5099_n ) capacitor c=0.0197567f \
 //x=56.24 //y=2.08 //x2=56.865 //y2=2.59
cc_3788 ( N_noxref_12_c_4853_n N_noxref_13_c_5149_n ) capacitor c=6.53213e-19 \
 //x=56.125 //y=3.7 //x2=51.545 //y2=2.59
cc_3789 ( N_noxref_12_c_4853_n N_noxref_13_c_5101_n ) capacitor c=0.0203405f \
 //x=56.125 //y=3.7 //x2=51.43 //y2=2.08
cc_3790 ( N_noxref_12_M130_noxref_g N_noxref_13_c_5112_n ) capacitor \
 c=0.0162556f //x=55.98 //y=6.02 //x2=56.115 //y2=5.155
cc_3791 ( N_noxref_12_M131_noxref_g N_noxref_13_c_5116_n ) capacitor \
 c=0.0183937f //x=56.42 //y=6.02 //x2=56.895 //y2=5.155
cc_3792 ( N_noxref_12_c_4808_n N_noxref_13_c_5116_n ) capacitor c=0.00201851f \
 //x=56.24 //y=4.7 //x2=56.895 //y2=5.155
cc_3793 ( N_noxref_12_c_4890_p N_noxref_13_c_5102_n ) capacitor c=0.00371277f \
 //x=56.605 //y=1.415 //x2=56.895 //y2=1.665
cc_3794 ( N_noxref_12_c_4891_p N_noxref_13_c_5102_n ) capacitor c=0.00457401f \
 //x=56.76 //y=1.26 //x2=56.895 //y2=1.665
cc_3795 ( N_noxref_12_c_4853_n N_noxref_13_c_5103_n ) capacitor c=0.00262125f \
 //x=56.125 //y=3.7 //x2=56.98 //y2=2.59
cc_3796 ( N_noxref_12_c_4748_n N_noxref_13_c_5103_n ) capacitor c=0.0724336f \
 //x=56.24 //y=2.08 //x2=56.98 //y2=2.59
cc_3797 ( N_noxref_12_c_4894_p N_noxref_13_c_5103_n ) capacitor c=0.00709342f \
 //x=56.24 //y=2.08 //x2=56.98 //y2=2.59
cc_3798 ( N_noxref_12_c_4895_p N_noxref_13_c_5103_n ) capacitor c=0.00283672f \
 //x=56.24 //y=1.915 //x2=56.98 //y2=2.59
cc_3799 ( N_noxref_12_c_4808_n N_noxref_13_c_5103_n ) capacitor c=0.0116291f \
 //x=56.24 //y=4.7 //x2=56.98 //y2=2.59
cc_3800 ( N_noxref_12_c_4748_n N_noxref_13_c_5161_n ) capacitor c=0.0126839f \
 //x=56.24 //y=2.08 //x2=56.2 //y2=5.155
cc_3801 ( N_noxref_12_c_4808_n N_noxref_13_c_5161_n ) capacitor c=0.00470675f \
 //x=56.24 //y=4.7 //x2=56.2 //y2=5.155
cc_3802 ( N_noxref_12_c_4899_p N_noxref_13_M35_noxref_d ) capacitor \
 c=0.00217566f //x=56.23 //y=0.915 //x2=56.305 //y2=0.915
cc_3803 ( N_noxref_12_c_4900_p N_noxref_13_M35_noxref_d ) capacitor \
 c=0.0034598f //x=56.23 //y=1.26 //x2=56.305 //y2=0.915
cc_3804 ( N_noxref_12_c_4901_p N_noxref_13_M35_noxref_d ) capacitor \
 c=0.00546784f //x=56.23 //y=1.57 //x2=56.305 //y2=0.915
cc_3805 ( N_noxref_12_c_4902_p N_noxref_13_M35_noxref_d ) capacitor \
 c=0.00241102f //x=56.605 //y=0.76 //x2=56.305 //y2=0.915
cc_3806 ( N_noxref_12_c_4890_p N_noxref_13_M35_noxref_d ) capacitor \
 c=0.0138621f //x=56.605 //y=1.415 //x2=56.305 //y2=0.915
cc_3807 ( N_noxref_12_c_4904_p N_noxref_13_M35_noxref_d ) capacitor \
 c=0.00219619f //x=56.76 //y=0.915 //x2=56.305 //y2=0.915
cc_3808 ( N_noxref_12_c_4891_p N_noxref_13_M35_noxref_d ) capacitor \
 c=0.00603828f //x=56.76 //y=1.26 //x2=56.305 //y2=0.915
cc_3809 ( N_noxref_12_c_4895_p N_noxref_13_M35_noxref_d ) capacitor \
 c=0.00661782f //x=56.24 //y=1.915 //x2=56.305 //y2=0.915
cc_3810 ( N_noxref_12_M130_noxref_g N_noxref_13_M130_noxref_d ) capacitor \
 c=0.0180032f //x=55.98 //y=6.02 //x2=56.055 //y2=5.02
cc_3811 ( N_noxref_12_M131_noxref_g N_noxref_13_M130_noxref_d ) capacitor \
 c=0.0194246f //x=56.42 //y=6.02 //x2=56.055 //y2=5.02
cc_3812 ( N_noxref_12_c_4809_n N_D_c_5328_n ) capacitor c=0.403974f //x=41.695 \
 //y=3.7 //x2=58.715 //y2=4.07
cc_3813 ( N_noxref_12_c_4849_n N_D_c_5328_n ) capacitor c=0.0292842f \
 //x=37.115 //y=3.7 //x2=58.715 //y2=4.07
cc_3814 ( N_noxref_12_c_4814_n N_D_c_5328_n ) capacitor c=0.468094f //x=47.245 \
 //y=3.7 //x2=58.715 //y2=4.07
cc_3815 ( N_noxref_12_c_4816_n N_D_c_5328_n ) capacitor c=0.026596f //x=41.925 \
 //y=3.7 //x2=58.715 //y2=4.07
cc_3816 ( N_noxref_12_c_4853_n N_D_c_5328_n ) capacitor c=0.792602f //x=56.125 \
 //y=3.7 //x2=58.715 //y2=4.07
cc_3817 ( N_noxref_12_c_4855_n N_D_c_5328_n ) capacitor c=0.026809f //x=47.475 \
 //y=3.7 //x2=58.715 //y2=4.07
cc_3818 ( N_noxref_12_c_4745_n N_D_c_5328_n ) capacitor c=0.0198068f //x=37 \
 //y=2.08 //x2=58.715 //y2=4.07
cc_3819 ( N_noxref_12_c_4746_n N_D_c_5328_n ) capacitor c=0.0198068f //x=41.81 \
 //y=2.08 //x2=58.715 //y2=4.07
cc_3820 ( N_noxref_12_c_4766_n N_D_c_5328_n ) capacitor c=0.0200135f //x=47.36 \
 //y=3.7 //x2=58.715 //y2=4.07
cc_3821 ( N_noxref_12_c_4748_n N_D_c_5328_n ) capacitor c=0.0198068f //x=56.24 \
 //y=2.08 //x2=58.715 //y2=4.07
cc_3822 ( N_noxref_12_c_4748_n N_D_c_5281_n ) capacitor c=9.22611e-19 \
 //x=56.24 //y=2.08 //x2=58.83 //y2=2.08
cc_3823 ( N_noxref_12_c_4809_n N_CLK_c_6068_n ) capacitor c=0.0344845f \
 //x=41.695 //y=3.7 //x2=45.395 //y2=4.44
cc_3824 ( N_noxref_12_c_4849_n N_CLK_c_6068_n ) capacitor c=7.0371e-19 \
 //x=37.115 //y=3.7 //x2=45.395 //y2=4.44
cc_3825 ( N_noxref_12_c_4814_n N_CLK_c_6068_n ) capacitor c=0.0246711f \
 //x=47.245 //y=3.7 //x2=45.395 //y2=4.44
cc_3826 ( N_noxref_12_c_4816_n N_CLK_c_6068_n ) capacitor c=4.78625e-19 \
 //x=41.925 //y=3.7 //x2=45.395 //y2=4.44
cc_3827 ( N_noxref_12_c_4745_n N_CLK_c_6068_n ) capacitor c=0.0178424f //x=37 \
 //y=2.08 //x2=45.395 //y2=4.44
cc_3828 ( N_noxref_12_c_4746_n N_CLK_c_6068_n ) capacitor c=0.0178424f \
 //x=41.81 //y=2.08 //x2=45.395 //y2=4.44
cc_3829 ( N_noxref_12_c_4806_n N_CLK_c_6068_n ) capacitor c=0.00731624f //x=37 \
 //y=4.7 //x2=45.395 //y2=4.44
cc_3830 ( N_noxref_12_c_4807_n N_CLK_c_6068_n ) capacitor c=0.00731624f \
 //x=41.81 //y=4.7 //x2=45.395 //y2=4.44
cc_3831 ( N_noxref_12_c_4745_n N_CLK_c_6190_n ) capacitor c=0.00153281f //x=37 \
 //y=2.08 //x2=36.005 //y2=4.44
cc_3832 ( N_noxref_12_c_4814_n N_CLK_c_6070_n ) capacitor c=0.014831f \
 //x=47.245 //y=3.7 //x2=64.635 //y2=4.44
cc_3833 ( N_noxref_12_c_4853_n N_CLK_c_6070_n ) capacitor c=0.0644712f \
 //x=56.125 //y=3.7 //x2=64.635 //y2=4.44
cc_3834 ( N_noxref_12_c_4855_n N_CLK_c_6070_n ) capacitor c=4.78746e-19 \
 //x=47.475 //y=3.7 //x2=64.635 //y2=4.44
cc_3835 ( N_noxref_12_c_4766_n N_CLK_c_6070_n ) capacitor c=0.0166101f \
 //x=47.36 //y=3.7 //x2=64.635 //y2=4.44
cc_3836 ( N_noxref_12_c_4748_n N_CLK_c_6070_n ) capacitor c=0.0178424f \
 //x=56.24 //y=2.08 //x2=64.635 //y2=4.44
cc_3837 ( N_noxref_12_c_4808_n N_CLK_c_6070_n ) capacitor c=0.00731624f \
 //x=56.24 //y=4.7 //x2=64.635 //y2=4.44
cc_3838 ( N_noxref_12_c_4814_n N_CLK_c_6192_n ) capacitor c=6.6036e-19 \
 //x=47.245 //y=3.7 //x2=45.625 //y2=4.44
cc_3839 ( N_noxref_12_c_4849_n N_CLK_c_6042_n ) capacitor c=0.00526349f \
 //x=37.115 //y=3.7 //x2=35.89 //y2=2.08
cc_3840 ( N_noxref_12_c_4745_n N_CLK_c_6042_n ) capacitor c=0.0402946f //x=37 \
 //y=2.08 //x2=35.89 //y2=2.08
cc_3841 ( N_noxref_12_c_4877_n N_CLK_c_6042_n ) capacitor c=0.00201097f //x=37 \
 //y=2.08 //x2=35.89 //y2=2.08
cc_3842 ( N_noxref_12_c_4806_n N_CLK_c_6042_n ) capacitor c=0.00196431f //x=37 \
 //y=4.7 //x2=35.89 //y2=2.08
cc_3843 ( N_noxref_12_c_4814_n N_CLK_c_6043_n ) capacitor c=0.0190398f \
 //x=47.245 //y=3.7 //x2=45.51 //y2=2.08
cc_3844 ( N_noxref_12_c_4752_n N_CLK_c_6043_n ) capacitor c=0.0121898f \
 //x=45.615 //y=5.155 //x2=45.51 //y2=2.08
cc_3845 ( N_noxref_12_c_4766_n N_CLK_c_6043_n ) capacitor c=0.00233004f \
 //x=47.36 //y=3.7 //x2=45.51 //y2=2.08
cc_3846 ( N_noxref_12_M106_noxref_g N_CLK_M104_noxref_g ) capacitor \
 c=0.0100903f //x=36.74 //y=6.02 //x2=35.86 //y2=6.02
cc_3847 ( N_noxref_12_M106_noxref_g N_CLK_M105_noxref_g ) capacitor \
 c=0.0600064f //x=36.74 //y=6.02 //x2=36.3 //y2=6.02
cc_3848 ( N_noxref_12_M107_noxref_g N_CLK_M105_noxref_g ) capacitor \
 c=0.0100903f //x=37.18 //y=6.02 //x2=36.3 //y2=6.02
cc_3849 ( N_noxref_12_c_4752_n N_CLK_M116_noxref_g ) capacitor c=0.0163793f \
 //x=45.615 //y=5.155 //x2=45.48 //y2=6.02
cc_3850 ( N_noxref_12_M116_noxref_d N_CLK_M116_noxref_g ) capacitor \
 c=0.0180032f //x=45.555 //y=5.02 //x2=45.48 //y2=6.02
cc_3851 ( N_noxref_12_c_4758_n N_CLK_M117_noxref_g ) capacitor c=0.0162556f \
 //x=46.495 //y=5.155 //x2=45.92 //y2=6.02
cc_3852 ( N_noxref_12_M116_noxref_d N_CLK_M117_noxref_g ) capacitor \
 c=0.0180032f //x=45.555 //y=5.02 //x2=45.92 //y2=6.02
cc_3853 ( N_noxref_12_c_4868_n N_CLK_c_6290_n ) capacitor c=0.00456962f \
 //x=36.99 //y=0.915 //x2=35.98 //y2=0.91
cc_3854 ( N_noxref_12_c_4869_n N_CLK_c_6291_n ) capacitor c=0.00438372f \
 //x=36.99 //y=1.26 //x2=35.98 //y2=1.22
cc_3855 ( N_noxref_12_c_4870_n N_CLK_c_6292_n ) capacitor c=0.00438372f \
 //x=36.99 //y=1.57 //x2=35.98 //y2=1.45
cc_3856 ( N_noxref_12_c_4745_n N_CLK_c_6293_n ) capacitor c=0.00205895f //x=37 \
 //y=2.08 //x2=35.98 //y2=1.915
cc_3857 ( N_noxref_12_c_4877_n N_CLK_c_6293_n ) capacitor c=0.00828003f //x=37 \
 //y=2.08 //x2=35.98 //y2=1.915
cc_3858 ( N_noxref_12_c_4878_n N_CLK_c_6293_n ) capacitor c=0.00438372f //x=37 \
 //y=1.915 //x2=35.98 //y2=1.915
cc_3859 ( N_noxref_12_c_4806_n N_CLK_c_6211_n ) capacitor c=0.0609323f //x=37 \
 //y=4.7 //x2=36.225 //y2=4.79
cc_3860 ( N_noxref_12_c_4957_p N_CLK_c_6212_n ) capacitor c=0.00392095f \
 //x=45.7 //y=5.155 //x2=45.845 //y2=4.79
cc_3861 ( N_noxref_12_c_4745_n N_CLK_c_6215_n ) capacitor c=0.00142741f //x=37 \
 //y=2.08 //x2=35.89 //y2=4.7
cc_3862 ( N_noxref_12_c_4806_n N_CLK_c_6215_n ) capacitor c=0.00487508f //x=37 \
 //y=4.7 //x2=35.89 //y2=4.7
cc_3863 ( N_noxref_12_c_4752_n N_CLK_c_6216_n ) capacitor c=0.00309994f \
 //x=45.615 //y=5.155 //x2=45.51 //y2=4.7
cc_3864 ( N_noxref_12_c_4745_n N_RN_c_7046_n ) capacitor c=0.0186201f //x=37 \
 //y=2.08 //x2=46.505 //y2=2.22
cc_3865 ( N_noxref_12_c_4746_n N_RN_c_7046_n ) capacitor c=0.0209607f \
 //x=41.81 //y=2.08 //x2=46.505 //y2=2.22
cc_3866 ( N_noxref_12_c_4872_n N_RN_c_7046_n ) capacitor c=3.13485e-19 \
 //x=37.365 //y=1.415 //x2=46.505 //y2=2.22
cc_3867 ( N_noxref_12_c_4833_n N_RN_c_7046_n ) capacitor c=3.13485e-19 \
 //x=42.175 //y=1.415 //x2=46.505 //y2=2.22
cc_3868 ( N_noxref_12_c_4877_n N_RN_c_7046_n ) capacitor c=0.00584491f //x=37 \
 //y=2.08 //x2=46.505 //y2=2.22
cc_3869 ( N_noxref_12_c_4838_n N_RN_c_7046_n ) capacitor c=0.00584491f \
 //x=41.81 //y=2.08 //x2=46.505 //y2=2.22
cc_3870 ( N_noxref_12_c_4853_n N_RN_c_7058_n ) capacitor c=0.00400452f \
 //x=56.125 //y=3.7 //x2=50.205 //y2=2.22
cc_3871 ( N_noxref_12_c_4968_p N_RN_c_7058_n ) capacitor c=0.016327f //x=46.96 \
 //y=1.665 //x2=50.205 //y2=2.22
cc_3872 ( N_noxref_12_c_4766_n N_RN_c_7058_n ) capacitor c=0.0220713f \
 //x=47.36 //y=3.7 //x2=50.205 //y2=2.22
cc_3873 ( N_noxref_12_c_4766_n N_RN_c_7062_n ) capacitor c=0.0012045f \
 //x=47.36 //y=3.7 //x2=46.735 //y2=2.22
cc_3874 ( N_noxref_12_c_4853_n N_RN_c_7063_n ) capacitor c=0.00433536f \
 //x=56.125 //y=3.7 //x2=59.825 //y2=2.22
cc_3875 ( N_noxref_12_c_4748_n N_RN_c_7063_n ) capacitor c=0.0186201f \
 //x=56.24 //y=2.08 //x2=59.825 //y2=2.22
cc_3876 ( N_noxref_12_c_4890_p N_RN_c_7063_n ) capacitor c=3.13485e-19 \
 //x=56.605 //y=1.415 //x2=59.825 //y2=2.22
cc_3877 ( N_noxref_12_c_4894_p N_RN_c_7063_n ) capacitor c=0.00584491f \
 //x=56.24 //y=2.08 //x2=59.825 //y2=2.22
cc_3878 ( N_noxref_12_c_4853_n N_RN_c_7070_n ) capacitor c=3.18831e-19 \
 //x=56.125 //y=3.7 //x2=50.435 //y2=2.22
cc_3879 ( N_noxref_12_c_4814_n N_RN_c_7092_n ) capacitor c=0.0179999f \
 //x=47.245 //y=3.7 //x2=46.62 //y2=2.08
cc_3880 ( N_noxref_12_c_4855_n N_RN_c_7092_n ) capacitor c=0.00179385f \
 //x=47.475 //y=3.7 //x2=46.62 //y2=2.08
cc_3881 ( N_noxref_12_c_4766_n N_RN_c_7092_n ) capacitor c=0.0757656f \
 //x=47.36 //y=3.7 //x2=46.62 //y2=2.08
cc_3882 ( N_noxref_12_c_4979_p N_RN_c_7092_n ) capacitor c=0.013297f //x=46.58 \
 //y=5.155 //x2=46.62 //y2=2.08
cc_3883 ( N_noxref_12_c_4853_n N_RN_c_7093_n ) capacitor c=0.0213788f \
 //x=56.125 //y=3.7 //x2=50.32 //y2=2.08
cc_3884 ( N_noxref_12_c_4766_n N_RN_c_7093_n ) capacitor c=5.91559e-19 \
 //x=47.36 //y=3.7 //x2=50.32 //y2=2.08
cc_3885 ( N_noxref_12_c_4758_n N_RN_M118_noxref_g ) capacitor c=0.0162556f \
 //x=46.495 //y=5.155 //x2=46.36 //y2=6.02
cc_3886 ( N_noxref_12_M118_noxref_d N_RN_M118_noxref_g ) capacitor \
 c=0.0180032f //x=46.435 //y=5.02 //x2=46.36 //y2=6.02
cc_3887 ( N_noxref_12_c_4762_n N_RN_M119_noxref_g ) capacitor c=0.0183937f \
 //x=47.275 //y=5.155 //x2=46.8 //y2=6.02
cc_3888 ( N_noxref_12_M118_noxref_d N_RN_M119_noxref_g ) capacitor \
 c=0.0194246f //x=46.435 //y=5.02 //x2=46.8 //y2=6.02
cc_3889 ( N_noxref_12_M29_noxref_d N_RN_c_7441_n ) capacitor c=0.00217566f \
 //x=46.685 //y=0.915 //x2=46.61 //y2=0.915
cc_3890 ( N_noxref_12_M29_noxref_d N_RN_c_7442_n ) capacitor c=0.0034598f \
 //x=46.685 //y=0.915 //x2=46.61 //y2=1.26
cc_3891 ( N_noxref_12_M29_noxref_d N_RN_c_7443_n ) capacitor c=0.00546784f \
 //x=46.685 //y=0.915 //x2=46.61 //y2=1.57
cc_3892 ( N_noxref_12_M29_noxref_d N_RN_c_7444_n ) capacitor c=0.00241102f \
 //x=46.685 //y=0.915 //x2=46.985 //y2=0.76
cc_3893 ( N_noxref_12_c_4747_n N_RN_c_7445_n ) capacitor c=0.00371277f \
 //x=47.275 //y=1.665 //x2=46.985 //y2=1.415
cc_3894 ( N_noxref_12_M29_noxref_d N_RN_c_7445_n ) capacitor c=0.0138621f \
 //x=46.685 //y=0.915 //x2=46.985 //y2=1.415
cc_3895 ( N_noxref_12_M29_noxref_d N_RN_c_7447_n ) capacitor c=0.00219619f \
 //x=46.685 //y=0.915 //x2=47.14 //y2=0.915
cc_3896 ( N_noxref_12_c_4747_n N_RN_c_7448_n ) capacitor c=0.00457401f \
 //x=47.275 //y=1.665 //x2=47.14 //y2=1.26
cc_3897 ( N_noxref_12_M29_noxref_d N_RN_c_7448_n ) capacitor c=0.00603828f \
 //x=46.685 //y=0.915 //x2=47.14 //y2=1.26
cc_3898 ( N_noxref_12_c_4766_n N_RN_c_7450_n ) capacitor c=0.00709342f \
 //x=47.36 //y=3.7 //x2=46.62 //y2=2.08
cc_3899 ( N_noxref_12_c_4766_n N_RN_c_7451_n ) capacitor c=0.00283672f \
 //x=47.36 //y=3.7 //x2=46.62 //y2=1.915
cc_3900 ( N_noxref_12_M29_noxref_d N_RN_c_7451_n ) capacitor c=0.00661782f \
 //x=46.685 //y=0.915 //x2=46.62 //y2=1.915
cc_3901 ( N_noxref_12_c_4762_n N_RN_c_7262_n ) capacitor c=0.00201851f \
 //x=47.275 //y=5.155 //x2=46.62 //y2=4.7
cc_3902 ( N_noxref_12_c_4766_n N_RN_c_7262_n ) capacitor c=0.0114782f \
 //x=47.36 //y=3.7 //x2=46.62 //y2=4.7
cc_3903 ( N_noxref_12_c_4979_p N_RN_c_7262_n ) capacitor c=0.00470675f \
 //x=46.58 //y=5.155 //x2=46.62 //y2=4.7
cc_3904 ( N_noxref_12_c_4809_n N_SN_c_8132_n ) capacitor c=0.0259591f \
 //x=41.695 //y=3.7 //x2=40.585 //y2=2.96
cc_3905 ( N_noxref_12_c_4849_n N_SN_c_8132_n ) capacitor c=8.32553e-19 \
 //x=37.115 //y=3.7 //x2=40.585 //y2=2.96
cc_3906 ( N_noxref_12_c_4745_n N_SN_c_8132_n ) capacitor c=0.0179917f //x=37 \
 //y=2.08 //x2=40.585 //y2=2.96
cc_3907 ( N_noxref_12_c_4809_n N_SN_c_8135_n ) capacitor c=0.0092394f \
 //x=41.695 //y=3.7 //x2=55.015 //y2=2.96
cc_3908 ( N_noxref_12_c_4814_n N_SN_c_8135_n ) capacitor c=0.041794f \
 //x=47.245 //y=3.7 //x2=55.015 //y2=2.96
cc_3909 ( N_noxref_12_c_4816_n N_SN_c_8135_n ) capacitor c=6.03896e-19 \
 //x=41.925 //y=3.7 //x2=55.015 //y2=2.96
cc_3910 ( N_noxref_12_c_4853_n N_SN_c_8135_n ) capacitor c=0.144271f \
 //x=56.125 //y=3.7 //x2=55.015 //y2=2.96
cc_3911 ( N_noxref_12_c_4855_n N_SN_c_8135_n ) capacitor c=4.80612e-19 \
 //x=47.475 //y=3.7 //x2=55.015 //y2=2.96
cc_3912 ( N_noxref_12_c_4746_n N_SN_c_8135_n ) capacitor c=0.0202855f \
 //x=41.81 //y=2.08 //x2=55.015 //y2=2.96
cc_3913 ( N_noxref_12_c_4766_n N_SN_c_8135_n ) capacitor c=0.0210712f \
 //x=47.36 //y=3.7 //x2=55.015 //y2=2.96
cc_3914 ( N_noxref_12_c_4809_n N_SN_c_8340_n ) capacitor c=6.65965e-19 \
 //x=41.695 //y=3.7 //x2=40.815 //y2=2.96
cc_3915 ( N_noxref_12_c_4746_n N_SN_c_8340_n ) capacitor c=0.00128547f \
 //x=41.81 //y=2.08 //x2=40.815 //y2=2.96
cc_3916 ( N_noxref_12_c_4853_n N_SN_c_8138_n ) capacitor c=0.0101624f \
 //x=56.125 //y=3.7 //x2=69.445 //y2=2.96
cc_3917 ( N_noxref_12_c_4748_n N_SN_c_8138_n ) capacitor c=0.0179917f \
 //x=56.24 //y=2.08 //x2=69.445 //y2=2.96
cc_3918 ( N_noxref_12_c_4853_n N_SN_c_8399_n ) capacitor c=6.65965e-19 \
 //x=56.125 //y=3.7 //x2=55.245 //y2=2.96
cc_3919 ( N_noxref_12_c_4748_n N_SN_c_8399_n ) capacitor c=0.00128547f \
 //x=56.24 //y=2.08 //x2=55.245 //y2=2.96
cc_3920 ( N_noxref_12_c_4809_n N_SN_c_8147_n ) capacitor c=0.0190398f \
 //x=41.695 //y=3.7 //x2=40.7 //y2=2.08
cc_3921 ( N_noxref_12_c_4816_n N_SN_c_8147_n ) capacitor c=0.00128547f \
 //x=41.925 //y=3.7 //x2=40.7 //y2=2.08
cc_3922 ( N_noxref_12_c_4746_n N_SN_c_8147_n ) capacitor c=0.0413563f \
 //x=41.81 //y=2.08 //x2=40.7 //y2=2.08
cc_3923 ( N_noxref_12_c_4838_n N_SN_c_8147_n ) capacitor c=0.00201097f \
 //x=41.81 //y=2.08 //x2=40.7 //y2=2.08
cc_3924 ( N_noxref_12_c_4807_n N_SN_c_8147_n ) capacitor c=0.00197875f \
 //x=41.81 //y=4.7 //x2=40.7 //y2=2.08
cc_3925 ( N_noxref_12_c_4853_n N_SN_c_8148_n ) capacitor c=0.0201805f \
 //x=56.125 //y=3.7 //x2=55.13 //y2=2.08
cc_3926 ( N_noxref_12_c_4748_n N_SN_c_8148_n ) capacitor c=0.0391831f \
 //x=56.24 //y=2.08 //x2=55.13 //y2=2.08
cc_3927 ( N_noxref_12_c_4894_p N_SN_c_8148_n ) capacitor c=0.00201097f \
 //x=56.24 //y=2.08 //x2=55.13 //y2=2.08
cc_3928 ( N_noxref_12_c_4808_n N_SN_c_8148_n ) capacitor c=0.00197875f \
 //x=56.24 //y=4.7 //x2=55.13 //y2=2.08
cc_3929 ( N_noxref_12_M112_noxref_g N_SN_M110_noxref_g ) capacitor \
 c=0.0100903f //x=41.55 //y=6.02 //x2=40.67 //y2=6.02
cc_3930 ( N_noxref_12_M112_noxref_g N_SN_M111_noxref_g ) capacitor \
 c=0.0600064f //x=41.55 //y=6.02 //x2=41.11 //y2=6.02
cc_3931 ( N_noxref_12_M113_noxref_g N_SN_M111_noxref_g ) capacitor \
 c=0.0100903f //x=41.99 //y=6.02 //x2=41.11 //y2=6.02
cc_3932 ( N_noxref_12_M130_noxref_g N_SN_M128_noxref_g ) capacitor \
 c=0.0100903f //x=55.98 //y=6.02 //x2=55.1 //y2=6.02
cc_3933 ( N_noxref_12_M130_noxref_g N_SN_M129_noxref_g ) capacitor \
 c=0.0600064f //x=55.98 //y=6.02 //x2=55.54 //y2=6.02
cc_3934 ( N_noxref_12_M131_noxref_g N_SN_M129_noxref_g ) capacitor \
 c=0.0100903f //x=56.42 //y=6.02 //x2=55.54 //y2=6.02
cc_3935 ( N_noxref_12_c_4829_n N_SN_c_8354_n ) capacitor c=0.00456962f \
 //x=41.8 //y=0.915 //x2=40.79 //y2=0.91
cc_3936 ( N_noxref_12_c_4830_n N_SN_c_8355_n ) capacitor c=0.00438372f \
 //x=41.8 //y=1.26 //x2=40.79 //y2=1.22
cc_3937 ( N_noxref_12_c_4831_n N_SN_c_8356_n ) capacitor c=0.00438372f \
 //x=41.8 //y=1.57 //x2=40.79 //y2=1.45
cc_3938 ( N_noxref_12_c_4746_n N_SN_c_8357_n ) capacitor c=0.00205895f \
 //x=41.81 //y=2.08 //x2=40.79 //y2=1.915
cc_3939 ( N_noxref_12_c_4838_n N_SN_c_8357_n ) capacitor c=0.00828003f \
 //x=41.81 //y=2.08 //x2=40.79 //y2=1.915
cc_3940 ( N_noxref_12_c_4839_n N_SN_c_8357_n ) capacitor c=0.00438372f \
 //x=41.81 //y=1.915 //x2=40.79 //y2=1.915
cc_3941 ( N_noxref_12_c_4807_n N_SN_c_8260_n ) capacitor c=0.0609323f \
 //x=41.81 //y=4.7 //x2=41.035 //y2=4.79
cc_3942 ( N_noxref_12_c_4899_p N_SN_c_8423_n ) capacitor c=0.00456962f \
 //x=56.23 //y=0.915 //x2=55.22 //y2=0.91
cc_3943 ( N_noxref_12_c_4900_p N_SN_c_8424_n ) capacitor c=0.00438372f \
 //x=56.23 //y=1.26 //x2=55.22 //y2=1.22
cc_3944 ( N_noxref_12_c_4901_p N_SN_c_8425_n ) capacitor c=0.00438372f \
 //x=56.23 //y=1.57 //x2=55.22 //y2=1.45
cc_3945 ( N_noxref_12_c_4748_n N_SN_c_8426_n ) capacitor c=0.00205895f \
 //x=56.24 //y=2.08 //x2=55.22 //y2=1.915
cc_3946 ( N_noxref_12_c_4894_p N_SN_c_8426_n ) capacitor c=0.00828003f \
 //x=56.24 //y=2.08 //x2=55.22 //y2=1.915
cc_3947 ( N_noxref_12_c_4895_p N_SN_c_8426_n ) capacitor c=0.00438372f \
 //x=56.24 //y=1.915 //x2=55.22 //y2=1.915
cc_3948 ( N_noxref_12_c_4808_n N_SN_c_8261_n ) capacitor c=0.0609323f \
 //x=56.24 //y=4.7 //x2=55.465 //y2=4.79
cc_3949 ( N_noxref_12_c_4746_n N_SN_c_8268_n ) capacitor c=0.00142741f \
 //x=41.81 //y=2.08 //x2=40.7 //y2=4.7
cc_3950 ( N_noxref_12_c_4807_n N_SN_c_8268_n ) capacitor c=0.00487508f \
 //x=41.81 //y=4.7 //x2=40.7 //y2=4.7
cc_3951 ( N_noxref_12_c_4748_n N_SN_c_8269_n ) capacitor c=0.00142741f \
 //x=56.24 //y=2.08 //x2=55.13 //y2=4.7
cc_3952 ( N_noxref_12_c_4808_n N_SN_c_8269_n ) capacitor c=0.00487508f \
 //x=56.24 //y=4.7 //x2=55.13 //y2=4.7
cc_3953 ( N_noxref_12_c_4853_n N_noxref_26_c_10048_n ) capacitor c=0.146536f \
 //x=56.125 //y=3.7 //x2=53.905 //y2=3.33
cc_3954 ( N_noxref_12_c_4853_n N_noxref_26_c_10043_n ) capacitor c=0.029467f \
 //x=56.125 //y=3.7 //x2=52.285 //y2=3.33
cc_3955 ( N_noxref_12_c_4853_n N_noxref_26_c_10050_n ) capacitor c=0.203691f \
 //x=56.125 //y=3.7 //x2=56.895 //y2=3.33
cc_3956 ( N_noxref_12_c_4748_n N_noxref_26_c_10050_n ) capacitor c=0.0198536f \
 //x=56.24 //y=2.08 //x2=56.895 //y2=3.33
cc_3957 ( N_noxref_12_c_4853_n N_noxref_26_c_10052_n ) capacitor c=0.0268338f \
 //x=56.125 //y=3.7 //x2=54.135 //y2=3.33
cc_3958 ( N_noxref_12_c_4853_n N_noxref_26_c_10053_n ) capacitor c=0.00137661f \
 //x=56.125 //y=3.7 //x2=56.98 //y2=3.615
cc_3959 ( N_noxref_12_c_4748_n N_noxref_26_c_10053_n ) capacitor c=0.00489438f \
 //x=56.24 //y=2.08 //x2=56.98 //y2=3.615
cc_3960 ( N_noxref_12_c_4853_n N_noxref_26_c_10055_n ) capacitor c=0.0145308f \
 //x=56.125 //y=3.7 //x2=57.065 //y2=3.7
cc_3961 ( N_noxref_12_c_4748_n N_noxref_26_c_10055_n ) capacitor c=4.93246e-19 \
 //x=56.24 //y=2.08 //x2=57.065 //y2=3.7
cc_3962 ( N_noxref_12_c_4762_n N_noxref_26_c_9948_n ) capacitor c=3.10026e-19 \
 //x=47.275 //y=5.155 //x2=49.715 //y2=5.155
cc_3963 ( N_noxref_12_c_4853_n N_noxref_26_c_9958_n ) capacitor c=0.0206044f \
 //x=56.125 //y=3.7 //x2=52.17 //y2=3.33
cc_3964 ( N_noxref_12_c_4853_n N_noxref_26_c_9916_n ) capacitor c=0.0216236f \
 //x=56.125 //y=3.7 //x2=54.02 //y2=2.08
cc_3965 ( N_noxref_12_c_4748_n N_noxref_26_c_9916_n ) capacitor c=0.00104576f \
 //x=56.24 //y=2.08 //x2=54.02 //y2=2.08
cc_3966 ( N_noxref_12_c_4745_n N_noxref_43_c_11310_n ) capacitor c=0.00204385f \
 //x=37 //y=2.08 //x2=37.655 //y2=0.54
cc_3967 ( N_noxref_12_c_4868_n N_noxref_43_c_11310_n ) capacitor c=0.0194423f \
 //x=36.99 //y=0.915 //x2=37.655 //y2=0.54
cc_3968 ( N_noxref_12_c_4874_n N_noxref_43_c_11310_n ) capacitor c=0.00656458f \
 //x=37.52 //y=0.915 //x2=37.655 //y2=0.54
cc_3969 ( N_noxref_12_c_4877_n N_noxref_43_c_11310_n ) capacitor c=2.20712e-19 \
 //x=37 //y=2.08 //x2=37.655 //y2=0.54
cc_3970 ( N_noxref_12_c_4869_n N_noxref_43_c_11320_n ) capacitor c=0.00538829f \
 //x=36.99 //y=1.26 //x2=36.77 //y2=0.995
cc_3971 ( N_noxref_12_c_4868_n N_noxref_43_M23_noxref_s ) capacitor \
 c=0.00538829f //x=36.99 //y=0.915 //x2=36.635 //y2=0.375
cc_3972 ( N_noxref_12_c_4870_n N_noxref_43_M23_noxref_s ) capacitor \
 c=0.00538829f //x=36.99 //y=1.57 //x2=36.635 //y2=0.375
cc_3973 ( N_noxref_12_c_4874_n N_noxref_43_M23_noxref_s ) capacitor \
 c=0.0143002f //x=37.52 //y=0.915 //x2=36.635 //y2=0.375
cc_3974 ( N_noxref_12_c_4875_n N_noxref_43_M23_noxref_s ) capacitor \
 c=0.00290153f //x=37.52 //y=1.26 //x2=36.635 //y2=0.375
cc_3975 ( N_noxref_12_c_4746_n N_noxref_45_c_11411_n ) capacitor c=0.00204385f \
 //x=41.81 //y=2.08 //x2=42.465 //y2=0.54
cc_3976 ( N_noxref_12_c_4829_n N_noxref_45_c_11411_n ) capacitor c=0.0194423f \
 //x=41.8 //y=0.915 //x2=42.465 //y2=0.54
cc_3977 ( N_noxref_12_c_4835_n N_noxref_45_c_11411_n ) capacitor c=0.00656458f \
 //x=42.33 //y=0.915 //x2=42.465 //y2=0.54
cc_3978 ( N_noxref_12_c_4838_n N_noxref_45_c_11411_n ) capacitor c=2.20712e-19 \
 //x=41.81 //y=2.08 //x2=42.465 //y2=0.54
cc_3979 ( N_noxref_12_c_4830_n N_noxref_45_c_11421_n ) capacitor c=0.00538829f \
 //x=41.8 //y=1.26 //x2=41.58 //y2=0.995
cc_3980 ( N_noxref_12_c_4829_n N_noxref_45_M26_noxref_s ) capacitor \
 c=0.00538829f //x=41.8 //y=0.915 //x2=41.445 //y2=0.375
cc_3981 ( N_noxref_12_c_4831_n N_noxref_45_M26_noxref_s ) capacitor \
 c=0.00538829f //x=41.8 //y=1.57 //x2=41.445 //y2=0.375
cc_3982 ( N_noxref_12_c_4835_n N_noxref_45_M26_noxref_s ) capacitor \
 c=0.0143002f //x=42.33 //y=0.915 //x2=41.445 //y2=0.375
cc_3983 ( N_noxref_12_c_4836_n N_noxref_45_M26_noxref_s ) capacitor \
 c=0.00290153f //x=42.33 //y=1.26 //x2=41.445 //y2=0.375
cc_3984 ( N_noxref_12_M29_noxref_d N_noxref_46_M27_noxref_s ) capacitor \
 c=0.00309936f //x=46.685 //y=0.915 //x2=43.745 //y2=0.375
cc_3985 ( N_noxref_12_c_4747_n N_noxref_47_c_11512_n ) capacitor c=0.00457167f \
 //x=47.275 //y=1.665 //x2=47.275 //y2=0.54
cc_3986 ( N_noxref_12_M29_noxref_d N_noxref_47_c_11512_n ) capacitor \
 c=0.0115903f //x=46.685 //y=0.915 //x2=47.275 //y2=0.54
cc_3987 ( N_noxref_12_c_4968_p N_noxref_47_c_11522_n ) capacitor c=0.0200405f \
 //x=46.96 //y=1.665 //x2=46.39 //y2=0.995
cc_3988 ( N_noxref_12_M29_noxref_d N_noxref_47_M28_noxref_d ) capacitor \
 c=5.27807e-19 //x=46.685 //y=0.915 //x2=45.15 //y2=0.91
cc_3989 ( N_noxref_12_c_4747_n N_noxref_47_M29_noxref_s ) capacitor \
 c=0.0196084f //x=47.275 //y=1.665 //x2=46.255 //y2=0.375
cc_3990 ( N_noxref_12_M29_noxref_d N_noxref_47_M29_noxref_s ) capacitor \
 c=0.0426368f //x=46.685 //y=0.915 //x2=46.255 //y2=0.375
cc_3991 ( N_noxref_12_c_4747_n N_noxref_48_c_11575_n ) capacitor c=3.84569e-19 \
 //x=47.275 //y=1.665 //x2=48.69 //y2=1.505
cc_3992 ( N_noxref_12_M29_noxref_d N_noxref_48_M30_noxref_s ) capacitor \
 c=2.55333e-19 //x=46.685 //y=0.915 //x2=48.555 //y2=0.375
cc_3993 ( N_noxref_12_c_4748_n N_noxref_51_c_11718_n ) capacitor c=0.00204385f \
 //x=56.24 //y=2.08 //x2=56.895 //y2=0.54
cc_3994 ( N_noxref_12_c_4899_p N_noxref_51_c_11718_n ) capacitor c=0.0194423f \
 //x=56.23 //y=0.915 //x2=56.895 //y2=0.54
cc_3995 ( N_noxref_12_c_4904_p N_noxref_51_c_11718_n ) capacitor c=0.00656458f \
 //x=56.76 //y=0.915 //x2=56.895 //y2=0.54
cc_3996 ( N_noxref_12_c_4894_p N_noxref_51_c_11718_n ) capacitor c=2.20712e-19 \
 //x=56.24 //y=2.08 //x2=56.895 //y2=0.54
cc_3997 ( N_noxref_12_c_4900_p N_noxref_51_c_11730_n ) capacitor c=0.00538829f \
 //x=56.23 //y=1.26 //x2=56.01 //y2=0.995
cc_3998 ( N_noxref_12_c_4899_p N_noxref_51_M35_noxref_s ) capacitor \
 c=0.00538829f //x=56.23 //y=0.915 //x2=55.875 //y2=0.375
cc_3999 ( N_noxref_12_c_4901_p N_noxref_51_M35_noxref_s ) capacitor \
 c=0.00538829f //x=56.23 //y=1.57 //x2=55.875 //y2=0.375
cc_4000 ( N_noxref_12_c_4904_p N_noxref_51_M35_noxref_s ) capacitor \
 c=0.0143002f //x=56.76 //y=0.915 //x2=55.875 //y2=0.375
cc_4001 ( N_noxref_12_c_4891_p N_noxref_51_M35_noxref_s ) capacitor \
 c=0.00290153f //x=56.76 //y=1.26 //x2=55.875 //y2=0.375
cc_4002 ( N_noxref_13_c_5101_n N_D_c_5328_n ) capacitor c=0.0179722f //x=51.43 \
 //y=2.08 //x2=58.715 //y2=4.07
cc_4003 ( N_noxref_13_c_5103_n N_D_c_5328_n ) capacitor c=0.0185296f //x=56.98 \
 //y=2.59 //x2=58.715 //y2=4.07
cc_4004 ( N_noxref_13_c_5103_n N_D_c_5281_n ) capacitor c=0.0105891f //x=56.98 \
 //y=2.59 //x2=58.83 //y2=2.08
cc_4005 ( N_noxref_13_c_5116_n N_noxref_15_c_5652_n ) capacitor c=3.10026e-19 \
 //x=56.895 //y=5.155 //x2=59.335 //y2=5.155
cc_4006 ( N_noxref_13_c_5101_n N_CLK_c_6070_n ) capacitor c=0.0178424f \
 //x=51.43 //y=2.08 //x2=64.635 //y2=4.44
cc_4007 ( N_noxref_13_c_5103_n N_CLK_c_6070_n ) capacitor c=0.0166101f \
 //x=56.98 //y=2.59 //x2=64.635 //y2=4.44
cc_4008 ( N_noxref_13_c_5145_n N_CLK_c_6070_n ) capacitor c=0.00731624f \
 //x=51.43 //y=4.7 //x2=64.635 //y2=4.44
cc_4009 ( N_noxref_13_c_5099_n N_RN_c_7063_n ) capacitor c=0.491184f \
 //x=56.865 //y=2.59 //x2=59.825 //y2=2.22
cc_4010 ( N_noxref_13_c_5149_n N_RN_c_7063_n ) capacitor c=0.0289738f \
 //x=51.545 //y=2.59 //x2=59.825 //y2=2.22
cc_4011 ( N_noxref_13_c_5101_n N_RN_c_7063_n ) capacitor c=0.0204547f \
 //x=51.43 //y=2.08 //x2=59.825 //y2=2.22
cc_4012 ( N_noxref_13_c_5183_p N_RN_c_7063_n ) capacitor c=0.016327f //x=56.58 \
 //y=1.665 //x2=59.825 //y2=2.22
cc_4013 ( N_noxref_13_c_5103_n N_RN_c_7063_n ) capacitor c=0.0215653f \
 //x=56.98 //y=2.59 //x2=59.825 //y2=2.22
cc_4014 ( N_noxref_13_c_5185_p N_RN_c_7063_n ) capacitor c=3.13485e-19 \
 //x=51.795 //y=1.415 //x2=59.825 //y2=2.22
cc_4015 ( N_noxref_13_c_5186_p N_RN_c_7063_n ) capacitor c=0.00584491f \
 //x=51.43 //y=2.08 //x2=59.825 //y2=2.22
cc_4016 ( N_noxref_13_c_5101_n N_RN_c_7070_n ) capacitor c=0.00165648f \
 //x=51.43 //y=2.08 //x2=50.435 //y2=2.22
cc_4017 ( N_noxref_13_c_5186_p N_RN_c_7070_n ) capacitor c=2.3323e-19 \
 //x=51.43 //y=2.08 //x2=50.435 //y2=2.22
cc_4018 ( N_noxref_13_c_5149_n N_RN_c_7093_n ) capacitor c=0.00526349f \
 //x=51.545 //y=2.59 //x2=50.32 //y2=2.08
cc_4019 ( N_noxref_13_c_5101_n N_RN_c_7093_n ) capacitor c=0.042257f //x=51.43 \
 //y=2.08 //x2=50.32 //y2=2.08
cc_4020 ( N_noxref_13_c_5186_p N_RN_c_7093_n ) capacitor c=0.0019893f \
 //x=51.43 //y=2.08 //x2=50.32 //y2=2.08
cc_4021 ( N_noxref_13_c_5145_n N_RN_c_7093_n ) capacitor c=0.00197875f \
 //x=51.43 //y=4.7 //x2=50.32 //y2=2.08
cc_4022 ( N_noxref_13_c_5103_n N_RN_c_7094_n ) capacitor c=8.03384e-19 \
 //x=56.98 //y=2.59 //x2=59.94 //y2=2.08
cc_4023 ( N_noxref_13_M124_noxref_g N_RN_M122_noxref_g ) capacitor \
 c=0.0100903f //x=51.17 //y=6.02 //x2=50.29 //y2=6.02
cc_4024 ( N_noxref_13_M124_noxref_g N_RN_M123_noxref_g ) capacitor \
 c=0.0600064f //x=51.17 //y=6.02 //x2=50.73 //y2=6.02
cc_4025 ( N_noxref_13_M125_noxref_g N_RN_M123_noxref_g ) capacitor \
 c=0.0100903f //x=51.61 //y=6.02 //x2=50.73 //y2=6.02
cc_4026 ( N_noxref_13_c_5197_p N_RN_c_7406_n ) capacitor c=0.00456962f \
 //x=51.42 //y=0.915 //x2=50.41 //y2=0.91
cc_4027 ( N_noxref_13_c_5198_p N_RN_c_7407_n ) capacitor c=0.00438372f \
 //x=51.42 //y=1.26 //x2=50.41 //y2=1.22
cc_4028 ( N_noxref_13_c_5199_p N_RN_c_7408_n ) capacitor c=0.00438372f \
 //x=51.42 //y=1.57 //x2=50.41 //y2=1.45
cc_4029 ( N_noxref_13_c_5101_n N_RN_c_7409_n ) capacitor c=0.00205895f \
 //x=51.43 //y=2.08 //x2=50.41 //y2=1.915
cc_4030 ( N_noxref_13_c_5186_p N_RN_c_7409_n ) capacitor c=0.00828003f \
 //x=51.43 //y=2.08 //x2=50.41 //y2=1.915
cc_4031 ( N_noxref_13_c_5202_p N_RN_c_7409_n ) capacitor c=0.00438372f \
 //x=51.43 //y=1.915 //x2=50.41 //y2=1.915
cc_4032 ( N_noxref_13_c_5145_n N_RN_c_7257_n ) capacitor c=0.0609323f \
 //x=51.43 //y=4.7 //x2=50.655 //y2=4.79
cc_4033 ( N_noxref_13_c_5101_n N_RN_c_7263_n ) capacitor c=0.00142741f \
 //x=51.43 //y=2.08 //x2=50.32 //y2=4.7
cc_4034 ( N_noxref_13_c_5145_n N_RN_c_7263_n ) capacitor c=0.00487508f \
 //x=51.43 //y=4.7 //x2=50.32 //y2=4.7
cc_4035 ( N_noxref_13_c_5099_n N_SN_c_8135_n ) capacitor c=0.303889f \
 //x=56.865 //y=2.59 //x2=55.015 //y2=2.96
cc_4036 ( N_noxref_13_c_5149_n N_SN_c_8135_n ) capacitor c=0.0291665f \
 //x=51.545 //y=2.59 //x2=55.015 //y2=2.96
cc_4037 ( N_noxref_13_c_5101_n N_SN_c_8135_n ) capacitor c=0.0221691f \
 //x=51.43 //y=2.08 //x2=55.015 //y2=2.96
cc_4038 ( N_noxref_13_c_5099_n N_SN_c_8138_n ) capacitor c=0.170173f \
 //x=56.865 //y=2.59 //x2=69.445 //y2=2.96
cc_4039 ( N_noxref_13_c_5103_n N_SN_c_8138_n ) capacitor c=0.0205746f \
 //x=56.98 //y=2.59 //x2=69.445 //y2=2.96
cc_4040 ( N_noxref_13_c_5099_n N_SN_c_8399_n ) capacitor c=0.0264232f \
 //x=56.865 //y=2.59 //x2=55.245 //y2=2.96
cc_4041 ( N_noxref_13_c_5099_n N_SN_c_8148_n ) capacitor c=0.0208352f \
 //x=56.865 //y=2.59 //x2=55.13 //y2=2.08
cc_4042 ( N_noxref_13_c_5106_n N_SN_c_8148_n ) capacitor c=0.0121898f \
 //x=55.235 //y=5.155 //x2=55.13 //y2=2.08
cc_4043 ( N_noxref_13_c_5103_n N_SN_c_8148_n ) capacitor c=0.00200263f \
 //x=56.98 //y=2.59 //x2=55.13 //y2=2.08
cc_4044 ( N_noxref_13_c_5106_n N_SN_M128_noxref_g ) capacitor c=0.0163793f \
 //x=55.235 //y=5.155 //x2=55.1 //y2=6.02
cc_4045 ( N_noxref_13_M128_noxref_d N_SN_M128_noxref_g ) capacitor \
 c=0.0180032f //x=55.175 //y=5.02 //x2=55.1 //y2=6.02
cc_4046 ( N_noxref_13_c_5112_n N_SN_M129_noxref_g ) capacitor c=0.0162556f \
 //x=56.115 //y=5.155 //x2=55.54 //y2=6.02
cc_4047 ( N_noxref_13_M128_noxref_d N_SN_M129_noxref_g ) capacitor \
 c=0.0180032f //x=55.175 //y=5.02 //x2=55.54 //y2=6.02
cc_4048 ( N_noxref_13_c_5219_p N_SN_c_8261_n ) capacitor c=0.00392095f \
 //x=55.32 //y=5.155 //x2=55.465 //y2=4.79
cc_4049 ( N_noxref_13_c_5106_n N_SN_c_8269_n ) capacitor c=0.00309994f \
 //x=55.235 //y=5.155 //x2=55.13 //y2=4.7
cc_4050 ( N_noxref_13_c_5099_n N_noxref_26_c_10048_n ) capacitor c=0.0111324f \
 //x=56.865 //y=2.59 //x2=53.905 //y2=3.33
cc_4051 ( N_noxref_13_c_5099_n N_noxref_26_c_10043_n ) capacitor c=8.93831e-19 \
 //x=56.865 //y=2.59 //x2=52.285 //y2=3.33
cc_4052 ( N_noxref_13_c_5101_n N_noxref_26_c_10043_n ) capacitor c=0.0044695f \
 //x=51.43 //y=2.08 //x2=52.285 //y2=3.33
cc_4053 ( N_noxref_13_c_5099_n N_noxref_26_c_10050_n ) capacitor c=0.025f \
 //x=56.865 //y=2.59 //x2=56.895 //y2=3.33
cc_4054 ( N_noxref_13_c_5103_n N_noxref_26_c_10050_n ) capacitor c=0.0140629f \
 //x=56.98 //y=2.59 //x2=56.895 //y2=3.33
cc_4055 ( N_noxref_13_c_5099_n N_noxref_26_c_10052_n ) capacitor c=5.41495e-19 \
 //x=56.865 //y=2.59 //x2=54.135 //y2=3.33
cc_4056 ( N_noxref_13_c_5103_n N_noxref_26_c_10053_n ) capacitor c=0.0100064f \
 //x=56.98 //y=2.59 //x2=56.98 //y2=3.615
cc_4057 ( N_noxref_13_c_5103_n N_noxref_26_c_10055_n ) capacitor c=0.0133081f \
 //x=56.98 //y=2.59 //x2=57.065 //y2=3.7
cc_4058 ( N_noxref_13_M124_noxref_g N_noxref_26_c_9950_n ) capacitor \
 c=0.0162556f //x=51.17 //y=6.02 //x2=51.305 //y2=5.155
cc_4059 ( N_noxref_13_c_5110_n N_noxref_26_c_9954_n ) capacitor c=3.10026e-19 \
 //x=54.525 //y=5.155 //x2=52.085 //y2=5.155
cc_4060 ( N_noxref_13_M125_noxref_g N_noxref_26_c_9954_n ) capacitor \
 c=0.0183937f //x=51.61 //y=6.02 //x2=52.085 //y2=5.155
cc_4061 ( N_noxref_13_c_5145_n N_noxref_26_c_9954_n ) capacitor c=0.00201851f \
 //x=51.43 //y=4.7 //x2=52.085 //y2=5.155
cc_4062 ( N_noxref_13_c_5185_p N_noxref_26_c_9915_n ) capacitor c=0.00371277f \
 //x=51.795 //y=1.415 //x2=52.085 //y2=1.665
cc_4063 ( N_noxref_13_c_5234_p N_noxref_26_c_9915_n ) capacitor c=0.00457401f \
 //x=51.95 //y=1.26 //x2=52.085 //y2=1.665
cc_4064 ( N_noxref_13_c_5099_n N_noxref_26_c_9958_n ) capacitor c=0.0165903f \
 //x=56.865 //y=2.59 //x2=52.17 //y2=3.33
cc_4065 ( N_noxref_13_c_5149_n N_noxref_26_c_9958_n ) capacitor c=0.00179385f \
 //x=51.545 //y=2.59 //x2=52.17 //y2=3.33
cc_4066 ( N_noxref_13_c_5101_n N_noxref_26_c_9958_n ) capacitor c=0.0751342f \
 //x=51.43 //y=2.08 //x2=52.17 //y2=3.33
cc_4067 ( N_noxref_13_c_5186_p N_noxref_26_c_9958_n ) capacitor c=0.00709342f \
 //x=51.43 //y=2.08 //x2=52.17 //y2=3.33
cc_4068 ( N_noxref_13_c_5202_p N_noxref_26_c_9958_n ) capacitor c=0.00283672f \
 //x=51.43 //y=1.915 //x2=52.17 //y2=3.33
cc_4069 ( N_noxref_13_c_5145_n N_noxref_26_c_9958_n ) capacitor c=0.0116291f \
 //x=51.43 //y=4.7 //x2=52.17 //y2=3.33
cc_4070 ( N_noxref_13_c_5099_n N_noxref_26_c_9916_n ) capacitor c=0.0188253f \
 //x=56.865 //y=2.59 //x2=54.02 //y2=2.08
cc_4071 ( N_noxref_13_c_5101_n N_noxref_26_c_9916_n ) capacitor c=8.50231e-19 \
 //x=51.43 //y=2.08 //x2=54.02 //y2=2.08
cc_4072 ( N_noxref_13_c_5101_n N_noxref_26_c_10083_n ) capacitor c=0.013297f \
 //x=51.43 //y=2.08 //x2=51.39 //y2=5.155
cc_4073 ( N_noxref_13_c_5145_n N_noxref_26_c_10083_n ) capacitor c=0.00470675f \
 //x=51.43 //y=4.7 //x2=51.39 //y2=5.155
cc_4074 ( N_noxref_13_c_5110_n N_noxref_26_M126_noxref_g ) capacitor \
 c=0.0213876f //x=54.525 //y=5.155 //x2=54.22 //y2=6.02
cc_4075 ( N_noxref_13_c_5106_n N_noxref_26_M127_noxref_g ) capacitor \
 c=0.0157304f //x=55.235 //y=5.155 //x2=54.66 //y2=6.02
cc_4076 ( N_noxref_13_M126_noxref_d N_noxref_26_M127_noxref_g ) capacitor \
 c=0.0180032f //x=54.295 //y=5.02 //x2=54.66 //y2=6.02
cc_4077 ( N_noxref_13_c_5110_n N_noxref_26_c_10024_n ) capacitor c=0.00393496f \
 //x=54.525 //y=5.155 //x2=54.585 //y2=4.79
cc_4078 ( N_noxref_13_c_5197_p N_noxref_26_M32_noxref_d ) capacitor \
 c=0.00217566f //x=51.42 //y=0.915 //x2=51.495 //y2=0.915
cc_4079 ( N_noxref_13_c_5198_p N_noxref_26_M32_noxref_d ) capacitor \
 c=0.0034598f //x=51.42 //y=1.26 //x2=51.495 //y2=0.915
cc_4080 ( N_noxref_13_c_5199_p N_noxref_26_M32_noxref_d ) capacitor \
 c=0.00546784f //x=51.42 //y=1.57 //x2=51.495 //y2=0.915
cc_4081 ( N_noxref_13_c_5252_p N_noxref_26_M32_noxref_d ) capacitor \
 c=0.00241102f //x=51.795 //y=0.76 //x2=51.495 //y2=0.915
cc_4082 ( N_noxref_13_c_5185_p N_noxref_26_M32_noxref_d ) capacitor \
 c=0.0138621f //x=51.795 //y=1.415 //x2=51.495 //y2=0.915
cc_4083 ( N_noxref_13_c_5254_p N_noxref_26_M32_noxref_d ) capacitor \
 c=0.00219619f //x=51.95 //y=0.915 //x2=51.495 //y2=0.915
cc_4084 ( N_noxref_13_c_5234_p N_noxref_26_M32_noxref_d ) capacitor \
 c=0.00603828f //x=51.95 //y=1.26 //x2=51.495 //y2=0.915
cc_4085 ( N_noxref_13_c_5202_p N_noxref_26_M32_noxref_d ) capacitor \
 c=0.00661782f //x=51.43 //y=1.915 //x2=51.495 //y2=0.915
cc_4086 ( N_noxref_13_M124_noxref_g N_noxref_26_M124_noxref_d ) capacitor \
 c=0.0180032f //x=51.17 //y=6.02 //x2=51.245 //y2=5.02
cc_4087 ( N_noxref_13_M125_noxref_g N_noxref_26_M124_noxref_d ) capacitor \
 c=0.0194246f //x=51.61 //y=6.02 //x2=51.245 //y2=5.02
cc_4088 ( N_noxref_13_c_5101_n N_noxref_49_c_11617_n ) capacitor c=0.00204385f \
 //x=51.43 //y=2.08 //x2=52.085 //y2=0.54
cc_4089 ( N_noxref_13_c_5197_p N_noxref_49_c_11617_n ) capacitor c=0.0194423f \
 //x=51.42 //y=0.915 //x2=52.085 //y2=0.54
cc_4090 ( N_noxref_13_c_5254_p N_noxref_49_c_11617_n ) capacitor c=0.00656458f \
 //x=51.95 //y=0.915 //x2=52.085 //y2=0.54
cc_4091 ( N_noxref_13_c_5186_p N_noxref_49_c_11617_n ) capacitor c=2.20712e-19 \
 //x=51.43 //y=2.08 //x2=52.085 //y2=0.54
cc_4092 ( N_noxref_13_c_5198_p N_noxref_49_c_11629_n ) capacitor c=0.00538829f \
 //x=51.42 //y=1.26 //x2=51.2 //y2=0.995
cc_4093 ( N_noxref_13_c_5197_p N_noxref_49_M32_noxref_s ) capacitor \
 c=0.00538829f //x=51.42 //y=0.915 //x2=51.065 //y2=0.375
cc_4094 ( N_noxref_13_c_5199_p N_noxref_49_M32_noxref_s ) capacitor \
 c=0.00538829f //x=51.42 //y=1.57 //x2=51.065 //y2=0.375
cc_4095 ( N_noxref_13_c_5254_p N_noxref_49_M32_noxref_s ) capacitor \
 c=0.0143002f //x=51.95 //y=0.915 //x2=51.065 //y2=0.375
cc_4096 ( N_noxref_13_c_5234_p N_noxref_49_M32_noxref_s ) capacitor \
 c=0.00290153f //x=51.95 //y=1.26 //x2=51.065 //y2=0.375
cc_4097 ( N_noxref_13_M35_noxref_d N_noxref_50_M33_noxref_s ) capacitor \
 c=0.00309936f //x=56.305 //y=0.915 //x2=53.365 //y2=0.375
cc_4098 ( N_noxref_13_c_5102_n N_noxref_51_c_11718_n ) capacitor c=0.00457167f \
 //x=56.895 //y=1.665 //x2=56.895 //y2=0.54
cc_4099 ( N_noxref_13_M35_noxref_d N_noxref_51_c_11718_n ) capacitor \
 c=0.0115903f //x=56.305 //y=0.915 //x2=56.895 //y2=0.54
cc_4100 ( N_noxref_13_c_5183_p N_noxref_51_c_11730_n ) capacitor c=0.0200405f \
 //x=56.58 //y=1.665 //x2=56.01 //y2=0.995
cc_4101 ( N_noxref_13_M35_noxref_d N_noxref_51_M34_noxref_d ) capacitor \
 c=5.27807e-19 //x=56.305 //y=0.915 //x2=54.77 //y2=0.91
cc_4102 ( N_noxref_13_c_5102_n N_noxref_51_M35_noxref_s ) capacitor \
 c=0.0184051f //x=56.895 //y=1.665 //x2=55.875 //y2=0.375
cc_4103 ( N_noxref_13_M35_noxref_d N_noxref_51_M35_noxref_s ) capacitor \
 c=0.0426368f //x=56.305 //y=0.915 //x2=55.875 //y2=0.375
cc_4104 ( N_noxref_13_c_5102_n N_noxref_52_c_11780_n ) capacitor c=3.84569e-19 \
 //x=56.895 //y=1.665 //x2=58.31 //y2=1.505
cc_4105 ( N_noxref_13_M35_noxref_d N_noxref_52_M36_noxref_s ) capacitor \
 c=2.55333e-19 //x=56.305 //y=0.915 //x2=58.175 //y2=0.375
cc_4106 ( N_D_M133_noxref_g N_noxref_15_c_5648_n ) capacitor c=0.0157304f \
 //x=59.47 //y=6.02 //x2=60.045 //y2=5.155
cc_4107 ( N_D_M132_noxref_g N_noxref_15_c_5652_n ) capacitor c=0.0213876f \
 //x=59.03 //y=6.02 //x2=59.335 //y2=5.155
cc_4108 ( N_D_c_5402_n N_noxref_15_c_5652_n ) capacitor c=0.00393496f \
 //x=59.395 //y=4.79 //x2=59.335 //y2=5.155
cc_4109 ( N_D_M133_noxref_g N_noxref_15_M132_noxref_d ) capacitor c=0.0180032f \
 //x=59.47 //y=6.02 //x2=59.105 //y2=5.02
cc_4110 ( N_D_c_5277_n N_CLK_c_6046_n ) capacitor c=0.816492f //x=29.855 \
 //y=4.07 //x2=16.535 //y2=4.44
cc_4111 ( N_D_c_5277_n N_CLK_c_6057_n ) capacitor c=0.0291328f //x=29.855 \
 //y=4.07 //x2=7.145 //y2=4.44
cc_4112 ( N_D_c_5277_n N_CLK_c_6058_n ) capacitor c=1.13884f //x=29.855 \
 //y=4.07 //x2=35.775 //y2=4.44
cc_4113 ( N_D_c_5328_n N_CLK_c_6058_n ) capacitor c=0.494146f //x=58.715 \
 //y=4.07 //x2=35.775 //y2=4.44
cc_4114 ( N_D_c_5334_n N_CLK_c_6058_n ) capacitor c=0.0263777f //x=30.085 \
 //y=4.07 //x2=35.775 //y2=4.44
cc_4115 ( N_D_c_5280_n N_CLK_c_6058_n ) capacitor c=0.0206206f //x=29.97 \
 //y=2.08 //x2=35.775 //y2=4.44
cc_4116 ( N_D_c_5358_n N_CLK_c_6058_n ) capacitor c=0.0112124f //x=30.245 \
 //y=4.79 //x2=35.775 //y2=4.44
cc_4117 ( N_D_c_5277_n N_CLK_c_6067_n ) capacitor c=0.026534f //x=29.855 \
 //y=4.07 //x2=16.765 //y2=4.44
cc_4118 ( N_D_c_5328_n N_CLK_c_6068_n ) capacitor c=0.816492f //x=58.715 \
 //y=4.07 //x2=45.395 //y2=4.44
cc_4119 ( N_D_c_5328_n N_CLK_c_6190_n ) capacitor c=0.026534f //x=58.715 \
 //y=4.07 //x2=36.005 //y2=4.44
cc_4120 ( N_D_c_5328_n N_CLK_c_6070_n ) capacitor c=1.16782f //x=58.715 \
 //y=4.07 //x2=64.635 //y2=4.44
cc_4121 ( N_D_c_5281_n N_CLK_c_6070_n ) capacitor c=0.0206206f //x=58.83 \
 //y=2.08 //x2=64.635 //y2=4.44
cc_4122 ( N_D_c_5360_n N_CLK_c_6070_n ) capacitor c=0.0112124f //x=59.105 \
 //y=4.79 //x2=64.635 //y2=4.44
cc_4123 ( N_D_c_5328_n N_CLK_c_6192_n ) capacitor c=0.026534f //x=58.715 \
 //y=4.07 //x2=45.625 //y2=4.44
cc_4124 ( N_D_c_5277_n N_CLK_c_6040_n ) capacitor c=0.0231929f //x=29.855 \
 //y=4.07 //x2=7.03 //y2=2.08
cc_4125 ( N_D_c_5277_n N_CLK_c_6041_n ) capacitor c=0.0208526f //x=29.855 \
 //y=4.07 //x2=16.65 //y2=2.08
cc_4126 ( N_D_c_5328_n N_CLK_c_6042_n ) capacitor c=0.0231929f //x=58.715 \
 //y=4.07 //x2=35.89 //y2=2.08
cc_4127 ( N_D_c_5328_n N_CLK_c_6043_n ) capacitor c=0.0208526f //x=58.715 \
 //y=4.07 //x2=45.51 //y2=2.08
cc_4128 ( N_D_c_5281_n N_noxref_18_c_6747_n ) capacitor c=0.001514f //x=58.83 \
 //y=2.08 //x2=61.05 //y2=2.08
cc_4129 ( N_D_c_5277_n N_RN_c_7021_n ) capacitor c=0.017478f //x=29.855 \
 //y=4.07 //x2=17.645 //y2=2.22
cc_4130 ( N_D_c_5277_n N_RN_c_7032_n ) capacitor c=0.00393113f //x=29.855 \
 //y=4.07 //x2=2.335 //y2=2.22
cc_4131 ( N_D_c_5279_n N_RN_c_7032_n ) capacitor c=0.00558344f //x=1.11 \
 //y=2.08 //x2=2.335 //y2=2.22
cc_4132 ( N_D_c_5286_n N_RN_c_7032_n ) capacitor c=0.00341397f //x=0.81 \
 //y=1.915 //x2=2.335 //y2=2.22
cc_4133 ( N_D_c_5277_n N_RN_c_7038_n ) capacitor c=0.00236788f //x=29.855 \
 //y=4.07 //x2=30.965 //y2=2.22
cc_4134 ( N_D_c_5328_n N_RN_c_7038_n ) capacitor c=0.00333858f //x=58.715 \
 //y=4.07 //x2=30.965 //y2=2.22
cc_4135 ( N_D_c_5280_n N_RN_c_7038_n ) capacitor c=0.0216101f //x=29.97 \
 //y=2.08 //x2=30.965 //y2=2.22
cc_4136 ( N_D_c_5296_n N_RN_c_7038_n ) capacitor c=0.011987f //x=29.67 \
 //y=1.915 //x2=30.965 //y2=2.22
cc_4137 ( N_D_c_5328_n N_RN_c_7046_n ) capacitor c=0.00359237f //x=58.715 \
 //y=4.07 //x2=46.505 //y2=2.22
cc_4138 ( N_D_c_5328_n N_RN_c_7057_n ) capacitor c=2.66524e-19 //x=58.715 \
 //y=4.07 //x2=31.195 //y2=2.22
cc_4139 ( N_D_c_5280_n N_RN_c_7057_n ) capacitor c=0.00165648f //x=29.97 \
 //y=2.08 //x2=31.195 //y2=2.22
cc_4140 ( N_D_c_5296_n N_RN_c_7057_n ) capacitor c=2.3323e-19 //x=29.67 \
 //y=1.915 //x2=31.195 //y2=2.22
cc_4141 ( N_D_c_5281_n N_RN_c_7063_n ) capacitor c=0.0216101f //x=58.83 \
 //y=2.08 //x2=59.825 //y2=2.22
cc_4142 ( N_D_c_5306_n N_RN_c_7063_n ) capacitor c=0.011987f //x=58.53 \
 //y=1.915 //x2=59.825 //y2=2.22
cc_4143 ( N_D_c_5281_n N_RN_c_7082_n ) capacitor c=0.00165648f //x=58.83 \
 //y=2.08 //x2=60.055 //y2=2.22
cc_4144 ( N_D_c_5306_n N_RN_c_7082_n ) capacitor c=2.3323e-19 //x=58.53 \
 //y=1.915 //x2=60.055 //y2=2.22
cc_4145 ( N_D_c_5277_n N_RN_c_7088_n ) capacitor c=0.0283962f //x=29.855 \
 //y=4.07 //x2=2.22 //y2=2.08
cc_4146 ( N_D_c_5278_n N_RN_c_7088_n ) capacitor c=0.00128547f //x=1.225 \
 //y=4.07 //x2=2.22 //y2=2.08
cc_4147 ( N_D_c_5279_n N_RN_c_7088_n ) capacitor c=0.0536972f //x=1.11 \
 //y=2.08 //x2=2.22 //y2=2.08
cc_4148 ( N_D_c_5286_n N_RN_c_7088_n ) capacitor c=0.00228225f //x=0.81 \
 //y=1.915 //x2=2.22 //y2=2.08
cc_4149 ( N_D_c_5376_n N_RN_c_7088_n ) capacitor c=0.00147352f //x=1.675 \
 //y=4.79 //x2=2.22 //y2=2.08
cc_4150 ( N_D_c_5356_n N_RN_c_7088_n ) capacitor c=0.00142741f //x=1.385 \
 //y=4.79 //x2=2.22 //y2=2.08
cc_4151 ( N_D_c_5277_n N_RN_c_7089_n ) capacitor c=0.0179722f //x=29.855 \
 //y=4.07 //x2=17.76 //y2=2.08
cc_4152 ( N_D_c_5277_n N_RN_c_7090_n ) capacitor c=0.0190126f //x=29.855 \
 //y=4.07 //x2=21.46 //y2=2.08
cc_4153 ( N_D_c_5328_n N_RN_c_7091_n ) capacitor c=0.0228716f //x=58.715 \
 //y=4.07 //x2=31.08 //y2=2.08
cc_4154 ( N_D_c_5334_n N_RN_c_7091_n ) capacitor c=0.00128547f //x=30.085 \
 //y=4.07 //x2=31.08 //y2=2.08
cc_4155 ( N_D_c_5280_n N_RN_c_7091_n ) capacitor c=0.0459779f //x=29.97 \
 //y=2.08 //x2=31.08 //y2=2.08
cc_4156 ( N_D_c_5296_n N_RN_c_7091_n ) capacitor c=0.00208635f //x=29.67 \
 //y=1.915 //x2=31.08 //y2=2.08
cc_4157 ( N_D_c_5400_n N_RN_c_7091_n ) capacitor c=0.00120758f //x=30.535 \
 //y=4.79 //x2=31.08 //y2=2.08
cc_4158 ( N_D_c_5358_n N_RN_c_7091_n ) capacitor c=0.00142741f //x=30.245 \
 //y=4.79 //x2=31.08 //y2=2.08
cc_4159 ( N_D_c_5328_n N_RN_c_7092_n ) capacitor c=0.0179722f //x=58.715 \
 //y=4.07 //x2=46.62 //y2=2.08
cc_4160 ( N_D_c_5328_n N_RN_c_7093_n ) capacitor c=0.0190126f //x=58.715 \
 //y=4.07 //x2=50.32 //y2=2.08
cc_4161 ( N_D_c_5328_n N_RN_c_7094_n ) capacitor c=0.00526349f //x=58.715 \
 //y=4.07 //x2=59.94 //y2=2.08
cc_4162 ( N_D_c_5281_n N_RN_c_7094_n ) capacitor c=0.0440868f //x=58.83 \
 //y=2.08 //x2=59.94 //y2=2.08
cc_4163 ( N_D_c_5306_n N_RN_c_7094_n ) capacitor c=0.00208635f //x=58.53 \
 //y=1.915 //x2=59.94 //y2=2.08
cc_4164 ( N_D_c_5402_n N_RN_c_7094_n ) capacitor c=0.00120758f //x=59.395 \
 //y=4.79 //x2=59.94 //y2=2.08
cc_4165 ( N_D_c_5360_n N_RN_c_7094_n ) capacitor c=0.00142741f //x=59.105 \
 //y=4.79 //x2=59.94 //y2=2.08
cc_4166 ( N_D_M60_noxref_g N_RN_M62_noxref_g ) capacitor c=0.0105869f //x=1.31 \
 //y=6.02 //x2=2.19 //y2=6.02
cc_4167 ( N_D_M61_noxref_g N_RN_M62_noxref_g ) capacitor c=0.10632f //x=1.75 \
 //y=6.02 //x2=2.19 //y2=6.02
cc_4168 ( N_D_M61_noxref_g N_RN_M63_noxref_g ) capacitor c=0.0101598f //x=1.75 \
 //y=6.02 //x2=2.63 //y2=6.02
cc_4169 ( N_D_M96_noxref_g N_RN_M98_noxref_g ) capacitor c=0.0105174f \
 //x=30.17 //y=6.02 //x2=31.05 //y2=6.02
cc_4170 ( N_D_M97_noxref_g N_RN_M98_noxref_g ) capacitor c=0.10624f //x=30.61 \
 //y=6.02 //x2=31.05 //y2=6.02
cc_4171 ( N_D_M97_noxref_g N_RN_M99_noxref_g ) capacitor c=0.0100903f \
 //x=30.61 //y=6.02 //x2=31.49 //y2=6.02
cc_4172 ( N_D_M132_noxref_g N_RN_M134_noxref_g ) capacitor c=0.0105174f \
 //x=59.03 //y=6.02 //x2=59.91 //y2=6.02
cc_4173 ( N_D_M133_noxref_g N_RN_M134_noxref_g ) capacitor c=0.10624f \
 //x=59.47 //y=6.02 //x2=59.91 //y2=6.02
cc_4174 ( N_D_M133_noxref_g N_RN_M135_noxref_g ) capacitor c=0.0100903f \
 //x=59.47 //y=6.02 //x2=60.35 //y2=6.02
cc_4175 ( N_D_c_5282_n N_RN_c_7528_n ) capacitor c=5.72482e-19 //x=0.81 \
 //y=0.875 //x2=1.785 //y2=0.91
cc_4176 ( N_D_c_5284_n N_RN_c_7528_n ) capacitor c=0.00149976f //x=0.81 \
 //y=1.22 //x2=1.785 //y2=0.91
cc_4177 ( N_D_c_5289_n N_RN_c_7528_n ) capacitor c=0.0160123f //x=1.34 \
 //y=0.875 //x2=1.785 //y2=0.91
cc_4178 ( N_D_c_5285_n N_RN_c_7531_n ) capacitor c=0.00111227f //x=0.81 \
 //y=1.53 //x2=1.785 //y2=1.22
cc_4179 ( N_D_c_5291_n N_RN_c_7531_n ) capacitor c=0.0124075f //x=1.34 \
 //y=1.22 //x2=1.785 //y2=1.22
cc_4180 ( N_D_c_5289_n N_RN_c_7204_n ) capacitor c=0.00103227f //x=1.34 \
 //y=0.875 //x2=2.31 //y2=0.91
cc_4181 ( N_D_c_5291_n N_RN_c_7205_n ) capacitor c=0.0010154f //x=1.34 \
 //y=1.22 //x2=2.31 //y2=1.22
cc_4182 ( N_D_c_5291_n N_RN_c_7206_n ) capacitor c=9.23422e-19 //x=1.34 \
 //y=1.22 //x2=2.31 //y2=1.45
cc_4183 ( N_D_c_5279_n N_RN_c_7207_n ) capacitor c=0.00211714f //x=1.11 \
 //y=2.08 //x2=2.31 //y2=1.915
cc_4184 ( N_D_c_5286_n N_RN_c_7207_n ) capacitor c=0.00909574f //x=0.81 \
 //y=1.915 //x2=2.31 //y2=1.915
cc_4185 ( N_D_c_5277_n N_RN_c_7161_n ) capacitor c=0.00495688f //x=29.855 \
 //y=4.07 //x2=2.555 //y2=4.79
cc_4186 ( N_D_c_5292_n N_RN_c_7539_n ) capacitor c=5.72482e-19 //x=29.67 \
 //y=0.875 //x2=30.645 //y2=0.91
cc_4187 ( N_D_c_5294_n N_RN_c_7539_n ) capacitor c=0.00149976f //x=29.67 \
 //y=1.22 //x2=30.645 //y2=0.91
cc_4188 ( N_D_c_5299_n N_RN_c_7539_n ) capacitor c=0.0160123f //x=30.2 \
 //y=0.875 //x2=30.645 //y2=0.91
cc_4189 ( N_D_c_5295_n N_RN_c_7542_n ) capacitor c=0.00111227f //x=29.67 \
 //y=1.53 //x2=30.645 //y2=1.22
cc_4190 ( N_D_c_5301_n N_RN_c_7542_n ) capacitor c=0.0124075f //x=30.2 \
 //y=1.22 //x2=30.645 //y2=1.22
cc_4191 ( N_D_c_5299_n N_RN_c_7394_n ) capacitor c=0.00103227f //x=30.2 \
 //y=0.875 //x2=31.17 //y2=0.91
cc_4192 ( N_D_c_5301_n N_RN_c_7395_n ) capacitor c=0.0010154f //x=30.2 \
 //y=1.22 //x2=31.17 //y2=1.22
cc_4193 ( N_D_c_5301_n N_RN_c_7396_n ) capacitor c=9.23422e-19 //x=30.2 \
 //y=1.22 //x2=31.17 //y2=1.45
cc_4194 ( N_D_c_5280_n N_RN_c_7397_n ) capacitor c=0.00203769f //x=29.97 \
 //y=2.08 //x2=31.17 //y2=1.915
cc_4195 ( N_D_c_5296_n N_RN_c_7397_n ) capacitor c=0.00834532f //x=29.67 \
 //y=1.915 //x2=31.17 //y2=1.915
cc_4196 ( N_D_c_5302_n N_RN_c_7549_n ) capacitor c=5.72482e-19 //x=58.53 \
 //y=0.875 //x2=59.505 //y2=0.91
cc_4197 ( N_D_c_5304_n N_RN_c_7549_n ) capacitor c=0.00149976f //x=58.53 \
 //y=1.22 //x2=59.505 //y2=0.91
cc_4198 ( N_D_c_5309_n N_RN_c_7549_n ) capacitor c=0.0160123f //x=59.06 \
 //y=0.875 //x2=59.505 //y2=0.91
cc_4199 ( N_D_c_5305_n N_RN_c_7552_n ) capacitor c=0.00111227f //x=58.53 \
 //y=1.53 //x2=59.505 //y2=1.22
cc_4200 ( N_D_c_5311_n N_RN_c_7552_n ) capacitor c=0.0124075f //x=59.06 \
 //y=1.22 //x2=59.505 //y2=1.22
cc_4201 ( N_D_c_5309_n N_RN_c_7554_n ) capacitor c=0.00103227f //x=59.06 \
 //y=0.875 //x2=60.03 //y2=0.91
cc_4202 ( N_D_c_5311_n N_RN_c_7555_n ) capacitor c=0.0010154f //x=59.06 \
 //y=1.22 //x2=60.03 //y2=1.22
cc_4203 ( N_D_c_5311_n N_RN_c_7556_n ) capacitor c=9.23422e-19 //x=59.06 \
 //y=1.22 //x2=60.03 //y2=1.45
cc_4204 ( N_D_c_5281_n N_RN_c_7557_n ) capacitor c=0.00203769f //x=58.83 \
 //y=2.08 //x2=60.03 //y2=1.915
cc_4205 ( N_D_c_5306_n N_RN_c_7557_n ) capacitor c=0.00834532f //x=58.53 \
 //y=1.915 //x2=60.03 //y2=1.915
cc_4206 ( N_D_c_5277_n N_RN_c_7162_n ) capacitor c=0.0018068f //x=29.855 \
 //y=4.07 //x2=2.22 //y2=4.7
cc_4207 ( N_D_c_5279_n N_RN_c_7162_n ) capacitor c=0.00183762f //x=1.11 \
 //y=2.08 //x2=2.22 //y2=4.7
cc_4208 ( N_D_c_5376_n N_RN_c_7162_n ) capacitor c=0.0168581f //x=1.675 \
 //y=4.79 //x2=2.22 //y2=4.7
cc_4209 ( N_D_c_5356_n N_RN_c_7162_n ) capacitor c=0.00484466f //x=1.385 \
 //y=4.79 //x2=2.22 //y2=4.7
cc_4210 ( N_D_c_5280_n N_RN_c_7261_n ) capacitor c=0.0017365f //x=29.97 \
 //y=2.08 //x2=31.08 //y2=4.7
cc_4211 ( N_D_c_5400_n N_RN_c_7261_n ) capacitor c=0.0170104f //x=30.535 \
 //y=4.79 //x2=31.08 //y2=4.7
cc_4212 ( N_D_c_5358_n N_RN_c_7261_n ) capacitor c=0.00484466f //x=30.245 \
 //y=4.79 //x2=31.08 //y2=4.7
cc_4213 ( N_D_c_5281_n N_RN_c_7264_n ) capacitor c=0.0017365f //x=58.83 \
 //y=2.08 //x2=59.94 //y2=4.7
cc_4214 ( N_D_c_5402_n N_RN_c_7264_n ) capacitor c=0.0170104f //x=59.395 \
 //y=4.79 //x2=59.94 //y2=4.7
cc_4215 ( N_D_c_5360_n N_RN_c_7264_n ) capacitor c=0.00484466f //x=59.105 \
 //y=4.79 //x2=59.94 //y2=4.7
cc_4216 ( N_D_c_5277_n N_SN_c_8129_n ) capacitor c=0.0135139f //x=29.855 \
 //y=4.07 //x2=26.155 //y2=2.96
cc_4217 ( N_D_c_5277_n N_SN_c_8132_n ) capacitor c=0.0546548f //x=29.855 \
 //y=4.07 //x2=40.585 //y2=2.96
cc_4218 ( N_D_c_5328_n N_SN_c_8132_n ) capacitor c=0.0790505f //x=58.715 \
 //y=4.07 //x2=40.585 //y2=2.96
cc_4219 ( N_D_c_5334_n N_SN_c_8132_n ) capacitor c=0.00684657f //x=30.085 \
 //y=4.07 //x2=40.585 //y2=2.96
cc_4220 ( N_D_c_5280_n N_SN_c_8132_n ) capacitor c=0.0260004f //x=29.97 \
 //y=2.08 //x2=40.585 //y2=2.96
cc_4221 ( N_D_c_5328_n N_SN_c_8135_n ) capacitor c=0.0175581f //x=58.715 \
 //y=4.07 //x2=55.015 //y2=2.96
cc_4222 ( N_D_c_5328_n N_SN_c_8138_n ) capacitor c=0.011813f //x=58.715 \
 //y=4.07 //x2=69.445 //y2=2.96
cc_4223 ( N_D_c_5281_n N_SN_c_8138_n ) capacitor c=0.0243892f //x=58.83 \
 //y=2.08 //x2=69.445 //y2=2.96
cc_4224 ( N_D_c_5277_n N_SN_c_8145_n ) capacitor c=0.0190126f //x=29.855 \
 //y=4.07 //x2=11.84 //y2=2.08
cc_4225 ( N_D_c_5277_n N_SN_c_8146_n ) capacitor c=0.0190126f //x=29.855 \
 //y=4.07 //x2=26.27 //y2=2.08
cc_4226 ( N_D_c_5328_n N_SN_c_8147_n ) capacitor c=0.0190126f //x=58.715 \
 //y=4.07 //x2=40.7 //y2=2.08
cc_4227 ( N_D_c_5328_n N_SN_c_8148_n ) capacitor c=0.0190126f //x=58.715 \
 //y=4.07 //x2=55.13 //y2=2.08
cc_4228 ( N_D_c_5328_n N_noxref_26_c_10048_n ) capacitor c=0.00990238f \
 //x=58.715 //y=4.07 //x2=53.905 //y2=3.33
cc_4229 ( N_D_c_5328_n N_noxref_26_c_10043_n ) capacitor c=7.97799e-19 \
 //x=58.715 //y=4.07 //x2=52.285 //y2=3.33
cc_4230 ( N_D_c_5328_n N_noxref_26_c_10050_n ) capacitor c=0.0408046f \
 //x=58.715 //y=4.07 //x2=56.895 //y2=3.33
cc_4231 ( N_D_c_5281_n N_noxref_26_c_10050_n ) capacitor c=0.00246861f \
 //x=58.83 //y=2.08 //x2=56.895 //y2=3.33
cc_4232 ( N_D_c_5328_n N_noxref_26_c_10052_n ) capacitor c=5.3905e-19 \
 //x=58.715 //y=4.07 //x2=54.135 //y2=3.33
cc_4233 ( N_D_c_5328_n N_noxref_26_c_9933_n ) capacitor c=0.0291659f \
 //x=58.715 //y=4.07 //x2=65.035 //y2=3.7
cc_4234 ( N_D_c_5281_n N_noxref_26_c_9933_n ) capacitor c=0.0239388f //x=58.83 \
 //y=2.08 //x2=65.035 //y2=3.7
cc_4235 ( N_D_c_5328_n N_noxref_26_c_10055_n ) capacitor c=0.164893f \
 //x=58.715 //y=4.07 //x2=57.065 //y2=3.7
cc_4236 ( N_D_c_5328_n N_noxref_26_c_9958_n ) capacitor c=0.0181982f \
 //x=58.715 //y=4.07 //x2=52.17 //y2=3.33
cc_4237 ( N_D_c_5328_n N_noxref_26_c_9916_n ) capacitor c=0.019517f //x=58.715 \
 //y=4.07 //x2=54.02 //y2=2.08
cc_4238 ( N_D_c_5286_n N_noxref_28_c_10558_n ) capacitor c=0.0034165f //x=0.81 \
 //y=1.915 //x2=0.59 //y2=1.505
cc_4239 ( N_D_c_5277_n N_noxref_28_c_10542_n ) capacitor c=0.00179505f \
 //x=29.855 //y=4.07 //x2=1.475 //y2=1.59
cc_4240 ( N_D_c_5278_n N_noxref_28_c_10542_n ) capacitor c=0.00254534f \
 //x=1.225 //y=4.07 //x2=1.475 //y2=1.59
cc_4241 ( N_D_c_5279_n N_noxref_28_c_10542_n ) capacitor c=0.0122033f //x=1.11 \
 //y=2.08 //x2=1.475 //y2=1.59
cc_4242 ( N_D_c_5285_n N_noxref_28_c_10542_n ) capacitor c=0.00703864f \
 //x=0.81 //y=1.53 //x2=1.475 //y2=1.59
cc_4243 ( N_D_c_5286_n N_noxref_28_c_10542_n ) capacitor c=0.0257397f //x=0.81 \
 //y=1.915 //x2=1.475 //y2=1.59
cc_4244 ( N_D_c_5288_n N_noxref_28_c_10542_n ) capacitor c=0.00708583f \
 //x=1.185 //y=1.375 //x2=1.475 //y2=1.59
cc_4245 ( N_D_c_5291_n N_noxref_28_c_10542_n ) capacitor c=0.00698822f \
 //x=1.34 //y=1.22 //x2=1.475 //y2=1.59
cc_4246 ( N_D_c_5277_n N_noxref_28_c_10566_n ) capacitor c=0.00316643f \
 //x=29.855 //y=4.07 //x2=2.445 //y2=1.59
cc_4247 ( N_D_c_5277_n N_noxref_28_M0_noxref_s ) capacitor c=0.00122424f \
 //x=29.855 //y=4.07 //x2=0.455 //y2=0.375
cc_4248 ( N_D_c_5282_n N_noxref_28_M0_noxref_s ) capacitor c=0.0327271f \
 //x=0.81 //y=0.875 //x2=0.455 //y2=0.375
cc_4249 ( N_D_c_5285_n N_noxref_28_M0_noxref_s ) capacitor c=7.99997e-19 \
 //x=0.81 //y=1.53 //x2=0.455 //y2=0.375
cc_4250 ( N_D_c_5286_n N_noxref_28_M0_noxref_s ) capacitor c=0.00122123f \
 //x=0.81 //y=1.915 //x2=0.455 //y2=0.375
cc_4251 ( N_D_c_5289_n N_noxref_28_M0_noxref_s ) capacitor c=0.0121427f \
 //x=1.34 //y=0.875 //x2=0.455 //y2=0.375
cc_4252 ( N_D_c_5296_n N_noxref_40_c_11167_n ) capacitor c=0.0034165f \
 //x=29.67 //y=1.915 //x2=29.45 //y2=1.505
cc_4253 ( N_D_c_5280_n N_noxref_40_c_11152_n ) capacitor c=0.0115578f \
 //x=29.97 //y=2.08 //x2=30.335 //y2=1.59
cc_4254 ( N_D_c_5295_n N_noxref_40_c_11152_n ) capacitor c=0.00697148f \
 //x=29.67 //y=1.53 //x2=30.335 //y2=1.59
cc_4255 ( N_D_c_5296_n N_noxref_40_c_11152_n ) capacitor c=0.0204849f \
 //x=29.67 //y=1.915 //x2=30.335 //y2=1.59
cc_4256 ( N_D_c_5298_n N_noxref_40_c_11152_n ) capacitor c=0.00610316f \
 //x=30.045 //y=1.375 //x2=30.335 //y2=1.59
cc_4257 ( N_D_c_5301_n N_noxref_40_c_11152_n ) capacitor c=0.00698822f \
 //x=30.2 //y=1.22 //x2=30.335 //y2=1.59
cc_4258 ( N_D_c_5292_n N_noxref_40_M18_noxref_s ) capacitor c=0.0327271f \
 //x=29.67 //y=0.875 //x2=29.315 //y2=0.375
cc_4259 ( N_D_c_5295_n N_noxref_40_M18_noxref_s ) capacitor c=7.99997e-19 \
 //x=29.67 //y=1.53 //x2=29.315 //y2=0.375
cc_4260 ( N_D_c_5296_n N_noxref_40_M18_noxref_s ) capacitor c=0.00122123f \
 //x=29.67 //y=1.915 //x2=29.315 //y2=0.375
cc_4261 ( N_D_c_5299_n N_noxref_40_M18_noxref_s ) capacitor c=0.0121427f \
 //x=30.2 //y=0.875 //x2=29.315 //y2=0.375
cc_4262 ( N_D_c_5306_n N_noxref_52_c_11780_n ) capacitor c=0.0034165f \
 //x=58.53 //y=1.915 //x2=58.31 //y2=1.505
cc_4263 ( N_D_c_5281_n N_noxref_52_c_11765_n ) capacitor c=0.0115578f \
 //x=58.83 //y=2.08 //x2=59.195 //y2=1.59
cc_4264 ( N_D_c_5305_n N_noxref_52_c_11765_n ) capacitor c=0.00697148f \
 //x=58.53 //y=1.53 //x2=59.195 //y2=1.59
cc_4265 ( N_D_c_5306_n N_noxref_52_c_11765_n ) capacitor c=0.0204849f \
 //x=58.53 //y=1.915 //x2=59.195 //y2=1.59
cc_4266 ( N_D_c_5308_n N_noxref_52_c_11765_n ) capacitor c=0.00610316f \
 //x=58.905 //y=1.375 //x2=59.195 //y2=1.59
cc_4267 ( N_D_c_5311_n N_noxref_52_c_11765_n ) capacitor c=0.00698822f \
 //x=59.06 //y=1.22 //x2=59.195 //y2=1.59
cc_4268 ( N_D_c_5302_n N_noxref_52_M36_noxref_s ) capacitor c=0.0327271f \
 //x=58.53 //y=0.875 //x2=58.175 //y2=0.375
cc_4269 ( N_D_c_5305_n N_noxref_52_M36_noxref_s ) capacitor c=7.99997e-19 \
 //x=58.53 //y=1.53 //x2=58.175 //y2=0.375
cc_4270 ( N_D_c_5306_n N_noxref_52_M36_noxref_s ) capacitor c=0.00122123f \
 //x=58.53 //y=1.915 //x2=58.175 //y2=0.375
cc_4271 ( N_D_c_5309_n N_noxref_52_M36_noxref_s ) capacitor c=0.0121427f \
 //x=59.06 //y=0.875 //x2=58.175 //y2=0.375
cc_4272 ( N_noxref_15_c_5621_n N_noxref_16_c_5873_n ) capacitor c=0.00564994f \
 //x=68.335 //y=2.59 //x2=71.525 //y2=2.59
cc_4273 ( N_noxref_15_M145_noxref_g N_noxref_16_c_5888_n ) capacitor \
 c=0.0157304f //x=69.09 //y=6.02 //x2=69.665 //y2=5.155
cc_4274 ( N_noxref_15_M144_noxref_g N_noxref_16_c_5892_n ) capacitor \
 c=0.0213876f //x=68.65 //y=6.02 //x2=68.955 //y2=5.155
cc_4275 ( N_noxref_15_c_5706_n N_noxref_16_c_5892_n ) capacitor c=0.00393496f \
 //x=69.015 //y=4.79 //x2=68.955 //y2=5.155
cc_4276 ( N_noxref_15_M145_noxref_g N_noxref_16_M144_noxref_d ) capacitor \
 c=0.0180032f //x=69.09 //y=6.02 //x2=68.725 //y2=5.02
cc_4277 ( N_noxref_15_c_5624_n N_CLK_c_6070_n ) capacitor c=0.0189507f \
 //x=61.79 //y=2.59 //x2=64.635 //y2=4.44
cc_4278 ( N_noxref_15_c_5625_n N_CLK_c_6070_n ) capacitor c=0.0211266f \
 //x=63.64 //y=2.08 //x2=64.635 //y2=4.44
cc_4279 ( N_noxref_15_c_5677_n N_CLK_c_6070_n ) capacitor c=0.0112124f \
 //x=63.915 //y=4.79 //x2=64.635 //y2=4.44
cc_4280 ( N_noxref_15_c_5626_n N_CLK_c_6074_n ) capacitor c=0.018786f \
 //x=68.45 //y=2.08 //x2=74.255 //y2=4.44
cc_4281 ( N_noxref_15_c_5679_n N_CLK_c_6074_n ) capacitor c=0.0112124f \
 //x=68.725 //y=4.79 //x2=74.255 //y2=4.44
cc_4282 ( N_noxref_15_c_5625_n N_CLK_c_6196_n ) capacitor c=0.00153281f \
 //x=63.64 //y=2.08 //x2=64.865 //y2=4.44
cc_4283 ( N_noxref_15_c_5621_n N_CLK_c_6044_n ) capacitor c=0.0190006f \
 //x=68.335 //y=2.59 //x2=64.75 //y2=2.08
cc_4284 ( N_noxref_15_c_5622_n N_CLK_c_6044_n ) capacitor c=9.95819e-19 \
 //x=63.755 //y=2.59 //x2=64.75 //y2=2.08
cc_4285 ( N_noxref_15_c_5624_n N_CLK_c_6044_n ) capacitor c=5.19237e-19 \
 //x=61.79 //y=2.59 //x2=64.75 //y2=2.08
cc_4286 ( N_noxref_15_c_5625_n N_CLK_c_6044_n ) capacitor c=0.0412985f \
 //x=63.64 //y=2.08 //x2=64.75 //y2=2.08
cc_4287 ( N_noxref_15_c_5631_n N_CLK_c_6044_n ) capacitor c=0.00210802f \
 //x=63.34 //y=1.915 //x2=64.75 //y2=2.08
cc_4288 ( N_noxref_15_c_5704_n N_CLK_c_6044_n ) capacitor c=0.00120758f \
 //x=64.205 //y=4.79 //x2=64.75 //y2=2.08
cc_4289 ( N_noxref_15_c_5677_n N_CLK_c_6044_n ) capacitor c=0.00141297f \
 //x=63.915 //y=4.79 //x2=64.75 //y2=2.08
cc_4290 ( N_noxref_15_M138_noxref_g N_CLK_M140_noxref_g ) capacitor \
 c=0.0105174f //x=63.84 //y=6.02 //x2=64.72 //y2=6.02
cc_4291 ( N_noxref_15_M139_noxref_g N_CLK_M140_noxref_g ) capacitor c=0.10624f \
 //x=64.28 //y=6.02 //x2=64.72 //y2=6.02
cc_4292 ( N_noxref_15_M139_noxref_g N_CLK_M141_noxref_g ) capacitor \
 c=0.0100903f //x=64.28 //y=6.02 //x2=65.16 //y2=6.02
cc_4293 ( N_noxref_15_c_5627_n N_CLK_c_6421_n ) capacitor c=5.72482e-19 \
 //x=63.34 //y=0.875 //x2=64.315 //y2=0.91
cc_4294 ( N_noxref_15_c_5629_n N_CLK_c_6421_n ) capacitor c=0.00149976f \
 //x=63.34 //y=1.22 //x2=64.315 //y2=0.91
cc_4295 ( N_noxref_15_c_5634_n N_CLK_c_6421_n ) capacitor c=0.0160123f \
 //x=63.87 //y=0.875 //x2=64.315 //y2=0.91
cc_4296 ( N_noxref_15_c_5630_n N_CLK_c_6424_n ) capacitor c=0.00111227f \
 //x=63.34 //y=1.53 //x2=64.315 //y2=1.22
cc_4297 ( N_noxref_15_c_5636_n N_CLK_c_6424_n ) capacitor c=0.0124075f \
 //x=63.87 //y=1.22 //x2=64.315 //y2=1.22
cc_4298 ( N_noxref_15_c_5634_n N_CLK_c_6426_n ) capacitor c=0.00103227f \
 //x=63.87 //y=0.875 //x2=64.84 //y2=0.91
cc_4299 ( N_noxref_15_c_5636_n N_CLK_c_6427_n ) capacitor c=0.0010154f \
 //x=63.87 //y=1.22 //x2=64.84 //y2=1.22
cc_4300 ( N_noxref_15_c_5636_n N_CLK_c_6428_n ) capacitor c=9.23422e-19 \
 //x=63.87 //y=1.22 //x2=64.84 //y2=1.45
cc_4301 ( N_noxref_15_c_5625_n N_CLK_c_6429_n ) capacitor c=0.00203769f \
 //x=63.64 //y=2.08 //x2=64.84 //y2=1.915
cc_4302 ( N_noxref_15_c_5631_n N_CLK_c_6429_n ) capacitor c=0.00834532f \
 //x=63.34 //y=1.915 //x2=64.84 //y2=1.915
cc_4303 ( N_noxref_15_c_5625_n N_CLK_c_6217_n ) capacitor c=0.0017365f \
 //x=63.64 //y=2.08 //x2=64.75 //y2=4.7
cc_4304 ( N_noxref_15_c_5704_n N_CLK_c_6217_n ) capacitor c=0.0170104f \
 //x=64.205 //y=4.79 //x2=64.75 //y2=4.7
cc_4305 ( N_noxref_15_c_5677_n N_CLK_c_6217_n ) capacitor c=0.00484466f \
 //x=63.915 //y=4.79 //x2=64.75 //y2=4.7
cc_4306 ( N_noxref_15_c_5619_n N_noxref_18_c_6814_n ) capacitor c=0.0111384f \
 //x=63.525 //y=2.59 //x2=66.485 //y2=3.33
cc_4307 ( N_noxref_15_c_5620_n N_noxref_18_c_6814_n ) capacitor c=8.87672e-19 \
 //x=61.905 //y=2.59 //x2=66.485 //y2=3.33
cc_4308 ( N_noxref_15_c_5621_n N_noxref_18_c_6814_n ) capacitor c=0.0246405f \
 //x=68.335 //y=2.59 //x2=66.485 //y2=3.33
cc_4309 ( N_noxref_15_c_5622_n N_noxref_18_c_6814_n ) capacitor c=5.36573e-19 \
 //x=63.755 //y=2.59 //x2=66.485 //y2=3.33
cc_4310 ( N_noxref_15_c_5624_n N_noxref_18_c_6814_n ) capacitor c=0.018769f \
 //x=61.79 //y=2.59 //x2=66.485 //y2=3.33
cc_4311 ( N_noxref_15_c_5625_n N_noxref_18_c_6814_n ) capacitor c=0.0197803f \
 //x=63.64 //y=2.08 //x2=66.485 //y2=3.33
cc_4312 ( N_noxref_15_c_5624_n N_noxref_18_c_6820_n ) capacitor c=0.00179385f \
 //x=61.79 //y=2.59 //x2=61.165 //y2=3.33
cc_4313 ( N_noxref_15_c_5621_n N_noxref_18_c_6821_n ) capacitor c=0.0118993f \
 //x=68.335 //y=2.59 //x2=77.955 //y2=3.33
cc_4314 ( N_noxref_15_c_5626_n N_noxref_18_c_6821_n ) capacitor c=0.0197803f \
 //x=68.45 //y=2.08 //x2=77.955 //y2=3.33
cc_4315 ( N_noxref_15_c_5621_n N_noxref_18_c_6823_n ) capacitor c=5.76706e-19 \
 //x=68.335 //y=2.59 //x2=66.715 //y2=3.33
cc_4316 ( N_noxref_15_c_5626_n N_noxref_18_c_6823_n ) capacitor c=7.01366e-19 \
 //x=68.45 //y=2.08 //x2=66.715 //y2=3.33
cc_4317 ( N_noxref_15_c_5620_n N_noxref_18_c_6747_n ) capacitor c=0.00687545f \
 //x=61.905 //y=2.59 //x2=61.05 //y2=2.08
cc_4318 ( N_noxref_15_c_5624_n N_noxref_18_c_6747_n ) capacitor c=0.0764456f \
 //x=61.79 //y=2.59 //x2=61.05 //y2=2.08
cc_4319 ( N_noxref_15_c_5625_n N_noxref_18_c_6747_n ) capacitor c=6.21485e-19 \
 //x=63.64 //y=2.08 //x2=61.05 //y2=2.08
cc_4320 ( N_noxref_15_c_5761_p N_noxref_18_c_6747_n ) capacitor c=0.013297f \
 //x=61.01 //y=5.155 //x2=61.05 //y2=2.08
cc_4321 ( N_noxref_15_M139_noxref_g N_noxref_18_c_6762_n ) capacitor \
 c=0.0157304f //x=64.28 //y=6.02 //x2=64.855 //y2=5.155
cc_4322 ( N_noxref_15_c_5658_n N_noxref_18_c_6766_n ) capacitor c=3.10026e-19 \
 //x=61.705 //y=5.155 //x2=64.145 //y2=5.155
cc_4323 ( N_noxref_15_M138_noxref_g N_noxref_18_c_6766_n ) capacitor \
 c=0.0213876f //x=63.84 //y=6.02 //x2=64.145 //y2=5.155
cc_4324 ( N_noxref_15_c_5704_n N_noxref_18_c_6766_n ) capacitor c=0.00393496f \
 //x=64.205 //y=4.79 //x2=64.145 //y2=5.155
cc_4325 ( N_noxref_15_c_5621_n N_noxref_18_c_6776_n ) capacitor c=0.0165903f \
 //x=68.335 //y=2.59 //x2=66.6 //y2=3.33
cc_4326 ( N_noxref_15_c_5626_n N_noxref_18_c_6776_n ) capacitor c=0.0104256f \
 //x=68.45 //y=2.08 //x2=66.6 //y2=3.33
cc_4327 ( N_noxref_15_c_5654_n N_noxref_18_M136_noxref_g ) capacitor \
 c=0.0162556f //x=60.925 //y=5.155 //x2=60.79 //y2=6.02
cc_4328 ( N_noxref_15_M136_noxref_d N_noxref_18_M136_noxref_g ) capacitor \
 c=0.0180032f //x=60.865 //y=5.02 //x2=60.79 //y2=6.02
cc_4329 ( N_noxref_15_c_5658_n N_noxref_18_M137_noxref_g ) capacitor \
 c=0.0183937f //x=61.705 //y=5.155 //x2=61.23 //y2=6.02
cc_4330 ( N_noxref_15_M136_noxref_d N_noxref_18_M137_noxref_g ) capacitor \
 c=0.0194246f //x=60.865 //y=5.02 //x2=61.23 //y2=6.02
cc_4331 ( N_noxref_15_M38_noxref_d N_noxref_18_c_6839_n ) capacitor \
 c=0.00217566f //x=61.115 //y=0.915 //x2=61.04 //y2=0.915
cc_4332 ( N_noxref_15_M38_noxref_d N_noxref_18_c_6840_n ) capacitor \
 c=0.0034598f //x=61.115 //y=0.915 //x2=61.04 //y2=1.26
cc_4333 ( N_noxref_15_M38_noxref_d N_noxref_18_c_6841_n ) capacitor \
 c=0.00546784f //x=61.115 //y=0.915 //x2=61.04 //y2=1.57
cc_4334 ( N_noxref_15_M38_noxref_d N_noxref_18_c_6842_n ) capacitor \
 c=0.00241102f //x=61.115 //y=0.915 //x2=61.415 //y2=0.76
cc_4335 ( N_noxref_15_c_5623_n N_noxref_18_c_6843_n ) capacitor c=0.00371277f \
 //x=61.705 //y=1.665 //x2=61.415 //y2=1.415
cc_4336 ( N_noxref_15_M38_noxref_d N_noxref_18_c_6843_n ) capacitor \
 c=0.0138621f //x=61.115 //y=0.915 //x2=61.415 //y2=1.415
cc_4337 ( N_noxref_15_M38_noxref_d N_noxref_18_c_6845_n ) capacitor \
 c=0.00219619f //x=61.115 //y=0.915 //x2=61.57 //y2=0.915
cc_4338 ( N_noxref_15_c_5623_n N_noxref_18_c_6846_n ) capacitor c=0.00457401f \
 //x=61.705 //y=1.665 //x2=61.57 //y2=1.26
cc_4339 ( N_noxref_15_M38_noxref_d N_noxref_18_c_6846_n ) capacitor \
 c=0.00603828f //x=61.115 //y=0.915 //x2=61.57 //y2=1.26
cc_4340 ( N_noxref_15_c_5624_n N_noxref_18_c_6848_n ) capacitor c=0.00709342f \
 //x=61.79 //y=2.59 //x2=61.05 //y2=2.08
cc_4341 ( N_noxref_15_c_5624_n N_noxref_18_c_6849_n ) capacitor c=0.00283672f \
 //x=61.79 //y=2.59 //x2=61.05 //y2=1.915
cc_4342 ( N_noxref_15_M38_noxref_d N_noxref_18_c_6849_n ) capacitor \
 c=0.00661782f //x=61.115 //y=0.915 //x2=61.05 //y2=1.915
cc_4343 ( N_noxref_15_c_5658_n N_noxref_18_c_6812_n ) capacitor c=0.00201851f \
 //x=61.705 //y=5.155 //x2=61.05 //y2=4.7
cc_4344 ( N_noxref_15_c_5624_n N_noxref_18_c_6812_n ) capacitor c=0.0114782f \
 //x=61.79 //y=2.59 //x2=61.05 //y2=4.7
cc_4345 ( N_noxref_15_c_5761_p N_noxref_18_c_6812_n ) capacitor c=0.00470675f \
 //x=61.01 //y=5.155 //x2=61.05 //y2=4.7
cc_4346 ( N_noxref_15_M139_noxref_g N_noxref_18_M138_noxref_d ) capacitor \
 c=0.0180032f //x=64.28 //y=6.02 //x2=63.915 //y2=5.02
cc_4347 ( N_noxref_15_c_5619_n N_RN_c_7071_n ) capacitor c=0.143487f \
 //x=63.525 //y=2.59 //x2=75.365 //y2=2.22
cc_4348 ( N_noxref_15_c_5620_n N_RN_c_7071_n ) capacitor c=0.0291301f \
 //x=61.905 //y=2.59 //x2=75.365 //y2=2.22
cc_4349 ( N_noxref_15_c_5621_n N_RN_c_7071_n ) capacitor c=0.42762f //x=68.335 \
 //y=2.59 //x2=75.365 //y2=2.22
cc_4350 ( N_noxref_15_c_5622_n N_RN_c_7071_n ) capacitor c=0.0264401f \
 //x=63.755 //y=2.59 //x2=75.365 //y2=2.22
cc_4351 ( N_noxref_15_c_5792_p N_RN_c_7071_n ) capacitor c=0.016327f //x=61.39 \
 //y=1.665 //x2=75.365 //y2=2.22
cc_4352 ( N_noxref_15_c_5624_n N_RN_c_7071_n ) capacitor c=0.0215653f \
 //x=61.79 //y=2.59 //x2=75.365 //y2=2.22
cc_4353 ( N_noxref_15_c_5625_n N_RN_c_7071_n ) capacitor c=0.021104f //x=63.64 \
 //y=2.08 //x2=75.365 //y2=2.22
cc_4354 ( N_noxref_15_c_5626_n N_RN_c_7071_n ) capacitor c=0.021104f //x=68.45 \
 //y=2.08 //x2=75.365 //y2=2.22
cc_4355 ( N_noxref_15_c_5631_n N_RN_c_7071_n ) capacitor c=0.011987f //x=63.34 \
 //y=1.915 //x2=75.365 //y2=2.22
cc_4356 ( N_noxref_15_c_5641_n N_RN_c_7071_n ) capacitor c=0.011987f //x=68.15 \
 //y=1.915 //x2=75.365 //y2=2.22
cc_4357 ( N_noxref_15_c_5648_n N_RN_c_7094_n ) capacitor c=0.0120276f \
 //x=60.045 //y=5.155 //x2=59.94 //y2=2.08
cc_4358 ( N_noxref_15_c_5624_n N_RN_c_7094_n ) capacitor c=0.00275195f \
 //x=61.79 //y=2.59 //x2=59.94 //y2=2.08
cc_4359 ( N_noxref_15_c_5648_n N_RN_M134_noxref_g ) capacitor c=0.0163793f \
 //x=60.045 //y=5.155 //x2=59.91 //y2=6.02
cc_4360 ( N_noxref_15_M134_noxref_d N_RN_M134_noxref_g ) capacitor \
 c=0.0180032f //x=59.985 //y=5.02 //x2=59.91 //y2=6.02
cc_4361 ( N_noxref_15_c_5654_n N_RN_M135_noxref_g ) capacitor c=0.0162556f \
 //x=60.925 //y=5.155 //x2=60.35 //y2=6.02
cc_4362 ( N_noxref_15_M134_noxref_d N_RN_M135_noxref_g ) capacitor \
 c=0.0180032f //x=59.985 //y=5.02 //x2=60.35 //y2=6.02
cc_4363 ( N_noxref_15_c_5804_p N_RN_c_7258_n ) capacitor c=0.00392095f \
 //x=60.13 //y=5.155 //x2=60.275 //y2=4.79
cc_4364 ( N_noxref_15_c_5648_n N_RN_c_7264_n ) capacitor c=0.00309994f \
 //x=60.045 //y=5.155 //x2=59.94 //y2=4.7
cc_4365 ( N_noxref_15_c_5619_n N_SN_c_8138_n ) capacitor c=0.143324f \
 //x=63.525 //y=2.59 //x2=69.445 //y2=2.96
cc_4366 ( N_noxref_15_c_5620_n N_SN_c_8138_n ) capacitor c=0.0293832f \
 //x=61.905 //y=2.59 //x2=69.445 //y2=2.96
cc_4367 ( N_noxref_15_c_5621_n N_SN_c_8138_n ) capacitor c=0.429547f \
 //x=68.335 //y=2.59 //x2=69.445 //y2=2.96
cc_4368 ( N_noxref_15_c_5622_n N_SN_c_8138_n ) capacitor c=0.0267736f \
 //x=63.755 //y=2.59 //x2=69.445 //y2=2.96
cc_4369 ( N_noxref_15_c_5624_n N_SN_c_8138_n ) capacitor c=0.0206007f \
 //x=61.79 //y=2.59 //x2=69.445 //y2=2.96
cc_4370 ( N_noxref_15_c_5625_n N_SN_c_8138_n ) capacitor c=0.0216195f \
 //x=63.64 //y=2.08 //x2=69.445 //y2=2.96
cc_4371 ( N_noxref_15_c_5626_n N_SN_c_8138_n ) capacitor c=0.0215933f \
 //x=68.45 //y=2.08 //x2=69.445 //y2=2.96
cc_4372 ( N_noxref_15_c_5626_n N_SN_c_8468_n ) capacitor c=0.00128547f \
 //x=68.45 //y=2.08 //x2=69.675 //y2=2.96
cc_4373 ( N_noxref_15_c_5621_n N_SN_c_8149_n ) capacitor c=0.00311593f \
 //x=68.335 //y=2.59 //x2=69.56 //y2=2.08
cc_4374 ( N_noxref_15_c_5626_n N_SN_c_8149_n ) capacitor c=0.0408822f \
 //x=68.45 //y=2.08 //x2=69.56 //y2=2.08
cc_4375 ( N_noxref_15_c_5641_n N_SN_c_8149_n ) capacitor c=0.00210802f \
 //x=68.15 //y=1.915 //x2=69.56 //y2=2.08
cc_4376 ( N_noxref_15_c_5706_n N_SN_c_8149_n ) capacitor c=0.00120758f \
 //x=69.015 //y=4.79 //x2=69.56 //y2=2.08
cc_4377 ( N_noxref_15_c_5679_n N_SN_c_8149_n ) capacitor c=0.00142741f \
 //x=68.725 //y=4.79 //x2=69.56 //y2=2.08
cc_4378 ( N_noxref_15_M144_noxref_g N_SN_M146_noxref_g ) capacitor \
 c=0.0105174f //x=68.65 //y=6.02 //x2=69.53 //y2=6.02
cc_4379 ( N_noxref_15_M145_noxref_g N_SN_M146_noxref_g ) capacitor c=0.10624f \
 //x=69.09 //y=6.02 //x2=69.53 //y2=6.02
cc_4380 ( N_noxref_15_M145_noxref_g N_SN_M147_noxref_g ) capacitor \
 c=0.0100903f //x=69.09 //y=6.02 //x2=69.97 //y2=6.02
cc_4381 ( N_noxref_15_c_5637_n N_SN_c_8477_n ) capacitor c=5.72482e-19 \
 //x=68.15 //y=0.875 //x2=69.125 //y2=0.91
cc_4382 ( N_noxref_15_c_5639_n N_SN_c_8477_n ) capacitor c=0.00149976f \
 //x=68.15 //y=1.22 //x2=69.125 //y2=0.91
cc_4383 ( N_noxref_15_c_5644_n N_SN_c_8477_n ) capacitor c=0.0160123f \
 //x=68.68 //y=0.875 //x2=69.125 //y2=0.91
cc_4384 ( N_noxref_15_c_5640_n N_SN_c_8480_n ) capacitor c=0.00111227f \
 //x=68.15 //y=1.53 //x2=69.125 //y2=1.22
cc_4385 ( N_noxref_15_c_5646_n N_SN_c_8480_n ) capacitor c=0.0124075f \
 //x=68.68 //y=1.22 //x2=69.125 //y2=1.22
cc_4386 ( N_noxref_15_c_5644_n N_SN_c_8482_n ) capacitor c=0.00103227f \
 //x=68.68 //y=0.875 //x2=69.65 //y2=0.91
cc_4387 ( N_noxref_15_c_5646_n N_SN_c_8483_n ) capacitor c=0.0010154f \
 //x=68.68 //y=1.22 //x2=69.65 //y2=1.22
cc_4388 ( N_noxref_15_c_5646_n N_SN_c_8484_n ) capacitor c=9.23422e-19 \
 //x=68.68 //y=1.22 //x2=69.65 //y2=1.45
cc_4389 ( N_noxref_15_c_5626_n N_SN_c_8485_n ) capacitor c=0.00203769f \
 //x=68.45 //y=2.08 //x2=69.65 //y2=1.915
cc_4390 ( N_noxref_15_c_5641_n N_SN_c_8485_n ) capacitor c=0.00834532f \
 //x=68.15 //y=1.915 //x2=69.65 //y2=1.915
cc_4391 ( N_noxref_15_c_5626_n N_SN_c_8270_n ) capacitor c=0.0017365f \
 //x=68.45 //y=2.08 //x2=69.56 //y2=4.7
cc_4392 ( N_noxref_15_c_5706_n N_SN_c_8270_n ) capacitor c=0.0170104f \
 //x=69.015 //y=4.79 //x2=69.56 //y2=4.7
cc_4393 ( N_noxref_15_c_5679_n N_SN_c_8270_n ) capacitor c=0.00484466f \
 //x=68.725 //y=4.79 //x2=69.56 //y2=4.7
cc_4394 ( N_noxref_15_c_5626_n N_noxref_21_c_8898_n ) capacitor c=0.0197627f \
 //x=68.45 //y=2.08 //x2=70.555 //y2=3.7
cc_4395 ( N_noxref_15_c_5621_n N_noxref_21_c_8828_n ) capacitor c=0.0179628f \
 //x=68.335 //y=2.59 //x2=65.86 //y2=2.08
cc_4396 ( N_noxref_15_c_5625_n N_noxref_21_c_8828_n ) capacitor c=0.00133811f \
 //x=63.64 //y=2.08 //x2=65.86 //y2=2.08
cc_4397 ( N_noxref_15_c_5626_n N_noxref_21_c_8828_n ) capacitor c=7.12947e-19 \
 //x=68.45 //y=2.08 //x2=65.86 //y2=2.08
cc_4398 ( N_noxref_15_c_5626_n N_noxref_21_c_8829_n ) capacitor c=0.00106679f \
 //x=68.45 //y=2.08 //x2=70.67 //y2=2.08
cc_4399 ( N_noxref_15_c_5624_n N_noxref_26_c_9933_n ) capacitor c=0.0211104f \
 //x=61.79 //y=2.59 //x2=65.035 //y2=3.7
cc_4400 ( N_noxref_15_c_5625_n N_noxref_26_c_9933_n ) capacitor c=0.022094f \
 //x=63.64 //y=2.08 //x2=65.035 //y2=3.7
cc_4401 ( N_noxref_15_c_5626_n N_noxref_26_c_9912_n ) capacitor c=0.0194977f \
 //x=68.45 //y=2.08 //x2=88.315 //y2=4.07
cc_4402 ( N_noxref_15_M38_noxref_d N_noxref_52_M36_noxref_s ) capacitor \
 c=0.00309936f //x=61.115 //y=0.915 //x2=58.175 //y2=0.375
cc_4403 ( N_noxref_15_c_5623_n N_noxref_53_c_11822_n ) capacitor c=0.00457167f \
 //x=61.705 //y=1.665 //x2=61.705 //y2=0.54
cc_4404 ( N_noxref_15_M38_noxref_d N_noxref_53_c_11822_n ) capacitor \
 c=0.0115903f //x=61.115 //y=0.915 //x2=61.705 //y2=0.54
cc_4405 ( N_noxref_15_c_5792_p N_noxref_53_c_11832_n ) capacitor c=0.0200405f \
 //x=61.39 //y=1.665 //x2=60.82 //y2=0.995
cc_4406 ( N_noxref_15_M38_noxref_d N_noxref_53_M37_noxref_d ) capacitor \
 c=5.27807e-19 //x=61.115 //y=0.915 //x2=59.58 //y2=0.91
cc_4407 ( N_noxref_15_c_5623_n N_noxref_53_M38_noxref_s ) capacitor \
 c=0.0184051f //x=61.705 //y=1.665 //x2=60.685 //y2=0.375
cc_4408 ( N_noxref_15_M38_noxref_d N_noxref_53_M38_noxref_s ) capacitor \
 c=0.0426368f //x=61.115 //y=0.915 //x2=60.685 //y2=0.375
cc_4409 ( N_noxref_15_c_5623_n N_noxref_54_c_11884_n ) capacitor c=3.84569e-19 \
 //x=61.705 //y=1.665 //x2=63.12 //y2=1.505
cc_4410 ( N_noxref_15_c_5631_n N_noxref_54_c_11884_n ) capacitor c=0.0034165f \
 //x=63.34 //y=1.915 //x2=63.12 //y2=1.505
cc_4411 ( N_noxref_15_c_5625_n N_noxref_54_c_11869_n ) capacitor c=0.0115578f \
 //x=63.64 //y=2.08 //x2=64.005 //y2=1.59
cc_4412 ( N_noxref_15_c_5630_n N_noxref_54_c_11869_n ) capacitor c=0.00697148f \
 //x=63.34 //y=1.53 //x2=64.005 //y2=1.59
cc_4413 ( N_noxref_15_c_5631_n N_noxref_54_c_11869_n ) capacitor c=0.0204849f \
 //x=63.34 //y=1.915 //x2=64.005 //y2=1.59
cc_4414 ( N_noxref_15_c_5633_n N_noxref_54_c_11869_n ) capacitor c=0.00610316f \
 //x=63.715 //y=1.375 //x2=64.005 //y2=1.59
cc_4415 ( N_noxref_15_c_5636_n N_noxref_54_c_11869_n ) capacitor c=0.00698822f \
 //x=63.87 //y=1.22 //x2=64.005 //y2=1.59
cc_4416 ( N_noxref_15_c_5627_n N_noxref_54_M39_noxref_s ) capacitor \
 c=0.0327271f //x=63.34 //y=0.875 //x2=62.985 //y2=0.375
cc_4417 ( N_noxref_15_c_5630_n N_noxref_54_M39_noxref_s ) capacitor \
 c=7.99997e-19 //x=63.34 //y=1.53 //x2=62.985 //y2=0.375
cc_4418 ( N_noxref_15_c_5631_n N_noxref_54_M39_noxref_s ) capacitor \
 c=0.00122123f //x=63.34 //y=1.915 //x2=62.985 //y2=0.375
cc_4419 ( N_noxref_15_c_5634_n N_noxref_54_M39_noxref_s ) capacitor \
 c=0.0121427f //x=63.87 //y=0.875 //x2=62.985 //y2=0.375
cc_4420 ( N_noxref_15_M38_noxref_d N_noxref_54_M39_noxref_s ) capacitor \
 c=2.55333e-19 //x=61.115 //y=0.915 //x2=62.985 //y2=0.375
cc_4421 ( N_noxref_15_c_5641_n N_noxref_56_c_11985_n ) capacitor c=0.0034165f \
 //x=68.15 //y=1.915 //x2=67.93 //y2=1.505
cc_4422 ( N_noxref_15_c_5626_n N_noxref_56_c_11970_n ) capacitor c=0.0115578f \
 //x=68.45 //y=2.08 //x2=68.815 //y2=1.59
cc_4423 ( N_noxref_15_c_5640_n N_noxref_56_c_11970_n ) capacitor c=0.00697148f \
 //x=68.15 //y=1.53 //x2=68.815 //y2=1.59
cc_4424 ( N_noxref_15_c_5641_n N_noxref_56_c_11970_n ) capacitor c=0.0204849f \
 //x=68.15 //y=1.915 //x2=68.815 //y2=1.59
cc_4425 ( N_noxref_15_c_5643_n N_noxref_56_c_11970_n ) capacitor c=0.00610316f \
 //x=68.525 //y=1.375 //x2=68.815 //y2=1.59
cc_4426 ( N_noxref_15_c_5646_n N_noxref_56_c_11970_n ) capacitor c=0.00698822f \
 //x=68.68 //y=1.22 //x2=68.815 //y2=1.59
cc_4427 ( N_noxref_15_c_5637_n N_noxref_56_M42_noxref_s ) capacitor \
 c=0.0327271f //x=68.15 //y=0.875 //x2=67.795 //y2=0.375
cc_4428 ( N_noxref_15_c_5640_n N_noxref_56_M42_noxref_s ) capacitor \
 c=7.99997e-19 //x=68.15 //y=1.53 //x2=67.795 //y2=0.375
cc_4429 ( N_noxref_15_c_5641_n N_noxref_56_M42_noxref_s ) capacitor \
 c=0.00122123f //x=68.15 //y=1.915 //x2=67.795 //y2=0.375
cc_4430 ( N_noxref_15_c_5644_n N_noxref_56_M42_noxref_s ) capacitor \
 c=0.0121427f //x=68.68 //y=0.875 //x2=67.795 //y2=0.375
cc_4431 ( N_noxref_16_c_5875_n N_CLK_c_6074_n ) capacitor c=0.0166101f \
 //x=71.41 //y=2.59 //x2=74.255 //y2=4.44
cc_4432 ( N_noxref_16_c_5876_n N_CLK_c_6074_n ) capacitor c=0.0202706f \
 //x=73.26 //y=2.08 //x2=74.255 //y2=4.44
cc_4433 ( N_noxref_16_c_5910_n N_CLK_c_6074_n ) capacitor c=0.0113679f \
 //x=73.535 //y=4.79 //x2=74.255 //y2=4.44
cc_4434 ( N_noxref_16_c_5872_n N_CLK_c_6045_n ) capacitor c=0.00520283f \
 //x=73.145 //y=2.59 //x2=74.37 //y2=2.08
cc_4435 ( N_noxref_16_c_5875_n N_CLK_c_6045_n ) capacitor c=2.96936e-19 \
 //x=71.41 //y=2.59 //x2=74.37 //y2=2.08
cc_4436 ( N_noxref_16_c_5876_n N_CLK_c_6045_n ) capacitor c=0.0401239f \
 //x=73.26 //y=2.08 //x2=74.37 //y2=2.08
cc_4437 ( N_noxref_16_c_5881_n N_CLK_c_6045_n ) capacitor c=0.00210802f \
 //x=72.96 //y=1.915 //x2=74.37 //y2=2.08
cc_4438 ( N_noxref_16_c_5932_n N_CLK_c_6045_n ) capacitor c=0.00120758f \
 //x=73.825 //y=4.79 //x2=74.37 //y2=2.08
cc_4439 ( N_noxref_16_c_5910_n N_CLK_c_6045_n ) capacitor c=0.00141297f \
 //x=73.535 //y=4.79 //x2=74.37 //y2=2.08
cc_4440 ( N_noxref_16_M150_noxref_g N_CLK_M152_noxref_g ) capacitor \
 c=0.0105174f //x=73.46 //y=6.02 //x2=74.34 //y2=6.02
cc_4441 ( N_noxref_16_M151_noxref_g N_CLK_M152_noxref_g ) capacitor c=0.10624f \
 //x=73.9 //y=6.02 //x2=74.34 //y2=6.02
cc_4442 ( N_noxref_16_M151_noxref_g N_CLK_M153_noxref_g ) capacitor \
 c=0.0100903f //x=73.9 //y=6.02 //x2=74.78 //y2=6.02
cc_4443 ( N_noxref_16_c_5877_n N_CLK_c_6446_n ) capacitor c=5.72482e-19 \
 //x=72.96 //y=0.875 //x2=73.935 //y2=0.91
cc_4444 ( N_noxref_16_c_5879_n N_CLK_c_6446_n ) capacitor c=0.00149976f \
 //x=72.96 //y=1.22 //x2=73.935 //y2=0.91
cc_4445 ( N_noxref_16_c_5884_n N_CLK_c_6446_n ) capacitor c=0.0160123f \
 //x=73.49 //y=0.875 //x2=73.935 //y2=0.91
cc_4446 ( N_noxref_16_c_5880_n N_CLK_c_6449_n ) capacitor c=0.00111227f \
 //x=72.96 //y=1.53 //x2=73.935 //y2=1.22
cc_4447 ( N_noxref_16_c_5886_n N_CLK_c_6449_n ) capacitor c=0.0124075f \
 //x=73.49 //y=1.22 //x2=73.935 //y2=1.22
cc_4448 ( N_noxref_16_c_5884_n N_CLK_c_6451_n ) capacitor c=0.00103227f \
 //x=73.49 //y=0.875 //x2=74.46 //y2=0.91
cc_4449 ( N_noxref_16_c_5886_n N_CLK_c_6452_n ) capacitor c=0.0010154f \
 //x=73.49 //y=1.22 //x2=74.46 //y2=1.22
cc_4450 ( N_noxref_16_c_5886_n N_CLK_c_6453_n ) capacitor c=9.23422e-19 \
 //x=73.49 //y=1.22 //x2=74.46 //y2=1.45
cc_4451 ( N_noxref_16_c_5876_n N_CLK_c_6454_n ) capacitor c=0.00203769f \
 //x=73.26 //y=2.08 //x2=74.46 //y2=1.915
cc_4452 ( N_noxref_16_c_5881_n N_CLK_c_6454_n ) capacitor c=0.00834532f \
 //x=72.96 //y=1.915 //x2=74.46 //y2=1.915
cc_4453 ( N_noxref_16_c_5876_n N_CLK_c_6218_n ) capacitor c=0.0017365f \
 //x=73.26 //y=2.08 //x2=74.37 //y2=4.7
cc_4454 ( N_noxref_16_c_5932_n N_CLK_c_6218_n ) capacitor c=0.0170104f \
 //x=73.825 //y=4.79 //x2=74.37 //y2=4.7
cc_4455 ( N_noxref_16_c_5910_n N_CLK_c_6218_n ) capacitor c=0.00484466f \
 //x=73.535 //y=4.79 //x2=74.37 //y2=4.7
cc_4456 ( N_noxref_16_c_5872_n N_noxref_18_c_6821_n ) capacitor c=0.0119023f \
 //x=73.145 //y=2.59 //x2=77.955 //y2=3.33
cc_4457 ( N_noxref_16_c_5873_n N_noxref_18_c_6821_n ) capacitor c=8.87672e-19 \
 //x=71.525 //y=2.59 //x2=77.955 //y2=3.33
cc_4458 ( N_noxref_16_c_5875_n N_noxref_18_c_6821_n ) capacitor c=0.018769f \
 //x=71.41 //y=2.59 //x2=77.955 //y2=3.33
cc_4459 ( N_noxref_16_c_5876_n N_noxref_18_c_6821_n ) capacitor c=0.0198064f \
 //x=73.26 //y=2.08 //x2=77.955 //y2=3.33
cc_4460 ( N_noxref_16_c_5892_n N_noxref_18_c_6772_n ) capacitor c=3.10026e-19 \
 //x=68.955 //y=5.155 //x2=66.515 //y2=5.155
cc_4461 ( N_noxref_16_c_5872_n N_RN_c_7071_n ) capacitor c=0.172592f \
 //x=73.145 //y=2.59 //x2=75.365 //y2=2.22
cc_4462 ( N_noxref_16_c_5873_n N_RN_c_7071_n ) capacitor c=0.0291301f \
 //x=71.525 //y=2.59 //x2=75.365 //y2=2.22
cc_4463 ( N_noxref_16_c_5971_p N_RN_c_7071_n ) capacitor c=0.016327f //x=71.01 \
 //y=1.665 //x2=75.365 //y2=2.22
cc_4464 ( N_noxref_16_c_5875_n N_RN_c_7071_n ) capacitor c=0.0215653f \
 //x=71.41 //y=2.59 //x2=75.365 //y2=2.22
cc_4465 ( N_noxref_16_c_5876_n N_RN_c_7071_n ) capacitor c=0.021104f //x=73.26 \
 //y=2.08 //x2=75.365 //y2=2.22
cc_4466 ( N_noxref_16_c_5881_n N_RN_c_7071_n ) capacitor c=0.011987f //x=72.96 \
 //y=1.915 //x2=75.365 //y2=2.22
cc_4467 ( N_noxref_16_c_5876_n N_RN_c_7095_n ) capacitor c=0.00107042f \
 //x=73.26 //y=2.08 //x2=75.48 //y2=2.08
cc_4468 ( N_noxref_16_c_5872_n N_SN_c_8141_n ) capacitor c=0.172781f \
 //x=73.145 //y=2.59 //x2=83.875 //y2=2.96
cc_4469 ( N_noxref_16_c_5873_n N_SN_c_8141_n ) capacitor c=0.0293832f \
 //x=71.525 //y=2.59 //x2=83.875 //y2=2.96
cc_4470 ( N_noxref_16_c_5875_n N_SN_c_8141_n ) capacitor c=0.0206007f \
 //x=71.41 //y=2.59 //x2=83.875 //y2=2.96
cc_4471 ( N_noxref_16_c_5876_n N_SN_c_8141_n ) capacitor c=0.0216195f \
 //x=73.26 //y=2.08 //x2=83.875 //y2=2.96
cc_4472 ( N_noxref_16_c_5888_n N_SN_c_8149_n ) capacitor c=0.0121898f \
 //x=69.665 //y=5.155 //x2=69.56 //y2=2.08
cc_4473 ( N_noxref_16_c_5875_n N_SN_c_8149_n ) capacitor c=0.00216737f \
 //x=71.41 //y=2.59 //x2=69.56 //y2=2.08
cc_4474 ( N_noxref_16_c_5888_n N_SN_M146_noxref_g ) capacitor c=0.0163793f \
 //x=69.665 //y=5.155 //x2=69.53 //y2=6.02
cc_4475 ( N_noxref_16_M146_noxref_d N_SN_M146_noxref_g ) capacitor \
 c=0.0180032f //x=69.605 //y=5.02 //x2=69.53 //y2=6.02
cc_4476 ( N_noxref_16_c_5894_n N_SN_M147_noxref_g ) capacitor c=0.0162556f \
 //x=70.545 //y=5.155 //x2=69.97 //y2=6.02
cc_4477 ( N_noxref_16_M146_noxref_d N_SN_M147_noxref_g ) capacitor \
 c=0.0180032f //x=69.605 //y=5.02 //x2=69.97 //y2=6.02
cc_4478 ( N_noxref_16_c_5986_p N_SN_c_8262_n ) capacitor c=0.00392095f \
 //x=69.75 //y=5.155 //x2=69.895 //y2=4.79
cc_4479 ( N_noxref_16_c_5888_n N_SN_c_8270_n ) capacitor c=0.00309994f \
 //x=69.665 //y=5.155 //x2=69.56 //y2=4.7
cc_4480 ( N_noxref_16_c_5875_n N_noxref_21_c_8878_n ) capacitor c=0.0187698f \
 //x=71.41 //y=2.59 //x2=76.105 //y2=3.7
cc_4481 ( N_noxref_16_c_5876_n N_noxref_21_c_8878_n ) capacitor c=0.0197889f \
 //x=73.26 //y=2.08 //x2=76.105 //y2=3.7
cc_4482 ( N_noxref_16_c_5875_n N_noxref_21_c_8905_n ) capacitor c=0.00179385f \
 //x=71.41 //y=2.59 //x2=70.785 //y2=3.7
cc_4483 ( N_noxref_16_c_5873_n N_noxref_21_c_8829_n ) capacitor c=0.00456439f \
 //x=71.525 //y=2.59 //x2=70.67 //y2=2.08
cc_4484 ( N_noxref_16_c_5875_n N_noxref_21_c_8829_n ) capacitor c=0.0750956f \
 //x=71.41 //y=2.59 //x2=70.67 //y2=2.08
cc_4485 ( N_noxref_16_c_5876_n N_noxref_21_c_8829_n ) capacitor c=5.32619e-19 \
 //x=73.26 //y=2.08 //x2=70.67 //y2=2.08
cc_4486 ( N_noxref_16_c_5994_p N_noxref_21_c_8829_n ) capacitor c=0.0126839f \
 //x=70.63 //y=5.155 //x2=70.67 //y2=2.08
cc_4487 ( N_noxref_16_M151_noxref_g N_noxref_21_c_8835_n ) capacitor \
 c=0.0157304f //x=73.9 //y=6.02 //x2=74.475 //y2=5.155
cc_4488 ( N_noxref_16_c_5898_n N_noxref_21_c_8839_n ) capacitor c=3.10026e-19 \
 //x=71.325 //y=5.155 //x2=73.765 //y2=5.155
cc_4489 ( N_noxref_16_M150_noxref_g N_noxref_21_c_8839_n ) capacitor \
 c=0.0213876f //x=73.46 //y=6.02 //x2=73.765 //y2=5.155
cc_4490 ( N_noxref_16_c_5932_n N_noxref_21_c_8839_n ) capacitor c=0.00393496f \
 //x=73.825 //y=4.79 //x2=73.765 //y2=5.155
cc_4491 ( N_noxref_16_c_5894_n N_noxref_21_M148_noxref_g ) capacitor \
 c=0.0162556f //x=70.545 //y=5.155 //x2=70.41 //y2=6.02
cc_4492 ( N_noxref_16_M148_noxref_d N_noxref_21_M148_noxref_g ) capacitor \
 c=0.0180032f //x=70.485 //y=5.02 //x2=70.41 //y2=6.02
cc_4493 ( N_noxref_16_c_5898_n N_noxref_21_M149_noxref_g ) capacitor \
 c=0.0183937f //x=71.325 //y=5.155 //x2=70.85 //y2=6.02
cc_4494 ( N_noxref_16_M148_noxref_d N_noxref_21_M149_noxref_g ) capacitor \
 c=0.0194246f //x=70.485 //y=5.02 //x2=70.85 //y2=6.02
cc_4495 ( N_noxref_16_M44_noxref_d N_noxref_21_c_8918_n ) capacitor \
 c=0.00217566f //x=70.735 //y=0.915 //x2=70.66 //y2=0.915
cc_4496 ( N_noxref_16_M44_noxref_d N_noxref_21_c_8919_n ) capacitor \
 c=0.0034598f //x=70.735 //y=0.915 //x2=70.66 //y2=1.26
cc_4497 ( N_noxref_16_M44_noxref_d N_noxref_21_c_8920_n ) capacitor \
 c=0.00546784f //x=70.735 //y=0.915 //x2=70.66 //y2=1.57
cc_4498 ( N_noxref_16_M44_noxref_d N_noxref_21_c_8921_n ) capacitor \
 c=0.00241102f //x=70.735 //y=0.915 //x2=71.035 //y2=0.76
cc_4499 ( N_noxref_16_c_5874_n N_noxref_21_c_8922_n ) capacitor c=0.00371277f \
 //x=71.325 //y=1.665 //x2=71.035 //y2=1.415
cc_4500 ( N_noxref_16_M44_noxref_d N_noxref_21_c_8922_n ) capacitor \
 c=0.0138621f //x=70.735 //y=0.915 //x2=71.035 //y2=1.415
cc_4501 ( N_noxref_16_M44_noxref_d N_noxref_21_c_8924_n ) capacitor \
 c=0.00219619f //x=70.735 //y=0.915 //x2=71.19 //y2=0.915
cc_4502 ( N_noxref_16_c_5874_n N_noxref_21_c_8925_n ) capacitor c=0.00457401f \
 //x=71.325 //y=1.665 //x2=71.19 //y2=1.26
cc_4503 ( N_noxref_16_M44_noxref_d N_noxref_21_c_8925_n ) capacitor \
 c=0.00603828f //x=70.735 //y=0.915 //x2=71.19 //y2=1.26
cc_4504 ( N_noxref_16_c_5875_n N_noxref_21_c_8927_n ) capacitor c=0.00731987f \
 //x=71.41 //y=2.59 //x2=70.67 //y2=2.08
cc_4505 ( N_noxref_16_c_5875_n N_noxref_21_c_8928_n ) capacitor c=0.00283672f \
 //x=71.41 //y=2.59 //x2=70.67 //y2=1.915
cc_4506 ( N_noxref_16_M44_noxref_d N_noxref_21_c_8928_n ) capacitor \
 c=0.00661782f //x=70.735 //y=0.915 //x2=70.67 //y2=1.915
cc_4507 ( N_noxref_16_c_5898_n N_noxref_21_c_8896_n ) capacitor c=0.00201851f \
 //x=71.325 //y=5.155 //x2=70.67 //y2=4.7
cc_4508 ( N_noxref_16_c_5875_n N_noxref_21_c_8896_n ) capacitor c=0.0114782f \
 //x=71.41 //y=2.59 //x2=70.67 //y2=4.7
cc_4509 ( N_noxref_16_c_5994_p N_noxref_21_c_8896_n ) capacitor c=0.00470675f \
 //x=70.63 //y=5.155 //x2=70.67 //y2=4.7
cc_4510 ( N_noxref_16_M151_noxref_g N_noxref_21_M150_noxref_d ) capacitor \
 c=0.0180032f //x=73.9 //y=6.02 //x2=73.535 //y2=5.02
cc_4511 ( N_noxref_16_c_5875_n N_noxref_26_c_9912_n ) capacitor c=0.0181982f \
 //x=71.41 //y=2.59 //x2=88.315 //y2=4.07
cc_4512 ( N_noxref_16_c_5876_n N_noxref_26_c_9912_n ) capacitor c=0.019517f \
 //x=73.26 //y=2.08 //x2=88.315 //y2=4.07
cc_4513 ( N_noxref_16_M44_noxref_d N_noxref_56_M42_noxref_s ) capacitor \
 c=0.00309936f //x=70.735 //y=0.915 //x2=67.795 //y2=0.375
cc_4514 ( N_noxref_16_c_5874_n N_noxref_57_c_12024_n ) capacitor c=0.00457167f \
 //x=71.325 //y=1.665 //x2=71.325 //y2=0.54
cc_4515 ( N_noxref_16_M44_noxref_d N_noxref_57_c_12024_n ) capacitor \
 c=0.0115903f //x=70.735 //y=0.915 //x2=71.325 //y2=0.54
cc_4516 ( N_noxref_16_c_5971_p N_noxref_57_c_12034_n ) capacitor c=0.0200405f \
 //x=71.01 //y=1.665 //x2=70.44 //y2=0.995
cc_4517 ( N_noxref_16_M44_noxref_d N_noxref_57_M43_noxref_d ) capacitor \
 c=5.27807e-19 //x=70.735 //y=0.915 //x2=69.2 //y2=0.91
cc_4518 ( N_noxref_16_c_5874_n N_noxref_57_M44_noxref_s ) capacitor \
 c=0.0184051f //x=71.325 //y=1.665 //x2=70.305 //y2=0.375
cc_4519 ( N_noxref_16_M44_noxref_d N_noxref_57_M44_noxref_s ) capacitor \
 c=0.0426368f //x=70.735 //y=0.915 //x2=70.305 //y2=0.375
cc_4520 ( N_noxref_16_c_5874_n N_noxref_58_c_12086_n ) capacitor c=3.84569e-19 \
 //x=71.325 //y=1.665 //x2=72.74 //y2=1.505
cc_4521 ( N_noxref_16_c_5881_n N_noxref_58_c_12086_n ) capacitor c=0.0034165f \
 //x=72.96 //y=1.915 //x2=72.74 //y2=1.505
cc_4522 ( N_noxref_16_c_5876_n N_noxref_58_c_12071_n ) capacitor c=0.0115578f \
 //x=73.26 //y=2.08 //x2=73.625 //y2=1.59
cc_4523 ( N_noxref_16_c_5880_n N_noxref_58_c_12071_n ) capacitor c=0.00697148f \
 //x=72.96 //y=1.53 //x2=73.625 //y2=1.59
cc_4524 ( N_noxref_16_c_5881_n N_noxref_58_c_12071_n ) capacitor c=0.0204849f \
 //x=72.96 //y=1.915 //x2=73.625 //y2=1.59
cc_4525 ( N_noxref_16_c_5883_n N_noxref_58_c_12071_n ) capacitor c=0.00610316f \
 //x=73.335 //y=1.375 //x2=73.625 //y2=1.59
cc_4526 ( N_noxref_16_c_5886_n N_noxref_58_c_12071_n ) capacitor c=0.00698822f \
 //x=73.49 //y=1.22 //x2=73.625 //y2=1.59
cc_4527 ( N_noxref_16_c_5877_n N_noxref_58_M45_noxref_s ) capacitor \
 c=0.0327271f //x=72.96 //y=0.875 //x2=72.605 //y2=0.375
cc_4528 ( N_noxref_16_c_5880_n N_noxref_58_M45_noxref_s ) capacitor \
 c=7.99997e-19 //x=72.96 //y=1.53 //x2=72.605 //y2=0.375
cc_4529 ( N_noxref_16_c_5881_n N_noxref_58_M45_noxref_s ) capacitor \
 c=0.00122123f //x=72.96 //y=1.915 //x2=72.605 //y2=0.375
cc_4530 ( N_noxref_16_c_5884_n N_noxref_58_M45_noxref_s ) capacitor \
 c=0.0121427f //x=73.49 //y=0.875 //x2=72.605 //y2=0.375
cc_4531 ( N_noxref_16_M44_noxref_d N_noxref_58_M45_noxref_s ) capacitor \
 c=2.55333e-19 //x=70.735 //y=0.915 //x2=72.605 //y2=0.375
cc_4532 ( N_CLK_c_6070_n N_noxref_18_c_6814_n ) capacitor c=0.0174051f \
 //x=64.635 //y=4.44 //x2=66.485 //y2=3.33
cc_4533 ( N_CLK_c_6074_n N_noxref_18_c_6814_n ) capacitor c=0.00713821f \
 //x=74.255 //y=4.44 //x2=66.485 //y2=3.33
cc_4534 ( N_CLK_c_6196_n N_noxref_18_c_6814_n ) capacitor c=4.82535e-19 \
 //x=64.865 //y=4.44 //x2=66.485 //y2=3.33
cc_4535 ( N_CLK_c_6044_n N_noxref_18_c_6814_n ) capacitor c=0.0190562f \
 //x=64.75 //y=2.08 //x2=66.485 //y2=3.33
cc_4536 ( N_CLK_c_6070_n N_noxref_18_c_6820_n ) capacitor c=5.79588e-19 \
 //x=64.635 //y=4.44 //x2=61.165 //y2=3.33
cc_4537 ( N_CLK_c_6045_n N_noxref_18_c_6821_n ) capacitor c=0.0190562f \
 //x=74.37 //y=2.08 //x2=77.955 //y2=3.33
cc_4538 ( N_CLK_c_6070_n N_noxref_18_c_6747_n ) capacitor c=0.020183f \
 //x=64.635 //y=4.44 //x2=61.05 //y2=2.08
cc_4539 ( N_CLK_c_6044_n N_noxref_18_c_6762_n ) capacitor c=0.0121898f \
 //x=64.75 //y=2.08 //x2=64.855 //y2=5.155
cc_4540 ( N_CLK_M140_noxref_g N_noxref_18_c_6762_n ) capacitor c=0.0163793f \
 //x=64.72 //y=6.02 //x2=64.855 //y2=5.155
cc_4541 ( N_CLK_c_6217_n N_noxref_18_c_6762_n ) capacitor c=0.00309994f \
 //x=64.75 //y=4.7 //x2=64.855 //y2=5.155
cc_4542 ( N_CLK_M141_noxref_g N_noxref_18_c_6768_n ) capacitor c=0.0162556f \
 //x=65.16 //y=6.02 //x2=65.735 //y2=5.155
cc_4543 ( N_CLK_c_6074_n N_noxref_18_c_6776_n ) capacitor c=0.0166101f \
 //x=74.255 //y=4.44 //x2=66.6 //y2=3.33
cc_4544 ( N_CLK_c_6044_n N_noxref_18_c_6776_n ) capacitor c=0.00248763f \
 //x=64.75 //y=2.08 //x2=66.6 //y2=3.33
cc_4545 ( N_CLK_c_6213_n N_noxref_18_c_6873_n ) capacitor c=0.00392095f \
 //x=65.085 //y=4.79 //x2=64.94 //y2=5.155
cc_4546 ( N_CLK_c_6070_n N_noxref_18_c_6812_n ) capacitor c=0.00731624f \
 //x=64.635 //y=4.44 //x2=61.05 //y2=4.7
cc_4547 ( N_CLK_M140_noxref_g N_noxref_18_M140_noxref_d ) capacitor \
 c=0.0180032f //x=64.72 //y=6.02 //x2=64.795 //y2=5.02
cc_4548 ( N_CLK_M141_noxref_g N_noxref_18_M140_noxref_d ) capacitor \
 c=0.0180032f //x=65.16 //y=6.02 //x2=64.795 //y2=5.02
cc_4549 ( N_CLK_c_6040_n N_RN_c_7021_n ) capacitor c=0.0193884f //x=7.03 \
 //y=2.08 //x2=17.645 //y2=2.22
cc_4550 ( N_CLK_c_6041_n N_RN_c_7021_n ) capacitor c=0.021729f //x=16.65 \
 //y=2.08 //x2=17.645 //y2=2.22
cc_4551 ( N_CLK_c_6129_n N_RN_c_7021_n ) capacitor c=0.00583058f //x=7.12 \
 //y=1.915 //x2=17.645 //y2=2.22
cc_4552 ( N_CLK_c_6158_n N_RN_c_7021_n ) capacitor c=0.00583058f //x=16.74 \
 //y=1.915 //x2=17.645 //y2=2.22
cc_4553 ( N_CLK_c_6041_n N_RN_c_7037_n ) capacitor c=0.00165648f //x=16.65 \
 //y=2.08 //x2=17.875 //y2=2.22
cc_4554 ( N_CLK_c_6158_n N_RN_c_7037_n ) capacitor c=2.3323e-19 //x=16.74 \
 //y=1.915 //x2=17.875 //y2=2.22
cc_4555 ( N_CLK_c_6042_n N_RN_c_7046_n ) capacitor c=0.0193884f //x=35.89 \
 //y=2.08 //x2=46.505 //y2=2.22
cc_4556 ( N_CLK_c_6043_n N_RN_c_7046_n ) capacitor c=0.021729f //x=45.51 \
 //y=2.08 //x2=46.505 //y2=2.22
cc_4557 ( N_CLK_c_6293_n N_RN_c_7046_n ) capacitor c=0.00583058f //x=35.98 \
 //y=1.915 //x2=46.505 //y2=2.22
cc_4558 ( N_CLK_c_6319_n N_RN_c_7046_n ) capacitor c=0.00583058f //x=45.6 \
 //y=1.915 //x2=46.505 //y2=2.22
cc_4559 ( N_CLK_c_6043_n N_RN_c_7062_n ) capacitor c=0.00165648f //x=45.51 \
 //y=2.08 //x2=46.735 //y2=2.22
cc_4560 ( N_CLK_c_6319_n N_RN_c_7062_n ) capacitor c=2.3323e-19 //x=45.6 \
 //y=1.915 //x2=46.735 //y2=2.22
cc_4561 ( N_CLK_c_6044_n N_RN_c_7071_n ) capacitor c=0.0193884f //x=64.75 \
 //y=2.08 //x2=75.365 //y2=2.22
cc_4562 ( N_CLK_c_6045_n N_RN_c_7071_n ) capacitor c=0.021729f //x=74.37 \
 //y=2.08 //x2=75.365 //y2=2.22
cc_4563 ( N_CLK_c_6429_n N_RN_c_7071_n ) capacitor c=0.00583058f //x=64.84 \
 //y=1.915 //x2=75.365 //y2=2.22
cc_4564 ( N_CLK_c_6454_n N_RN_c_7071_n ) capacitor c=0.00583058f //x=74.46 \
 //y=1.915 //x2=75.365 //y2=2.22
cc_4565 ( N_CLK_c_6045_n N_RN_c_7087_n ) capacitor c=0.00165648f //x=74.37 \
 //y=2.08 //x2=75.595 //y2=2.22
cc_4566 ( N_CLK_c_6454_n N_RN_c_7087_n ) capacitor c=2.3323e-19 //x=74.46 \
 //y=1.915 //x2=75.595 //y2=2.22
cc_4567 ( N_CLK_c_6058_n N_RN_c_7089_n ) capacitor c=0.0200057f //x=35.775 \
 //y=4.44 //x2=17.76 //y2=2.08
cc_4568 ( N_CLK_c_6067_n N_RN_c_7089_n ) capacitor c=0.00153281f //x=16.765 \
 //y=4.44 //x2=17.76 //y2=2.08
cc_4569 ( N_CLK_c_6041_n N_RN_c_7089_n ) capacitor c=0.0435729f //x=16.65 \
 //y=2.08 //x2=17.76 //y2=2.08
cc_4570 ( N_CLK_c_6158_n N_RN_c_7089_n ) capacitor c=0.00203728f //x=16.74 \
 //y=1.915 //x2=17.76 //y2=2.08
cc_4571 ( N_CLK_c_6160_n N_RN_c_7089_n ) capacitor c=0.00142741f //x=16.65 \
 //y=4.7 //x2=17.76 //y2=2.08
cc_4572 ( N_CLK_c_6058_n N_RN_c_7090_n ) capacitor c=0.0210462f //x=35.775 \
 //y=4.44 //x2=21.46 //y2=2.08
cc_4573 ( N_CLK_c_6058_n N_RN_c_7091_n ) capacitor c=0.0188829f //x=35.775 \
 //y=4.44 //x2=31.08 //y2=2.08
cc_4574 ( N_CLK_c_6070_n N_RN_c_7092_n ) capacitor c=0.0178424f //x=64.635 \
 //y=4.44 //x2=46.62 //y2=2.08
cc_4575 ( N_CLK_c_6192_n N_RN_c_7092_n ) capacitor c=0.00153281f //x=45.625 \
 //y=4.44 //x2=46.62 //y2=2.08
cc_4576 ( N_CLK_c_6043_n N_RN_c_7092_n ) capacitor c=0.0416369f //x=45.51 \
 //y=2.08 //x2=46.62 //y2=2.08
cc_4577 ( N_CLK_c_6319_n N_RN_c_7092_n ) capacitor c=0.00203728f //x=45.6 \
 //y=1.915 //x2=46.62 //y2=2.08
cc_4578 ( N_CLK_c_6216_n N_RN_c_7092_n ) capacitor c=0.00142741f //x=45.51 \
 //y=4.7 //x2=46.62 //y2=2.08
cc_4579 ( N_CLK_c_6070_n N_RN_c_7093_n ) capacitor c=0.0188829f //x=64.635 \
 //y=4.44 //x2=50.32 //y2=2.08
cc_4580 ( N_CLK_c_6070_n N_RN_c_7094_n ) capacitor c=0.0212234f //x=64.635 \
 //y=4.44 //x2=59.94 //y2=2.08
cc_4581 ( N_CLK_c_6074_n N_RN_c_7095_n ) capacitor c=0.00163971f //x=74.255 \
 //y=4.44 //x2=75.48 //y2=2.08
cc_4582 ( N_CLK_c_6045_n N_RN_c_7095_n ) capacitor c=0.0407128f //x=74.37 \
 //y=2.08 //x2=75.48 //y2=2.08
cc_4583 ( N_CLK_c_6454_n N_RN_c_7095_n ) capacitor c=0.00203728f //x=74.46 \
 //y=1.915 //x2=75.48 //y2=2.08
cc_4584 ( N_CLK_c_6218_n N_RN_c_7095_n ) capacitor c=0.00142741f //x=74.37 \
 //y=4.7 //x2=75.48 //y2=2.08
cc_4585 ( N_CLK_M80_noxref_g N_RN_M82_noxref_g ) capacitor c=0.0101598f \
 //x=16.62 //y=6.02 //x2=17.5 //y2=6.02
cc_4586 ( N_CLK_M81_noxref_g N_RN_M82_noxref_g ) capacitor c=0.0602553f \
 //x=17.06 //y=6.02 //x2=17.5 //y2=6.02
cc_4587 ( N_CLK_M81_noxref_g N_RN_M83_noxref_g ) capacitor c=0.0101598f \
 //x=17.06 //y=6.02 //x2=17.94 //y2=6.02
cc_4588 ( N_CLK_M116_noxref_g N_RN_M118_noxref_g ) capacitor c=0.0100903f \
 //x=45.48 //y=6.02 //x2=46.36 //y2=6.02
cc_4589 ( N_CLK_M117_noxref_g N_RN_M118_noxref_g ) capacitor c=0.0600064f \
 //x=45.92 //y=6.02 //x2=46.36 //y2=6.02
cc_4590 ( N_CLK_M117_noxref_g N_RN_M119_noxref_g ) capacitor c=0.0100903f \
 //x=45.92 //y=6.02 //x2=46.8 //y2=6.02
cc_4591 ( N_CLK_M152_noxref_g N_RN_M154_noxref_g ) capacitor c=0.0100903f \
 //x=74.34 //y=6.02 //x2=75.22 //y2=6.02
cc_4592 ( N_CLK_M153_noxref_g N_RN_M154_noxref_g ) capacitor c=0.0599334f \
 //x=74.78 //y=6.02 //x2=75.22 //y2=6.02
cc_4593 ( N_CLK_M153_noxref_g N_RN_M155_noxref_g ) capacitor c=0.0101723f \
 //x=74.78 //y=6.02 //x2=75.66 //y2=6.02
cc_4594 ( N_CLK_c_6155_n N_RN_c_7295_n ) capacitor c=0.00456962f //x=16.74 \
 //y=0.91 //x2=17.75 //y2=0.915
cc_4595 ( N_CLK_c_6156_n N_RN_c_7296_n ) capacitor c=0.00438372f //x=16.74 \
 //y=1.22 //x2=17.75 //y2=1.26
cc_4596 ( N_CLK_c_6157_n N_RN_c_7297_n ) capacitor c=0.00438372f //x=16.74 \
 //y=1.45 //x2=17.75 //y2=1.57
cc_4597 ( N_CLK_c_6058_n N_RN_c_7255_n ) capacitor c=0.0085986f //x=35.775 \
 //y=4.44 //x2=21.795 //y2=4.79
cc_4598 ( N_CLK_c_6058_n N_RN_c_7256_n ) capacitor c=0.00554824f //x=35.775 \
 //y=4.44 //x2=31.415 //y2=4.79
cc_4599 ( N_CLK_c_6316_n N_RN_c_7441_n ) capacitor c=0.00456962f //x=45.6 \
 //y=0.91 //x2=46.61 //y2=0.915
cc_4600 ( N_CLK_c_6317_n N_RN_c_7442_n ) capacitor c=0.00438372f //x=45.6 \
 //y=1.22 //x2=46.61 //y2=1.26
cc_4601 ( N_CLK_c_6318_n N_RN_c_7443_n ) capacitor c=0.00438372f //x=45.6 \
 //y=1.45 //x2=46.61 //y2=1.57
cc_4602 ( N_CLK_c_6070_n N_RN_c_7257_n ) capacitor c=0.00554824f //x=64.635 \
 //y=4.44 //x2=50.655 //y2=4.79
cc_4603 ( N_CLK_c_6070_n N_RN_c_7258_n ) capacitor c=0.00554824f //x=64.635 \
 //y=4.44 //x2=60.275 //y2=4.79
cc_4604 ( N_CLK_c_6451_n N_RN_c_7649_n ) capacitor c=0.00456962f //x=74.46 \
 //y=0.91 //x2=75.47 //y2=0.915
cc_4605 ( N_CLK_c_6452_n N_RN_c_7650_n ) capacitor c=0.00438372f //x=74.46 \
 //y=1.22 //x2=75.47 //y2=1.26
cc_4606 ( N_CLK_c_6453_n N_RN_c_7651_n ) capacitor c=0.00438372f //x=74.46 \
 //y=1.45 //x2=75.47 //y2=1.57
cc_4607 ( N_CLK_c_6041_n N_RN_c_7304_n ) capacitor c=0.00201097f //x=16.65 \
 //y=2.08 //x2=17.76 //y2=2.08
cc_4608 ( N_CLK_c_6158_n N_RN_c_7304_n ) capacitor c=0.00828003f //x=16.74 \
 //y=1.915 //x2=17.76 //y2=2.08
cc_4609 ( N_CLK_c_6158_n N_RN_c_7305_n ) capacitor c=0.00438372f //x=16.74 \
 //y=1.915 //x2=17.76 //y2=1.915
cc_4610 ( N_CLK_c_6058_n N_RN_c_7307_n ) capacitor c=0.0111881f //x=35.775 \
 //y=4.44 //x2=17.76 //y2=4.7
cc_4611 ( N_CLK_c_6041_n N_RN_c_7307_n ) capacitor c=0.00218014f //x=16.65 \
 //y=2.08 //x2=17.76 //y2=4.7
cc_4612 ( N_CLK_c_6261_n N_RN_c_7307_n ) capacitor c=0.0611812f //x=16.985 \
 //y=4.79 //x2=17.76 //y2=4.7
cc_4613 ( N_CLK_c_6160_n N_RN_c_7307_n ) capacitor c=0.00487508f //x=16.65 \
 //y=4.7 //x2=17.76 //y2=4.7
cc_4614 ( N_CLK_c_6058_n N_RN_c_7223_n ) capacitor c=0.00293313f //x=35.775 \
 //y=4.44 //x2=21.46 //y2=4.7
cc_4615 ( N_CLK_c_6058_n N_RN_c_7261_n ) capacitor c=0.00187486f //x=35.775 \
 //y=4.44 //x2=31.08 //y2=4.7
cc_4616 ( N_CLK_c_6043_n N_RN_c_7450_n ) capacitor c=0.00201097f //x=45.51 \
 //y=2.08 //x2=46.62 //y2=2.08
cc_4617 ( N_CLK_c_6319_n N_RN_c_7450_n ) capacitor c=0.00828003f //x=45.6 \
 //y=1.915 //x2=46.62 //y2=2.08
cc_4618 ( N_CLK_c_6319_n N_RN_c_7451_n ) capacitor c=0.00438372f //x=45.6 \
 //y=1.915 //x2=46.62 //y2=1.915
cc_4619 ( N_CLK_c_6070_n N_RN_c_7262_n ) capacitor c=0.00731624f //x=64.635 \
 //y=4.44 //x2=46.62 //y2=4.7
cc_4620 ( N_CLK_c_6043_n N_RN_c_7262_n ) capacitor c=0.00196431f //x=45.51 \
 //y=2.08 //x2=46.62 //y2=4.7
cc_4621 ( N_CLK_c_6212_n N_RN_c_7262_n ) capacitor c=0.0609323f //x=45.845 \
 //y=4.79 //x2=46.62 //y2=4.7
cc_4622 ( N_CLK_c_6216_n N_RN_c_7262_n ) capacitor c=0.00487508f //x=45.51 \
 //y=4.7 //x2=46.62 //y2=4.7
cc_4623 ( N_CLK_c_6070_n N_RN_c_7263_n ) capacitor c=0.00187486f //x=64.635 \
 //y=4.44 //x2=50.32 //y2=4.7
cc_4624 ( N_CLK_c_6070_n N_RN_c_7264_n ) capacitor c=0.00187486f //x=64.635 \
 //y=4.44 //x2=59.94 //y2=4.7
cc_4625 ( N_CLK_c_6045_n N_RN_c_7670_n ) capacitor c=0.00201097f //x=74.37 \
 //y=2.08 //x2=75.48 //y2=2.08
cc_4626 ( N_CLK_c_6454_n N_RN_c_7670_n ) capacitor c=0.00828003f //x=74.46 \
 //y=1.915 //x2=75.48 //y2=2.08
cc_4627 ( N_CLK_c_6454_n N_RN_c_7672_n ) capacitor c=0.00438372f //x=74.46 \
 //y=1.915 //x2=75.48 //y2=1.915
cc_4628 ( N_CLK_c_6045_n N_RN_c_7265_n ) capacitor c=0.0019552f //x=74.37 \
 //y=2.08 //x2=75.48 //y2=4.7
cc_4629 ( N_CLK_c_6214_n N_RN_c_7265_n ) capacitor c=0.0608593f //x=74.705 \
 //y=4.79 //x2=75.48 //y2=4.7
cc_4630 ( N_CLK_c_6218_n N_RN_c_7265_n ) capacitor c=0.00484771f //x=74.37 \
 //y=4.7 //x2=75.48 //y2=4.7
cc_4631 ( N_CLK_c_6041_n N_SN_c_8129_n ) capacitor c=0.021326f //x=16.65 \
 //y=2.08 //x2=26.155 //y2=2.96
cc_4632 ( N_CLK_c_6058_n N_SN_c_8132_n ) capacitor c=0.0181287f //x=35.775 \
 //y=4.44 //x2=40.585 //y2=2.96
cc_4633 ( N_CLK_c_6042_n N_SN_c_8132_n ) capacitor c=0.0190322f //x=35.89 \
 //y=2.08 //x2=40.585 //y2=2.96
cc_4634 ( N_CLK_c_6043_n N_SN_c_8135_n ) capacitor c=0.021326f //x=45.51 \
 //y=2.08 //x2=55.015 //y2=2.96
cc_4635 ( N_CLK_c_6070_n N_SN_c_8138_n ) capacitor c=0.0086541f //x=64.635 \
 //y=4.44 //x2=69.445 //y2=2.96
cc_4636 ( N_CLK_c_6044_n N_SN_c_8138_n ) capacitor c=0.0190322f //x=64.75 \
 //y=2.08 //x2=69.445 //y2=2.96
cc_4637 ( N_CLK_c_6045_n N_SN_c_8141_n ) capacitor c=0.021326f //x=74.37 \
 //y=2.08 //x2=83.875 //y2=2.96
cc_4638 ( N_CLK_c_6046_n N_SN_c_8145_n ) capacitor c=0.0210462f //x=16.535 \
 //y=4.44 //x2=11.84 //y2=2.08
cc_4639 ( N_CLK_c_6058_n N_SN_c_8146_n ) capacitor c=0.0188829f //x=35.775 \
 //y=4.44 //x2=26.27 //y2=2.08
cc_4640 ( N_CLK_c_6068_n N_SN_c_8147_n ) capacitor c=0.0188829f //x=45.395 \
 //y=4.44 //x2=40.7 //y2=2.08
cc_4641 ( N_CLK_c_6070_n N_SN_c_8148_n ) capacitor c=0.0188829f //x=64.635 \
 //y=4.44 //x2=55.13 //y2=2.08
cc_4642 ( N_CLK_c_6074_n N_SN_c_8149_n ) capacitor c=0.0188829f //x=74.255 \
 //y=4.44 //x2=69.56 //y2=2.08
cc_4643 ( N_CLK_c_6046_n N_SN_c_8215_n ) capacitor c=0.0085986f //x=16.535 \
 //y=4.44 //x2=12.175 //y2=4.79
cc_4644 ( N_CLK_c_6058_n N_SN_c_8259_n ) capacitor c=0.00554824f //x=35.775 \
 //y=4.44 //x2=26.605 //y2=4.79
cc_4645 ( N_CLK_c_6068_n N_SN_c_8260_n ) capacitor c=0.00554824f //x=45.395 \
 //y=4.44 //x2=41.035 //y2=4.79
cc_4646 ( N_CLK_c_6070_n N_SN_c_8261_n ) capacitor c=0.00554824f //x=64.635 \
 //y=4.44 //x2=55.465 //y2=4.79
cc_4647 ( N_CLK_c_6074_n N_SN_c_8262_n ) capacitor c=0.00554824f //x=74.255 \
 //y=4.44 //x2=69.895 //y2=4.79
cc_4648 ( N_CLK_c_6046_n N_SN_c_8202_n ) capacitor c=0.00293313f //x=16.535 \
 //y=4.44 //x2=11.84 //y2=4.7
cc_4649 ( N_CLK_c_6058_n N_SN_c_8264_n ) capacitor c=0.00187486f //x=35.775 \
 //y=4.44 //x2=26.27 //y2=4.7
cc_4650 ( N_CLK_c_6068_n N_SN_c_8268_n ) capacitor c=0.00187486f //x=45.395 \
 //y=4.44 //x2=40.7 //y2=4.7
cc_4651 ( N_CLK_c_6070_n N_SN_c_8269_n ) capacitor c=0.00187486f //x=64.635 \
 //y=4.44 //x2=55.13 //y2=4.7
cc_4652 ( N_CLK_c_6074_n N_SN_c_8270_n ) capacitor c=0.00187486f //x=74.255 \
 //y=4.44 //x2=69.56 //y2=4.7
cc_4653 ( N_CLK_c_6074_n N_noxref_21_c_8898_n ) capacitor c=0.0344845f \
 //x=74.255 //y=4.44 //x2=70.555 //y2=3.7
cc_4654 ( N_CLK_c_6074_n N_noxref_21_c_8935_n ) capacitor c=7.0371e-19 \
 //x=74.255 //y=4.44 //x2=65.975 //y2=3.7
cc_4655 ( N_CLK_c_6044_n N_noxref_21_c_8935_n ) capacitor c=0.00163582f \
 //x=64.75 //y=2.08 //x2=65.975 //y2=3.7
cc_4656 ( N_CLK_c_6074_n N_noxref_21_c_8878_n ) capacitor c=0.0256468f \
 //x=74.255 //y=4.44 //x2=76.105 //y2=3.7
cc_4657 ( N_CLK_c_6045_n N_noxref_21_c_8878_n ) capacitor c=0.0190398f \
 //x=74.37 //y=2.08 //x2=76.105 //y2=3.7
cc_4658 ( N_CLK_c_6074_n N_noxref_21_c_8905_n ) capacitor c=4.78625e-19 \
 //x=74.255 //y=4.44 //x2=70.785 //y2=3.7
cc_4659 ( N_CLK_c_6074_n N_noxref_21_c_8828_n ) capacitor c=0.0178424f \
 //x=74.255 //y=4.44 //x2=65.86 //y2=2.08
cc_4660 ( N_CLK_c_6196_n N_noxref_21_c_8828_n ) capacitor c=0.00153281f \
 //x=64.865 //y=4.44 //x2=65.86 //y2=2.08
cc_4661 ( N_CLK_c_6044_n N_noxref_21_c_8828_n ) capacitor c=0.0396012f \
 //x=64.75 //y=2.08 //x2=65.86 //y2=2.08
cc_4662 ( N_CLK_c_6429_n N_noxref_21_c_8828_n ) capacitor c=0.00205895f \
 //x=64.84 //y=1.915 //x2=65.86 //y2=2.08
cc_4663 ( N_CLK_c_6217_n N_noxref_21_c_8828_n ) capacitor c=0.00142741f \
 //x=64.75 //y=4.7 //x2=65.86 //y2=2.08
cc_4664 ( N_CLK_c_6074_n N_noxref_21_c_8829_n ) capacitor c=0.0178424f \
 //x=74.255 //y=4.44 //x2=70.67 //y2=2.08
cc_4665 ( N_CLK_c_6045_n N_noxref_21_c_8835_n ) capacitor c=0.0121898f \
 //x=74.37 //y=2.08 //x2=74.475 //y2=5.155
cc_4666 ( N_CLK_M152_noxref_g N_noxref_21_c_8835_n ) capacitor c=0.0163793f \
 //x=74.34 //y=6.02 //x2=74.475 //y2=5.155
cc_4667 ( N_CLK_c_6218_n N_noxref_21_c_8835_n ) capacitor c=0.00309994f \
 //x=74.37 //y=4.7 //x2=74.475 //y2=5.155
cc_4668 ( N_CLK_M153_noxref_g N_noxref_21_c_8841_n ) capacitor c=0.0162556f \
 //x=74.78 //y=6.02 //x2=75.355 //y2=5.155
cc_4669 ( N_CLK_c_6045_n N_noxref_21_c_8849_n ) capacitor c=0.00251642f \
 //x=74.37 //y=2.08 //x2=76.22 //y2=3.7
cc_4670 ( N_CLK_c_6214_n N_noxref_21_c_8951_n ) capacitor c=0.00392095f \
 //x=74.705 //y=4.79 //x2=74.56 //y2=5.155
cc_4671 ( N_CLK_M140_noxref_g N_noxref_21_M142_noxref_g ) capacitor \
 c=0.0100903f //x=64.72 //y=6.02 //x2=65.6 //y2=6.02
cc_4672 ( N_CLK_M141_noxref_g N_noxref_21_M142_noxref_g ) capacitor \
 c=0.0600064f //x=65.16 //y=6.02 //x2=65.6 //y2=6.02
cc_4673 ( N_CLK_M141_noxref_g N_noxref_21_M143_noxref_g ) capacitor \
 c=0.0100903f //x=65.16 //y=6.02 //x2=66.04 //y2=6.02
cc_4674 ( N_CLK_c_6426_n N_noxref_21_c_8955_n ) capacitor c=0.00456962f \
 //x=64.84 //y=0.91 //x2=65.85 //y2=0.915
cc_4675 ( N_CLK_c_6427_n N_noxref_21_c_8956_n ) capacitor c=0.00438372f \
 //x=64.84 //y=1.22 //x2=65.85 //y2=1.26
cc_4676 ( N_CLK_c_6428_n N_noxref_21_c_8957_n ) capacitor c=0.00438372f \
 //x=64.84 //y=1.45 //x2=65.85 //y2=1.57
cc_4677 ( N_CLK_c_6044_n N_noxref_21_c_8958_n ) capacitor c=0.00201097f \
 //x=64.75 //y=2.08 //x2=65.86 //y2=2.08
cc_4678 ( N_CLK_c_6429_n N_noxref_21_c_8958_n ) capacitor c=0.00828003f \
 //x=64.84 //y=1.915 //x2=65.86 //y2=2.08
cc_4679 ( N_CLK_c_6429_n N_noxref_21_c_8960_n ) capacitor c=0.00438372f \
 //x=64.84 //y=1.915 //x2=65.86 //y2=1.915
cc_4680 ( N_CLK_c_6074_n N_noxref_21_c_8895_n ) capacitor c=0.00731624f \
 //x=74.255 //y=4.44 //x2=65.86 //y2=4.7
cc_4681 ( N_CLK_c_6044_n N_noxref_21_c_8895_n ) capacitor c=0.00196431f \
 //x=64.75 //y=2.08 //x2=65.86 //y2=4.7
cc_4682 ( N_CLK_c_6213_n N_noxref_21_c_8895_n ) capacitor c=0.0609323f \
 //x=65.085 //y=4.79 //x2=65.86 //y2=4.7
cc_4683 ( N_CLK_c_6217_n N_noxref_21_c_8895_n ) capacitor c=0.00487508f \
 //x=64.75 //y=4.7 //x2=65.86 //y2=4.7
cc_4684 ( N_CLK_c_6074_n N_noxref_21_c_8896_n ) capacitor c=0.00731624f \
 //x=74.255 //y=4.44 //x2=70.67 //y2=4.7
cc_4685 ( N_CLK_M152_noxref_g N_noxref_21_M152_noxref_d ) capacitor \
 c=0.0180032f //x=74.34 //y=6.02 //x2=74.415 //y2=5.02
cc_4686 ( N_CLK_M153_noxref_g N_noxref_21_M152_noxref_d ) capacitor \
 c=0.0180032f //x=74.78 //y=6.02 //x2=74.415 //y2=5.02
cc_4687 ( N_CLK_c_6070_n N_noxref_26_c_10050_n ) capacitor c=0.00392792f \
 //x=64.635 //y=4.44 //x2=56.895 //y2=3.33
cc_4688 ( N_CLK_c_6070_n N_noxref_26_c_9933_n ) capacitor c=0.249854f \
 //x=64.635 //y=4.44 //x2=65.035 //y2=3.7
cc_4689 ( N_CLK_c_6074_n N_noxref_26_c_9933_n ) capacitor c=0.00708979f \
 //x=74.255 //y=4.44 //x2=65.035 //y2=3.7
cc_4690 ( N_CLK_c_6196_n N_noxref_26_c_9933_n ) capacitor c=0.0120266f \
 //x=64.865 //y=4.44 //x2=65.035 //y2=3.7
cc_4691 ( N_CLK_c_6044_n N_noxref_26_c_9933_n ) capacitor c=0.0208267f \
 //x=64.75 //y=2.08 //x2=65.035 //y2=3.7
cc_4692 ( N_CLK_c_6044_n N_noxref_26_c_10119_n ) capacitor c=0.0165481f \
 //x=64.75 //y=2.08 //x2=65.12 //y2=3.985
cc_4693 ( N_CLK_c_6074_n N_noxref_26_c_9912_n ) capacitor c=0.0291328f \
 //x=74.255 //y=4.44 //x2=88.315 //y2=4.07
cc_4694 ( N_CLK_c_6045_n N_noxref_26_c_9912_n ) capacitor c=0.0208526f \
 //x=74.37 //y=2.08 //x2=88.315 //y2=4.07
cc_4695 ( N_CLK_c_6214_n N_noxref_26_c_9912_n ) capacitor c=0.00478828f \
 //x=74.705 //y=4.79 //x2=88.315 //y2=4.07
cc_4696 ( N_CLK_c_6074_n N_noxref_26_c_10001_n ) capacitor c=0.802413f \
 //x=74.255 //y=4.44 //x2=65.205 //y2=4.07
cc_4697 ( N_CLK_c_6070_n N_noxref_26_c_9958_n ) capacitor c=0.0166101f \
 //x=64.635 //y=4.44 //x2=52.17 //y2=3.33
cc_4698 ( N_CLK_c_6070_n N_noxref_26_c_9916_n ) capacitor c=0.018786f \
 //x=64.635 //y=4.44 //x2=54.02 //y2=2.08
cc_4699 ( N_CLK_c_6070_n N_noxref_26_c_9977_n ) capacitor c=0.0112124f \
 //x=64.635 //y=4.44 //x2=54.295 //y2=4.79
cc_4700 ( N_CLK_c_6121_n N_noxref_30_c_10650_n ) capacitor c=0.0167228f \
 //x=6.595 //y=0.91 //x2=7.255 //y2=0.54
cc_4701 ( N_CLK_c_6126_n N_noxref_30_c_10650_n ) capacitor c=0.00534519f \
 //x=7.12 //y=0.91 //x2=7.255 //y2=0.54
cc_4702 ( N_CLK_c_6040_n N_noxref_30_c_10673_n ) capacitor c=0.0117694f \
 //x=7.03 //y=2.08 //x2=7.255 //y2=1.59
cc_4703 ( N_CLK_c_6124_n N_noxref_30_c_10673_n ) capacitor c=0.0157358f \
 //x=6.595 //y=1.22 //x2=7.255 //y2=1.59
cc_4704 ( N_CLK_c_6129_n N_noxref_30_c_10673_n ) capacitor c=0.021347f \
 //x=7.12 //y=1.915 //x2=7.255 //y2=1.59
cc_4705 ( N_CLK_c_6121_n N_noxref_30_M3_noxref_s ) capacitor c=0.00798959f \
 //x=6.595 //y=0.91 //x2=5.265 //y2=0.375
cc_4706 ( N_CLK_c_6128_n N_noxref_30_M3_noxref_s ) capacitor c=0.00212176f \
 //x=7.12 //y=1.45 //x2=5.265 //y2=0.375
cc_4707 ( N_CLK_c_6129_n N_noxref_30_M3_noxref_s ) capacitor c=0.00298115f \
 //x=7.12 //y=1.915 //x2=5.265 //y2=0.375
cc_4708 ( N_CLK_c_6635_p N_noxref_31_c_10692_n ) capacitor c=2.14837e-19 \
 //x=6.965 //y=0.755 //x2=7.825 //y2=0.995
cc_4709 ( N_CLK_c_6126_n N_noxref_31_c_10692_n ) capacitor c=0.00123426f \
 //x=7.12 //y=0.91 //x2=7.825 //y2=0.995
cc_4710 ( N_CLK_c_6127_n N_noxref_31_c_10692_n ) capacitor c=0.0129288f \
 //x=7.12 //y=1.22 //x2=7.825 //y2=0.995
cc_4711 ( N_CLK_c_6128_n N_noxref_31_c_10692_n ) capacitor c=0.00142359f \
 //x=7.12 //y=1.45 //x2=7.825 //y2=0.995
cc_4712 ( N_CLK_c_6121_n N_noxref_31_M4_noxref_d ) capacitor c=0.00223875f \
 //x=6.595 //y=0.91 //x2=6.67 //y2=0.91
cc_4713 ( N_CLK_c_6124_n N_noxref_31_M4_noxref_d ) capacitor c=0.00262485f \
 //x=6.595 //y=1.22 //x2=6.67 //y2=0.91
cc_4714 ( N_CLK_c_6635_p N_noxref_31_M4_noxref_d ) capacitor c=0.00220746f \
 //x=6.965 //y=0.755 //x2=6.67 //y2=0.91
cc_4715 ( N_CLK_c_6642_p N_noxref_31_M4_noxref_d ) capacitor c=0.00194798f \
 //x=6.965 //y=1.375 //x2=6.67 //y2=0.91
cc_4716 ( N_CLK_c_6126_n N_noxref_31_M4_noxref_d ) capacitor c=0.00198465f \
 //x=7.12 //y=0.91 //x2=6.67 //y2=0.91
cc_4717 ( N_CLK_c_6127_n N_noxref_31_M4_noxref_d ) capacitor c=0.00128384f \
 //x=7.12 //y=1.22 //x2=6.67 //y2=0.91
cc_4718 ( N_CLK_c_6126_n N_noxref_31_M5_noxref_s ) capacitor c=7.21316e-19 \
 //x=7.12 //y=0.91 //x2=7.775 //y2=0.375
cc_4719 ( N_CLK_c_6127_n N_noxref_31_M5_noxref_s ) capacitor c=0.00348171f \
 //x=7.12 //y=1.22 //x2=7.775 //y2=0.375
cc_4720 ( N_CLK_c_6150_n N_noxref_34_c_10852_n ) capacitor c=0.0167228f \
 //x=16.215 //y=0.91 //x2=16.875 //y2=0.54
cc_4721 ( N_CLK_c_6155_n N_noxref_34_c_10852_n ) capacitor c=0.00534519f \
 //x=16.74 //y=0.91 //x2=16.875 //y2=0.54
cc_4722 ( N_CLK_c_6041_n N_noxref_34_c_10875_n ) capacitor c=0.0117694f \
 //x=16.65 //y=2.08 //x2=16.875 //y2=1.59
cc_4723 ( N_CLK_c_6153_n N_noxref_34_c_10875_n ) capacitor c=0.0157358f \
 //x=16.215 //y=1.22 //x2=16.875 //y2=1.59
cc_4724 ( N_CLK_c_6158_n N_noxref_34_c_10875_n ) capacitor c=0.021347f \
 //x=16.74 //y=1.915 //x2=16.875 //y2=1.59
cc_4725 ( N_CLK_c_6150_n N_noxref_34_M9_noxref_s ) capacitor c=0.00798959f \
 //x=16.215 //y=0.91 //x2=14.885 //y2=0.375
cc_4726 ( N_CLK_c_6157_n N_noxref_34_M9_noxref_s ) capacitor c=0.00212176f \
 //x=16.74 //y=1.45 //x2=14.885 //y2=0.375
cc_4727 ( N_CLK_c_6158_n N_noxref_34_M9_noxref_s ) capacitor c=0.00298115f \
 //x=16.74 //y=1.915 //x2=14.885 //y2=0.375
cc_4728 ( N_CLK_c_6655_p N_noxref_35_c_10894_n ) capacitor c=2.14837e-19 \
 //x=16.585 //y=0.755 //x2=17.445 //y2=0.995
cc_4729 ( N_CLK_c_6155_n N_noxref_35_c_10894_n ) capacitor c=0.00123426f \
 //x=16.74 //y=0.91 //x2=17.445 //y2=0.995
cc_4730 ( N_CLK_c_6156_n N_noxref_35_c_10894_n ) capacitor c=0.0129288f \
 //x=16.74 //y=1.22 //x2=17.445 //y2=0.995
cc_4731 ( N_CLK_c_6157_n N_noxref_35_c_10894_n ) capacitor c=0.00142359f \
 //x=16.74 //y=1.45 //x2=17.445 //y2=0.995
cc_4732 ( N_CLK_c_6150_n N_noxref_35_M10_noxref_d ) capacitor c=0.00223875f \
 //x=16.215 //y=0.91 //x2=16.29 //y2=0.91
cc_4733 ( N_CLK_c_6153_n N_noxref_35_M10_noxref_d ) capacitor c=0.00262485f \
 //x=16.215 //y=1.22 //x2=16.29 //y2=0.91
cc_4734 ( N_CLK_c_6655_p N_noxref_35_M10_noxref_d ) capacitor c=0.00220746f \
 //x=16.585 //y=0.755 //x2=16.29 //y2=0.91
cc_4735 ( N_CLK_c_6662_p N_noxref_35_M10_noxref_d ) capacitor c=0.00194798f \
 //x=16.585 //y=1.375 //x2=16.29 //y2=0.91
cc_4736 ( N_CLK_c_6155_n N_noxref_35_M10_noxref_d ) capacitor c=0.00198465f \
 //x=16.74 //y=0.91 //x2=16.29 //y2=0.91
cc_4737 ( N_CLK_c_6156_n N_noxref_35_M10_noxref_d ) capacitor c=0.00128384f \
 //x=16.74 //y=1.22 //x2=16.29 //y2=0.91
cc_4738 ( N_CLK_c_6155_n N_noxref_35_M11_noxref_s ) capacitor c=7.21316e-19 \
 //x=16.74 //y=0.91 //x2=17.395 //y2=0.375
cc_4739 ( N_CLK_c_6156_n N_noxref_35_M11_noxref_s ) capacitor c=0.00348171f \
 //x=16.74 //y=1.22 //x2=17.395 //y2=0.375
cc_4740 ( N_CLK_c_6285_n N_noxref_42_c_11263_n ) capacitor c=0.0167228f \
 //x=35.455 //y=0.91 //x2=36.115 //y2=0.54
cc_4741 ( N_CLK_c_6290_n N_noxref_42_c_11263_n ) capacitor c=0.00534519f \
 //x=35.98 //y=0.91 //x2=36.115 //y2=0.54
cc_4742 ( N_CLK_c_6042_n N_noxref_42_c_11286_n ) capacitor c=0.0120267f \
 //x=35.89 //y=2.08 //x2=36.115 //y2=1.59
cc_4743 ( N_CLK_c_6288_n N_noxref_42_c_11286_n ) capacitor c=0.0157358f \
 //x=35.455 //y=1.22 //x2=36.115 //y2=1.59
cc_4744 ( N_CLK_c_6293_n N_noxref_42_c_11286_n ) capacitor c=0.021347f \
 //x=35.98 //y=1.915 //x2=36.115 //y2=1.59
cc_4745 ( N_CLK_c_6285_n N_noxref_42_M21_noxref_s ) capacitor c=0.00798959f \
 //x=35.455 //y=0.91 //x2=34.125 //y2=0.375
cc_4746 ( N_CLK_c_6292_n N_noxref_42_M21_noxref_s ) capacitor c=0.00212176f \
 //x=35.98 //y=1.45 //x2=34.125 //y2=0.375
cc_4747 ( N_CLK_c_6293_n N_noxref_42_M21_noxref_s ) capacitor c=0.00298115f \
 //x=35.98 //y=1.915 //x2=34.125 //y2=0.375
cc_4748 ( N_CLK_c_6675_p N_noxref_43_c_11305_n ) capacitor c=2.14837e-19 \
 //x=35.825 //y=0.755 //x2=36.685 //y2=0.995
cc_4749 ( N_CLK_c_6290_n N_noxref_43_c_11305_n ) capacitor c=0.00123426f \
 //x=35.98 //y=0.91 //x2=36.685 //y2=0.995
cc_4750 ( N_CLK_c_6291_n N_noxref_43_c_11305_n ) capacitor c=0.0129288f \
 //x=35.98 //y=1.22 //x2=36.685 //y2=0.995
cc_4751 ( N_CLK_c_6292_n N_noxref_43_c_11305_n ) capacitor c=0.00142359f \
 //x=35.98 //y=1.45 //x2=36.685 //y2=0.995
cc_4752 ( N_CLK_c_6285_n N_noxref_43_M22_noxref_d ) capacitor c=0.00223875f \
 //x=35.455 //y=0.91 //x2=35.53 //y2=0.91
cc_4753 ( N_CLK_c_6288_n N_noxref_43_M22_noxref_d ) capacitor c=0.00262485f \
 //x=35.455 //y=1.22 //x2=35.53 //y2=0.91
cc_4754 ( N_CLK_c_6675_p N_noxref_43_M22_noxref_d ) capacitor c=0.00220746f \
 //x=35.825 //y=0.755 //x2=35.53 //y2=0.91
cc_4755 ( N_CLK_c_6682_p N_noxref_43_M22_noxref_d ) capacitor c=0.00194798f \
 //x=35.825 //y=1.375 //x2=35.53 //y2=0.91
cc_4756 ( N_CLK_c_6290_n N_noxref_43_M22_noxref_d ) capacitor c=0.00198465f \
 //x=35.98 //y=0.91 //x2=35.53 //y2=0.91
cc_4757 ( N_CLK_c_6291_n N_noxref_43_M22_noxref_d ) capacitor c=0.00128384f \
 //x=35.98 //y=1.22 //x2=35.53 //y2=0.91
cc_4758 ( N_CLK_c_6290_n N_noxref_43_M23_noxref_s ) capacitor c=7.21316e-19 \
 //x=35.98 //y=0.91 //x2=36.635 //y2=0.375
cc_4759 ( N_CLK_c_6291_n N_noxref_43_M23_noxref_s ) capacitor c=0.00348171f \
 //x=35.98 //y=1.22 //x2=36.635 //y2=0.375
cc_4760 ( N_CLK_c_6311_n N_noxref_46_c_11465_n ) capacitor c=0.0167228f \
 //x=45.075 //y=0.91 //x2=45.735 //y2=0.54
cc_4761 ( N_CLK_c_6316_n N_noxref_46_c_11465_n ) capacitor c=0.00534519f \
 //x=45.6 //y=0.91 //x2=45.735 //y2=0.54
cc_4762 ( N_CLK_c_6043_n N_noxref_46_c_11488_n ) capacitor c=0.0120267f \
 //x=45.51 //y=2.08 //x2=45.735 //y2=1.59
cc_4763 ( N_CLK_c_6314_n N_noxref_46_c_11488_n ) capacitor c=0.0157358f \
 //x=45.075 //y=1.22 //x2=45.735 //y2=1.59
cc_4764 ( N_CLK_c_6319_n N_noxref_46_c_11488_n ) capacitor c=0.021347f \
 //x=45.6 //y=1.915 //x2=45.735 //y2=1.59
cc_4765 ( N_CLK_c_6311_n N_noxref_46_M27_noxref_s ) capacitor c=0.00798959f \
 //x=45.075 //y=0.91 //x2=43.745 //y2=0.375
cc_4766 ( N_CLK_c_6318_n N_noxref_46_M27_noxref_s ) capacitor c=0.00212176f \
 //x=45.6 //y=1.45 //x2=43.745 //y2=0.375
cc_4767 ( N_CLK_c_6319_n N_noxref_46_M27_noxref_s ) capacitor c=0.00298115f \
 //x=45.6 //y=1.915 //x2=43.745 //y2=0.375
cc_4768 ( N_CLK_c_6695_p N_noxref_47_c_11507_n ) capacitor c=2.14837e-19 \
 //x=45.445 //y=0.755 //x2=46.305 //y2=0.995
cc_4769 ( N_CLK_c_6316_n N_noxref_47_c_11507_n ) capacitor c=0.00123426f \
 //x=45.6 //y=0.91 //x2=46.305 //y2=0.995
cc_4770 ( N_CLK_c_6317_n N_noxref_47_c_11507_n ) capacitor c=0.0129288f \
 //x=45.6 //y=1.22 //x2=46.305 //y2=0.995
cc_4771 ( N_CLK_c_6318_n N_noxref_47_c_11507_n ) capacitor c=0.00142359f \
 //x=45.6 //y=1.45 //x2=46.305 //y2=0.995
cc_4772 ( N_CLK_c_6311_n N_noxref_47_M28_noxref_d ) capacitor c=0.00223875f \
 //x=45.075 //y=0.91 //x2=45.15 //y2=0.91
cc_4773 ( N_CLK_c_6314_n N_noxref_47_M28_noxref_d ) capacitor c=0.00262485f \
 //x=45.075 //y=1.22 //x2=45.15 //y2=0.91
cc_4774 ( N_CLK_c_6695_p N_noxref_47_M28_noxref_d ) capacitor c=0.00220746f \
 //x=45.445 //y=0.755 //x2=45.15 //y2=0.91
cc_4775 ( N_CLK_c_6702_p N_noxref_47_M28_noxref_d ) capacitor c=0.00194798f \
 //x=45.445 //y=1.375 //x2=45.15 //y2=0.91
cc_4776 ( N_CLK_c_6316_n N_noxref_47_M28_noxref_d ) capacitor c=0.00198465f \
 //x=45.6 //y=0.91 //x2=45.15 //y2=0.91
cc_4777 ( N_CLK_c_6317_n N_noxref_47_M28_noxref_d ) capacitor c=0.00128384f \
 //x=45.6 //y=1.22 //x2=45.15 //y2=0.91
cc_4778 ( N_CLK_c_6316_n N_noxref_47_M29_noxref_s ) capacitor c=7.21316e-19 \
 //x=45.6 //y=0.91 //x2=46.255 //y2=0.375
cc_4779 ( N_CLK_c_6317_n N_noxref_47_M29_noxref_s ) capacitor c=0.00348171f \
 //x=45.6 //y=1.22 //x2=46.255 //y2=0.375
cc_4780 ( N_CLK_c_6421_n N_noxref_54_c_11876_n ) capacitor c=0.0167228f \
 //x=64.315 //y=0.91 //x2=64.975 //y2=0.54
cc_4781 ( N_CLK_c_6426_n N_noxref_54_c_11876_n ) capacitor c=0.00534519f \
 //x=64.84 //y=0.91 //x2=64.975 //y2=0.54
cc_4782 ( N_CLK_c_6044_n N_noxref_54_c_11898_n ) capacitor c=0.0120267f \
 //x=64.75 //y=2.08 //x2=64.975 //y2=1.59
cc_4783 ( N_CLK_c_6424_n N_noxref_54_c_11898_n ) capacitor c=0.0157358f \
 //x=64.315 //y=1.22 //x2=64.975 //y2=1.59
cc_4784 ( N_CLK_c_6429_n N_noxref_54_c_11898_n ) capacitor c=0.021347f \
 //x=64.84 //y=1.915 //x2=64.975 //y2=1.59
cc_4785 ( N_CLK_c_6421_n N_noxref_54_M39_noxref_s ) capacitor c=0.00798959f \
 //x=64.315 //y=0.91 //x2=62.985 //y2=0.375
cc_4786 ( N_CLK_c_6428_n N_noxref_54_M39_noxref_s ) capacitor c=0.00212176f \
 //x=64.84 //y=1.45 //x2=62.985 //y2=0.375
cc_4787 ( N_CLK_c_6429_n N_noxref_54_M39_noxref_s ) capacitor c=0.00298115f \
 //x=64.84 //y=1.915 //x2=62.985 //y2=0.375
cc_4788 ( N_CLK_c_6715_p N_noxref_55_c_11918_n ) capacitor c=2.14837e-19 \
 //x=64.685 //y=0.755 //x2=65.545 //y2=0.995
cc_4789 ( N_CLK_c_6426_n N_noxref_55_c_11918_n ) capacitor c=0.00123426f \
 //x=64.84 //y=0.91 //x2=65.545 //y2=0.995
cc_4790 ( N_CLK_c_6427_n N_noxref_55_c_11918_n ) capacitor c=0.0129288f \
 //x=64.84 //y=1.22 //x2=65.545 //y2=0.995
cc_4791 ( N_CLK_c_6428_n N_noxref_55_c_11918_n ) capacitor c=0.00142359f \
 //x=64.84 //y=1.45 //x2=65.545 //y2=0.995
cc_4792 ( N_CLK_c_6421_n N_noxref_55_M40_noxref_d ) capacitor c=0.00223875f \
 //x=64.315 //y=0.91 //x2=64.39 //y2=0.91
cc_4793 ( N_CLK_c_6424_n N_noxref_55_M40_noxref_d ) capacitor c=0.00262485f \
 //x=64.315 //y=1.22 //x2=64.39 //y2=0.91
cc_4794 ( N_CLK_c_6715_p N_noxref_55_M40_noxref_d ) capacitor c=0.00220746f \
 //x=64.685 //y=0.755 //x2=64.39 //y2=0.91
cc_4795 ( N_CLK_c_6722_p N_noxref_55_M40_noxref_d ) capacitor c=0.00194798f \
 //x=64.685 //y=1.375 //x2=64.39 //y2=0.91
cc_4796 ( N_CLK_c_6426_n N_noxref_55_M40_noxref_d ) capacitor c=0.00198465f \
 //x=64.84 //y=0.91 //x2=64.39 //y2=0.91
cc_4797 ( N_CLK_c_6427_n N_noxref_55_M40_noxref_d ) capacitor c=0.00128384f \
 //x=64.84 //y=1.22 //x2=64.39 //y2=0.91
cc_4798 ( N_CLK_c_6426_n N_noxref_55_M41_noxref_s ) capacitor c=7.21316e-19 \
 //x=64.84 //y=0.91 //x2=65.495 //y2=0.375
cc_4799 ( N_CLK_c_6427_n N_noxref_55_M41_noxref_s ) capacitor c=0.00348171f \
 //x=64.84 //y=1.22 //x2=65.495 //y2=0.375
cc_4800 ( N_CLK_c_6446_n N_noxref_58_c_12078_n ) capacitor c=0.0167228f \
 //x=73.935 //y=0.91 //x2=74.595 //y2=0.54
cc_4801 ( N_CLK_c_6451_n N_noxref_58_c_12078_n ) capacitor c=0.00534519f \
 //x=74.46 //y=0.91 //x2=74.595 //y2=0.54
cc_4802 ( N_CLK_c_6045_n N_noxref_58_c_12100_n ) capacitor c=0.0120267f \
 //x=74.37 //y=2.08 //x2=74.595 //y2=1.59
cc_4803 ( N_CLK_c_6449_n N_noxref_58_c_12100_n ) capacitor c=0.0157358f \
 //x=73.935 //y=1.22 //x2=74.595 //y2=1.59
cc_4804 ( N_CLK_c_6454_n N_noxref_58_c_12100_n ) capacitor c=0.021347f \
 //x=74.46 //y=1.915 //x2=74.595 //y2=1.59
cc_4805 ( N_CLK_c_6446_n N_noxref_58_M45_noxref_s ) capacitor c=0.00798959f \
 //x=73.935 //y=0.91 //x2=72.605 //y2=0.375
cc_4806 ( N_CLK_c_6453_n N_noxref_58_M45_noxref_s ) capacitor c=0.00212176f \
 //x=74.46 //y=1.45 //x2=72.605 //y2=0.375
cc_4807 ( N_CLK_c_6454_n N_noxref_58_M45_noxref_s ) capacitor c=0.00298115f \
 //x=74.46 //y=1.915 //x2=72.605 //y2=0.375
cc_4808 ( N_CLK_c_6735_p N_noxref_59_c_12120_n ) capacitor c=2.14837e-19 \
 //x=74.305 //y=0.755 //x2=75.165 //y2=0.995
cc_4809 ( N_CLK_c_6451_n N_noxref_59_c_12120_n ) capacitor c=0.00123426f \
 //x=74.46 //y=0.91 //x2=75.165 //y2=0.995
cc_4810 ( N_CLK_c_6452_n N_noxref_59_c_12120_n ) capacitor c=0.0129288f \
 //x=74.46 //y=1.22 //x2=75.165 //y2=0.995
cc_4811 ( N_CLK_c_6453_n N_noxref_59_c_12120_n ) capacitor c=0.00142359f \
 //x=74.46 //y=1.45 //x2=75.165 //y2=0.995
cc_4812 ( N_CLK_c_6446_n N_noxref_59_M46_noxref_d ) capacitor c=0.00223875f \
 //x=73.935 //y=0.91 //x2=74.01 //y2=0.91
cc_4813 ( N_CLK_c_6449_n N_noxref_59_M46_noxref_d ) capacitor c=0.00262485f \
 //x=73.935 //y=1.22 //x2=74.01 //y2=0.91
cc_4814 ( N_CLK_c_6735_p N_noxref_59_M46_noxref_d ) capacitor c=0.00220746f \
 //x=74.305 //y=0.755 //x2=74.01 //y2=0.91
cc_4815 ( N_CLK_c_6742_p N_noxref_59_M46_noxref_d ) capacitor c=0.00194798f \
 //x=74.305 //y=1.375 //x2=74.01 //y2=0.91
cc_4816 ( N_CLK_c_6451_n N_noxref_59_M46_noxref_d ) capacitor c=0.00198465f \
 //x=74.46 //y=0.91 //x2=74.01 //y2=0.91
cc_4817 ( N_CLK_c_6452_n N_noxref_59_M46_noxref_d ) capacitor c=0.00128384f \
 //x=74.46 //y=1.22 //x2=74.01 //y2=0.91
cc_4818 ( N_CLK_c_6451_n N_noxref_59_M47_noxref_s ) capacitor c=7.21316e-19 \
 //x=74.46 //y=0.91 //x2=75.115 //y2=0.375
cc_4819 ( N_CLK_c_6452_n N_noxref_59_M47_noxref_s ) capacitor c=0.00348171f \
 //x=74.46 //y=1.22 //x2=75.115 //y2=0.375
cc_4820 ( N_noxref_18_c_6814_n N_RN_c_7071_n ) capacitor c=0.00374603f \
 //x=66.485 //y=3.33 //x2=75.365 //y2=2.22
cc_4821 ( N_noxref_18_c_6820_n N_RN_c_7071_n ) capacitor c=7.32243e-19 \
 //x=61.165 //y=3.33 //x2=75.365 //y2=2.22
cc_4822 ( N_noxref_18_c_6821_n N_RN_c_7071_n ) capacitor c=0.0316113f \
 //x=77.955 //y=3.33 //x2=75.365 //y2=2.22
cc_4823 ( N_noxref_18_c_6747_n N_RN_c_7071_n ) capacitor c=0.0209607f \
 //x=61.05 //y=2.08 //x2=75.365 //y2=2.22
cc_4824 ( N_noxref_18_c_6881_p N_RN_c_7071_n ) capacitor c=0.016327f //x=66.2 \
 //y=1.665 //x2=75.365 //y2=2.22
cc_4825 ( N_noxref_18_c_6776_n N_RN_c_7071_n ) capacitor c=0.0197307f //x=66.6 \
 //y=3.33 //x2=75.365 //y2=2.22
cc_4826 ( N_noxref_18_c_6843_n N_RN_c_7071_n ) capacitor c=3.13485e-19 \
 //x=61.415 //y=1.415 //x2=75.365 //y2=2.22
cc_4827 ( N_noxref_18_c_6848_n N_RN_c_7071_n ) capacitor c=0.00584491f \
 //x=61.05 //y=2.08 //x2=75.365 //y2=2.22
cc_4828 ( N_noxref_18_c_6747_n N_RN_c_7082_n ) capacitor c=0.00165648f \
 //x=61.05 //y=2.08 //x2=60.055 //y2=2.22
cc_4829 ( N_noxref_18_c_6848_n N_RN_c_7082_n ) capacitor c=2.3323e-19 \
 //x=61.05 //y=2.08 //x2=60.055 //y2=2.22
cc_4830 ( N_noxref_18_c_6821_n N_RN_c_7083_n ) capacitor c=0.014255f \
 //x=77.955 //y=3.33 //x2=79.065 //y2=2.22
cc_4831 ( N_noxref_18_c_6749_n N_RN_c_7083_n ) capacitor c=0.0226137f \
 //x=78.07 //y=2.08 //x2=79.065 //y2=2.22
cc_4832 ( N_noxref_18_c_6754_n N_RN_c_7083_n ) capacitor c=0.0121989f \
 //x=77.77 //y=1.915 //x2=79.065 //y2=2.22
cc_4833 ( N_noxref_18_c_6821_n N_RN_c_7087_n ) capacitor c=4.86139e-19 \
 //x=77.955 //y=3.33 //x2=75.595 //y2=2.22
cc_4834 ( N_noxref_18_c_6820_n N_RN_c_7094_n ) capacitor c=0.00373989f \
 //x=61.165 //y=3.33 //x2=59.94 //y2=2.08
cc_4835 ( N_noxref_18_c_6747_n N_RN_c_7094_n ) capacitor c=0.0446367f \
 //x=61.05 //y=2.08 //x2=59.94 //y2=2.08
cc_4836 ( N_noxref_18_c_6848_n N_RN_c_7094_n ) capacitor c=0.0019893f \
 //x=61.05 //y=2.08 //x2=59.94 //y2=2.08
cc_4837 ( N_noxref_18_c_6812_n N_RN_c_7094_n ) capacitor c=0.00197875f \
 //x=61.05 //y=4.7 //x2=59.94 //y2=2.08
cc_4838 ( N_noxref_18_c_6821_n N_RN_c_7095_n ) capacitor c=0.0180187f \
 //x=77.955 //y=3.33 //x2=75.48 //y2=2.08
cc_4839 ( N_noxref_18_c_6749_n N_RN_c_7095_n ) capacitor c=6.89573e-19 \
 //x=78.07 //y=2.08 //x2=75.48 //y2=2.08
cc_4840 ( N_noxref_18_c_6821_n N_RN_c_7096_n ) capacitor c=0.00526349f \
 //x=77.955 //y=3.33 //x2=79.18 //y2=2.08
cc_4841 ( N_noxref_18_c_6749_n N_RN_c_7096_n ) capacitor c=0.0444055f \
 //x=78.07 //y=2.08 //x2=79.18 //y2=2.08
cc_4842 ( N_noxref_18_c_6754_n N_RN_c_7096_n ) capacitor c=0.00208635f \
 //x=77.77 //y=1.915 //x2=79.18 //y2=2.08
cc_4843 ( N_noxref_18_c_6900_p N_RN_c_7096_n ) capacitor c=0.00147352f \
 //x=78.635 //y=4.79 //x2=79.18 //y2=2.08
cc_4844 ( N_noxref_18_c_6788_n N_RN_c_7096_n ) capacitor c=0.00142741f \
 //x=78.345 //y=4.79 //x2=79.18 //y2=2.08
cc_4845 ( N_noxref_18_M136_noxref_g N_RN_M134_noxref_g ) capacitor \
 c=0.0100903f //x=60.79 //y=6.02 //x2=59.91 //y2=6.02
cc_4846 ( N_noxref_18_M136_noxref_g N_RN_M135_noxref_g ) capacitor \
 c=0.0600064f //x=60.79 //y=6.02 //x2=60.35 //y2=6.02
cc_4847 ( N_noxref_18_M137_noxref_g N_RN_M135_noxref_g ) capacitor \
 c=0.0100903f //x=61.23 //y=6.02 //x2=60.35 //y2=6.02
cc_4848 ( N_noxref_18_M156_noxref_g N_RN_M158_noxref_g ) capacitor \
 c=0.0105869f //x=78.27 //y=6.02 //x2=79.15 //y2=6.02
cc_4849 ( N_noxref_18_M157_noxref_g N_RN_M158_noxref_g ) capacitor c=0.10632f \
 //x=78.71 //y=6.02 //x2=79.15 //y2=6.02
cc_4850 ( N_noxref_18_M157_noxref_g N_RN_M159_noxref_g ) capacitor \
 c=0.0101598f //x=78.71 //y=6.02 //x2=79.59 //y2=6.02
cc_4851 ( N_noxref_18_c_6839_n N_RN_c_7554_n ) capacitor c=0.00456962f \
 //x=61.04 //y=0.915 //x2=60.03 //y2=0.91
cc_4852 ( N_noxref_18_c_6840_n N_RN_c_7555_n ) capacitor c=0.00438372f \
 //x=61.04 //y=1.26 //x2=60.03 //y2=1.22
cc_4853 ( N_noxref_18_c_6841_n N_RN_c_7556_n ) capacitor c=0.00438372f \
 //x=61.04 //y=1.57 //x2=60.03 //y2=1.45
cc_4854 ( N_noxref_18_c_6747_n N_RN_c_7557_n ) capacitor c=0.00205895f \
 //x=61.05 //y=2.08 //x2=60.03 //y2=1.915
cc_4855 ( N_noxref_18_c_6848_n N_RN_c_7557_n ) capacitor c=0.00828003f \
 //x=61.05 //y=2.08 //x2=60.03 //y2=1.915
cc_4856 ( N_noxref_18_c_6849_n N_RN_c_7557_n ) capacitor c=0.00438372f \
 //x=61.05 //y=1.915 //x2=60.03 //y2=1.915
cc_4857 ( N_noxref_18_c_6812_n N_RN_c_7258_n ) capacitor c=0.0609323f \
 //x=61.05 //y=4.7 //x2=60.275 //y2=4.79
cc_4858 ( N_noxref_18_c_6750_n N_RN_c_7714_n ) capacitor c=5.72482e-19 \
 //x=77.77 //y=0.875 //x2=78.745 //y2=0.91
cc_4859 ( N_noxref_18_c_6752_n N_RN_c_7714_n ) capacitor c=0.00149976f \
 //x=77.77 //y=1.22 //x2=78.745 //y2=0.91
cc_4860 ( N_noxref_18_c_6757_n N_RN_c_7714_n ) capacitor c=0.0160123f //x=78.3 \
 //y=0.875 //x2=78.745 //y2=0.91
cc_4861 ( N_noxref_18_c_6753_n N_RN_c_7717_n ) capacitor c=0.00111227f \
 //x=77.77 //y=1.53 //x2=78.745 //y2=1.22
cc_4862 ( N_noxref_18_c_6759_n N_RN_c_7717_n ) capacitor c=0.0124075f //x=78.3 \
 //y=1.22 //x2=78.745 //y2=1.22
cc_4863 ( N_noxref_18_c_6757_n N_RN_c_7719_n ) capacitor c=0.00103227f \
 //x=78.3 //y=0.875 //x2=79.27 //y2=0.91
cc_4864 ( N_noxref_18_c_6759_n N_RN_c_7720_n ) capacitor c=0.0010154f //x=78.3 \
 //y=1.22 //x2=79.27 //y2=1.22
cc_4865 ( N_noxref_18_c_6759_n N_RN_c_7721_n ) capacitor c=9.23422e-19 \
 //x=78.3 //y=1.22 //x2=79.27 //y2=1.45
cc_4866 ( N_noxref_18_c_6749_n N_RN_c_7722_n ) capacitor c=0.00203769f \
 //x=78.07 //y=2.08 //x2=79.27 //y2=1.915
cc_4867 ( N_noxref_18_c_6754_n N_RN_c_7722_n ) capacitor c=0.00834532f \
 //x=77.77 //y=1.915 //x2=79.27 //y2=1.915
cc_4868 ( N_noxref_18_c_6747_n N_RN_c_7264_n ) capacitor c=0.00142741f \
 //x=61.05 //y=2.08 //x2=59.94 //y2=4.7
cc_4869 ( N_noxref_18_c_6812_n N_RN_c_7264_n ) capacitor c=0.00487508f \
 //x=61.05 //y=4.7 //x2=59.94 //y2=4.7
cc_4870 ( N_noxref_18_c_6749_n N_RN_c_7268_n ) capacitor c=0.00183762f \
 //x=78.07 //y=2.08 //x2=79.18 //y2=4.7
cc_4871 ( N_noxref_18_c_6900_p N_RN_c_7268_n ) capacitor c=0.0168581f \
 //x=78.635 //y=4.79 //x2=79.18 //y2=4.7
cc_4872 ( N_noxref_18_c_6788_n N_RN_c_7268_n ) capacitor c=0.00484466f \
 //x=78.345 //y=4.79 //x2=79.18 //y2=4.7
cc_4873 ( N_noxref_18_c_6814_n N_SN_c_8138_n ) capacitor c=0.466581f \
 //x=66.485 //y=3.33 //x2=69.445 //y2=2.96
cc_4874 ( N_noxref_18_c_6820_n N_SN_c_8138_n ) capacitor c=0.0291389f \
 //x=61.165 //y=3.33 //x2=69.445 //y2=2.96
cc_4875 ( N_noxref_18_c_6821_n N_SN_c_8138_n ) capacitor c=0.241804f \
 //x=77.955 //y=3.33 //x2=69.445 //y2=2.96
cc_4876 ( N_noxref_18_c_6823_n N_SN_c_8138_n ) capacitor c=0.0266688f \
 //x=66.715 //y=3.33 //x2=69.445 //y2=2.96
cc_4877 ( N_noxref_18_c_6747_n N_SN_c_8138_n ) capacitor c=0.0221202f \
 //x=61.05 //y=2.08 //x2=69.445 //y2=2.96
cc_4878 ( N_noxref_18_c_6776_n N_SN_c_8138_n ) capacitor c=0.020574f //x=66.6 \
 //y=3.33 //x2=69.445 //y2=2.96
cc_4879 ( N_noxref_18_c_6821_n N_SN_c_8141_n ) capacitor c=0.756732f \
 //x=77.955 //y=3.33 //x2=83.875 //y2=2.96
cc_4880 ( N_noxref_18_c_6749_n N_SN_c_8141_n ) capacitor c=0.0238838f \
 //x=78.07 //y=2.08 //x2=83.875 //y2=2.96
cc_4881 ( N_noxref_18_c_6821_n N_SN_c_8468_n ) capacitor c=0.0265806f \
 //x=77.955 //y=3.33 //x2=69.675 //y2=2.96
cc_4882 ( N_noxref_18_c_6821_n N_SN_c_8149_n ) capacitor c=0.0208912f \
 //x=77.955 //y=3.33 //x2=69.56 //y2=2.08
cc_4883 ( N_noxref_18_c_6776_n N_SN_c_8149_n ) capacitor c=3.55725e-19 \
 //x=66.6 //y=3.33 //x2=69.56 //y2=2.08
cc_4884 ( N_noxref_18_c_6814_n N_noxref_21_c_8898_n ) capacitor c=0.0446157f \
 //x=66.485 //y=3.33 //x2=70.555 //y2=3.7
cc_4885 ( N_noxref_18_c_6821_n N_noxref_21_c_8898_n ) capacitor c=0.340407f \
 //x=77.955 //y=3.33 //x2=70.555 //y2=3.7
cc_4886 ( N_noxref_18_c_6823_n N_noxref_21_c_8898_n ) capacitor c=0.0268386f \
 //x=66.715 //y=3.33 //x2=70.555 //y2=3.7
cc_4887 ( N_noxref_18_c_6776_n N_noxref_21_c_8898_n ) capacitor c=0.0205782f \
 //x=66.6 //y=3.33 //x2=70.555 //y2=3.7
cc_4888 ( N_noxref_18_c_6814_n N_noxref_21_c_8935_n ) capacitor c=0.029444f \
 //x=66.485 //y=3.33 //x2=65.975 //y2=3.7
cc_4889 ( N_noxref_18_c_6776_n N_noxref_21_c_8935_n ) capacitor c=0.00155359f \
 //x=66.6 //y=3.33 //x2=65.975 //y2=3.7
cc_4890 ( N_noxref_18_c_6821_n N_noxref_21_c_8878_n ) capacitor c=0.468734f \
 //x=77.955 //y=3.33 //x2=76.105 //y2=3.7
cc_4891 ( N_noxref_18_c_6821_n N_noxref_21_c_8905_n ) capacitor c=0.026734f \
 //x=77.955 //y=3.33 //x2=70.785 //y2=3.7
cc_4892 ( N_noxref_18_c_6821_n N_noxref_21_c_8880_n ) capacitor c=0.176086f \
 //x=77.955 //y=3.33 //x2=84.985 //y2=3.7
cc_4893 ( N_noxref_18_c_6749_n N_noxref_21_c_8880_n ) capacitor c=0.0215974f \
 //x=78.07 //y=2.08 //x2=84.985 //y2=3.7
cc_4894 ( N_noxref_18_c_6821_n N_noxref_21_c_8881_n ) capacitor c=0.0268461f \
 //x=77.955 //y=3.33 //x2=76.335 //y2=3.7
cc_4895 ( N_noxref_18_c_6749_n N_noxref_21_c_8881_n ) capacitor c=7.01366e-19 \
 //x=78.07 //y=2.08 //x2=76.335 //y2=3.7
cc_4896 ( N_noxref_18_c_6814_n N_noxref_21_c_8828_n ) capacitor c=0.0198536f \
 //x=66.485 //y=3.33 //x2=65.86 //y2=2.08
cc_4897 ( N_noxref_18_c_6823_n N_noxref_21_c_8828_n ) capacitor c=0.00179385f \
 //x=66.715 //y=3.33 //x2=65.86 //y2=2.08
cc_4898 ( N_noxref_18_c_6776_n N_noxref_21_c_8828_n ) capacitor c=0.0730663f \
 //x=66.6 //y=3.33 //x2=65.86 //y2=2.08
cc_4899 ( N_noxref_18_c_6956_p N_noxref_21_c_8828_n ) capacitor c=0.0126839f \
 //x=65.82 //y=5.155 //x2=65.86 //y2=2.08
cc_4900 ( N_noxref_18_c_6821_n N_noxref_21_c_8829_n ) capacitor c=0.0198536f \
 //x=77.955 //y=3.33 //x2=70.67 //y2=2.08
cc_4901 ( N_noxref_18_c_6821_n N_noxref_21_c_8849_n ) capacitor c=0.0212788f \
 //x=77.955 //y=3.33 //x2=76.22 //y2=3.7
cc_4902 ( N_noxref_18_c_6749_n N_noxref_21_c_8849_n ) capacitor c=0.0106001f \
 //x=78.07 //y=2.08 //x2=76.22 //y2=3.7
cc_4903 ( N_noxref_18_c_6768_n N_noxref_21_M142_noxref_g ) capacitor \
 c=0.0162556f //x=65.735 //y=5.155 //x2=65.6 //y2=6.02
cc_4904 ( N_noxref_18_M142_noxref_d N_noxref_21_M142_noxref_g ) capacitor \
 c=0.0180032f //x=65.675 //y=5.02 //x2=65.6 //y2=6.02
cc_4905 ( N_noxref_18_c_6772_n N_noxref_21_M143_noxref_g ) capacitor \
 c=0.0183937f //x=66.515 //y=5.155 //x2=66.04 //y2=6.02
cc_4906 ( N_noxref_18_M142_noxref_d N_noxref_21_M143_noxref_g ) capacitor \
 c=0.0194246f //x=65.675 //y=5.02 //x2=66.04 //y2=6.02
cc_4907 ( N_noxref_18_M41_noxref_d N_noxref_21_c_8955_n ) capacitor \
 c=0.00217566f //x=65.925 //y=0.915 //x2=65.85 //y2=0.915
cc_4908 ( N_noxref_18_M41_noxref_d N_noxref_21_c_8956_n ) capacitor \
 c=0.0034598f //x=65.925 //y=0.915 //x2=65.85 //y2=1.26
cc_4909 ( N_noxref_18_M41_noxref_d N_noxref_21_c_8957_n ) capacitor \
 c=0.00546784f //x=65.925 //y=0.915 //x2=65.85 //y2=1.57
cc_4910 ( N_noxref_18_M41_noxref_d N_noxref_21_c_8994_n ) capacitor \
 c=0.00241102f //x=65.925 //y=0.915 //x2=66.225 //y2=0.76
cc_4911 ( N_noxref_18_c_6748_n N_noxref_21_c_8995_n ) capacitor c=0.00371277f \
 //x=66.515 //y=1.665 //x2=66.225 //y2=1.415
cc_4912 ( N_noxref_18_M41_noxref_d N_noxref_21_c_8995_n ) capacitor \
 c=0.0138621f //x=65.925 //y=0.915 //x2=66.225 //y2=1.415
cc_4913 ( N_noxref_18_M41_noxref_d N_noxref_21_c_8997_n ) capacitor \
 c=0.00219619f //x=65.925 //y=0.915 //x2=66.38 //y2=0.915
cc_4914 ( N_noxref_18_c_6748_n N_noxref_21_c_8998_n ) capacitor c=0.00457401f \
 //x=66.515 //y=1.665 //x2=66.38 //y2=1.26
cc_4915 ( N_noxref_18_M41_noxref_d N_noxref_21_c_8998_n ) capacitor \
 c=0.00603828f //x=65.925 //y=0.915 //x2=66.38 //y2=1.26
cc_4916 ( N_noxref_18_c_6776_n N_noxref_21_c_8958_n ) capacitor c=0.00731987f \
 //x=66.6 //y=3.33 //x2=65.86 //y2=2.08
cc_4917 ( N_noxref_18_c_6776_n N_noxref_21_c_8960_n ) capacitor c=0.00283672f \
 //x=66.6 //y=3.33 //x2=65.86 //y2=1.915
cc_4918 ( N_noxref_18_M41_noxref_d N_noxref_21_c_8960_n ) capacitor \
 c=0.00661782f //x=65.925 //y=0.915 //x2=65.86 //y2=1.915
cc_4919 ( N_noxref_18_c_6772_n N_noxref_21_c_8895_n ) capacitor c=0.00201851f \
 //x=66.515 //y=5.155 //x2=65.86 //y2=4.7
cc_4920 ( N_noxref_18_c_6776_n N_noxref_21_c_8895_n ) capacitor c=0.0114782f \
 //x=66.6 //y=3.33 //x2=65.86 //y2=4.7
cc_4921 ( N_noxref_18_c_6956_p N_noxref_21_c_8895_n ) capacitor c=0.00470675f \
 //x=65.82 //y=5.155 //x2=65.86 //y2=4.7
cc_4922 ( N_noxref_18_c_6749_n N_noxref_22_c_9175_n ) capacitor c=0.00127817f \
 //x=78.07 //y=2.08 //x2=80.29 //y2=2.08
cc_4923 ( N_noxref_18_M157_noxref_g N_noxref_24_c_9478_n ) capacitor \
 c=0.0168349f //x=78.71 //y=6.02 //x2=79.285 //y2=5.155
cc_4924 ( N_noxref_18_M156_noxref_g N_noxref_24_c_9482_n ) capacitor \
 c=0.0213876f //x=78.27 //y=6.02 //x2=78.575 //y2=5.155
cc_4925 ( N_noxref_18_c_6900_p N_noxref_24_c_9482_n ) capacitor c=0.00428486f \
 //x=78.635 //y=4.79 //x2=78.575 //y2=5.155
cc_4926 ( N_noxref_18_M157_noxref_g N_noxref_24_M156_noxref_d ) capacitor \
 c=0.0180032f //x=78.71 //y=6.02 //x2=78.345 //y2=5.02
cc_4927 ( N_noxref_18_c_6820_n N_noxref_26_c_10050_n ) capacitor c=0.0018493f \
 //x=61.165 //y=3.33 //x2=56.895 //y2=3.33
cc_4928 ( N_noxref_18_c_6814_n N_noxref_26_c_9933_n ) capacitor c=0.35768f \
 //x=66.485 //y=3.33 //x2=65.035 //y2=3.7
cc_4929 ( N_noxref_18_c_6820_n N_noxref_26_c_9933_n ) capacitor c=0.0293356f \
 //x=61.165 //y=3.33 //x2=65.035 //y2=3.7
cc_4930 ( N_noxref_18_c_6747_n N_noxref_26_c_9933_n ) capacitor c=0.0221397f \
 //x=61.05 //y=2.08 //x2=65.035 //y2=3.7
cc_4931 ( N_noxref_18_c_6814_n N_noxref_26_c_9912_n ) capacitor c=0.0274571f \
 //x=66.485 //y=3.33 //x2=88.315 //y2=4.07
cc_4932 ( N_noxref_18_c_6821_n N_noxref_26_c_9912_n ) capacitor c=0.0809428f \
 //x=77.955 //y=3.33 //x2=88.315 //y2=4.07
cc_4933 ( N_noxref_18_c_6823_n N_noxref_26_c_9912_n ) capacitor c=4.80262e-19 \
 //x=66.715 //y=3.33 //x2=88.315 //y2=4.07
cc_4934 ( N_noxref_18_c_6776_n N_noxref_26_c_9912_n ) capacitor c=0.0181789f \
 //x=66.6 //y=3.33 //x2=88.315 //y2=4.07
cc_4935 ( N_noxref_18_c_6749_n N_noxref_26_c_9912_n ) capacitor c=0.0194977f \
 //x=78.07 //y=2.08 //x2=88.315 //y2=4.07
cc_4936 ( N_noxref_18_c_6747_n N_noxref_53_c_11822_n ) capacitor c=0.00204385f \
 //x=61.05 //y=2.08 //x2=61.705 //y2=0.54
cc_4937 ( N_noxref_18_c_6839_n N_noxref_53_c_11822_n ) capacitor c=0.0194423f \
 //x=61.04 //y=0.915 //x2=61.705 //y2=0.54
cc_4938 ( N_noxref_18_c_6845_n N_noxref_53_c_11822_n ) capacitor c=0.00656458f \
 //x=61.57 //y=0.915 //x2=61.705 //y2=0.54
cc_4939 ( N_noxref_18_c_6848_n N_noxref_53_c_11822_n ) capacitor c=2.20712e-19 \
 //x=61.05 //y=2.08 //x2=61.705 //y2=0.54
cc_4940 ( N_noxref_18_c_6840_n N_noxref_53_c_11832_n ) capacitor c=0.00538829f \
 //x=61.04 //y=1.26 //x2=60.82 //y2=0.995
cc_4941 ( N_noxref_18_c_6839_n N_noxref_53_M38_noxref_s ) capacitor \
 c=0.00538829f //x=61.04 //y=0.915 //x2=60.685 //y2=0.375
cc_4942 ( N_noxref_18_c_6841_n N_noxref_53_M38_noxref_s ) capacitor \
 c=0.00538829f //x=61.04 //y=1.57 //x2=60.685 //y2=0.375
cc_4943 ( N_noxref_18_c_6845_n N_noxref_53_M38_noxref_s ) capacitor \
 c=0.0143002f //x=61.57 //y=0.915 //x2=60.685 //y2=0.375
cc_4944 ( N_noxref_18_c_6846_n N_noxref_53_M38_noxref_s ) capacitor \
 c=0.00290153f //x=61.57 //y=1.26 //x2=60.685 //y2=0.375
cc_4945 ( N_noxref_18_M41_noxref_d N_noxref_54_M39_noxref_s ) capacitor \
 c=0.00309936f //x=65.925 //y=0.915 //x2=62.985 //y2=0.375
cc_4946 ( N_noxref_18_c_6748_n N_noxref_55_c_11923_n ) capacitor c=0.00457167f \
 //x=66.515 //y=1.665 //x2=66.515 //y2=0.54
cc_4947 ( N_noxref_18_M41_noxref_d N_noxref_55_c_11923_n ) capacitor \
 c=0.0115903f //x=65.925 //y=0.915 //x2=66.515 //y2=0.54
cc_4948 ( N_noxref_18_c_6881_p N_noxref_55_c_11945_n ) capacitor c=0.0200405f \
 //x=66.2 //y=1.665 //x2=65.63 //y2=0.995
cc_4949 ( N_noxref_18_M41_noxref_d N_noxref_55_M40_noxref_d ) capacitor \
 c=5.27807e-19 //x=65.925 //y=0.915 //x2=64.39 //y2=0.91
cc_4950 ( N_noxref_18_c_6748_n N_noxref_55_M41_noxref_s ) capacitor \
 c=0.0196084f //x=66.515 //y=1.665 //x2=65.495 //y2=0.375
cc_4951 ( N_noxref_18_M41_noxref_d N_noxref_55_M41_noxref_s ) capacitor \
 c=0.0426368f //x=65.925 //y=0.915 //x2=65.495 //y2=0.375
cc_4952 ( N_noxref_18_c_6748_n N_noxref_56_c_11985_n ) capacitor c=3.84569e-19 \
 //x=66.515 //y=1.665 //x2=67.93 //y2=1.505
cc_4953 ( N_noxref_18_M41_noxref_d N_noxref_56_M42_noxref_s ) capacitor \
 c=2.55333e-19 //x=65.925 //y=0.915 //x2=67.795 //y2=0.375
cc_4954 ( N_noxref_18_c_6754_n N_noxref_60_c_12188_n ) capacitor c=0.0034165f \
 //x=77.77 //y=1.915 //x2=77.55 //y2=1.505
cc_4955 ( N_noxref_18_c_6749_n N_noxref_60_c_12173_n ) capacitor c=0.0115578f \
 //x=78.07 //y=2.08 //x2=78.435 //y2=1.59
cc_4956 ( N_noxref_18_c_6753_n N_noxref_60_c_12173_n ) capacitor c=0.00697148f \
 //x=77.77 //y=1.53 //x2=78.435 //y2=1.59
cc_4957 ( N_noxref_18_c_6754_n N_noxref_60_c_12173_n ) capacitor c=0.0204849f \
 //x=77.77 //y=1.915 //x2=78.435 //y2=1.59
cc_4958 ( N_noxref_18_c_6756_n N_noxref_60_c_12173_n ) capacitor c=0.00610316f \
 //x=78.145 //y=1.375 //x2=78.435 //y2=1.59
cc_4959 ( N_noxref_18_c_6759_n N_noxref_60_c_12173_n ) capacitor c=0.00698822f \
 //x=78.3 //y=1.22 //x2=78.435 //y2=1.59
cc_4960 ( N_noxref_18_c_6750_n N_noxref_60_M48_noxref_s ) capacitor \
 c=0.0327271f //x=77.77 //y=0.875 //x2=77.415 //y2=0.375
cc_4961 ( N_noxref_18_c_6753_n N_noxref_60_M48_noxref_s ) capacitor \
 c=7.99997e-19 //x=77.77 //y=1.53 //x2=77.415 //y2=0.375
cc_4962 ( N_noxref_18_c_6754_n N_noxref_60_M48_noxref_s ) capacitor \
 c=0.00122123f //x=77.77 //y=1.915 //x2=77.415 //y2=0.375
cc_4963 ( N_noxref_18_c_6757_n N_noxref_60_M48_noxref_s ) capacitor \
 c=0.0121427f //x=78.3 //y=0.875 //x2=77.415 //y2=0.375
cc_4964 ( N_RN_c_7021_n N_SN_c_8129_n ) capacitor c=0.16065f //x=17.645 \
 //y=2.22 //x2=26.155 //y2=2.96
cc_4965 ( N_RN_c_7033_n N_SN_c_8129_n ) capacitor c=0.147213f //x=21.345 \
 //y=2.22 //x2=26.155 //y2=2.96
cc_4966 ( N_RN_c_7037_n N_SN_c_8129_n ) capacitor c=0.0120222f //x=17.875 \
 //y=2.22 //x2=26.155 //y2=2.96
cc_4967 ( N_RN_c_7038_n N_SN_c_8129_n ) capacitor c=0.114788f //x=30.965 \
 //y=2.22 //x2=26.155 //y2=2.96
cc_4968 ( N_RN_c_7045_n N_SN_c_8129_n ) capacitor c=0.0120222f //x=21.575 \
 //y=2.22 //x2=26.155 //y2=2.96
cc_4969 ( N_RN_c_7089_n N_SN_c_8129_n ) capacitor c=0.0206071f //x=17.76 \
 //y=2.08 //x2=26.155 //y2=2.96
cc_4970 ( N_RN_c_7090_n N_SN_c_8129_n ) capacitor c=0.0239871f //x=21.46 \
 //y=2.08 //x2=26.155 //y2=2.96
cc_4971 ( N_RN_c_7021_n N_SN_c_8183_n ) capacitor c=0.0132253f //x=17.645 \
 //y=2.22 //x2=11.955 //y2=2.96
cc_4972 ( N_RN_c_7038_n N_SN_c_8132_n ) capacitor c=0.193077f //x=30.965 \
 //y=2.22 //x2=40.585 //y2=2.96
cc_4973 ( N_RN_c_7046_n N_SN_c_8132_n ) capacitor c=0.151423f //x=46.505 \
 //y=2.22 //x2=40.585 //y2=2.96
cc_4974 ( N_RN_c_7057_n N_SN_c_8132_n ) capacitor c=0.0120222f //x=31.195 \
 //y=2.22 //x2=40.585 //y2=2.96
cc_4975 ( N_RN_c_7091_n N_SN_c_8132_n ) capacitor c=0.0255045f //x=31.08 \
 //y=2.08 //x2=40.585 //y2=2.96
cc_4976 ( N_RN_c_7038_n N_SN_c_8226_n ) capacitor c=0.0119704f //x=30.965 \
 //y=2.22 //x2=26.385 //y2=2.96
cc_4977 ( N_RN_c_7046_n N_SN_c_8135_n ) capacitor c=0.16065f //x=46.505 \
 //y=2.22 //x2=55.015 //y2=2.96
cc_4978 ( N_RN_c_7058_n N_SN_c_8135_n ) capacitor c=0.147213f //x=50.205 \
 //y=2.22 //x2=55.015 //y2=2.96
cc_4979 ( N_RN_c_7062_n N_SN_c_8135_n ) capacitor c=0.0120222f //x=46.735 \
 //y=2.22 //x2=55.015 //y2=2.96
cc_4980 ( N_RN_c_7063_n N_SN_c_8135_n ) capacitor c=0.062775f //x=59.825 \
 //y=2.22 //x2=55.015 //y2=2.96
cc_4981 ( N_RN_c_7070_n N_SN_c_8135_n ) capacitor c=0.0120222f //x=50.435 \
 //y=2.22 //x2=55.015 //y2=2.96
cc_4982 ( N_RN_c_7092_n N_SN_c_8135_n ) capacitor c=0.0206071f //x=46.62 \
 //y=2.08 //x2=55.015 //y2=2.96
cc_4983 ( N_RN_c_7093_n N_SN_c_8135_n ) capacitor c=0.0239871f //x=50.32 \
 //y=2.08 //x2=55.015 //y2=2.96
cc_4984 ( N_RN_c_7046_n N_SN_c_8340_n ) capacitor c=0.0119704f //x=46.505 \
 //y=2.22 //x2=40.815 //y2=2.96
cc_4985 ( N_RN_c_7063_n N_SN_c_8138_n ) capacitor c=0.131652f //x=59.825 \
 //y=2.22 //x2=69.445 //y2=2.96
cc_4986 ( N_RN_c_7071_n N_SN_c_8138_n ) capacitor c=0.151423f //x=75.365 \
 //y=2.22 //x2=69.445 //y2=2.96
cc_4987 ( N_RN_c_7082_n N_SN_c_8138_n ) capacitor c=0.0120222f //x=60.055 \
 //y=2.22 //x2=69.445 //y2=2.96
cc_4988 ( N_RN_c_7094_n N_SN_c_8138_n ) capacitor c=0.0239871f //x=59.94 \
 //y=2.08 //x2=69.445 //y2=2.96
cc_4989 ( N_RN_c_7063_n N_SN_c_8399_n ) capacitor c=6.57895e-19 //x=59.825 \
 //y=2.22 //x2=55.245 //y2=2.96
cc_4990 ( N_RN_c_7071_n N_SN_c_8141_n ) capacitor c=0.16065f //x=75.365 \
 //y=2.22 //x2=83.875 //y2=2.96
cc_4991 ( N_RN_c_7083_n N_SN_c_8141_n ) capacitor c=0.16049f //x=79.065 \
 //y=2.22 //x2=83.875 //y2=2.96
cc_4992 ( N_RN_c_7087_n N_SN_c_8141_n ) capacitor c=0.0120222f //x=75.595 \
 //y=2.22 //x2=83.875 //y2=2.96
cc_4993 ( N_RN_c_7095_n N_SN_c_8141_n ) capacitor c=0.0206071f //x=75.48 \
 //y=2.08 //x2=83.875 //y2=2.96
cc_4994 ( N_RN_c_7096_n N_SN_c_8141_n ) capacitor c=0.0239871f //x=79.18 \
 //y=2.08 //x2=83.875 //y2=2.96
cc_4995 ( N_RN_c_7722_n N_SN_c_8141_n ) capacitor c=4.10467e-19 //x=79.27 \
 //y=1.915 //x2=83.875 //y2=2.96
cc_4996 ( N_RN_c_7071_n N_SN_c_8468_n ) capacitor c=0.0119704f //x=75.365 \
 //y=2.22 //x2=69.675 //y2=2.96
cc_4997 ( N_RN_c_7021_n N_SN_c_8145_n ) capacitor c=0.0220464f //x=17.645 \
 //y=2.22 //x2=11.84 //y2=2.08
cc_4998 ( N_RN_c_7038_n N_SN_c_8146_n ) capacitor c=0.0220464f //x=30.965 \
 //y=2.22 //x2=26.27 //y2=2.08
cc_4999 ( N_RN_c_7046_n N_SN_c_8147_n ) capacitor c=0.0220464f //x=46.505 \
 //y=2.22 //x2=40.7 //y2=2.08
cc_5000 ( N_RN_c_7063_n N_SN_c_8148_n ) capacitor c=0.0193884f //x=59.825 \
 //y=2.22 //x2=55.13 //y2=2.08
cc_5001 ( N_RN_c_7071_n N_SN_c_8149_n ) capacitor c=0.0220464f //x=75.365 \
 //y=2.22 //x2=69.56 //y2=2.08
cc_5002 ( N_RN_c_7021_n N_SN_c_8200_n ) capacitor c=0.00583058f //x=17.645 \
 //y=2.22 //x2=11.93 //y2=1.915
cc_5003 ( N_RN_c_7038_n N_SN_c_8257_n ) capacitor c=0.00583058f //x=30.965 \
 //y=2.22 //x2=26.36 //y2=1.915
cc_5004 ( N_RN_c_7046_n N_SN_c_8357_n ) capacitor c=0.00583058f //x=46.505 \
 //y=2.22 //x2=40.79 //y2=1.915
cc_5005 ( N_RN_c_7063_n N_SN_c_8426_n ) capacitor c=0.00583058f //x=59.825 \
 //y=2.22 //x2=55.22 //y2=1.915
cc_5006 ( N_RN_c_7071_n N_SN_c_8485_n ) capacitor c=0.00583058f //x=75.365 \
 //y=2.22 //x2=69.65 //y2=1.915
cc_5007 ( N_RN_c_7095_n N_noxref_21_c_8878_n ) capacitor c=0.0179999f \
 //x=75.48 //y=2.08 //x2=76.105 //y2=3.7
cc_5008 ( N_RN_c_7083_n N_noxref_21_c_8880_n ) capacitor c=0.0044763f \
 //x=79.065 //y=2.22 //x2=84.985 //y2=3.7
cc_5009 ( N_RN_c_7096_n N_noxref_21_c_8880_n ) capacitor c=0.0213788f \
 //x=79.18 //y=2.08 //x2=84.985 //y2=3.7
cc_5010 ( N_RN_c_7095_n N_noxref_21_c_8881_n ) capacitor c=0.00179385f \
 //x=75.48 //y=2.08 //x2=76.335 //y2=3.7
cc_5011 ( N_RN_c_7071_n N_noxref_21_c_8828_n ) capacitor c=0.0186201f \
 //x=75.365 //y=2.22 //x2=65.86 //y2=2.08
cc_5012 ( N_RN_c_7071_n N_noxref_21_c_8829_n ) capacitor c=0.0209607f \
 //x=75.365 //y=2.22 //x2=70.67 //y2=2.08
cc_5013 ( N_RN_M154_noxref_g N_noxref_21_c_8841_n ) capacitor c=0.0169919f \
 //x=75.22 //y=6.02 //x2=75.355 //y2=5.155
cc_5014 ( N_RN_M155_noxref_g N_noxref_21_c_8845_n ) capacitor c=0.0194981f \
 //x=75.66 //y=6.02 //x2=76.135 //y2=5.155
cc_5015 ( N_RN_c_7265_n N_noxref_21_c_8845_n ) capacitor c=0.00201851f \
 //x=75.48 //y=4.7 //x2=76.135 //y2=5.155
cc_5016 ( N_RN_c_7781_p N_noxref_21_c_8830_n ) capacitor c=0.00371277f \
 //x=75.845 //y=1.415 //x2=76.135 //y2=1.665
cc_5017 ( N_RN_c_7782_p N_noxref_21_c_8830_n ) capacitor c=0.00457401f //x=76 \
 //y=1.26 //x2=76.135 //y2=1.665
cc_5018 ( N_RN_c_7083_n N_noxref_21_c_9017_n ) capacitor c=0.016327f \
 //x=79.065 //y=2.22 //x2=75.82 //y2=1.665
cc_5019 ( N_RN_c_7083_n N_noxref_21_c_8849_n ) capacitor c=0.0220713f \
 //x=79.065 //y=2.22 //x2=76.22 //y2=3.7
cc_5020 ( N_RN_c_7087_n N_noxref_21_c_8849_n ) capacitor c=0.0012045f \
 //x=75.595 //y=2.22 //x2=76.22 //y2=3.7
cc_5021 ( N_RN_c_7095_n N_noxref_21_c_8849_n ) capacitor c=0.0771911f \
 //x=75.48 //y=2.08 //x2=76.22 //y2=3.7
cc_5022 ( N_RN_c_7096_n N_noxref_21_c_8849_n ) capacitor c=5.91559e-19 \
 //x=79.18 //y=2.08 //x2=76.22 //y2=3.7
cc_5023 ( N_RN_c_7670_n N_noxref_21_c_8849_n ) capacitor c=0.00709342f \
 //x=75.48 //y=2.08 //x2=76.22 //y2=3.7
cc_5024 ( N_RN_c_7672_n N_noxref_21_c_8849_n ) capacitor c=0.00283672f \
 //x=75.48 //y=1.915 //x2=76.22 //y2=3.7
cc_5025 ( N_RN_c_7265_n N_noxref_21_c_8849_n ) capacitor c=0.0112909f \
 //x=75.48 //y=4.7 //x2=76.22 //y2=3.7
cc_5026 ( N_RN_c_7095_n N_noxref_21_c_9025_n ) capacitor c=0.0171303f \
 //x=75.48 //y=2.08 //x2=75.44 //y2=5.155
cc_5027 ( N_RN_c_7265_n N_noxref_21_c_9025_n ) capacitor c=0.00475601f \
 //x=75.48 //y=4.7 //x2=75.44 //y2=5.155
cc_5028 ( N_RN_c_7071_n N_noxref_21_c_8995_n ) capacitor c=3.13485e-19 \
 //x=75.365 //y=2.22 //x2=66.225 //y2=1.415
cc_5029 ( N_RN_c_7071_n N_noxref_21_c_8922_n ) capacitor c=3.13485e-19 \
 //x=75.365 //y=2.22 //x2=71.035 //y2=1.415
cc_5030 ( N_RN_c_7071_n N_noxref_21_c_8958_n ) capacitor c=0.00584491f \
 //x=75.365 //y=2.22 //x2=65.86 //y2=2.08
cc_5031 ( N_RN_c_7071_n N_noxref_21_c_8927_n ) capacitor c=0.00584491f \
 //x=75.365 //y=2.22 //x2=70.67 //y2=2.08
cc_5032 ( N_RN_c_7649_n N_noxref_21_M47_noxref_d ) capacitor c=0.00217566f \
 //x=75.47 //y=0.915 //x2=75.545 //y2=0.915
cc_5033 ( N_RN_c_7650_n N_noxref_21_M47_noxref_d ) capacitor c=0.0034598f \
 //x=75.47 //y=1.26 //x2=75.545 //y2=0.915
cc_5034 ( N_RN_c_7651_n N_noxref_21_M47_noxref_d ) capacitor c=0.00546784f \
 //x=75.47 //y=1.57 //x2=75.545 //y2=0.915
cc_5035 ( N_RN_c_7800_p N_noxref_21_M47_noxref_d ) capacitor c=0.00241102f \
 //x=75.845 //y=0.76 //x2=75.545 //y2=0.915
cc_5036 ( N_RN_c_7781_p N_noxref_21_M47_noxref_d ) capacitor c=0.0138621f \
 //x=75.845 //y=1.415 //x2=75.545 //y2=0.915
cc_5037 ( N_RN_c_7802_p N_noxref_21_M47_noxref_d ) capacitor c=0.00219619f \
 //x=76 //y=0.915 //x2=75.545 //y2=0.915
cc_5038 ( N_RN_c_7782_p N_noxref_21_M47_noxref_d ) capacitor c=0.00603828f \
 //x=76 //y=1.26 //x2=75.545 //y2=0.915
cc_5039 ( N_RN_c_7672_n N_noxref_21_M47_noxref_d ) capacitor c=0.00661782f \
 //x=75.48 //y=1.915 //x2=75.545 //y2=0.915
cc_5040 ( N_RN_M154_noxref_g N_noxref_21_M154_noxref_d ) capacitor \
 c=0.0180032f //x=75.22 //y=6.02 //x2=75.295 //y2=5.02
cc_5041 ( N_RN_M155_noxref_g N_noxref_21_M154_noxref_d ) capacitor \
 c=0.0194246f //x=75.66 //y=6.02 //x2=75.295 //y2=5.02
cc_5042 ( N_RN_c_7096_n N_noxref_22_c_9174_n ) capacitor c=0.00526349f \
 //x=79.18 //y=2.08 //x2=80.405 //y2=2.59
cc_5043 ( N_RN_c_7083_n N_noxref_22_c_9175_n ) capacitor c=0.00319026f \
 //x=79.065 //y=2.22 //x2=80.29 //y2=2.08
cc_5044 ( N_RN_c_7096_n N_noxref_22_c_9175_n ) capacitor c=0.045311f //x=79.18 \
 //y=2.08 //x2=80.29 //y2=2.08
cc_5045 ( N_RN_c_7722_n N_noxref_22_c_9175_n ) capacitor c=0.00213841f \
 //x=79.27 //y=1.915 //x2=80.29 //y2=2.08
cc_5046 ( N_RN_c_7268_n N_noxref_22_c_9175_n ) capacitor c=0.00142741f \
 //x=79.18 //y=4.7 //x2=80.29 //y2=2.08
cc_5047 ( N_RN_M158_noxref_g N_noxref_22_M160_noxref_g ) capacitor \
 c=0.0101598f //x=79.15 //y=6.02 //x2=80.03 //y2=6.02
cc_5048 ( N_RN_M159_noxref_g N_noxref_22_M160_noxref_g ) capacitor \
 c=0.0602553f //x=79.59 //y=6.02 //x2=80.03 //y2=6.02
cc_5049 ( N_RN_M159_noxref_g N_noxref_22_M161_noxref_g ) capacitor \
 c=0.0101598f //x=79.59 //y=6.02 //x2=80.47 //y2=6.02
cc_5050 ( N_RN_c_7719_n N_noxref_22_c_9232_n ) capacitor c=0.00456962f \
 //x=79.27 //y=0.91 //x2=80.28 //y2=0.915
cc_5051 ( N_RN_c_7720_n N_noxref_22_c_9233_n ) capacitor c=0.00438372f \
 //x=79.27 //y=1.22 //x2=80.28 //y2=1.26
cc_5052 ( N_RN_c_7721_n N_noxref_22_c_9234_n ) capacitor c=0.00438372f \
 //x=79.27 //y=1.45 //x2=80.28 //y2=1.57
cc_5053 ( N_RN_c_7083_n N_noxref_22_c_9235_n ) capacitor c=0.00192686f \
 //x=79.065 //y=2.22 //x2=80.29 //y2=2.08
cc_5054 ( N_RN_c_7096_n N_noxref_22_c_9235_n ) capacitor c=0.0021852f \
 //x=79.18 //y=2.08 //x2=80.29 //y2=2.08
cc_5055 ( N_RN_c_7722_n N_noxref_22_c_9235_n ) capacitor c=0.00896806f \
 //x=79.27 //y=1.915 //x2=80.29 //y2=2.08
cc_5056 ( N_RN_c_7722_n N_noxref_22_c_9238_n ) capacitor c=0.00438372f \
 //x=79.27 //y=1.915 //x2=80.29 //y2=1.915
cc_5057 ( N_RN_c_7096_n N_noxref_22_c_9222_n ) capacitor c=0.00219458f \
 //x=79.18 //y=2.08 //x2=80.29 //y2=4.7
cc_5058 ( N_RN_c_7259_n N_noxref_22_c_9222_n ) capacitor c=0.0611812f \
 //x=79.515 //y=4.79 //x2=80.29 //y2=4.7
cc_5059 ( N_RN_c_7268_n N_noxref_22_c_9222_n ) capacitor c=0.00487508f \
 //x=79.18 //y=4.7 //x2=80.29 //y2=4.7
cc_5060 ( N_RN_c_7083_n N_noxref_24_c_9437_n ) capacitor c=0.00935733f \
 //x=79.065 //y=2.22 //x2=81.145 //y2=2.22
cc_5061 ( N_RN_c_7096_n N_noxref_24_c_9478_n ) capacitor c=0.0144268f \
 //x=79.18 //y=2.08 //x2=79.285 //y2=5.155
cc_5062 ( N_RN_M158_noxref_g N_noxref_24_c_9478_n ) capacitor c=0.0165266f \
 //x=79.15 //y=6.02 //x2=79.285 //y2=5.155
cc_5063 ( N_RN_c_7268_n N_noxref_24_c_9478_n ) capacitor c=0.00322054f \
 //x=79.18 //y=4.7 //x2=79.285 //y2=5.155
cc_5064 ( N_RN_M159_noxref_g N_noxref_24_c_9484_n ) capacitor c=0.01736f \
 //x=79.59 //y=6.02 //x2=80.165 //y2=5.155
cc_5065 ( N_RN_c_7096_n N_noxref_24_c_9451_n ) capacitor c=0.00268303f \
 //x=79.18 //y=2.08 //x2=81.03 //y2=2.22
cc_5066 ( N_RN_c_7259_n N_noxref_24_c_9574_n ) capacitor c=0.00426767f \
 //x=79.515 //y=4.79 //x2=79.37 //y2=5.155
cc_5067 ( N_RN_M158_noxref_g N_noxref_24_M158_noxref_d ) capacitor \
 c=0.0180032f //x=79.15 //y=6.02 //x2=79.225 //y2=5.02
cc_5068 ( N_RN_M159_noxref_g N_noxref_24_M158_noxref_d ) capacitor \
 c=0.0180032f //x=79.59 //y=6.02 //x2=79.225 //y2=5.02
cc_5069 ( N_RN_c_7063_n N_noxref_26_c_9933_n ) capacitor c=0.00811391f \
 //x=59.825 //y=2.22 //x2=65.035 //y2=3.7
cc_5070 ( N_RN_c_7071_n N_noxref_26_c_9933_n ) capacitor c=0.00433536f \
 //x=75.365 //y=2.22 //x2=65.035 //y2=3.7
cc_5071 ( N_RN_c_7082_n N_noxref_26_c_9933_n ) capacitor c=3.18831e-19 \
 //x=60.055 //y=2.22 //x2=65.035 //y2=3.7
cc_5072 ( N_RN_c_7094_n N_noxref_26_c_9933_n ) capacitor c=0.023684f //x=59.94 \
 //y=2.08 //x2=65.035 //y2=3.7
cc_5073 ( N_RN_c_7095_n N_noxref_26_c_9912_n ) capacitor c=0.0179722f \
 //x=75.48 //y=2.08 //x2=88.315 //y2=4.07
cc_5074 ( N_RN_c_7096_n N_noxref_26_c_9912_n ) capacitor c=0.0190126f \
 //x=79.18 //y=2.08 //x2=88.315 //y2=4.07
cc_5075 ( N_RN_c_7093_n N_noxref_26_c_9944_n ) capacitor c=0.0121898f \
 //x=50.32 //y=2.08 //x2=50.425 //y2=5.155
cc_5076 ( N_RN_M122_noxref_g N_noxref_26_c_9944_n ) capacitor c=0.0163793f \
 //x=50.29 //y=6.02 //x2=50.425 //y2=5.155
cc_5077 ( N_RN_c_7263_n N_noxref_26_c_9944_n ) capacitor c=0.00309994f \
 //x=50.32 //y=4.7 //x2=50.425 //y2=5.155
cc_5078 ( N_RN_M123_noxref_g N_noxref_26_c_9950_n ) capacitor c=0.0162556f \
 //x=50.73 //y=6.02 //x2=51.305 //y2=5.155
cc_5079 ( N_RN_c_7063_n N_noxref_26_c_10146_n ) capacitor c=0.016327f \
 //x=59.825 //y=2.22 //x2=51.77 //y2=1.665
cc_5080 ( N_RN_c_7063_n N_noxref_26_c_9958_n ) capacitor c=0.0197307f \
 //x=59.825 //y=2.22 //x2=52.17 //y2=3.33
cc_5081 ( N_RN_c_7093_n N_noxref_26_c_9958_n ) capacitor c=0.00231968f \
 //x=50.32 //y=2.08 //x2=52.17 //y2=3.33
cc_5082 ( N_RN_c_7063_n N_noxref_26_c_9916_n ) capacitor c=0.0192695f \
 //x=59.825 //y=2.22 //x2=54.02 //y2=2.08
cc_5083 ( N_RN_c_7257_n N_noxref_26_c_10150_n ) capacitor c=0.00392095f \
 //x=50.655 //y=4.79 //x2=50.51 //y2=5.155
cc_5084 ( N_RN_c_7063_n N_noxref_26_c_9925_n ) capacitor c=0.011987f \
 //x=59.825 //y=2.22 //x2=53.72 //y2=1.915
cc_5085 ( N_RN_M122_noxref_g N_noxref_26_M122_noxref_d ) capacitor \
 c=0.0180032f //x=50.29 //y=6.02 //x2=50.365 //y2=5.02
cc_5086 ( N_RN_M123_noxref_g N_noxref_26_M122_noxref_d ) capacitor \
 c=0.0180032f //x=50.73 //y=6.02 //x2=50.365 //y2=5.02
cc_5087 ( N_RN_c_7528_n N_noxref_28_c_10549_n ) capacitor c=0.0167228f \
 //x=1.785 //y=0.91 //x2=2.445 //y2=0.54
cc_5088 ( N_RN_c_7204_n N_noxref_28_c_10549_n ) capacitor c=0.00534519f \
 //x=2.31 //y=0.91 //x2=2.445 //y2=0.54
cc_5089 ( N_RN_c_7021_n N_noxref_28_c_10566_n ) capacitor c=0.00387656f \
 //x=17.645 //y=2.22 //x2=2.445 //y2=1.59
cc_5090 ( N_RN_c_7032_n N_noxref_28_c_10566_n ) capacitor c=0.00354473f \
 //x=2.335 //y=2.22 //x2=2.445 //y2=1.59
cc_5091 ( N_RN_c_7088_n N_noxref_28_c_10566_n ) capacitor c=0.011736f //x=2.22 \
 //y=2.08 //x2=2.445 //y2=1.59
cc_5092 ( N_RN_c_7531_n N_noxref_28_c_10566_n ) capacitor c=0.0153695f \
 //x=1.785 //y=1.22 //x2=2.445 //y2=1.59
cc_5093 ( N_RN_c_7207_n N_noxref_28_c_10566_n ) capacitor c=0.0213278f \
 //x=2.31 //y=1.915 //x2=2.445 //y2=1.59
cc_5094 ( N_RN_c_7021_n N_noxref_28_M0_noxref_s ) capacitor c=0.00599513f \
 //x=17.645 //y=2.22 //x2=0.455 //y2=0.375
cc_5095 ( N_RN_c_7528_n N_noxref_28_M0_noxref_s ) capacitor c=0.00798959f \
 //x=1.785 //y=0.91 //x2=0.455 //y2=0.375
cc_5096 ( N_RN_c_7206_n N_noxref_28_M0_noxref_s ) capacitor c=0.00212176f \
 //x=2.31 //y=1.45 //x2=0.455 //y2=0.375
cc_5097 ( N_RN_c_7207_n N_noxref_28_M0_noxref_s ) capacitor c=0.00298115f \
 //x=2.31 //y=1.915 //x2=0.455 //y2=0.375
cc_5098 ( N_RN_c_7021_n N_noxref_29_c_10591_n ) capacitor c=0.00657782f \
 //x=17.645 //y=2.22 //x2=3.015 //y2=0.995
cc_5099 ( N_RN_c_7864_p N_noxref_29_c_10591_n ) capacitor c=2.14837e-19 \
 //x=2.155 //y=0.755 //x2=3.015 //y2=0.995
cc_5100 ( N_RN_c_7204_n N_noxref_29_c_10591_n ) capacitor c=0.00123426f \
 //x=2.31 //y=0.91 //x2=3.015 //y2=0.995
cc_5101 ( N_RN_c_7205_n N_noxref_29_c_10591_n ) capacitor c=0.0129288f \
 //x=2.31 //y=1.22 //x2=3.015 //y2=0.995
cc_5102 ( N_RN_c_7206_n N_noxref_29_c_10591_n ) capacitor c=0.00142359f \
 //x=2.31 //y=1.45 //x2=3.015 //y2=0.995
cc_5103 ( N_RN_c_7021_n N_noxref_29_c_10596_n ) capacitor c=0.00147946f \
 //x=17.645 //y=2.22 //x2=3.985 //y2=0.54
cc_5104 ( N_RN_c_7528_n N_noxref_29_M1_noxref_d ) capacitor c=0.00223875f \
 //x=1.785 //y=0.91 //x2=1.86 //y2=0.91
cc_5105 ( N_RN_c_7531_n N_noxref_29_M1_noxref_d ) capacitor c=0.00262485f \
 //x=1.785 //y=1.22 //x2=1.86 //y2=0.91
cc_5106 ( N_RN_c_7864_p N_noxref_29_M1_noxref_d ) capacitor c=0.00220746f \
 //x=2.155 //y=0.755 //x2=1.86 //y2=0.91
cc_5107 ( N_RN_c_7872_p N_noxref_29_M1_noxref_d ) capacitor c=0.00194798f \
 //x=2.155 //y=1.375 //x2=1.86 //y2=0.91
cc_5108 ( N_RN_c_7204_n N_noxref_29_M1_noxref_d ) capacitor c=0.00198465f \
 //x=2.31 //y=0.91 //x2=1.86 //y2=0.91
cc_5109 ( N_RN_c_7205_n N_noxref_29_M1_noxref_d ) capacitor c=0.00128384f \
 //x=2.31 //y=1.22 //x2=1.86 //y2=0.91
cc_5110 ( N_RN_c_7021_n N_noxref_29_M2_noxref_s ) capacitor c=0.00642985f \
 //x=17.645 //y=2.22 //x2=2.965 //y2=0.375
cc_5111 ( N_RN_c_7204_n N_noxref_29_M2_noxref_s ) capacitor c=7.21316e-19 \
 //x=2.31 //y=0.91 //x2=2.965 //y2=0.375
cc_5112 ( N_RN_c_7205_n N_noxref_29_M2_noxref_s ) capacitor c=0.00348171f \
 //x=2.31 //y=1.22 //x2=2.965 //y2=0.375
cc_5113 ( N_RN_c_7021_n N_noxref_30_c_10658_n ) capacitor c=0.00642985f \
 //x=17.645 //y=2.22 //x2=5.4 //y2=1.505
cc_5114 ( N_RN_c_7021_n N_noxref_30_c_10643_n ) capacitor c=0.0225733f \
 //x=17.645 //y=2.22 //x2=6.285 //y2=1.59
cc_5115 ( N_RN_c_7021_n N_noxref_30_c_10673_n ) capacitor c=0.0203655f \
 //x=17.645 //y=2.22 //x2=7.255 //y2=1.59
cc_5116 ( N_RN_c_7021_n N_noxref_30_M3_noxref_s ) capacitor c=0.012425f \
 //x=17.645 //y=2.22 //x2=5.265 //y2=0.375
cc_5117 ( N_RN_c_7021_n N_noxref_31_c_10692_n ) capacitor c=0.00657782f \
 //x=17.645 //y=2.22 //x2=7.825 //y2=0.995
cc_5118 ( N_RN_c_7021_n N_noxref_31_c_10697_n ) capacitor c=0.00147946f \
 //x=17.645 //y=2.22 //x2=8.795 //y2=0.54
cc_5119 ( N_RN_c_7021_n N_noxref_31_M5_noxref_s ) capacitor c=0.00642985f \
 //x=17.645 //y=2.22 //x2=7.775 //y2=0.375
cc_5120 ( N_RN_c_7021_n N_noxref_32_c_10759_n ) capacitor c=0.00642985f \
 //x=17.645 //y=2.22 //x2=10.21 //y2=1.505
cc_5121 ( N_RN_c_7021_n N_noxref_32_c_10744_n ) capacitor c=0.0225733f \
 //x=17.645 //y=2.22 //x2=11.095 //y2=1.59
cc_5122 ( N_RN_c_7021_n N_noxref_32_c_10774_n ) capacitor c=0.0203655f \
 //x=17.645 //y=2.22 //x2=12.065 //y2=1.59
cc_5123 ( N_RN_c_7021_n N_noxref_32_M6_noxref_s ) capacitor c=0.012425f \
 //x=17.645 //y=2.22 //x2=10.075 //y2=0.375
cc_5124 ( N_RN_c_7021_n N_noxref_33_c_10793_n ) capacitor c=0.00657782f \
 //x=17.645 //y=2.22 //x2=12.635 //y2=0.995
cc_5125 ( N_RN_c_7021_n N_noxref_33_c_10798_n ) capacitor c=0.00147946f \
 //x=17.645 //y=2.22 //x2=13.605 //y2=0.54
cc_5126 ( N_RN_c_7021_n N_noxref_33_M8_noxref_s ) capacitor c=0.00642985f \
 //x=17.645 //y=2.22 //x2=12.585 //y2=0.375
cc_5127 ( N_RN_c_7021_n N_noxref_34_c_10860_n ) capacitor c=0.00642985f \
 //x=17.645 //y=2.22 //x2=15.02 //y2=1.505
cc_5128 ( N_RN_c_7021_n N_noxref_34_c_10845_n ) capacitor c=0.0225733f \
 //x=17.645 //y=2.22 //x2=15.905 //y2=1.59
cc_5129 ( N_RN_c_7021_n N_noxref_34_c_10875_n ) capacitor c=0.0203655f \
 //x=17.645 //y=2.22 //x2=16.875 //y2=1.59
cc_5130 ( N_RN_c_7021_n N_noxref_34_M9_noxref_s ) capacitor c=0.012425f \
 //x=17.645 //y=2.22 //x2=14.885 //y2=0.375
cc_5131 ( N_RN_c_7021_n N_noxref_35_c_10894_n ) capacitor c=0.00657782f \
 //x=17.645 //y=2.22 //x2=17.445 //y2=0.995
cc_5132 ( N_RN_c_7033_n N_noxref_35_c_10899_n ) capacitor c=7.41833e-19 \
 //x=21.345 //y=2.22 //x2=18.415 //y2=0.54
cc_5133 ( N_RN_c_7037_n N_noxref_35_c_10899_n ) capacitor c=7.4531e-19 \
 //x=17.875 //y=2.22 //x2=18.415 //y2=0.54
cc_5134 ( N_RN_c_7089_n N_noxref_35_c_10899_n ) capacitor c=0.00204178f \
 //x=17.76 //y=2.08 //x2=18.415 //y2=0.54
cc_5135 ( N_RN_c_7295_n N_noxref_35_c_10899_n ) capacitor c=0.0194423f \
 //x=17.75 //y=0.915 //x2=18.415 //y2=0.54
cc_5136 ( N_RN_c_7301_n N_noxref_35_c_10899_n ) capacitor c=0.00656458f \
 //x=18.28 //y=0.915 //x2=18.415 //y2=0.54
cc_5137 ( N_RN_c_7304_n N_noxref_35_c_10899_n ) capacitor c=2.20712e-19 \
 //x=17.76 //y=2.08 //x2=18.415 //y2=0.54
cc_5138 ( N_RN_c_7296_n N_noxref_35_c_10909_n ) capacitor c=0.00538829f \
 //x=17.75 //y=1.26 //x2=17.53 //y2=0.995
cc_5139 ( N_RN_c_7021_n N_noxref_35_M11_noxref_s ) capacitor c=0.00642985f \
 //x=17.645 //y=2.22 //x2=17.395 //y2=0.375
cc_5140 ( N_RN_c_7295_n N_noxref_35_M11_noxref_s ) capacitor c=0.00538829f \
 //x=17.75 //y=0.915 //x2=17.395 //y2=0.375
cc_5141 ( N_RN_c_7297_n N_noxref_35_M11_noxref_s ) capacitor c=0.00538829f \
 //x=17.75 //y=1.57 //x2=17.395 //y2=0.375
cc_5142 ( N_RN_c_7301_n N_noxref_35_M11_noxref_s ) capacitor c=0.0143002f \
 //x=18.28 //y=0.915 //x2=17.395 //y2=0.375
cc_5143 ( N_RN_c_7302_n N_noxref_35_M11_noxref_s ) capacitor c=0.00290153f \
 //x=18.28 //y=1.26 //x2=17.395 //y2=0.375
cc_5144 ( N_RN_c_7033_n N_noxref_36_c_10962_n ) capacitor c=0.00642985f \
 //x=21.345 //y=2.22 //x2=19.83 //y2=1.505
cc_5145 ( N_RN_c_7033_n N_noxref_36_c_10947_n ) capacitor c=0.0225733f \
 //x=21.345 //y=2.22 //x2=20.715 //y2=1.59
cc_5146 ( N_RN_c_7211_n N_noxref_36_c_10954_n ) capacitor c=0.0167228f \
 //x=21.025 //y=0.91 //x2=21.685 //y2=0.54
cc_5147 ( N_RN_c_7216_n N_noxref_36_c_10954_n ) capacitor c=0.00534519f \
 //x=21.55 //y=0.91 //x2=21.685 //y2=0.54
cc_5148 ( N_RN_c_7033_n N_noxref_36_c_10979_n ) capacitor c=0.0139868f \
 //x=21.345 //y=2.22 //x2=21.685 //y2=1.59
cc_5149 ( N_RN_c_7038_n N_noxref_36_c_10979_n ) capacitor c=0.00387656f \
 //x=30.965 //y=2.22 //x2=21.685 //y2=1.59
cc_5150 ( N_RN_c_7045_n N_noxref_36_c_10979_n ) capacitor c=0.00251375f \
 //x=21.575 //y=2.22 //x2=21.685 //y2=1.59
cc_5151 ( N_RN_c_7090_n N_noxref_36_c_10979_n ) capacitor c=0.011736f \
 //x=21.46 //y=2.08 //x2=21.685 //y2=1.59
cc_5152 ( N_RN_c_7214_n N_noxref_36_c_10979_n ) capacitor c=0.0157358f \
 //x=21.025 //y=1.22 //x2=21.685 //y2=1.59
cc_5153 ( N_RN_c_7219_n N_noxref_36_c_10979_n ) capacitor c=0.0213278f \
 //x=21.55 //y=1.915 //x2=21.685 //y2=1.59
cc_5154 ( N_RN_c_7033_n N_noxref_36_M12_noxref_s ) capacitor c=0.00642985f \
 //x=21.345 //y=2.22 //x2=19.695 //y2=0.375
cc_5155 ( N_RN_c_7038_n N_noxref_36_M12_noxref_s ) capacitor c=0.00599513f \
 //x=30.965 //y=2.22 //x2=19.695 //y2=0.375
cc_5156 ( N_RN_c_7211_n N_noxref_36_M12_noxref_s ) capacitor c=0.00798959f \
 //x=21.025 //y=0.91 //x2=19.695 //y2=0.375
cc_5157 ( N_RN_c_7218_n N_noxref_36_M12_noxref_s ) capacitor c=0.00212176f \
 //x=21.55 //y=1.45 //x2=19.695 //y2=0.375
cc_5158 ( N_RN_c_7219_n N_noxref_36_M12_noxref_s ) capacitor c=0.00298115f \
 //x=21.55 //y=1.915 //x2=19.695 //y2=0.375
cc_5159 ( N_RN_c_7038_n N_noxref_37_c_10999_n ) capacitor c=0.00657782f \
 //x=30.965 //y=2.22 //x2=22.255 //y2=0.995
cc_5160 ( N_RN_c_7925_p N_noxref_37_c_10999_n ) capacitor c=2.14837e-19 \
 //x=21.395 //y=0.755 //x2=22.255 //y2=0.995
cc_5161 ( N_RN_c_7216_n N_noxref_37_c_10999_n ) capacitor c=0.00123426f \
 //x=21.55 //y=0.91 //x2=22.255 //y2=0.995
cc_5162 ( N_RN_c_7217_n N_noxref_37_c_10999_n ) capacitor c=0.0129288f \
 //x=21.55 //y=1.22 //x2=22.255 //y2=0.995
cc_5163 ( N_RN_c_7218_n N_noxref_37_c_10999_n ) capacitor c=0.00142359f \
 //x=21.55 //y=1.45 //x2=22.255 //y2=0.995
cc_5164 ( N_RN_c_7038_n N_noxref_37_c_11004_n ) capacitor c=0.00147946f \
 //x=30.965 //y=2.22 //x2=23.225 //y2=0.54
cc_5165 ( N_RN_c_7211_n N_noxref_37_M13_noxref_d ) capacitor c=0.00223875f \
 //x=21.025 //y=0.91 //x2=21.1 //y2=0.91
cc_5166 ( N_RN_c_7214_n N_noxref_37_M13_noxref_d ) capacitor c=0.00262485f \
 //x=21.025 //y=1.22 //x2=21.1 //y2=0.91
cc_5167 ( N_RN_c_7925_p N_noxref_37_M13_noxref_d ) capacitor c=0.00220746f \
 //x=21.395 //y=0.755 //x2=21.1 //y2=0.91
cc_5168 ( N_RN_c_7933_p N_noxref_37_M13_noxref_d ) capacitor c=0.00194798f \
 //x=21.395 //y=1.375 //x2=21.1 //y2=0.91
cc_5169 ( N_RN_c_7216_n N_noxref_37_M13_noxref_d ) capacitor c=0.00198465f \
 //x=21.55 //y=0.91 //x2=21.1 //y2=0.91
cc_5170 ( N_RN_c_7217_n N_noxref_37_M13_noxref_d ) capacitor c=0.00128384f \
 //x=21.55 //y=1.22 //x2=21.1 //y2=0.91
cc_5171 ( N_RN_c_7038_n N_noxref_37_M14_noxref_s ) capacitor c=0.00642985f \
 //x=30.965 //y=2.22 //x2=22.205 //y2=0.375
cc_5172 ( N_RN_c_7216_n N_noxref_37_M14_noxref_s ) capacitor c=7.21316e-19 \
 //x=21.55 //y=0.91 //x2=22.205 //y2=0.375
cc_5173 ( N_RN_c_7217_n N_noxref_37_M14_noxref_s ) capacitor c=0.00348171f \
 //x=21.55 //y=1.22 //x2=22.205 //y2=0.375
cc_5174 ( N_RN_c_7038_n N_noxref_38_c_11066_n ) capacitor c=0.00642985f \
 //x=30.965 //y=2.22 //x2=24.64 //y2=1.505
cc_5175 ( N_RN_c_7038_n N_noxref_38_c_11051_n ) capacitor c=0.0225733f \
 //x=30.965 //y=2.22 //x2=25.525 //y2=1.59
cc_5176 ( N_RN_c_7038_n N_noxref_38_c_11081_n ) capacitor c=0.0203655f \
 //x=30.965 //y=2.22 //x2=26.495 //y2=1.59
cc_5177 ( N_RN_c_7038_n N_noxref_38_M15_noxref_s ) capacitor c=0.012425f \
 //x=30.965 //y=2.22 //x2=24.505 //y2=0.375
cc_5178 ( N_RN_c_7038_n N_noxref_39_c_11100_n ) capacitor c=0.00657782f \
 //x=30.965 //y=2.22 //x2=27.065 //y2=0.995
cc_5179 ( N_RN_c_7038_n N_noxref_39_c_11105_n ) capacitor c=0.00147946f \
 //x=30.965 //y=2.22 //x2=28.035 //y2=0.54
cc_5180 ( N_RN_c_7038_n N_noxref_39_M17_noxref_s ) capacitor c=0.00642985f \
 //x=30.965 //y=2.22 //x2=27.015 //y2=0.375
cc_5181 ( N_RN_c_7038_n N_noxref_40_c_11167_n ) capacitor c=0.00642985f \
 //x=30.965 //y=2.22 //x2=29.45 //y2=1.505
cc_5182 ( N_RN_c_7038_n N_noxref_40_c_11152_n ) capacitor c=0.0225733f \
 //x=30.965 //y=2.22 //x2=30.335 //y2=1.59
cc_5183 ( N_RN_c_7539_n N_noxref_40_c_11159_n ) capacitor c=0.0167228f \
 //x=30.645 //y=0.91 //x2=31.305 //y2=0.54
cc_5184 ( N_RN_c_7394_n N_noxref_40_c_11159_n ) capacitor c=0.00534519f \
 //x=31.17 //y=0.91 //x2=31.305 //y2=0.54
cc_5185 ( N_RN_c_7038_n N_noxref_40_c_11184_n ) capacitor c=0.0139868f \
 //x=30.965 //y=2.22 //x2=31.305 //y2=1.59
cc_5186 ( N_RN_c_7046_n N_noxref_40_c_11184_n ) capacitor c=0.00387656f \
 //x=46.505 //y=2.22 //x2=31.305 //y2=1.59
cc_5187 ( N_RN_c_7057_n N_noxref_40_c_11184_n ) capacitor c=0.00251375f \
 //x=31.195 //y=2.22 //x2=31.305 //y2=1.59
cc_5188 ( N_RN_c_7091_n N_noxref_40_c_11184_n ) capacitor c=0.011736f \
 //x=31.08 //y=2.08 //x2=31.305 //y2=1.59
cc_5189 ( N_RN_c_7542_n N_noxref_40_c_11184_n ) capacitor c=0.0157358f \
 //x=30.645 //y=1.22 //x2=31.305 //y2=1.59
cc_5190 ( N_RN_c_7397_n N_noxref_40_c_11184_n ) capacitor c=0.0213278f \
 //x=31.17 //y=1.915 //x2=31.305 //y2=1.59
cc_5191 ( N_RN_c_7038_n N_noxref_40_M18_noxref_s ) capacitor c=0.00642985f \
 //x=30.965 //y=2.22 //x2=29.315 //y2=0.375
cc_5192 ( N_RN_c_7046_n N_noxref_40_M18_noxref_s ) capacitor c=0.00599513f \
 //x=46.505 //y=2.22 //x2=29.315 //y2=0.375
cc_5193 ( N_RN_c_7539_n N_noxref_40_M18_noxref_s ) capacitor c=0.00798959f \
 //x=30.645 //y=0.91 //x2=29.315 //y2=0.375
cc_5194 ( N_RN_c_7396_n N_noxref_40_M18_noxref_s ) capacitor c=0.00212176f \
 //x=31.17 //y=1.45 //x2=29.315 //y2=0.375
cc_5195 ( N_RN_c_7397_n N_noxref_40_M18_noxref_s ) capacitor c=0.00298115f \
 //x=31.17 //y=1.915 //x2=29.315 //y2=0.375
cc_5196 ( N_RN_c_7046_n N_noxref_41_c_11204_n ) capacitor c=0.00657782f \
 //x=46.505 //y=2.22 //x2=31.875 //y2=0.995
cc_5197 ( N_RN_c_7962_p N_noxref_41_c_11204_n ) capacitor c=2.14837e-19 \
 //x=31.015 //y=0.755 //x2=31.875 //y2=0.995
cc_5198 ( N_RN_c_7394_n N_noxref_41_c_11204_n ) capacitor c=0.00123426f \
 //x=31.17 //y=0.91 //x2=31.875 //y2=0.995
cc_5199 ( N_RN_c_7395_n N_noxref_41_c_11204_n ) capacitor c=0.0129288f \
 //x=31.17 //y=1.22 //x2=31.875 //y2=0.995
cc_5200 ( N_RN_c_7396_n N_noxref_41_c_11204_n ) capacitor c=0.00142359f \
 //x=31.17 //y=1.45 //x2=31.875 //y2=0.995
cc_5201 ( N_RN_c_7046_n N_noxref_41_c_11209_n ) capacitor c=0.00147946f \
 //x=46.505 //y=2.22 //x2=32.845 //y2=0.54
cc_5202 ( N_RN_c_7539_n N_noxref_41_M19_noxref_d ) capacitor c=0.00223875f \
 //x=30.645 //y=0.91 //x2=30.72 //y2=0.91
cc_5203 ( N_RN_c_7542_n N_noxref_41_M19_noxref_d ) capacitor c=0.00262485f \
 //x=30.645 //y=1.22 //x2=30.72 //y2=0.91
cc_5204 ( N_RN_c_7962_p N_noxref_41_M19_noxref_d ) capacitor c=0.00220746f \
 //x=31.015 //y=0.755 //x2=30.72 //y2=0.91
cc_5205 ( N_RN_c_7970_p N_noxref_41_M19_noxref_d ) capacitor c=0.00194798f \
 //x=31.015 //y=1.375 //x2=30.72 //y2=0.91
cc_5206 ( N_RN_c_7394_n N_noxref_41_M19_noxref_d ) capacitor c=0.00198465f \
 //x=31.17 //y=0.91 //x2=30.72 //y2=0.91
cc_5207 ( N_RN_c_7395_n N_noxref_41_M19_noxref_d ) capacitor c=0.00128384f \
 //x=31.17 //y=1.22 //x2=30.72 //y2=0.91
cc_5208 ( N_RN_c_7046_n N_noxref_41_M20_noxref_s ) capacitor c=0.00642985f \
 //x=46.505 //y=2.22 //x2=31.825 //y2=0.375
cc_5209 ( N_RN_c_7394_n N_noxref_41_M20_noxref_s ) capacitor c=7.21316e-19 \
 //x=31.17 //y=0.91 //x2=31.825 //y2=0.375
cc_5210 ( N_RN_c_7395_n N_noxref_41_M20_noxref_s ) capacitor c=0.00348171f \
 //x=31.17 //y=1.22 //x2=31.825 //y2=0.375
cc_5211 ( N_RN_c_7046_n N_noxref_42_c_11271_n ) capacitor c=0.00642985f \
 //x=46.505 //y=2.22 //x2=34.26 //y2=1.505
cc_5212 ( N_RN_c_7046_n N_noxref_42_c_11256_n ) capacitor c=0.0225733f \
 //x=46.505 //y=2.22 //x2=35.145 //y2=1.59
cc_5213 ( N_RN_c_7046_n N_noxref_42_c_11286_n ) capacitor c=0.0203655f \
 //x=46.505 //y=2.22 //x2=36.115 //y2=1.59
cc_5214 ( N_RN_c_7046_n N_noxref_42_M21_noxref_s ) capacitor c=0.012425f \
 //x=46.505 //y=2.22 //x2=34.125 //y2=0.375
cc_5215 ( N_RN_c_7046_n N_noxref_43_c_11305_n ) capacitor c=0.00657782f \
 //x=46.505 //y=2.22 //x2=36.685 //y2=0.995
cc_5216 ( N_RN_c_7046_n N_noxref_43_c_11310_n ) capacitor c=0.00147946f \
 //x=46.505 //y=2.22 //x2=37.655 //y2=0.54
cc_5217 ( N_RN_c_7046_n N_noxref_43_M23_noxref_s ) capacitor c=0.00642985f \
 //x=46.505 //y=2.22 //x2=36.635 //y2=0.375
cc_5218 ( N_RN_c_7046_n N_noxref_44_c_11372_n ) capacitor c=0.00642985f \
 //x=46.505 //y=2.22 //x2=39.07 //y2=1.505
cc_5219 ( N_RN_c_7046_n N_noxref_44_c_11357_n ) capacitor c=0.0225733f \
 //x=46.505 //y=2.22 //x2=39.955 //y2=1.59
cc_5220 ( N_RN_c_7046_n N_noxref_44_c_11387_n ) capacitor c=0.0203655f \
 //x=46.505 //y=2.22 //x2=40.925 //y2=1.59
cc_5221 ( N_RN_c_7046_n N_noxref_44_M24_noxref_s ) capacitor c=0.012425f \
 //x=46.505 //y=2.22 //x2=38.935 //y2=0.375
cc_5222 ( N_RN_c_7046_n N_noxref_45_c_11406_n ) capacitor c=0.00657782f \
 //x=46.505 //y=2.22 //x2=41.495 //y2=0.995
cc_5223 ( N_RN_c_7046_n N_noxref_45_c_11411_n ) capacitor c=0.00147946f \
 //x=46.505 //y=2.22 //x2=42.465 //y2=0.54
cc_5224 ( N_RN_c_7046_n N_noxref_45_M26_noxref_s ) capacitor c=0.00642985f \
 //x=46.505 //y=2.22 //x2=41.445 //y2=0.375
cc_5225 ( N_RN_c_7046_n N_noxref_46_c_11473_n ) capacitor c=0.00642985f \
 //x=46.505 //y=2.22 //x2=43.88 //y2=1.505
cc_5226 ( N_RN_c_7046_n N_noxref_46_c_11458_n ) capacitor c=0.0225733f \
 //x=46.505 //y=2.22 //x2=44.765 //y2=1.59
cc_5227 ( N_RN_c_7046_n N_noxref_46_c_11488_n ) capacitor c=0.0203655f \
 //x=46.505 //y=2.22 //x2=45.735 //y2=1.59
cc_5228 ( N_RN_c_7046_n N_noxref_46_M27_noxref_s ) capacitor c=0.012425f \
 //x=46.505 //y=2.22 //x2=43.745 //y2=0.375
cc_5229 ( N_RN_c_7046_n N_noxref_47_c_11507_n ) capacitor c=0.00657782f \
 //x=46.505 //y=2.22 //x2=46.305 //y2=0.995
cc_5230 ( N_RN_c_7058_n N_noxref_47_c_11512_n ) capacitor c=7.41833e-19 \
 //x=50.205 //y=2.22 //x2=47.275 //y2=0.54
cc_5231 ( N_RN_c_7062_n N_noxref_47_c_11512_n ) capacitor c=7.4531e-19 \
 //x=46.735 //y=2.22 //x2=47.275 //y2=0.54
cc_5232 ( N_RN_c_7092_n N_noxref_47_c_11512_n ) capacitor c=0.00204178f \
 //x=46.62 //y=2.08 //x2=47.275 //y2=0.54
cc_5233 ( N_RN_c_7441_n N_noxref_47_c_11512_n ) capacitor c=0.0194423f \
 //x=46.61 //y=0.915 //x2=47.275 //y2=0.54
cc_5234 ( N_RN_c_7447_n N_noxref_47_c_11512_n ) capacitor c=0.00656458f \
 //x=47.14 //y=0.915 //x2=47.275 //y2=0.54
cc_5235 ( N_RN_c_7450_n N_noxref_47_c_11512_n ) capacitor c=2.20712e-19 \
 //x=46.62 //y=2.08 //x2=47.275 //y2=0.54
cc_5236 ( N_RN_c_7442_n N_noxref_47_c_11522_n ) capacitor c=0.00538829f \
 //x=46.61 //y=1.26 //x2=46.39 //y2=0.995
cc_5237 ( N_RN_c_7046_n N_noxref_47_M29_noxref_s ) capacitor c=0.00642985f \
 //x=46.505 //y=2.22 //x2=46.255 //y2=0.375
cc_5238 ( N_RN_c_7441_n N_noxref_47_M29_noxref_s ) capacitor c=0.00538829f \
 //x=46.61 //y=0.915 //x2=46.255 //y2=0.375
cc_5239 ( N_RN_c_7443_n N_noxref_47_M29_noxref_s ) capacitor c=0.00538829f \
 //x=46.61 //y=1.57 //x2=46.255 //y2=0.375
cc_5240 ( N_RN_c_7447_n N_noxref_47_M29_noxref_s ) capacitor c=0.0143002f \
 //x=47.14 //y=0.915 //x2=46.255 //y2=0.375
cc_5241 ( N_RN_c_7448_n N_noxref_47_M29_noxref_s ) capacitor c=0.00290153f \
 //x=47.14 //y=1.26 //x2=46.255 //y2=0.375
cc_5242 ( N_RN_c_7058_n N_noxref_48_c_11575_n ) capacitor c=0.00642985f \
 //x=50.205 //y=2.22 //x2=48.69 //y2=1.505
cc_5243 ( N_RN_c_7058_n N_noxref_48_c_11560_n ) capacitor c=0.0225733f \
 //x=50.205 //y=2.22 //x2=49.575 //y2=1.59
cc_5244 ( N_RN_c_7401_n N_noxref_48_c_11567_n ) capacitor c=0.0167228f \
 //x=49.885 //y=0.91 //x2=50.545 //y2=0.54
cc_5245 ( N_RN_c_7406_n N_noxref_48_c_11567_n ) capacitor c=0.00534519f \
 //x=50.41 //y=0.91 //x2=50.545 //y2=0.54
cc_5246 ( N_RN_c_7058_n N_noxref_48_c_11591_n ) capacitor c=0.0139868f \
 //x=50.205 //y=2.22 //x2=50.545 //y2=1.59
cc_5247 ( N_RN_c_7063_n N_noxref_48_c_11591_n ) capacitor c=0.00387656f \
 //x=59.825 //y=2.22 //x2=50.545 //y2=1.59
cc_5248 ( N_RN_c_7070_n N_noxref_48_c_11591_n ) capacitor c=0.00251375f \
 //x=50.435 //y=2.22 //x2=50.545 //y2=1.59
cc_5249 ( N_RN_c_7093_n N_noxref_48_c_11591_n ) capacitor c=0.011736f \
 //x=50.32 //y=2.08 //x2=50.545 //y2=1.59
cc_5250 ( N_RN_c_7404_n N_noxref_48_c_11591_n ) capacitor c=0.0157358f \
 //x=49.885 //y=1.22 //x2=50.545 //y2=1.59
cc_5251 ( N_RN_c_7409_n N_noxref_48_c_11591_n ) capacitor c=0.0213278f \
 //x=50.41 //y=1.915 //x2=50.545 //y2=1.59
cc_5252 ( N_RN_c_7058_n N_noxref_48_M30_noxref_s ) capacitor c=0.00642985f \
 //x=50.205 //y=2.22 //x2=48.555 //y2=0.375
cc_5253 ( N_RN_c_7063_n N_noxref_48_M30_noxref_s ) capacitor c=0.00599513f \
 //x=59.825 //y=2.22 //x2=48.555 //y2=0.375
cc_5254 ( N_RN_c_7401_n N_noxref_48_M30_noxref_s ) capacitor c=0.00798959f \
 //x=49.885 //y=0.91 //x2=48.555 //y2=0.375
cc_5255 ( N_RN_c_7408_n N_noxref_48_M30_noxref_s ) capacitor c=0.00212176f \
 //x=50.41 //y=1.45 //x2=48.555 //y2=0.375
cc_5256 ( N_RN_c_7409_n N_noxref_48_M30_noxref_s ) capacitor c=0.00298115f \
 //x=50.41 //y=1.915 //x2=48.555 //y2=0.375
cc_5257 ( N_RN_c_7063_n N_noxref_49_c_11612_n ) capacitor c=0.00657782f \
 //x=59.825 //y=2.22 //x2=51.115 //y2=0.995
cc_5258 ( N_RN_c_8023_p N_noxref_49_c_11612_n ) capacitor c=2.14837e-19 \
 //x=50.255 //y=0.755 //x2=51.115 //y2=0.995
cc_5259 ( N_RN_c_7406_n N_noxref_49_c_11612_n ) capacitor c=0.00123426f \
 //x=50.41 //y=0.91 //x2=51.115 //y2=0.995
cc_5260 ( N_RN_c_7407_n N_noxref_49_c_11612_n ) capacitor c=0.0129288f \
 //x=50.41 //y=1.22 //x2=51.115 //y2=0.995
cc_5261 ( N_RN_c_7408_n N_noxref_49_c_11612_n ) capacitor c=0.00142359f \
 //x=50.41 //y=1.45 //x2=51.115 //y2=0.995
cc_5262 ( N_RN_c_7063_n N_noxref_49_c_11617_n ) capacitor c=0.00147946f \
 //x=59.825 //y=2.22 //x2=52.085 //y2=0.54
cc_5263 ( N_RN_c_7401_n N_noxref_49_M31_noxref_d ) capacitor c=0.00223875f \
 //x=49.885 //y=0.91 //x2=49.96 //y2=0.91
cc_5264 ( N_RN_c_7404_n N_noxref_49_M31_noxref_d ) capacitor c=0.00262485f \
 //x=49.885 //y=1.22 //x2=49.96 //y2=0.91
cc_5265 ( N_RN_c_8023_p N_noxref_49_M31_noxref_d ) capacitor c=0.00220746f \
 //x=50.255 //y=0.755 //x2=49.96 //y2=0.91
cc_5266 ( N_RN_c_8031_p N_noxref_49_M31_noxref_d ) capacitor c=0.00194798f \
 //x=50.255 //y=1.375 //x2=49.96 //y2=0.91
cc_5267 ( N_RN_c_7406_n N_noxref_49_M31_noxref_d ) capacitor c=0.00198465f \
 //x=50.41 //y=0.91 //x2=49.96 //y2=0.91
cc_5268 ( N_RN_c_7407_n N_noxref_49_M31_noxref_d ) capacitor c=0.00128384f \
 //x=50.41 //y=1.22 //x2=49.96 //y2=0.91
cc_5269 ( N_RN_c_7063_n N_noxref_49_M32_noxref_s ) capacitor c=0.00642985f \
 //x=59.825 //y=2.22 //x2=51.065 //y2=0.375
cc_5270 ( N_RN_c_7406_n N_noxref_49_M32_noxref_s ) capacitor c=7.21316e-19 \
 //x=50.41 //y=0.91 //x2=51.065 //y2=0.375
cc_5271 ( N_RN_c_7407_n N_noxref_49_M32_noxref_s ) capacitor c=0.00348171f \
 //x=50.41 //y=1.22 //x2=51.065 //y2=0.375
cc_5272 ( N_RN_c_7063_n N_noxref_50_c_11680_n ) capacitor c=0.00642985f \
 //x=59.825 //y=2.22 //x2=53.5 //y2=1.505
cc_5273 ( N_RN_c_7063_n N_noxref_50_c_11664_n ) capacitor c=0.0225733f \
 //x=59.825 //y=2.22 //x2=54.385 //y2=1.59
cc_5274 ( N_RN_c_7063_n N_noxref_50_c_11682_n ) capacitor c=0.0203655f \
 //x=59.825 //y=2.22 //x2=55.355 //y2=1.59
cc_5275 ( N_RN_c_7063_n N_noxref_50_M33_noxref_s ) capacitor c=0.012425f \
 //x=59.825 //y=2.22 //x2=53.365 //y2=0.375
cc_5276 ( N_RN_c_7063_n N_noxref_51_c_11713_n ) capacitor c=0.00657782f \
 //x=59.825 //y=2.22 //x2=55.925 //y2=0.995
cc_5277 ( N_RN_c_7063_n N_noxref_51_c_11718_n ) capacitor c=0.00147946f \
 //x=59.825 //y=2.22 //x2=56.895 //y2=0.54
cc_5278 ( N_RN_c_7063_n N_noxref_51_M35_noxref_s ) capacitor c=0.00642985f \
 //x=59.825 //y=2.22 //x2=55.875 //y2=0.375
cc_5279 ( N_RN_c_7063_n N_noxref_52_c_11780_n ) capacitor c=0.00642985f \
 //x=59.825 //y=2.22 //x2=58.31 //y2=1.505
cc_5280 ( N_RN_c_7063_n N_noxref_52_c_11765_n ) capacitor c=0.0225733f \
 //x=59.825 //y=2.22 //x2=59.195 //y2=1.59
cc_5281 ( N_RN_c_7549_n N_noxref_52_c_11772_n ) capacitor c=0.0167228f \
 //x=59.505 //y=0.91 //x2=60.165 //y2=0.54
cc_5282 ( N_RN_c_7554_n N_noxref_52_c_11772_n ) capacitor c=0.00534519f \
 //x=60.03 //y=0.91 //x2=60.165 //y2=0.54
cc_5283 ( N_RN_c_7063_n N_noxref_52_c_11797_n ) capacitor c=0.0139868f \
 //x=59.825 //y=2.22 //x2=60.165 //y2=1.59
cc_5284 ( N_RN_c_7071_n N_noxref_52_c_11797_n ) capacitor c=0.00387656f \
 //x=75.365 //y=2.22 //x2=60.165 //y2=1.59
cc_5285 ( N_RN_c_7082_n N_noxref_52_c_11797_n ) capacitor c=0.00251375f \
 //x=60.055 //y=2.22 //x2=60.165 //y2=1.59
cc_5286 ( N_RN_c_7094_n N_noxref_52_c_11797_n ) capacitor c=0.011736f \
 //x=59.94 //y=2.08 //x2=60.165 //y2=1.59
cc_5287 ( N_RN_c_7552_n N_noxref_52_c_11797_n ) capacitor c=0.0157358f \
 //x=59.505 //y=1.22 //x2=60.165 //y2=1.59
cc_5288 ( N_RN_c_7557_n N_noxref_52_c_11797_n ) capacitor c=0.0213278f \
 //x=60.03 //y=1.915 //x2=60.165 //y2=1.59
cc_5289 ( N_RN_c_7063_n N_noxref_52_M36_noxref_s ) capacitor c=0.00642985f \
 //x=59.825 //y=2.22 //x2=58.175 //y2=0.375
cc_5290 ( N_RN_c_7071_n N_noxref_52_M36_noxref_s ) capacitor c=0.00599513f \
 //x=75.365 //y=2.22 //x2=58.175 //y2=0.375
cc_5291 ( N_RN_c_7549_n N_noxref_52_M36_noxref_s ) capacitor c=0.00798959f \
 //x=59.505 //y=0.91 //x2=58.175 //y2=0.375
cc_5292 ( N_RN_c_7556_n N_noxref_52_M36_noxref_s ) capacitor c=0.00212176f \
 //x=60.03 //y=1.45 //x2=58.175 //y2=0.375
cc_5293 ( N_RN_c_7557_n N_noxref_52_M36_noxref_s ) capacitor c=0.00298115f \
 //x=60.03 //y=1.915 //x2=58.175 //y2=0.375
cc_5294 ( N_RN_c_7071_n N_noxref_53_c_11817_n ) capacitor c=0.00657782f \
 //x=75.365 //y=2.22 //x2=60.735 //y2=0.995
cc_5295 ( N_RN_c_8060_p N_noxref_53_c_11817_n ) capacitor c=2.14837e-19 \
 //x=59.875 //y=0.755 //x2=60.735 //y2=0.995
cc_5296 ( N_RN_c_7554_n N_noxref_53_c_11817_n ) capacitor c=0.00123426f \
 //x=60.03 //y=0.91 //x2=60.735 //y2=0.995
cc_5297 ( N_RN_c_7555_n N_noxref_53_c_11817_n ) capacitor c=0.0129288f \
 //x=60.03 //y=1.22 //x2=60.735 //y2=0.995
cc_5298 ( N_RN_c_7556_n N_noxref_53_c_11817_n ) capacitor c=0.00142359f \
 //x=60.03 //y=1.45 //x2=60.735 //y2=0.995
cc_5299 ( N_RN_c_7071_n N_noxref_53_c_11822_n ) capacitor c=0.00147946f \
 //x=75.365 //y=2.22 //x2=61.705 //y2=0.54
cc_5300 ( N_RN_c_7549_n N_noxref_53_M37_noxref_d ) capacitor c=0.00223875f \
 //x=59.505 //y=0.91 //x2=59.58 //y2=0.91
cc_5301 ( N_RN_c_7552_n N_noxref_53_M37_noxref_d ) capacitor c=0.00262485f \
 //x=59.505 //y=1.22 //x2=59.58 //y2=0.91
cc_5302 ( N_RN_c_8060_p N_noxref_53_M37_noxref_d ) capacitor c=0.00220746f \
 //x=59.875 //y=0.755 //x2=59.58 //y2=0.91
cc_5303 ( N_RN_c_8068_p N_noxref_53_M37_noxref_d ) capacitor c=0.00194798f \
 //x=59.875 //y=1.375 //x2=59.58 //y2=0.91
cc_5304 ( N_RN_c_7554_n N_noxref_53_M37_noxref_d ) capacitor c=0.00198465f \
 //x=60.03 //y=0.91 //x2=59.58 //y2=0.91
cc_5305 ( N_RN_c_7555_n N_noxref_53_M37_noxref_d ) capacitor c=0.00128384f \
 //x=60.03 //y=1.22 //x2=59.58 //y2=0.91
cc_5306 ( N_RN_c_7071_n N_noxref_53_M38_noxref_s ) capacitor c=0.00642985f \
 //x=75.365 //y=2.22 //x2=60.685 //y2=0.375
cc_5307 ( N_RN_c_7554_n N_noxref_53_M38_noxref_s ) capacitor c=7.21316e-19 \
 //x=60.03 //y=0.91 //x2=60.685 //y2=0.375
cc_5308 ( N_RN_c_7555_n N_noxref_53_M38_noxref_s ) capacitor c=0.00348171f \
 //x=60.03 //y=1.22 //x2=60.685 //y2=0.375
cc_5309 ( N_RN_c_7071_n N_noxref_54_c_11884_n ) capacitor c=0.00642985f \
 //x=75.365 //y=2.22 //x2=63.12 //y2=1.505
cc_5310 ( N_RN_c_7071_n N_noxref_54_c_11869_n ) capacitor c=0.0225733f \
 //x=75.365 //y=2.22 //x2=64.005 //y2=1.59
cc_5311 ( N_RN_c_7071_n N_noxref_54_c_11898_n ) capacitor c=0.0203655f \
 //x=75.365 //y=2.22 //x2=64.975 //y2=1.59
cc_5312 ( N_RN_c_7071_n N_noxref_54_M39_noxref_s ) capacitor c=0.012425f \
 //x=75.365 //y=2.22 //x2=62.985 //y2=0.375
cc_5313 ( N_RN_c_7071_n N_noxref_55_c_11918_n ) capacitor c=0.00657782f \
 //x=75.365 //y=2.22 //x2=65.545 //y2=0.995
cc_5314 ( N_RN_c_7071_n N_noxref_55_c_11923_n ) capacitor c=0.00147946f \
 //x=75.365 //y=2.22 //x2=66.515 //y2=0.54
cc_5315 ( N_RN_c_7071_n N_noxref_55_M41_noxref_s ) capacitor c=0.00642985f \
 //x=75.365 //y=2.22 //x2=65.495 //y2=0.375
cc_5316 ( N_RN_c_7071_n N_noxref_56_c_11985_n ) capacitor c=0.00642985f \
 //x=75.365 //y=2.22 //x2=67.93 //y2=1.505
cc_5317 ( N_RN_c_7071_n N_noxref_56_c_11970_n ) capacitor c=0.0225733f \
 //x=75.365 //y=2.22 //x2=68.815 //y2=1.59
cc_5318 ( N_RN_c_7071_n N_noxref_56_c_12000_n ) capacitor c=0.0203655f \
 //x=75.365 //y=2.22 //x2=69.785 //y2=1.59
cc_5319 ( N_RN_c_7071_n N_noxref_56_M42_noxref_s ) capacitor c=0.012425f \
 //x=75.365 //y=2.22 //x2=67.795 //y2=0.375
cc_5320 ( N_RN_c_7071_n N_noxref_57_c_12019_n ) capacitor c=0.00657782f \
 //x=75.365 //y=2.22 //x2=70.355 //y2=0.995
cc_5321 ( N_RN_c_7071_n N_noxref_57_c_12024_n ) capacitor c=0.00147946f \
 //x=75.365 //y=2.22 //x2=71.325 //y2=0.54
cc_5322 ( N_RN_c_7071_n N_noxref_57_M44_noxref_s ) capacitor c=0.00642985f \
 //x=75.365 //y=2.22 //x2=70.305 //y2=0.375
cc_5323 ( N_RN_c_7071_n N_noxref_58_c_12086_n ) capacitor c=0.00642985f \
 //x=75.365 //y=2.22 //x2=72.74 //y2=1.505
cc_5324 ( N_RN_c_7071_n N_noxref_58_c_12071_n ) capacitor c=0.0225733f \
 //x=75.365 //y=2.22 //x2=73.625 //y2=1.59
cc_5325 ( N_RN_c_7071_n N_noxref_58_c_12100_n ) capacitor c=0.0203655f \
 //x=75.365 //y=2.22 //x2=74.595 //y2=1.59
cc_5326 ( N_RN_c_7071_n N_noxref_58_M45_noxref_s ) capacitor c=0.012425f \
 //x=75.365 //y=2.22 //x2=72.605 //y2=0.375
cc_5327 ( N_RN_c_7071_n N_noxref_59_c_12120_n ) capacitor c=0.00657782f \
 //x=75.365 //y=2.22 //x2=75.165 //y2=0.995
cc_5328 ( N_RN_c_7083_n N_noxref_59_c_12125_n ) capacitor c=7.41833e-19 \
 //x=79.065 //y=2.22 //x2=76.135 //y2=0.54
cc_5329 ( N_RN_c_7087_n N_noxref_59_c_12125_n ) capacitor c=7.4531e-19 \
 //x=75.595 //y=2.22 //x2=76.135 //y2=0.54
cc_5330 ( N_RN_c_7095_n N_noxref_59_c_12125_n ) capacitor c=0.00204178f \
 //x=75.48 //y=2.08 //x2=76.135 //y2=0.54
cc_5331 ( N_RN_c_7649_n N_noxref_59_c_12125_n ) capacitor c=0.0194423f \
 //x=75.47 //y=0.915 //x2=76.135 //y2=0.54
cc_5332 ( N_RN_c_7802_p N_noxref_59_c_12125_n ) capacitor c=0.00656458f //x=76 \
 //y=0.915 //x2=76.135 //y2=0.54
cc_5333 ( N_RN_c_7670_n N_noxref_59_c_12125_n ) capacitor c=2.20712e-19 \
 //x=75.48 //y=2.08 //x2=76.135 //y2=0.54
cc_5334 ( N_RN_c_7650_n N_noxref_59_c_12152_n ) capacitor c=0.00538829f \
 //x=75.47 //y=1.26 //x2=75.25 //y2=0.995
cc_5335 ( N_RN_c_7071_n N_noxref_59_M47_noxref_s ) capacitor c=0.00642985f \
 //x=75.365 //y=2.22 //x2=75.115 //y2=0.375
cc_5336 ( N_RN_c_7649_n N_noxref_59_M47_noxref_s ) capacitor c=0.00538829f \
 //x=75.47 //y=0.915 //x2=75.115 //y2=0.375
cc_5337 ( N_RN_c_7651_n N_noxref_59_M47_noxref_s ) capacitor c=0.00538829f \
 //x=75.47 //y=1.57 //x2=75.115 //y2=0.375
cc_5338 ( N_RN_c_7802_p N_noxref_59_M47_noxref_s ) capacitor c=0.0143002f \
 //x=76 //y=0.915 //x2=75.115 //y2=0.375
cc_5339 ( N_RN_c_7782_p N_noxref_59_M47_noxref_s ) capacitor c=0.00290153f \
 //x=76 //y=1.26 //x2=75.115 //y2=0.375
cc_5340 ( N_RN_c_7083_n N_noxref_60_c_12188_n ) capacitor c=0.00642985f \
 //x=79.065 //y=2.22 //x2=77.55 //y2=1.505
cc_5341 ( N_RN_c_7083_n N_noxref_60_c_12173_n ) capacitor c=0.0225733f \
 //x=79.065 //y=2.22 //x2=78.435 //y2=1.59
cc_5342 ( N_RN_c_7714_n N_noxref_60_c_12180_n ) capacitor c=0.0167228f \
 //x=78.745 //y=0.91 //x2=79.405 //y2=0.54
cc_5343 ( N_RN_c_7719_n N_noxref_60_c_12180_n ) capacitor c=0.00534519f \
 //x=79.27 //y=0.91 //x2=79.405 //y2=0.54
cc_5344 ( N_RN_c_7083_n N_noxref_60_c_12202_n ) capacitor c=0.0178105f \
 //x=79.065 //y=2.22 //x2=79.405 //y2=1.59
cc_5345 ( N_RN_c_7096_n N_noxref_60_c_12202_n ) capacitor c=0.011736f \
 //x=79.18 //y=2.08 //x2=79.405 //y2=1.59
cc_5346 ( N_RN_c_7717_n N_noxref_60_c_12202_n ) capacitor c=0.0157358f \
 //x=78.745 //y=1.22 //x2=79.405 //y2=1.59
cc_5347 ( N_RN_c_7722_n N_noxref_60_c_12202_n ) capacitor c=0.0215856f \
 //x=79.27 //y=1.915 //x2=79.405 //y2=1.59
cc_5348 ( N_RN_c_7083_n N_noxref_60_M48_noxref_s ) capacitor c=0.00642985f \
 //x=79.065 //y=2.22 //x2=77.415 //y2=0.375
cc_5349 ( N_RN_c_7714_n N_noxref_60_M48_noxref_s ) capacitor c=0.00798959f \
 //x=78.745 //y=0.91 //x2=77.415 //y2=0.375
cc_5350 ( N_RN_c_7721_n N_noxref_60_M48_noxref_s ) capacitor c=0.00212176f \
 //x=79.27 //y=1.45 //x2=77.415 //y2=0.375
cc_5351 ( N_RN_c_7722_n N_noxref_60_M48_noxref_s ) capacitor c=0.00298115f \
 //x=79.27 //y=1.915 //x2=77.415 //y2=0.375
cc_5352 ( N_RN_c_8117_p N_noxref_61_c_12224_n ) capacitor c=2.14837e-19 \
 //x=79.115 //y=0.755 //x2=79.975 //y2=0.995
cc_5353 ( N_RN_c_7719_n N_noxref_61_c_12224_n ) capacitor c=0.00123426f \
 //x=79.27 //y=0.91 //x2=79.975 //y2=0.995
cc_5354 ( N_RN_c_7720_n N_noxref_61_c_12224_n ) capacitor c=0.0129288f \
 //x=79.27 //y=1.22 //x2=79.975 //y2=0.995
cc_5355 ( N_RN_c_7721_n N_noxref_61_c_12224_n ) capacitor c=0.00142359f \
 //x=79.27 //y=1.45 //x2=79.975 //y2=0.995
cc_5356 ( N_RN_c_7714_n N_noxref_61_M49_noxref_d ) capacitor c=0.00223875f \
 //x=78.745 //y=0.91 //x2=78.82 //y2=0.91
cc_5357 ( N_RN_c_7717_n N_noxref_61_M49_noxref_d ) capacitor c=0.00262485f \
 //x=78.745 //y=1.22 //x2=78.82 //y2=0.91
cc_5358 ( N_RN_c_8117_p N_noxref_61_M49_noxref_d ) capacitor c=0.00220746f \
 //x=79.115 //y=0.755 //x2=78.82 //y2=0.91
cc_5359 ( N_RN_c_8124_p N_noxref_61_M49_noxref_d ) capacitor c=0.00194798f \
 //x=79.115 //y=1.375 //x2=78.82 //y2=0.91
cc_5360 ( N_RN_c_7719_n N_noxref_61_M49_noxref_d ) capacitor c=0.00198465f \
 //x=79.27 //y=0.91 //x2=78.82 //y2=0.91
cc_5361 ( N_RN_c_7720_n N_noxref_61_M49_noxref_d ) capacitor c=0.00128384f \
 //x=79.27 //y=1.22 //x2=78.82 //y2=0.91
cc_5362 ( N_RN_c_7719_n N_noxref_61_M50_noxref_s ) capacitor c=7.21316e-19 \
 //x=79.27 //y=0.91 //x2=79.925 //y2=0.375
cc_5363 ( N_RN_c_7720_n N_noxref_61_M50_noxref_s ) capacitor c=0.00348171f \
 //x=79.27 //y=1.22 //x2=79.925 //y2=0.375
cc_5364 ( N_SN_c_8138_n N_noxref_21_c_8898_n ) capacitor c=0.0259591f \
 //x=69.445 //y=2.96 //x2=70.555 //y2=3.7
cc_5365 ( N_SN_c_8141_n N_noxref_21_c_8898_n ) capacitor c=0.0092394f \
 //x=83.875 //y=2.96 //x2=70.555 //y2=3.7
cc_5366 ( N_SN_c_8468_n N_noxref_21_c_8898_n ) capacitor c=6.65965e-19 \
 //x=69.675 //y=2.96 //x2=70.555 //y2=3.7
cc_5367 ( N_SN_c_8149_n N_noxref_21_c_8898_n ) capacitor c=0.0190398f \
 //x=69.56 //y=2.08 //x2=70.555 //y2=3.7
cc_5368 ( N_SN_c_8138_n N_noxref_21_c_8935_n ) capacitor c=8.32553e-19 \
 //x=69.445 //y=2.96 //x2=65.975 //y2=3.7
cc_5369 ( N_SN_c_8141_n N_noxref_21_c_8878_n ) capacitor c=0.041794f \
 //x=83.875 //y=2.96 //x2=76.105 //y2=3.7
cc_5370 ( N_SN_c_8141_n N_noxref_21_c_8905_n ) capacitor c=6.03896e-19 \
 //x=83.875 //y=2.96 //x2=70.785 //y2=3.7
cc_5371 ( N_SN_c_8149_n N_noxref_21_c_8905_n ) capacitor c=0.00128547f \
 //x=69.56 //y=2.08 //x2=70.785 //y2=3.7
cc_5372 ( N_SN_c_8141_n N_noxref_21_c_8880_n ) capacitor c=0.267326f \
 //x=83.875 //y=2.96 //x2=84.985 //y2=3.7
cc_5373 ( N_SN_c_8150_n N_noxref_21_c_8880_n ) capacitor c=0.0229819f \
 //x=83.99 //y=2.08 //x2=84.985 //y2=3.7
cc_5374 ( N_SN_c_8141_n N_noxref_21_c_8881_n ) capacitor c=4.80612e-19 \
 //x=83.875 //y=2.96 //x2=76.335 //y2=3.7
cc_5375 ( N_SN_c_8138_n N_noxref_21_c_8828_n ) capacitor c=0.0179917f \
 //x=69.445 //y=2.96 //x2=65.86 //y2=2.08
cc_5376 ( N_SN_c_8141_n N_noxref_21_c_8829_n ) capacitor c=0.0202855f \
 //x=83.875 //y=2.96 //x2=70.67 //y2=2.08
cc_5377 ( N_SN_c_8468_n N_noxref_21_c_8829_n ) capacitor c=0.00128547f \
 //x=69.675 //y=2.96 //x2=70.67 //y2=2.08
cc_5378 ( N_SN_c_8149_n N_noxref_21_c_8829_n ) capacitor c=0.0413563f \
 //x=69.56 //y=2.08 //x2=70.67 //y2=2.08
cc_5379 ( N_SN_c_8485_n N_noxref_21_c_8829_n ) capacitor c=0.00205895f \
 //x=69.65 //y=1.915 //x2=70.67 //y2=2.08
cc_5380 ( N_SN_c_8270_n N_noxref_21_c_8829_n ) capacitor c=0.00142741f \
 //x=69.56 //y=4.7 //x2=70.67 //y2=2.08
cc_5381 ( N_SN_c_8141_n N_noxref_21_c_8849_n ) capacitor c=0.0210712f \
 //x=83.875 //y=2.96 //x2=76.22 //y2=3.7
cc_5382 ( N_SN_c_8141_n N_noxref_21_c_8831_n ) capacitor c=0.00526349f \
 //x=83.875 //y=2.96 //x2=85.1 //y2=2.08
cc_5383 ( N_SN_c_8150_n N_noxref_21_c_8831_n ) capacitor c=0.044554f //x=83.99 \
 //y=2.08 //x2=85.1 //y2=2.08
cc_5384 ( N_SN_c_8598_p N_noxref_21_c_8831_n ) capacitor c=0.00205895f \
 //x=84.08 //y=1.915 //x2=85.1 //y2=2.08
cc_5385 ( N_SN_c_8271_n N_noxref_21_c_8831_n ) capacitor c=0.00142741f \
 //x=83.99 //y=4.7 //x2=85.1 //y2=2.08
cc_5386 ( N_SN_M146_noxref_g N_noxref_21_M148_noxref_g ) capacitor \
 c=0.0100903f //x=69.53 //y=6.02 //x2=70.41 //y2=6.02
cc_5387 ( N_SN_M147_noxref_g N_noxref_21_M148_noxref_g ) capacitor \
 c=0.0600064f //x=69.97 //y=6.02 //x2=70.41 //y2=6.02
cc_5388 ( N_SN_M147_noxref_g N_noxref_21_M149_noxref_g ) capacitor \
 c=0.0100903f //x=69.97 //y=6.02 //x2=70.85 //y2=6.02
cc_5389 ( N_SN_M164_noxref_g N_noxref_21_M166_noxref_g ) capacitor \
 c=0.0101598f //x=83.96 //y=6.02 //x2=84.84 //y2=6.02
cc_5390 ( N_SN_M165_noxref_g N_noxref_21_M166_noxref_g ) capacitor \
 c=0.0602553f //x=84.4 //y=6.02 //x2=84.84 //y2=6.02
cc_5391 ( N_SN_M165_noxref_g N_noxref_21_M167_noxref_g ) capacitor \
 c=0.0101598f //x=84.4 //y=6.02 //x2=85.28 //y2=6.02
cc_5392 ( N_SN_c_8482_n N_noxref_21_c_8918_n ) capacitor c=0.00456962f \
 //x=69.65 //y=0.91 //x2=70.66 //y2=0.915
cc_5393 ( N_SN_c_8483_n N_noxref_21_c_8919_n ) capacitor c=0.00438372f \
 //x=69.65 //y=1.22 //x2=70.66 //y2=1.26
cc_5394 ( N_SN_c_8484_n N_noxref_21_c_8920_n ) capacitor c=0.00438372f \
 //x=69.65 //y=1.45 //x2=70.66 //y2=1.57
cc_5395 ( N_SN_c_8609_p N_noxref_21_c_9072_n ) capacitor c=0.00456962f \
 //x=84.08 //y=0.91 //x2=85.09 //y2=0.915
cc_5396 ( N_SN_c_8610_p N_noxref_21_c_9073_n ) capacitor c=0.00438372f \
 //x=84.08 //y=1.22 //x2=85.09 //y2=1.26
cc_5397 ( N_SN_c_8611_p N_noxref_21_c_9074_n ) capacitor c=0.00438372f \
 //x=84.08 //y=1.45 //x2=85.09 //y2=1.57
cc_5398 ( N_SN_c_8149_n N_noxref_21_c_8927_n ) capacitor c=0.00201097f \
 //x=69.56 //y=2.08 //x2=70.67 //y2=2.08
cc_5399 ( N_SN_c_8485_n N_noxref_21_c_8927_n ) capacitor c=0.00828003f \
 //x=69.65 //y=1.915 //x2=70.67 //y2=2.08
cc_5400 ( N_SN_c_8485_n N_noxref_21_c_8928_n ) capacitor c=0.00438372f \
 //x=69.65 //y=1.915 //x2=70.67 //y2=1.915
cc_5401 ( N_SN_c_8149_n N_noxref_21_c_8896_n ) capacitor c=0.00197875f \
 //x=69.56 //y=2.08 //x2=70.67 //y2=4.7
cc_5402 ( N_SN_c_8262_n N_noxref_21_c_8896_n ) capacitor c=0.0609323f \
 //x=69.895 //y=4.79 //x2=70.67 //y2=4.7
cc_5403 ( N_SN_c_8270_n N_noxref_21_c_8896_n ) capacitor c=0.00487508f \
 //x=69.56 //y=4.7 //x2=70.67 //y2=4.7
cc_5404 ( N_SN_c_8150_n N_noxref_21_c_9081_n ) capacitor c=0.00201097f \
 //x=83.99 //y=2.08 //x2=85.1 //y2=2.08
cc_5405 ( N_SN_c_8598_p N_noxref_21_c_9081_n ) capacitor c=0.00828003f \
 //x=84.08 //y=1.915 //x2=85.1 //y2=2.08
cc_5406 ( N_SN_c_8598_p N_noxref_21_c_9083_n ) capacitor c=0.00438372f \
 //x=84.08 //y=1.915 //x2=85.1 //y2=1.915
cc_5407 ( N_SN_c_8150_n N_noxref_21_c_8897_n ) capacitor c=0.00219458f \
 //x=83.99 //y=2.08 //x2=85.1 //y2=4.7
cc_5408 ( N_SN_c_8263_n N_noxref_21_c_8897_n ) capacitor c=0.0611812f \
 //x=84.325 //y=4.79 //x2=85.1 //y2=4.7
cc_5409 ( N_SN_c_8271_n N_noxref_21_c_8897_n ) capacitor c=0.00487508f \
 //x=83.99 //y=4.7 //x2=85.1 //y2=4.7
cc_5410 ( N_SN_c_8141_n N_noxref_22_c_9171_n ) capacitor c=0.332921f \
 //x=83.875 //y=2.96 //x2=85.725 //y2=2.59
cc_5411 ( N_SN_c_8150_n N_noxref_22_c_9171_n ) capacitor c=0.0208352f \
 //x=83.99 //y=2.08 //x2=85.725 //y2=2.59
cc_5412 ( N_SN_c_8141_n N_noxref_22_c_9174_n ) capacitor c=0.0291665f \
 //x=83.875 //y=2.96 //x2=80.405 //y2=2.59
cc_5413 ( N_SN_c_8141_n N_noxref_22_c_9175_n ) capacitor c=0.0221691f \
 //x=83.875 //y=2.96 //x2=80.29 //y2=2.08
cc_5414 ( N_SN_c_8150_n N_noxref_22_c_9180_n ) capacitor c=0.0146f //x=83.99 \
 //y=2.08 //x2=84.095 //y2=5.155
cc_5415 ( N_SN_M164_noxref_g N_noxref_22_c_9180_n ) capacitor c=0.0165266f \
 //x=83.96 //y=6.02 //x2=84.095 //y2=5.155
cc_5416 ( N_SN_c_8271_n N_noxref_22_c_9180_n ) capacitor c=0.00322054f \
 //x=83.99 //y=4.7 //x2=84.095 //y2=5.155
cc_5417 ( N_SN_M165_noxref_g N_noxref_22_c_9186_n ) capacitor c=0.01736f \
 //x=84.4 //y=6.02 //x2=84.975 //y2=5.155
cc_5418 ( N_SN_c_8150_n N_noxref_22_c_9177_n ) capacitor c=0.00300507f \
 //x=83.99 //y=2.08 //x2=85.84 //y2=2.59
cc_5419 ( N_SN_c_8263_n N_noxref_22_c_9251_n ) capacitor c=0.00426767f \
 //x=84.325 //y=4.79 //x2=84.18 //y2=5.155
cc_5420 ( N_SN_M164_noxref_g N_noxref_22_M164_noxref_d ) capacitor \
 c=0.0180032f //x=83.96 //y=6.02 //x2=84.035 //y2=5.02
cc_5421 ( N_SN_M165_noxref_g N_noxref_22_M164_noxref_d ) capacitor \
 c=0.0180032f //x=84.4 //y=6.02 //x2=84.035 //y2=5.02
cc_5422 ( N_SN_c_8141_n N_noxref_24_c_9433_n ) capacitor c=0.0110334f \
 //x=83.875 //y=2.96 //x2=82.765 //y2=2.22
cc_5423 ( N_SN_c_8141_n N_noxref_24_c_9437_n ) capacitor c=8.83918e-19 \
 //x=83.875 //y=2.96 //x2=81.145 //y2=2.22
cc_5424 ( N_SN_c_8141_n N_noxref_24_c_9440_n ) capacitor c=0.00956254f \
 //x=83.875 //y=2.96 //x2=92.355 //y2=2.22
cc_5425 ( N_SN_c_8150_n N_noxref_24_c_9440_n ) capacitor c=0.0193884f \
 //x=83.99 //y=2.08 //x2=92.355 //y2=2.22
cc_5426 ( N_SN_c_8598_p N_noxref_24_c_9440_n ) capacitor c=0.00583058f \
 //x=84.08 //y=1.915 //x2=92.355 //y2=2.22
cc_5427 ( N_SN_c_8141_n N_noxref_24_c_9446_n ) capacitor c=5.30243e-19 \
 //x=83.875 //y=2.96 //x2=82.995 //y2=2.22
cc_5428 ( N_SN_c_8150_n N_noxref_24_c_9446_n ) capacitor c=0.00151165f \
 //x=83.99 //y=2.08 //x2=82.995 //y2=2.22
cc_5429 ( N_SN_c_8598_p N_noxref_24_c_9446_n ) capacitor c=2.3323e-19 \
 //x=84.08 //y=1.915 //x2=82.995 //y2=2.22
cc_5430 ( N_SN_c_8141_n N_noxref_24_c_9451_n ) capacitor c=0.0210801f \
 //x=83.875 //y=2.96 //x2=81.03 //y2=2.22
cc_5431 ( N_SN_c_8150_n N_noxref_24_c_9451_n ) capacitor c=3.78301e-19 \
 //x=83.99 //y=2.08 //x2=81.03 //y2=2.22
cc_5432 ( N_SN_c_8141_n N_noxref_24_c_9452_n ) capacitor c=0.0234071f \
 //x=83.875 //y=2.96 //x2=82.88 //y2=2.08
cc_5433 ( N_SN_c_8150_n N_noxref_24_c_9452_n ) capacitor c=0.043739f //x=83.99 \
 //y=2.08 //x2=82.88 //y2=2.08
cc_5434 ( N_SN_c_8598_p N_noxref_24_c_9452_n ) capacitor c=0.00201602f \
 //x=84.08 //y=1.915 //x2=82.88 //y2=2.08
cc_5435 ( N_SN_c_8271_n N_noxref_24_c_9452_n ) capacitor c=0.00183762f \
 //x=83.99 //y=4.7 //x2=82.88 //y2=2.08
cc_5436 ( N_SN_M164_noxref_g N_noxref_24_M162_noxref_g ) capacitor \
 c=0.0105869f //x=83.96 //y=6.02 //x2=83.08 //y2=6.02
cc_5437 ( N_SN_M164_noxref_g N_noxref_24_M163_noxref_g ) capacitor c=0.10632f \
 //x=83.96 //y=6.02 //x2=83.52 //y2=6.02
cc_5438 ( N_SN_M165_noxref_g N_noxref_24_M163_noxref_g ) capacitor \
 c=0.0101598f //x=84.4 //y=6.02 //x2=83.52 //y2=6.02
cc_5439 ( N_SN_c_8653_p N_noxref_24_c_9456_n ) capacitor c=5.72482e-19 \
 //x=83.555 //y=0.91 //x2=82.58 //y2=0.875
cc_5440 ( N_SN_c_8653_p N_noxref_24_c_9458_n ) capacitor c=0.00149976f \
 //x=83.555 //y=0.91 //x2=82.58 //y2=1.22
cc_5441 ( N_SN_c_8655_p N_noxref_24_c_9459_n ) capacitor c=0.00111227f \
 //x=83.555 //y=1.22 //x2=82.58 //y2=1.53
cc_5442 ( N_SN_c_8150_n N_noxref_24_c_9460_n ) capacitor c=0.00210802f \
 //x=83.99 //y=2.08 //x2=82.58 //y2=1.915
cc_5443 ( N_SN_c_8598_p N_noxref_24_c_9460_n ) capacitor c=0.00834532f \
 //x=84.08 //y=1.915 //x2=82.58 //y2=1.915
cc_5444 ( N_SN_c_8653_p N_noxref_24_c_9463_n ) capacitor c=0.0160123f \
 //x=83.555 //y=0.91 //x2=83.11 //y2=0.875
cc_5445 ( N_SN_c_8609_p N_noxref_24_c_9463_n ) capacitor c=0.00103227f \
 //x=84.08 //y=0.91 //x2=83.11 //y2=0.875
cc_5446 ( N_SN_c_8655_p N_noxref_24_c_9465_n ) capacitor c=0.0124075f \
 //x=83.555 //y=1.22 //x2=83.11 //y2=1.22
cc_5447 ( N_SN_c_8610_p N_noxref_24_c_9465_n ) capacitor c=0.0010154f \
 //x=84.08 //y=1.22 //x2=83.11 //y2=1.22
cc_5448 ( N_SN_c_8611_p N_noxref_24_c_9465_n ) capacitor c=9.23422e-19 \
 //x=84.08 //y=1.45 //x2=83.11 //y2=1.22
cc_5449 ( N_SN_c_8150_n N_noxref_24_c_9604_n ) capacitor c=0.00147352f \
 //x=83.99 //y=2.08 //x2=83.445 //y2=4.79
cc_5450 ( N_SN_c_8271_n N_noxref_24_c_9604_n ) capacitor c=0.0168581f \
 //x=83.99 //y=4.7 //x2=83.445 //y2=4.79
cc_5451 ( N_SN_c_8150_n N_noxref_24_c_9509_n ) capacitor c=0.00142741f \
 //x=83.99 //y=2.08 //x2=83.155 //y2=4.79
cc_5452 ( N_SN_c_8271_n N_noxref_24_c_9509_n ) capacitor c=0.00484466f \
 //x=83.99 //y=4.7 //x2=83.155 //y2=4.79
cc_5453 ( N_SN_c_8135_n N_noxref_26_c_10048_n ) capacitor c=0.144685f \
 //x=55.015 //y=2.96 //x2=53.905 //y2=3.33
cc_5454 ( N_SN_c_8135_n N_noxref_26_c_10043_n ) capacitor c=0.0292951f \
 //x=55.015 //y=2.96 //x2=52.285 //y2=3.33
cc_5455 ( N_SN_c_8135_n N_noxref_26_c_10050_n ) capacitor c=0.0775856f \
 //x=55.015 //y=2.96 //x2=56.895 //y2=3.33
cc_5456 ( N_SN_c_8138_n N_noxref_26_c_10050_n ) capacitor c=0.158511f \
 //x=69.445 //y=2.96 //x2=56.895 //y2=3.33
cc_5457 ( N_SN_c_8399_n N_noxref_26_c_10050_n ) capacitor c=0.0265806f \
 //x=55.245 //y=2.96 //x2=56.895 //y2=3.33
cc_5458 ( N_SN_c_8148_n N_noxref_26_c_10050_n ) capacitor c=0.0208912f \
 //x=55.13 //y=2.08 //x2=56.895 //y2=3.33
cc_5459 ( N_SN_c_8135_n N_noxref_26_c_10052_n ) capacitor c=0.0265971f \
 //x=55.015 //y=2.96 //x2=54.135 //y2=3.33
cc_5460 ( N_SN_c_8148_n N_noxref_26_c_10052_n ) capacitor c=8.75907e-19 \
 //x=55.13 //y=2.08 //x2=54.135 //y2=3.33
cc_5461 ( N_SN_c_8138_n N_noxref_26_c_9933_n ) capacitor c=0.197778f \
 //x=69.445 //y=2.96 //x2=65.035 //y2=3.7
cc_5462 ( N_SN_c_8138_n N_noxref_26_c_9912_n ) capacitor c=0.00400427f \
 //x=69.445 //y=2.96 //x2=88.315 //y2=4.07
cc_5463 ( N_SN_c_8141_n N_noxref_26_c_9912_n ) capacitor c=0.0329309f \
 //x=83.875 //y=2.96 //x2=88.315 //y2=4.07
cc_5464 ( N_SN_c_8149_n N_noxref_26_c_9912_n ) capacitor c=0.0190126f \
 //x=69.56 //y=2.08 //x2=88.315 //y2=4.07
cc_5465 ( N_SN_c_8150_n N_noxref_26_c_9912_n ) capacitor c=0.0190126f \
 //x=83.99 //y=2.08 //x2=88.315 //y2=4.07
cc_5466 ( N_SN_c_8135_n N_noxref_26_c_9958_n ) capacitor c=0.0206002f \
 //x=55.015 //y=2.96 //x2=52.17 //y2=3.33
cc_5467 ( N_SN_c_8148_n N_noxref_26_c_9958_n ) capacitor c=3.49835e-19 \
 //x=55.13 //y=2.08 //x2=52.17 //y2=3.33
cc_5468 ( N_SN_c_8135_n N_noxref_26_c_9916_n ) capacitor c=0.0216162f \
 //x=55.015 //y=2.96 //x2=54.02 //y2=2.08
cc_5469 ( N_SN_c_8399_n N_noxref_26_c_9916_n ) capacitor c=0.00128547f \
 //x=55.245 //y=2.96 //x2=54.02 //y2=2.08
cc_5470 ( N_SN_c_8148_n N_noxref_26_c_9916_n ) capacitor c=0.0393552f \
 //x=55.13 //y=2.08 //x2=54.02 //y2=2.08
cc_5471 ( N_SN_c_8426_n N_noxref_26_c_9916_n ) capacitor c=0.00203769f \
 //x=55.22 //y=1.915 //x2=54.02 //y2=2.08
cc_5472 ( N_SN_c_8269_n N_noxref_26_c_9916_n ) capacitor c=0.0017365f \
 //x=55.13 //y=4.7 //x2=54.02 //y2=2.08
cc_5473 ( N_SN_M128_noxref_g N_noxref_26_M126_noxref_g ) capacitor \
 c=0.0105174f //x=55.1 //y=6.02 //x2=54.22 //y2=6.02
cc_5474 ( N_SN_M128_noxref_g N_noxref_26_M127_noxref_g ) capacitor c=0.10624f \
 //x=55.1 //y=6.02 //x2=54.66 //y2=6.02
cc_5475 ( N_SN_M129_noxref_g N_noxref_26_M127_noxref_g ) capacitor \
 c=0.0100903f //x=55.54 //y=6.02 //x2=54.66 //y2=6.02
cc_5476 ( N_SN_c_8690_p N_noxref_26_c_9921_n ) capacitor c=5.72482e-19 \
 //x=54.695 //y=0.91 //x2=53.72 //y2=0.875
cc_5477 ( N_SN_c_8690_p N_noxref_26_c_9923_n ) capacitor c=0.00149976f \
 //x=54.695 //y=0.91 //x2=53.72 //y2=1.22
cc_5478 ( N_SN_c_8692_p N_noxref_26_c_9924_n ) capacitor c=0.00111227f \
 //x=54.695 //y=1.22 //x2=53.72 //y2=1.53
cc_5479 ( N_SN_c_8148_n N_noxref_26_c_9925_n ) capacitor c=0.00210802f \
 //x=55.13 //y=2.08 //x2=53.72 //y2=1.915
cc_5480 ( N_SN_c_8426_n N_noxref_26_c_9925_n ) capacitor c=0.00834532f \
 //x=55.22 //y=1.915 //x2=53.72 //y2=1.915
cc_5481 ( N_SN_c_8690_p N_noxref_26_c_9928_n ) capacitor c=0.0160123f \
 //x=54.695 //y=0.91 //x2=54.25 //y2=0.875
cc_5482 ( N_SN_c_8423_n N_noxref_26_c_9928_n ) capacitor c=0.00103227f \
 //x=55.22 //y=0.91 //x2=54.25 //y2=0.875
cc_5483 ( N_SN_c_8692_p N_noxref_26_c_9930_n ) capacitor c=0.0124075f \
 //x=54.695 //y=1.22 //x2=54.25 //y2=1.22
cc_5484 ( N_SN_c_8424_n N_noxref_26_c_9930_n ) capacitor c=0.0010154f \
 //x=55.22 //y=1.22 //x2=54.25 //y2=1.22
cc_5485 ( N_SN_c_8425_n N_noxref_26_c_9930_n ) capacitor c=9.23422e-19 \
 //x=55.22 //y=1.45 //x2=54.25 //y2=1.22
cc_5486 ( N_SN_c_8148_n N_noxref_26_c_10024_n ) capacitor c=0.00120758f \
 //x=55.13 //y=2.08 //x2=54.585 //y2=4.79
cc_5487 ( N_SN_c_8269_n N_noxref_26_c_10024_n ) capacitor c=0.0170104f \
 //x=55.13 //y=4.7 //x2=54.585 //y2=4.79
cc_5488 ( N_SN_c_8148_n N_noxref_26_c_9977_n ) capacitor c=0.00142741f \
 //x=55.13 //y=2.08 //x2=54.295 //y2=4.79
cc_5489 ( N_SN_c_8269_n N_noxref_26_c_9977_n ) capacitor c=0.00484466f \
 //x=55.13 //y=4.7 //x2=54.295 //y2=4.79
cc_5490 ( N_SN_c_8192_n N_noxref_32_c_10751_n ) capacitor c=0.0167228f \
 //x=11.405 //y=0.91 //x2=12.065 //y2=0.54
cc_5491 ( N_SN_c_8197_n N_noxref_32_c_10751_n ) capacitor c=0.00534519f \
 //x=11.93 //y=0.91 //x2=12.065 //y2=0.54
cc_5492 ( N_SN_c_8145_n N_noxref_32_c_10774_n ) capacitor c=0.0117694f \
 //x=11.84 //y=2.08 //x2=12.065 //y2=1.59
cc_5493 ( N_SN_c_8195_n N_noxref_32_c_10774_n ) capacitor c=0.0157358f \
 //x=11.405 //y=1.22 //x2=12.065 //y2=1.59
cc_5494 ( N_SN_c_8200_n N_noxref_32_c_10774_n ) capacitor c=0.021347f \
 //x=11.93 //y=1.915 //x2=12.065 //y2=1.59
cc_5495 ( N_SN_c_8192_n N_noxref_32_M6_noxref_s ) capacitor c=0.00798959f \
 //x=11.405 //y=0.91 //x2=10.075 //y2=0.375
cc_5496 ( N_SN_c_8199_n N_noxref_32_M6_noxref_s ) capacitor c=0.00212176f \
 //x=11.93 //y=1.45 //x2=10.075 //y2=0.375
cc_5497 ( N_SN_c_8200_n N_noxref_32_M6_noxref_s ) capacitor c=0.00298115f \
 //x=11.93 //y=1.915 //x2=10.075 //y2=0.375
cc_5498 ( N_SN_c_8712_p N_noxref_33_c_10793_n ) capacitor c=2.14837e-19 \
 //x=11.775 //y=0.755 //x2=12.635 //y2=0.995
cc_5499 ( N_SN_c_8197_n N_noxref_33_c_10793_n ) capacitor c=0.00123426f \
 //x=11.93 //y=0.91 //x2=12.635 //y2=0.995
cc_5500 ( N_SN_c_8198_n N_noxref_33_c_10793_n ) capacitor c=0.0129288f \
 //x=11.93 //y=1.22 //x2=12.635 //y2=0.995
cc_5501 ( N_SN_c_8199_n N_noxref_33_c_10793_n ) capacitor c=0.00142359f \
 //x=11.93 //y=1.45 //x2=12.635 //y2=0.995
cc_5502 ( N_SN_c_8192_n N_noxref_33_M7_noxref_d ) capacitor c=0.00223875f \
 //x=11.405 //y=0.91 //x2=11.48 //y2=0.91
cc_5503 ( N_SN_c_8195_n N_noxref_33_M7_noxref_d ) capacitor c=0.00262485f \
 //x=11.405 //y=1.22 //x2=11.48 //y2=0.91
cc_5504 ( N_SN_c_8712_p N_noxref_33_M7_noxref_d ) capacitor c=0.00220746f \
 //x=11.775 //y=0.755 //x2=11.48 //y2=0.91
cc_5505 ( N_SN_c_8719_p N_noxref_33_M7_noxref_d ) capacitor c=0.00194798f \
 //x=11.775 //y=1.375 //x2=11.48 //y2=0.91
cc_5506 ( N_SN_c_8197_n N_noxref_33_M7_noxref_d ) capacitor c=0.00198465f \
 //x=11.93 //y=0.91 //x2=11.48 //y2=0.91
cc_5507 ( N_SN_c_8198_n N_noxref_33_M7_noxref_d ) capacitor c=0.00128384f \
 //x=11.93 //y=1.22 //x2=11.48 //y2=0.91
cc_5508 ( N_SN_c_8197_n N_noxref_33_M8_noxref_s ) capacitor c=7.21316e-19 \
 //x=11.93 //y=0.91 //x2=12.585 //y2=0.375
cc_5509 ( N_SN_c_8198_n N_noxref_33_M8_noxref_s ) capacitor c=0.00348171f \
 //x=11.93 //y=1.22 //x2=12.585 //y2=0.375
cc_5510 ( N_SN_c_8249_n N_noxref_38_c_11058_n ) capacitor c=0.0167228f \
 //x=25.835 //y=0.91 //x2=26.495 //y2=0.54
cc_5511 ( N_SN_c_8254_n N_noxref_38_c_11058_n ) capacitor c=0.00534519f \
 //x=26.36 //y=0.91 //x2=26.495 //y2=0.54
cc_5512 ( N_SN_c_8146_n N_noxref_38_c_11081_n ) capacitor c=0.0117694f \
 //x=26.27 //y=2.08 //x2=26.495 //y2=1.59
cc_5513 ( N_SN_c_8252_n N_noxref_38_c_11081_n ) capacitor c=0.0157358f \
 //x=25.835 //y=1.22 //x2=26.495 //y2=1.59
cc_5514 ( N_SN_c_8257_n N_noxref_38_c_11081_n ) capacitor c=0.021347f \
 //x=26.36 //y=1.915 //x2=26.495 //y2=1.59
cc_5515 ( N_SN_c_8249_n N_noxref_38_M15_noxref_s ) capacitor c=0.00798959f \
 //x=25.835 //y=0.91 //x2=24.505 //y2=0.375
cc_5516 ( N_SN_c_8256_n N_noxref_38_M15_noxref_s ) capacitor c=0.00212176f \
 //x=26.36 //y=1.45 //x2=24.505 //y2=0.375
cc_5517 ( N_SN_c_8257_n N_noxref_38_M15_noxref_s ) capacitor c=0.00298115f \
 //x=26.36 //y=1.915 //x2=24.505 //y2=0.375
cc_5518 ( N_SN_c_8732_p N_noxref_39_c_11100_n ) capacitor c=2.14837e-19 \
 //x=26.205 //y=0.755 //x2=27.065 //y2=0.995
cc_5519 ( N_SN_c_8254_n N_noxref_39_c_11100_n ) capacitor c=0.00123426f \
 //x=26.36 //y=0.91 //x2=27.065 //y2=0.995
cc_5520 ( N_SN_c_8255_n N_noxref_39_c_11100_n ) capacitor c=0.0129288f \
 //x=26.36 //y=1.22 //x2=27.065 //y2=0.995
cc_5521 ( N_SN_c_8256_n N_noxref_39_c_11100_n ) capacitor c=0.00142359f \
 //x=26.36 //y=1.45 //x2=27.065 //y2=0.995
cc_5522 ( N_SN_c_8249_n N_noxref_39_M16_noxref_d ) capacitor c=0.00223875f \
 //x=25.835 //y=0.91 //x2=25.91 //y2=0.91
cc_5523 ( N_SN_c_8252_n N_noxref_39_M16_noxref_d ) capacitor c=0.00262485f \
 //x=25.835 //y=1.22 //x2=25.91 //y2=0.91
cc_5524 ( N_SN_c_8732_p N_noxref_39_M16_noxref_d ) capacitor c=0.00220746f \
 //x=26.205 //y=0.755 //x2=25.91 //y2=0.91
cc_5525 ( N_SN_c_8739_p N_noxref_39_M16_noxref_d ) capacitor c=0.00194798f \
 //x=26.205 //y=1.375 //x2=25.91 //y2=0.91
cc_5526 ( N_SN_c_8254_n N_noxref_39_M16_noxref_d ) capacitor c=0.00198465f \
 //x=26.36 //y=0.91 //x2=25.91 //y2=0.91
cc_5527 ( N_SN_c_8255_n N_noxref_39_M16_noxref_d ) capacitor c=0.00128384f \
 //x=26.36 //y=1.22 //x2=25.91 //y2=0.91
cc_5528 ( N_SN_c_8254_n N_noxref_39_M17_noxref_s ) capacitor c=7.21316e-19 \
 //x=26.36 //y=0.91 //x2=27.015 //y2=0.375
cc_5529 ( N_SN_c_8255_n N_noxref_39_M17_noxref_s ) capacitor c=0.00348171f \
 //x=26.36 //y=1.22 //x2=27.015 //y2=0.375
cc_5530 ( N_SN_c_8349_n N_noxref_44_c_11364_n ) capacitor c=0.0167228f \
 //x=40.265 //y=0.91 //x2=40.925 //y2=0.54
cc_5531 ( N_SN_c_8354_n N_noxref_44_c_11364_n ) capacitor c=0.00534519f \
 //x=40.79 //y=0.91 //x2=40.925 //y2=0.54
cc_5532 ( N_SN_c_8147_n N_noxref_44_c_11387_n ) capacitor c=0.0117694f \
 //x=40.7 //y=2.08 //x2=40.925 //y2=1.59
cc_5533 ( N_SN_c_8352_n N_noxref_44_c_11387_n ) capacitor c=0.0157358f \
 //x=40.265 //y=1.22 //x2=40.925 //y2=1.59
cc_5534 ( N_SN_c_8357_n N_noxref_44_c_11387_n ) capacitor c=0.021347f \
 //x=40.79 //y=1.915 //x2=40.925 //y2=1.59
cc_5535 ( N_SN_c_8349_n N_noxref_44_M24_noxref_s ) capacitor c=0.00798959f \
 //x=40.265 //y=0.91 //x2=38.935 //y2=0.375
cc_5536 ( N_SN_c_8356_n N_noxref_44_M24_noxref_s ) capacitor c=0.00212176f \
 //x=40.79 //y=1.45 //x2=38.935 //y2=0.375
cc_5537 ( N_SN_c_8357_n N_noxref_44_M24_noxref_s ) capacitor c=0.00298115f \
 //x=40.79 //y=1.915 //x2=38.935 //y2=0.375
cc_5538 ( N_SN_c_8752_p N_noxref_45_c_11406_n ) capacitor c=2.14837e-19 \
 //x=40.635 //y=0.755 //x2=41.495 //y2=0.995
cc_5539 ( N_SN_c_8354_n N_noxref_45_c_11406_n ) capacitor c=0.00123426f \
 //x=40.79 //y=0.91 //x2=41.495 //y2=0.995
cc_5540 ( N_SN_c_8355_n N_noxref_45_c_11406_n ) capacitor c=0.0129288f \
 //x=40.79 //y=1.22 //x2=41.495 //y2=0.995
cc_5541 ( N_SN_c_8356_n N_noxref_45_c_11406_n ) capacitor c=0.00142359f \
 //x=40.79 //y=1.45 //x2=41.495 //y2=0.995
cc_5542 ( N_SN_c_8349_n N_noxref_45_M25_noxref_d ) capacitor c=0.00223875f \
 //x=40.265 //y=0.91 //x2=40.34 //y2=0.91
cc_5543 ( N_SN_c_8352_n N_noxref_45_M25_noxref_d ) capacitor c=0.00262485f \
 //x=40.265 //y=1.22 //x2=40.34 //y2=0.91
cc_5544 ( N_SN_c_8752_p N_noxref_45_M25_noxref_d ) capacitor c=0.00220746f \
 //x=40.635 //y=0.755 //x2=40.34 //y2=0.91
cc_5545 ( N_SN_c_8759_p N_noxref_45_M25_noxref_d ) capacitor c=0.00194798f \
 //x=40.635 //y=1.375 //x2=40.34 //y2=0.91
cc_5546 ( N_SN_c_8354_n N_noxref_45_M25_noxref_d ) capacitor c=0.00198465f \
 //x=40.79 //y=0.91 //x2=40.34 //y2=0.91
cc_5547 ( N_SN_c_8355_n N_noxref_45_M25_noxref_d ) capacitor c=0.00128384f \
 //x=40.79 //y=1.22 //x2=40.34 //y2=0.91
cc_5548 ( N_SN_c_8354_n N_noxref_45_M26_noxref_s ) capacitor c=7.21316e-19 \
 //x=40.79 //y=0.91 //x2=41.445 //y2=0.375
cc_5549 ( N_SN_c_8355_n N_noxref_45_M26_noxref_s ) capacitor c=0.00348171f \
 //x=40.79 //y=1.22 //x2=41.445 //y2=0.375
cc_5550 ( N_SN_c_8690_p N_noxref_50_c_11671_n ) capacitor c=0.0167228f \
 //x=54.695 //y=0.91 //x2=55.355 //y2=0.54
cc_5551 ( N_SN_c_8423_n N_noxref_50_c_11671_n ) capacitor c=0.00534519f \
 //x=55.22 //y=0.91 //x2=55.355 //y2=0.54
cc_5552 ( N_SN_c_8148_n N_noxref_50_c_11682_n ) capacitor c=0.0117694f \
 //x=55.13 //y=2.08 //x2=55.355 //y2=1.59
cc_5553 ( N_SN_c_8692_p N_noxref_50_c_11682_n ) capacitor c=0.0157358f \
 //x=54.695 //y=1.22 //x2=55.355 //y2=1.59
cc_5554 ( N_SN_c_8426_n N_noxref_50_c_11682_n ) capacitor c=0.021347f \
 //x=55.22 //y=1.915 //x2=55.355 //y2=1.59
cc_5555 ( N_SN_c_8690_p N_noxref_50_M33_noxref_s ) capacitor c=0.00798959f \
 //x=54.695 //y=0.91 //x2=53.365 //y2=0.375
cc_5556 ( N_SN_c_8425_n N_noxref_50_M33_noxref_s ) capacitor c=0.00212176f \
 //x=55.22 //y=1.45 //x2=53.365 //y2=0.375
cc_5557 ( N_SN_c_8426_n N_noxref_50_M33_noxref_s ) capacitor c=0.00298115f \
 //x=55.22 //y=1.915 //x2=53.365 //y2=0.375
cc_5558 ( N_SN_c_8772_p N_noxref_51_c_11713_n ) capacitor c=2.14837e-19 \
 //x=55.065 //y=0.755 //x2=55.925 //y2=0.995
cc_5559 ( N_SN_c_8423_n N_noxref_51_c_11713_n ) capacitor c=0.00123426f \
 //x=55.22 //y=0.91 //x2=55.925 //y2=0.995
cc_5560 ( N_SN_c_8424_n N_noxref_51_c_11713_n ) capacitor c=0.0129288f \
 //x=55.22 //y=1.22 //x2=55.925 //y2=0.995
cc_5561 ( N_SN_c_8425_n N_noxref_51_c_11713_n ) capacitor c=0.00142359f \
 //x=55.22 //y=1.45 //x2=55.925 //y2=0.995
cc_5562 ( N_SN_c_8690_p N_noxref_51_M34_noxref_d ) capacitor c=0.00223875f \
 //x=54.695 //y=0.91 //x2=54.77 //y2=0.91
cc_5563 ( N_SN_c_8692_p N_noxref_51_M34_noxref_d ) capacitor c=0.00262485f \
 //x=54.695 //y=1.22 //x2=54.77 //y2=0.91
cc_5564 ( N_SN_c_8772_p N_noxref_51_M34_noxref_d ) capacitor c=0.00220746f \
 //x=55.065 //y=0.755 //x2=54.77 //y2=0.91
cc_5565 ( N_SN_c_8779_p N_noxref_51_M34_noxref_d ) capacitor c=0.00194798f \
 //x=55.065 //y=1.375 //x2=54.77 //y2=0.91
cc_5566 ( N_SN_c_8423_n N_noxref_51_M34_noxref_d ) capacitor c=0.00198465f \
 //x=55.22 //y=0.91 //x2=54.77 //y2=0.91
cc_5567 ( N_SN_c_8424_n N_noxref_51_M34_noxref_d ) capacitor c=0.00128384f \
 //x=55.22 //y=1.22 //x2=54.77 //y2=0.91
cc_5568 ( N_SN_c_8423_n N_noxref_51_M35_noxref_s ) capacitor c=7.21316e-19 \
 //x=55.22 //y=0.91 //x2=55.875 //y2=0.375
cc_5569 ( N_SN_c_8424_n N_noxref_51_M35_noxref_s ) capacitor c=0.00348171f \
 //x=55.22 //y=1.22 //x2=55.875 //y2=0.375
cc_5570 ( N_SN_c_8477_n N_noxref_56_c_11977_n ) capacitor c=0.0167228f \
 //x=69.125 //y=0.91 //x2=69.785 //y2=0.54
cc_5571 ( N_SN_c_8482_n N_noxref_56_c_11977_n ) capacitor c=0.00534519f \
 //x=69.65 //y=0.91 //x2=69.785 //y2=0.54
cc_5572 ( N_SN_c_8149_n N_noxref_56_c_12000_n ) capacitor c=0.0117694f \
 //x=69.56 //y=2.08 //x2=69.785 //y2=1.59
cc_5573 ( N_SN_c_8480_n N_noxref_56_c_12000_n ) capacitor c=0.0157358f \
 //x=69.125 //y=1.22 //x2=69.785 //y2=1.59
cc_5574 ( N_SN_c_8485_n N_noxref_56_c_12000_n ) capacitor c=0.021347f \
 //x=69.65 //y=1.915 //x2=69.785 //y2=1.59
cc_5575 ( N_SN_c_8477_n N_noxref_56_M42_noxref_s ) capacitor c=0.00798959f \
 //x=69.125 //y=0.91 //x2=67.795 //y2=0.375
cc_5576 ( N_SN_c_8484_n N_noxref_56_M42_noxref_s ) capacitor c=0.00212176f \
 //x=69.65 //y=1.45 //x2=67.795 //y2=0.375
cc_5577 ( N_SN_c_8485_n N_noxref_56_M42_noxref_s ) capacitor c=0.00298115f \
 //x=69.65 //y=1.915 //x2=67.795 //y2=0.375
cc_5578 ( N_SN_c_8792_p N_noxref_57_c_12019_n ) capacitor c=2.14837e-19 \
 //x=69.495 //y=0.755 //x2=70.355 //y2=0.995
cc_5579 ( N_SN_c_8482_n N_noxref_57_c_12019_n ) capacitor c=0.00123426f \
 //x=69.65 //y=0.91 //x2=70.355 //y2=0.995
cc_5580 ( N_SN_c_8483_n N_noxref_57_c_12019_n ) capacitor c=0.0129288f \
 //x=69.65 //y=1.22 //x2=70.355 //y2=0.995
cc_5581 ( N_SN_c_8484_n N_noxref_57_c_12019_n ) capacitor c=0.00142359f \
 //x=69.65 //y=1.45 //x2=70.355 //y2=0.995
cc_5582 ( N_SN_c_8477_n N_noxref_57_M43_noxref_d ) capacitor c=0.00223875f \
 //x=69.125 //y=0.91 //x2=69.2 //y2=0.91
cc_5583 ( N_SN_c_8480_n N_noxref_57_M43_noxref_d ) capacitor c=0.00262485f \
 //x=69.125 //y=1.22 //x2=69.2 //y2=0.91
cc_5584 ( N_SN_c_8792_p N_noxref_57_M43_noxref_d ) capacitor c=0.00220746f \
 //x=69.495 //y=0.755 //x2=69.2 //y2=0.91
cc_5585 ( N_SN_c_8799_p N_noxref_57_M43_noxref_d ) capacitor c=0.00194798f \
 //x=69.495 //y=1.375 //x2=69.2 //y2=0.91
cc_5586 ( N_SN_c_8482_n N_noxref_57_M43_noxref_d ) capacitor c=0.00198465f \
 //x=69.65 //y=0.91 //x2=69.2 //y2=0.91
cc_5587 ( N_SN_c_8483_n N_noxref_57_M43_noxref_d ) capacitor c=0.00128384f \
 //x=69.65 //y=1.22 //x2=69.2 //y2=0.91
cc_5588 ( N_SN_c_8482_n N_noxref_57_M44_noxref_s ) capacitor c=7.21316e-19 \
 //x=69.65 //y=0.91 //x2=70.305 //y2=0.375
cc_5589 ( N_SN_c_8483_n N_noxref_57_M44_noxref_s ) capacitor c=0.00348171f \
 //x=69.65 //y=1.22 //x2=70.305 //y2=0.375
cc_5590 ( N_SN_c_8141_n N_noxref_60_c_12202_n ) capacitor c=0.00152987f \
 //x=83.875 //y=2.96 //x2=79.405 //y2=1.59
cc_5591 ( N_SN_c_8141_n N_noxref_60_M48_noxref_s ) capacitor c=0.00302917f \
 //x=83.875 //y=2.96 //x2=77.415 //y2=0.375
cc_5592 ( N_SN_c_8141_n N_noxref_61_c_12224_n ) capacitor c=0.00383675f \
 //x=83.875 //y=2.96 //x2=79.975 //y2=0.995
cc_5593 ( N_SN_c_8141_n N_noxref_61_M50_noxref_s ) capacitor c=0.00324882f \
 //x=83.875 //y=2.96 //x2=79.925 //y2=0.375
cc_5594 ( N_SN_c_8653_p N_noxref_62_c_12285_n ) capacitor c=0.0167228f \
 //x=83.555 //y=0.91 //x2=84.215 //y2=0.54
cc_5595 ( N_SN_c_8609_p N_noxref_62_c_12285_n ) capacitor c=0.00534519f \
 //x=84.08 //y=0.91 //x2=84.215 //y2=0.54
cc_5596 ( N_SN_c_8150_n N_noxref_62_c_12295_n ) capacitor c=0.0117694f \
 //x=83.99 //y=2.08 //x2=84.215 //y2=1.59
cc_5597 ( N_SN_c_8655_p N_noxref_62_c_12295_n ) capacitor c=0.0157358f \
 //x=83.555 //y=1.22 //x2=84.215 //y2=1.59
cc_5598 ( N_SN_c_8598_p N_noxref_62_c_12295_n ) capacitor c=0.021347f \
 //x=84.08 //y=1.915 //x2=84.215 //y2=1.59
cc_5599 ( N_SN_c_8653_p N_noxref_62_M51_noxref_s ) capacitor c=0.00798959f \
 //x=83.555 //y=0.91 //x2=82.225 //y2=0.375
cc_5600 ( N_SN_c_8611_p N_noxref_62_M51_noxref_s ) capacitor c=0.00212176f \
 //x=84.08 //y=1.45 //x2=82.225 //y2=0.375
cc_5601 ( N_SN_c_8598_p N_noxref_62_M51_noxref_s ) capacitor c=0.00298115f \
 //x=84.08 //y=1.915 //x2=82.225 //y2=0.375
cc_5602 ( N_SN_c_8816_p N_noxref_63_c_12329_n ) capacitor c=2.14837e-19 \
 //x=83.925 //y=0.755 //x2=84.785 //y2=0.995
cc_5603 ( N_SN_c_8609_p N_noxref_63_c_12329_n ) capacitor c=0.00123426f \
 //x=84.08 //y=0.91 //x2=84.785 //y2=0.995
cc_5604 ( N_SN_c_8610_p N_noxref_63_c_12329_n ) capacitor c=0.0129288f \
 //x=84.08 //y=1.22 //x2=84.785 //y2=0.995
cc_5605 ( N_SN_c_8611_p N_noxref_63_c_12329_n ) capacitor c=0.00142359f \
 //x=84.08 //y=1.45 //x2=84.785 //y2=0.995
cc_5606 ( N_SN_c_8653_p N_noxref_63_M52_noxref_d ) capacitor c=0.00223875f \
 //x=83.555 //y=0.91 //x2=83.63 //y2=0.91
cc_5607 ( N_SN_c_8655_p N_noxref_63_M52_noxref_d ) capacitor c=0.00262485f \
 //x=83.555 //y=1.22 //x2=83.63 //y2=0.91
cc_5608 ( N_SN_c_8816_p N_noxref_63_M52_noxref_d ) capacitor c=0.00220746f \
 //x=83.925 //y=0.755 //x2=83.63 //y2=0.91
cc_5609 ( N_SN_c_8823_p N_noxref_63_M52_noxref_d ) capacitor c=0.00194798f \
 //x=83.925 //y=1.375 //x2=83.63 //y2=0.91
cc_5610 ( N_SN_c_8609_p N_noxref_63_M52_noxref_d ) capacitor c=0.00198465f \
 //x=84.08 //y=0.91 //x2=83.63 //y2=0.91
cc_5611 ( N_SN_c_8610_p N_noxref_63_M52_noxref_d ) capacitor c=0.00128384f \
 //x=84.08 //y=1.22 //x2=83.63 //y2=0.91
cc_5612 ( N_SN_c_8609_p N_noxref_63_M53_noxref_s ) capacitor c=7.21316e-19 \
 //x=84.08 //y=0.91 //x2=84.735 //y2=0.375
cc_5613 ( N_SN_c_8610_p N_noxref_63_M53_noxref_s ) capacitor c=0.00348171f \
 //x=84.08 //y=1.22 //x2=84.735 //y2=0.375
cc_5614 ( N_noxref_21_c_8880_n N_noxref_22_c_9171_n ) capacitor c=0.04877f \
 //x=84.985 //y=3.7 //x2=85.725 //y2=2.59
cc_5615 ( N_noxref_21_c_8831_n N_noxref_22_c_9171_n ) capacitor c=0.0237087f \
 //x=85.1 //y=2.08 //x2=85.725 //y2=2.59
cc_5616 ( N_noxref_21_c_8880_n N_noxref_22_c_9174_n ) capacitor c=6.53213e-19 \
 //x=84.985 //y=3.7 //x2=80.405 //y2=2.59
cc_5617 ( N_noxref_21_c_8880_n N_noxref_22_c_9175_n ) capacitor c=0.0203405f \
 //x=84.985 //y=3.7 //x2=80.29 //y2=2.08
cc_5618 ( N_noxref_21_M166_noxref_g N_noxref_22_c_9186_n ) capacitor \
 c=0.01736f //x=84.84 //y=6.02 //x2=84.975 //y2=5.155
cc_5619 ( N_noxref_21_M167_noxref_g N_noxref_22_c_9190_n ) capacitor \
 c=0.0194981f //x=85.28 //y=6.02 //x2=85.755 //y2=5.155
cc_5620 ( N_noxref_21_c_8897_n N_noxref_22_c_9190_n ) capacitor c=0.00201851f \
 //x=85.1 //y=4.7 //x2=85.755 //y2=5.155
cc_5621 ( N_noxref_21_c_9094_p N_noxref_22_c_9176_n ) capacitor c=0.00371277f \
 //x=85.465 //y=1.415 //x2=85.755 //y2=1.665
cc_5622 ( N_noxref_21_c_9095_p N_noxref_22_c_9176_n ) capacitor c=0.00457401f \
 //x=85.62 //y=1.26 //x2=85.755 //y2=1.665
cc_5623 ( N_noxref_21_c_8880_n N_noxref_22_c_9177_n ) capacitor c=0.00735597f \
 //x=84.985 //y=3.7 //x2=85.84 //y2=2.59
cc_5624 ( N_noxref_21_c_8831_n N_noxref_22_c_9177_n ) capacitor c=0.0805664f \
 //x=85.1 //y=2.08 //x2=85.84 //y2=2.59
cc_5625 ( N_noxref_21_c_9081_n N_noxref_22_c_9177_n ) capacitor c=0.00709342f \
 //x=85.1 //y=2.08 //x2=85.84 //y2=2.59
cc_5626 ( N_noxref_21_c_9083_n N_noxref_22_c_9177_n ) capacitor c=0.00283672f \
 //x=85.1 //y=1.915 //x2=85.84 //y2=2.59
cc_5627 ( N_noxref_21_c_8897_n N_noxref_22_c_9177_n ) capacitor c=0.013693f \
 //x=85.1 //y=4.7 //x2=85.84 //y2=2.59
cc_5628 ( N_noxref_21_c_8831_n N_noxref_22_c_9268_n ) capacitor c=0.016476f \
 //x=85.1 //y=2.08 //x2=85.06 //y2=5.155
cc_5629 ( N_noxref_21_c_8897_n N_noxref_22_c_9268_n ) capacitor c=0.00475601f \
 //x=85.1 //y=4.7 //x2=85.06 //y2=5.155
cc_5630 ( N_noxref_21_c_9072_n N_noxref_22_M53_noxref_d ) capacitor \
 c=0.00217566f //x=85.09 //y=0.915 //x2=85.165 //y2=0.915
cc_5631 ( N_noxref_21_c_9073_n N_noxref_22_M53_noxref_d ) capacitor \
 c=0.0034598f //x=85.09 //y=1.26 //x2=85.165 //y2=0.915
cc_5632 ( N_noxref_21_c_9074_n N_noxref_22_M53_noxref_d ) capacitor \
 c=0.00546784f //x=85.09 //y=1.57 //x2=85.165 //y2=0.915
cc_5633 ( N_noxref_21_c_9106_p N_noxref_22_M53_noxref_d ) capacitor \
 c=0.00241102f //x=85.465 //y=0.76 //x2=85.165 //y2=0.915
cc_5634 ( N_noxref_21_c_9094_p N_noxref_22_M53_noxref_d ) capacitor \
 c=0.0138621f //x=85.465 //y=1.415 //x2=85.165 //y2=0.915
cc_5635 ( N_noxref_21_c_9108_p N_noxref_22_M53_noxref_d ) capacitor \
 c=0.00219619f //x=85.62 //y=0.915 //x2=85.165 //y2=0.915
cc_5636 ( N_noxref_21_c_9095_p N_noxref_22_M53_noxref_d ) capacitor \
 c=0.00603828f //x=85.62 //y=1.26 //x2=85.165 //y2=0.915
cc_5637 ( N_noxref_21_c_9083_n N_noxref_22_M53_noxref_d ) capacitor \
 c=0.00661782f //x=85.1 //y=1.915 //x2=85.165 //y2=0.915
cc_5638 ( N_noxref_21_M166_noxref_g N_noxref_22_M166_noxref_d ) capacitor \
 c=0.0180032f //x=84.84 //y=6.02 //x2=84.915 //y2=5.02
cc_5639 ( N_noxref_21_M167_noxref_g N_noxref_22_M166_noxref_d ) capacitor \
 c=0.0194246f //x=85.28 //y=6.02 //x2=84.915 //y2=5.02
cc_5640 ( N_noxref_21_c_8880_n N_noxref_24_c_9440_n ) capacitor c=0.00651954f \
 //x=84.985 //y=3.7 //x2=92.355 //y2=2.22
cc_5641 ( N_noxref_21_c_8831_n N_noxref_24_c_9440_n ) capacitor c=0.0186201f \
 //x=85.1 //y=2.08 //x2=92.355 //y2=2.22
cc_5642 ( N_noxref_21_c_9094_p N_noxref_24_c_9440_n ) capacitor c=3.13485e-19 \
 //x=85.465 //y=1.415 //x2=92.355 //y2=2.22
cc_5643 ( N_noxref_21_c_9081_n N_noxref_24_c_9440_n ) capacitor c=0.00584491f \
 //x=85.1 //y=2.08 //x2=92.355 //y2=2.22
cc_5644 ( N_noxref_21_c_8845_n N_noxref_24_c_9482_n ) capacitor c=3.10026e-19 \
 //x=76.135 //y=5.155 //x2=78.575 //y2=5.155
cc_5645 ( N_noxref_21_c_8880_n N_noxref_24_c_9451_n ) capacitor c=0.0211098f \
 //x=84.985 //y=3.7 //x2=81.03 //y2=2.22
cc_5646 ( N_noxref_21_c_8880_n N_noxref_24_c_9452_n ) capacitor c=0.0221279f \
 //x=84.985 //y=3.7 //x2=82.88 //y2=2.08
cc_5647 ( N_noxref_21_c_8831_n N_noxref_24_c_9452_n ) capacitor c=0.00118806f \
 //x=85.1 //y=2.08 //x2=82.88 //y2=2.08
cc_5648 ( N_noxref_21_c_8935_n N_noxref_26_c_9933_n ) capacitor c=0.0158317f \
 //x=65.975 //y=3.7 //x2=65.035 //y2=3.7
cc_5649 ( N_noxref_21_c_8828_n N_noxref_26_c_9933_n ) capacitor c=0.00222024f \
 //x=65.86 //y=2.08 //x2=65.035 //y2=3.7
cc_5650 ( N_noxref_21_c_8935_n N_noxref_26_c_10119_n ) capacitor c=0.00147396f \
 //x=65.975 //y=3.7 //x2=65.12 //y2=3.985
cc_5651 ( N_noxref_21_c_8828_n N_noxref_26_c_10119_n ) capacitor c=0.00494521f \
 //x=65.86 //y=2.08 //x2=65.12 //y2=3.985
cc_5652 ( N_noxref_21_c_8898_n N_noxref_26_c_9912_n ) capacitor c=0.403974f \
 //x=70.555 //y=3.7 //x2=88.315 //y2=4.07
cc_5653 ( N_noxref_21_c_8935_n N_noxref_26_c_9912_n ) capacitor c=0.0292842f \
 //x=65.975 //y=3.7 //x2=88.315 //y2=4.07
cc_5654 ( N_noxref_21_c_8878_n N_noxref_26_c_9912_n ) capacitor c=0.468094f \
 //x=76.105 //y=3.7 //x2=88.315 //y2=4.07
cc_5655 ( N_noxref_21_c_8905_n N_noxref_26_c_9912_n ) capacitor c=0.026596f \
 //x=70.785 //y=3.7 //x2=88.315 //y2=4.07
cc_5656 ( N_noxref_21_c_8880_n N_noxref_26_c_9912_n ) capacitor c=0.792602f \
 //x=84.985 //y=3.7 //x2=88.315 //y2=4.07
cc_5657 ( N_noxref_21_c_8881_n N_noxref_26_c_9912_n ) capacitor c=0.026809f \
 //x=76.335 //y=3.7 //x2=88.315 //y2=4.07
cc_5658 ( N_noxref_21_c_8828_n N_noxref_26_c_9912_n ) capacitor c=0.0197551f \
 //x=65.86 //y=2.08 //x2=88.315 //y2=4.07
cc_5659 ( N_noxref_21_c_8829_n N_noxref_26_c_9912_n ) capacitor c=0.0198068f \
 //x=70.67 //y=2.08 //x2=88.315 //y2=4.07
cc_5660 ( N_noxref_21_c_8849_n N_noxref_26_c_9912_n ) capacitor c=0.0200135f \
 //x=76.22 //y=3.7 //x2=88.315 //y2=4.07
cc_5661 ( N_noxref_21_c_8831_n N_noxref_26_c_9912_n ) capacitor c=0.0198068f \
 //x=85.1 //y=2.08 //x2=88.315 //y2=4.07
cc_5662 ( N_noxref_21_c_8828_n N_noxref_55_c_11923_n ) capacitor c=0.00204385f \
 //x=65.86 //y=2.08 //x2=66.515 //y2=0.54
cc_5663 ( N_noxref_21_c_8955_n N_noxref_55_c_11923_n ) capacitor c=0.0194423f \
 //x=65.85 //y=0.915 //x2=66.515 //y2=0.54
cc_5664 ( N_noxref_21_c_8997_n N_noxref_55_c_11923_n ) capacitor c=0.00656458f \
 //x=66.38 //y=0.915 //x2=66.515 //y2=0.54
cc_5665 ( N_noxref_21_c_8958_n N_noxref_55_c_11923_n ) capacitor c=2.20712e-19 \
 //x=65.86 //y=2.08 //x2=66.515 //y2=0.54
cc_5666 ( N_noxref_21_c_8956_n N_noxref_55_c_11945_n ) capacitor c=0.00538829f \
 //x=65.85 //y=1.26 //x2=65.63 //y2=0.995
cc_5667 ( N_noxref_21_c_8955_n N_noxref_55_M41_noxref_s ) capacitor \
 c=0.00538829f //x=65.85 //y=0.915 //x2=65.495 //y2=0.375
cc_5668 ( N_noxref_21_c_8957_n N_noxref_55_M41_noxref_s ) capacitor \
 c=0.00538829f //x=65.85 //y=1.57 //x2=65.495 //y2=0.375
cc_5669 ( N_noxref_21_c_8997_n N_noxref_55_M41_noxref_s ) capacitor \
 c=0.0143002f //x=66.38 //y=0.915 //x2=65.495 //y2=0.375
cc_5670 ( N_noxref_21_c_8998_n N_noxref_55_M41_noxref_s ) capacitor \
 c=0.00290153f //x=66.38 //y=1.26 //x2=65.495 //y2=0.375
cc_5671 ( N_noxref_21_c_8829_n N_noxref_57_c_12024_n ) capacitor c=0.00204385f \
 //x=70.67 //y=2.08 //x2=71.325 //y2=0.54
cc_5672 ( N_noxref_21_c_8918_n N_noxref_57_c_12024_n ) capacitor c=0.0194423f \
 //x=70.66 //y=0.915 //x2=71.325 //y2=0.54
cc_5673 ( N_noxref_21_c_8924_n N_noxref_57_c_12024_n ) capacitor c=0.00656458f \
 //x=71.19 //y=0.915 //x2=71.325 //y2=0.54
cc_5674 ( N_noxref_21_c_8927_n N_noxref_57_c_12024_n ) capacitor c=2.20712e-19 \
 //x=70.67 //y=2.08 //x2=71.325 //y2=0.54
cc_5675 ( N_noxref_21_c_8919_n N_noxref_57_c_12034_n ) capacitor c=0.00538829f \
 //x=70.66 //y=1.26 //x2=70.44 //y2=0.995
cc_5676 ( N_noxref_21_c_8918_n N_noxref_57_M44_noxref_s ) capacitor \
 c=0.00538829f //x=70.66 //y=0.915 //x2=70.305 //y2=0.375
cc_5677 ( N_noxref_21_c_8920_n N_noxref_57_M44_noxref_s ) capacitor \
 c=0.00538829f //x=70.66 //y=1.57 //x2=70.305 //y2=0.375
cc_5678 ( N_noxref_21_c_8924_n N_noxref_57_M44_noxref_s ) capacitor \
 c=0.0143002f //x=71.19 //y=0.915 //x2=70.305 //y2=0.375
cc_5679 ( N_noxref_21_c_8925_n N_noxref_57_M44_noxref_s ) capacitor \
 c=0.00290153f //x=71.19 //y=1.26 //x2=70.305 //y2=0.375
cc_5680 ( N_noxref_21_M47_noxref_d N_noxref_58_M45_noxref_s ) capacitor \
 c=0.00309936f //x=75.545 //y=0.915 //x2=72.605 //y2=0.375
cc_5681 ( N_noxref_21_c_8830_n N_noxref_59_c_12125_n ) capacitor c=0.00457167f \
 //x=76.135 //y=1.665 //x2=76.135 //y2=0.54
cc_5682 ( N_noxref_21_M47_noxref_d N_noxref_59_c_12125_n ) capacitor \
 c=0.0115903f //x=75.545 //y=0.915 //x2=76.135 //y2=0.54
cc_5683 ( N_noxref_21_c_9017_n N_noxref_59_c_12152_n ) capacitor c=0.0200405f \
 //x=75.82 //y=1.665 //x2=75.25 //y2=0.995
cc_5684 ( N_noxref_21_M47_noxref_d N_noxref_59_M46_noxref_d ) capacitor \
 c=5.27807e-19 //x=75.545 //y=0.915 //x2=74.01 //y2=0.91
cc_5685 ( N_noxref_21_c_8830_n N_noxref_59_M47_noxref_s ) capacitor \
 c=0.0196084f //x=76.135 //y=1.665 //x2=75.115 //y2=0.375
cc_5686 ( N_noxref_21_M47_noxref_d N_noxref_59_M47_noxref_s ) capacitor \
 c=0.0426368f //x=75.545 //y=0.915 //x2=75.115 //y2=0.375
cc_5687 ( N_noxref_21_c_8830_n N_noxref_60_c_12188_n ) capacitor c=3.84569e-19 \
 //x=76.135 //y=1.665 //x2=77.55 //y2=1.505
cc_5688 ( N_noxref_21_M47_noxref_d N_noxref_60_M48_noxref_s ) capacitor \
 c=2.55333e-19 //x=75.545 //y=0.915 //x2=77.415 //y2=0.375
cc_5689 ( N_noxref_21_c_8831_n N_noxref_63_c_12334_n ) capacitor c=0.00204385f \
 //x=85.1 //y=2.08 //x2=85.755 //y2=0.54
cc_5690 ( N_noxref_21_c_9072_n N_noxref_63_c_12334_n ) capacitor c=0.0194423f \
 //x=85.09 //y=0.915 //x2=85.755 //y2=0.54
cc_5691 ( N_noxref_21_c_9108_p N_noxref_63_c_12334_n ) capacitor c=0.00656458f \
 //x=85.62 //y=0.915 //x2=85.755 //y2=0.54
cc_5692 ( N_noxref_21_c_9081_n N_noxref_63_c_12334_n ) capacitor c=2.20712e-19 \
 //x=85.1 //y=2.08 //x2=85.755 //y2=0.54
cc_5693 ( N_noxref_21_c_9073_n N_noxref_63_c_12358_n ) capacitor c=0.00538829f \
 //x=85.09 //y=1.26 //x2=84.87 //y2=0.995
cc_5694 ( N_noxref_21_c_9072_n N_noxref_63_M53_noxref_s ) capacitor \
 c=0.00538829f //x=85.09 //y=0.915 //x2=84.735 //y2=0.375
cc_5695 ( N_noxref_21_c_9074_n N_noxref_63_M53_noxref_s ) capacitor \
 c=0.00538829f //x=85.09 //y=1.57 //x2=84.735 //y2=0.375
cc_5696 ( N_noxref_21_c_9108_p N_noxref_63_M53_noxref_s ) capacitor \
 c=0.0143002f //x=85.62 //y=0.915 //x2=84.735 //y2=0.375
cc_5697 ( N_noxref_21_c_9095_p N_noxref_63_M53_noxref_s ) capacitor \
 c=0.00290153f //x=85.62 //y=1.26 //x2=84.735 //y2=0.375
cc_5698 ( N_noxref_22_c_9171_n N_noxref_24_c_9433_n ) capacitor c=0.14348f \
 //x=85.725 //y=2.59 //x2=82.765 //y2=2.22
cc_5699 ( N_noxref_22_c_9171_n N_noxref_24_c_9437_n ) capacitor c=0.029328f \
 //x=85.725 //y=2.59 //x2=81.145 //y2=2.22
cc_5700 ( N_noxref_22_c_9175_n N_noxref_24_c_9437_n ) capacitor c=0.00397358f \
 //x=80.29 //y=2.08 //x2=81.145 //y2=2.22
cc_5701 ( N_noxref_22_c_9235_n N_noxref_24_c_9437_n ) capacitor c=0.00289405f \
 //x=80.29 //y=2.08 //x2=81.145 //y2=2.22
cc_5702 ( N_noxref_22_c_9171_n N_noxref_24_c_9440_n ) capacitor c=0.264813f \
 //x=85.725 //y=2.59 //x2=92.355 //y2=2.22
cc_5703 ( N_noxref_22_c_9285_p N_noxref_24_c_9440_n ) capacitor c=0.016327f \
 //x=85.44 //y=1.665 //x2=92.355 //y2=2.22
cc_5704 ( N_noxref_22_c_9177_n N_noxref_24_c_9440_n ) capacitor c=0.0215653f \
 //x=85.84 //y=2.59 //x2=92.355 //y2=2.22
cc_5705 ( N_noxref_22_c_9171_n N_noxref_24_c_9446_n ) capacitor c=0.0267441f \
 //x=85.725 //y=2.59 //x2=82.995 //y2=2.22
cc_5706 ( N_noxref_22_M160_noxref_g N_noxref_24_c_9484_n ) capacitor \
 c=0.01736f //x=80.03 //y=6.02 //x2=80.165 //y2=5.155
cc_5707 ( N_noxref_22_c_9184_n N_noxref_24_c_9488_n ) capacitor c=3.10026e-19 \
 //x=83.385 //y=5.155 //x2=80.945 //y2=5.155
cc_5708 ( N_noxref_22_M161_noxref_g N_noxref_24_c_9488_n ) capacitor \
 c=0.0194981f //x=80.47 //y=6.02 //x2=80.945 //y2=5.155
cc_5709 ( N_noxref_22_c_9222_n N_noxref_24_c_9488_n ) capacitor c=0.00201851f \
 //x=80.29 //y=4.7 //x2=80.945 //y2=5.155
cc_5710 ( N_noxref_22_c_9292_p N_noxref_24_c_9450_n ) capacitor c=0.00359704f \
 //x=80.655 //y=1.415 //x2=80.945 //y2=1.665
cc_5711 ( N_noxref_22_c_9293_p N_noxref_24_c_9450_n ) capacitor c=0.00457401f \
 //x=80.81 //y=1.26 //x2=80.945 //y2=1.665
cc_5712 ( N_noxref_22_c_9171_n N_noxref_24_c_9630_n ) capacitor c=0.0102157f \
 //x=85.725 //y=2.59 //x2=80.63 //y2=1.665
cc_5713 ( N_noxref_22_c_9171_n N_noxref_24_c_9451_n ) capacitor c=0.0184272f \
 //x=85.725 //y=2.59 //x2=81.03 //y2=2.22
cc_5714 ( N_noxref_22_c_9174_n N_noxref_24_c_9451_n ) capacitor c=0.00179385f \
 //x=80.405 //y=2.59 //x2=81.03 //y2=2.22
cc_5715 ( N_noxref_22_c_9175_n N_noxref_24_c_9451_n ) capacitor c=0.0785134f \
 //x=80.29 //y=2.08 //x2=81.03 //y2=2.22
cc_5716 ( N_noxref_22_c_9235_n N_noxref_24_c_9451_n ) capacitor c=0.00768602f \
 //x=80.29 //y=2.08 //x2=81.03 //y2=2.22
cc_5717 ( N_noxref_22_c_9238_n N_noxref_24_c_9451_n ) capacitor c=0.00283672f \
 //x=80.29 //y=1.915 //x2=81.03 //y2=2.22
cc_5718 ( N_noxref_22_c_9222_n N_noxref_24_c_9451_n ) capacitor c=0.013844f \
 //x=80.29 //y=4.7 //x2=81.03 //y2=2.22
cc_5719 ( N_noxref_22_c_9171_n N_noxref_24_c_9452_n ) capacitor c=0.0206666f \
 //x=85.725 //y=2.59 //x2=82.88 //y2=2.08
cc_5720 ( N_noxref_22_c_9175_n N_noxref_24_c_9452_n ) capacitor c=6.57608e-19 \
 //x=80.29 //y=2.08 //x2=82.88 //y2=2.08
cc_5721 ( N_noxref_22_c_9175_n N_noxref_24_c_9639_n ) capacitor c=0.0166016f \
 //x=80.29 //y=2.08 //x2=80.25 //y2=5.155
cc_5722 ( N_noxref_22_c_9222_n N_noxref_24_c_9639_n ) capacitor c=0.00475601f \
 //x=80.29 //y=4.7 //x2=80.25 //y2=5.155
cc_5723 ( N_noxref_22_c_9184_n N_noxref_24_M162_noxref_g ) capacitor \
 c=0.0213876f //x=83.385 //y=5.155 //x2=83.08 //y2=6.02
cc_5724 ( N_noxref_22_c_9180_n N_noxref_24_M163_noxref_g ) capacitor \
 c=0.0168349f //x=84.095 //y=5.155 //x2=83.52 //y2=6.02
cc_5725 ( N_noxref_22_M162_noxref_d N_noxref_24_M163_noxref_g ) capacitor \
 c=0.0180032f //x=83.155 //y=5.02 //x2=83.52 //y2=6.02
cc_5726 ( N_noxref_22_c_9184_n N_noxref_24_c_9604_n ) capacitor c=0.00428486f \
 //x=83.385 //y=5.155 //x2=83.445 //y2=4.79
cc_5727 ( N_noxref_22_c_9232_n N_noxref_24_M50_noxref_d ) capacitor \
 c=0.00217566f //x=80.28 //y=0.915 //x2=80.355 //y2=0.915
cc_5728 ( N_noxref_22_c_9233_n N_noxref_24_M50_noxref_d ) capacitor \
 c=0.0034598f //x=80.28 //y=1.26 //x2=80.355 //y2=0.915
cc_5729 ( N_noxref_22_c_9234_n N_noxref_24_M50_noxref_d ) capacitor \
 c=0.00544291f //x=80.28 //y=1.57 //x2=80.355 //y2=0.915
cc_5730 ( N_noxref_22_c_9312_p N_noxref_24_M50_noxref_d ) capacitor \
 c=0.00241102f //x=80.655 //y=0.76 //x2=80.355 //y2=0.915
cc_5731 ( N_noxref_22_c_9292_p N_noxref_24_M50_noxref_d ) capacitor \
 c=0.0140297f //x=80.655 //y=1.415 //x2=80.355 //y2=0.915
cc_5732 ( N_noxref_22_c_9314_p N_noxref_24_M50_noxref_d ) capacitor \
 c=0.00219619f //x=80.81 //y=0.915 //x2=80.355 //y2=0.915
cc_5733 ( N_noxref_22_c_9293_p N_noxref_24_M50_noxref_d ) capacitor \
 c=0.00603828f //x=80.81 //y=1.26 //x2=80.355 //y2=0.915
cc_5734 ( N_noxref_22_c_9238_n N_noxref_24_M50_noxref_d ) capacitor \
 c=0.00661782f //x=80.29 //y=1.915 //x2=80.355 //y2=0.915
cc_5735 ( N_noxref_22_M160_noxref_g N_noxref_24_M160_noxref_d ) capacitor \
 c=0.0180032f //x=80.03 //y=6.02 //x2=80.105 //y2=5.02
cc_5736 ( N_noxref_22_M161_noxref_g N_noxref_24_M160_noxref_d ) capacitor \
 c=0.0194246f //x=80.47 //y=6.02 //x2=80.105 //y2=5.02
cc_5737 ( N_noxref_22_c_9171_n N_noxref_26_c_9912_n ) capacitor c=0.0217211f \
 //x=85.725 //y=2.59 //x2=88.315 //y2=4.07
cc_5738 ( N_noxref_22_c_9175_n N_noxref_26_c_9912_n ) capacitor c=0.0179722f \
 //x=80.29 //y=2.08 //x2=88.315 //y2=4.07
cc_5739 ( N_noxref_22_c_9177_n N_noxref_26_c_9912_n ) capacitor c=0.0228844f \
 //x=85.84 //y=2.59 //x2=88.315 //y2=4.07
cc_5740 ( N_noxref_22_c_9177_n N_noxref_26_c_9917_n ) capacitor c=7.99399e-19 \
 //x=85.84 //y=2.59 //x2=88.43 //y2=2.08
cc_5741 ( N_noxref_22_c_9171_n N_noxref_61_c_12229_n ) capacitor c=4.77662e-19 \
 //x=85.725 //y=2.59 //x2=80.945 //y2=0.54
cc_5742 ( N_noxref_22_c_9174_n N_noxref_61_c_12229_n ) capacitor c=3.67738e-19 \
 //x=80.405 //y=2.59 //x2=80.945 //y2=0.54
cc_5743 ( N_noxref_22_c_9175_n N_noxref_61_c_12229_n ) capacitor c=0.00206286f \
 //x=80.29 //y=2.08 //x2=80.945 //y2=0.54
cc_5744 ( N_noxref_22_c_9232_n N_noxref_61_c_12229_n ) capacitor c=0.0194423f \
 //x=80.28 //y=0.915 //x2=80.945 //y2=0.54
cc_5745 ( N_noxref_22_c_9314_p N_noxref_61_c_12229_n ) capacitor c=0.00656458f \
 //x=80.81 //y=0.915 //x2=80.945 //y2=0.54
cc_5746 ( N_noxref_22_c_9235_n N_noxref_61_c_12229_n ) capacitor c=2.20712e-19 \
 //x=80.29 //y=2.08 //x2=80.945 //y2=0.54
cc_5747 ( N_noxref_22_c_9233_n N_noxref_61_c_12257_n ) capacitor c=0.00538829f \
 //x=80.28 //y=1.26 //x2=80.06 //y2=0.995
cc_5748 ( N_noxref_22_c_9232_n N_noxref_61_M50_noxref_s ) capacitor \
 c=0.00538829f //x=80.28 //y=0.915 //x2=79.925 //y2=0.375
cc_5749 ( N_noxref_22_c_9234_n N_noxref_61_M50_noxref_s ) capacitor \
 c=0.00538829f //x=80.28 //y=1.57 //x2=79.925 //y2=0.375
cc_5750 ( N_noxref_22_c_9314_p N_noxref_61_M50_noxref_s ) capacitor \
 c=0.0143002f //x=80.81 //y=0.915 //x2=79.925 //y2=0.375
cc_5751 ( N_noxref_22_c_9293_p N_noxref_61_M50_noxref_s ) capacitor \
 c=0.00290153f //x=80.81 //y=1.26 //x2=79.925 //y2=0.375
cc_5752 ( N_noxref_22_M53_noxref_d N_noxref_62_M51_noxref_s ) capacitor \
 c=0.00309936f //x=85.165 //y=0.915 //x2=82.225 //y2=0.375
cc_5753 ( N_noxref_22_c_9176_n N_noxref_63_c_12334_n ) capacitor c=0.00457167f \
 //x=85.755 //y=1.665 //x2=85.755 //y2=0.54
cc_5754 ( N_noxref_22_M53_noxref_d N_noxref_63_c_12334_n ) capacitor \
 c=0.0115903f //x=85.165 //y=0.915 //x2=85.755 //y2=0.54
cc_5755 ( N_noxref_22_c_9285_p N_noxref_63_c_12358_n ) capacitor c=0.020048f \
 //x=85.44 //y=1.665 //x2=84.87 //y2=0.995
cc_5756 ( N_noxref_22_M53_noxref_d N_noxref_63_M52_noxref_d ) capacitor \
 c=5.27807e-19 //x=85.165 //y=0.915 //x2=83.63 //y2=0.91
cc_5757 ( N_noxref_22_c_9176_n N_noxref_63_M53_noxref_s ) capacitor \
 c=0.0184051f //x=85.755 //y=1.665 //x2=84.735 //y2=0.375
cc_5758 ( N_noxref_22_M53_noxref_d N_noxref_63_M53_noxref_s ) capacitor \
 c=0.0426134f //x=85.165 //y=0.915 //x2=84.735 //y2=0.375
cc_5759 ( N_noxref_22_c_9176_n N_noxref_64_c_12399_n ) capacitor c=3.04182e-19 \
 //x=85.755 //y=1.665 //x2=87.275 //y2=1.495
cc_5760 ( N_noxref_23_M175_noxref_d N_noxref_24_c_9453_n ) capacitor \
 c=0.00511793f //x=92.305 //y=5.025 //x2=92.5 //y2=2.08
cc_5761 ( N_noxref_23_c_9395_p N_noxref_24_M174_noxref_g ) capacitor \
 c=0.0150104f //x=92.365 //y=6.91 //x2=91.79 //y2=6.025
cc_5762 ( N_noxref_23_M173_noxref_d N_noxref_24_M174_noxref_g ) capacitor \
 c=0.0130327f //x=91.425 //y=5.025 //x2=91.79 //y2=6.025
cc_5763 ( N_noxref_23_c_9395_p N_noxref_24_M175_noxref_g ) capacitor \
 c=0.0155183f //x=92.365 //y=6.91 //x2=92.23 //y2=6.025
cc_5764 ( N_noxref_23_M175_noxref_d N_noxref_24_M175_noxref_g ) capacitor \
 c=0.0398886f //x=92.305 //y=5.025 //x2=92.23 //y2=6.025
cc_5765 ( N_noxref_23_M175_noxref_d N_noxref_24_c_9511_n ) capacitor \
 c=0.00411435f //x=92.305 //y=5.025 //x2=92.23 //y2=4.87
cc_5766 ( N_noxref_23_c_9395_p N_noxref_25_c_9823_n ) capacitor c=0.00546043f \
 //x=92.365 //y=6.91 //x2=93.915 //y2=5.21
cc_5767 ( N_noxref_23_M175_noxref_d N_noxref_25_c_9823_n ) capacitor \
 c=0.00675852f //x=92.305 //y=5.025 //x2=93.915 //y2=5.21
cc_5768 ( N_noxref_23_c_9342_n N_noxref_25_c_9827_n ) capacitor c=0.0086908f \
 //x=90.575 //y=5.21 //x2=92.125 //y2=5.21
cc_5769 ( N_noxref_23_c_9395_p N_noxref_25_c_9827_n ) capacitor c=9.39989e-19 \
 //x=92.365 //y=6.91 //x2=92.125 //y2=5.21
cc_5770 ( N_noxref_23_c_9388_n N_noxref_25_c_9838_n ) capacitor c=0.00102709f \
 //x=91.485 //y=6.91 //x2=91.925 //y2=5.21
cc_5771 ( N_noxref_23_c_9395_p N_noxref_25_c_9838_n ) capacitor c=9.89472e-19 \
 //x=92.365 //y=6.91 //x2=91.925 //y2=5.21
cc_5772 ( N_noxref_23_M173_noxref_d N_noxref_25_c_9838_n ) capacitor \
 c=0.0124612f //x=91.425 //y=5.025 //x2=91.925 //y2=5.21
cc_5773 ( N_noxref_23_c_9342_n N_noxref_25_c_9829_n ) capacitor c=0.00638395f \
 //x=90.575 //y=5.21 //x2=91.215 //y2=5.21
cc_5774 ( N_noxref_23_c_9362_n N_noxref_25_c_9829_n ) capacitor c=0.0682565f \
 //x=90.69 //y=5.21 //x2=91.215 //y2=5.21
cc_5775 ( N_noxref_23_c_9362_n N_noxref_25_c_9830_n ) capacitor c=9.46973e-19 \
 //x=90.69 //y=5.21 //x2=92.01 //y2=5.295
cc_5776 ( N_noxref_23_M175_noxref_d N_noxref_25_c_9831_n ) capacitor \
 c=0.001104f //x=92.305 //y=5.025 //x2=94.03 //y2=5.21
cc_5777 ( N_noxref_23_c_9395_p N_noxref_25_c_9833_n ) capacitor c=0.001104f \
 //x=92.365 //y=6.91 //x2=94.115 //y2=6.91
cc_5778 ( N_noxref_23_c_9342_n N_noxref_25_M172_noxref_d ) capacitor \
 c=4.76678e-19 //x=90.575 //y=5.21 //x2=90.985 //y2=5.025
cc_5779 ( N_noxref_23_c_9388_n N_noxref_25_M172_noxref_d ) capacitor \
 c=0.0115421f //x=91.485 //y=6.91 //x2=90.985 //y2=5.025
cc_5780 ( N_noxref_23_M173_noxref_d N_noxref_25_M172_noxref_d ) capacitor \
 c=0.0458293f //x=91.425 //y=5.025 //x2=90.985 //y2=5.025
cc_5781 ( N_noxref_23_M175_noxref_d N_noxref_25_M172_noxref_d ) capacitor \
 c=7.47391e-19 //x=92.305 //y=5.025 //x2=90.985 //y2=5.025
cc_5782 ( N_noxref_23_c_9362_n N_noxref_25_M174_noxref_d ) capacitor \
 c=9.55e-19 //x=90.69 //y=5.21 //x2=91.865 //y2=5.025
cc_5783 ( N_noxref_23_c_9395_p N_noxref_25_M174_noxref_d ) capacitor \
 c=0.0115693f //x=92.365 //y=6.91 //x2=91.865 //y2=5.025
cc_5784 ( N_noxref_23_M173_noxref_d N_noxref_25_M174_noxref_d ) capacitor \
 c=0.0458293f //x=91.425 //y=5.025 //x2=91.865 //y2=5.025
cc_5785 ( N_noxref_23_M175_noxref_d N_noxref_25_M174_noxref_d ) capacitor \
 c=0.0550393f //x=92.305 //y=5.025 //x2=91.865 //y2=5.025
cc_5786 ( N_noxref_23_c_9342_n N_noxref_26_c_9913_n ) capacitor c=0.00923886f \
 //x=90.575 //y=5.21 //x2=94.975 //y2=4.07
cc_5787 ( N_noxref_23_c_9348_n N_noxref_26_c_9913_n ) capacitor c=0.00122833f \
 //x=88.805 //y=5.21 //x2=94.975 //y2=4.07
cc_5788 ( N_noxref_23_c_9353_n N_noxref_26_c_9962_n ) capacitor c=0.012748f \
 //x=88.605 //y=5.21 //x2=88.43 //y2=4.54
cc_5789 ( N_noxref_23_c_9348_n N_noxref_26_M170_noxref_g ) capacitor \
 c=0.0010118f //x=88.805 //y=5.21 //x2=88.47 //y2=6.025
cc_5790 ( N_noxref_23_c_9353_n N_noxref_26_M170_noxref_g ) capacitor \
 c=0.0161605f //x=88.605 //y=5.21 //x2=88.47 //y2=6.025
cc_5791 ( N_noxref_23_c_9359_n N_noxref_26_M170_noxref_g ) capacitor \
 c=0.00226657f //x=88.69 //y=5.295 //x2=88.47 //y2=6.025
cc_5792 ( N_noxref_23_M170_noxref_d N_noxref_26_M170_noxref_g ) capacitor \
 c=0.016914f //x=88.545 //y=5.025 //x2=88.47 //y2=6.025
cc_5793 ( N_noxref_23_c_9342_n N_noxref_26_M171_noxref_g ) capacitor \
 c=0.0104371f //x=90.575 //y=5.21 //x2=88.91 //y2=6.025
cc_5794 ( N_noxref_23_c_9348_n N_noxref_26_M171_noxref_g ) capacitor \
 c=8.30848e-19 //x=88.805 //y=5.21 //x2=88.91 //y2=6.025
cc_5795 ( N_noxref_23_c_9359_n N_noxref_26_M171_noxref_g ) capacitor \
 c=0.0197448f //x=88.69 //y=5.295 //x2=88.91 //y2=6.025
cc_5796 ( N_noxref_23_c_9359_n N_noxref_26_c_9979_n ) capacitor c=0.00458101f \
 //x=88.69 //y=5.295 //x2=88.835 //y2=4.795
cc_5797 ( N_noxref_23_c_9353_n N_noxref_26_c_9980_n ) capacitor c=0.00307538f \
 //x=88.605 //y=5.21 //x2=88.47 //y2=4.705
cc_5798 ( N_noxref_23_c_9362_n N_noxref_65_c_12455_n ) capacitor c=0.00104325f \
 //x=90.69 //y=5.21 //x2=90.605 //y2=1.495
cc_5799 ( N_noxref_24_c_9440_n N_noxref_25_c_9823_n ) capacitor c=5.84148e-19 \
 //x=92.355 //y=2.22 //x2=93.915 //y2=5.21
cc_5800 ( N_noxref_24_c_9448_n N_noxref_25_c_9823_n ) capacitor c=5.85064e-19 \
 //x=93.865 //y=2.08 //x2=93.915 //y2=5.21
cc_5801 ( N_noxref_24_c_9453_n N_noxref_25_c_9823_n ) capacitor c=0.00419026f \
 //x=92.5 //y=2.08 //x2=93.915 //y2=5.21
cc_5802 ( N_noxref_24_c_9455_n N_noxref_25_c_9823_n ) capacitor c=0.0031527f \
 //x=93.98 //y=2.08 //x2=93.915 //y2=5.21
cc_5803 ( N_noxref_24_M175_noxref_g N_noxref_25_c_9823_n ) capacitor \
 c=0.0109874f //x=92.23 //y=6.025 //x2=93.915 //y2=5.21
cc_5804 ( N_noxref_24_M176_noxref_g N_noxref_25_c_9823_n ) capacitor \
 c=0.00645933f //x=94.25 //y=6.025 //x2=93.915 //y2=5.21
cc_5805 ( N_noxref_24_c_9511_n N_noxref_25_c_9823_n ) capacitor c=0.00270424f \
 //x=92.23 //y=4.87 //x2=93.915 //y2=5.21
cc_5806 ( N_noxref_24_c_9512_n N_noxref_25_c_9823_n ) capacitor c=0.00176728f \
 //x=94.325 //y=4.795 //x2=93.915 //y2=5.21
cc_5807 ( N_noxref_24_c_9440_n N_noxref_25_c_9827_n ) capacitor c=2.38143e-19 \
 //x=92.355 //y=2.22 //x2=92.125 //y2=5.21
cc_5808 ( N_noxref_24_M174_noxref_g N_noxref_25_c_9827_n ) capacitor \
 c=6.87102e-19 //x=91.79 //y=6.025 //x2=92.125 //y2=5.21
cc_5809 ( N_noxref_24_M175_noxref_g N_noxref_25_c_9827_n ) capacitor \
 c=8.33934e-19 //x=92.23 //y=6.025 //x2=92.125 //y2=5.21
cc_5810 ( N_noxref_24_M174_noxref_g N_noxref_25_c_9838_n ) capacitor \
 c=0.0179287f //x=91.79 //y=6.025 //x2=91.925 //y2=5.21
cc_5811 ( N_noxref_24_M174_noxref_g N_noxref_25_c_9830_n ) capacitor \
 c=0.0019882f //x=91.79 //y=6.025 //x2=92.01 //y2=5.295
cc_5812 ( N_noxref_24_M175_noxref_g N_noxref_25_c_9830_n ) capacitor \
 c=0.0159381f //x=92.23 //y=6.025 //x2=92.01 //y2=5.295
cc_5813 ( N_noxref_24_c_9675_p N_noxref_25_c_9830_n ) capacitor c=0.00456817f \
 //x=92.155 //y=4.795 //x2=92.01 //y2=5.295
cc_5814 ( N_noxref_24_c_9455_n N_noxref_25_c_9831_n ) capacitor c=0.0184695f \
 //x=93.98 //y=2.08 //x2=94.03 //y2=5.21
cc_5815 ( N_noxref_24_M176_noxref_g N_noxref_25_c_9831_n ) capacitor \
 c=0.0484795f //x=94.25 //y=6.025 //x2=94.03 //y2=5.21
cc_5816 ( N_noxref_24_c_9512_n N_noxref_25_c_9831_n ) capacitor c=0.0078825f \
 //x=94.325 //y=4.795 //x2=94.03 //y2=5.21
cc_5817 ( N_noxref_24_M176_noxref_g N_noxref_25_c_9882_n ) capacitor \
 c=0.0164606f //x=94.25 //y=6.025 //x2=94.825 //y2=6.91
cc_5818 ( N_noxref_24_M177_noxref_g N_noxref_25_c_9882_n ) capacitor \
 c=0.0150104f //x=94.69 //y=6.025 //x2=94.825 //y2=6.91
cc_5819 ( N_noxref_24_M174_noxref_g N_noxref_25_M174_noxref_d ) capacitor \
 c=0.0129738f //x=91.79 //y=6.025 //x2=91.865 //y2=5.025
cc_5820 ( N_noxref_24_M177_noxref_g N_noxref_25_M177_noxref_d ) capacitor \
 c=0.0130327f //x=94.69 //y=6.025 //x2=94.765 //y2=5.025
cc_5821 ( N_noxref_24_c_9440_n N_noxref_26_c_9912_n ) capacitor c=0.0437933f \
 //x=92.355 //y=2.22 //x2=88.315 //y2=4.07
cc_5822 ( N_noxref_24_c_9451_n N_noxref_26_c_9912_n ) capacitor c=0.0181982f \
 //x=81.03 //y=2.22 //x2=88.315 //y2=4.07
cc_5823 ( N_noxref_24_c_9452_n N_noxref_26_c_9912_n ) capacitor c=0.019517f \
 //x=82.88 //y=2.08 //x2=88.315 //y2=4.07
cc_5824 ( N_noxref_24_c_9440_n N_noxref_26_c_9913_n ) capacitor c=0.0716681f \
 //x=92.355 //y=2.22 //x2=94.975 //y2=4.07
cc_5825 ( N_noxref_24_c_9448_n N_noxref_26_c_9913_n ) capacitor c=0.0238267f \
 //x=93.865 //y=2.08 //x2=94.975 //y2=4.07
cc_5826 ( N_noxref_24_c_9453_n N_noxref_26_c_9913_n ) capacitor c=0.0276725f \
 //x=92.5 //y=2.08 //x2=94.975 //y2=4.07
cc_5827 ( N_noxref_24_c_9455_n N_noxref_26_c_9913_n ) capacitor c=0.0282853f \
 //x=93.98 //y=2.08 //x2=94.975 //y2=4.07
cc_5828 ( N_noxref_24_c_9555_n N_noxref_26_c_9913_n ) capacitor c=0.00791694f \
 //x=91.865 //y=4.795 //x2=94.975 //y2=4.07
cc_5829 ( N_noxref_24_c_9511_n N_noxref_26_c_9913_n ) capacitor c=0.0014567f \
 //x=92.23 //y=4.87 //x2=94.975 //y2=4.07
cc_5830 ( N_noxref_24_c_9512_n N_noxref_26_c_9913_n ) capacitor c=0.0117386f \
 //x=94.325 //y=4.795 //x2=94.975 //y2=4.07
cc_5831 ( N_noxref_24_c_9440_n N_noxref_26_c_9943_n ) capacitor c=0.00342879f \
 //x=92.355 //y=2.22 //x2=88.545 //y2=4.07
cc_5832 ( N_noxref_24_c_9440_n N_noxref_26_c_9917_n ) capacitor c=0.0250901f \
 //x=92.355 //y=2.22 //x2=88.43 //y2=2.08
cc_5833 ( N_noxref_24_c_9448_n N_noxref_26_c_9919_n ) capacitor c=0.00669222f \
 //x=93.865 //y=2.08 //x2=95.09 //y2=2.08
cc_5834 ( N_noxref_24_c_9453_n N_noxref_26_c_9919_n ) capacitor c=6.01206e-19 \
 //x=92.5 //y=2.08 //x2=95.09 //y2=2.08
cc_5835 ( N_noxref_24_c_9455_n N_noxref_26_c_9919_n ) capacitor c=0.0539835f \
 //x=93.98 //y=2.08 //x2=95.09 //y2=2.08
cc_5836 ( N_noxref_24_c_9476_n N_noxref_26_c_9919_n ) capacitor c=0.00218919f \
 //x=93.98 //y=2.08 //x2=95.09 //y2=2.08
cc_5837 ( N_noxref_24_c_9699_p N_noxref_26_c_10237_n ) capacitor c=0.00168516f \
 //x=94.615 //y=4.795 //x2=95.11 //y2=4.705
cc_5838 ( N_noxref_24_c_9512_n N_noxref_26_c_10237_n ) capacitor c=0.00143876f \
 //x=94.325 //y=4.795 //x2=95.11 //y2=4.705
cc_5839 ( N_noxref_24_M176_noxref_g N_noxref_26_M178_noxref_g ) capacitor \
 c=0.00932631f //x=94.25 //y=6.025 //x2=95.13 //y2=6.025
cc_5840 ( N_noxref_24_M177_noxref_g N_noxref_26_M178_noxref_g ) capacitor \
 c=0.110179f //x=94.69 //y=6.025 //x2=95.13 //y2=6.025
cc_5841 ( N_noxref_24_M177_noxref_g N_noxref_26_M179_noxref_g ) capacitor \
 c=0.00876656f //x=94.69 //y=6.025 //x2=95.57 //y2=6.025
cc_5842 ( N_noxref_24_c_9440_n N_noxref_26_c_10242_n ) capacitor c=0.0026659f \
 //x=92.355 //y=2.22 //x2=88.84 //y2=1.405
cc_5843 ( N_noxref_24_c_9467_n N_noxref_26_c_10243_n ) capacitor c=4.86506e-19 \
 //x=94.155 //y=0.865 //x2=95.125 //y2=0.905
cc_5844 ( N_noxref_24_c_9469_n N_noxref_26_c_10243_n ) capacitor c=0.00101233f \
 //x=94.155 //y=1.21 //x2=95.125 //y2=0.905
cc_5845 ( N_noxref_24_c_9473_n N_noxref_26_c_10243_n ) capacitor c=0.0161138f \
 //x=94.685 //y=0.865 //x2=95.125 //y2=0.905
cc_5846 ( N_noxref_24_c_9475_n N_noxref_26_c_10246_n ) capacitor c=0.0120728f \
 //x=94.685 //y=1.21 //x2=95.125 //y2=1.255
cc_5847 ( N_noxref_24_c_9709_p N_noxref_26_c_10247_n ) capacitor c=0.00257836f \
 //x=94.155 //y=1.52 //x2=95.125 //y2=1.56
cc_5848 ( N_noxref_24_c_9470_n N_noxref_26_c_10247_n ) capacitor c=0.00662747f \
 //x=94.155 //y=1.915 //x2=95.125 //y2=1.56
cc_5849 ( N_noxref_24_c_9475_n N_noxref_26_c_10247_n ) capacitor c=0.00862358f \
 //x=94.685 //y=1.21 //x2=95.125 //y2=1.56
cc_5850 ( N_noxref_24_c_9475_n N_noxref_26_c_10250_n ) capacitor c=4.4593e-19 \
 //x=94.685 //y=1.21 //x2=95.5 //y2=1.405
cc_5851 ( N_noxref_24_c_9473_n N_noxref_26_c_10251_n ) capacitor c=0.00130607f \
 //x=94.685 //y=0.865 //x2=95.655 //y2=0.905
cc_5852 ( N_noxref_24_c_9475_n N_noxref_26_c_10252_n ) capacitor c=0.00111855f \
 //x=94.685 //y=1.21 //x2=95.655 //y2=1.255
cc_5853 ( N_noxref_24_c_9440_n N_noxref_26_c_9931_n ) capacitor c=0.00615545f \
 //x=92.355 //y=2.22 //x2=88.43 //y2=2.08
cc_5854 ( N_noxref_24_c_9448_n N_noxref_26_c_10254_n ) capacitor c=0.00341891f \
 //x=93.865 //y=2.08 //x2=95.09 //y2=2.08
cc_5855 ( N_noxref_24_c_9455_n N_noxref_26_c_10254_n ) capacitor c=0.00207994f \
 //x=93.98 //y=2.08 //x2=95.09 //y2=2.08
cc_5856 ( N_noxref_24_c_9476_n N_noxref_26_c_10254_n ) capacitor c=0.00908973f \
 //x=93.98 //y=2.08 //x2=95.09 //y2=2.08
cc_5857 ( N_noxref_24_c_9455_n N_noxref_26_c_10257_n ) capacitor c=0.00196222f \
 //x=93.98 //y=2.08 //x2=95.11 //y2=4.705
cc_5858 ( N_noxref_24_c_9699_p N_noxref_26_c_10257_n ) capacitor c=0.0225854f \
 //x=94.615 //y=4.795 //x2=95.11 //y2=4.705
cc_5859 ( N_noxref_24_c_9512_n N_noxref_26_c_10257_n ) capacitor c=0.00469886f \
 //x=94.325 //y=4.795 //x2=95.11 //y2=4.705
cc_5860 ( N_noxref_24_c_9440_n N_Q_c_10368_n ) capacitor c=0.0874774f \
 //x=92.355 //y=2.22 //x2=91.945 //y2=1.18
cc_5861 ( N_noxref_24_c_9550_n N_Q_c_10368_n ) capacitor c=5.17481e-19 \
 //x=91.795 //y=0.905 //x2=91.945 //y2=1.18
cc_5862 ( N_noxref_24_c_9553_n N_Q_c_10368_n ) capacitor c=0.00560566f \
 //x=91.795 //y=1.25 //x2=91.945 //y2=1.18
cc_5863 ( N_noxref_24_c_9440_n N_Q_c_10375_n ) capacitor c=0.00876802f \
 //x=92.355 //y=2.22 //x2=88.845 //y2=1.18
cc_5864 ( N_noxref_24_c_9440_n N_Q_c_10376_n ) capacitor c=0.0053658f \
 //x=92.355 //y=2.22 //x2=95.275 //y2=1.18
cc_5865 ( N_noxref_24_c_9448_n N_Q_c_10376_n ) capacitor c=0.053129f \
 //x=93.865 //y=2.08 //x2=95.275 //y2=1.18
cc_5866 ( N_noxref_24_c_9449_n N_Q_c_10376_n ) capacitor c=0.0103746f //x=92.5 \
 //y=2.08 //x2=95.275 //y2=1.18
cc_5867 ( N_noxref_24_c_9453_n N_Q_c_10376_n ) capacitor c=0.00189559f \
 //x=92.5 //y=2.08 //x2=95.275 //y2=1.18
cc_5868 ( N_noxref_24_c_9455_n N_Q_c_10376_n ) capacitor c=0.00134607f \
 //x=93.98 //y=2.08 //x2=95.275 //y2=1.18
cc_5869 ( N_noxref_24_c_9559_n N_Q_c_10376_n ) capacitor c=4.67724e-19 \
 //x=92.325 //y=0.905 //x2=95.275 //y2=1.18
cc_5870 ( N_noxref_24_c_9560_n N_Q_c_10376_n ) capacitor c=0.00591245f \
 //x=92.325 //y=1.25 //x2=95.275 //y2=1.18
cc_5871 ( N_noxref_24_c_9561_n N_Q_c_10376_n ) capacitor c=0.00282482f \
 //x=92.325 //y=1.56 //x2=95.275 //y2=1.18
cc_5872 ( N_noxref_24_c_9466_n N_Q_c_10376_n ) capacitor c=2.04565e-19 \
 //x=92.325 //y=1.915 //x2=95.275 //y2=1.18
cc_5873 ( N_noxref_24_c_9469_n N_Q_c_10376_n ) capacitor c=0.00500281f \
 //x=94.155 //y=1.21 //x2=95.275 //y2=1.18
cc_5874 ( N_noxref_24_c_9709_p N_Q_c_10376_n ) capacitor c=0.00361177f \
 //x=94.155 //y=1.52 //x2=95.275 //y2=1.18
cc_5875 ( N_noxref_24_c_9471_n N_Q_c_10376_n ) capacitor c=4.02408e-19 \
 //x=94.53 //y=0.71 //x2=95.275 //y2=1.18
cc_5876 ( N_noxref_24_c_9472_n N_Q_c_10376_n ) capacitor c=0.0036677f \
 //x=94.53 //y=1.365 //x2=95.275 //y2=1.18
cc_5877 ( N_noxref_24_c_9475_n N_Q_c_10376_n ) capacitor c=0.00776505f \
 //x=94.685 //y=1.21 //x2=95.275 //y2=1.18
cc_5878 ( N_noxref_24_c_9440_n N_Q_c_10382_n ) capacitor c=0.00786826f \
 //x=92.355 //y=2.22 //x2=92.175 //y2=1.18
cc_5879 ( N_noxref_24_c_9553_n N_Q_c_10382_n ) capacitor c=0.00152807f \
 //x=91.795 //y=1.25 //x2=92.175 //y2=1.18
cc_5880 ( N_noxref_24_c_9742_p N_Q_c_10382_n ) capacitor c=4.52813e-19 \
 //x=92.17 //y=0.75 //x2=92.175 //y2=1.18
cc_5881 ( N_noxref_24_c_9743_p N_Q_c_10382_n ) capacitor c=5.84553e-19 \
 //x=92.17 //y=1.405 //x2=92.175 //y2=1.18
cc_5882 ( N_noxref_24_c_9560_n N_Q_c_10382_n ) capacitor c=4.79299e-19 \
 //x=92.325 //y=1.25 //x2=92.175 //y2=1.18
cc_5883 ( N_noxref_24_c_9561_n N_Q_c_10382_n ) capacitor c=9.48308e-19 \
 //x=92.325 //y=1.56 //x2=92.175 //y2=1.18
cc_5884 ( N_noxref_24_M177_noxref_g N_Q_c_10433_n ) capacitor c=0.0179287f \
 //x=94.69 //y=6.025 //x2=95.265 //y2=5.21
cc_5885 ( N_noxref_24_M176_noxref_g N_Q_c_10397_n ) capacitor c=0.0132916f \
 //x=94.25 //y=6.025 //x2=94.555 //y2=5.21
cc_5886 ( N_noxref_24_c_9699_p N_Q_c_10397_n ) capacitor c=0.00405122f \
 //x=94.615 //y=4.795 //x2=94.555 //y2=5.21
cc_5887 ( N_noxref_24_c_9455_n N_Q_c_10384_n ) capacitor c=0.00314046f \
 //x=93.98 //y=2.08 //x2=95.83 //y2=4.07
cc_5888 ( N_noxref_24_c_9440_n N_Q_M55_noxref_d ) capacitor c=0.00540518f \
 //x=92.355 //y=2.22 //x2=88.54 //y2=0.905
cc_5889 ( N_noxref_24_c_9440_n N_Q_M57_noxref_d ) capacitor c=0.0054066f \
 //x=92.355 //y=2.22 //x2=91.87 //y2=0.905
cc_5890 ( N_noxref_24_c_9550_n N_Q_M57_noxref_d ) capacitor c=0.00217566f \
 //x=91.795 //y=0.905 //x2=91.87 //y2=0.905
cc_5891 ( N_noxref_24_c_9553_n N_Q_M57_noxref_d ) capacitor c=0.00711747f \
 //x=91.795 //y=1.25 //x2=91.87 //y2=0.905
cc_5892 ( N_noxref_24_c_9742_p N_Q_M57_noxref_d ) capacitor c=0.00234223f \
 //x=92.17 //y=0.75 //x2=91.87 //y2=0.905
cc_5893 ( N_noxref_24_c_9743_p N_Q_M57_noxref_d ) capacitor c=0.00602848f \
 //x=92.17 //y=1.405 //x2=91.87 //y2=0.905
cc_5894 ( N_noxref_24_c_9559_n N_Q_M57_noxref_d ) capacitor c=0.00132245f \
 //x=92.325 //y=0.905 //x2=91.87 //y2=0.905
cc_5895 ( N_noxref_24_c_9560_n N_Q_M57_noxref_d ) capacitor c=0.004434f \
 //x=92.325 //y=1.25 //x2=91.87 //y2=0.905
cc_5896 ( N_noxref_24_c_9561_n N_Q_M57_noxref_d ) capacitor c=0.00270197f \
 //x=92.325 //y=1.56 //x2=91.87 //y2=0.905
cc_5897 ( N_noxref_24_M177_noxref_g N_Q_M176_noxref_d ) capacitor c=0.0130327f \
 //x=94.69 //y=6.025 //x2=94.325 //y2=5.025
cc_5898 ( N_noxref_24_M50_noxref_d N_noxref_60_M48_noxref_s ) capacitor \
 c=0.00309936f //x=80.355 //y=0.915 //x2=77.415 //y2=0.375
cc_5899 ( N_noxref_24_c_9450_n N_noxref_61_c_12229_n ) capacitor c=0.00461316f \
 //x=80.945 //y=1.665 //x2=80.945 //y2=0.54
cc_5900 ( N_noxref_24_M50_noxref_d N_noxref_61_c_12229_n ) capacitor \
 c=0.0116817f //x=80.355 //y=0.915 //x2=80.945 //y2=0.54
cc_5901 ( N_noxref_24_c_9630_n N_noxref_61_c_12257_n ) capacitor c=0.0200405f \
 //x=80.63 //y=1.665 //x2=80.06 //y2=0.995
cc_5902 ( N_noxref_24_M50_noxref_d N_noxref_61_M49_noxref_d ) capacitor \
 c=5.27807e-19 //x=80.355 //y=0.915 //x2=78.82 //y2=0.91
cc_5903 ( N_noxref_24_c_9450_n N_noxref_61_M50_noxref_s ) capacitor \
 c=0.0195547f //x=80.945 //y=1.665 //x2=79.925 //y2=0.375
cc_5904 ( N_noxref_24_c_9451_n N_noxref_61_M50_noxref_s ) capacitor \
 c=2.38752e-19 //x=81.03 //y=2.22 //x2=79.925 //y2=0.375
cc_5905 ( N_noxref_24_M50_noxref_d N_noxref_61_M50_noxref_s ) capacitor \
 c=0.0426368f //x=80.355 //y=0.915 //x2=79.925 //y2=0.375
cc_5906 ( N_noxref_24_c_9433_n N_noxref_62_c_12302_n ) capacitor c=0.00642985f \
 //x=82.765 //y=2.22 //x2=82.36 //y2=1.505
cc_5907 ( N_noxref_24_c_9450_n N_noxref_62_c_12302_n ) capacitor c=3.84569e-19 \
 //x=80.945 //y=1.665 //x2=82.36 //y2=1.505
cc_5908 ( N_noxref_24_c_9460_n N_noxref_62_c_12302_n ) capacitor c=0.0034165f \
 //x=82.58 //y=1.915 //x2=82.36 //y2=1.505
cc_5909 ( N_noxref_24_c_9433_n N_noxref_62_c_12278_n ) capacitor c=0.0112993f \
 //x=82.765 //y=2.22 //x2=83.245 //y2=1.59
cc_5910 ( N_noxref_24_c_9440_n N_noxref_62_c_12278_n ) capacitor c=0.00784493f \
 //x=92.355 //y=2.22 //x2=83.245 //y2=1.59
cc_5911 ( N_noxref_24_c_9446_n N_noxref_62_c_12278_n ) capacitor c=0.00350496f \
 //x=82.995 //y=2.22 //x2=83.245 //y2=1.59
cc_5912 ( N_noxref_24_c_9452_n N_noxref_62_c_12278_n ) capacitor c=0.0115361f \
 //x=82.88 //y=2.08 //x2=83.245 //y2=1.59
cc_5913 ( N_noxref_24_c_9459_n N_noxref_62_c_12278_n ) capacitor c=0.00697148f \
 //x=82.58 //y=1.53 //x2=83.245 //y2=1.59
cc_5914 ( N_noxref_24_c_9460_n N_noxref_62_c_12278_n ) capacitor c=0.0204849f \
 //x=82.58 //y=1.915 //x2=83.245 //y2=1.59
cc_5915 ( N_noxref_24_c_9462_n N_noxref_62_c_12278_n ) capacitor c=0.00610316f \
 //x=82.955 //y=1.375 //x2=83.245 //y2=1.59
cc_5916 ( N_noxref_24_c_9465_n N_noxref_62_c_12278_n ) capacitor c=0.00698822f \
 //x=83.11 //y=1.22 //x2=83.245 //y2=1.59
cc_5917 ( N_noxref_24_c_9440_n N_noxref_62_c_12295_n ) capacitor c=0.0203655f \
 //x=92.355 //y=2.22 //x2=84.215 //y2=1.59
cc_5918 ( N_noxref_24_c_9440_n N_noxref_62_M51_noxref_s ) capacitor \
 c=0.012425f //x=92.355 //y=2.22 //x2=82.225 //y2=0.375
cc_5919 ( N_noxref_24_c_9456_n N_noxref_62_M51_noxref_s ) capacitor \
 c=0.0327271f //x=82.58 //y=0.875 //x2=82.225 //y2=0.375
cc_5920 ( N_noxref_24_c_9459_n N_noxref_62_M51_noxref_s ) capacitor \
 c=7.99997e-19 //x=82.58 //y=1.53 //x2=82.225 //y2=0.375
cc_5921 ( N_noxref_24_c_9460_n N_noxref_62_M51_noxref_s ) capacitor \
 c=0.00122123f //x=82.58 //y=1.915 //x2=82.225 //y2=0.375
cc_5922 ( N_noxref_24_c_9463_n N_noxref_62_M51_noxref_s ) capacitor \
 c=0.0121427f //x=83.11 //y=0.875 //x2=82.225 //y2=0.375
cc_5923 ( N_noxref_24_M50_noxref_d N_noxref_62_M51_noxref_s ) capacitor \
 c=2.55333e-19 //x=80.355 //y=0.915 //x2=82.225 //y2=0.375
cc_5924 ( N_noxref_24_c_9440_n N_noxref_63_c_12329_n ) capacitor c=0.00657782f \
 //x=92.355 //y=2.22 //x2=84.785 //y2=0.995
cc_5925 ( N_noxref_24_c_9440_n N_noxref_63_c_12334_n ) capacitor c=0.00147946f \
 //x=92.355 //y=2.22 //x2=85.755 //y2=0.54
cc_5926 ( N_noxref_24_c_9440_n N_noxref_63_M53_noxref_s ) capacitor \
 c=0.00642985f //x=92.355 //y=2.22 //x2=84.735 //y2=0.375
cc_5927 ( N_noxref_24_c_9440_n N_noxref_64_c_12399_n ) capacitor c=0.0018561f \
 //x=92.355 //y=2.22 //x2=87.275 //y2=1.495
cc_5928 ( N_noxref_24_c_9440_n N_noxref_64_c_12381_n ) capacitor c=0.024432f \
 //x=92.355 //y=2.22 //x2=88.16 //y2=1.58
cc_5929 ( N_noxref_24_c_9440_n N_noxref_64_c_12388_n ) capacitor c=0.00649228f \
 //x=92.355 //y=2.22 //x2=88.245 //y2=1.495
cc_5930 ( N_noxref_24_c_9440_n N_noxref_64_c_12389_n ) capacitor c=0.00102132f \
 //x=92.355 //y=2.22 //x2=89.13 //y2=0.53
cc_5931 ( N_noxref_24_c_9440_n N_noxref_64_M54_noxref_s ) capacitor \
 c=0.00528401f //x=92.355 //y=2.22 //x2=87.14 //y2=0.365
cc_5932 ( N_noxref_24_c_9440_n N_noxref_65_c_12455_n ) capacitor c=0.00502209f \
 //x=92.355 //y=2.22 //x2=90.605 //y2=1.495
cc_5933 ( N_noxref_24_c_9440_n N_noxref_65_c_12438_n ) capacitor c=0.018617f \
 //x=92.355 //y=2.22 //x2=91.49 //y2=1.58
cc_5934 ( N_noxref_24_c_9440_n N_noxref_65_c_12444_n ) capacitor c=0.00528401f \
 //x=92.355 //y=2.22 //x2=91.575 //y2=1.495
cc_5935 ( N_noxref_24_c_9466_n N_noxref_65_c_12444_n ) capacitor c=0.0028747f \
 //x=92.325 //y=1.915 //x2=91.575 //y2=1.495
cc_5936 ( N_noxref_24_c_9550_n N_noxref_65_c_12445_n ) capacitor c=0.021566f \
 //x=91.795 //y=0.905 //x2=92.46 //y2=0.53
cc_5937 ( N_noxref_24_c_9559_n N_noxref_65_c_12445_n ) capacitor c=0.00781103f \
 //x=92.325 //y=0.905 //x2=92.46 //y2=0.53
cc_5938 ( N_noxref_24_c_9448_n N_noxref_65_M56_noxref_s ) capacitor \
 c=5.34178e-19 //x=93.865 //y=2.08 //x2=90.47 //y2=0.365
cc_5939 ( N_noxref_24_c_9449_n N_noxref_65_M56_noxref_s ) capacitor \
 c=0.00122678f //x=92.5 //y=2.08 //x2=90.47 //y2=0.365
cc_5940 ( N_noxref_24_c_9453_n N_noxref_65_M56_noxref_s ) capacitor \
 c=0.0156825f //x=92.5 //y=2.08 //x2=90.47 //y2=0.365
cc_5941 ( N_noxref_24_c_9550_n N_noxref_65_M56_noxref_s ) capacitor \
 c=0.0064603f //x=91.795 //y=0.905 //x2=90.47 //y2=0.365
cc_5942 ( N_noxref_24_c_9553_n N_noxref_65_M56_noxref_s ) capacitor \
 c=0.00629878f //x=91.795 //y=1.25 //x2=90.47 //y2=0.365
cc_5943 ( N_noxref_24_c_9559_n N_noxref_65_M56_noxref_s ) capacitor \
 c=0.0321601f //x=92.325 //y=0.905 //x2=90.47 //y2=0.365
cc_5944 ( N_noxref_24_c_9561_n N_noxref_65_M56_noxref_s ) capacitor \
 c=0.00244207f //x=92.325 //y=1.56 //x2=90.47 //y2=0.365
cc_5945 ( N_noxref_24_c_9466_n N_noxref_65_M56_noxref_s ) capacitor \
 c=0.00784558f //x=92.325 //y=1.915 //x2=90.47 //y2=0.365
cc_5946 ( N_noxref_24_c_9448_n N_noxref_66_c_12509_n ) capacitor c=0.00169534f \
 //x=93.865 //y=2.08 //x2=93.935 //y2=1.495
cc_5947 ( N_noxref_24_c_9455_n N_noxref_66_c_12509_n ) capacitor c=0.016698f \
 //x=93.98 //y=2.08 //x2=93.935 //y2=1.495
cc_5948 ( N_noxref_24_c_9470_n N_noxref_66_c_12509_n ) capacitor c=0.0034165f \
 //x=94.155 //y=1.915 //x2=93.935 //y2=1.495
cc_5949 ( N_noxref_24_c_9476_n N_noxref_66_c_12509_n ) capacitor c=0.00531095f \
 //x=93.98 //y=2.08 //x2=93.935 //y2=1.495
cc_5950 ( N_noxref_24_c_9448_n N_noxref_66_c_12493_n ) capacitor c=0.00222439f \
 //x=93.865 //y=2.08 //x2=94.82 //y2=1.58
cc_5951 ( N_noxref_24_c_9455_n N_noxref_66_c_12493_n ) capacitor c=0.00587616f \
 //x=93.98 //y=2.08 //x2=94.82 //y2=1.58
cc_5952 ( N_noxref_24_c_9709_p N_noxref_66_c_12493_n ) capacitor c=0.0061593f \
 //x=94.155 //y=1.52 //x2=94.82 //y2=1.58
cc_5953 ( N_noxref_24_c_9470_n N_noxref_66_c_12493_n ) capacitor c=0.0142098f \
 //x=94.155 //y=1.915 //x2=94.82 //y2=1.58
cc_5954 ( N_noxref_24_c_9472_n N_noxref_66_c_12493_n ) capacitor c=0.00991953f \
 //x=94.53 //y=1.365 //x2=94.82 //y2=1.58
cc_5955 ( N_noxref_24_c_9475_n N_noxref_66_c_12493_n ) capacitor c=0.00339872f \
 //x=94.685 //y=1.21 //x2=94.82 //y2=1.58
cc_5956 ( N_noxref_24_c_9476_n N_noxref_66_c_12493_n ) capacitor c=0.00147967f \
 //x=93.98 //y=2.08 //x2=94.82 //y2=1.58
cc_5957 ( N_noxref_24_c_9470_n N_noxref_66_c_12499_n ) capacitor c=6.71402e-19 \
 //x=94.155 //y=1.915 //x2=94.905 //y2=1.495
cc_5958 ( N_noxref_24_c_9467_n N_noxref_66_M58_noxref_s ) capacitor \
 c=0.0314164f //x=94.155 //y=0.865 //x2=93.8 //y2=0.365
cc_5959 ( N_noxref_24_c_9709_p N_noxref_66_M58_noxref_s ) capacitor \
 c=0.00110192f //x=94.155 //y=1.52 //x2=93.8 //y2=0.365
cc_5960 ( N_noxref_24_c_9473_n N_noxref_66_M58_noxref_s ) capacitor \
 c=0.0132463f //x=94.685 //y=0.865 //x2=93.8 //y2=0.365
cc_5961 ( N_noxref_25_c_9823_n N_noxref_26_c_9913_n ) capacitor c=0.0535575f \
 //x=93.915 //y=5.21 //x2=94.975 //y2=4.07
cc_5962 ( N_noxref_25_c_9827_n N_noxref_26_c_9913_n ) capacitor c=0.008149f \
 //x=92.125 //y=5.21 //x2=94.975 //y2=4.07
cc_5963 ( N_noxref_25_c_9838_n N_noxref_26_c_9913_n ) capacitor c=3.2507e-19 \
 //x=91.925 //y=5.21 //x2=94.975 //y2=4.07
cc_5964 ( N_noxref_25_c_9829_n N_noxref_26_c_9913_n ) capacitor c=0.0181202f \
 //x=91.215 //y=5.21 //x2=94.975 //y2=4.07
cc_5965 ( N_noxref_25_c_9830_n N_noxref_26_c_9913_n ) capacitor c=0.00337443f \
 //x=92.01 //y=5.295 //x2=94.975 //y2=4.07
cc_5966 ( N_noxref_25_c_9831_n N_noxref_26_c_9913_n ) capacitor c=0.0011253f \
 //x=94.03 //y=5.21 //x2=94.975 //y2=4.07
cc_5967 ( N_noxref_25_c_9882_n N_noxref_26_c_9913_n ) capacitor c=0.00358031f \
 //x=94.825 //y=6.91 //x2=94.975 //y2=4.07
cc_5968 ( N_noxref_25_c_9893_p N_noxref_26_M178_noxref_g ) capacitor \
 c=0.0150104f //x=95.705 //y=6.91 //x2=95.13 //y2=6.025
cc_5969 ( N_noxref_25_M177_noxref_d N_noxref_26_M178_noxref_g ) capacitor \
 c=0.0130327f //x=94.765 //y=5.025 //x2=95.13 //y2=6.025
cc_5970 ( N_noxref_25_c_9893_p N_noxref_26_M179_noxref_g ) capacitor \
 c=0.0163361f //x=95.705 //y=6.91 //x2=95.57 //y2=6.025
cc_5971 ( N_noxref_25_M179_noxref_d N_noxref_26_M179_noxref_g ) capacitor \
 c=0.0351101f //x=95.645 //y=5.025 //x2=95.57 //y2=6.025
cc_5972 ( N_noxref_25_c_9882_n N_Q_c_10433_n ) capacitor c=0.00102709f \
 //x=94.825 //y=6.91 //x2=95.265 //y2=5.21
cc_5973 ( N_noxref_25_c_9893_p N_Q_c_10433_n ) capacitor c=0.00101874f \
 //x=95.705 //y=6.91 //x2=95.265 //y2=5.21
cc_5974 ( N_noxref_25_M177_noxref_d N_Q_c_10433_n ) capacitor c=0.012404f \
 //x=94.765 //y=5.025 //x2=95.265 //y2=5.21
cc_5975 ( N_noxref_25_c_9823_n N_Q_c_10397_n ) capacitor c=0.00602307f \
 //x=93.915 //y=5.21 //x2=94.555 //y2=5.21
cc_5976 ( N_noxref_25_c_9831_n N_Q_c_10397_n ) capacitor c=0.0683084f \
 //x=94.03 //y=5.21 //x2=94.555 //y2=5.21
cc_5977 ( N_noxref_25_c_9893_p N_Q_c_10398_n ) capacitor c=0.00173777f \
 //x=95.705 //y=6.91 //x2=95.745 //y2=5.21
cc_5978 ( N_noxref_25_M179_noxref_d N_Q_c_10398_n ) capacitor c=0.0154399f \
 //x=95.645 //y=5.025 //x2=95.745 //y2=5.21
cc_5979 ( N_noxref_25_c_9831_n N_Q_c_10384_n ) capacitor c=3.02032e-19 \
 //x=94.03 //y=5.21 //x2=95.83 //y2=4.07
cc_5980 ( N_noxref_25_c_9823_n N_Q_M176_noxref_d ) capacitor c=8.04912e-19 \
 //x=93.915 //y=5.21 //x2=94.325 //y2=5.025
cc_5981 ( N_noxref_25_c_9882_n N_Q_M176_noxref_d ) capacitor c=0.0117542f \
 //x=94.825 //y=6.91 //x2=94.325 //y2=5.025
cc_5982 ( N_noxref_25_M177_noxref_d N_Q_M176_noxref_d ) capacitor c=0.0458293f \
 //x=94.765 //y=5.025 //x2=94.325 //y2=5.025
cc_5983 ( N_noxref_25_c_9831_n N_Q_M178_noxref_d ) capacitor c=9.91979e-19 \
 //x=94.03 //y=5.21 //x2=95.205 //y2=5.025
cc_5984 ( N_noxref_25_c_9893_p N_Q_M178_noxref_d ) capacitor c=0.0118172f \
 //x=95.705 //y=6.91 //x2=95.205 //y2=5.025
cc_5985 ( N_noxref_25_M177_noxref_d N_Q_M178_noxref_d ) capacitor c=0.0458293f \
 //x=94.765 //y=5.025 //x2=95.205 //y2=5.025
cc_5986 ( N_noxref_25_M179_noxref_d N_Q_M178_noxref_d ) capacitor c=0.0458293f \
 //x=95.645 //y=5.025 //x2=95.205 //y2=5.025
cc_5987 ( N_noxref_26_c_9913_n Q ) capacitor c=0.0244534f //x=94.975 //y=4.07 \
 //x2=95.83 //y2=4.07
cc_5988 ( N_noxref_26_c_9919_n Q ) capacitor c=0.00238921f //x=95.09 //y=2.08 \
 //x2=95.83 //y2=4.07
cc_5989 ( N_noxref_26_c_9913_n N_Q_c_10368_n ) capacitor c=0.00257374f \
 //x=94.975 //y=4.07 //x2=91.945 //y2=1.18
cc_5990 ( N_noxref_26_c_10035_n N_Q_c_10368_n ) capacitor c=4.67724e-19 \
 //x=88.995 //y=0.905 //x2=91.945 //y2=1.18
cc_5991 ( N_noxref_26_c_10036_n N_Q_c_10368_n ) capacitor c=0.00683548f \
 //x=88.995 //y=1.25 //x2=91.945 //y2=1.18
cc_5992 ( N_noxref_26_c_9913_n N_Q_c_10375_n ) capacitor c=3.47851e-19 \
 //x=94.975 //y=4.07 //x2=88.845 //y2=1.18
cc_5993 ( N_noxref_26_c_10026_n N_Q_c_10375_n ) capacitor c=3.66947e-19 \
 //x=88.465 //y=0.905 //x2=88.845 //y2=1.18
cc_5994 ( N_noxref_26_c_10029_n N_Q_c_10375_n ) capacitor c=0.00353233f \
 //x=88.465 //y=1.25 //x2=88.845 //y2=1.18
cc_5995 ( N_noxref_26_c_10031_n N_Q_c_10375_n ) capacitor c=0.00278363f \
 //x=88.465 //y=1.56 //x2=88.845 //y2=1.18
cc_5996 ( N_noxref_26_c_10280_p N_Q_c_10375_n ) capacitor c=4.06815e-19 \
 //x=88.84 //y=0.75 //x2=88.845 //y2=1.18
cc_5997 ( N_noxref_26_c_10242_n N_Q_c_10375_n ) capacitor c=5.84553e-19 \
 //x=88.84 //y=1.405 //x2=88.845 //y2=1.18
cc_5998 ( N_noxref_26_c_10036_n N_Q_c_10375_n ) capacitor c=0.00132321f \
 //x=88.995 //y=1.25 //x2=88.845 //y2=1.18
cc_5999 ( N_noxref_26_c_9913_n N_Q_c_10376_n ) capacitor c=0.011537f \
 //x=94.975 //y=4.07 //x2=95.275 //y2=1.18
cc_6000 ( N_noxref_26_c_9919_n N_Q_c_10376_n ) capacitor c=0.00449159f \
 //x=95.09 //y=2.08 //x2=95.275 //y2=1.18
cc_6001 ( N_noxref_26_c_10243_n N_Q_c_10376_n ) capacitor c=6.33948e-19 \
 //x=95.125 //y=0.905 //x2=95.275 //y2=1.18
cc_6002 ( N_noxref_26_c_10246_n N_Q_c_10376_n ) capacitor c=0.0043333f \
 //x=95.125 //y=1.255 //x2=95.275 //y2=1.18
cc_6003 ( N_noxref_26_c_10247_n N_Q_c_10376_n ) capacitor c=0.0040799f \
 //x=95.125 //y=1.56 //x2=95.275 //y2=1.18
cc_6004 ( N_noxref_26_c_10288_p N_Q_c_10376_n ) capacitor c=4.52813e-19 \
 //x=95.5 //y=0.75 //x2=95.275 //y2=1.18
cc_6005 ( N_noxref_26_c_10250_n N_Q_c_10376_n ) capacitor c=0.00296491f \
 //x=95.5 //y=1.405 //x2=95.275 //y2=1.18
cc_6006 ( N_noxref_26_c_10251_n N_Q_c_10376_n ) capacitor c=2.65983e-19 \
 //x=95.655 //y=0.905 //x2=95.275 //y2=1.18
cc_6007 ( N_noxref_26_c_10252_n N_Q_c_10376_n ) capacitor c=0.00362989f \
 //x=95.655 //y=1.255 //x2=95.275 //y2=1.18
cc_6008 ( N_noxref_26_c_10254_n N_Q_c_10376_n ) capacitor c=5.89141e-19 \
 //x=95.09 //y=2.08 //x2=95.275 //y2=1.18
cc_6009 ( N_noxref_26_c_9913_n N_Q_c_10382_n ) capacitor c=2.93491e-19 \
 //x=94.975 //y=4.07 //x2=92.175 //y2=1.18
cc_6010 ( N_noxref_26_c_9913_n N_Q_c_10433_n ) capacitor c=0.00154966f \
 //x=94.975 //y=4.07 //x2=95.265 //y2=5.21
cc_6011 ( N_noxref_26_c_10237_n N_Q_c_10433_n ) capacitor c=0.0128151f \
 //x=95.11 //y=4.705 //x2=95.265 //y2=5.21
cc_6012 ( N_noxref_26_M178_noxref_g N_Q_c_10433_n ) capacitor c=0.0167296f \
 //x=95.13 //y=6.025 //x2=95.265 //y2=5.21
cc_6013 ( N_noxref_26_c_10257_n N_Q_c_10433_n ) capacitor c=0.00368327f \
 //x=95.11 //y=4.705 //x2=95.265 //y2=5.21
cc_6014 ( N_noxref_26_c_9913_n N_Q_c_10397_n ) capacitor c=0.0138451f \
 //x=94.975 //y=4.07 //x2=94.555 //y2=5.21
cc_6015 ( N_noxref_26_M179_noxref_g N_Q_c_10398_n ) capacitor c=0.0222938f \
 //x=95.57 //y=6.025 //x2=95.745 //y2=5.21
cc_6016 ( N_noxref_26_c_10250_n N_Q_c_10383_n ) capacitor c=0.00810194f \
 //x=95.5 //y=1.405 //x2=95.745 //y2=1.645
cc_6017 ( N_noxref_26_c_10301_p N_Q_c_10492_n ) capacitor c=0.00671029f \
 //x=95.09 //y=1.915 //x2=95.475 //y2=1.645
cc_6018 ( N_noxref_26_c_9913_n N_Q_c_10384_n ) capacitor c=0.00246068f \
 //x=94.975 //y=4.07 //x2=95.83 //y2=4.07
cc_6019 ( N_noxref_26_c_9919_n N_Q_c_10384_n ) capacitor c=0.082481f //x=95.09 \
 //y=2.08 //x2=95.83 //y2=4.07
cc_6020 ( N_noxref_26_c_10237_n N_Q_c_10384_n ) capacitor c=0.00998395f \
 //x=95.11 //y=4.705 //x2=95.83 //y2=4.07
cc_6021 ( N_noxref_26_c_10305_p N_Q_c_10384_n ) capacitor c=0.0143966f \
 //x=95.495 //y=4.795 //x2=95.83 //y2=4.07
cc_6022 ( N_noxref_26_c_10254_n N_Q_c_10384_n ) capacitor c=0.00666633f \
 //x=95.09 //y=2.08 //x2=95.83 //y2=4.07
cc_6023 ( N_noxref_26_c_10301_p N_Q_c_10384_n ) capacitor c=0.0033061f \
 //x=95.09 //y=1.915 //x2=95.83 //y2=4.07
cc_6024 ( N_noxref_26_c_10257_n N_Q_c_10384_n ) capacitor c=0.00526987f \
 //x=95.11 //y=4.705 //x2=95.83 //y2=4.07
cc_6025 ( N_noxref_26_c_10305_p N_Q_c_10500_n ) capacitor c=0.00410596f \
 //x=95.495 //y=4.795 //x2=95.35 //y2=5.21
cc_6026 ( N_noxref_26_c_10026_n N_Q_M55_noxref_d ) capacitor c=0.00218556f \
 //x=88.465 //y=0.905 //x2=88.54 //y2=0.905
cc_6027 ( N_noxref_26_c_10029_n N_Q_M55_noxref_d ) capacitor c=0.00327871f \
 //x=88.465 //y=1.25 //x2=88.54 //y2=0.905
cc_6028 ( N_noxref_26_c_10031_n N_Q_M55_noxref_d ) capacitor c=0.00292542f \
 //x=88.465 //y=1.56 //x2=88.54 //y2=0.905
cc_6029 ( N_noxref_26_c_10280_p N_Q_M55_noxref_d ) capacitor c=0.00235569f \
 //x=88.84 //y=0.75 //x2=88.54 //y2=0.905
cc_6030 ( N_noxref_26_c_10242_n N_Q_M55_noxref_d ) capacitor c=0.00613695f \
 //x=88.84 //y=1.405 //x2=88.54 //y2=0.905
cc_6031 ( N_noxref_26_c_10035_n N_Q_M55_noxref_d ) capacitor c=0.00131413f \
 //x=88.995 //y=0.905 //x2=88.54 //y2=0.905
cc_6032 ( N_noxref_26_c_10036_n N_Q_M55_noxref_d ) capacitor c=0.00676348f \
 //x=88.995 //y=1.25 //x2=88.54 //y2=0.905
cc_6033 ( N_noxref_26_c_10243_n N_Q_M59_noxref_d ) capacitor c=0.00226395f \
 //x=95.125 //y=0.905 //x2=95.2 //y2=0.905
cc_6034 ( N_noxref_26_c_10246_n N_Q_M59_noxref_d ) capacitor c=0.004517f \
 //x=95.125 //y=1.255 //x2=95.2 //y2=0.905
cc_6035 ( N_noxref_26_c_10247_n N_Q_M59_noxref_d ) capacitor c=0.00655125f \
 //x=95.125 //y=1.56 //x2=95.2 //y2=0.905
cc_6036 ( N_noxref_26_c_10288_p N_Q_M59_noxref_d ) capacitor c=0.00241003f \
 //x=95.5 //y=0.75 //x2=95.2 //y2=0.905
cc_6037 ( N_noxref_26_c_10250_n N_Q_M59_noxref_d ) capacitor c=0.0159024f \
 //x=95.5 //y=1.405 //x2=95.2 //y2=0.905
cc_6038 ( N_noxref_26_c_10251_n N_Q_M59_noxref_d ) capacitor c=0.00132831f \
 //x=95.655 //y=0.905 //x2=95.2 //y2=0.905
cc_6039 ( N_noxref_26_c_10252_n N_Q_M59_noxref_d ) capacitor c=0.00330743f \
 //x=95.655 //y=1.255 //x2=95.2 //y2=0.905
cc_6040 ( N_noxref_26_M178_noxref_g N_Q_M178_noxref_d ) capacitor c=0.0130327f \
 //x=95.13 //y=6.025 //x2=95.205 //y2=5.025
cc_6041 ( N_noxref_26_M179_noxref_g N_Q_M178_noxref_d ) capacitor c=0.0136385f \
 //x=95.57 //y=6.025 //x2=95.205 //y2=5.025
cc_6042 ( N_noxref_26_M32_noxref_d N_noxref_48_M30_noxref_s ) capacitor \
 c=0.00309936f //x=51.495 //y=0.915 //x2=48.555 //y2=0.375
cc_6043 ( N_noxref_26_c_9915_n N_noxref_49_c_11617_n ) capacitor c=0.00457167f \
 //x=52.085 //y=1.665 //x2=52.085 //y2=0.54
cc_6044 ( N_noxref_26_M32_noxref_d N_noxref_49_c_11617_n ) capacitor \
 c=0.0115903f //x=51.495 //y=0.915 //x2=52.085 //y2=0.54
cc_6045 ( N_noxref_26_c_10146_n N_noxref_49_c_11629_n ) capacitor c=0.0200405f \
 //x=51.77 //y=1.665 //x2=51.2 //y2=0.995
cc_6046 ( N_noxref_26_M32_noxref_d N_noxref_49_M31_noxref_d ) capacitor \
 c=5.27807e-19 //x=51.495 //y=0.915 //x2=49.96 //y2=0.91
cc_6047 ( N_noxref_26_c_9915_n N_noxref_49_M32_noxref_s ) capacitor \
 c=0.0196084f //x=52.085 //y=1.665 //x2=51.065 //y2=0.375
cc_6048 ( N_noxref_26_M32_noxref_d N_noxref_49_M32_noxref_s ) capacitor \
 c=0.0426368f //x=51.495 //y=0.915 //x2=51.065 //y2=0.375
cc_6049 ( N_noxref_26_c_9915_n N_noxref_50_c_11680_n ) capacitor c=3.84569e-19 \
 //x=52.085 //y=1.665 //x2=53.5 //y2=1.505
cc_6050 ( N_noxref_26_c_9925_n N_noxref_50_c_11680_n ) capacitor c=0.0034165f \
 //x=53.72 //y=1.915 //x2=53.5 //y2=1.505
cc_6051 ( N_noxref_26_c_9916_n N_noxref_50_c_11664_n ) capacitor c=0.0115578f \
 //x=54.02 //y=2.08 //x2=54.385 //y2=1.59
cc_6052 ( N_noxref_26_c_9924_n N_noxref_50_c_11664_n ) capacitor c=0.00697148f \
 //x=53.72 //y=1.53 //x2=54.385 //y2=1.59
cc_6053 ( N_noxref_26_c_9925_n N_noxref_50_c_11664_n ) capacitor c=0.0204849f \
 //x=53.72 //y=1.915 //x2=54.385 //y2=1.59
cc_6054 ( N_noxref_26_c_9927_n N_noxref_50_c_11664_n ) capacitor c=0.00610316f \
 //x=54.095 //y=1.375 //x2=54.385 //y2=1.59
cc_6055 ( N_noxref_26_c_9930_n N_noxref_50_c_11664_n ) capacitor c=0.00698822f \
 //x=54.25 //y=1.22 //x2=54.385 //y2=1.59
cc_6056 ( N_noxref_26_c_9921_n N_noxref_50_M33_noxref_s ) capacitor \
 c=0.0327271f //x=53.72 //y=0.875 //x2=53.365 //y2=0.375
cc_6057 ( N_noxref_26_c_9924_n N_noxref_50_M33_noxref_s ) capacitor \
 c=7.99997e-19 //x=53.72 //y=1.53 //x2=53.365 //y2=0.375
cc_6058 ( N_noxref_26_c_9925_n N_noxref_50_M33_noxref_s ) capacitor \
 c=0.00122123f //x=53.72 //y=1.915 //x2=53.365 //y2=0.375
cc_6059 ( N_noxref_26_c_9928_n N_noxref_50_M33_noxref_s ) capacitor \
 c=0.0121427f //x=54.25 //y=0.875 //x2=53.365 //y2=0.375
cc_6060 ( N_noxref_26_M32_noxref_d N_noxref_50_M33_noxref_s ) capacitor \
 c=2.55333e-19 //x=51.495 //y=0.915 //x2=53.365 //y2=0.375
cc_6061 ( N_noxref_26_c_10031_n N_noxref_64_c_12388_n ) capacitor \
 c=0.00746306f //x=88.465 //y=1.56 //x2=88.245 //y2=1.495
cc_6062 ( N_noxref_26_c_9931_n N_noxref_64_c_12388_n ) capacitor c=0.00173579f \
 //x=88.43 //y=2.08 //x2=88.245 //y2=1.495
cc_6063 ( N_noxref_26_c_9917_n N_noxref_64_c_12389_n ) capacitor c=0.00156604f \
 //x=88.43 //y=2.08 //x2=89.13 //y2=0.53
cc_6064 ( N_noxref_26_c_10026_n N_noxref_64_c_12389_n ) capacitor c=0.0200006f \
 //x=88.465 //y=0.905 //x2=89.13 //y2=0.53
cc_6065 ( N_noxref_26_c_10035_n N_noxref_64_c_12389_n ) capacitor \
 c=0.00825432f //x=88.995 //y=0.905 //x2=89.13 //y2=0.53
cc_6066 ( N_noxref_26_c_9931_n N_noxref_64_c_12389_n ) capacitor c=2.1838e-19 \
 //x=88.43 //y=2.08 //x2=89.13 //y2=0.53
cc_6067 ( N_noxref_26_c_10026_n N_noxref_64_M54_noxref_s ) capacitor \
 c=0.00746306f //x=88.465 //y=0.905 //x2=87.14 //y2=0.365
cc_6068 ( N_noxref_26_c_10031_n N_noxref_64_M54_noxref_s ) capacitor \
 c=0.0021955f //x=88.465 //y=1.56 //x2=87.14 //y2=0.365
cc_6069 ( N_noxref_26_c_10035_n N_noxref_64_M54_noxref_s ) capacitor \
 c=0.0133026f //x=88.995 //y=0.905 //x2=87.14 //y2=0.365
cc_6070 ( N_noxref_26_c_10036_n N_noxref_64_M54_noxref_s ) capacitor \
 c=0.00793126f //x=88.995 //y=1.25 //x2=87.14 //y2=0.365
cc_6071 ( N_noxref_26_c_10355_p N_noxref_64_M54_noxref_s ) capacitor \
 c=0.00392195f //x=88.43 //y=1.915 //x2=87.14 //y2=0.365
cc_6072 ( N_noxref_26_c_9913_n N_noxref_66_c_12493_n ) capacitor c=0.00631223f \
 //x=94.975 //y=4.07 //x2=94.82 //y2=1.58
cc_6073 ( N_noxref_26_c_9913_n N_noxref_66_c_12499_n ) capacitor c=0.00108825f \
 //x=94.975 //y=4.07 //x2=94.905 //y2=1.495
cc_6074 ( N_noxref_26_c_10247_n N_noxref_66_c_12499_n ) capacitor \
 c=0.00698471f //x=95.125 //y=1.56 //x2=94.905 //y2=1.495
cc_6075 ( N_noxref_26_c_10254_n N_noxref_66_c_12499_n ) capacitor \
 c=0.00171785f //x=95.09 //y=2.08 //x2=94.905 //y2=1.495
cc_6076 ( N_noxref_26_c_9919_n N_noxref_66_c_12500_n ) capacitor c=0.00118117f \
 //x=95.09 //y=2.08 //x2=95.79 //y2=0.53
cc_6077 ( N_noxref_26_c_10243_n N_noxref_66_c_12500_n ) capacitor c=0.0191024f \
 //x=95.125 //y=0.905 //x2=95.79 //y2=0.53
cc_6078 ( N_noxref_26_c_10251_n N_noxref_66_c_12500_n ) capacitor \
 c=0.00655165f //x=95.655 //y=0.905 //x2=95.79 //y2=0.53
cc_6079 ( N_noxref_26_c_10254_n N_noxref_66_c_12500_n ) capacitor c=2.1838e-19 \
 //x=95.09 //y=2.08 //x2=95.79 //y2=0.53
cc_6080 ( N_noxref_26_c_10243_n N_noxref_66_M58_noxref_s ) capacitor \
 c=0.00698471f //x=95.125 //y=0.905 //x2=93.8 //y2=0.365
cc_6081 ( N_noxref_26_c_10250_n N_noxref_66_M58_noxref_s ) capacitor \
 c=0.00316186f //x=95.5 //y=1.405 //x2=93.8 //y2=0.365
cc_6082 ( N_noxref_26_c_10251_n N_noxref_66_M58_noxref_s ) capacitor \
 c=0.0142835f //x=95.655 //y=0.905 //x2=93.8 //y2=0.365
cc_6083 ( N_Q_c_10368_n N_noxref_64_c_12389_n ) capacitor c=0.00641749f \
 //x=91.945 //y=1.18 //x2=89.13 //y2=0.53
cc_6084 ( N_Q_c_10375_n N_noxref_64_c_12389_n ) capacitor c=0.00219859f \
 //x=88.845 //y=1.18 //x2=89.13 //y2=0.53
cc_6085 ( N_Q_M55_noxref_d N_noxref_64_c_12389_n ) capacitor c=0.0136817f \
 //x=88.54 //y=0.905 //x2=89.13 //y2=0.53
cc_6086 ( N_Q_c_10368_n N_noxref_64_M54_noxref_s ) capacitor c=0.0197032f \
 //x=91.945 //y=1.18 //x2=87.14 //y2=0.365
cc_6087 ( N_Q_c_10375_n N_noxref_64_M54_noxref_s ) capacitor c=0.00804471f \
 //x=88.845 //y=1.18 //x2=87.14 //y2=0.365
cc_6088 ( N_Q_M55_noxref_d N_noxref_64_M54_noxref_s ) capacitor c=0.0458734f \
 //x=88.54 //y=0.905 //x2=87.14 //y2=0.365
cc_6089 ( N_Q_c_10368_n N_noxref_65_c_12438_n ) capacitor c=0.0202902f \
 //x=91.945 //y=1.18 //x2=91.49 //y2=1.58
cc_6090 ( N_Q_c_10368_n N_noxref_65_c_12445_n ) capacitor c=0.00641749f \
 //x=91.945 //y=1.18 //x2=92.46 //y2=0.53
cc_6091 ( N_Q_c_10376_n N_noxref_65_c_12445_n ) capacitor c=0.00641749f \
 //x=95.275 //y=1.18 //x2=92.46 //y2=0.53
cc_6092 ( N_Q_c_10382_n N_noxref_65_c_12445_n ) capacitor c=0.0015838f \
 //x=92.175 //y=1.18 //x2=92.46 //y2=0.53
cc_6093 ( N_Q_M57_noxref_d N_noxref_65_c_12445_n ) capacitor c=0.0130616f \
 //x=91.87 //y=0.905 //x2=92.46 //y2=0.53
cc_6094 ( N_Q_c_10368_n N_noxref_65_M56_noxref_s ) capacitor c=0.0422002f \
 //x=91.945 //y=1.18 //x2=90.47 //y2=0.365
cc_6095 ( N_Q_c_10376_n N_noxref_65_M56_noxref_s ) capacitor c=0.019112f \
 //x=95.275 //y=1.18 //x2=90.47 //y2=0.365
cc_6096 ( N_Q_c_10382_n N_noxref_65_M56_noxref_s ) capacitor c=0.00279707f \
 //x=92.175 //y=1.18 //x2=90.47 //y2=0.365
cc_6097 ( N_Q_M57_noxref_d N_noxref_65_M56_noxref_s ) capacitor c=0.0444718f \
 //x=91.87 //y=0.905 //x2=90.47 //y2=0.365
cc_6098 ( N_Q_c_10492_n N_noxref_66_c_12509_n ) capacitor c=2.73698e-19 \
 //x=95.475 //y=1.645 //x2=93.935 //y2=1.495
cc_6099 ( N_Q_c_10376_n N_noxref_66_c_12493_n ) capacitor c=0.0234642f \
 //x=95.275 //y=1.18 //x2=94.82 //y2=1.58
cc_6100 ( N_Q_c_10492_n N_noxref_66_c_12499_n ) capacitor c=0.0195484f \
 //x=95.475 //y=1.645 //x2=94.905 //y2=1.495
cc_6101 ( N_Q_c_10376_n N_noxref_66_c_12500_n ) capacitor c=0.0069137f \
 //x=95.275 //y=1.18 //x2=95.79 //y2=0.53
cc_6102 ( N_Q_c_10383_n N_noxref_66_c_12500_n ) capacitor c=0.00458011f \
 //x=95.745 //y=1.645 //x2=95.79 //y2=0.53
cc_6103 ( N_Q_M59_noxref_d N_noxref_66_c_12500_n ) capacitor c=0.0132979f \
 //x=95.2 //y=0.905 //x2=95.79 //y2=0.53
cc_6104 ( Q N_noxref_66_M58_noxref_s ) capacitor c=2.62341e-19 //x=95.83 \
 //y=4.07 //x2=93.8 //y2=0.365
cc_6105 ( N_Q_c_10376_n N_noxref_66_M58_noxref_s ) capacitor c=0.0513705f \
 //x=95.275 //y=1.18 //x2=93.8 //y2=0.365
cc_6106 ( N_Q_c_10383_n N_noxref_66_M58_noxref_s ) capacitor c=0.0154295f \
 //x=95.745 //y=1.645 //x2=93.8 //y2=0.365
cc_6107 ( N_Q_M59_noxref_d N_noxref_66_M58_noxref_s ) capacitor c=0.0438441f \
 //x=95.2 //y=0.905 //x2=93.8 //y2=0.365
cc_6108 ( N_noxref_28_c_10549_n N_noxref_29_c_10591_n ) capacitor c=0.0131801f \
 //x=2.445 //y=0.54 //x2=3.015 //y2=0.995
cc_6109 ( N_noxref_28_c_10566_n N_noxref_29_c_10591_n ) capacitor \
 c=0.00980353f //x=2.445 //y=1.59 //x2=3.015 //y2=0.995
cc_6110 ( N_noxref_28_M0_noxref_s N_noxref_29_c_10591_n ) capacitor \
 c=0.0221661f //x=0.455 //y=0.375 //x2=3.015 //y2=0.995
cc_6111 ( N_noxref_28_M0_noxref_s N_noxref_29_c_10593_n ) capacitor \
 c=0.0180035f //x=0.455 //y=0.375 //x2=3.1 //y2=0.625
cc_6112 ( N_noxref_28_c_10549_n N_noxref_29_M1_noxref_d ) capacitor \
 c=0.0128687f //x=2.445 //y=0.54 //x2=1.86 //y2=0.91
cc_6113 ( N_noxref_28_c_10566_n N_noxref_29_M1_noxref_d ) capacitor \
 c=0.00888766f //x=2.445 //y=1.59 //x2=1.86 //y2=0.91
cc_6114 ( N_noxref_28_M0_noxref_s N_noxref_29_M1_noxref_d ) capacitor \
 c=0.0159202f //x=0.455 //y=0.375 //x2=1.86 //y2=0.91
cc_6115 ( N_noxref_28_M0_noxref_s N_noxref_29_M2_noxref_s ) capacitor \
 c=0.0213553f //x=0.455 //y=0.375 //x2=2.965 //y2=0.375
cc_6116 ( N_noxref_29_c_10598_n N_noxref_30_M3_noxref_s ) capacitor \
 c=0.00191848f //x=4.07 //y=0.625 //x2=5.265 //y2=0.375
cc_6117 ( N_noxref_30_c_10650_n N_noxref_31_c_10692_n ) capacitor c=0.0131877f \
 //x=7.255 //y=0.54 //x2=7.825 //y2=0.995
cc_6118 ( N_noxref_30_c_10673_n N_noxref_31_c_10692_n ) capacitor \
 c=0.00981707f //x=7.255 //y=1.59 //x2=7.825 //y2=0.995
cc_6119 ( N_noxref_30_M3_noxref_s N_noxref_31_c_10692_n ) capacitor \
 c=0.0221661f //x=5.265 //y=0.375 //x2=7.825 //y2=0.995
cc_6120 ( N_noxref_30_M3_noxref_s N_noxref_31_c_10694_n ) capacitor \
 c=0.0180035f //x=5.265 //y=0.375 //x2=7.91 //y2=0.625
cc_6121 ( N_noxref_30_c_10650_n N_noxref_31_M4_noxref_d ) capacitor \
 c=0.0127191f //x=7.255 //y=0.54 //x2=6.67 //y2=0.91
cc_6122 ( N_noxref_30_c_10673_n N_noxref_31_M4_noxref_d ) capacitor \
 c=0.00861161f //x=7.255 //y=1.59 //x2=6.67 //y2=0.91
cc_6123 ( N_noxref_30_M3_noxref_s N_noxref_31_M4_noxref_d ) capacitor \
 c=0.0159202f //x=5.265 //y=0.375 //x2=6.67 //y2=0.91
cc_6124 ( N_noxref_30_M3_noxref_s N_noxref_31_M5_noxref_s ) capacitor \
 c=0.0213553f //x=5.265 //y=0.375 //x2=7.775 //y2=0.375
cc_6125 ( N_noxref_31_c_10699_n N_noxref_32_M6_noxref_s ) capacitor \
 c=0.00191848f //x=8.88 //y=0.625 //x2=10.075 //y2=0.375
cc_6126 ( N_noxref_32_c_10751_n N_noxref_33_c_10793_n ) capacitor c=0.0131877f \
 //x=12.065 //y=0.54 //x2=12.635 //y2=0.995
cc_6127 ( N_noxref_32_c_10774_n N_noxref_33_c_10793_n ) capacitor \
 c=0.00981707f //x=12.065 //y=1.59 //x2=12.635 //y2=0.995
cc_6128 ( N_noxref_32_M6_noxref_s N_noxref_33_c_10793_n ) capacitor \
 c=0.0221661f //x=10.075 //y=0.375 //x2=12.635 //y2=0.995
cc_6129 ( N_noxref_32_M6_noxref_s N_noxref_33_c_10795_n ) capacitor \
 c=0.0180035f //x=10.075 //y=0.375 //x2=12.72 //y2=0.625
cc_6130 ( N_noxref_32_c_10751_n N_noxref_33_M7_noxref_d ) capacitor \
 c=0.0127191f //x=12.065 //y=0.54 //x2=11.48 //y2=0.91
cc_6131 ( N_noxref_32_c_10774_n N_noxref_33_M7_noxref_d ) capacitor \
 c=0.00861161f //x=12.065 //y=1.59 //x2=11.48 //y2=0.91
cc_6132 ( N_noxref_32_M6_noxref_s N_noxref_33_M7_noxref_d ) capacitor \
 c=0.0159202f //x=10.075 //y=0.375 //x2=11.48 //y2=0.91
cc_6133 ( N_noxref_32_M6_noxref_s N_noxref_33_M8_noxref_s ) capacitor \
 c=0.0213553f //x=10.075 //y=0.375 //x2=12.585 //y2=0.375
cc_6134 ( N_noxref_33_c_10800_n N_noxref_34_M9_noxref_s ) capacitor \
 c=0.00191848f //x=13.69 //y=0.625 //x2=14.885 //y2=0.375
cc_6135 ( N_noxref_34_c_10852_n N_noxref_35_c_10894_n ) capacitor c=0.0131877f \
 //x=16.875 //y=0.54 //x2=17.445 //y2=0.995
cc_6136 ( N_noxref_34_c_10875_n N_noxref_35_c_10894_n ) capacitor \
 c=0.00981707f //x=16.875 //y=1.59 //x2=17.445 //y2=0.995
cc_6137 ( N_noxref_34_M9_noxref_s N_noxref_35_c_10894_n ) capacitor \
 c=0.0221661f //x=14.885 //y=0.375 //x2=17.445 //y2=0.995
cc_6138 ( N_noxref_34_M9_noxref_s N_noxref_35_c_10896_n ) capacitor \
 c=0.0180035f //x=14.885 //y=0.375 //x2=17.53 //y2=0.625
cc_6139 ( N_noxref_34_c_10852_n N_noxref_35_M10_noxref_d ) capacitor \
 c=0.0127191f //x=16.875 //y=0.54 //x2=16.29 //y2=0.91
cc_6140 ( N_noxref_34_c_10875_n N_noxref_35_M10_noxref_d ) capacitor \
 c=0.00861161f //x=16.875 //y=1.59 //x2=16.29 //y2=0.91
cc_6141 ( N_noxref_34_M9_noxref_s N_noxref_35_M10_noxref_d ) capacitor \
 c=0.0159202f //x=14.885 //y=0.375 //x2=16.29 //y2=0.91
cc_6142 ( N_noxref_34_M9_noxref_s N_noxref_35_M11_noxref_s ) capacitor \
 c=0.0213553f //x=14.885 //y=0.375 //x2=17.395 //y2=0.375
cc_6143 ( N_noxref_35_c_10901_n N_noxref_36_M12_noxref_s ) capacitor \
 c=0.00191848f //x=18.5 //y=0.625 //x2=19.695 //y2=0.375
cc_6144 ( N_noxref_36_c_10954_n N_noxref_37_c_10999_n ) capacitor c=0.0131801f \
 //x=21.685 //y=0.54 //x2=22.255 //y2=0.995
cc_6145 ( N_noxref_36_c_10979_n N_noxref_37_c_10999_n ) capacitor \
 c=0.00980353f //x=21.685 //y=1.59 //x2=22.255 //y2=0.995
cc_6146 ( N_noxref_36_M12_noxref_s N_noxref_37_c_10999_n ) capacitor \
 c=0.0221661f //x=19.695 //y=0.375 //x2=22.255 //y2=0.995
cc_6147 ( N_noxref_36_M12_noxref_s N_noxref_37_c_11001_n ) capacitor \
 c=0.0180035f //x=19.695 //y=0.375 //x2=22.34 //y2=0.625
cc_6148 ( N_noxref_36_c_10954_n N_noxref_37_M13_noxref_d ) capacitor \
 c=0.0127176f //x=21.685 //y=0.54 //x2=21.1 //y2=0.91
cc_6149 ( N_noxref_36_c_10979_n N_noxref_37_M13_noxref_d ) capacitor \
 c=0.0086073f //x=21.685 //y=1.59 //x2=21.1 //y2=0.91
cc_6150 ( N_noxref_36_M12_noxref_s N_noxref_37_M13_noxref_d ) capacitor \
 c=0.0159202f //x=19.695 //y=0.375 //x2=21.1 //y2=0.91
cc_6151 ( N_noxref_36_M12_noxref_s N_noxref_37_M14_noxref_s ) capacitor \
 c=0.0213553f //x=19.695 //y=0.375 //x2=22.205 //y2=0.375
cc_6152 ( N_noxref_37_c_11006_n N_noxref_38_M15_noxref_s ) capacitor \
 c=0.00191848f //x=23.31 //y=0.625 //x2=24.505 //y2=0.375
cc_6153 ( N_noxref_38_c_11058_n N_noxref_39_c_11100_n ) capacitor c=0.0131877f \
 //x=26.495 //y=0.54 //x2=27.065 //y2=0.995
cc_6154 ( N_noxref_38_c_11081_n N_noxref_39_c_11100_n ) capacitor \
 c=0.00981707f //x=26.495 //y=1.59 //x2=27.065 //y2=0.995
cc_6155 ( N_noxref_38_M15_noxref_s N_noxref_39_c_11100_n ) capacitor \
 c=0.0221661f //x=24.505 //y=0.375 //x2=27.065 //y2=0.995
cc_6156 ( N_noxref_38_M15_noxref_s N_noxref_39_c_11102_n ) capacitor \
 c=0.0180035f //x=24.505 //y=0.375 //x2=27.15 //y2=0.625
cc_6157 ( N_noxref_38_c_11058_n N_noxref_39_M16_noxref_d ) capacitor \
 c=0.0127191f //x=26.495 //y=0.54 //x2=25.91 //y2=0.91
cc_6158 ( N_noxref_38_c_11081_n N_noxref_39_M16_noxref_d ) capacitor \
 c=0.00861161f //x=26.495 //y=1.59 //x2=25.91 //y2=0.91
cc_6159 ( N_noxref_38_M15_noxref_s N_noxref_39_M16_noxref_d ) capacitor \
 c=0.0159202f //x=24.505 //y=0.375 //x2=25.91 //y2=0.91
cc_6160 ( N_noxref_38_M15_noxref_s N_noxref_39_M17_noxref_s ) capacitor \
 c=0.0213553f //x=24.505 //y=0.375 //x2=27.015 //y2=0.375
cc_6161 ( N_noxref_39_c_11107_n N_noxref_40_M18_noxref_s ) capacitor \
 c=0.00191848f //x=28.12 //y=0.625 //x2=29.315 //y2=0.375
cc_6162 ( N_noxref_40_c_11159_n N_noxref_41_c_11204_n ) capacitor c=0.0131801f \
 //x=31.305 //y=0.54 //x2=31.875 //y2=0.995
cc_6163 ( N_noxref_40_c_11184_n N_noxref_41_c_11204_n ) capacitor \
 c=0.00980353f //x=31.305 //y=1.59 //x2=31.875 //y2=0.995
cc_6164 ( N_noxref_40_M18_noxref_s N_noxref_41_c_11204_n ) capacitor \
 c=0.0221661f //x=29.315 //y=0.375 //x2=31.875 //y2=0.995
cc_6165 ( N_noxref_40_M18_noxref_s N_noxref_41_c_11206_n ) capacitor \
 c=0.0180035f //x=29.315 //y=0.375 //x2=31.96 //y2=0.625
cc_6166 ( N_noxref_40_c_11159_n N_noxref_41_M19_noxref_d ) capacitor \
 c=0.0127176f //x=31.305 //y=0.54 //x2=30.72 //y2=0.91
cc_6167 ( N_noxref_40_c_11184_n N_noxref_41_M19_noxref_d ) capacitor \
 c=0.0086073f //x=31.305 //y=1.59 //x2=30.72 //y2=0.91
cc_6168 ( N_noxref_40_M18_noxref_s N_noxref_41_M19_noxref_d ) capacitor \
 c=0.0159202f //x=29.315 //y=0.375 //x2=30.72 //y2=0.91
cc_6169 ( N_noxref_40_M18_noxref_s N_noxref_41_M20_noxref_s ) capacitor \
 c=0.0213553f //x=29.315 //y=0.375 //x2=31.825 //y2=0.375
cc_6170 ( N_noxref_41_c_11211_n N_noxref_42_M21_noxref_s ) capacitor \
 c=0.00191848f //x=32.93 //y=0.625 //x2=34.125 //y2=0.375
cc_6171 ( N_noxref_42_c_11263_n N_noxref_43_c_11305_n ) capacitor c=0.0131877f \
 //x=36.115 //y=0.54 //x2=36.685 //y2=0.995
cc_6172 ( N_noxref_42_c_11286_n N_noxref_43_c_11305_n ) capacitor \
 c=0.00981707f //x=36.115 //y=1.59 //x2=36.685 //y2=0.995
cc_6173 ( N_noxref_42_M21_noxref_s N_noxref_43_c_11305_n ) capacitor \
 c=0.0221661f //x=34.125 //y=0.375 //x2=36.685 //y2=0.995
cc_6174 ( N_noxref_42_M21_noxref_s N_noxref_43_c_11307_n ) capacitor \
 c=0.0180035f //x=34.125 //y=0.375 //x2=36.77 //y2=0.625
cc_6175 ( N_noxref_42_c_11263_n N_noxref_43_M22_noxref_d ) capacitor \
 c=0.0127191f //x=36.115 //y=0.54 //x2=35.53 //y2=0.91
cc_6176 ( N_noxref_42_c_11286_n N_noxref_43_M22_noxref_d ) capacitor \
 c=0.00861161f //x=36.115 //y=1.59 //x2=35.53 //y2=0.91
cc_6177 ( N_noxref_42_M21_noxref_s N_noxref_43_M22_noxref_d ) capacitor \
 c=0.0159202f //x=34.125 //y=0.375 //x2=35.53 //y2=0.91
cc_6178 ( N_noxref_42_M21_noxref_s N_noxref_43_M23_noxref_s ) capacitor \
 c=0.0213553f //x=34.125 //y=0.375 //x2=36.635 //y2=0.375
cc_6179 ( N_noxref_43_c_11312_n N_noxref_44_M24_noxref_s ) capacitor \
 c=0.00191848f //x=37.74 //y=0.625 //x2=38.935 //y2=0.375
cc_6180 ( N_noxref_44_c_11364_n N_noxref_45_c_11406_n ) capacitor c=0.0131877f \
 //x=40.925 //y=0.54 //x2=41.495 //y2=0.995
cc_6181 ( N_noxref_44_c_11387_n N_noxref_45_c_11406_n ) capacitor \
 c=0.00981707f //x=40.925 //y=1.59 //x2=41.495 //y2=0.995
cc_6182 ( N_noxref_44_M24_noxref_s N_noxref_45_c_11406_n ) capacitor \
 c=0.0221661f //x=38.935 //y=0.375 //x2=41.495 //y2=0.995
cc_6183 ( N_noxref_44_M24_noxref_s N_noxref_45_c_11408_n ) capacitor \
 c=0.0180035f //x=38.935 //y=0.375 //x2=41.58 //y2=0.625
cc_6184 ( N_noxref_44_c_11364_n N_noxref_45_M25_noxref_d ) capacitor \
 c=0.0127191f //x=40.925 //y=0.54 //x2=40.34 //y2=0.91
cc_6185 ( N_noxref_44_c_11387_n N_noxref_45_M25_noxref_d ) capacitor \
 c=0.00861161f //x=40.925 //y=1.59 //x2=40.34 //y2=0.91
cc_6186 ( N_noxref_44_M24_noxref_s N_noxref_45_M25_noxref_d ) capacitor \
 c=0.0159202f //x=38.935 //y=0.375 //x2=40.34 //y2=0.91
cc_6187 ( N_noxref_44_M24_noxref_s N_noxref_45_M26_noxref_s ) capacitor \
 c=0.0213553f //x=38.935 //y=0.375 //x2=41.445 //y2=0.375
cc_6188 ( N_noxref_45_c_11413_n N_noxref_46_M27_noxref_s ) capacitor \
 c=0.00191848f //x=42.55 //y=0.625 //x2=43.745 //y2=0.375
cc_6189 ( N_noxref_46_c_11465_n N_noxref_47_c_11507_n ) capacitor c=0.0131877f \
 //x=45.735 //y=0.54 //x2=46.305 //y2=0.995
cc_6190 ( N_noxref_46_c_11488_n N_noxref_47_c_11507_n ) capacitor \
 c=0.00981707f //x=45.735 //y=1.59 //x2=46.305 //y2=0.995
cc_6191 ( N_noxref_46_M27_noxref_s N_noxref_47_c_11507_n ) capacitor \
 c=0.0221661f //x=43.745 //y=0.375 //x2=46.305 //y2=0.995
cc_6192 ( N_noxref_46_M27_noxref_s N_noxref_47_c_11509_n ) capacitor \
 c=0.0180035f //x=43.745 //y=0.375 //x2=46.39 //y2=0.625
cc_6193 ( N_noxref_46_c_11465_n N_noxref_47_M28_noxref_d ) capacitor \
 c=0.0127191f //x=45.735 //y=0.54 //x2=45.15 //y2=0.91
cc_6194 ( N_noxref_46_c_11488_n N_noxref_47_M28_noxref_d ) capacitor \
 c=0.00861161f //x=45.735 //y=1.59 //x2=45.15 //y2=0.91
cc_6195 ( N_noxref_46_M27_noxref_s N_noxref_47_M28_noxref_d ) capacitor \
 c=0.0159202f //x=43.745 //y=0.375 //x2=45.15 //y2=0.91
cc_6196 ( N_noxref_46_M27_noxref_s N_noxref_47_M29_noxref_s ) capacitor \
 c=0.0213553f //x=43.745 //y=0.375 //x2=46.255 //y2=0.375
cc_6197 ( N_noxref_47_c_11514_n N_noxref_48_M30_noxref_s ) capacitor \
 c=0.00191848f //x=47.36 //y=0.625 //x2=48.555 //y2=0.375
cc_6198 ( N_noxref_48_c_11567_n N_noxref_49_c_11612_n ) capacitor c=0.0131801f \
 //x=50.545 //y=0.54 //x2=51.115 //y2=0.995
cc_6199 ( N_noxref_48_c_11591_n N_noxref_49_c_11612_n ) capacitor \
 c=0.00980353f //x=50.545 //y=1.59 //x2=51.115 //y2=0.995
cc_6200 ( N_noxref_48_M30_noxref_s N_noxref_49_c_11612_n ) capacitor \
 c=0.0221661f //x=48.555 //y=0.375 //x2=51.115 //y2=0.995
cc_6201 ( N_noxref_48_M30_noxref_s N_noxref_49_c_11614_n ) capacitor \
 c=0.0180035f //x=48.555 //y=0.375 //x2=51.2 //y2=0.625
cc_6202 ( N_noxref_48_c_11567_n N_noxref_49_M31_noxref_d ) capacitor \
 c=0.0127176f //x=50.545 //y=0.54 //x2=49.96 //y2=0.91
cc_6203 ( N_noxref_48_c_11591_n N_noxref_49_M31_noxref_d ) capacitor \
 c=0.0086073f //x=50.545 //y=1.59 //x2=49.96 //y2=0.91
cc_6204 ( N_noxref_48_M30_noxref_s N_noxref_49_M31_noxref_d ) capacitor \
 c=0.0159202f //x=48.555 //y=0.375 //x2=49.96 //y2=0.91
cc_6205 ( N_noxref_48_M30_noxref_s N_noxref_49_M32_noxref_s ) capacitor \
 c=0.0213553f //x=48.555 //y=0.375 //x2=51.065 //y2=0.375
cc_6206 ( N_noxref_49_c_11619_n N_noxref_50_M33_noxref_s ) capacitor \
 c=0.00191848f //x=52.17 //y=0.625 //x2=53.365 //y2=0.375
cc_6207 ( N_noxref_50_c_11671_n N_noxref_51_c_11713_n ) capacitor c=0.0131877f \
 //x=55.355 //y=0.54 //x2=55.925 //y2=0.995
cc_6208 ( N_noxref_50_c_11682_n N_noxref_51_c_11713_n ) capacitor \
 c=0.00981707f //x=55.355 //y=1.59 //x2=55.925 //y2=0.995
cc_6209 ( N_noxref_50_M33_noxref_s N_noxref_51_c_11713_n ) capacitor \
 c=0.0221661f //x=53.365 //y=0.375 //x2=55.925 //y2=0.995
cc_6210 ( N_noxref_50_M33_noxref_s N_noxref_51_c_11715_n ) capacitor \
 c=0.0180035f //x=53.365 //y=0.375 //x2=56.01 //y2=0.625
cc_6211 ( N_noxref_50_c_11671_n N_noxref_51_M34_noxref_d ) capacitor \
 c=0.0127191f //x=55.355 //y=0.54 //x2=54.77 //y2=0.91
cc_6212 ( N_noxref_50_c_11682_n N_noxref_51_M34_noxref_d ) capacitor \
 c=0.00861161f //x=55.355 //y=1.59 //x2=54.77 //y2=0.91
cc_6213 ( N_noxref_50_M33_noxref_s N_noxref_51_M34_noxref_d ) capacitor \
 c=0.0159202f //x=53.365 //y=0.375 //x2=54.77 //y2=0.91
cc_6214 ( N_noxref_50_M33_noxref_s N_noxref_51_M35_noxref_s ) capacitor \
 c=0.0213553f //x=53.365 //y=0.375 //x2=55.875 //y2=0.375
cc_6215 ( N_noxref_51_c_11720_n N_noxref_52_M36_noxref_s ) capacitor \
 c=0.00191848f //x=56.98 //y=0.625 //x2=58.175 //y2=0.375
cc_6216 ( N_noxref_52_c_11772_n N_noxref_53_c_11817_n ) capacitor c=0.0131801f \
 //x=60.165 //y=0.54 //x2=60.735 //y2=0.995
cc_6217 ( N_noxref_52_c_11797_n N_noxref_53_c_11817_n ) capacitor \
 c=0.00980353f //x=60.165 //y=1.59 //x2=60.735 //y2=0.995
cc_6218 ( N_noxref_52_M36_noxref_s N_noxref_53_c_11817_n ) capacitor \
 c=0.0221661f //x=58.175 //y=0.375 //x2=60.735 //y2=0.995
cc_6219 ( N_noxref_52_M36_noxref_s N_noxref_53_c_11819_n ) capacitor \
 c=0.0180035f //x=58.175 //y=0.375 //x2=60.82 //y2=0.625
cc_6220 ( N_noxref_52_c_11772_n N_noxref_53_M37_noxref_d ) capacitor \
 c=0.0127176f //x=60.165 //y=0.54 //x2=59.58 //y2=0.91
cc_6221 ( N_noxref_52_c_11797_n N_noxref_53_M37_noxref_d ) capacitor \
 c=0.0086073f //x=60.165 //y=1.59 //x2=59.58 //y2=0.91
cc_6222 ( N_noxref_52_M36_noxref_s N_noxref_53_M37_noxref_d ) capacitor \
 c=0.0159202f //x=58.175 //y=0.375 //x2=59.58 //y2=0.91
cc_6223 ( N_noxref_52_M36_noxref_s N_noxref_53_M38_noxref_s ) capacitor \
 c=0.0213553f //x=58.175 //y=0.375 //x2=60.685 //y2=0.375
cc_6224 ( N_noxref_53_c_11824_n N_noxref_54_M39_noxref_s ) capacitor \
 c=0.00191848f //x=61.79 //y=0.625 //x2=62.985 //y2=0.375
cc_6225 ( N_noxref_54_c_11876_n N_noxref_55_c_11918_n ) capacitor c=0.0131877f \
 //x=64.975 //y=0.54 //x2=65.545 //y2=0.995
cc_6226 ( N_noxref_54_c_11898_n N_noxref_55_c_11918_n ) capacitor \
 c=0.00981707f //x=64.975 //y=1.59 //x2=65.545 //y2=0.995
cc_6227 ( N_noxref_54_M39_noxref_s N_noxref_55_c_11918_n ) capacitor \
 c=0.0221661f //x=62.985 //y=0.375 //x2=65.545 //y2=0.995
cc_6228 ( N_noxref_54_M39_noxref_s N_noxref_55_c_11920_n ) capacitor \
 c=0.0180035f //x=62.985 //y=0.375 //x2=65.63 //y2=0.625
cc_6229 ( N_noxref_54_c_11876_n N_noxref_55_M40_noxref_d ) capacitor \
 c=0.0127191f //x=64.975 //y=0.54 //x2=64.39 //y2=0.91
cc_6230 ( N_noxref_54_c_11898_n N_noxref_55_M40_noxref_d ) capacitor \
 c=0.00861161f //x=64.975 //y=1.59 //x2=64.39 //y2=0.91
cc_6231 ( N_noxref_54_M39_noxref_s N_noxref_55_M40_noxref_d ) capacitor \
 c=0.0159202f //x=62.985 //y=0.375 //x2=64.39 //y2=0.91
cc_6232 ( N_noxref_54_M39_noxref_s N_noxref_55_M41_noxref_s ) capacitor \
 c=0.0213553f //x=62.985 //y=0.375 //x2=65.495 //y2=0.375
cc_6233 ( N_noxref_55_c_11925_n N_noxref_56_M42_noxref_s ) capacitor \
 c=0.00191848f //x=66.6 //y=0.625 //x2=67.795 //y2=0.375
cc_6234 ( N_noxref_56_c_11977_n N_noxref_57_c_12019_n ) capacitor c=0.0131877f \
 //x=69.785 //y=0.54 //x2=70.355 //y2=0.995
cc_6235 ( N_noxref_56_c_12000_n N_noxref_57_c_12019_n ) capacitor \
 c=0.00981707f //x=69.785 //y=1.59 //x2=70.355 //y2=0.995
cc_6236 ( N_noxref_56_M42_noxref_s N_noxref_57_c_12019_n ) capacitor \
 c=0.0221661f //x=67.795 //y=0.375 //x2=70.355 //y2=0.995
cc_6237 ( N_noxref_56_M42_noxref_s N_noxref_57_c_12021_n ) capacitor \
 c=0.0180035f //x=67.795 //y=0.375 //x2=70.44 //y2=0.625
cc_6238 ( N_noxref_56_c_11977_n N_noxref_57_M43_noxref_d ) capacitor \
 c=0.0127191f //x=69.785 //y=0.54 //x2=69.2 //y2=0.91
cc_6239 ( N_noxref_56_c_12000_n N_noxref_57_M43_noxref_d ) capacitor \
 c=0.00861161f //x=69.785 //y=1.59 //x2=69.2 //y2=0.91
cc_6240 ( N_noxref_56_M42_noxref_s N_noxref_57_M43_noxref_d ) capacitor \
 c=0.0159202f //x=67.795 //y=0.375 //x2=69.2 //y2=0.91
cc_6241 ( N_noxref_56_M42_noxref_s N_noxref_57_M44_noxref_s ) capacitor \
 c=0.0213553f //x=67.795 //y=0.375 //x2=70.305 //y2=0.375
cc_6242 ( N_noxref_57_c_12026_n N_noxref_58_M45_noxref_s ) capacitor \
 c=0.00191848f //x=71.41 //y=0.625 //x2=72.605 //y2=0.375
cc_6243 ( N_noxref_58_c_12078_n N_noxref_59_c_12120_n ) capacitor c=0.0131877f \
 //x=74.595 //y=0.54 //x2=75.165 //y2=0.995
cc_6244 ( N_noxref_58_c_12100_n N_noxref_59_c_12120_n ) capacitor \
 c=0.00981707f //x=74.595 //y=1.59 //x2=75.165 //y2=0.995
cc_6245 ( N_noxref_58_M45_noxref_s N_noxref_59_c_12120_n ) capacitor \
 c=0.0221661f //x=72.605 //y=0.375 //x2=75.165 //y2=0.995
cc_6246 ( N_noxref_58_M45_noxref_s N_noxref_59_c_12122_n ) capacitor \
 c=0.0180035f //x=72.605 //y=0.375 //x2=75.25 //y2=0.625
cc_6247 ( N_noxref_58_c_12078_n N_noxref_59_M46_noxref_d ) capacitor \
 c=0.0127191f //x=74.595 //y=0.54 //x2=74.01 //y2=0.91
cc_6248 ( N_noxref_58_c_12100_n N_noxref_59_M46_noxref_d ) capacitor \
 c=0.00861161f //x=74.595 //y=1.59 //x2=74.01 //y2=0.91
cc_6249 ( N_noxref_58_M45_noxref_s N_noxref_59_M46_noxref_d ) capacitor \
 c=0.0159202f //x=72.605 //y=0.375 //x2=74.01 //y2=0.91
cc_6250 ( N_noxref_58_M45_noxref_s N_noxref_59_M47_noxref_s ) capacitor \
 c=0.0213553f //x=72.605 //y=0.375 //x2=75.115 //y2=0.375
cc_6251 ( N_noxref_59_c_12127_n N_noxref_60_M48_noxref_s ) capacitor \
 c=0.00191848f //x=76.22 //y=0.625 //x2=77.415 //y2=0.375
cc_6252 ( N_noxref_60_c_12180_n N_noxref_61_c_12224_n ) capacitor c=0.0132328f \
 //x=79.405 //y=0.54 //x2=79.975 //y2=0.995
cc_6253 ( N_noxref_60_c_12202_n N_noxref_61_c_12224_n ) capacitor \
 c=0.00988406f //x=79.405 //y=1.59 //x2=79.975 //y2=0.995
cc_6254 ( N_noxref_60_M48_noxref_s N_noxref_61_c_12224_n ) capacitor \
 c=0.0226274f //x=77.415 //y=0.375 //x2=79.975 //y2=0.995
cc_6255 ( N_noxref_60_M48_noxref_s N_noxref_61_c_12226_n ) capacitor \
 c=0.0180035f //x=77.415 //y=0.375 //x2=80.06 //y2=0.625
cc_6256 ( N_noxref_60_c_12180_n N_noxref_61_M49_noxref_d ) capacitor \
 c=0.0127176f //x=79.405 //y=0.54 //x2=78.82 //y2=0.91
cc_6257 ( N_noxref_60_c_12202_n N_noxref_61_M49_noxref_d ) capacitor \
 c=0.0086073f //x=79.405 //y=1.59 //x2=78.82 //y2=0.91
cc_6258 ( N_noxref_60_M48_noxref_s N_noxref_61_M49_noxref_d ) capacitor \
 c=0.0159202f //x=77.415 //y=0.375 //x2=78.82 //y2=0.91
cc_6259 ( N_noxref_60_M48_noxref_s N_noxref_61_M50_noxref_s ) capacitor \
 c=0.0213553f //x=77.415 //y=0.375 //x2=79.925 //y2=0.375
cc_6260 ( N_noxref_61_c_12231_n N_noxref_62_M51_noxref_s ) capacitor \
 c=0.00191848f //x=81.03 //y=0.625 //x2=82.225 //y2=0.375
cc_6261 ( N_noxref_62_c_12285_n N_noxref_63_c_12329_n ) capacitor c=0.0131877f \
 //x=84.215 //y=0.54 //x2=84.785 //y2=0.995
cc_6262 ( N_noxref_62_c_12295_n N_noxref_63_c_12329_n ) capacitor \
 c=0.00981707f //x=84.215 //y=1.59 //x2=84.785 //y2=0.995
cc_6263 ( N_noxref_62_M51_noxref_s N_noxref_63_c_12329_n ) capacitor \
 c=0.0221661f //x=82.225 //y=0.375 //x2=84.785 //y2=0.995
cc_6264 ( N_noxref_62_M51_noxref_s N_noxref_63_c_12331_n ) capacitor \
 c=0.0180035f //x=82.225 //y=0.375 //x2=84.87 //y2=0.625
cc_6265 ( N_noxref_62_c_12285_n N_noxref_63_M52_noxref_d ) capacitor \
 c=0.0127191f //x=84.215 //y=0.54 //x2=83.63 //y2=0.91
cc_6266 ( N_noxref_62_c_12295_n N_noxref_63_M52_noxref_d ) capacitor \
 c=0.00861161f //x=84.215 //y=1.59 //x2=83.63 //y2=0.91
cc_6267 ( N_noxref_62_M51_noxref_s N_noxref_63_M52_noxref_d ) capacitor \
 c=0.0159202f //x=82.225 //y=0.375 //x2=83.63 //y2=0.91
cc_6268 ( N_noxref_62_M51_noxref_s N_noxref_63_M53_noxref_s ) capacitor \
 c=0.0213553f //x=82.225 //y=0.375 //x2=84.735 //y2=0.375
cc_6269 ( N_noxref_63_c_12336_n N_noxref_64_M54_noxref_s ) capacitor \
 c=0.00195059f //x=85.84 //y=0.625 //x2=87.14 //y2=0.365
cc_6270 ( N_noxref_64_M54_noxref_s N_noxref_65_c_12455_n ) capacitor \
 c=0.0011299f //x=87.14 //y=0.365 //x2=90.605 //y2=1.495
cc_6271 ( N_noxref_64_c_12391_n N_noxref_65_M56_noxref_s ) capacitor \
 c=0.0011299f //x=89.215 //y=0.615 //x2=90.47 //y2=0.365
cc_6272 ( N_noxref_65_M56_noxref_s N_noxref_66_c_12509_n ) capacitor \
 c=0.0011299f //x=90.47 //y=0.365 //x2=93.935 //y2=1.495
cc_6273 ( N_noxref_65_c_12447_n N_noxref_66_M58_noxref_s ) capacitor \
 c=0.0011299f //x=92.545 //y=0.615 //x2=93.8 //y2=0.365
