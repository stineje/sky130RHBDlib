magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -66 377 1122 897
<< pwell >>
rect 4 43 914 283
rect -26 -43 1082 43
<< locali >>
rect 25 99 76 751
rect 284 355 430 411
rect 396 314 430 355
rect 466 350 551 424
rect 591 316 650 424
rect 697 316 839 382
rect 396 280 555 314
rect 910 280 976 403
rect 521 246 976 280
rect 607 242 742 246
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 112 735 650 751
rect 146 701 184 735
rect 218 701 256 735
rect 290 701 328 735
rect 362 701 400 735
rect 434 701 472 735
rect 506 701 544 735
rect 578 701 616 735
rect 112 530 650 701
rect 686 494 736 751
rect 117 460 736 494
rect 117 319 183 460
rect 686 435 736 460
rect 772 735 1034 747
rect 772 701 778 735
rect 812 701 850 735
rect 884 701 922 735
rect 956 701 994 735
rect 1028 701 1034 735
rect 772 439 1034 701
rect 117 285 360 319
rect 112 113 290 249
rect 326 244 360 285
rect 326 210 485 244
rect 451 176 571 210
rect 146 79 184 113
rect 218 79 256 113
rect 112 73 290 79
rect 349 87 415 174
rect 505 123 571 176
rect 670 87 736 206
rect 349 53 736 87
rect 778 113 1038 210
rect 778 79 783 113
rect 817 79 855 113
rect 889 79 927 113
rect 961 79 999 113
rect 1033 79 1038 113
rect 778 73 1038 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 112 701 146 735
rect 184 701 218 735
rect 256 701 290 735
rect 328 701 362 735
rect 400 701 434 735
rect 472 701 506 735
rect 544 701 578 735
rect 616 701 650 735
rect 778 701 812 735
rect 850 701 884 735
rect 922 701 956 735
rect 994 701 1028 735
rect 112 79 146 113
rect 184 79 218 113
rect 256 79 290 113
rect 783 79 817 113
rect 855 79 889 113
rect 927 79 961 113
rect 999 79 1033 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 831 1056 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 0 791 1056 797
rect 0 735 1056 763
rect 0 701 112 735
rect 146 701 184 735
rect 218 701 256 735
rect 290 701 328 735
rect 362 701 400 735
rect 434 701 472 735
rect 506 701 544 735
rect 578 701 616 735
rect 650 701 778 735
rect 812 701 850 735
rect 884 701 922 735
rect 956 701 994 735
rect 1028 701 1056 735
rect 0 689 1056 701
rect 0 113 1056 125
rect 0 79 112 113
rect 146 79 184 113
rect 218 79 256 113
rect 290 79 783 113
rect 817 79 855 113
rect 889 79 927 113
rect 961 79 999 113
rect 1033 79 1056 113
rect 0 51 1056 79
rect 0 17 1056 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -23 1056 -17
<< labels >>
rlabel locali s 607 242 742 246 6 A1
port 1 nsew signal input
rlabel locali s 521 246 976 280 6 A1
port 1 nsew signal input
rlabel locali s 910 280 976 403 6 A1
port 1 nsew signal input
rlabel locali s 396 280 555 314 6 A1
port 1 nsew signal input
rlabel locali s 396 314 430 355 6 A1
port 1 nsew signal input
rlabel locali s 284 355 430 411 6 A1
port 1 nsew signal input
rlabel locali s 697 316 839 382 6 A2
port 2 nsew signal input
rlabel locali s 466 350 551 424 6 B1
port 3 nsew signal input
rlabel locali s 591 316 650 424 6 B2
port 4 nsew signal input
rlabel metal1 s 0 51 1056 125 6 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 -23 1056 23 8 VNB
port 6 nsew ground bidirectional
rlabel pwell s -26 -43 1082 43 8 VNB
port 6 nsew ground bidirectional
rlabel pwell s 4 43 914 283 6 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 791 1056 837 6 VPB
port 7 nsew power bidirectional
rlabel nwell s -66 377 1122 897 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 689 1056 763 6 VPWR
port 8 nsew power bidirectional
rlabel locali s 25 99 76 751 6 X
port 9 nsew signal output
<< properties >>
string LEFsite unithv
string LEFclass CORE
string FIXED_BBOX 0 0 1056 814
string LEFsymmetry X Y
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_END 398928
string GDS_START 386192
<< end >>
