* SPICE3 file created from VOTERN3X1.ext - technology: sky130A

.subckt VOTERN3X1 YN A B C VDD GND
M1000 a_217_1051.t5 B.t0 a_881_1051.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_881_1051.t7 A.t0 YN.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 GND B.t1 a_778_101.t0 nshort w=-1.605u l=1.765u
+  ad=0.5373p pd=4.71u as=0p ps=0u
M1003 a_217_1051.t3 A.t1 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_217_1051.t2 C.t0 a_881_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 YN.t4 C.t1 a_881_1051.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 GND B.t2 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1007 GND C.t2 a_1444_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1008 YN A.t2 a_1444_101.t0 nshort w=-1.83u l=2.06u
+  ad=0.5373p pd=4.72u as=0p ps=0u
M1009 YN A.t4 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1010 VDD.t3 B.t3 a_217_1051.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 YN.t0 A.t3 a_881_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 YN C.t5 a_778_101.t0 nshort w=-1.235u l=1.535u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_881_1051.t1 C.t3 a_217_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t0 A.t5 a_217_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_881_1051.t4 C.t4 YN.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_881_1051.t5 B.t4 a_217_1051.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_217_1051.t7 B.t5 VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 B A 0.96fF
C1 B YN 0.05fF
C2 B VDD 0.28fF
C3 B C 0.15fF
C4 A YN 0.30fF
C5 A VDD 0.85fF
C6 C A 0.26fF
C7 YN VDD 0.29fF
C8 C YN 0.27fF
C9 C VDD 0.18fF
R0 B.n2 B.t3 512.525
R1 B.n0 B.t0 477.179
R2 B.n0 B.t4 406.485
R3 B.n2 B.t5 371.139
R4 B.n1 B.t1 363.924
R5 B.n3 B.t2 357.498
R6 B.n3 B.n2 71.88
R7 B.n4 B.n1 52.017
R8 B.n4 B.n3 49.342
R9 B.n1 B.n0 15.776
R10 B.n4 B 0.046
R11 a_881_1051.n3 a_881_1051.n2 196.002
R12 a_881_1051.n4 a_881_1051.t7 89.553
R13 a_881_1051.n2 a_881_1051.n1 75.271
R14 a_881_1051.n4 a_881_1051.n3 75.214
R15 a_881_1051.n2 a_881_1051.n0 36.52
R16 a_881_1051.n3 a_881_1051.t3 14.338
R17 a_881_1051.n0 a_881_1051.t2 14.282
R18 a_881_1051.n0 a_881_1051.t1 14.282
R19 a_881_1051.n1 a_881_1051.t6 14.282
R20 a_881_1051.n1 a_881_1051.t5 14.282
R21 a_881_1051.t0 a_881_1051.n5 14.282
R22 a_881_1051.n5 a_881_1051.t4 14.282
R23 a_881_1051.n5 a_881_1051.n4 12.122
R24 a_217_1051.n3 a_217_1051.n2 195.987
R25 a_217_1051.n4 a_217_1051.t2 89.553
R26 a_217_1051.n2 a_217_1051.n1 75.271
R27 a_217_1051.n4 a_217_1051.n3 75.214
R28 a_217_1051.n2 a_217_1051.n0 36.519
R29 a_217_1051.n3 a_217_1051.t4 14.338
R30 a_217_1051.n0 a_217_1051.t0 14.282
R31 a_217_1051.n0 a_217_1051.t3 14.282
R32 a_217_1051.n1 a_217_1051.t6 14.282
R33 a_217_1051.n1 a_217_1051.t7 14.282
R34 a_217_1051.n5 a_217_1051.t1 14.282
R35 a_217_1051.t5 a_217_1051.n5 14.282
R36 a_217_1051.n5 a_217_1051.n4 12.122
R37 A.n0 A.t0 475.572
R38 A.n2 A.t5 469.145
R39 A.n2 A.t1 384.527
R40 A.n0 A.t3 384.527
R41 A.n3 A.t4 294.278
R42 A.n1 A.t2 294.278
R43 A.n4 A.n1 80.851
R44 A.n4 A.n3 76
R45 A.n1 A.n0 57.842
R46 A.n3 A.n2 56.833
R47 A.n4 A 0.046
R48 YN.n15 YN.n14 216.728
R49 YN.n15 YN.n2 126.664
R50 YN.n10 YN.n5 111.94
R51 YN.n10 YN.n9 98.501
R52 YN.n13 YN.n11 80.526
R53 YN.n14 YN.n10 78.403
R54 YN.n16 YN.n15 76
R55 YN.n2 YN.n1 75.271
R56 YN.n9 YN.n8 30
R57 YN.n13 YN.n12 30
R58 YN.n7 YN.n6 24.383
R59 YN.n9 YN.n7 23.684
R60 YN.n5 YN.n4 22.578
R61 YN.n14 YN.n13 20.417
R62 YN.n0 YN.t1 14.282
R63 YN.n0 YN.t0 14.282
R64 YN.n1 YN.t5 14.282
R65 YN.n1 YN.t4 14.282
R66 YN.n2 YN.n0 12.119
R67 YN.n5 YN.n3 8.58
R68 YN.n16 YN 0.046
R69 VDD.n76 VDD.n74 144.705
R70 VDD.n173 VDD.n171 144.705
R71 VDD.n39 VDD.n38 76
R72 VDD.n43 VDD.n42 76
R73 VDD.n47 VDD.n46 76
R74 VDD.n51 VDD.n50 76
R75 VDD.n78 VDD.n77 76
R76 VDD.n82 VDD.n81 76
R77 VDD.n86 VDD.n85 76
R78 VDD.n90 VDD.n89 76
R79 VDD.n187 VDD.n186 76
R80 VDD.n183 VDD.n182 76
R81 VDD.n179 VDD.n178 76
R82 VDD.n175 VDD.n174 76
R83 VDD.n148 VDD.n147 76
R84 VDD.n144 VDD.n143 76
R85 VDD.n139 VDD.n138 76
R86 VDD.n134 VDD.n133 76
R87 VDD.n128 VDD.n127 76
R88 VDD.n123 VDD.n122 76
R89 VDD.n118 VDD.n117 76
R90 VDD.n113 VDD.n112 76
R91 VDD.n114 VDD.t2 55.465
R92 VDD.n140 VDD.t0 55.465
R93 VDD.n130 VDD.n129 41.183
R94 VDD.n56 VDD.n55 36.774
R95 VDD.n164 VDD.n163 36.774
R96 VDD.n136 VDD.n135 36.608
R97 VDD.n34 VDD.n33 34.942
R98 VDD.n120 VDD.n119 32.032
R99 VDD.n112 VDD.n109 21.841
R100 VDD.n23 VDD.n20 21.841
R101 VDD.n129 VDD.t1 14.282
R102 VDD.n129 VDD.t3 14.282
R103 VDD.n109 VDD.n92 14.167
R104 VDD.n92 VDD.n91 14.167
R105 VDD.n72 VDD.n53 14.167
R106 VDD.n53 VDD.n52 14.167
R107 VDD.n169 VDD.n150 14.167
R108 VDD.n150 VDD.n149 14.167
R109 VDD.n20 VDD.n19 14.167
R110 VDD.n19 VDD.n17 14.167
R111 VDD.n32 VDD.n29 14.167
R112 VDD.n29 VDD.n28 14.167
R113 VDD.n77 VDD.n73 14.167
R114 VDD.n174 VDD.n170 14.167
R115 VDD.n23 VDD.n22 13.653
R116 VDD.n22 VDD.n21 13.653
R117 VDD.n32 VDD.n31 13.653
R118 VDD.n31 VDD.n30 13.653
R119 VDD.n29 VDD.n25 13.653
R120 VDD.n25 VDD.n24 13.653
R121 VDD.n28 VDD.n27 13.653
R122 VDD.n27 VDD.n26 13.653
R123 VDD.n38 VDD.n37 13.653
R124 VDD.n37 VDD.n36 13.653
R125 VDD.n42 VDD.n41 13.653
R126 VDD.n41 VDD.n40 13.653
R127 VDD.n46 VDD.n45 13.653
R128 VDD.n45 VDD.n44 13.653
R129 VDD.n50 VDD.n49 13.653
R130 VDD.n49 VDD.n48 13.653
R131 VDD.n77 VDD.n76 13.653
R132 VDD.n76 VDD.n75 13.653
R133 VDD.n81 VDD.n80 13.653
R134 VDD.n80 VDD.n79 13.653
R135 VDD.n85 VDD.n84 13.653
R136 VDD.n84 VDD.n83 13.653
R137 VDD.n89 VDD.n88 13.653
R138 VDD.n88 VDD.n87 13.653
R139 VDD.n186 VDD.n185 13.653
R140 VDD.n185 VDD.n184 13.653
R141 VDD.n182 VDD.n181 13.653
R142 VDD.n181 VDD.n180 13.653
R143 VDD.n178 VDD.n177 13.653
R144 VDD.n177 VDD.n176 13.653
R145 VDD.n174 VDD.n173 13.653
R146 VDD.n173 VDD.n172 13.653
R147 VDD.n147 VDD.n146 13.653
R148 VDD.n146 VDD.n145 13.653
R149 VDD.n143 VDD.n142 13.653
R150 VDD.n142 VDD.n141 13.653
R151 VDD.n138 VDD.n137 13.653
R152 VDD.n137 VDD.n136 13.653
R153 VDD.n133 VDD.n132 13.653
R154 VDD.n132 VDD.n131 13.653
R155 VDD.n127 VDD.n126 13.653
R156 VDD.n126 VDD.n125 13.653
R157 VDD.n122 VDD.n121 13.653
R158 VDD.n121 VDD.n120 13.653
R159 VDD.n117 VDD.n116 13.653
R160 VDD.n116 VDD.n115 13.653
R161 VDD.n112 VDD.n111 13.653
R162 VDD.n111 VDD.n110 13.653
R163 VDD.n4 VDD.n2 12.915
R164 VDD.n4 VDD.n3 12.66
R165 VDD.n12 VDD.n11 12.343
R166 VDD.n12 VDD.n9 12.343
R167 VDD.n7 VDD.n6 12.343
R168 VDD.n133 VDD.n130 8.658
R169 VDD.n73 VDD.n72 7.674
R170 VDD.n170 VDD.n169 7.674
R171 VDD.n67 VDD.n66 7.5
R172 VDD.n61 VDD.n60 7.5
R173 VDD.n63 VDD.n62 7.5
R174 VDD.n58 VDD.n57 7.5
R175 VDD.n72 VDD.n71 7.5
R176 VDD.n154 VDD.n153 7.5
R177 VDD.n157 VDD.n156 7.5
R178 VDD.n159 VDD.n158 7.5
R179 VDD.n162 VDD.n161 7.5
R180 VDD.n169 VDD.n168 7.5
R181 VDD.n104 VDD.n103 7.5
R182 VDD.n98 VDD.n97 7.5
R183 VDD.n100 VDD.n99 7.5
R184 VDD.n106 VDD.n96 7.5
R185 VDD.n106 VDD.n94 7.5
R186 VDD.n109 VDD.n108 7.5
R187 VDD.n20 VDD.n16 7.5
R188 VDD.n2 VDD.n1 7.5
R189 VDD.n6 VDD.n5 7.5
R190 VDD.n11 VDD.n10 7.5
R191 VDD.n19 VDD.n18 7.5
R192 VDD.n14 VDD.n0 7.5
R193 VDD.n59 VDD.n56 6.772
R194 VDD.n70 VDD.n54 6.772
R195 VDD.n68 VDD.n65 6.772
R196 VDD.n64 VDD.n61 6.772
R197 VDD.n107 VDD.n93 6.772
R198 VDD.n105 VDD.n102 6.772
R199 VDD.n101 VDD.n98 6.772
R200 VDD.n59 VDD.n58 6.772
R201 VDD.n64 VDD.n63 6.772
R202 VDD.n68 VDD.n67 6.772
R203 VDD.n71 VDD.n70 6.772
R204 VDD.n101 VDD.n100 6.772
R205 VDD.n105 VDD.n104 6.772
R206 VDD.n108 VDD.n107 6.772
R207 VDD.n168 VDD.n167 6.772
R208 VDD.n155 VDD.n152 6.772
R209 VDD.n160 VDD.n157 6.772
R210 VDD.n165 VDD.n162 6.772
R211 VDD.n165 VDD.n164 6.772
R212 VDD.n160 VDD.n159 6.772
R213 VDD.n155 VDD.n154 6.772
R214 VDD.n167 VDD.n151 6.772
R215 VDD.n33 VDD.n23 6.487
R216 VDD.n33 VDD.n32 6.475
R217 VDD.n16 VDD.n15 6.458
R218 VDD.n96 VDD.n95 6.202
R219 VDD.n125 VDD.n124 4.576
R220 VDD.n117 VDD.n114 2.754
R221 VDD.n143 VDD.n140 2.361
R222 VDD.n14 VDD.n7 1.329
R223 VDD.n14 VDD.n8 1.329
R224 VDD.n14 VDD.n12 1.329
R225 VDD.n14 VDD.n13 1.329
R226 VDD.n15 VDD.n14 0.696
R227 VDD.n14 VDD.n4 0.696
R228 VDD.n69 VDD.n68 0.365
R229 VDD.n69 VDD.n64 0.365
R230 VDD.n69 VDD.n59 0.365
R231 VDD.n70 VDD.n69 0.365
R232 VDD.n106 VDD.n105 0.365
R233 VDD.n106 VDD.n101 0.365
R234 VDD.n107 VDD.n106 0.365
R235 VDD.n166 VDD.n165 0.365
R236 VDD.n166 VDD.n160 0.365
R237 VDD.n166 VDD.n155 0.365
R238 VDD.n167 VDD.n166 0.365
R239 VDD.n78 VDD.n51 0.29
R240 VDD.n175 VDD.n148 0.29
R241 VDD.n113 VDD 0.207
R242 VDD.n39 VDD.n35 0.181
R243 VDD.n134 VDD.n128 0.181
R244 VDD.n35 VDD.n34 0.145
R245 VDD.n43 VDD.n39 0.145
R246 VDD.n47 VDD.n43 0.145
R247 VDD.n51 VDD.n47 0.145
R248 VDD.n82 VDD.n78 0.145
R249 VDD.n86 VDD.n82 0.145
R250 VDD.n90 VDD.n86 0.145
R251 VDD.n187 VDD.n183 0.145
R252 VDD.n183 VDD.n179 0.145
R253 VDD.n179 VDD.n175 0.145
R254 VDD.n148 VDD.n144 0.145
R255 VDD.n144 VDD.n139 0.145
R256 VDD.n139 VDD.n134 0.145
R257 VDD.n128 VDD.n123 0.145
R258 VDD.n123 VDD.n118 0.145
R259 VDD.n118 VDD.n113 0.145
R260 VDD VDD.n90 0.09
R261 VDD VDD.n187 0.09
R262 C.n2 C.t3 512.525
R263 C.n0 C.t4 512.525
R264 C.n2 C.t0 371.139
R265 C.n0 C.t1 371.139
R266 C.n3 C.n2 265.439
R267 C.n1 C.n0 265.439
R268 C.n1 C.t2 176.995
R269 C.n3 C.t5 170.569
R270 C.n4 C.n1 77.043
R271 C.n4 C.n3 76
R272 C.n4 C 0.046
R273 a_778_101.t0 a_778_101.n0 93.333
R274 a_778_101.n3 a_778_101.n1 55.048
R275 a_778_101.n3 a_778_101.n2 2.097
R276 a_778_101.t0 a_778_101.n3 0.11
R277 GND.n29 GND.n27 219.745
R278 GND.n75 GND.n74 219.745
R279 GND.n29 GND.n28 85.529
R280 GND.n75 GND.n73 85.529
R281 GND.n83 GND.n82 84.842
R282 GND.n45 GND.n44 76
R283 GND.n42 GND.n41 76
R284 GND.n89 GND.n88 76
R285 GND.n86 GND.n85 76
R286 GND.n81 GND.n80 76
R287 GND.n78 GND.n77 76
R288 GND.n71 GND.n70 76
R289 GND.n68 GND.n67 76
R290 GND.n65 GND.n64 76
R291 GND.n62 GND.n61 76
R292 GND.n59 GND.n58 76
R293 GND.n56 GND.n55 76
R294 GND.n48 GND.n47 76
R295 GND.n12 GND.n11 76
R296 GND.n20 GND.n19 76
R297 GND.n23 GND.n22 76
R298 GND.n26 GND.n25 76
R299 GND.n33 GND.n32 76
R300 GND.n36 GND.n35 76
R301 GND.n39 GND.n38 76
R302 GND.n53 GND.n52 63.835
R303 GND.n17 GND.n16 63.835
R304 GND.n8 GND.n7 34.942
R305 GND.n52 GND.n51 28.421
R306 GND.n16 GND.n15 28.421
R307 GND.n52 GND.n50 25.263
R308 GND.n16 GND.n14 25.263
R309 GND.n50 GND.n49 24.383
R310 GND.n14 GND.n13 24.383
R311 GND.n5 GND.n4 14.167
R312 GND.n4 GND.n2 14.167
R313 GND.n32 GND.n30 14.167
R314 GND.n77 GND.n76 14.167
R315 GND.n47 GND.n46 13.653
R316 GND.n55 GND.n54 13.653
R317 GND.n58 GND.n57 13.653
R318 GND.n61 GND.n60 13.653
R319 GND.n64 GND.n63 13.653
R320 GND.n67 GND.n66 13.653
R321 GND.n70 GND.n69 13.653
R322 GND.n77 GND.n72 13.653
R323 GND.n80 GND.n79 13.653
R324 GND.n85 GND.n84 13.653
R325 GND.n88 GND.n87 13.653
R326 GND.n41 GND.n40 13.653
R327 GND.n5 GND.n0 13.653
R328 GND.n4 GND.n3 13.653
R329 GND.n2 GND.n1 13.653
R330 GND.n11 GND.n10 13.653
R331 GND.n19 GND.n18 13.653
R332 GND.n22 GND.n21 13.653
R333 GND.n25 GND.n24 13.653
R334 GND.n32 GND.n31 13.653
R335 GND.n35 GND.n34 13.653
R336 GND.n38 GND.n37 13.653
R337 GND.n30 GND.n29 7.312
R338 GND.n76 GND.n75 7.312
R339 GND.n7 GND.n6 7.084
R340 GND.n7 GND.n5 6.475
R341 GND.n19 GND.n17 3.935
R342 GND.n85 GND.n83 3.935
R343 GND.n55 GND.n53 3.935
R344 GND.n44 GND.n43 0.596
R345 GND.n33 GND.n26 0.29
R346 GND.n78 GND.n71 0.29
R347 GND.n45 GND 0.207
R348 GND.n12 GND.n9 0.181
R349 GND.n62 GND.n59 0.181
R350 GND.n9 GND.n8 0.145
R351 GND.n20 GND.n12 0.145
R352 GND.n23 GND.n20 0.145
R353 GND.n26 GND.n23 0.145
R354 GND.n36 GND.n33 0.145
R355 GND.n39 GND.n36 0.145
R356 GND.n42 GND.n39 0.145
R357 GND.n89 GND.n86 0.145
R358 GND.n86 GND.n81 0.145
R359 GND.n81 GND.n78 0.145
R360 GND.n71 GND.n68 0.145
R361 GND.n68 GND.n65 0.145
R362 GND.n65 GND.n62 0.145
R363 GND.n59 GND.n56 0.145
R364 GND.n56 GND.n48 0.145
R365 GND.n48 GND.n45 0.145
R366 GND GND.n42 0.09
R367 GND GND.n89 0.09
R368 a_112_101.n1 a_112_101.n0 32.249
R369 a_112_101.t0 a_112_101.n5 7.911
R370 a_112_101.n4 a_112_101.n2 4.032
R371 a_112_101.n4 a_112_101.n3 3.644
R372 a_112_101.t0 a_112_101.n1 2.534
R373 a_112_101.t0 a_112_101.n4 1.099
R374 a_1444_101.t0 a_1444_101.n1 34.62
R375 a_1444_101.t0 a_1444_101.n0 8.137
R376 a_1444_101.t0 a_1444_101.n2 4.69
C10 VDD GND 8.11fF
C11 a_1444_101.n0 GND 0.06fF
C12 a_1444_101.n1 GND 0.13fF
C13 a_1444_101.n2 GND 0.04fF
C14 a_112_101.n0 GND 0.10fF
C15 a_112_101.n1 GND 0.09fF
C16 a_112_101.n2 GND 0.08fF
C17 a_112_101.n3 GND 0.02fF
C18 a_112_101.n4 GND 0.01fF
C19 a_112_101.n5 GND 0.06fF
C20 a_778_101.n0 GND 0.03fF
C21 a_778_101.n1 GND 0.13fF
C22 a_778_101.n2 GND 0.13fF
C23 a_778_101.n3 GND 0.15fF
C24 VDD.n0 GND 0.15fF
C25 VDD.n1 GND 0.02fF
C26 VDD.n2 GND 0.02fF
C27 VDD.n3 GND 0.04fF
C28 VDD.n4 GND 0.01fF
C29 VDD.n5 GND 0.02fF
C30 VDD.n6 GND 0.02fF
C31 VDD.n9 GND 0.02fF
C32 VDD.n10 GND 0.02fF
C33 VDD.n11 GND 0.02fF
C34 VDD.n14 GND 0.45fF
C35 VDD.n16 GND 0.03fF
C36 VDD.n17 GND 0.02fF
C37 VDD.n18 GND 0.02fF
C38 VDD.n19 GND 0.02fF
C39 VDD.n20 GND 0.04fF
C40 VDD.n21 GND 0.27fF
C41 VDD.n22 GND 0.02fF
C42 VDD.n23 GND 0.03fF
C43 VDD.n24 GND 0.27fF
C44 VDD.n25 GND 0.01fF
C45 VDD.n26 GND 0.31fF
C46 VDD.n27 GND 0.01fF
C47 VDD.n28 GND 0.03fF
C48 VDD.n29 GND 0.02fF
C49 VDD.n30 GND 0.27fF
C50 VDD.n31 GND 0.01fF
C51 VDD.n32 GND 0.02fF
C52 VDD.n33 GND 0.00fF
C53 VDD.n34 GND 0.09fF
C54 VDD.n35 GND 0.03fF
C55 VDD.n36 GND 0.31fF
C56 VDD.n37 GND 0.01fF
C57 VDD.n38 GND 0.03fF
C58 VDD.n39 GND 0.03fF
C59 VDD.n40 GND 0.27fF
C60 VDD.n41 GND 0.01fF
C61 VDD.n42 GND 0.02fF
C62 VDD.n43 GND 0.02fF
C63 VDD.n44 GND 0.27fF
C64 VDD.n45 GND 0.01fF
C65 VDD.n46 GND 0.02fF
C66 VDD.n47 GND 0.02fF
C67 VDD.n48 GND 0.27fF
C68 VDD.n49 GND 0.01fF
C69 VDD.n50 GND 0.02fF
C70 VDD.n51 GND 0.03fF
C71 VDD.n52 GND 0.02fF
C72 VDD.n53 GND 0.02fF
C73 VDD.n54 GND 0.02fF
C74 VDD.n55 GND 0.22fF
C75 VDD.n56 GND 0.04fF
C76 VDD.n57 GND 0.04fF
C77 VDD.n58 GND 0.02fF
C78 VDD.n60 GND 0.02fF
C79 VDD.n61 GND 0.02fF
C80 VDD.n62 GND 0.02fF
C81 VDD.n63 GND 0.02fF
C82 VDD.n65 GND 0.02fF
C83 VDD.n66 GND 0.02fF
C84 VDD.n67 GND 0.02fF
C85 VDD.n69 GND 0.27fF
C86 VDD.n71 GND 0.02fF
C87 VDD.n72 GND 0.02fF
C88 VDD.n73 GND 0.03fF
C89 VDD.n74 GND 0.02fF
C90 VDD.n75 GND 0.27fF
C91 VDD.n76 GND 0.01fF
C92 VDD.n77 GND 0.02fF
C93 VDD.n78 GND 0.03fF
C94 VDD.n79 GND 0.27fF
C95 VDD.n80 GND 0.01fF
C96 VDD.n81 GND 0.02fF
C97 VDD.n82 GND 0.02fF
C98 VDD.n83 GND 0.27fF
C99 VDD.n84 GND 0.01fF
C100 VDD.n85 GND 0.02fF
C101 VDD.n86 GND 0.02fF
C102 VDD.n87 GND 0.31fF
C103 VDD.n88 GND 0.01fF
C104 VDD.n89 GND 0.03fF
C105 VDD.n90 GND 0.02fF
C106 VDD.n91 GND 0.02fF
C107 VDD.n92 GND 0.02fF
C108 VDD.n93 GND 0.02fF
C109 VDD.n94 GND 0.15fF
C110 VDD.n95 GND 0.03fF
C111 VDD.n96 GND 0.02fF
C112 VDD.n97 GND 0.02fF
C113 VDD.n98 GND 0.02fF
C114 VDD.n99 GND 0.02fF
C115 VDD.n100 GND 0.02fF
C116 VDD.n102 GND 0.02fF
C117 VDD.n103 GND 0.02fF
C118 VDD.n104 GND 0.02fF
C119 VDD.n106 GND 0.45fF
C120 VDD.n108 GND 0.03fF
C121 VDD.n109 GND 0.04fF
C122 VDD.n110 GND 0.27fF
C123 VDD.n111 GND 0.02fF
C124 VDD.n112 GND 0.03fF
C125 VDD.n113 GND 0.03fF
C126 VDD.n114 GND 0.06fF
C127 VDD.n115 GND 0.25fF
C128 VDD.n116 GND 0.01fF
C129 VDD.n117 GND 0.01fF
C130 VDD.n118 GND 0.02fF
C131 VDD.n119 GND 0.14fF
C132 VDD.n120 GND 0.16fF
C133 VDD.n121 GND 0.01fF
C134 VDD.n122 GND 0.02fF
C135 VDD.n123 GND 0.02fF
C136 VDD.n124 GND 0.17fF
C137 VDD.n125 GND 0.14fF
C138 VDD.n126 GND 0.01fF
C139 VDD.n127 GND 0.02fF
C140 VDD.n128 GND 0.03fF
C141 VDD.n129 GND 0.11fF
C142 VDD.n130 GND 0.03fF
C143 VDD.n131 GND 0.30fF
C144 VDD.n132 GND 0.01fF
C145 VDD.n133 GND 0.02fF
C146 VDD.n134 GND 0.03fF
C147 VDD.n135 GND 0.14fF
C148 VDD.n136 GND 0.17fF
C149 VDD.n137 GND 0.01fF
C150 VDD.n138 GND 0.02fF
C151 VDD.n139 GND 0.02fF
C152 VDD.n140 GND 0.06fF
C153 VDD.n141 GND 0.24fF
C154 VDD.n142 GND 0.01fF
C155 VDD.n143 GND 0.01fF
C156 VDD.n144 GND 0.02fF
C157 VDD.n145 GND 0.27fF
C158 VDD.n146 GND 0.01fF
C159 VDD.n147 GND 0.02fF
C160 VDD.n148 GND 0.03fF
C161 VDD.n149 GND 0.02fF
C162 VDD.n150 GND 0.02fF
C163 VDD.n151 GND 0.02fF
C164 VDD.n152 GND 0.02fF
C165 VDD.n153 GND 0.02fF
C166 VDD.n154 GND 0.02fF
C167 VDD.n156 GND 0.02fF
C168 VDD.n157 GND 0.02fF
C169 VDD.n158 GND 0.02fF
C170 VDD.n159 GND 0.02fF
C171 VDD.n161 GND 0.04fF
C172 VDD.n162 GND 0.02fF
C173 VDD.n163 GND 0.22fF
C174 VDD.n164 GND 0.04fF
C175 VDD.n166 GND 0.27fF
C176 VDD.n168 GND 0.02fF
C177 VDD.n169 GND 0.02fF
C178 VDD.n170 GND 0.03fF
C179 VDD.n171 GND 0.02fF
C180 VDD.n172 GND 0.27fF
C181 VDD.n173 GND 0.01fF
C182 VDD.n174 GND 0.02fF
C183 VDD.n175 GND 0.03fF
C184 VDD.n176 GND 0.27fF
C185 VDD.n177 GND 0.01fF
C186 VDD.n178 GND 0.02fF
C187 VDD.n179 GND 0.02fF
C188 VDD.n180 GND 0.27fF
C189 VDD.n181 GND 0.01fF
C190 VDD.n182 GND 0.02fF
C191 VDD.n183 GND 0.02fF
C192 VDD.n184 GND 0.31fF
C193 VDD.n185 GND 0.01fF
C194 VDD.n186 GND 0.03fF
C195 VDD.n187 GND 0.02fF
C196 YN.n0 GND 0.41fF
C197 YN.n1 GND 0.49fF
C198 YN.n2 GND 0.25fF
C199 YN.n3 GND 0.04fF
C200 YN.n4 GND 0.05fF
C201 YN.n5 GND 0.10fF
C202 YN.n6 GND 0.04fF
C203 YN.n7 GND 0.05fF
C204 YN.n8 GND 0.03fF
C205 YN.n9 GND 0.10fF
C206 YN.n10 GND 1.05fF
C207 YN.n11 GND 0.06fF
C208 YN.n12 GND 0.03fF
C209 YN.n13 GND 0.08fF
C210 YN.n14 GND 0.27fF
C211 YN.n15 GND 0.36fF
C212 YN.n16 GND 0.01fF
C213 a_217_1051.n0 GND 0.36fF
C214 a_217_1051.n1 GND 0.40fF
C215 a_217_1051.n2 GND 0.28fF
C216 a_217_1051.n3 GND 0.62fF
C217 a_217_1051.n4 GND 0.23fF
C218 a_217_1051.n5 GND 0.32fF
C219 a_881_1051.n0 GND 0.27fF
C220 a_881_1051.n1 GND 0.35fF
C221 a_881_1051.n2 GND 0.24fF
C222 a_881_1051.n3 GND 0.55fF
C223 a_881_1051.n4 GND 0.20fF
C224 a_881_1051.n5 GND 0.28fF
.ends
