* SPICE3 file created from AOI3X1.ext - technology: sky130A

.subckt AOI3X1 YN A B C VDD GND
X0 GND A aoi3x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X1 aoi3x1_pcell_0/m1_537_501# B aoi3x1_pcell_0/nand2x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X2 VDD A aoi3x1_pcell_0/m1_537_501# VDD pshort w=2 l=0.15
X3 VDD B aoi3x1_pcell_0/m1_537_501# VDD pshort w=2 l=0.15
X4 VDD aoi3x1_pcell_0/m1_537_501# aoi3x1_pcell_0/nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X5 YN C aoi3x1_pcell_0/nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X6 YN aoi3x1_pcell_0/m1_537_501# GND GND nshort w=3 l=0.15
X7 YN C GND GND nshort w=3 l=0.15
C0 VDD GND 2.54fF
.ends
