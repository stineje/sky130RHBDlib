magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 133 157 919 203
rect 36 21 919 157
rect 36 17 58 21
rect 24 -17 58 17
<< scnmos >>
rect 114 47 144 131
rect 209 47 239 177
rect 397 47 427 131
rect 492 47 522 177
rect 716 47 746 131
rect 811 47 841 177
<< scpmoshvt >>
rect 114 413 144 497
rect 209 297 239 497
rect 397 413 427 497
rect 492 297 522 497
rect 716 413 746 497
rect 811 297 841 497
<< ndiff >>
rect 159 131 209 177
rect 62 106 114 131
rect 62 72 70 106
rect 104 72 114 106
rect 62 47 114 72
rect 144 93 209 131
rect 144 59 159 93
rect 193 59 209 93
rect 144 47 209 59
rect 239 105 291 177
rect 442 131 492 177
rect 239 71 249 105
rect 283 71 291 105
rect 239 47 291 71
rect 345 105 397 131
rect 345 71 353 105
rect 387 71 397 105
rect 345 47 397 71
rect 427 93 492 131
rect 427 59 442 93
rect 476 59 492 93
rect 427 47 492 59
rect 522 105 574 177
rect 761 131 811 177
rect 522 71 532 105
rect 566 71 574 105
rect 522 47 574 71
rect 664 105 716 131
rect 664 71 672 105
rect 706 71 716 105
rect 664 47 716 71
rect 746 93 811 131
rect 746 59 761 93
rect 795 59 811 93
rect 746 47 811 59
rect 841 105 893 177
rect 841 71 851 105
rect 885 71 893 105
rect 841 47 893 71
<< pdiff >>
rect 62 472 114 497
rect 62 438 70 472
rect 104 438 114 472
rect 62 413 114 438
rect 144 489 209 497
rect 144 455 160 489
rect 194 455 209 489
rect 144 413 209 455
rect 159 297 209 413
rect 239 477 291 497
rect 239 443 249 477
rect 283 443 291 477
rect 239 409 291 443
rect 345 472 397 497
rect 345 438 353 472
rect 387 438 397 472
rect 345 413 397 438
rect 427 489 492 497
rect 427 455 443 489
rect 477 455 492 489
rect 427 413 492 455
rect 239 375 249 409
rect 283 375 291 409
rect 239 297 291 375
rect 442 297 492 413
rect 522 477 574 497
rect 522 443 532 477
rect 566 443 574 477
rect 522 409 574 443
rect 664 472 716 497
rect 664 438 672 472
rect 706 438 716 472
rect 664 413 716 438
rect 746 489 811 497
rect 746 455 762 489
rect 796 455 811 489
rect 746 413 811 455
rect 522 375 532 409
rect 566 375 574 409
rect 522 297 574 375
rect 761 297 811 413
rect 841 477 893 497
rect 841 443 851 477
rect 885 443 893 477
rect 841 409 893 443
rect 841 375 851 409
rect 885 375 893 409
rect 841 297 893 375
<< ndiffc >>
rect 70 72 104 106
rect 159 59 193 93
rect 249 71 283 105
rect 353 71 387 105
rect 442 59 476 93
rect 532 71 566 105
rect 672 71 706 105
rect 761 59 795 93
rect 851 71 885 105
<< pdiffc >>
rect 70 438 104 472
rect 160 455 194 489
rect 249 443 283 477
rect 353 438 387 472
rect 443 455 477 489
rect 249 375 283 409
rect 532 443 566 477
rect 672 438 706 472
rect 762 455 796 489
rect 532 375 566 409
rect 851 443 885 477
rect 851 375 885 409
<< poly >>
rect 114 497 144 523
rect 209 497 239 523
rect 397 497 427 523
rect 492 497 522 523
rect 716 497 746 523
rect 811 497 841 523
rect 114 265 144 413
rect 209 265 239 297
rect 397 265 427 413
rect 492 265 522 297
rect 716 265 746 413
rect 811 265 841 297
rect 57 249 144 265
rect 57 215 67 249
rect 101 215 144 249
rect 57 199 144 215
rect 186 249 240 265
rect 186 215 196 249
rect 230 215 240 249
rect 186 199 240 215
rect 340 249 427 265
rect 340 215 350 249
rect 384 215 427 249
rect 340 199 427 215
rect 469 249 523 265
rect 469 215 479 249
rect 513 215 523 249
rect 469 199 523 215
rect 659 249 746 265
rect 659 215 669 249
rect 703 215 746 249
rect 659 199 746 215
rect 788 249 842 265
rect 788 215 798 249
rect 832 215 842 249
rect 788 199 842 215
rect 114 131 144 199
rect 209 177 239 199
rect 397 131 427 199
rect 492 177 522 199
rect 716 131 746 199
rect 811 177 841 199
rect 114 21 144 47
rect 209 21 239 47
rect 397 21 427 47
rect 492 21 522 47
rect 716 21 746 47
rect 811 21 841 47
<< polycont >>
rect 67 215 101 249
rect 196 215 230 249
rect 350 215 384 249
rect 479 215 513 249
rect 669 215 703 249
rect 798 215 832 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 472 104 493
rect 17 438 70 472
rect 138 489 215 527
rect 138 455 160 489
rect 194 455 215 489
rect 138 442 215 455
rect 249 477 303 493
rect 283 443 303 477
rect 17 408 104 438
rect 249 409 303 443
rect 17 374 215 408
rect 17 249 114 340
rect 17 215 67 249
rect 101 215 114 249
rect 17 199 114 215
rect 148 265 215 374
rect 283 375 303 409
rect 249 335 303 375
rect 337 472 387 493
rect 337 438 353 472
rect 421 489 498 527
rect 421 455 443 489
rect 477 455 498 489
rect 421 442 498 455
rect 532 477 621 493
rect 566 443 621 477
rect 337 408 387 438
rect 532 409 621 443
rect 337 369 498 408
rect 249 299 394 335
rect 148 249 230 265
rect 148 215 196 249
rect 148 199 230 215
rect 264 249 394 299
rect 264 215 350 249
rect 384 215 394 249
rect 264 199 394 215
rect 428 265 498 369
rect 566 375 621 409
rect 532 335 621 375
rect 655 472 706 493
rect 655 438 672 472
rect 740 489 817 527
rect 740 455 762 489
rect 796 455 817 489
rect 740 442 817 455
rect 851 477 903 493
rect 885 443 903 477
rect 655 408 706 438
rect 851 409 903 443
rect 655 369 817 408
rect 532 299 713 335
rect 428 249 513 265
rect 428 215 479 249
rect 428 199 513 215
rect 547 249 713 299
rect 547 215 669 249
rect 703 215 713 249
rect 547 199 713 215
rect 747 265 817 369
rect 885 375 903 409
rect 851 299 903 375
rect 747 249 832 265
rect 747 215 798 249
rect 747 199 832 215
rect 148 165 215 199
rect 264 165 303 199
rect 428 165 498 199
rect 547 165 621 199
rect 747 165 817 199
rect 866 165 903 299
rect 17 131 215 165
rect 17 106 104 131
rect 17 72 70 106
rect 249 105 303 165
rect 17 51 104 72
rect 138 93 215 97
rect 138 59 159 93
rect 193 59 215 93
rect 138 17 215 59
rect 283 71 303 105
rect 249 51 303 71
rect 337 131 498 165
rect 337 105 387 131
rect 337 71 353 105
rect 532 105 621 165
rect 337 51 387 71
rect 421 93 498 97
rect 421 59 442 93
rect 476 59 498 93
rect 421 17 498 59
rect 566 71 621 105
rect 532 51 621 71
rect 655 131 817 165
rect 655 105 706 131
rect 655 71 672 105
rect 851 105 903 165
rect 655 51 706 71
rect 740 93 817 97
rect 740 59 761 93
rect 795 59 817 93
rect 740 17 817 59
rect 885 71 903 105
rect 851 51 903 71
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel metal1 s 24 527 58 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 24 -17 58 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel nwell s 24 527 58 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 24 -17 58 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel locali s 24 221 58 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 580 289 614 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 24 289 58 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 580 357 614 391 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 580 425 614 459 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 580 221 614 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 580 153 614 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 580 85 614 119 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 672 221 706 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 672 289 706 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
rlabel comment s 0 0 0 0 4 dlymetal6s4s_1
rlabel metal1 s 0 -48 920 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 920 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string LEFsymmetry X Y R90
string GDS_END 2909810
string GDS_START 2902034
string path 0.000 13.600 23.000 13.600 
<< end >>
