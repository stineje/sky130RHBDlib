* SPICE3 file created from INVX1.ext - technology: sky130A

.subckt INVX1 Y A VDD VSS
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0058 pd=4.58 as=0.0011 ps=9.1 w=2 l=0.15 M=2
X1 Y A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.001791 pd=1.57 as=0.0011408 ps=8.1 w=3 l=0.15
.ends
