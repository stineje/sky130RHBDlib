* SPICE3 file created from TIEHI.ext - technology: sky130A

.subckt TIEHI Y VPB VNB
M1000 a_121_383# a_121_383# VNB VNB nshort w=3u l=0.15u
+  ad=0p pd=0u as=1.1408p ps=8.1u

R0 VPB.n44 VPB.n43 13.653
R1 VPB.n43 VPB.n42 13.653
R2 VPB.n51 VPB.n50 13.653
R3 VPB.n50 VPB.n49 13.653
R4 VPB.n48 VPB.n47 13.653
R5 VPB.n47 VPB.n46 13.653
R6 VPB.n55 VPB.n0 13.653
R7 VPB VPB.n0 13.653
R8 VPB.n59 VPB.n58 13.276
R9 VPB.n58 VPB.n56 13.276
R10 VPB.n51 VPB.n44 13.276
R11 VPB.n51 VPB.n48 13.276
R12 VPB.n36 VPB.n18 13.276
R13 VPB.n18 VPB.n16 13.276
R14 VPB.n23 VPB.n21 12.796
R15 VPB.n23 VPB.n22 12.564
R16 VPB.n31 VPB.n30 12.198
R17 VPB.n27 VPB.n26 12.198
R18 VPB.n31 VPB.n28 12.198
R19 VPB.n40 VPB.n39 10.764
R20 VPB.n55 VPB.n14 10.764
R21 VPB.n36 VPB.n35 7.5
R22 VPB.n21 VPB.n20 7.5
R23 VPB.n26 VPB.n25 7.5
R24 VPB.n30 VPB.n29 7.5
R25 VPB.n18 VPB.n17 7.5
R26 VPB.n33 VPB.n19 7.5
R27 VPB.n58 VPB.n57 7.5
R28 VPB.n12 VPB.n11 7.5
R29 VPB.n6 VPB.n5 7.5
R30 VPB.n8 VPB.n7 7.5
R31 VPB.n2 VPB.n1 7.5
R32 VPB.n60 VPB.n59 7.5
R33 VPB.n13 VPB.n10 6.729
R34 VPB.n9 VPB.n6 6.729
R35 VPB.n4 VPB.n2 6.729
R36 VPB.n4 VPB.n3 6.728
R37 VPB.n9 VPB.n8 6.728
R38 VPB.n13 VPB.n12 6.728
R39 VPB.n61 VPB.n60 6.728
R40 VPB.n35 VPB.n34 6.398
R41 VPB.n44 VPB.n40 2.511
R42 VPB.n48 VPB.n14 2.511
R43 VPB.n33 VPB.n24 1.402
R44 VPB.n33 VPB.n27 1.402
R45 VPB.n33 VPB.n31 1.402
R46 VPB.n33 VPB.n32 1.402
R47 VPB.n34 VPB.n33 0.735
R48 VPB.n33 VPB.n23 0.735
R49 VPB.n62 VPB.n13 0.387
R50 VPB.n62 VPB.n9 0.387
R51 VPB.n62 VPB.n4 0.387
R52 VPB.n62 VPB.n61 0.387
R53 VPB.n54 VPB 0.198
R54 VPB.n52 VPB.n15 0.136
R55 VPB.n53 VPB.n52 0.136
R56 VPB.n54 VPB.n53 0.136
R57 a_193_1004.t0 a_193_1004.t1 28.564
R58 VNB VNB.n56 1525
R59 VNB.n56 VNB 1525
R60 VNB.n31 VNB.n7 76
R61 VNB.n36 VNB.n35 76
R62 VNB.n54 VNB.n38 76
R63 VNB.n11 VNB.n10 35.01
R64 VNB.t0 VNB.n2 32.601
R65 VNB.n28 VNB.n26 20.452
R66 VNB.n54 VNB.n53 20.452
R67 VNB.n35 VNB.n8 19.735
R68 VNB.n29 VNB.n11 19.735
R69 VNB.n6 VNB.n5 19.735
R70 VNB.n11 VNB.n9 19.017
R71 VNB.n15 VNB.n12 18.356
R72 VNB.n42 VNB.n39 18.356
R73 VNB.n4 VNB.t0 17.353
R74 VNB.n18 VNB.n15 13.919
R75 VNB.n45 VNB.n42 13.919
R76 VNB.n34 VNB.n33 13.653
R77 VNB.n35 VNB.n32 13.653
R78 VNB.n31 VNB.n30 13.653
R79 VNB.n28 VNB.n27 13.653
R80 VNB.n55 VNB.n54 13.653
R81 VNB.n56 VNB.n55 13.653
R82 VNB.n21 VNB.n18 13.276
R83 VNB.n24 VNB.n21 13.276
R84 VNB.n26 VNB.n24 13.276
R85 VNB.n48 VNB.n45 13.276
R86 VNB.n51 VNB.n48 13.276
R87 VNB.n53 VNB.n51 13.276
R88 VNB.n35 VNB.n31 13.276
R89 VNB.n35 VNB.n34 13.276
R90 VNB.n5 VNB.n4 12.837
R91 VNB.n54 VNB.n6 9.329
R92 VNB.n29 VNB.n28 8.97
R93 VNB.n4 VNB.n3 7.566
R94 VNB.n26 VNB.n25 7.5
R95 VNB.n14 VNB.n13 7.5
R96 VNB.n18 VNB.n17 7.5
R97 VNB.n17 VNB.n16 7.5
R98 VNB.n21 VNB.n20 7.5
R99 VNB.n20 VNB.n19 7.5
R100 VNB.n24 VNB.n23 7.5
R101 VNB.n41 VNB.n40 7.5
R102 VNB.n53 VNB.n52 7.5
R103 VNB.n51 VNB.n50 7.5
R104 VNB.n48 VNB.n47 7.5
R105 VNB.n47 VNB.n46 7.5
R106 VNB.n45 VNB.n44 7.5
R107 VNB.n44 VNB.n43 7.5
R108 VNB.n15 VNB.n14 6.627
R109 VNB.n42 VNB.n41 6.627
R110 VNB.n1 VNB.n0 4.551
R111 VNB.n31 VNB.n29 4.305
R112 VNB.n34 VNB.n6 3.947
R113 VNB.t0 VNB.n1 2.238
R114 VNB.n23 VNB.n22 0.454
R115 VNB.n50 VNB.n49 0.454
R116 VNB.n38 VNB 0.198
R117 VNB.n36 VNB.n7 0.136
R118 VNB.n37 VNB.n36 0.136
R119 VNB.n38 VNB.n37 0.136





















































.ends
