// File: nmos_top.spi.NMOS_TOP.pxi
// Created: Tue Oct 15 15:58:44 2024
// 
simulator lang=spectre
cc_1 ( noxref_1 noxref_2 ) capacitor c=0.046371f //x=0.42 //y=0.54 //x2=0 //y2=0
cc_2 ( noxref_1 noxref_3 ) capacitor c=0.016062f //x=0.42 //y=0.54 //x2=0.61 \
 //y2=0.965
cc_3 ( noxref_2 noxref_3 ) capacitor c=0.0904498f //x=0 //y=0 //x2=0.61 \
 //y2=0.965
