magic
tech sky130A
magscale 1 2
timestamp 1645210163
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 2 21 1839 203
rect 30 -17 64 21
<< locali >>
rect 22 215 89 273
rect 191 215 259 265
rect 368 283 637 341
rect 603 181 637 283
rect 1030 215 1421 257
rect 1475 215 1822 257
rect 387 145 1733 181
rect 387 51 453 145
rect 555 51 621 145
rect 723 51 789 145
rect 891 51 957 145
rect 1163 51 1229 145
rect 1331 51 1397 145
rect 1499 51 1565 145
rect 1667 51 1733 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 17 409 73 493
rect 107 443 173 527
rect 303 459 1039 493
rect 303 443 705 459
rect 17 375 705 409
rect 17 307 157 375
rect 191 307 327 341
rect 123 179 157 307
rect 293 249 327 307
rect 293 215 569 249
rect 293 181 327 215
rect 671 257 705 375
rect 739 325 781 425
rect 815 359 865 459
rect 899 325 949 425
rect 983 359 1039 459
rect 1076 459 1473 493
rect 1076 359 1137 459
rect 1171 325 1221 425
rect 1255 359 1305 459
rect 1339 325 1389 425
rect 739 291 1389 325
rect 1423 325 1473 459
rect 1507 359 1557 527
rect 1591 325 1641 493
rect 1675 359 1725 527
rect 1759 325 1822 493
rect 1423 291 1822 325
rect 671 215 981 257
rect 17 145 157 179
rect 191 147 327 181
rect 17 51 89 145
rect 123 17 157 111
rect 191 51 257 147
rect 319 17 353 111
rect 487 17 521 111
rect 655 17 689 111
rect 823 17 857 111
rect 991 17 1129 111
rect 1263 17 1297 111
rect 1431 17 1465 111
rect 1599 17 1633 111
rect 1767 17 1822 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
rlabel locali s 1475 215 1822 257 6 A
port 1 nsew signal input
rlabel locali s 1030 215 1421 257 6 B
port 2 nsew signal input
rlabel locali s 22 215 89 273 6 C_N
port 3 nsew signal input
rlabel locali s 191 215 259 265 6 D_N
port 4 nsew signal input
rlabel metal1 s 0 -48 1840 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 2 21 1839 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1878 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1840 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1667 51 1733 145 6 Y
port 9 nsew signal output
rlabel locali s 1499 51 1565 145 6 Y
port 9 nsew signal output
rlabel locali s 1331 51 1397 145 6 Y
port 9 nsew signal output
rlabel locali s 1163 51 1229 145 6 Y
port 9 nsew signal output
rlabel locali s 891 51 957 145 6 Y
port 9 nsew signal output
rlabel locali s 723 51 789 145 6 Y
port 9 nsew signal output
rlabel locali s 555 51 621 145 6 Y
port 9 nsew signal output
rlabel locali s 387 51 453 145 6 Y
port 9 nsew signal output
rlabel locali s 387 145 1733 181 6 Y
port 9 nsew signal output
rlabel locali s 603 181 637 283 6 Y
port 9 nsew signal output
rlabel locali s 368 283 637 341 6 Y
port 9 nsew signal output
<< properties >>
string LEFsite unithd
string LEFclass CORE
string FIXED_BBOX 0 0 1840 544
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_END 1229000
string GDS_START 1215476
<< end >>
