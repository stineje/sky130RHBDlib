* SPICE3 file created from AOI3X1.ext - technology: sky130A

.subckt AOI3X1 YN A B C VDD VSS
X0 VDD A a_217_1050 VDD sky130_fd_pr__pfet_01v8 ad=0.00226 pd=1.826 as=0 ps=0 w=2 l=0.15 M=2
X1 VDD a_217_1050 a_797_1051 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X2 VDD B a_217_1050 VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.15 M=2
X3 a_797_1051 C YN VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.0058 ps=4.58 w=2 l=0.15 M=2
X4 VSS A a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0.0021157 pd=1.451 as=0 ps=0 w=3 l=0.15
X5 YN a_217_1050 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.003582 pd=3.15 as=0 ps=0 w=3 l=0.15
X6 a_217_1050 B a_112_101 VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
X7 YN C VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=3 l=0.15
C0 VDD a_217_1050 2.17f
C1 VDD VSS 2.67f
.ends
