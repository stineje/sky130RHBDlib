magic
tech sky130A
magscale 1 2
timestamp 1652514973
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 427 871 461 905
rect 3017 871 3051 905
rect 5607 871 5641 905
rect 8197 871 8231 905
rect 10787 871 10821 905
rect 13377 871 13411 905
rect 17817 871 17851 905
rect 17817 797 17851 831
rect 427 723 461 757
rect 5607 723 5641 757
rect 9159 723 9193 757
rect 10787 723 10821 757
rect 14339 723 14373 757
rect 17817 723 17851 757
rect 427 649 461 683
rect 3017 649 3051 683
rect 3239 649 3273 683
rect 3979 649 4013 683
rect 5607 649 5641 683
rect 8197 649 8231 683
rect 8419 649 8453 683
rect 9159 649 9193 683
rect 17817 649 17851 683
rect 427 575 461 609
rect 1389 575 1423 609
rect 1611 575 1645 609
rect 3017 575 3051 609
rect 3239 575 3273 609
rect 3979 575 4013 609
rect 17817 575 17851 609
rect 427 501 461 535
rect 1389 501 1423 535
rect 17817 501 17851 535
rect 1611 427 1645 461
rect 17817 427 17851 461
<< metal1 >>
rect -34 1446 18016 1514
rect 2906 871 13416 905
rect 4419 797 4683 831
rect 14779 797 15043 831
rect 9599 723 9863 757
rect 14631 723 15339 757
rect 15421 723 15857 757
rect 9451 649 10159 683
rect 10241 649 15635 683
rect 4271 575 4979 609
rect 5061 575 16671 609
rect 1459 501 6557 535
rect 6639 501 11737 535
rect 3891 427 14375 461
rect -34 -34 18016 34
use li1_M1_contact  li1_M1_contact_4 pcells
timestamp 1648061256
transform -1 0 1406 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 4366 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 4736 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_8
timestamp 1648061256
transform -1 0 4218 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform 1 0 5032 0 1 592
box -53 -33 29 33
use dffrnx1_pcell  dffrnx1_pcell_1 pcells
timestamp 1652425808
transform 1 0 5180 0 1 0
box -87 -34 5267 1550
use dffrnx1_pcell  dffrnx1_pcell_0
timestamp 1652425808
transform 1 0 0 0 1 0
box -87 -34 5267 1550
use li1_M1_contact  li1_M1_contact_16
timestamp 1648061256
transform -1 0 6586 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform 1 0 9916 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform -1 0 9546 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform -1 0 9398 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 10212 0 1 666
box -53 -33 29 33
use dffrnx1_pcell  dffrnx1_pcell_2
timestamp 1652425808
transform 1 0 10360 0 1 0
box -87 -34 5267 1550
use voter3x1_pcell  voter3x1_pcell_0 pcells
timestamp 1652393968
transform 1 0 15540 0 1 0
box -87 -34 2529 1550
use li1_M1_contact  li1_M1_contact_17
timestamp 1648061256
transform -1 0 11766 0 -1 518
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_15
timestamp 1648061256
transform 1 0 15688 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_14
timestamp 1648061256
transform 1 0 15910 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_12
timestamp 1648061256
transform 1 0 15392 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_9
timestamp 1648061256
transform 1 0 15096 0 1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_10
timestamp 1648061256
transform -1 0 14726 0 -1 814
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_11
timestamp 1648061256
transform -1 0 14578 0 -1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 16724 0 1 592
box -53 -33 29 33
<< labels >>
rlabel locali 17817 871 17851 905 1 Q
port 1 nsew signal output
rlabel locali 17817 797 17851 831 1 Q
port 1 nsew signal output
rlabel locali 17817 723 17851 757 1 Q
port 1 nsew signal output
rlabel locali 17817 649 17851 683 1 Q
port 1 nsew signal output
rlabel locali 17817 575 17851 609 1 Q
port 1 nsew signal output
rlabel locali 17817 501 17851 535 1 Q
port 1 nsew signal output
rlabel locali 17817 427 17851 461 1 Q
port 1 nsew signal output
rlabel locali 1389 501 1423 535 1 D
port 2 nsew signal input
rlabel locali 1389 575 1423 609 1 D
port 2 nsew signal input
rlabel locali 427 871 461 905 1 CLK
port 3 nsew signal input
rlabel locali 427 723 461 757 1 CLK
port 3 nsew signal input
rlabel locali 427 649 461 683 1 CLK
port 3 nsew signal input
rlabel locali 427 575 461 609 1 CLK
port 3 nsew signal input
rlabel locali 427 501 461 535 1 CLK
port 3 nsew signal input
rlabel locali 3017 575 3051 609 1 CLK
port 3 nsew signal input
rlabel locali 3017 649 3051 683 1 CLK
port 3 nsew signal input
rlabel locali 5607 649 5641 683 1 CLK
port 3 nsew signal input
rlabel locali 5607 723 5641 757 1 CLK
port 3 nsew signal input
rlabel locali 8197 649 8231 683 1 CLK
port 3 nsew signal input
rlabel locali 10787 723 10821 757 1 CLK
port 3 nsew signal input
rlabel locali 3017 871 3051 905 1 CLK
port 3 nsew signal input
rlabel locali 5607 871 5641 905 1 CLK
port 3 nsew signal input
rlabel locali 8197 871 8231 905 1 CLK
port 3 nsew signal input
rlabel locali 10787 871 10821 905 1 CLK
port 3 nsew signal input
rlabel locali 13377 871 13411 905 1 CLK
port 3 nsew signal input
rlabel locali 1611 575 1645 609 1 RN
port 4 nsew signal input
rlabel locali 1611 427 1645 461 1 RN
port 4 nsew signal input
rlabel locali 3239 575 3273 609 1 RN
port 4 nsew signal input
rlabel locali 3239 649 3273 683 1 RN
port 4 nsew signal input
rlabel locali 3979 649 4013 683 1 RN
port 4 nsew signal input
rlabel locali 3979 575 4013 609 1 RN
port 4 nsew signal input
rlabel locali 8419 649 8453 683 1 RN
port 4 nsew signal input
rlabel locali 9159 649 9193 683 1 RN
port 4 nsew signal input
rlabel locali 9159 723 9193 757 1 RN
port 4 nsew signal input
rlabel locali 14339 723 14373 757 1 RN
port 4 nsew signal input
rlabel metal1 -34 -34 18016 34 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 -34 1446 18016 1514 1 VPWR
port 5 nsew power bidirectional abutment
rlabel nwell 57 1463 91 1497 1 VPB
port 7 nsew power bidirectional
rlabel pwell 57 -17 91 17 1 VNB
port 8 nsew ground bidirectional
<< properties >>
string LEFclass CORE
string LEFsite unithd
string FIXED_BBOX 0 0 17982 1480
string LEFsymmetry X Y R90
<< end >>
