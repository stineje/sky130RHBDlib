// File: NOR3X1.spi.pex
// Created: Tue Oct 15 15:50:29 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_NOR3X1\%GND ( 1 11 23 27 35 39 47 51 62 65 92 )
c51 ( 92 0 ) capacitor c=0.0964353f //x=0.56 //y=0.365
c52 ( 65 0 ) capacitor c=0.203672f //x=0.695 //y=0
c53 ( 62 0 ) capacitor c=0.250916f //x=4.07 //y=0
c54 ( 60 0 ) capacitor c=0.095941f //x=3.69 //y=0
c55 ( 54 0 ) capacitor c=0.00803396f //x=3.605 //y=0.445
c56 ( 51 0 ) capacitor c=0.00510317f //x=3.52 //y=0.53
c57 ( 50 0 ) capacitor c=0.00468234f //x=3.12 //y=0.445
c58 ( 47 0 ) capacitor c=0.00514697f //x=3.035 //y=0.53
c59 ( 42 0 ) capacitor c=0.00468234f //x=2.635 //y=0.445
c60 ( 39 0 ) capacitor c=0.00556167f //x=2.55 //y=0.53
c61 ( 38 0 ) capacitor c=0.00468234f //x=2.15 //y=0.445
c62 ( 35 0 ) capacitor c=0.00556167f //x=2.065 //y=0.53
c63 ( 30 0 ) capacitor c=0.00468234f //x=1.665 //y=0.445
c64 ( 27 0 ) capacitor c=0.00556167f //x=1.58 //y=0.53
c65 ( 26 0 ) capacitor c=0.00468234f //x=1.18 //y=0.445
c66 ( 23 0 ) capacitor c=0.00709092f //x=1.095 //y=0.53
c67 ( 18 0 ) capacitor c=0.00609805f //x=0.695 //y=0.445
c68 ( 11 0 ) capacitor c=0.207649f //x=4.07 //y=0
r69 (  76 77 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.12 //y=0 //x2=3.605 //y2=0
r70 (  75 76 ) resistor r=5.73669 //w=0.357 //l=0.16 //layer=li \
 //thickness=0.1 //x=2.96 //y=0 //x2=3.12 //y2=0
r71 (  73 75 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=2.635 //y=0 //x2=2.96 //y2=0
r72 (  72 73 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.15 //y=0 //x2=2.635 //y2=0
r73 (  71 72 ) resistor r=10.7563 //w=0.357 //l=0.3 //layer=li //thickness=0.1 \
 //x=1.85 //y=0 //x2=2.15 //y2=0
r74 (  69 71 ) resistor r=6.63305 //w=0.357 //l=0.185 //layer=li \
 //thickness=0.1 //x=1.665 //y=0 //x2=1.85 //y2=0
r75 (  68 69 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.18 //y=0 //x2=1.665 //y2=0
r76 (  67 68 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.18 //y2=0
r77 (  65 67 ) resistor r=1.61345 //w=0.357 //l=0.045 //layer=li \
 //thickness=0.1 //x=0.695 //y=0 //x2=0.74 //y2=0
r78 (  60 77 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.69 //y=0 //x2=3.605 //y2=0
r79 (  60 62 ) resistor r=13.6247 //w=0.357 //l=0.38 //layer=li \
 //thickness=0.1 //x=3.69 //y=0 //x2=4.07 //y2=0
r80 (  55 92 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.605 //y=0.615 //x2=3.605 //y2=0.53
r81 (  55 92 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=3.605 //y=0.615 //x2=3.605 //y2=0.88
r82 (  54 92 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.605 //y=0.445 //x2=3.605 //y2=0.53
r83 (  53 77 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.605 //y=0.17 //x2=3.605 //y2=0
r84 (  53 54 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=3.605 //y=0.17 //x2=3.605 //y2=0.445
r85 (  52 92 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.205 //y=0.53 //x2=3.12 //y2=0.53
r86 (  51 92 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.52 //y=0.53 //x2=3.605 //y2=0.53
r87 (  51 52 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.52 //y=0.53 //x2=3.205 //y2=0.53
r88 (  50 92 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.12 //y=0.445 //x2=3.12 //y2=0.53
r89 (  49 76 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.12 //y=0.17 //x2=3.12 //y2=0
r90 (  49 50 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=3.12 //y=0.17 //x2=3.12 //y2=0.445
r91 (  48 92 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.72 //y=0.53 //x2=2.635 //y2=0.53
r92 (  47 92 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.035 //y=0.53 //x2=3.12 //y2=0.53
r93 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.035 //y=0.53 //x2=2.72 //y2=0.53
r94 (  43 92 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.635 //y=0.615 //x2=2.635 //y2=0.53
r95 (  43 92 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r96 (  42 92 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.635 //y=0.445 //x2=2.635 //y2=0.53
r97 (  41 73 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.635 //y=0.17 //x2=2.635 //y2=0
r98 (  41 42 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.17 //x2=2.635 //y2=0.445
r99 (  40 92 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.235 //y=0.53 //x2=2.15 //y2=0.53
r100 (  39 92 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.55 //y=0.53 //x2=2.635 //y2=0.53
r101 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.235 //y2=0.53
r102 (  38 92 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.445 //x2=2.15 //y2=0.53
r103 (  37 72 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.17 //x2=2.15 //y2=0
r104 (  37 38 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.17 //x2=2.15 //y2=0.445
r105 (  36 92 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=1.665 //y2=0.53
r106 (  35 92 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.065 //y=0.53 //x2=2.15 //y2=0.53
r107 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=2.065 //y=0.53 //x2=1.75 //y2=0.53
r108 (  31 92 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.53
r109 (  31 92 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r110 (  30 92 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.445 //x2=1.665 //y2=0.53
r111 (  29 69 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.17 //x2=1.665 //y2=0
r112 (  29 30 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.17 //x2=1.665 //y2=0.445
r113 (  28 92 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0.53 //x2=1.18 //y2=0.53
r114 (  27 92 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.58 //y=0.53 //x2=1.665 //y2=0.53
r115 (  27 28 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.58 //y=0.53 //x2=1.265 //y2=0.53
r116 (  26 92 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.445 //x2=1.18 //y2=0.53
r117 (  25 68 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r118 (  25 26 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.445
r119 (  24 92 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.78 //y=0.53 //x2=0.695 //y2=0.53
r120 (  23 92 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0.53 //x2=1.18 //y2=0.53
r121 (  23 24 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.095 //y=0.53 //x2=0.78 //y2=0.53
r122 (  19 92 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.615 //x2=0.695 //y2=0.53
r123 (  19 92 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.615 //x2=0.695 //y2=1.22
r124 (  18 92 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.445 //x2=0.695 //y2=0.53
r125 (  17 65 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.17 //x2=0.695 //y2=0
r126 (  17 18 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.17 //x2=0.695 //y2=0.445
r127 (  11 62 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r128 (  9 75 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r129 (  9 11 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.07 //y2=0
r130 (  6 71 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r131 (  3 67 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r132 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r133 (  1 9 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=2.405 //y=0 //x2=2.96 //y2=0
r134 (  1 6 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=2.405 //y=0 //x2=1.85 //y2=0
ends PM_NOR3X1\%GND

subckt PM_NOR3X1\%VDD ( 1 11 15 18 32 36 )
c42 ( 36 0 ) capacitor c=0.0267864f //x=1.085 //y=5.025
c43 ( 35 0 ) capacitor c=0.00591168f //x=1.23 //y=7.4
c44 ( 32 0 ) capacitor c=0.351373f //x=4.07 //y=7.4
c45 ( 18 0 ) capacitor c=0.211583f //x=0.74 //y=7.4
c46 ( 15 0 ) capacitor c=0.0465804f //x=1.145 //y=7.4
c47 ( 11 0 ) capacitor c=0.203056f //x=4.07 //y=7.4
r48 (  30 32 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r49 (  28 30 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r50 (  26 35 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.315 //y=7.4 //x2=1.23 //y2=7.4
r51 (  26 28 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=1.315 //y=7.4 //x2=1.85 //y2=7.4
r52 (  19 35 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.23 //y=7.23 //x2=1.23 //y2=7.4
r53 (  19 36 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=1.23 //y=7.23 //x2=1.23 //y2=6.74
r54 (  15 35 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.145 //y=7.4 //x2=1.23 //y2=7.4
r55 (  15 18 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=1.145 //y=7.4 //x2=0.74 //y2=7.4
r56 (  11 32 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=7.4 //x2=4.07 //y2=7.4
r57 (  9 30 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=2.96 \
 //y=7.4 //x2=2.96 //y2=7.4
r58 (  9 11 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r59 (  6 28 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=1.85 \
 //y=7.4 //x2=1.85 //y2=7.4
r60 (  3 18 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=0.74 \
 //y=7.4 //x2=0.74 //y2=7.4
r61 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r62 (  1 9 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=2.405 //y=7.4 //x2=2.96 //y2=7.4
r63 (  1 6 ) resistor r=0.230482 //w=0.301 //l=0.555 //layer=m1 \
 //thickness=0.36 //x=2.405 //y=7.4 //x2=1.85 //y2=7.4
ends PM_NOR3X1\%VDD

subckt PM_NOR3X1\%A ( 1 2 3 4 5 6 7 10 20 22 23 24 25 26 27 28 32 34 37 39 40 \
 45 )
c65 ( 45 0 ) capacitor c=0.04214f //x=0.955 //y=4.705
c66 ( 40 0 ) capacitor c=0.0321911f //x=1.445 //y=1.25
c67 ( 39 0 ) capacitor c=0.0185201f //x=1.445 //y=0.905
c68 ( 37 0 ) capacitor c=0.0344254f //x=1.375 //y=4.795
c69 ( 34 0 ) capacitor c=0.0133656f //x=1.29 //y=1.405
c70 ( 32 0 ) capacitor c=0.0157804f //x=1.29 //y=0.75
c71 ( 28 0 ) capacitor c=0.0828832f //x=0.915 //y=1.915
c72 ( 27 0 ) capacitor c=0.022867f //x=0.915 //y=1.56
c73 ( 26 0 ) capacitor c=0.0234318f //x=0.915 //y=1.25
c74 ( 25 0 ) capacitor c=0.0192004f //x=0.915 //y=0.905
c75 ( 24 0 ) capacitor c=0.110795f //x=1.45 //y=6.025
c76 ( 23 0 ) capacitor c=0.153847f //x=1.01 //y=6.025
c77 ( 20 0 ) capacitor c=0.00995068f //x=0.955 //y=4.705
c78 ( 10 0 ) capacitor c=0.112895f //x=1.11 //y=2.08
r79 (  47 48 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=0.955 //y=4.795 //x2=0.955 //y2=4.87
r80 (  45 47 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=0.955 //y=4.705 //x2=0.955 //y2=4.795
r81 (  40 54 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.25 //x2=1.405 //y2=1.405
r82 (  39 53 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.905 //x2=1.405 //y2=0.75
r83 (  39 40 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.905 //x2=1.445 //y2=1.25
r84 (  38 47 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=1.09 //y=4.795 //x2=0.955 //y2=4.795
r85 (  37 41 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.375 //y=4.795 //x2=1.45 //y2=4.87
r86 (  37 38 ) resistor r=146.138 //w=0.094 //l=0.285 //layer=ply \
 //thickness=0.18 //x=1.375 //y=4.795 //x2=1.09 //y2=4.795
r87 (  35 52 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.405 //x2=0.955 //y2=1.405
r88 (  34 54 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.405 //x2=1.405 //y2=1.405
r89 (  33 51 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.75 //x2=0.955 //y2=0.75
r90 (  32 53 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.75 //x2=1.405 //y2=0.75
r91 (  32 33 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.75 //x2=1.07 //y2=0.75
r92 (  28 50 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r93 (  27 52 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.56 //x2=0.955 //y2=1.405
r94 (  27 28 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.56 //x2=0.915 //y2=1.915
r95 (  26 52 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.25 //x2=0.955 //y2=1.405
r96 (  25 51 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.905 //x2=0.955 //y2=0.75
r97 (  25 26 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.905 //x2=0.915 //y2=1.25
r98 (  24 41 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.025 //x2=1.45 //y2=4.87
r99 (  23 48 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.025 //x2=1.01 //y2=4.87
r100 (  22 34 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.405 //x2=1.29 //y2=1.405
r101 (  22 35 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.405 //x2=1.07 //y2=1.405
r102 (  20 45 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.955 //y=4.705 //x2=0.955 //y2=4.705
r103 (  20 21 ) resistor r=7.81102 //w=0.254 //l=0.155 //layer=li \
 //thickness=0.1 //x=0.955 //y=4.705 //x2=1.11 //y2=4.705
r104 (  10 50 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r105 (  8 21 ) resistor r=3.23951 //w=0.254 //l=0.165 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.54 //x2=1.11 //y2=4.705
r106 (  7 8 ) resistor r=6.84492 //w=0.187 //l=0.1 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.44 //x2=1.11 //y2=4.54
r107 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.44
r108 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=3.7 //x2=1.11 //y2=4.07
r109 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=3.33 //x2=1.11 //y2=3.7
r110 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.96 //x2=1.11 //y2=3.33
r111 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.59 //x2=1.11 //y2=2.96
r112 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.22 //x2=1.11 //y2=2.59
r113 (  1 10 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.22 //x2=1.11 //y2=2.08
ends PM_NOR3X1\%A

subckt PM_NOR3X1\%B ( 1 2 3 4 5 6 7 8 10 21 22 23 24 25 26 31 33 35 41 42 44 \
 45 48 )
c80 ( 48 0 ) capacitor c=0.0366246f //x=1.885 //y=4.705
c81 ( 45 0 ) capacitor c=0.0260062f //x=1.85 //y=1.915
c82 ( 44 0 ) capacitor c=0.0407292f //x=1.85 //y=2.08
c83 ( 42 0 ) capacitor c=0.0170937f //x=2.415 //y=1.255
c84 ( 41 0 ) capacitor c=0.0176605f //x=2.415 //y=0.905
c85 ( 35 0 ) capacitor c=0.0305703f //x=2.26 //y=1.405
c86 ( 33 0 ) capacitor c=0.0157804f //x=2.26 //y=0.75
c87 ( 31 0 ) capacitor c=0.0337811f //x=2.255 //y=4.795
c88 ( 26 0 ) capacitor c=0.0189312f //x=1.885 //y=1.56
c89 ( 25 0 ) capacitor c=0.0169608f //x=1.885 //y=1.255
c90 ( 24 0 ) capacitor c=0.0176782f //x=1.885 //y=0.905
c91 ( 23 0 ) capacitor c=0.13968f //x=2.33 //y=6.025
c92 ( 22 0 ) capacitor c=0.110232f //x=1.89 //y=6.025
c93 ( 10 0 ) capacitor c=0.092194f //x=1.85 //y=2.08
c94 ( 8 0 ) capacitor c=0.00580576f //x=1.85 //y=4.54
r95 (  50 51 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.885 //y=4.795 //x2=1.885 //y2=4.87
r96 (  48 50 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.885 //y=4.705 //x2=1.885 //y2=4.795
r97 (  44 45 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r98 (  42 55 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.255 //x2=2.415 //y2=1.367
r99 (  41 54 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r100 (  41 42 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.255
r101 (  36 53 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r102 (  35 55 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.415 //y2=1.367
r103 (  34 52 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r104 (  33 54 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r105 (  33 34 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r106 (  32 50 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.02 //y=4.795 //x2=1.885 //y2=4.795
r107 (  31 38 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.795 //x2=2.33 //y2=4.87
r108 (  31 32 ) resistor r=120.5 //w=0.094 //l=0.235 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.795 //x2=2.02 //y2=4.795
r109 (  26 53 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r110 (  26 45 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r111 (  25 53 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.255 //x2=1.925 //y2=1.405
r112 (  24 52 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r113 (  24 25 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.255
r114 (  23 38 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.025 //x2=2.33 //y2=4.87
r115 (  22 51 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.025 //x2=1.89 //y2=4.87
r116 (  21 35 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r117 (  21 36 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r118 (  20 48 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.885 //y=4.705 //x2=1.885 //y2=4.705
r119 (  10 44 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r120 (  8 20 ) resistor r=11.332 //w=0.189 //l=0.173292 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.54 //x2=1.867 //y2=4.705
r121 (  7 8 ) resistor r=6.84492 //w=0.187 //l=0.1 //layer=li //thickness=0.1 \
 //x=1.85 //y=4.44 //x2=1.85 //y2=4.54
r122 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=4.07 //x2=1.85 //y2=4.44
r123 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=3.7 //x2=1.85 //y2=4.07
r124 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=3.33 //x2=1.85 //y2=3.7
r125 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=2.96 //x2=1.85 //y2=3.33
r126 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=2.59 //x2=1.85 //y2=2.96
r127 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=2.22 //x2=1.85 //y2=2.59
r128 (  1 10 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=1.85 //y=2.22 //x2=1.85 //y2=2.08
ends PM_NOR3X1\%B

subckt PM_NOR3X1\%noxref_5 ( 7 8 15 16 23 24 25 )
c43 ( 25 0 ) capacitor c=0.0202519f //x=2.405 //y=5.025
c44 ( 24 0 ) capacitor c=0.0185379f //x=1.525 //y=5.025
c45 ( 23 0 ) capacitor c=0.0408953f //x=0.655 //y=5.025
c46 ( 16 0 ) capacitor c=0.00193672f //x=1.755 //y=6.91
c47 ( 15 0 ) capacitor c=0.0126253f //x=2.465 //y=6.91
c48 ( 8 0 ) capacitor c=0.00844339f //x=0.875 //y=5.21
c49 ( 7 0 ) capacitor c=0.0252644f //x=1.585 //y=5.21
r50 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.55 //y=6.825 //x2=2.55 //y2=6.74
r51 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.465 //y=6.91 //x2=2.55 //y2=6.825
r52 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.465 //y=6.91 //x2=1.755 //y2=6.91
r53 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.67 //y=6.825 //x2=1.755 //y2=6.91
r54 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.67 //y=6.825 //x2=1.67 //y2=6.4
r55 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.67 //y=5.295 //x2=1.67 //y2=5.72
r56 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.585 //y=5.21 //x2=1.67 //y2=5.295
r57 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=1.585 //y=5.21 //x2=0.875 //y2=5.21
r58 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=0.79 //y=5.295 //x2=0.875 //y2=5.21
r59 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=0.79 //y=5.295 //x2=0.79 //y2=5.72
ends PM_NOR3X1\%noxref_5

subckt PM_NOR3X1\%C ( 1 2 3 4 5 6 7 9 21 22 23 24 25 26 27 28 30 38 39 40 45 \
 49 )
c67 ( 55 0 ) capacitor c=0.011077f //x=3.37 //y=4.795
c68 ( 49 0 ) capacitor c=0.0431417f //x=2.96 //y=4.705
c69 ( 45 0 ) capacitor c=0.0492905f //x=2.855 //y=2.08
c70 ( 40 0 ) capacitor c=0.0363749f //x=3.735 //y=4.795
c71 ( 39 0 ) capacitor c=0.0237734f //x=3.385 //y=1.255
c72 ( 38 0 ) capacitor c=0.0191782f //x=3.385 //y=0.905
c73 ( 33 0 ) capacitor c=0.0202859f //x=3.295 //y=4.795
c74 ( 30 0 ) capacitor c=0.033152f //x=3.23 //y=1.405
c75 ( 28 0 ) capacitor c=0.0157803f //x=3.23 //y=0.75
c76 ( 27 0 ) capacitor c=0.0280515f //x=2.855 //y=1.915
c77 ( 26 0 ) capacitor c=0.0189445f //x=2.855 //y=1.56
c78 ( 25 0 ) capacitor c=0.0170937f //x=2.855 //y=1.255
c79 ( 24 0 ) capacitor c=0.0185081f //x=2.855 //y=0.905
c80 ( 23 0 ) capacitor c=0.154473f //x=3.81 //y=6.025
c81 ( 22 0 ) capacitor c=0.139411f //x=3.37 //y=6.025
c82 ( 9 0 ) capacitor c=0.0965855f //x=2.96 //y=2.08
r83 (  49 51 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.96 //y=4.705 //x2=2.96 //y2=4.795
r84 (  45 47 ) resistor r=16.5934 //w=0.305 //l=0.105 //layer=ply \
 //thickness=0.18 //x=2.855 //y=2.08 //x2=2.96 //y2=2.08
r85 (  41 55 ) resistor r=20.4101 //w=0.15 //l=0.075 //layer=ply \
 //thickness=0.18 //x=3.445 //y=4.795 //x2=3.37 //y2=4.795
r86 (  40 42 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=3.735 //y=4.795 //x2=3.81 //y2=4.87
r87 (  40 41 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=3.735 //y=4.795 //x2=3.445 //y2=4.795
r88 (  39 57 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=3.385 //y=1.255 //x2=3.385 //y2=1.367
r89 (  38 56 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.385 //y=0.905 //x2=3.345 //y2=0.75
r90 (  38 39 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=3.385 //y=0.905 //x2=3.385 //y2=1.255
r91 (  35 55 ) resistor r=5.30422 //w=0.3 //l=0.075 //layer=ply \
 //thickness=0.18 //x=3.37 //y=4.87 //x2=3.37 //y2=4.795
r92 (  34 51 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=3.095 //y=4.795 //x2=2.96 //y2=4.795
r93 (  33 55 ) resistor r=20.4101 //w=0.15 //l=0.075 //layer=ply \
 //thickness=0.18 //x=3.295 //y=4.795 //x2=3.37 //y2=4.795
r94 (  33 34 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=3.295 //y=4.795 //x2=3.095 //y2=4.795
r95 (  31 54 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.01 //y=1.405 //x2=2.895 //y2=1.405
r96 (  30 57 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=3.23 //y=1.405 //x2=3.385 //y2=1.367
r97 (  29 53 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.01 //y=0.75 //x2=2.895 //y2=0.75
r98 (  28 56 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.23 //y=0.75 //x2=3.345 //y2=0.75
r99 (  28 29 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.23 //y=0.75 //x2=3.01 //y2=0.75
r100 (  27 45 ) resistor r=19.3576 //w=0.305 //l=0.165 //layer=ply \
 //thickness=0.18 //x=2.855 //y=1.915 //x2=2.855 //y2=2.08
r101 (  26 54 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.855 //y=1.56 //x2=2.895 //y2=1.405
r102 (  26 27 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=2.855 //y=1.56 //x2=2.855 //y2=1.915
r103 (  25 54 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=2.855 //y=1.255 //x2=2.895 //y2=1.405
r104 (  24 53 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.855 //y=0.905 //x2=2.895 //y2=0.75
r105 (  24 25 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=2.855 //y=0.905 //x2=2.855 //y2=1.255
r106 (  23 42 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.81 //y=6.025 //x2=3.81 //y2=4.87
r107 (  22 35 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.37 //y=6.025 //x2=3.37 //y2=4.87
r108 (  21 30 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.12 //y=1.405 //x2=3.23 //y2=1.405
r109 (  21 31 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.12 //y=1.405 //x2=3.01 //y2=1.405
r110 (  19 49 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.96 //y=4.705 //x2=2.96 //y2=4.705
r111 (  9 47 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.96 //y=2.08 //x2=2.96 //y2=2.08
r112 (  7 19 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.96 //y=4.44 //x2=2.96 //y2=4.705
r113 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=2.96 //y=4.07 //x2=2.96 //y2=4.44
r114 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=2.96 //y=3.7 //x2=2.96 //y2=4.07
r115 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=2.96 //y=3.33 //x2=2.96 //y2=3.7
r116 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=2.96 //y=2.96 //x2=2.96 //y2=3.33
r117 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=2.96 //y=2.59 //x2=2.96 //y2=2.96
r118 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=2.96 //y=2.22 //x2=2.96 //y2=2.59
r119 (  1 9 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li //thickness=0.1 \
 //x=2.96 //y=2.22 //x2=2.96 //y2=2.08
ends PM_NOR3X1\%C

subckt PM_NOR3X1\%Y ( 1 2 3 4 5 6 7 12 13 18 24 40 43 45 46 47 51 )
c83 ( 51 0 ) capacitor c=0.0159625f //x=3.445 //y=5.025
c84 ( 47 0 ) capacitor c=0.00969064f //x=2.93 //y=0.905
c85 ( 46 0 ) capacitor c=0.00860823f //x=1.96 //y=0.905
c86 ( 45 0 ) capacitor c=0.007684f //x=0.99 //y=0.905
c87 ( 43 0 ) capacitor c=0.00603509f //x=3.7 //y=5.21
c88 ( 40 0 ) capacitor c=0.00544799f //x=3.12 //y=1.655
c89 ( 39 0 ) capacitor c=0.00710337f //x=2.15 //y=1.655
c90 ( 24 0 ) capacitor c=0.0260487f //x=3.615 //y=1.655
c91 ( 18 0 ) capacitor c=0.0281501f //x=3.035 //y=1.655
c92 ( 13 0 ) capacitor c=0.00277859f //x=1.265 //y=1.655
c93 ( 12 0 ) capacitor c=0.0280953f //x=2.065 //y=1.655
c94 ( 1 0 ) capacitor c=0.14166f //x=3.7 //y=2.22
r95 (  41 43 ) resistor r=7.52941 //w=0.187 //l=0.11 //layer=li \
 //thickness=0.1 //x=3.59 //y=5.21 //x2=3.7 //y2=5.21
r96 (  31 43 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.7 //y=5.125 //x2=3.7 //y2=5.21
r97 (  26 41 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.59 //y=5.295 //x2=3.59 //y2=5.21
r98 (  26 51 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=3.59 //y=5.295 //x2=3.59 //y2=6.06
r99 (  25 40 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.205 //y=1.655 //x2=3.12 //y2=1.655
r100 (  24 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.615 //y=1.655 //x2=3.7 //y2=1.74
r101 (  24 25 ) resistor r=28.0642 //w=0.187 //l=0.41 //layer=li \
 //thickness=0.1 //x=3.615 //y=1.655 //x2=3.205 //y2=1.655
r102 (  20 40 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.12 //y=1.57 //x2=3.12 //y2=1.655
r103 (  20 47 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=3.12 //y=1.57 //x2=3.12 //y2=1
r104 (  19 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.235 //y=1.655 //x2=2.15 //y2=1.655
r105 (  18 40 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.035 //y=1.655 //x2=3.12 //y2=1.655
r106 (  18 19 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li \
 //thickness=0.1 //x=3.035 //y=1.655 //x2=2.235 //y2=1.655
r107 (  14 39 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1.655
r108 (  14 46 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r109 (  12 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.065 //y=1.655 //x2=2.15 //y2=1.655
r110 (  12 13 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li \
 //thickness=0.1 //x=2.065 //y=1.655 //x2=1.265 //y2=1.655
r111 (  8 13 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.18 //y=1.57 //x2=1.265 //y2=1.655
r112 (  8 45 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=1.18 //y=1.57 //x2=1.18 //y2=1
r113 (  7 31 ) resistor r=46.8877 //w=0.187 //l=0.685 //layer=li \
 //thickness=0.1 //x=3.7 //y=4.44 //x2=3.7 //y2=5.125
r114 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=3.7 //y=4.07 //x2=3.7 //y2=4.44
r115 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=3.7 //y=3.7 //x2=3.7 //y2=4.07
r116 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=3.7 //y=3.33 //x2=3.7 //y2=3.7
r117 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=3.7 //y=2.96 //x2=3.7 //y2=3.33
r118 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=3.7 //y=2.59 //x2=3.7 //y2=2.96
r119 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=3.7 //y=2.22 //x2=3.7 //y2=2.59
r120 (  1 30 ) resistor r=32.8556 //w=0.187 //l=0.48 //layer=li \
 //thickness=0.1 //x=3.7 //y=2.22 //x2=3.7 //y2=1.74
ends PM_NOR3X1\%Y

subckt PM_NOR3X1\%noxref_8 ( 7 8 15 16 23 24 25 )
c37 ( 25 0 ) capacitor c=0.0362595f //x=3.885 //y=5.025
c38 ( 24 0 ) capacitor c=0.023843f //x=3.015 //y=5.025
c39 ( 23 0 ) capacitor c=0.0167469f //x=1.965 //y=5.025
c40 ( 16 0 ) capacitor c=0.00239377f //x=3.235 //y=6.91
c41 ( 15 0 ) capacitor c=0.0145111f //x=3.945 //y=6.91
c42 ( 8 0 ) capacitor c=0.00499653f //x=2.195 //y=5.21
c43 ( 7 0 ) capacitor c=0.0417267f //x=3.065 //y=5.21
r44 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.03 //y=6.825 //x2=4.03 //y2=6.74
r45 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.945 //y=6.91 //x2=4.03 //y2=6.825
r46 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.945 //y=6.91 //x2=3.235 //y2=6.91
r47 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.15 //y=6.825 //x2=3.235 //y2=6.91
r48 (  10 24 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.15 //y=6.825 //x2=3.15 //y2=6.74
r49 (  9 24 ) resistor r=52.3636 //w=0.187 //l=0.765 //layer=li \
 //thickness=0.1 //x=3.15 //y=5.295 //x2=3.15 //y2=6.06
r50 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.065 //y=5.21 //x2=3.15 //y2=5.295
r51 (  7 8 ) resistor r=59.5508 //w=0.187 //l=0.87 //layer=li //thickness=0.1 \
 //x=3.065 //y=5.21 //x2=2.195 //y2=5.21
r52 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.295 //x2=2.195 //y2=5.21
r53 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.295 //x2=2.11 //y2=5.72
ends PM_NOR3X1\%noxref_8

