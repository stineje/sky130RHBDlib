* SPICE3 file created from NOR2X1.ext - technology: sky130A

.subckt NOR2X1 Y A B VDD GND
X0 VDD A nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X1 Y B nor2x1_pcell_0/a_317_1331# VDD pshort w=2 l=0.15
X2 Y A GND GND nshort w=3 l=0.15
X3 Y B GND GND nshort w=3 l=0.15
.ends
