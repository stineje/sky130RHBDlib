// File: xnor2x1_pcell.spi.XNOR2X1_PCELL.pxi
// Created: Tue Oct 15 16:01:15 2024
// 
simulator lang=spectre
x_PM_XNOR2X1_PCELL\%noxref_1 ( N_noxref_1_c_6_p N_noxref_1_c_11_p \
 N_noxref_1_c_20_p N_noxref_1_c_138_p N_noxref_1_c_36_p N_noxref_1_c_23_p \
 N_noxref_1_c_29_p N_noxref_1_c_39_p N_noxref_1_c_40_p N_noxref_1_c_75_p \
 N_noxref_1_c_158_p N_noxref_1_c_84_p N_noxref_1_c_96_p N_noxref_1_c_1_p \
 N_noxref_1_c_2_p N_noxref_1_c_3_p N_noxref_1_c_4_p N_noxref_1_c_5_p \
 N_noxref_1_M0_noxref_s N_noxref_1_M1_noxref_d N_noxref_1_M3_noxref_d \
 N_noxref_1_M5_noxref_s )  PM_XNOR2X1_PCELL\%noxref_1
x_PM_XNOR2X1_PCELL\%noxref_2 ( N_noxref_2_c_173_p N_noxref_2_c_174_p \
 N_noxref_2_c_175_p N_noxref_2_c_176_p N_noxref_2_c_195_p N_noxref_2_c_250_p \
 N_noxref_2_c_210_p N_noxref_2_c_236_p N_noxref_2_c_237_p N_noxref_2_c_168_n \
 N_noxref_2_c_169_n N_noxref_2_c_170_n N_noxref_2_c_171_n N_noxref_2_c_172_n \
 N_noxref_2_M6_noxref_s N_noxref_2_M7_noxref_d N_noxref_2_M8_noxref_d \
 N_noxref_2_M12_noxref_d N_noxref_2_M16_noxref_s N_noxref_2_M17_noxref_d )  \
 PM_XNOR2X1_PCELL\%noxref_2
x_PM_XNOR2X1_PCELL\%noxref_3 ( N_noxref_3_c_326_n N_noxref_3_c_328_n \
 N_noxref_3_c_330_n N_noxref_3_c_335_n N_noxref_3_M0_noxref_g \
 N_noxref_3_M1_noxref_g N_noxref_3_M6_noxref_g N_noxref_3_M7_noxref_g \
 N_noxref_3_M8_noxref_g N_noxref_3_M9_noxref_g N_noxref_3_c_336_n \
 N_noxref_3_c_402_p N_noxref_3_c_403_p N_noxref_3_c_338_n N_noxref_3_c_379_n \
 N_noxref_3_c_380_n N_noxref_3_c_339_n N_noxref_3_c_389_p N_noxref_3_c_340_n \
 N_noxref_3_c_342_n N_noxref_3_c_343_n N_noxref_3_c_345_n N_noxref_3_c_421_p \
 N_noxref_3_c_346_n N_noxref_3_c_347_n N_noxref_3_c_348_n N_noxref_3_c_349_n \
 N_noxref_3_c_351_n N_noxref_3_c_352_n N_noxref_3_c_382_n )  \
 PM_XNOR2X1_PCELL\%noxref_3
x_PM_XNOR2X1_PCELL\%noxref_4 ( N_noxref_4_c_459_n N_noxref_4_c_468_n \
 N_noxref_4_c_471_n N_noxref_4_c_510_n N_noxref_4_c_486_n N_noxref_4_c_489_n \
 N_noxref_4_c_474_n N_noxref_4_c_477_n N_noxref_4_M4_noxref_g \
 N_noxref_4_M14_noxref_g N_noxref_4_M15_noxref_g N_noxref_4_c_559_p \
 N_noxref_4_c_560_p N_noxref_4_c_561_p N_noxref_4_c_549_p N_noxref_4_c_563_p \
 N_noxref_4_c_550_p N_noxref_4_c_565_p N_noxref_4_c_551_p N_noxref_4_c_544_p \
 N_noxref_4_M0_noxref_d N_noxref_4_M6_noxref_d )  PM_XNOR2X1_PCELL\%noxref_4
x_PM_XNOR2X1_PCELL\%noxref_5 ( N_noxref_5_c_657_n N_noxref_5_c_655_n \
 N_noxref_5_c_640_n N_noxref_5_c_642_n N_noxref_5_c_628_n N_noxref_5_c_663_n \
 N_noxref_5_c_629_n N_noxref_5_c_645_n N_noxref_5_c_647_n N_noxref_5_c_630_n \
 N_noxref_5_c_676_n N_noxref_5_c_632_n N_noxref_5_M2_noxref_d \
 N_noxref_5_M4_noxref_d N_noxref_5_M10_noxref_d N_noxref_5_M14_noxref_d )  \
 PM_XNOR2X1_PCELL\%noxref_5
x_PM_XNOR2X1_PCELL\%noxref_6 ( N_noxref_6_c_777_n N_noxref_6_c_823_n \
 N_noxref_6_c_795_n N_noxref_6_c_801_n N_noxref_6_c_783_n N_noxref_6_c_803_n \
 N_noxref_6_c_785_n N_noxref_6_c_786_n N_noxref_6_c_787_n N_noxref_6_c_806_n \
 N_noxref_6_c_807_n N_noxref_6_M2_noxref_g N_noxref_6_M12_noxref_g \
 N_noxref_6_M13_noxref_g N_noxref_6_c_826_n N_noxref_6_c_829_n \
 N_noxref_6_c_831_n N_noxref_6_c_834_n N_noxref_6_c_879_n N_noxref_6_c_880_n \
 N_noxref_6_c_836_n N_noxref_6_c_837_n N_noxref_6_c_816_n \
 N_noxref_6_M5_noxref_d N_noxref_6_M16_noxref_d )  PM_XNOR2X1_PCELL\%noxref_6
x_PM_XNOR2X1_PCELL\%noxref_7 ( N_noxref_7_c_976_n N_noxref_7_c_984_n \
 N_noxref_7_c_947_n N_noxref_7_c_1018_n N_noxref_7_c_985_n N_noxref_7_c_950_n \
 N_noxref_7_c_951_n N_noxref_7_M3_noxref_g N_noxref_7_M5_noxref_g \
 N_noxref_7_M10_noxref_g N_noxref_7_M11_noxref_g N_noxref_7_M16_noxref_g \
 N_noxref_7_M17_noxref_g N_noxref_7_c_956_n N_noxref_7_c_958_n \
 N_noxref_7_c_959_n N_noxref_7_c_960_n N_noxref_7_c_961_n N_noxref_7_c_962_n \
 N_noxref_7_c_963_n N_noxref_7_c_965_n N_noxref_7_c_966_n N_noxref_7_c_968_n \
 N_noxref_7_c_1091_n N_noxref_7_c_999_n N_noxref_7_c_969_n N_noxref_7_c_1095_n \
 N_noxref_7_c_1000_n N_noxref_7_c_970_n N_noxref_7_c_1099_n \
 N_noxref_7_c_1100_n N_noxref_7_c_972_n N_noxref_7_c_1011_n N_noxref_7_c_973_n \
 )  PM_XNOR2X1_PCELL\%noxref_7
x_PM_XNOR2X1_PCELL\%noxref_8 ( N_noxref_8_c_1119_n N_noxref_8_c_1124_n \
 N_noxref_8_c_1126_n N_noxref_8_c_1127_n N_noxref_8_M8_noxref_s \
 N_noxref_8_M9_noxref_d N_noxref_8_M11_noxref_d )  PM_XNOR2X1_PCELL\%noxref_8
x_PM_XNOR2X1_PCELL\%noxref_9 ( N_noxref_9_c_1159_n N_noxref_9_c_1160_n \
 N_noxref_9_c_1164_n N_noxref_9_c_1168_n N_noxref_9_c_1169_n \
 N_noxref_9_c_1172_n N_noxref_9_M1_noxref_s )  PM_XNOR2X1_PCELL\%noxref_9
x_PM_XNOR2X1_PCELL\%noxref_10 ( N_noxref_10_c_1211_n N_noxref_10_c_1216_n \
 N_noxref_10_c_1217_n N_noxref_10_c_1218_n N_noxref_10_M12_noxref_s \
 N_noxref_10_M13_noxref_d N_noxref_10_M15_noxref_d )  \
 PM_XNOR2X1_PCELL\%noxref_10
x_PM_XNOR2X1_PCELL\%noxref_11 ( N_noxref_11_c_1278_n N_noxref_11_c_1254_n \
 N_noxref_11_c_1258_n N_noxref_11_c_1262_n N_noxref_11_c_1263_n \
 N_noxref_11_c_1266_n N_noxref_11_M3_noxref_s )  PM_XNOR2X1_PCELL\%noxref_11
cc_1 ( N_noxref_1_c_1_p N_noxref_2_c_168_n ) capacitor c=0.00989031f //x=0.63 \
 //y=0 //x2=0.74 //y2=7.4
cc_2 ( N_noxref_1_c_2_p N_noxref_2_c_169_n ) capacitor c=0.00582097f //x=2.22 \
 //y=0 //x2=2.22 //y2=7.4
cc_3 ( N_noxref_1_c_3_p N_noxref_2_c_170_n ) capacitor c=0.0057235f //x=5.55 \
 //y=0 //x2=5.55 //y2=7.4
cc_4 ( N_noxref_1_c_4_p N_noxref_2_c_171_n ) capacitor c=0.00478842f //x=8.88 \
 //y=0 //x2=8.88 //y2=7.4
cc_5 ( N_noxref_1_c_5_p N_noxref_2_c_172_n ) capacitor c=0.00989031f //x=10.47 \
 //y=0 //x2=10.36 //y2=7.4
cc_6 ( N_noxref_1_c_6_p N_noxref_3_c_326_n ) capacitor c=0.00375416f //x=10.36 \
 //y=0 //x2=3.215 //y2=4.07
cc_7 ( N_noxref_1_c_2_p N_noxref_3_c_326_n ) capacitor c=0.00249386f //x=2.22 \
 //y=0 //x2=3.215 //y2=4.07
cc_8 ( N_noxref_1_c_6_p N_noxref_3_c_328_n ) capacitor c=0.00155455f //x=10.36 \
 //y=0 //x2=0.855 //y2=4.07
cc_9 ( N_noxref_1_M0_noxref_s N_noxref_3_c_328_n ) capacitor c=5.91312e-19 \
 //x=0.495 //y=0.37 //x2=0.855 //y2=4.07
cc_10 ( N_noxref_1_c_6_p N_noxref_3_c_330_n ) capacitor c=0.00187124f \
 //x=10.36 //y=0 //x2=0.74 //y2=2.085
cc_11 ( N_noxref_1_c_11_p N_noxref_3_c_330_n ) capacitor c=8.01092e-19 \
 //x=1.03 //y=0.535 //x2=0.74 //y2=2.085
cc_12 ( N_noxref_1_c_1_p N_noxref_3_c_330_n ) capacitor c=0.028767f //x=0.63 \
 //y=0 //x2=0.74 //y2=2.085
cc_13 ( N_noxref_1_c_2_p N_noxref_3_c_330_n ) capacitor c=0.00133655f //x=2.22 \
 //y=0 //x2=0.74 //y2=2.085
cc_14 ( N_noxref_1_M0_noxref_s N_noxref_3_c_330_n ) capacitor c=0.0110965f \
 //x=0.495 //y=0.37 //x2=0.74 //y2=2.085
cc_15 ( N_noxref_1_c_2_p N_noxref_3_c_335_n ) capacitor c=0.0152607f //x=2.22 \
 //y=0 //x2=3.33 //y2=2.08
cc_16 ( N_noxref_1_c_11_p N_noxref_3_c_336_n ) capacitor c=0.0120496f //x=1.03 \
 //y=0.535 //x2=0.85 //y2=0.91
cc_17 ( N_noxref_1_M0_noxref_s N_noxref_3_c_336_n ) capacitor c=0.0316657f \
 //x=0.495 //y=0.37 //x2=0.85 //y2=0.91
cc_18 ( N_noxref_1_c_1_p N_noxref_3_c_338_n ) capacitor c=0.0124051f //x=0.63 \
 //y=0 //x2=0.85 //y2=1.92
cc_19 ( N_noxref_1_M0_noxref_s N_noxref_3_c_339_n ) capacitor c=0.00483274f \
 //x=0.495 //y=0.37 //x2=1.225 //y2=0.755
cc_20 ( N_noxref_1_c_20_p N_noxref_3_c_340_n ) capacitor c=0.0118602f \
 //x=1.515 //y=0.535 //x2=1.38 //y2=0.91
cc_21 ( N_noxref_1_M0_noxref_s N_noxref_3_c_340_n ) capacitor c=0.0143355f \
 //x=0.495 //y=0.37 //x2=1.38 //y2=0.91
cc_22 ( N_noxref_1_M0_noxref_s N_noxref_3_c_342_n ) capacitor c=0.0074042f \
 //x=0.495 //y=0.37 //x2=1.38 //y2=1.255
cc_23 ( N_noxref_1_c_23_p N_noxref_3_c_343_n ) capacitor c=0.00135046f \
 //x=3.315 //y=0 //x2=3.135 //y2=0.865
cc_24 ( N_noxref_1_M1_noxref_d N_noxref_3_c_343_n ) capacitor c=0.00220047f \
 //x=3.21 //y=0.865 //x2=3.135 //y2=0.865
cc_25 ( N_noxref_1_M1_noxref_d N_noxref_3_c_345_n ) capacitor c=0.00255985f \
 //x=3.21 //y=0.865 //x2=3.135 //y2=1.21
cc_26 ( N_noxref_1_c_2_p N_noxref_3_c_346_n ) capacitor c=0.0114882f //x=2.22 \
 //y=0 //x2=3.135 //y2=1.915
cc_27 ( N_noxref_1_M1_noxref_d N_noxref_3_c_347_n ) capacitor c=0.0131326f \
 //x=3.21 //y=0.865 //x2=3.51 //y2=0.71
cc_28 ( N_noxref_1_M1_noxref_d N_noxref_3_c_348_n ) capacitor c=0.00193127f \
 //x=3.21 //y=0.865 //x2=3.51 //y2=1.365
cc_29 ( N_noxref_1_c_29_p N_noxref_3_c_349_n ) capacitor c=0.00130622f \
 //x=5.38 //y=0 //x2=3.665 //y2=0.865
cc_30 ( N_noxref_1_M1_noxref_d N_noxref_3_c_349_n ) capacitor c=0.00257848f \
 //x=3.21 //y=0.865 //x2=3.665 //y2=0.865
cc_31 ( N_noxref_1_M1_noxref_d N_noxref_3_c_351_n ) capacitor c=0.00255985f \
 //x=3.21 //y=0.865 //x2=3.665 //y2=1.21
cc_32 ( N_noxref_1_c_11_p N_noxref_3_c_352_n ) capacitor c=2.1838e-19 //x=1.03 \
 //y=0.535 //x2=0.74 //y2=2.085
cc_33 ( N_noxref_1_c_1_p N_noxref_3_c_352_n ) capacitor c=0.0108179f //x=0.63 \
 //y=0 //x2=0.74 //y2=2.085
cc_34 ( N_noxref_1_M0_noxref_s N_noxref_3_c_352_n ) capacitor c=0.00655738f \
 //x=0.495 //y=0.37 //x2=0.74 //y2=2.085
cc_35 ( N_noxref_1_c_6_p N_noxref_4_c_459_n ) capacitor c=0.0533435f //x=10.36 \
 //y=0 //x2=7.655 //y2=2.59
cc_36 ( N_noxref_1_c_36_p N_noxref_4_c_459_n ) capacitor c=0.0015622f //x=2.05 \
 //y=0 //x2=7.655 //y2=2.59
cc_37 ( N_noxref_1_c_23_p N_noxref_4_c_459_n ) capacitor c=0.00280978f \
 //x=3.315 //y=0 //x2=7.655 //y2=2.59
cc_38 ( N_noxref_1_c_29_p N_noxref_4_c_459_n ) capacitor c=0.00345949f \
 //x=5.38 //y=0 //x2=7.655 //y2=2.59
cc_39 ( N_noxref_1_c_39_p N_noxref_4_c_459_n ) capacitor c=0.00280978f \
 //x=6.645 //y=0 //x2=7.655 //y2=2.59
cc_40 ( N_noxref_1_c_40_p N_noxref_4_c_459_n ) capacitor c=9.24405e-19 \
 //x=8.71 //y=0 //x2=7.655 //y2=2.59
cc_41 ( N_noxref_1_c_2_p N_noxref_4_c_459_n ) capacitor c=0.038878f //x=2.22 \
 //y=0 //x2=7.655 //y2=2.59
cc_42 ( N_noxref_1_c_3_p N_noxref_4_c_459_n ) capacitor c=0.0338055f //x=5.55 \
 //y=0 //x2=7.655 //y2=2.59
cc_43 ( N_noxref_1_M0_noxref_s N_noxref_4_c_459_n ) capacitor c=0.00248261f \
 //x=0.495 //y=0.37 //x2=7.655 //y2=2.59
cc_44 ( N_noxref_1_c_6_p N_noxref_4_c_468_n ) capacitor c=0.00231366f \
 //x=10.36 //y=0 //x2=1.595 //y2=2.59
cc_45 ( N_noxref_1_c_2_p N_noxref_4_c_468_n ) capacitor c=0.00209945f //x=2.22 \
 //y=0 //x2=1.595 //y2=2.59
cc_46 ( N_noxref_1_M0_noxref_s N_noxref_4_c_468_n ) capacitor c=0.00120637f \
 //x=0.495 //y=0.37 //x2=1.595 //y2=2.59
cc_47 ( N_noxref_1_c_6_p N_noxref_4_c_471_n ) capacitor c=0.00129718f \
 //x=10.36 //y=0 //x2=1.395 //y2=2.08
cc_48 ( N_noxref_1_c_2_p N_noxref_4_c_471_n ) capacitor c=0.0263587f //x=2.22 \
 //y=0 //x2=1.395 //y2=2.08
cc_49 ( N_noxref_1_M0_noxref_s N_noxref_4_c_471_n ) capacitor c=0.00949589f \
 //x=0.495 //y=0.37 //x2=1.395 //y2=2.08
cc_50 ( N_noxref_1_c_1_p N_noxref_4_c_474_n ) capacitor c=9.71e-19 //x=0.63 \
 //y=0 //x2=1.48 //y2=2.59
cc_51 ( N_noxref_1_c_2_p N_noxref_4_c_474_n ) capacitor c=5.56859e-19 //x=2.22 \
 //y=0 //x2=1.48 //y2=2.59
cc_52 ( N_noxref_1_M0_noxref_s N_noxref_4_c_474_n ) capacitor c=2.30929e-19 \
 //x=0.495 //y=0.37 //x2=1.48 //y2=2.59
cc_53 ( N_noxref_1_c_3_p N_noxref_4_c_477_n ) capacitor c=6.92592e-19 //x=5.55 \
 //y=0 //x2=7.77 //y2=2.08
cc_54 ( N_noxref_1_c_4_p N_noxref_4_c_477_n ) capacitor c=0.00185226f //x=8.88 \
 //y=0 //x2=7.77 //y2=2.08
cc_55 ( N_noxref_1_c_6_p N_noxref_4_M0_noxref_d ) capacitor c=0.00136354f \
 //x=10.36 //y=0 //x2=0.925 //y2=0.91
cc_56 ( N_noxref_1_c_11_p N_noxref_4_M0_noxref_d ) capacitor c=0.0151737f \
 //x=1.03 //y=0.535 //x2=0.925 //y2=0.91
cc_57 ( N_noxref_1_c_1_p N_noxref_4_M0_noxref_d ) capacitor c=0.0094373f \
 //x=0.63 //y=0 //x2=0.925 //y2=0.91
cc_58 ( N_noxref_1_c_2_p N_noxref_4_M0_noxref_d ) capacitor c=0.00949241f \
 //x=2.22 //y=0 //x2=0.925 //y2=0.91
cc_59 ( N_noxref_1_c_5_p N_noxref_4_M0_noxref_d ) capacitor c=2.29264e-19 \
 //x=10.47 //y=0 //x2=0.925 //y2=0.91
cc_60 ( N_noxref_1_M0_noxref_s N_noxref_4_M0_noxref_d ) capacitor c=0.076995f \
 //x=0.495 //y=0.37 //x2=0.925 //y2=0.91
cc_61 ( N_noxref_1_c_3_p N_noxref_5_c_628_n ) capacitor c=0.0430893f //x=5.55 \
 //y=0 //x2=4.725 //y2=1.65
cc_62 ( N_noxref_1_c_2_p N_noxref_5_c_629_n ) capacitor c=0.00105873f //x=2.22 \
 //y=0 //x2=4.81 //y2=3.7
cc_63 ( N_noxref_1_c_4_p N_noxref_5_c_630_n ) capacitor c=0.0448856f //x=8.88 \
 //y=0 //x2=8.055 //y2=1.65
cc_64 ( N_noxref_1_M5_noxref_s N_noxref_5_c_630_n ) capacitor c=3.53049e-19 \
 //x=9.375 //y=0.37 //x2=8.055 //y2=1.65
cc_65 ( N_noxref_1_c_3_p N_noxref_5_c_632_n ) capacitor c=0.00100332f //x=5.55 \
 //y=0 //x2=8.14 //y2=3.7
cc_66 ( N_noxref_1_c_2_p N_noxref_5_M2_noxref_d ) capacitor c=8.60262e-19 \
 //x=2.22 //y=0 //x2=4.18 //y2=0.905
cc_67 ( N_noxref_1_c_3_p N_noxref_5_M2_noxref_d ) capacitor c=0.00605305f \
 //x=5.55 //y=0 //x2=4.18 //y2=0.905
cc_68 ( N_noxref_1_M1_noxref_d N_noxref_5_M2_noxref_d ) capacitor \
 c=0.00143464f //x=3.21 //y=0.865 //x2=4.18 //y2=0.905
cc_69 ( N_noxref_1_c_3_p N_noxref_5_M4_noxref_d ) capacitor c=8.60262e-19 \
 //x=5.55 //y=0 //x2=7.51 //y2=0.905
cc_70 ( N_noxref_1_c_4_p N_noxref_5_M4_noxref_d ) capacitor c=0.00605305f \
 //x=8.88 //y=0 //x2=7.51 //y2=0.905
cc_71 ( N_noxref_1_M3_noxref_d N_noxref_5_M4_noxref_d ) capacitor \
 c=0.00143464f //x=6.54 //y=0.865 //x2=7.51 //y2=0.905
cc_72 ( N_noxref_1_M5_noxref_s N_noxref_5_M4_noxref_d ) capacitor \
 c=2.07711e-19 //x=9.375 //y=0.37 //x2=7.51 //y2=0.905
cc_73 ( N_noxref_1_c_6_p N_noxref_6_c_777_n ) capacitor c=0.0292011f //x=10.36 \
 //y=0 //x2=9.505 //y2=2.96
cc_74 ( N_noxref_1_c_40_p N_noxref_6_c_777_n ) capacitor c=0.00208984f \
 //x=8.71 //y=0 //x2=9.505 //y2=2.96
cc_75 ( N_noxref_1_c_75_p N_noxref_6_c_777_n ) capacitor c=0.00129597f \
 //x=9.415 //y=0 //x2=9.505 //y2=2.96
cc_76 ( N_noxref_1_c_3_p N_noxref_6_c_777_n ) capacitor c=0.00750857f //x=5.55 \
 //y=0 //x2=9.505 //y2=2.96
cc_77 ( N_noxref_1_c_4_p N_noxref_6_c_777_n ) capacitor c=0.0144849f //x=8.88 \
 //y=0 //x2=9.505 //y2=2.96
cc_78 ( N_noxref_1_M5_noxref_s N_noxref_6_c_777_n ) capacitor c=0.00263458f \
 //x=9.375 //y=0.37 //x2=9.505 //y2=2.96
cc_79 ( N_noxref_1_c_2_p N_noxref_6_c_783_n ) capacitor c=7.03122e-19 //x=2.22 \
 //y=0 //x2=4.44 //y2=2.08
cc_80 ( N_noxref_1_c_3_p N_noxref_6_c_783_n ) capacitor c=0.00165751f //x=5.55 \
 //y=0 //x2=4.44 //y2=2.08
cc_81 ( N_noxref_1_c_5_p N_noxref_6_c_785_n ) capacitor c=0.00114558f \
 //x=10.47 //y=0 //x2=9.62 //y2=2.96
cc_82 ( N_noxref_1_M5_noxref_s N_noxref_6_c_786_n ) capacitor c=0.00178664f \
 //x=9.375 //y=0.37 //x2=9.905 //y2=2.08
cc_83 ( N_noxref_1_c_6_p N_noxref_6_c_787_n ) capacitor c=0.00128871f \
 //x=10.36 //y=0 //x2=9.705 //y2=2.08
cc_84 ( N_noxref_1_c_84_p N_noxref_6_c_787_n ) capacitor c=0.00178664f //x=9.9 \
 //y=0.535 //x2=9.705 //y2=2.08
cc_85 ( N_noxref_1_c_4_p N_noxref_6_c_787_n ) capacitor c=0.0291959f //x=8.88 \
 //y=0 //x2=9.705 //y2=2.08
cc_86 ( N_noxref_1_M5_noxref_s N_noxref_6_c_787_n ) capacitor c=0.00570196f \
 //x=9.375 //y=0.37 //x2=9.705 //y2=2.08
cc_87 ( N_noxref_1_c_6_p N_noxref_6_M5_noxref_d ) capacitor c=0.00128496f \
 //x=10.36 //y=0 //x2=9.795 //y2=0.91
cc_88 ( N_noxref_1_c_4_p N_noxref_6_M5_noxref_d ) capacitor c=0.00945919f \
 //x=8.88 //y=0 //x2=9.795 //y2=0.91
cc_89 ( N_noxref_1_c_5_p N_noxref_6_M5_noxref_d ) capacitor c=0.00966656f \
 //x=10.47 //y=0 //x2=9.795 //y2=0.91
cc_90 ( N_noxref_1_M5_noxref_s N_noxref_6_M5_noxref_d ) capacitor c=0.0920885f \
 //x=9.375 //y=0.37 //x2=9.795 //y2=0.91
cc_91 ( N_noxref_1_c_6_p N_noxref_7_c_947_n ) capacitor c=0.0127184f //x=10.36 \
 //y=0 //x2=10.245 //y2=3.33
cc_92 ( N_noxref_1_c_84_p N_noxref_7_c_947_n ) capacitor c=8.90535e-19 //x=9.9 \
 //y=0.535 //x2=10.245 //y2=3.33
cc_93 ( N_noxref_1_M5_noxref_s N_noxref_7_c_947_n ) capacitor c=0.00106019f \
 //x=9.375 //y=0.37 //x2=10.245 //y2=3.33
cc_94 ( N_noxref_1_c_3_p N_noxref_7_c_950_n ) capacitor c=0.0152684f //x=5.55 \
 //y=0 //x2=6.66 //y2=2.08
cc_95 ( N_noxref_1_c_6_p N_noxref_7_c_951_n ) capacitor c=0.00184963f \
 //x=10.36 //y=0 //x2=10.36 //y2=2.085
cc_96 ( N_noxref_1_c_96_p N_noxref_7_c_951_n ) capacitor c=7.87839e-19 \
 //x=10.385 //y=0.535 //x2=10.36 //y2=2.085
cc_97 ( N_noxref_1_c_4_p N_noxref_7_c_951_n ) capacitor c=0.00146529f //x=8.88 \
 //y=0 //x2=10.36 //y2=2.085
cc_98 ( N_noxref_1_c_5_p N_noxref_7_c_951_n ) capacitor c=0.0290276f //x=10.47 \
 //y=0 //x2=10.36 //y2=2.085
cc_99 ( N_noxref_1_M5_noxref_s N_noxref_7_c_951_n ) capacitor c=0.0109271f \
 //x=9.375 //y=0.37 //x2=10.36 //y2=2.085
cc_100 ( N_noxref_1_c_39_p N_noxref_7_c_956_n ) capacitor c=0.00135046f \
 //x=6.645 //y=0 //x2=6.465 //y2=0.865
cc_101 ( N_noxref_1_M3_noxref_d N_noxref_7_c_956_n ) capacitor c=0.00220047f \
 //x=6.54 //y=0.865 //x2=6.465 //y2=0.865
cc_102 ( N_noxref_1_M3_noxref_d N_noxref_7_c_958_n ) capacitor c=0.00255985f \
 //x=6.54 //y=0.865 //x2=6.465 //y2=1.21
cc_103 ( N_noxref_1_c_3_p N_noxref_7_c_959_n ) capacitor c=0.00176175f \
 //x=5.55 //y=0 //x2=6.465 //y2=1.52
cc_104 ( N_noxref_1_c_3_p N_noxref_7_c_960_n ) capacitor c=0.0114882f //x=5.55 \
 //y=0 //x2=6.465 //y2=1.915
cc_105 ( N_noxref_1_M3_noxref_d N_noxref_7_c_961_n ) capacitor c=0.0131326f \
 //x=6.54 //y=0.865 //x2=6.84 //y2=0.71
cc_106 ( N_noxref_1_M3_noxref_d N_noxref_7_c_962_n ) capacitor c=0.00193127f \
 //x=6.54 //y=0.865 //x2=6.84 //y2=1.365
cc_107 ( N_noxref_1_c_40_p N_noxref_7_c_963_n ) capacitor c=0.00130622f \
 //x=8.71 //y=0 //x2=6.995 //y2=0.865
cc_108 ( N_noxref_1_M3_noxref_d N_noxref_7_c_963_n ) capacitor c=0.00257848f \
 //x=6.54 //y=0.865 //x2=6.995 //y2=0.865
cc_109 ( N_noxref_1_M3_noxref_d N_noxref_7_c_965_n ) capacitor c=0.00255985f \
 //x=6.54 //y=0.865 //x2=6.995 //y2=1.21
cc_110 ( N_noxref_1_c_84_p N_noxref_7_c_966_n ) capacitor c=0.0119174f //x=9.9 \
 //y=0.535 //x2=9.72 //y2=0.91
cc_111 ( N_noxref_1_M5_noxref_s N_noxref_7_c_966_n ) capacitor c=0.0143355f \
 //x=9.375 //y=0.37 //x2=9.72 //y2=0.91
cc_112 ( N_noxref_1_M5_noxref_s N_noxref_7_c_968_n ) capacitor c=0.0074042f \
 //x=9.375 //y=0.37 //x2=9.72 //y2=1.255
cc_113 ( N_noxref_1_M5_noxref_s N_noxref_7_c_969_n ) capacitor c=0.00489f \
 //x=9.375 //y=0.37 //x2=10.095 //y2=0.755
cc_114 ( N_noxref_1_c_96_p N_noxref_7_c_970_n ) capacitor c=0.0123171f \
 //x=10.385 //y=0.535 //x2=10.25 //y2=0.91
cc_115 ( N_noxref_1_M5_noxref_s N_noxref_7_c_970_n ) capacitor c=0.0318096f \
 //x=9.375 //y=0.37 //x2=10.25 //y2=0.91
cc_116 ( N_noxref_1_c_5_p N_noxref_7_c_972_n ) capacitor c=0.0124811f \
 //x=10.47 //y=0 //x2=10.25 //y2=1.92
cc_117 ( N_noxref_1_c_96_p N_noxref_7_c_973_n ) capacitor c=2.1838e-19 \
 //x=10.385 //y=0.535 //x2=10.25 //y2=2.085
cc_118 ( N_noxref_1_c_5_p N_noxref_7_c_973_n ) capacitor c=0.0108179f \
 //x=10.47 //y=0 //x2=10.25 //y2=2.085
cc_119 ( N_noxref_1_M5_noxref_s N_noxref_7_c_973_n ) capacitor c=0.00655738f \
 //x=9.375 //y=0.37 //x2=10.25 //y2=2.085
cc_120 ( N_noxref_1_M0_noxref_s N_noxref_9_c_1159_n ) capacitor c=0.0013253f \
 //x=0.495 //y=0.37 //x2=2.915 //y2=1.495
cc_121 ( N_noxref_1_c_6_p N_noxref_9_c_1160_n ) capacitor c=0.00530453f \
 //x=10.36 //y=0 //x2=3.8 //y2=1.58
cc_122 ( N_noxref_1_c_23_p N_noxref_9_c_1160_n ) capacitor c=0.00112921f \
 //x=3.315 //y=0 //x2=3.8 //y2=1.58
cc_123 ( N_noxref_1_c_29_p N_noxref_9_c_1160_n ) capacitor c=0.00182339f \
 //x=5.38 //y=0 //x2=3.8 //y2=1.58
cc_124 ( N_noxref_1_M1_noxref_d N_noxref_9_c_1160_n ) capacitor c=0.00879185f \
 //x=3.21 //y=0.865 //x2=3.8 //y2=1.58
cc_125 ( N_noxref_1_c_6_p N_noxref_9_c_1164_n ) capacitor c=0.00271584f \
 //x=10.36 //y=0 //x2=3.885 //y2=0.615
cc_126 ( N_noxref_1_c_29_p N_noxref_9_c_1164_n ) capacitor c=0.014783f \
 //x=5.38 //y=0 //x2=3.885 //y2=0.615
cc_127 ( N_noxref_1_c_5_p N_noxref_9_c_1164_n ) capacitor c=0.00145873f \
 //x=10.47 //y=0 //x2=3.885 //y2=0.615
cc_128 ( N_noxref_1_M1_noxref_d N_noxref_9_c_1164_n ) capacitor c=0.033812f \
 //x=3.21 //y=0.865 //x2=3.885 //y2=0.615
cc_129 ( N_noxref_1_c_2_p N_noxref_9_c_1168_n ) capacitor c=2.91423e-19 \
 //x=2.22 //y=0 //x2=3.885 //y2=1.495
cc_130 ( N_noxref_1_c_6_p N_noxref_9_c_1169_n ) capacitor c=0.0111902f \
 //x=10.36 //y=0 //x2=4.77 //y2=0.53
cc_131 ( N_noxref_1_c_29_p N_noxref_9_c_1169_n ) capacitor c=0.0375381f \
 //x=5.38 //y=0 //x2=4.77 //y2=0.53
cc_132 ( N_noxref_1_c_5_p N_noxref_9_c_1169_n ) capacitor c=0.00199432f \
 //x=10.47 //y=0 //x2=4.77 //y2=0.53
cc_133 ( N_noxref_1_c_6_p N_noxref_9_c_1172_n ) capacitor c=0.00271457f \
 //x=10.36 //y=0 //x2=4.855 //y2=0.615
cc_134 ( N_noxref_1_c_29_p N_noxref_9_c_1172_n ) capacitor c=0.0147189f \
 //x=5.38 //y=0 //x2=4.855 //y2=0.615
cc_135 ( N_noxref_1_c_3_p N_noxref_9_c_1172_n ) capacitor c=0.0431718f \
 //x=5.55 //y=0 //x2=4.855 //y2=0.615
cc_136 ( N_noxref_1_c_5_p N_noxref_9_c_1172_n ) capacitor c=0.00145015f \
 //x=10.47 //y=0 //x2=4.855 //y2=0.615
cc_137 ( N_noxref_1_c_6_p N_noxref_9_M1_noxref_s ) capacitor c=0.00271584f \
 //x=10.36 //y=0 //x2=2.78 //y2=0.365
cc_138 ( N_noxref_1_c_138_p N_noxref_9_M1_noxref_s ) capacitor c=0.0013253f \
 //x=1.6 //y=0.45 //x2=2.78 //y2=0.365
cc_139 ( N_noxref_1_c_23_p N_noxref_9_M1_noxref_s ) capacitor c=0.014783f \
 //x=3.315 //y=0 //x2=2.78 //y2=0.365
cc_140 ( N_noxref_1_c_2_p N_noxref_9_M1_noxref_s ) capacitor c=0.058339f \
 //x=2.22 //y=0 //x2=2.78 //y2=0.365
cc_141 ( N_noxref_1_c_3_p N_noxref_9_M1_noxref_s ) capacitor c=0.00200438f \
 //x=5.55 //y=0 //x2=2.78 //y2=0.365
cc_142 ( N_noxref_1_c_5_p N_noxref_9_M1_noxref_s ) capacitor c=0.00145873f \
 //x=10.47 //y=0 //x2=2.78 //y2=0.365
cc_143 ( N_noxref_1_M1_noxref_d N_noxref_9_M1_noxref_s ) capacitor \
 c=0.0334197f //x=3.21 //y=0.865 //x2=2.78 //y2=0.365
cc_144 ( N_noxref_1_c_6_p N_noxref_11_c_1254_n ) capacitor c=0.00530453f \
 //x=10.36 //y=0 //x2=7.13 //y2=1.58
cc_145 ( N_noxref_1_c_39_p N_noxref_11_c_1254_n ) capacitor c=0.00112921f \
 //x=6.645 //y=0 //x2=7.13 //y2=1.58
cc_146 ( N_noxref_1_c_40_p N_noxref_11_c_1254_n ) capacitor c=0.00182339f \
 //x=8.71 //y=0 //x2=7.13 //y2=1.58
cc_147 ( N_noxref_1_M3_noxref_d N_noxref_11_c_1254_n ) capacitor c=0.00879185f \
 //x=6.54 //y=0.865 //x2=7.13 //y2=1.58
cc_148 ( N_noxref_1_c_6_p N_noxref_11_c_1258_n ) capacitor c=0.00271584f \
 //x=10.36 //y=0 //x2=7.215 //y2=0.615
cc_149 ( N_noxref_1_c_40_p N_noxref_11_c_1258_n ) capacitor c=0.014783f \
 //x=8.71 //y=0 //x2=7.215 //y2=0.615
cc_150 ( N_noxref_1_c_5_p N_noxref_11_c_1258_n ) capacitor c=0.00145873f \
 //x=10.47 //y=0 //x2=7.215 //y2=0.615
cc_151 ( N_noxref_1_M3_noxref_d N_noxref_11_c_1258_n ) capacitor c=0.033812f \
 //x=6.54 //y=0.865 //x2=7.215 //y2=0.615
cc_152 ( N_noxref_1_c_3_p N_noxref_11_c_1262_n ) capacitor c=2.91423e-19 \
 //x=5.55 //y=0 //x2=7.215 //y2=1.495
cc_153 ( N_noxref_1_c_6_p N_noxref_11_c_1263_n ) capacitor c=0.0112826f \
 //x=10.36 //y=0 //x2=8.1 //y2=0.53
cc_154 ( N_noxref_1_c_40_p N_noxref_11_c_1263_n ) capacitor c=0.037559f \
 //x=8.71 //y=0 //x2=8.1 //y2=0.53
cc_155 ( N_noxref_1_c_5_p N_noxref_11_c_1263_n ) capacitor c=0.00199432f \
 //x=10.47 //y=0 //x2=8.1 //y2=0.53
cc_156 ( N_noxref_1_c_6_p N_noxref_11_c_1266_n ) capacitor c=0.00282863f \
 //x=10.36 //y=0 //x2=8.185 //y2=0.615
cc_157 ( N_noxref_1_c_40_p N_noxref_11_c_1266_n ) capacitor c=0.0148003f \
 //x=8.71 //y=0 //x2=8.185 //y2=0.615
cc_158 ( N_noxref_1_c_158_p N_noxref_11_c_1266_n ) capacitor c=9.92084e-19 \
 //x=9.5 //y=0.45 //x2=8.185 //y2=0.615
cc_159 ( N_noxref_1_c_4_p N_noxref_11_c_1266_n ) capacitor c=0.0431718f \
 //x=8.88 //y=0 //x2=8.185 //y2=0.615
cc_160 ( N_noxref_1_c_5_p N_noxref_11_c_1266_n ) capacitor c=0.00145015f \
 //x=10.47 //y=0 //x2=8.185 //y2=0.615
cc_161 ( N_noxref_1_c_6_p N_noxref_11_M3_noxref_s ) capacitor c=0.00271584f \
 //x=10.36 //y=0 //x2=6.11 //y2=0.365
cc_162 ( N_noxref_1_c_39_p N_noxref_11_M3_noxref_s ) capacitor c=0.014783f \
 //x=6.645 //y=0 //x2=6.11 //y2=0.365
cc_163 ( N_noxref_1_c_3_p N_noxref_11_M3_noxref_s ) capacitor c=0.058339f \
 //x=5.55 //y=0 //x2=6.11 //y2=0.365
cc_164 ( N_noxref_1_c_4_p N_noxref_11_M3_noxref_s ) capacitor c=0.00200548f \
 //x=8.88 //y=0 //x2=6.11 //y2=0.365
cc_165 ( N_noxref_1_c_5_p N_noxref_11_M3_noxref_s ) capacitor c=0.00145873f \
 //x=10.47 //y=0 //x2=6.11 //y2=0.365
cc_166 ( N_noxref_1_M3_noxref_d N_noxref_11_M3_noxref_s ) capacitor \
 c=0.0334197f //x=6.54 //y=0.865 //x2=6.11 //y2=0.365
cc_167 ( N_noxref_1_M5_noxref_s N_noxref_11_M3_noxref_s ) capacitor \
 c=9.92084e-19 //x=9.375 //y=0.37 //x2=6.11 //y2=0.365
cc_168 ( N_noxref_2_c_173_p N_noxref_3_c_326_n ) capacitor c=0.0179155f \
 //x=10.36 //y=7.4 //x2=3.215 //y2=4.07
cc_169 ( N_noxref_2_c_174_p N_noxref_3_c_326_n ) capacitor c=9.77842e-19 \
 //x=1.47 //y=7.4 //x2=3.215 //y2=4.07
cc_170 ( N_noxref_2_c_175_p N_noxref_3_c_326_n ) capacitor c=0.00124367f \
 //x=2.05 //y=7.4 //x2=3.215 //y2=4.07
cc_171 ( N_noxref_2_c_176_p N_noxref_3_c_326_n ) capacitor c=0.00216965f \
 //x=3.365 //y=7.4 //x2=3.215 //y2=4.07
cc_172 ( N_noxref_2_c_169_n N_noxref_3_c_326_n ) capacitor c=0.0280406f \
 //x=2.22 //y=7.4 //x2=3.215 //y2=4.07
cc_173 ( N_noxref_2_M7_noxref_d N_noxref_3_c_326_n ) capacitor c=0.00213856f \
 //x=1.41 //y=5.02 //x2=3.215 //y2=4.07
cc_174 ( N_noxref_2_c_173_p N_noxref_3_c_328_n ) capacitor c=0.00188164f \
 //x=10.36 //y=7.4 //x2=0.855 //y2=4.07
cc_175 ( N_noxref_2_c_168_n N_noxref_3_c_328_n ) capacitor c=0.00208272f \
 //x=0.74 //y=7.4 //x2=0.855 //y2=4.07
cc_176 ( N_noxref_2_M6_noxref_s N_noxref_3_c_328_n ) capacitor c=0.00185024f \
 //x=0.54 //y=5.02 //x2=0.855 //y2=4.07
cc_177 ( N_noxref_2_c_173_p N_noxref_3_c_330_n ) capacitor c=0.00157744f \
 //x=10.36 //y=7.4 //x2=0.74 //y2=2.085
cc_178 ( N_noxref_2_c_168_n N_noxref_3_c_330_n ) capacitor c=0.0272385f \
 //x=0.74 //y=7.4 //x2=0.74 //y2=2.085
cc_179 ( N_noxref_2_c_169_n N_noxref_3_c_330_n ) capacitor c=0.00139956f \
 //x=2.22 //y=7.4 //x2=0.74 //y2=2.085
cc_180 ( N_noxref_2_M6_noxref_s N_noxref_3_c_330_n ) capacitor c=0.00896093f \
 //x=0.54 //y=5.02 //x2=0.74 //y2=2.085
cc_181 ( N_noxref_2_c_169_n N_noxref_3_c_335_n ) capacitor c=0.0160048f \
 //x=2.22 //y=7.4 //x2=3.33 //y2=2.08
cc_182 ( N_noxref_2_c_174_p N_noxref_3_M6_noxref_g ) capacitor c=0.00748034f \
 //x=1.47 //y=7.4 //x2=0.895 //y2=6.02
cc_183 ( N_noxref_2_c_168_n N_noxref_3_M6_noxref_g ) capacitor c=0.0241676f \
 //x=0.74 //y=7.4 //x2=0.895 //y2=6.02
cc_184 ( N_noxref_2_M6_noxref_s N_noxref_3_M6_noxref_g ) capacitor \
 c=0.0528676f //x=0.54 //y=5.02 //x2=0.895 //y2=6.02
cc_185 ( N_noxref_2_c_174_p N_noxref_3_M7_noxref_g ) capacitor c=0.00697478f \
 //x=1.47 //y=7.4 //x2=1.335 //y2=6.02
cc_186 ( N_noxref_2_M7_noxref_d N_noxref_3_M7_noxref_g ) capacitor \
 c=0.0528676f //x=1.41 //y=5.02 //x2=1.335 //y2=6.02
cc_187 ( N_noxref_2_c_176_p N_noxref_3_M8_noxref_g ) capacitor c=0.00673447f \
 //x=3.365 //y=7.4 //x2=3.23 //y2=6.02
cc_188 ( N_noxref_2_c_169_n N_noxref_3_M8_noxref_g ) capacitor c=0.00449901f \
 //x=2.22 //y=7.4 //x2=3.23 //y2=6.02
cc_189 ( N_noxref_2_M8_noxref_d N_noxref_3_M8_noxref_g ) capacitor \
 c=0.0166176f //x=3.305 //y=5.02 //x2=3.23 //y2=6.02
cc_190 ( N_noxref_2_c_195_p N_noxref_3_M9_noxref_g ) capacitor c=0.006727f \
 //x=5.38 //y=7.4 //x2=3.67 //y2=6.02
cc_191 ( N_noxref_2_M8_noxref_d N_noxref_3_M9_noxref_g ) capacitor \
 c=0.0186652f //x=3.305 //y=5.02 //x2=3.67 //y2=6.02
cc_192 ( N_noxref_2_c_169_n N_noxref_3_c_379_n ) capacitor c=0.0132667f \
 //x=2.22 //y=7.4 //x2=1.26 //y2=4.79
cc_193 ( N_noxref_2_c_168_n N_noxref_3_c_380_n ) capacitor c=0.011132f \
 //x=0.74 //y=7.4 //x2=0.97 //y2=4.79
cc_194 ( N_noxref_2_M6_noxref_s N_noxref_3_c_380_n ) capacitor c=0.00524527f \
 //x=0.54 //y=5.02 //x2=0.97 //y2=4.79
cc_195 ( N_noxref_2_c_169_n N_noxref_3_c_382_n ) capacitor c=0.0125867f \
 //x=2.22 //y=7.4 //x2=3.33 //y2=4.7
cc_196 ( N_noxref_2_c_169_n N_noxref_4_c_459_n ) capacitor c=0.00137387f \
 //x=2.22 //y=7.4 //x2=7.655 //y2=2.59
cc_197 ( N_noxref_2_c_173_p N_noxref_4_c_486_n ) capacitor c=0.0012271f \
 //x=10.36 //y=7.4 //x2=1.395 //y2=4.58
cc_198 ( N_noxref_2_c_174_p N_noxref_4_c_486_n ) capacitor c=9.08147e-19 \
 //x=1.47 //y=7.4 //x2=1.395 //y2=4.58
cc_199 ( N_noxref_2_M7_noxref_d N_noxref_4_c_486_n ) capacitor c=0.00609088f \
 //x=1.41 //y=5.02 //x2=1.395 //y2=4.58
cc_200 ( N_noxref_2_c_168_n N_noxref_4_c_489_n ) capacitor c=0.0179238f \
 //x=0.74 //y=7.4 //x2=1.2 //y2=4.58
cc_201 ( N_noxref_2_c_168_n N_noxref_4_c_474_n ) capacitor c=5.65246e-19 \
 //x=0.74 //y=7.4 //x2=1.48 //y2=2.59
cc_202 ( N_noxref_2_c_169_n N_noxref_4_c_474_n ) capacitor c=0.0220651f \
 //x=2.22 //y=7.4 //x2=1.48 //y2=2.59
cc_203 ( N_noxref_2_c_170_n N_noxref_4_c_477_n ) capacitor c=0.00210246f \
 //x=5.55 //y=7.4 //x2=7.77 //y2=2.08
cc_204 ( N_noxref_2_c_171_n N_noxref_4_c_477_n ) capacitor c=0.00147437f \
 //x=8.88 //y=7.4 //x2=7.77 //y2=2.08
cc_205 ( N_noxref_2_c_210_p N_noxref_4_M14_noxref_g ) capacitor c=0.00510247f \
 //x=8.71 //y=7.4 //x2=7.44 //y2=6.02
cc_206 ( N_noxref_2_c_210_p N_noxref_4_M15_noxref_g ) capacitor c=0.00510919f \
 //x=8.71 //y=7.4 //x2=7.88 //y2=6.02
cc_207 ( N_noxref_2_c_171_n N_noxref_4_M15_noxref_g ) capacitor c=0.00788519f \
 //x=8.88 //y=7.4 //x2=7.88 //y2=6.02
cc_208 ( N_noxref_2_c_173_p N_noxref_4_M6_noxref_d ) capacitor c=0.00285171f \
 //x=10.36 //y=7.4 //x2=0.97 //y2=5.02
cc_209 ( N_noxref_2_c_174_p N_noxref_4_M6_noxref_d ) capacitor c=0.0141332f \
 //x=1.47 //y=7.4 //x2=0.97 //y2=5.02
cc_210 ( N_noxref_2_c_169_n N_noxref_4_M6_noxref_d ) capacitor c=0.0204646f \
 //x=2.22 //y=7.4 //x2=0.97 //y2=5.02
cc_211 ( N_noxref_2_c_172_n N_noxref_4_M6_noxref_d ) capacitor c=0.00135976f \
 //x=10.36 //y=7.4 //x2=0.97 //y2=5.02
cc_212 ( N_noxref_2_M6_noxref_s N_noxref_4_M6_noxref_d ) capacitor \
 c=0.0843065f //x=0.54 //y=5.02 //x2=0.97 //y2=5.02
cc_213 ( N_noxref_2_M7_noxref_d N_noxref_4_M6_noxref_d ) capacitor \
 c=0.0832641f //x=1.41 //y=5.02 //x2=0.97 //y2=5.02
cc_214 ( N_noxref_2_c_173_p N_noxref_5_c_640_n ) capacitor c=0.00114116f \
 //x=10.36 //y=7.4 //x2=4.725 //y2=5.205
cc_215 ( N_noxref_2_c_195_p N_noxref_5_c_640_n ) capacitor c=0.0013904f \
 //x=5.38 //y=7.4 //x2=4.725 //y2=5.205
cc_216 ( N_noxref_2_c_169_n N_noxref_5_c_642_n ) capacitor c=8.9933e-19 \
 //x=2.22 //y=7.4 //x2=4.415 //y2=5.205
cc_217 ( N_noxref_2_c_169_n N_noxref_5_c_629_n ) capacitor c=0.00163766f \
 //x=2.22 //y=7.4 //x2=4.81 //y2=3.7
cc_218 ( N_noxref_2_c_170_n N_noxref_5_c_629_n ) capacitor c=0.0445615f \
 //x=5.55 //y=7.4 //x2=4.81 //y2=3.7
cc_219 ( N_noxref_2_c_173_p N_noxref_5_c_645_n ) capacitor c=0.00113725f \
 //x=10.36 //y=7.4 //x2=8.055 //y2=5.205
cc_220 ( N_noxref_2_c_210_p N_noxref_5_c_645_n ) capacitor c=0.00138981f \
 //x=8.71 //y=7.4 //x2=8.055 //y2=5.205
cc_221 ( N_noxref_2_c_170_n N_noxref_5_c_647_n ) capacitor c=8.9933e-19 \
 //x=5.55 //y=7.4 //x2=7.745 //y2=5.205
cc_222 ( N_noxref_2_c_170_n N_noxref_5_c_632_n ) capacitor c=0.00177938f \
 //x=5.55 //y=7.4 //x2=8.14 //y2=3.7
cc_223 ( N_noxref_2_c_171_n N_noxref_5_c_632_n ) capacitor c=0.0420694f \
 //x=8.88 //y=7.4 //x2=8.14 //y2=3.7
cc_224 ( N_noxref_2_c_170_n N_noxref_5_M10_noxref_d ) capacitor c=0.00966019f \
 //x=5.55 //y=7.4 //x2=4.185 //y2=5.02
cc_225 ( N_noxref_2_M8_noxref_d N_noxref_5_M10_noxref_d ) capacitor \
 c=0.00561178f //x=3.305 //y=5.02 //x2=4.185 //y2=5.02
cc_226 ( N_noxref_2_c_171_n N_noxref_5_M14_noxref_d ) capacitor c=0.00966019f \
 //x=8.88 //y=7.4 //x2=7.515 //y2=5.02
cc_227 ( N_noxref_2_M12_noxref_d N_noxref_5_M14_noxref_d ) capacitor \
 c=0.00561178f //x=6.635 //y=5.02 //x2=7.515 //y2=5.02
cc_228 ( N_noxref_2_M16_noxref_s N_noxref_5_M14_noxref_d ) capacitor \
 c=5.00921e-19 //x=9.42 //y=5.02 //x2=7.515 //y2=5.02
cc_229 ( N_noxref_2_c_173_p N_noxref_6_c_795_n ) capacitor c=0.0213498f \
 //x=10.36 //y=7.4 //x2=9.505 //y2=4.44
cc_230 ( N_noxref_2_c_210_p N_noxref_6_c_795_n ) capacitor c=0.00304371f \
 //x=8.71 //y=7.4 //x2=9.505 //y2=4.44
cc_231 ( N_noxref_2_c_236_p N_noxref_6_c_795_n ) capacitor c=0.00151604f \
 //x=9.46 //y=7.4 //x2=9.505 //y2=4.44
cc_232 ( N_noxref_2_c_237_p N_noxref_6_c_795_n ) capacitor c=2.37111e-19 \
 //x=10.34 //y=7.4 //x2=9.505 //y2=4.44
cc_233 ( N_noxref_2_c_171_n N_noxref_6_c_795_n ) capacitor c=0.0389665f \
 //x=8.88 //y=7.4 //x2=9.505 //y2=4.44
cc_234 ( N_noxref_2_M16_noxref_s N_noxref_6_c_795_n ) capacitor c=0.00329872f \
 //x=9.42 //y=5.02 //x2=9.505 //y2=4.44
cc_235 ( N_noxref_2_c_173_p N_noxref_6_c_801_n ) capacitor c=0.00150124f \
 //x=10.36 //y=7.4 //x2=6.775 //y2=4.44
cc_236 ( N_noxref_2_c_170_n N_noxref_6_c_801_n ) capacitor c=0.00663859f \
 //x=5.55 //y=7.4 //x2=6.775 //y2=4.44
cc_237 ( N_noxref_2_c_170_n N_noxref_6_c_803_n ) capacitor c=0.0112651f \
 //x=5.55 //y=7.4 //x2=6.66 //y2=4.44
cc_238 ( N_noxref_2_c_171_n N_noxref_6_c_785_n ) capacitor c=0.0189497f \
 //x=8.88 //y=7.4 //x2=9.62 //y2=2.96
cc_239 ( N_noxref_2_c_172_n N_noxref_6_c_785_n ) capacitor c=6.49092e-19 \
 //x=10.36 //y=7.4 //x2=9.62 //y2=2.96
cc_240 ( N_noxref_2_c_172_n N_noxref_6_c_806_n ) capacitor c=0.0179734f \
 //x=10.36 //y=7.4 //x2=9.9 //y2=4.58
cc_241 ( N_noxref_2_c_173_p N_noxref_6_c_807_n ) capacitor c=0.00120205f \
 //x=10.36 //y=7.4 //x2=9.705 //y2=4.58
cc_242 ( N_noxref_2_c_237_p N_noxref_6_c_807_n ) capacitor c=9.4426e-19 \
 //x=10.34 //y=7.4 //x2=9.705 //y2=4.58
cc_243 ( N_noxref_2_c_171_n N_noxref_6_c_807_n ) capacitor c=0.00111372f \
 //x=8.88 //y=7.4 //x2=9.705 //y2=4.58
cc_244 ( N_noxref_2_M16_noxref_s N_noxref_6_c_807_n ) capacitor c=0.00613507f \
 //x=9.42 //y=5.02 //x2=9.705 //y2=4.58
cc_245 ( N_noxref_2_c_250_p N_noxref_6_M12_noxref_g ) capacitor c=0.00673447f \
 //x=6.695 //y=7.4 //x2=6.56 //y2=6.02
cc_246 ( N_noxref_2_c_170_n N_noxref_6_M12_noxref_g ) capacitor c=0.00661226f \
 //x=5.55 //y=7.4 //x2=6.56 //y2=6.02
cc_247 ( N_noxref_2_M12_noxref_d N_noxref_6_M12_noxref_g ) capacitor \
 c=0.0166176f //x=6.635 //y=5.02 //x2=6.56 //y2=6.02
cc_248 ( N_noxref_2_c_210_p N_noxref_6_M13_noxref_g ) capacitor c=0.006727f \
 //x=8.71 //y=7.4 //x2=7 //y2=6.02
cc_249 ( N_noxref_2_M12_noxref_d N_noxref_6_M13_noxref_g ) capacitor \
 c=0.0186652f //x=6.635 //y=5.02 //x2=7 //y2=6.02
cc_250 ( N_noxref_2_c_170_n N_noxref_6_c_816_n ) capacitor c=0.0124704f \
 //x=5.55 //y=7.4 //x2=6.66 //y2=4.7
cc_251 ( N_noxref_2_c_173_p N_noxref_6_M16_noxref_d ) capacitor c=0.00285171f \
 //x=10.36 //y=7.4 //x2=9.84 //y2=5.02
cc_252 ( N_noxref_2_c_237_p N_noxref_6_M16_noxref_d ) capacitor c=0.0141332f \
 //x=10.34 //y=7.4 //x2=9.84 //y2=5.02
cc_253 ( N_noxref_2_c_171_n N_noxref_6_M16_noxref_d ) capacitor c=0.0201812f \
 //x=8.88 //y=7.4 //x2=9.84 //y2=5.02
cc_254 ( N_noxref_2_c_172_n N_noxref_6_M16_noxref_d ) capacitor c=0.00135976f \
 //x=10.36 //y=7.4 //x2=9.84 //y2=5.02
cc_255 ( N_noxref_2_M16_noxref_s N_noxref_6_M16_noxref_d ) capacitor \
 c=0.0832641f //x=9.42 //y=5.02 //x2=9.84 //y2=5.02
cc_256 ( N_noxref_2_M17_noxref_d N_noxref_6_M16_noxref_d ) capacitor \
 c=0.0843065f //x=10.28 //y=5.02 //x2=9.84 //y2=5.02
cc_257 ( N_noxref_2_c_173_p N_noxref_7_c_976_n ) capacitor c=0.03033f \
 //x=10.36 //y=7.4 //x2=10.245 //y2=4.07
cc_258 ( N_noxref_2_c_195_p N_noxref_7_c_976_n ) capacitor c=0.00187833f \
 //x=5.38 //y=7.4 //x2=10.245 //y2=4.07
cc_259 ( N_noxref_2_c_250_p N_noxref_7_c_976_n ) capacitor c=0.00213804f \
 //x=6.695 //y=7.4 //x2=10.245 //y2=4.07
cc_260 ( N_noxref_2_c_237_p N_noxref_7_c_976_n ) capacitor c=9.9102e-19 \
 //x=10.34 //y=7.4 //x2=10.245 //y2=4.07
cc_261 ( N_noxref_2_c_170_n N_noxref_7_c_976_n ) capacitor c=0.0272145f \
 //x=5.55 //y=7.4 //x2=10.245 //y2=4.07
cc_262 ( N_noxref_2_c_171_n N_noxref_7_c_976_n ) capacitor c=0.0140095f \
 //x=8.88 //y=7.4 //x2=10.245 //y2=4.07
cc_263 ( N_noxref_2_c_172_n N_noxref_7_c_976_n ) capacitor c=0.00238507f \
 //x=10.36 //y=7.4 //x2=10.245 //y2=4.07
cc_264 ( N_noxref_2_M17_noxref_d N_noxref_7_c_976_n ) capacitor c=0.00188659f \
 //x=10.28 //y=5.02 //x2=10.245 //y2=4.07
cc_265 ( N_noxref_2_c_173_p N_noxref_7_c_984_n ) capacitor c=0.00164816f \
 //x=10.36 //y=7.4 //x2=4.555 //y2=4.07
cc_266 ( N_noxref_2_c_169_n N_noxref_7_c_985_n ) capacitor c=7.20931e-19 \
 //x=2.22 //y=7.4 //x2=4.44 //y2=4.07
cc_267 ( N_noxref_2_c_170_n N_noxref_7_c_985_n ) capacitor c=0.00211919f \
 //x=5.55 //y=7.4 //x2=4.44 //y2=4.07
cc_268 ( N_noxref_2_c_173_p N_noxref_7_c_951_n ) capacitor c=0.00157744f \
 //x=10.36 //y=7.4 //x2=10.36 //y2=2.085
cc_269 ( N_noxref_2_c_171_n N_noxref_7_c_951_n ) capacitor c=0.00126456f \
 //x=8.88 //y=7.4 //x2=10.36 //y2=2.085
cc_270 ( N_noxref_2_c_172_n N_noxref_7_c_951_n ) capacitor c=0.0266578f \
 //x=10.36 //y=7.4 //x2=10.36 //y2=2.085
cc_271 ( N_noxref_2_M17_noxref_d N_noxref_7_c_951_n ) capacitor c=0.00896093f \
 //x=10.28 //y=5.02 //x2=10.36 //y2=2.085
cc_272 ( N_noxref_2_c_195_p N_noxref_7_M10_noxref_g ) capacitor c=0.00510247f \
 //x=5.38 //y=7.4 //x2=4.11 //y2=6.02
cc_273 ( N_noxref_2_c_195_p N_noxref_7_M11_noxref_g ) capacitor c=0.00510919f \
 //x=5.38 //y=7.4 //x2=4.55 //y2=6.02
cc_274 ( N_noxref_2_c_170_n N_noxref_7_M11_noxref_g ) capacitor c=0.0122307f \
 //x=5.55 //y=7.4 //x2=4.55 //y2=6.02
cc_275 ( N_noxref_2_c_237_p N_noxref_7_M16_noxref_g ) capacitor c=0.00697478f \
 //x=10.34 //y=7.4 //x2=9.765 //y2=6.02
cc_276 ( N_noxref_2_M16_noxref_s N_noxref_7_M16_noxref_g ) capacitor \
 c=0.0528676f //x=9.42 //y=5.02 //x2=9.765 //y2=6.02
cc_277 ( N_noxref_2_c_237_p N_noxref_7_M17_noxref_g ) capacitor c=0.00748034f \
 //x=10.34 //y=7.4 //x2=10.205 //y2=6.02
cc_278 ( N_noxref_2_c_172_n N_noxref_7_M17_noxref_g ) capacitor c=0.0241676f \
 //x=10.36 //y=7.4 //x2=10.205 //y2=6.02
cc_279 ( N_noxref_2_M17_noxref_d N_noxref_7_M17_noxref_g ) capacitor \
 c=0.0528676f //x=10.28 //y=5.02 //x2=10.205 //y2=6.02
cc_280 ( N_noxref_2_c_171_n N_noxref_7_c_999_n ) capacitor c=0.0148045f \
 //x=8.88 //y=7.4 //x2=9.84 //y2=4.79
cc_281 ( N_noxref_2_c_172_n N_noxref_7_c_1000_n ) capacitor c=0.0109438f \
 //x=10.36 //y=7.4 //x2=10.205 //y2=4.865
cc_282 ( N_noxref_2_M17_noxref_d N_noxref_7_c_1000_n ) capacitor c=0.00524527f \
 //x=10.28 //y=5.02 //x2=10.205 //y2=4.865
cc_283 ( N_noxref_2_c_173_p N_noxref_8_c_1119_n ) capacitor c=0.00494742f \
 //x=10.36 //y=7.4 //x2=3.805 //y2=5.205
cc_284 ( N_noxref_2_c_176_p N_noxref_8_c_1119_n ) capacitor c=4.50595e-19 \
 //x=3.365 //y=7.4 //x2=3.805 //y2=5.205
cc_285 ( N_noxref_2_c_195_p N_noxref_8_c_1119_n ) capacitor c=4.35755e-19 \
 //x=5.38 //y=7.4 //x2=3.805 //y2=5.205
cc_286 ( N_noxref_2_c_170_n N_noxref_8_c_1119_n ) capacitor c=0.00289291f \
 //x=5.55 //y=7.4 //x2=3.805 //y2=5.205
cc_287 ( N_noxref_2_M8_noxref_d N_noxref_8_c_1119_n ) capacitor c=0.0127094f \
 //x=3.305 //y=5.02 //x2=3.805 //y2=5.205
cc_288 ( N_noxref_2_c_169_n N_noxref_8_c_1124_n ) capacitor c=0.0628444f \
 //x=2.22 //y=7.4 //x2=3.095 //y2=5.205
cc_289 ( N_noxref_2_M7_noxref_d N_noxref_8_c_1124_n ) capacitor c=0.00269577f \
 //x=1.41 //y=5.02 //x2=3.095 //y2=5.205
cc_290 ( N_noxref_2_c_172_n N_noxref_8_c_1126_n ) capacitor c=0.00351514f \
 //x=10.36 //y=7.4 //x2=4.685 //y2=6.905
cc_291 ( N_noxref_2_c_173_p N_noxref_8_c_1127_n ) capacitor c=0.0260915f \
 //x=10.36 //y=7.4 //x2=3.975 //y2=6.905
cc_292 ( N_noxref_2_c_195_p N_noxref_8_c_1127_n ) capacitor c=0.0593394f \
 //x=5.38 //y=7.4 //x2=3.975 //y2=6.905
cc_293 ( N_noxref_2_c_172_n N_noxref_8_c_1127_n ) capacitor c=0.00115705f \
 //x=10.36 //y=7.4 //x2=3.975 //y2=6.905
cc_294 ( N_noxref_2_c_173_p N_noxref_8_M8_noxref_s ) capacitor c=0.00242367f \
 //x=10.36 //y=7.4 //x2=2.875 //y2=5.02
cc_295 ( N_noxref_2_c_176_p N_noxref_8_M8_noxref_s ) capacitor c=0.0100244f \
 //x=3.365 //y=7.4 //x2=2.875 //y2=5.02
cc_296 ( N_noxref_2_c_172_n N_noxref_8_M8_noxref_s ) capacitor c=7.63704e-19 \
 //x=10.36 //y=7.4 //x2=2.875 //y2=5.02
cc_297 ( N_noxref_2_M8_noxref_d N_noxref_8_M8_noxref_s ) capacitor c=0.061257f \
 //x=3.305 //y=5.02 //x2=2.875 //y2=5.02
cc_298 ( N_noxref_2_c_169_n N_noxref_8_M9_noxref_d ) capacitor c=0.00130916f \
 //x=2.22 //y=7.4 //x2=3.745 //y2=5.02
cc_299 ( N_noxref_2_M8_noxref_d N_noxref_8_M9_noxref_d ) capacitor \
 c=0.0659925f //x=3.305 //y=5.02 //x2=3.745 //y2=5.02
cc_300 ( N_noxref_2_c_170_n N_noxref_8_M11_noxref_d ) capacitor c=0.0520312f \
 //x=5.55 //y=7.4 //x2=4.625 //y2=5.02
cc_301 ( N_noxref_2_M8_noxref_d N_noxref_8_M11_noxref_d ) capacitor \
 c=0.00107819f //x=3.305 //y=5.02 //x2=4.625 //y2=5.02
cc_302 ( N_noxref_2_c_173_p N_noxref_10_c_1211_n ) capacitor c=0.00445614f \
 //x=10.36 //y=7.4 //x2=7.135 //y2=5.205
cc_303 ( N_noxref_2_c_250_p N_noxref_10_c_1211_n ) capacitor c=4.50436e-19 \
 //x=6.695 //y=7.4 //x2=7.135 //y2=5.205
cc_304 ( N_noxref_2_c_210_p N_noxref_10_c_1211_n ) capacitor c=4.50291e-19 \
 //x=8.71 //y=7.4 //x2=7.135 //y2=5.205
cc_305 ( N_noxref_2_c_171_n N_noxref_10_c_1211_n ) capacitor c=0.00289291f \
 //x=8.88 //y=7.4 //x2=7.135 //y2=5.205
cc_306 ( N_noxref_2_M12_noxref_d N_noxref_10_c_1211_n ) capacitor c=0.0123249f \
 //x=6.635 //y=5.02 //x2=7.135 //y2=5.205
cc_307 ( N_noxref_2_c_170_n N_noxref_10_c_1216_n ) capacitor c=0.0628444f \
 //x=5.55 //y=7.4 //x2=6.425 //y2=5.205
cc_308 ( N_noxref_2_c_172_n N_noxref_10_c_1217_n ) capacitor c=0.00351514f \
 //x=10.36 //y=7.4 //x2=8.015 //y2=6.905
cc_309 ( N_noxref_2_c_173_p N_noxref_10_c_1218_n ) capacitor c=0.0164961f \
 //x=10.36 //y=7.4 //x2=7.305 //y2=6.905
cc_310 ( N_noxref_2_c_210_p N_noxref_10_c_1218_n ) capacitor c=0.0608014f \
 //x=8.71 //y=7.4 //x2=7.305 //y2=6.905
cc_311 ( N_noxref_2_c_172_n N_noxref_10_c_1218_n ) capacitor c=0.00115705f \
 //x=10.36 //y=7.4 //x2=7.305 //y2=6.905
cc_312 ( N_noxref_2_c_173_p N_noxref_10_M12_noxref_s ) capacitor c=0.00242367f \
 //x=10.36 //y=7.4 //x2=6.205 //y2=5.02
cc_313 ( N_noxref_2_c_250_p N_noxref_10_M12_noxref_s ) capacitor c=0.0100244f \
 //x=6.695 //y=7.4 //x2=6.205 //y2=5.02
cc_314 ( N_noxref_2_c_172_n N_noxref_10_M12_noxref_s ) capacitor c=7.63704e-19 \
 //x=10.36 //y=7.4 //x2=6.205 //y2=5.02
cc_315 ( N_noxref_2_M12_noxref_d N_noxref_10_M12_noxref_s ) capacitor \
 c=0.061257f //x=6.635 //y=5.02 //x2=6.205 //y2=5.02
cc_316 ( N_noxref_2_c_170_n N_noxref_10_M13_noxref_d ) capacitor c=0.00130916f \
 //x=5.55 //y=7.4 //x2=7.075 //y2=5.02
cc_317 ( N_noxref_2_M12_noxref_d N_noxref_10_M13_noxref_d ) capacitor \
 c=0.0659925f //x=6.635 //y=5.02 //x2=7.075 //y2=5.02
cc_318 ( N_noxref_2_c_171_n N_noxref_10_M15_noxref_d ) capacitor c=0.0520312f \
 //x=8.88 //y=7.4 //x2=7.955 //y2=5.02
cc_319 ( N_noxref_2_M12_noxref_d N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00107819f //x=6.635 //y=5.02 //x2=7.955 //y2=5.02
cc_320 ( N_noxref_2_M16_noxref_s N_noxref_10_M15_noxref_d ) capacitor \
 c=0.00230193f //x=9.42 //y=5.02 //x2=7.955 //y2=5.02
cc_321 ( N_noxref_3_c_326_n N_noxref_4_c_459_n ) capacitor c=0.0423764f \
 //x=3.215 //y=4.07 //x2=7.655 //y2=2.59
cc_322 ( N_noxref_3_c_335_n N_noxref_4_c_459_n ) capacitor c=0.0272395f \
 //x=3.33 //y=2.08 //x2=7.655 //y2=2.59
cc_323 ( N_noxref_3_c_346_n N_noxref_4_c_459_n ) capacitor c=0.0039674f \
 //x=3.135 //y=1.915 //x2=7.655 //y2=2.59
cc_324 ( N_noxref_3_c_326_n N_noxref_4_c_468_n ) capacitor c=0.00521938f \
 //x=3.215 //y=4.07 //x2=1.595 //y2=2.59
cc_325 ( N_noxref_3_c_330_n N_noxref_4_c_468_n ) capacitor c=0.00735597f \
 //x=0.74 //y=2.085 //x2=1.595 //y2=2.59
cc_326 ( N_noxref_3_c_335_n N_noxref_4_c_471_n ) capacitor c=0.0160792f \
 //x=3.33 //y=2.08 //x2=1.395 //y2=2.08
cc_327 ( N_noxref_3_c_389_p N_noxref_4_c_471_n ) capacitor c=0.0023507f \
 //x=1.225 //y=1.41 //x2=1.395 //y2=2.08
cc_328 ( N_noxref_3_c_326_n N_noxref_4_c_510_n ) capacitor c=0.0023373f \
 //x=3.215 //y=4.07 //x2=1.195 //y2=2.08
cc_329 ( N_noxref_3_c_352_n N_noxref_4_c_510_n ) capacitor c=0.0167852f \
 //x=0.74 //y=2.085 //x2=1.195 //y2=2.08
cc_330 ( N_noxref_3_c_379_n N_noxref_4_c_486_n ) capacitor c=0.0099173f \
 //x=1.26 //y=4.79 //x2=1.395 //y2=4.58
cc_331 ( N_noxref_3_c_326_n N_noxref_4_c_489_n ) capacitor c=0.0123666f \
 //x=3.215 //y=4.07 //x2=1.2 //y2=4.58
cc_332 ( N_noxref_3_c_330_n N_noxref_4_c_489_n ) capacitor c=0.0250789f \
 //x=0.74 //y=2.085 //x2=1.2 //y2=4.58
cc_333 ( N_noxref_3_c_380_n N_noxref_4_c_489_n ) capacitor c=0.00962086f \
 //x=0.97 //y=4.79 //x2=1.2 //y2=4.58
cc_334 ( N_noxref_3_c_326_n N_noxref_4_c_474_n ) capacitor c=0.0269755f \
 //x=3.215 //y=4.07 //x2=1.48 //y2=2.59
cc_335 ( N_noxref_3_c_328_n N_noxref_4_c_474_n ) capacitor c=0.00101501f \
 //x=0.855 //y=4.07 //x2=1.48 //y2=2.59
cc_336 ( N_noxref_3_c_330_n N_noxref_4_c_474_n ) capacitor c=0.068675f \
 //x=0.74 //y=2.085 //x2=1.48 //y2=2.59
cc_337 ( N_noxref_3_c_352_n N_noxref_4_c_474_n ) capacitor c=8.49451e-19 \
 //x=0.74 //y=2.085 //x2=1.48 //y2=2.59
cc_338 ( N_noxref_3_c_330_n N_noxref_4_M0_noxref_d ) capacitor c=0.0175773f \
 //x=0.74 //y=2.085 //x2=0.925 //y2=0.91
cc_339 ( N_noxref_3_c_336_n N_noxref_4_M0_noxref_d ) capacitor c=0.00218556f \
 //x=0.85 //y=0.91 //x2=0.925 //y2=0.91
cc_340 ( N_noxref_3_c_402_p N_noxref_4_M0_noxref_d ) capacitor c=0.00347355f \
 //x=0.85 //y=1.255 //x2=0.925 //y2=0.91
cc_341 ( N_noxref_3_c_403_p N_noxref_4_M0_noxref_d ) capacitor c=0.00742431f \
 //x=0.85 //y=1.565 //x2=0.925 //y2=0.91
cc_342 ( N_noxref_3_c_338_n N_noxref_4_M0_noxref_d ) capacitor c=0.00957707f \
 //x=0.85 //y=1.92 //x2=0.925 //y2=0.91
cc_343 ( N_noxref_3_c_339_n N_noxref_4_M0_noxref_d ) capacitor c=0.00220879f \
 //x=1.225 //y=0.755 //x2=0.925 //y2=0.91
cc_344 ( N_noxref_3_c_389_p N_noxref_4_M0_noxref_d ) capacitor c=0.0138447f \
 //x=1.225 //y=1.41 //x2=0.925 //y2=0.91
cc_345 ( N_noxref_3_c_340_n N_noxref_4_M0_noxref_d ) capacitor c=0.00218624f \
 //x=1.38 //y=0.91 //x2=0.925 //y2=0.91
cc_346 ( N_noxref_3_c_342_n N_noxref_4_M0_noxref_d ) capacitor c=0.00601286f \
 //x=1.38 //y=1.255 //x2=0.925 //y2=0.91
cc_347 ( N_noxref_3_M6_noxref_g N_noxref_4_M6_noxref_d ) capacitor \
 c=0.0219309f //x=0.895 //y=6.02 //x2=0.97 //y2=5.02
cc_348 ( N_noxref_3_M7_noxref_g N_noxref_4_M6_noxref_d ) capacitor c=0.021902f \
 //x=1.335 //y=6.02 //x2=0.97 //y2=5.02
cc_349 ( N_noxref_3_c_379_n N_noxref_4_M6_noxref_d ) capacitor c=0.0146106f \
 //x=1.26 //y=4.79 //x2=0.97 //y2=5.02
cc_350 ( N_noxref_3_c_380_n N_noxref_4_M6_noxref_d ) capacitor c=0.00307344f \
 //x=0.97 //y=4.79 //x2=0.97 //y2=5.02
cc_351 ( N_noxref_3_c_335_n N_noxref_5_c_655_n ) capacitor c=0.00382062f \
 //x=3.33 //y=2.08 //x2=4.925 //y2=3.7
cc_352 ( N_noxref_3_c_335_n N_noxref_5_c_629_n ) capacitor c=0.015408f \
 //x=3.33 //y=2.08 //x2=4.81 //y2=3.7
cc_353 ( N_noxref_3_c_335_n N_noxref_6_c_823_n ) capacitor c=0.00526349f \
 //x=3.33 //y=2.08 //x2=4.555 //y2=2.96
cc_354 ( N_noxref_3_c_335_n N_noxref_6_c_783_n ) capacitor c=0.0198069f \
 //x=3.33 //y=2.08 //x2=4.44 //y2=2.08
cc_355 ( N_noxref_3_c_346_n N_noxref_6_c_783_n ) capacitor c=0.00220284f \
 //x=3.135 //y=1.915 //x2=4.44 //y2=2.08
cc_356 ( N_noxref_3_c_343_n N_noxref_6_c_826_n ) capacitor c=4.86506e-19 \
 //x=3.135 //y=0.865 //x2=4.105 //y2=0.905
cc_357 ( N_noxref_3_c_345_n N_noxref_6_c_826_n ) capacitor c=0.00152104f \
 //x=3.135 //y=1.21 //x2=4.105 //y2=0.905
cc_358 ( N_noxref_3_c_349_n N_noxref_6_c_826_n ) capacitor c=0.0157772f \
 //x=3.665 //y=0.865 //x2=4.105 //y2=0.905
cc_359 ( N_noxref_3_c_421_p N_noxref_6_c_829_n ) capacitor c=0.00109982f \
 //x=3.135 //y=1.52 //x2=4.105 //y2=1.25
cc_360 ( N_noxref_3_c_351_n N_noxref_6_c_829_n ) capacitor c=0.0117362f \
 //x=3.665 //y=1.21 //x2=4.105 //y2=1.25
cc_361 ( N_noxref_3_c_421_p N_noxref_6_c_831_n ) capacitor c=9.57794e-19 \
 //x=3.135 //y=1.52 //x2=4.105 //y2=1.56
cc_362 ( N_noxref_3_c_346_n N_noxref_6_c_831_n ) capacitor c=0.00662747f \
 //x=3.135 //y=1.915 //x2=4.105 //y2=1.56
cc_363 ( N_noxref_3_c_351_n N_noxref_6_c_831_n ) capacitor c=0.00862358f \
 //x=3.665 //y=1.21 //x2=4.105 //y2=1.56
cc_364 ( N_noxref_3_c_335_n N_noxref_6_c_834_n ) capacitor c=0.00251238f \
 //x=3.33 //y=2.08 //x2=4.105 //y2=1.915
cc_365 ( N_noxref_3_c_346_n N_noxref_6_c_834_n ) capacitor c=0.012079f \
 //x=3.135 //y=1.915 //x2=4.105 //y2=1.915
cc_366 ( N_noxref_3_c_349_n N_noxref_6_c_836_n ) capacitor c=0.00124821f \
 //x=3.665 //y=0.865 //x2=4.635 //y2=0.905
cc_367 ( N_noxref_3_c_351_n N_noxref_6_c_837_n ) capacitor c=0.00200715f \
 //x=3.665 //y=1.21 //x2=4.635 //y2=1.25
cc_368 ( N_noxref_3_c_326_n N_noxref_7_c_984_n ) capacitor c=0.0159617f \
 //x=3.215 //y=4.07 //x2=4.555 //y2=4.07
cc_369 ( N_noxref_3_c_335_n N_noxref_7_c_984_n ) capacitor c=0.00187343f \
 //x=3.33 //y=2.08 //x2=4.555 //y2=4.07
cc_370 ( N_noxref_3_c_326_n N_noxref_7_c_985_n ) capacitor c=0.00186775f \
 //x=3.215 //y=4.07 //x2=4.44 //y2=4.07
cc_371 ( N_noxref_3_c_335_n N_noxref_7_c_985_n ) capacitor c=0.0166316f \
 //x=3.33 //y=2.08 //x2=4.44 //y2=4.07
cc_372 ( N_noxref_3_c_382_n N_noxref_7_c_985_n ) capacitor c=0.0022916f \
 //x=3.33 //y=4.7 //x2=4.44 //y2=4.07
cc_373 ( N_noxref_3_c_335_n N_noxref_7_c_950_n ) capacitor c=2.12957e-19 \
 //x=3.33 //y=2.08 //x2=6.66 //y2=2.08
cc_374 ( N_noxref_3_M8_noxref_g N_noxref_7_M10_noxref_g ) capacitor \
 c=0.0100243f //x=3.23 //y=6.02 //x2=4.11 //y2=6.02
cc_375 ( N_noxref_3_M9_noxref_g N_noxref_7_M10_noxref_g ) capacitor \
 c=0.0610135f //x=3.67 //y=6.02 //x2=4.11 //y2=6.02
cc_376 ( N_noxref_3_M9_noxref_g N_noxref_7_M11_noxref_g ) capacitor \
 c=0.0094155f //x=3.67 //y=6.02 //x2=4.55 //y2=6.02
cc_377 ( N_noxref_3_c_335_n N_noxref_7_c_1011_n ) capacitor c=0.00227843f \
 //x=3.33 //y=2.08 //x2=4.44 //y2=4.7
cc_378 ( N_noxref_3_c_382_n N_noxref_7_c_1011_n ) capacitor c=0.066749f \
 //x=3.33 //y=4.7 //x2=4.44 //y2=4.7
cc_379 ( N_noxref_3_c_326_n N_noxref_8_c_1119_n ) capacitor c=0.00305144f \
 //x=3.215 //y=4.07 //x2=3.805 //y2=5.205
cc_380 ( N_noxref_3_c_335_n N_noxref_8_c_1119_n ) capacitor c=0.0120072f \
 //x=3.33 //y=2.08 //x2=3.805 //y2=5.205
cc_381 ( N_noxref_3_M8_noxref_g N_noxref_8_c_1119_n ) capacitor c=0.019052f \
 //x=3.23 //y=6.02 //x2=3.805 //y2=5.205
cc_382 ( N_noxref_3_M9_noxref_g N_noxref_8_c_1119_n ) capacitor c=0.0198429f \
 //x=3.67 //y=6.02 //x2=3.805 //y2=5.205
cc_383 ( N_noxref_3_c_382_n N_noxref_8_c_1119_n ) capacitor c=0.00525548f \
 //x=3.33 //y=4.7 //x2=3.805 //y2=5.205
cc_384 ( N_noxref_3_c_326_n N_noxref_8_c_1124_n ) capacitor c=0.00704018f \
 //x=3.215 //y=4.07 //x2=3.095 //y2=5.205
cc_385 ( N_noxref_3_M8_noxref_g N_noxref_8_M8_noxref_s ) capacitor \
 c=0.0441361f //x=3.23 //y=6.02 //x2=2.875 //y2=5.02
cc_386 ( N_noxref_3_M9_noxref_g N_noxref_8_M9_noxref_d ) capacitor \
 c=0.0170604f //x=3.67 //y=6.02 //x2=3.745 //y2=5.02
cc_387 ( N_noxref_3_c_346_n N_noxref_9_c_1159_n ) capacitor c=0.0034165f \
 //x=3.135 //y=1.915 //x2=2.915 //y2=1.495
cc_388 ( N_noxref_3_c_335_n N_noxref_9_c_1160_n ) capacitor c=0.011424f \
 //x=3.33 //y=2.08 //x2=3.8 //y2=1.58
cc_389 ( N_noxref_3_c_421_p N_noxref_9_c_1160_n ) capacitor c=0.00703567f \
 //x=3.135 //y=1.52 //x2=3.8 //y2=1.58
cc_390 ( N_noxref_3_c_346_n N_noxref_9_c_1160_n ) capacitor c=0.018562f \
 //x=3.135 //y=1.915 //x2=3.8 //y2=1.58
cc_391 ( N_noxref_3_c_348_n N_noxref_9_c_1160_n ) capacitor c=0.00780629f \
 //x=3.51 //y=1.365 //x2=3.8 //y2=1.58
cc_392 ( N_noxref_3_c_351_n N_noxref_9_c_1160_n ) capacitor c=0.00339872f \
 //x=3.665 //y=1.21 //x2=3.8 //y2=1.58
cc_393 ( N_noxref_3_c_346_n N_noxref_9_c_1168_n ) capacitor c=6.71402e-19 \
 //x=3.135 //y=1.915 //x2=3.885 //y2=1.495
cc_394 ( N_noxref_3_c_343_n N_noxref_9_M1_noxref_s ) capacitor c=0.0326577f \
 //x=3.135 //y=0.865 //x2=2.78 //y2=0.365
cc_395 ( N_noxref_3_c_421_p N_noxref_9_M1_noxref_s ) capacitor c=3.48408e-19 \
 //x=3.135 //y=1.52 //x2=2.78 //y2=0.365
cc_396 ( N_noxref_3_c_349_n N_noxref_9_M1_noxref_s ) capacitor c=0.0120759f \
 //x=3.665 //y=0.865 //x2=2.78 //y2=0.365
cc_397 ( N_noxref_4_c_459_n N_noxref_5_c_657_n ) capacitor c=0.00619192f \
 //x=7.655 //y=2.59 //x2=8.025 //y2=3.7
cc_398 ( N_noxref_4_c_477_n N_noxref_5_c_657_n ) capacitor c=0.0182358f \
 //x=7.77 //y=2.08 //x2=8.025 //y2=3.7
cc_399 ( N_noxref_4_c_459_n N_noxref_5_c_655_n ) capacitor c=6.30522e-19 \
 //x=7.655 //y=2.59 //x2=4.925 //y2=3.7
cc_400 ( N_noxref_4_c_477_n N_noxref_5_c_655_n ) capacitor c=2.02744e-19 \
 //x=7.77 //y=2.08 //x2=4.925 //y2=3.7
cc_401 ( N_noxref_4_c_459_n N_noxref_5_c_642_n ) capacitor c=4.14375e-19 \
 //x=7.655 //y=2.59 //x2=4.415 //y2=5.205
cc_402 ( N_noxref_4_c_459_n N_noxref_5_c_628_n ) capacitor c=0.00450697f \
 //x=7.655 //y=2.59 //x2=4.725 //y2=1.65
cc_403 ( N_noxref_4_c_459_n N_noxref_5_c_663_n ) capacitor c=0.00178688f \
 //x=7.655 //y=2.59 //x2=4.455 //y2=1.65
cc_404 ( N_noxref_4_c_459_n N_noxref_5_c_629_n ) capacitor c=0.0188708f \
 //x=7.655 //y=2.59 //x2=4.81 //y2=3.7
cc_405 ( N_noxref_4_c_474_n N_noxref_5_c_629_n ) capacitor c=2.79968e-19 \
 //x=1.48 //y=2.59 //x2=4.81 //y2=3.7
cc_406 ( N_noxref_4_c_477_n N_noxref_5_c_629_n ) capacitor c=0.00277451f \
 //x=7.77 //y=2.08 //x2=4.81 //y2=3.7
cc_407 ( N_noxref_4_M15_noxref_g N_noxref_5_c_645_n ) capacitor c=0.0180846f \
 //x=7.88 //y=6.02 //x2=8.055 //y2=5.205
cc_408 ( N_noxref_4_c_544_p N_noxref_5_c_645_n ) capacitor c=0.00161455f \
 //x=7.77 //y=4.7 //x2=8.055 //y2=5.205
cc_409 ( N_noxref_4_c_477_n N_noxref_5_c_647_n ) capacitor c=0.012972f \
 //x=7.77 //y=2.08 //x2=7.745 //y2=5.205
cc_410 ( N_noxref_4_M14_noxref_g N_noxref_5_c_647_n ) capacitor c=0.0132788f \
 //x=7.44 //y=6.02 //x2=7.745 //y2=5.205
cc_411 ( N_noxref_4_c_544_p N_noxref_5_c_647_n ) capacitor c=0.00554627f \
 //x=7.77 //y=4.7 //x2=7.745 //y2=5.205
cc_412 ( N_noxref_4_c_459_n N_noxref_5_c_630_n ) capacitor c=0.00139832f \
 //x=7.655 //y=2.59 //x2=8.055 //y2=1.65
cc_413 ( N_noxref_4_c_549_p N_noxref_5_c_630_n ) capacitor c=0.00363601f \
 //x=7.435 //y=1.915 //x2=8.055 //y2=1.65
cc_414 ( N_noxref_4_c_550_p N_noxref_5_c_630_n ) capacitor c=0.00196666f \
 //x=7.81 //y=1.405 //x2=8.055 //y2=1.65
cc_415 ( N_noxref_4_c_551_p N_noxref_5_c_630_n ) capacitor c=0.00423452f \
 //x=7.965 //y=1.25 //x2=8.055 //y2=1.65
cc_416 ( N_noxref_4_c_459_n N_noxref_5_c_676_n ) capacitor c=0.00184518f \
 //x=7.655 //y=2.59 //x2=7.785 //y2=1.65
cc_417 ( N_noxref_4_c_477_n N_noxref_5_c_676_n ) capacitor c=0.0171043f \
 //x=7.77 //y=2.08 //x2=7.785 //y2=1.65
cc_418 ( N_noxref_4_c_549_p N_noxref_5_c_676_n ) capacitor c=0.00637984f \
 //x=7.435 //y=1.915 //x2=7.785 //y2=1.65
cc_419 ( N_noxref_4_c_459_n N_noxref_5_c_632_n ) capacitor c=0.0100753f \
 //x=7.655 //y=2.59 //x2=8.14 //y2=3.7
cc_420 ( N_noxref_4_c_477_n N_noxref_5_c_632_n ) capacitor c=0.187581f \
 //x=7.77 //y=2.08 //x2=8.14 //y2=3.7
cc_421 ( N_noxref_4_c_549_p N_noxref_5_c_632_n ) capacitor c=0.0185661f \
 //x=7.435 //y=1.915 //x2=8.14 //y2=3.7
cc_422 ( N_noxref_4_c_544_p N_noxref_5_c_632_n ) capacitor c=0.0232466f \
 //x=7.77 //y=4.7 //x2=8.14 //y2=3.7
cc_423 ( N_noxref_4_c_559_p N_noxref_5_M4_noxref_d ) capacitor c=0.00217566f \
 //x=7.435 //y=0.905 //x2=7.51 //y2=0.905
cc_424 ( N_noxref_4_c_560_p N_noxref_5_M4_noxref_d ) capacitor c=0.0034598f \
 //x=7.435 //y=1.25 //x2=7.51 //y2=0.905
cc_425 ( N_noxref_4_c_561_p N_noxref_5_M4_noxref_d ) capacitor c=0.00522042f \
 //x=7.435 //y=1.56 //x2=7.51 //y2=0.905
cc_426 ( N_noxref_4_c_549_p N_noxref_5_M4_noxref_d ) capacitor c=0.00643086f \
 //x=7.435 //y=1.915 //x2=7.51 //y2=0.905
cc_427 ( N_noxref_4_c_563_p N_noxref_5_M4_noxref_d ) capacitor c=0.00241053f \
 //x=7.81 //y=0.75 //x2=7.51 //y2=0.905
cc_428 ( N_noxref_4_c_550_p N_noxref_5_M4_noxref_d ) capacitor c=0.0124466f \
 //x=7.81 //y=1.405 //x2=7.51 //y2=0.905
cc_429 ( N_noxref_4_c_565_p N_noxref_5_M4_noxref_d ) capacitor c=0.00132245f \
 //x=7.965 //y=0.905 //x2=7.51 //y2=0.905
cc_430 ( N_noxref_4_c_551_p N_noxref_5_M4_noxref_d ) capacitor c=0.00566463f \
 //x=7.965 //y=1.25 //x2=7.51 //y2=0.905
cc_431 ( N_noxref_4_M15_noxref_g N_noxref_5_M14_noxref_d ) capacitor \
 c=0.0136385f //x=7.88 //y=6.02 //x2=7.515 //y2=5.02
cc_432 ( N_noxref_4_c_459_n N_noxref_6_c_777_n ) capacitor c=0.300248f \
 //x=7.655 //y=2.59 //x2=9.505 //y2=2.96
cc_433 ( N_noxref_4_c_477_n N_noxref_6_c_777_n ) capacitor c=0.017634f \
 //x=7.77 //y=2.08 //x2=9.505 //y2=2.96
cc_434 ( N_noxref_4_c_459_n N_noxref_6_c_823_n ) capacitor c=0.0290334f \
 //x=7.655 //y=2.59 //x2=4.555 //y2=2.96
cc_435 ( N_noxref_4_c_477_n N_noxref_6_c_795_n ) capacitor c=0.01781f //x=7.77 \
 //y=2.08 //x2=9.505 //y2=4.44
cc_436 ( N_noxref_4_c_544_p N_noxref_6_c_795_n ) capacitor c=0.0105048f \
 //x=7.77 //y=4.7 //x2=9.505 //y2=4.44
cc_437 ( N_noxref_4_c_477_n N_noxref_6_c_801_n ) capacitor c=8.88124e-19 \
 //x=7.77 //y=2.08 //x2=6.775 //y2=4.44
cc_438 ( N_noxref_4_c_459_n N_noxref_6_c_783_n ) capacitor c=0.0210269f \
 //x=7.655 //y=2.59 //x2=4.44 //y2=2.08
cc_439 ( N_noxref_4_c_474_n N_noxref_6_c_783_n ) capacitor c=2.14844e-19 \
 //x=1.48 //y=2.59 //x2=4.44 //y2=2.08
cc_440 ( N_noxref_4_c_477_n N_noxref_6_c_803_n ) capacitor c=0.00835507f \
 //x=7.77 //y=2.08 //x2=6.66 //y2=4.44
cc_441 ( N_noxref_4_c_544_p N_noxref_6_c_803_n ) capacitor c=0.00226398f \
 //x=7.77 //y=4.7 //x2=6.66 //y2=4.44
cc_442 ( N_noxref_4_c_477_n N_noxref_6_c_785_n ) capacitor c=0.00205806f \
 //x=7.77 //y=2.08 //x2=9.62 //y2=2.96
cc_443 ( N_noxref_4_M14_noxref_g N_noxref_6_M12_noxref_g ) capacitor \
 c=0.0100243f //x=7.44 //y=6.02 //x2=6.56 //y2=6.02
cc_444 ( N_noxref_4_M14_noxref_g N_noxref_6_M13_noxref_g ) capacitor \
 c=0.0610135f //x=7.44 //y=6.02 //x2=7 //y2=6.02
cc_445 ( N_noxref_4_M15_noxref_g N_noxref_6_M13_noxref_g ) capacitor \
 c=0.0094155f //x=7.88 //y=6.02 //x2=7 //y2=6.02
cc_446 ( N_noxref_4_c_459_n N_noxref_6_c_834_n ) capacitor c=0.0077361f \
 //x=7.655 //y=2.59 //x2=4.105 //y2=1.915
cc_447 ( N_noxref_4_c_477_n N_noxref_6_c_816_n ) capacitor c=0.0022916f \
 //x=7.77 //y=2.08 //x2=6.66 //y2=4.7
cc_448 ( N_noxref_4_c_544_p N_noxref_6_c_816_n ) capacitor c=0.066749f \
 //x=7.77 //y=4.7 //x2=6.66 //y2=4.7
cc_449 ( N_noxref_4_c_459_n N_noxref_7_c_976_n ) capacitor c=7.67053e-19 \
 //x=7.655 //y=2.59 //x2=10.245 //y2=4.07
cc_450 ( N_noxref_4_c_477_n N_noxref_7_c_976_n ) capacitor c=0.0166527f \
 //x=7.77 //y=2.08 //x2=10.245 //y2=4.07
cc_451 ( N_noxref_4_c_459_n N_noxref_7_c_984_n ) capacitor c=6.56379e-19 \
 //x=7.655 //y=2.59 //x2=4.555 //y2=4.07
cc_452 ( N_noxref_4_c_459_n N_noxref_7_c_947_n ) capacitor c=0.00949333f \
 //x=7.655 //y=2.59 //x2=10.245 //y2=3.33
cc_453 ( N_noxref_4_c_477_n N_noxref_7_c_947_n ) capacitor c=0.0158196f \
 //x=7.77 //y=2.08 //x2=10.245 //y2=3.33
cc_454 ( N_noxref_4_c_459_n N_noxref_7_c_1018_n ) capacitor c=9.79061e-19 \
 //x=7.655 //y=2.59 //x2=6.775 //y2=3.33
cc_455 ( N_noxref_4_c_477_n N_noxref_7_c_1018_n ) capacitor c=8.17135e-19 \
 //x=7.77 //y=2.08 //x2=6.775 //y2=3.33
cc_456 ( N_noxref_4_c_459_n N_noxref_7_c_950_n ) capacitor c=0.0236477f \
 //x=7.655 //y=2.59 //x2=6.66 //y2=2.08
cc_457 ( N_noxref_4_c_477_n N_noxref_7_c_950_n ) capacitor c=0.0239362f \
 //x=7.77 //y=2.08 //x2=6.66 //y2=2.08
cc_458 ( N_noxref_4_c_549_p N_noxref_7_c_950_n ) capacitor c=0.00251238f \
 //x=7.435 //y=1.915 //x2=6.66 //y2=2.08
cc_459 ( N_noxref_4_c_559_p N_noxref_7_c_956_n ) capacitor c=4.86506e-19 \
 //x=7.435 //y=0.905 //x2=6.465 //y2=0.865
cc_460 ( N_noxref_4_c_559_p N_noxref_7_c_958_n ) capacitor c=0.00152104f \
 //x=7.435 //y=0.905 //x2=6.465 //y2=1.21
cc_461 ( N_noxref_4_c_560_p N_noxref_7_c_959_n ) capacitor c=0.00109982f \
 //x=7.435 //y=1.25 //x2=6.465 //y2=1.52
cc_462 ( N_noxref_4_c_561_p N_noxref_7_c_959_n ) capacitor c=9.57794e-19 \
 //x=7.435 //y=1.56 //x2=6.465 //y2=1.52
cc_463 ( N_noxref_4_c_459_n N_noxref_7_c_960_n ) capacitor c=0.0052136f \
 //x=7.655 //y=2.59 //x2=6.465 //y2=1.915
cc_464 ( N_noxref_4_c_477_n N_noxref_7_c_960_n ) capacitor c=0.00220284f \
 //x=7.77 //y=2.08 //x2=6.465 //y2=1.915
cc_465 ( N_noxref_4_c_561_p N_noxref_7_c_960_n ) capacitor c=0.00662747f \
 //x=7.435 //y=1.56 //x2=6.465 //y2=1.915
cc_466 ( N_noxref_4_c_549_p N_noxref_7_c_960_n ) capacitor c=0.012079f \
 //x=7.435 //y=1.915 //x2=6.465 //y2=1.915
cc_467 ( N_noxref_4_c_559_p N_noxref_7_c_963_n ) capacitor c=0.0157772f \
 //x=7.435 //y=0.905 //x2=6.995 //y2=0.865
cc_468 ( N_noxref_4_c_565_p N_noxref_7_c_963_n ) capacitor c=0.00124821f \
 //x=7.965 //y=0.905 //x2=6.995 //y2=0.865
cc_469 ( N_noxref_4_c_560_p N_noxref_7_c_965_n ) capacitor c=0.0117362f \
 //x=7.435 //y=1.25 //x2=6.995 //y2=1.21
cc_470 ( N_noxref_4_c_561_p N_noxref_7_c_965_n ) capacitor c=0.00862358f \
 //x=7.435 //y=1.56 //x2=6.995 //y2=1.21
cc_471 ( N_noxref_4_c_551_p N_noxref_7_c_965_n ) capacitor c=0.00200715f \
 //x=7.965 //y=1.25 //x2=6.995 //y2=1.21
cc_472 ( N_noxref_4_c_459_n N_noxref_8_c_1119_n ) capacitor c=0.00649136f \
 //x=7.655 //y=2.59 //x2=3.805 //y2=5.205
cc_473 ( N_noxref_4_c_459_n N_noxref_9_c_1159_n ) capacitor c=0.00444239f \
 //x=7.655 //y=2.59 //x2=2.915 //y2=1.495
cc_474 ( N_noxref_4_c_459_n N_noxref_9_c_1160_n ) capacitor c=0.0161747f \
 //x=7.655 //y=2.59 //x2=3.8 //y2=1.58
cc_475 ( N_noxref_4_c_459_n N_noxref_9_c_1168_n ) capacitor c=0.00432969f \
 //x=7.655 //y=2.59 //x2=3.885 //y2=1.495
cc_476 ( N_noxref_4_c_459_n N_noxref_9_c_1169_n ) capacitor c=0.00191775f \
 //x=7.655 //y=2.59 //x2=4.77 //y2=0.53
cc_477 ( N_noxref_4_c_459_n N_noxref_9_M1_noxref_s ) capacitor c=8.24206e-19 \
 //x=7.655 //y=2.59 //x2=2.78 //y2=0.365
cc_478 ( N_noxref_4_M14_noxref_g N_noxref_10_c_1211_n ) capacitor c=0.0170604f \
 //x=7.44 //y=6.02 //x2=7.135 //y2=5.205
cc_479 ( N_noxref_4_M14_noxref_g N_noxref_10_c_1217_n ) capacitor c=0.0144401f \
 //x=7.44 //y=6.02 //x2=8.015 //y2=6.905
cc_480 ( N_noxref_4_M15_noxref_g N_noxref_10_c_1217_n ) capacitor c=0.0163317f \
 //x=7.88 //y=6.02 //x2=8.015 //y2=6.905
cc_481 ( N_noxref_4_M15_noxref_g N_noxref_10_M15_noxref_d ) capacitor \
 c=0.0351101f //x=7.88 //y=6.02 //x2=7.955 //y2=5.02
cc_482 ( N_noxref_4_c_459_n N_noxref_11_c_1278_n ) capacitor c=0.00444239f \
 //x=7.655 //y=2.59 //x2=6.245 //y2=1.495
cc_483 ( N_noxref_4_c_459_n N_noxref_11_c_1254_n ) capacitor c=0.0162171f \
 //x=7.655 //y=2.59 //x2=7.13 //y2=1.58
cc_484 ( N_noxref_4_c_459_n N_noxref_11_c_1262_n ) capacitor c=0.00444239f \
 //x=7.655 //y=2.59 //x2=7.215 //y2=1.495
cc_485 ( N_noxref_4_c_561_p N_noxref_11_c_1262_n ) capacitor c=0.00628626f \
 //x=7.435 //y=1.56 //x2=7.215 //y2=1.495
cc_486 ( N_noxref_4_c_459_n N_noxref_11_c_1263_n ) capacitor c=0.00229834f \
 //x=7.655 //y=2.59 //x2=8.1 //y2=0.53
cc_487 ( N_noxref_4_c_559_p N_noxref_11_c_1263_n ) capacitor c=0.0197889f \
 //x=7.435 //y=0.905 //x2=8.1 //y2=0.53
cc_488 ( N_noxref_4_c_565_p N_noxref_11_c_1263_n ) capacitor c=0.00655813f \
 //x=7.965 //y=0.905 //x2=8.1 //y2=0.53
cc_489 ( N_noxref_4_c_559_p N_noxref_11_M3_noxref_s ) capacitor c=0.00628626f \
 //x=7.435 //y=0.905 //x2=6.11 //y2=0.365
cc_490 ( N_noxref_4_c_565_p N_noxref_11_M3_noxref_s ) capacitor c=0.0143002f \
 //x=7.965 //y=0.905 //x2=6.11 //y2=0.365
cc_491 ( N_noxref_4_c_551_p N_noxref_11_M3_noxref_s ) capacitor c=0.00290153f \
 //x=7.965 //y=1.25 //x2=6.11 //y2=0.365
cc_492 ( N_noxref_5_c_657_n N_noxref_6_c_777_n ) capacitor c=0.085017f \
 //x=8.025 //y=3.7 //x2=9.505 //y2=2.96
cc_493 ( N_noxref_5_c_655_n N_noxref_6_c_777_n ) capacitor c=0.0133599f \
 //x=4.925 //y=3.7 //x2=9.505 //y2=2.96
cc_494 ( N_noxref_5_c_629_n N_noxref_6_c_777_n ) capacitor c=0.0192028f \
 //x=4.81 //y=3.7 //x2=9.505 //y2=2.96
cc_495 ( N_noxref_5_c_630_n N_noxref_6_c_777_n ) capacitor c=0.00228574f \
 //x=8.055 //y=1.65 //x2=9.505 //y2=2.96
cc_496 ( N_noxref_5_c_632_n N_noxref_6_c_777_n ) capacitor c=0.022345f \
 //x=8.14 //y=3.7 //x2=9.505 //y2=2.96
cc_497 ( N_noxref_5_c_629_n N_noxref_6_c_823_n ) capacitor c=0.00244604f \
 //x=4.81 //y=3.7 //x2=4.555 //y2=2.96
cc_498 ( N_noxref_5_c_657_n N_noxref_6_c_795_n ) capacitor c=0.0110295f \
 //x=8.025 //y=3.7 //x2=9.505 //y2=4.44
cc_499 ( N_noxref_5_c_645_n N_noxref_6_c_795_n ) capacitor c=0.00665427f \
 //x=8.055 //y=5.205 //x2=9.505 //y2=4.44
cc_500 ( N_noxref_5_c_647_n N_noxref_6_c_795_n ) capacitor c=0.00351988f \
 //x=7.745 //y=5.205 //x2=9.505 //y2=4.44
cc_501 ( N_noxref_5_c_632_n N_noxref_6_c_795_n ) capacitor c=0.0186188f \
 //x=8.14 //y=3.7 //x2=9.505 //y2=4.44
cc_502 ( N_noxref_5_c_657_n N_noxref_6_c_801_n ) capacitor c=0.00181513f \
 //x=8.025 //y=3.7 //x2=6.775 //y2=4.44
cc_503 ( N_noxref_5_c_663_n N_noxref_6_c_783_n ) capacitor c=0.0163956f \
 //x=4.455 //y=1.65 //x2=4.44 //y2=2.08
cc_504 ( N_noxref_5_c_629_n N_noxref_6_c_783_n ) capacitor c=0.0793595f \
 //x=4.81 //y=3.7 //x2=4.44 //y2=2.08
cc_505 ( N_noxref_5_c_629_n N_noxref_6_c_803_n ) capacitor c=7.44407e-19 \
 //x=4.81 //y=3.7 //x2=6.66 //y2=4.44
cc_506 ( N_noxref_5_c_632_n N_noxref_6_c_803_n ) capacitor c=0.00138227f \
 //x=8.14 //y=3.7 //x2=6.66 //y2=4.44
cc_507 ( N_noxref_5_c_657_n N_noxref_6_c_785_n ) capacitor c=0.00382062f \
 //x=8.025 //y=3.7 //x2=9.62 //y2=2.96
cc_508 ( N_noxref_5_c_632_n N_noxref_6_c_787_n ) capacitor c=0.0154636f \
 //x=8.14 //y=3.7 //x2=9.705 //y2=2.08
cc_509 ( N_noxref_5_M2_noxref_d N_noxref_6_c_826_n ) capacitor c=0.00217566f \
 //x=4.18 //y=0.905 //x2=4.105 //y2=0.905
cc_510 ( N_noxref_5_M2_noxref_d N_noxref_6_c_829_n ) capacitor c=0.0034598f \
 //x=4.18 //y=0.905 //x2=4.105 //y2=1.25
cc_511 ( N_noxref_5_M2_noxref_d N_noxref_6_c_831_n ) capacitor c=0.00522042f \
 //x=4.18 //y=0.905 //x2=4.105 //y2=1.56
cc_512 ( N_noxref_5_c_628_n N_noxref_6_c_834_n ) capacitor c=0.00363601f \
 //x=4.725 //y=1.65 //x2=4.105 //y2=1.915
cc_513 ( N_noxref_5_c_663_n N_noxref_6_c_834_n ) capacitor c=0.00637984f \
 //x=4.455 //y=1.65 //x2=4.105 //y2=1.915
cc_514 ( N_noxref_5_c_629_n N_noxref_6_c_834_n ) capacitor c=0.0185661f \
 //x=4.81 //y=3.7 //x2=4.105 //y2=1.915
cc_515 ( N_noxref_5_M2_noxref_d N_noxref_6_c_834_n ) capacitor c=0.00643086f \
 //x=4.18 //y=0.905 //x2=4.105 //y2=1.915
cc_516 ( N_noxref_5_M2_noxref_d N_noxref_6_c_879_n ) capacitor c=0.00241053f \
 //x=4.18 //y=0.905 //x2=4.48 //y2=0.75
cc_517 ( N_noxref_5_c_628_n N_noxref_6_c_880_n ) capacitor c=0.00196666f \
 //x=4.725 //y=1.65 //x2=4.48 //y2=1.405
cc_518 ( N_noxref_5_M2_noxref_d N_noxref_6_c_880_n ) capacitor c=0.0124466f \
 //x=4.18 //y=0.905 //x2=4.48 //y2=1.405
cc_519 ( N_noxref_5_M2_noxref_d N_noxref_6_c_836_n ) capacitor c=0.00132245f \
 //x=4.18 //y=0.905 //x2=4.635 //y2=0.905
cc_520 ( N_noxref_5_c_628_n N_noxref_6_c_837_n ) capacitor c=0.00423452f \
 //x=4.725 //y=1.65 //x2=4.635 //y2=1.25
cc_521 ( N_noxref_5_M2_noxref_d N_noxref_6_c_837_n ) capacitor c=0.00566463f \
 //x=4.18 //y=0.905 //x2=4.635 //y2=1.25
cc_522 ( N_noxref_5_c_632_n N_noxref_6_M5_noxref_d ) capacitor c=2.77389e-19 \
 //x=8.14 //y=3.7 //x2=9.795 //y2=0.91
cc_523 ( N_noxref_5_c_632_n N_noxref_6_M16_noxref_d ) capacitor c=7.99492e-19 \
 //x=8.14 //y=3.7 //x2=9.84 //y2=5.02
cc_524 ( N_noxref_5_c_657_n N_noxref_7_c_976_n ) capacitor c=0.304761f \
 //x=8.025 //y=3.7 //x2=10.245 //y2=4.07
cc_525 ( N_noxref_5_c_655_n N_noxref_7_c_976_n ) capacitor c=0.0293665f \
 //x=4.925 //y=3.7 //x2=10.245 //y2=4.07
cc_526 ( N_noxref_5_c_640_n N_noxref_7_c_976_n ) capacitor c=0.00431193f \
 //x=4.725 //y=5.205 //x2=10.245 //y2=4.07
cc_527 ( N_noxref_5_c_629_n N_noxref_7_c_976_n ) capacitor c=0.0229481f \
 //x=4.81 //y=3.7 //x2=10.245 //y2=4.07
cc_528 ( N_noxref_5_c_632_n N_noxref_7_c_976_n ) capacitor c=0.0176431f \
 //x=8.14 //y=3.7 //x2=10.245 //y2=4.07
cc_529 ( N_noxref_5_c_640_n N_noxref_7_c_984_n ) capacitor c=0.00102585f \
 //x=4.725 //y=5.205 //x2=4.555 //y2=4.07
cc_530 ( N_noxref_5_c_642_n N_noxref_7_c_984_n ) capacitor c=0.00142608f \
 //x=4.415 //y=5.205 //x2=4.555 //y2=4.07
cc_531 ( N_noxref_5_c_629_n N_noxref_7_c_984_n ) capacitor c=0.00168517f \
 //x=4.81 //y=3.7 //x2=4.555 //y2=4.07
cc_532 ( N_noxref_5_c_657_n N_noxref_7_c_947_n ) capacitor c=0.139121f \
 //x=8.025 //y=3.7 //x2=10.245 //y2=3.33
cc_533 ( N_noxref_5_c_632_n N_noxref_7_c_947_n ) capacitor c=0.0181506f \
 //x=8.14 //y=3.7 //x2=10.245 //y2=3.33
cc_534 ( N_noxref_5_c_657_n N_noxref_7_c_1018_n ) capacitor c=0.0286718f \
 //x=8.025 //y=3.7 //x2=6.775 //y2=3.33
cc_535 ( N_noxref_5_c_629_n N_noxref_7_c_1018_n ) capacitor c=0.00286475f \
 //x=4.81 //y=3.7 //x2=6.775 //y2=3.33
cc_536 ( N_noxref_5_c_642_n N_noxref_7_c_985_n ) capacitor c=0.0123412f \
 //x=4.415 //y=5.205 //x2=4.44 //y2=4.07
cc_537 ( N_noxref_5_c_629_n N_noxref_7_c_985_n ) capacitor c=0.0637046f \
 //x=4.81 //y=3.7 //x2=4.44 //y2=4.07
cc_538 ( N_noxref_5_c_657_n N_noxref_7_c_950_n ) capacitor c=0.00490285f \
 //x=8.025 //y=3.7 //x2=6.66 //y2=2.08
cc_539 ( N_noxref_5_c_629_n N_noxref_7_c_950_n ) capacitor c=0.00705644f \
 //x=4.81 //y=3.7 //x2=6.66 //y2=2.08
cc_540 ( N_noxref_5_c_632_n N_noxref_7_c_950_n ) capacitor c=0.00348039f \
 //x=8.14 //y=3.7 //x2=6.66 //y2=2.08
cc_541 ( N_noxref_5_c_632_n N_noxref_7_c_951_n ) capacitor c=0.00139461f \
 //x=8.14 //y=3.7 //x2=10.36 //y2=2.085
cc_542 ( N_noxref_5_c_642_n N_noxref_7_M10_noxref_g ) capacitor c=0.0132788f \
 //x=4.415 //y=5.205 //x2=4.11 //y2=6.02
cc_543 ( N_noxref_5_c_640_n N_noxref_7_M11_noxref_g ) capacitor c=0.0187432f \
 //x=4.725 //y=5.205 //x2=4.55 //y2=6.02
cc_544 ( N_noxref_5_M10_noxref_d N_noxref_7_M11_noxref_g ) capacitor \
 c=0.0136385f //x=4.185 //y=5.02 //x2=4.55 //y2=6.02
cc_545 ( N_noxref_5_c_640_n N_noxref_7_c_1011_n ) capacitor c=0.00161455f \
 //x=4.725 //y=5.205 //x2=4.44 //y2=4.7
cc_546 ( N_noxref_5_c_642_n N_noxref_7_c_1011_n ) capacitor c=0.00557817f \
 //x=4.415 //y=5.205 //x2=4.44 //y2=4.7
cc_547 ( N_noxref_5_c_629_n N_noxref_7_c_1011_n ) capacitor c=0.0232466f \
 //x=4.81 //y=3.7 //x2=4.44 //y2=4.7
cc_548 ( N_noxref_5_c_642_n N_noxref_8_c_1119_n ) capacitor c=0.0348754f \
 //x=4.415 //y=5.205 //x2=3.805 //y2=5.205
cc_549 ( N_noxref_5_c_640_n N_noxref_8_c_1126_n ) capacitor c=0.0015978f \
 //x=4.725 //y=5.205 //x2=4.685 //y2=6.905
cc_550 ( N_noxref_5_M10_noxref_d N_noxref_8_c_1126_n ) capacitor c=0.01159f \
 //x=4.185 //y=5.02 //x2=4.685 //y2=6.905
cc_551 ( N_noxref_5_M10_noxref_d N_noxref_8_M8_noxref_s ) capacitor \
 c=0.00107541f //x=4.185 //y=5.02 //x2=2.875 //y2=5.02
cc_552 ( N_noxref_5_M10_noxref_d N_noxref_8_M9_noxref_d ) capacitor \
 c=0.0348754f //x=4.185 //y=5.02 //x2=3.745 //y2=5.02
cc_553 ( N_noxref_5_c_640_n N_noxref_8_M11_noxref_d ) capacitor c=0.0154558f \
 //x=4.725 //y=5.205 //x2=4.625 //y2=5.02
cc_554 ( N_noxref_5_M10_noxref_d N_noxref_8_M11_noxref_d ) capacitor \
 c=0.0458293f //x=4.185 //y=5.02 //x2=4.625 //y2=5.02
cc_555 ( N_noxref_5_c_663_n N_noxref_9_c_1159_n ) capacitor c=2.94752e-19 \
 //x=4.455 //y=1.65 //x2=2.915 //y2=1.495
cc_556 ( N_noxref_5_c_663_n N_noxref_9_c_1168_n ) capacitor c=0.0200666f \
 //x=4.455 //y=1.65 //x2=3.885 //y2=1.495
cc_557 ( N_noxref_5_c_628_n N_noxref_9_c_1169_n ) capacitor c=0.00457164f \
 //x=4.725 //y=1.65 //x2=4.77 //y2=0.53
cc_558 ( N_noxref_5_M2_noxref_d N_noxref_9_c_1169_n ) capacitor c=0.0113664f \
 //x=4.18 //y=0.905 //x2=4.77 //y2=0.53
cc_559 ( N_noxref_5_c_628_n N_noxref_9_M1_noxref_s ) capacitor c=0.0141104f \
 //x=4.725 //y=1.65 //x2=2.78 //y2=0.365
cc_560 ( N_noxref_5_M2_noxref_d N_noxref_9_M1_noxref_s ) capacitor \
 c=0.0436902f //x=4.18 //y=0.905 //x2=2.78 //y2=0.365
cc_561 ( N_noxref_5_c_647_n N_noxref_10_c_1211_n ) capacitor c=0.0348754f \
 //x=7.745 //y=5.205 //x2=7.135 //y2=5.205
cc_562 ( N_noxref_5_c_640_n N_noxref_10_c_1216_n ) capacitor c=2.91997e-19 \
 //x=4.725 //y=5.205 //x2=6.425 //y2=5.205
cc_563 ( N_noxref_5_c_645_n N_noxref_10_c_1217_n ) capacitor c=0.00157156f \
 //x=8.055 //y=5.205 //x2=8.015 //y2=6.905
cc_564 ( N_noxref_5_M14_noxref_d N_noxref_10_c_1217_n ) capacitor c=0.011538f \
 //x=7.515 //y=5.02 //x2=8.015 //y2=6.905
cc_565 ( N_noxref_5_M10_noxref_d N_noxref_10_M12_noxref_s ) capacitor \
 c=4.36987e-19 //x=4.185 //y=5.02 //x2=6.205 //y2=5.02
cc_566 ( N_noxref_5_M14_noxref_d N_noxref_10_M12_noxref_s ) capacitor \
 c=0.00107541f //x=7.515 //y=5.02 //x2=6.205 //y2=5.02
cc_567 ( N_noxref_5_M14_noxref_d N_noxref_10_M13_noxref_d ) capacitor \
 c=0.0348754f //x=7.515 //y=5.02 //x2=7.075 //y2=5.02
cc_568 ( N_noxref_5_c_645_n N_noxref_10_M15_noxref_d ) capacitor c=0.0151541f \
 //x=8.055 //y=5.205 //x2=7.955 //y2=5.02
cc_569 ( N_noxref_5_M14_noxref_d N_noxref_10_M15_noxref_d ) capacitor \
 c=0.0458293f //x=7.515 //y=5.02 //x2=7.955 //y2=5.02
cc_570 ( N_noxref_5_c_628_n N_noxref_11_c_1278_n ) capacitor c=3.32751e-19 \
 //x=4.725 //y=1.65 //x2=6.245 //y2=1.495
cc_571 ( N_noxref_5_c_676_n N_noxref_11_c_1278_n ) capacitor c=2.94752e-19 \
 //x=7.785 //y=1.65 //x2=6.245 //y2=1.495
cc_572 ( N_noxref_5_c_676_n N_noxref_11_c_1262_n ) capacitor c=0.0202508f \
 //x=7.785 //y=1.65 //x2=7.215 //y2=1.495
cc_573 ( N_noxref_5_c_630_n N_noxref_11_c_1263_n ) capacitor c=0.00458486f \
 //x=8.055 //y=1.65 //x2=8.1 //y2=0.53
cc_574 ( N_noxref_5_M4_noxref_d N_noxref_11_c_1263_n ) capacitor c=0.0113622f \
 //x=7.51 //y=0.905 //x2=8.1 //y2=0.53
cc_575 ( N_noxref_5_c_630_n N_noxref_11_M3_noxref_s ) capacitor c=0.0143541f \
 //x=8.055 //y=1.65 //x2=6.11 //y2=0.365
cc_576 ( N_noxref_5_M4_noxref_d N_noxref_11_M3_noxref_s ) capacitor \
 c=0.0438744f //x=7.51 //y=0.905 //x2=6.11 //y2=0.365
cc_577 ( N_noxref_6_c_777_n N_noxref_7_c_976_n ) capacitor c=0.016678f \
 //x=9.505 //y=2.96 //x2=10.245 //y2=4.07
cc_578 ( N_noxref_6_c_795_n N_noxref_7_c_976_n ) capacitor c=0.267882f \
 //x=9.505 //y=4.44 //x2=10.245 //y2=4.07
cc_579 ( N_noxref_6_c_801_n N_noxref_7_c_976_n ) capacitor c=0.0286084f \
 //x=6.775 //y=4.44 //x2=10.245 //y2=4.07
cc_580 ( N_noxref_6_c_803_n N_noxref_7_c_976_n ) capacitor c=0.00480464f \
 //x=6.66 //y=4.44 //x2=10.245 //y2=4.07
cc_581 ( N_noxref_6_c_785_n N_noxref_7_c_976_n ) capacitor c=0.0218892f \
 //x=9.62 //y=2.96 //x2=10.245 //y2=4.07
cc_582 ( N_noxref_6_c_806_n N_noxref_7_c_976_n ) capacitor c=0.0104128f \
 //x=9.9 //y=4.58 //x2=10.245 //y2=4.07
cc_583 ( N_noxref_6_c_807_n N_noxref_7_c_976_n ) capacitor c=0.00207246f \
 //x=9.705 //y=4.58 //x2=10.245 //y2=4.07
cc_584 ( N_noxref_6_c_816_n N_noxref_7_c_976_n ) capacitor c=6.08197e-19 \
 //x=6.66 //y=4.7 //x2=10.245 //y2=4.07
cc_585 ( N_noxref_6_c_823_n N_noxref_7_c_984_n ) capacitor c=0.00956039f \
 //x=4.555 //y=2.96 //x2=4.555 //y2=4.07
cc_586 ( N_noxref_6_c_783_n N_noxref_7_c_984_n ) capacitor c=2.06418e-19 \
 //x=4.44 //y=2.08 //x2=4.555 //y2=4.07
cc_587 ( N_noxref_6_c_777_n N_noxref_7_c_947_n ) capacitor c=0.269451f \
 //x=9.505 //y=2.96 //x2=10.245 //y2=3.33
cc_588 ( N_noxref_6_c_795_n N_noxref_7_c_947_n ) capacitor c=0.00458832f \
 //x=9.505 //y=4.44 //x2=10.245 //y2=3.33
cc_589 ( N_noxref_6_c_785_n N_noxref_7_c_947_n ) capacitor c=0.023832f \
 //x=9.62 //y=2.96 //x2=10.245 //y2=3.33
cc_590 ( N_noxref_6_c_786_n N_noxref_7_c_947_n ) capacitor c=0.00433609f \
 //x=9.905 //y=2.08 //x2=10.245 //y2=3.33
cc_591 ( N_noxref_6_c_777_n N_noxref_7_c_1018_n ) capacitor c=0.029123f \
 //x=9.505 //y=2.96 //x2=6.775 //y2=3.33
cc_592 ( N_noxref_6_c_823_n N_noxref_7_c_985_n ) capacitor c=2.06418e-19 \
 //x=4.555 //y=2.96 //x2=4.44 //y2=4.07
cc_593 ( N_noxref_6_c_783_n N_noxref_7_c_985_n ) capacitor c=0.0091252f \
 //x=4.44 //y=2.08 //x2=4.44 //y2=4.07
cc_594 ( N_noxref_6_c_777_n N_noxref_7_c_950_n ) capacitor c=0.0215795f \
 //x=9.505 //y=2.96 //x2=6.66 //y2=2.08
cc_595 ( N_noxref_6_c_783_n N_noxref_7_c_950_n ) capacitor c=3.72011e-19 \
 //x=4.44 //y=2.08 //x2=6.66 //y2=2.08
cc_596 ( N_noxref_6_c_803_n N_noxref_7_c_950_n ) capacitor c=0.00883256f \
 //x=6.66 //y=4.44 //x2=6.66 //y2=2.08
cc_597 ( N_noxref_6_c_777_n N_noxref_7_c_951_n ) capacitor c=0.00599141f \
 //x=9.505 //y=2.96 //x2=10.36 //y2=2.085
cc_598 ( N_noxref_6_c_795_n N_noxref_7_c_951_n ) capacitor c=0.00569864f \
 //x=9.505 //y=4.44 //x2=10.36 //y2=2.085
cc_599 ( N_noxref_6_c_785_n N_noxref_7_c_951_n ) capacitor c=0.0635926f \
 //x=9.62 //y=2.96 //x2=10.36 //y2=2.085
cc_600 ( N_noxref_6_c_806_n N_noxref_7_c_951_n ) capacitor c=0.0248426f \
 //x=9.9 //y=4.58 //x2=10.36 //y2=2.085
cc_601 ( N_noxref_6_c_807_n N_noxref_7_c_951_n ) capacitor c=8.0359e-19 \
 //x=9.705 //y=4.58 //x2=10.36 //y2=2.085
cc_602 ( N_noxref_6_M5_noxref_d N_noxref_7_c_951_n ) capacitor c=0.0175773f \
 //x=9.795 //y=0.91 //x2=10.36 //y2=2.085
cc_603 ( N_noxref_6_M16_noxref_d N_noxref_7_M16_noxref_g ) capacitor \
 c=0.021902f //x=9.84 //y=5.02 //x2=9.765 //y2=6.02
cc_604 ( N_noxref_6_M16_noxref_d N_noxref_7_M17_noxref_g ) capacitor \
 c=0.0219309f //x=9.84 //y=5.02 //x2=10.205 //y2=6.02
cc_605 ( N_noxref_6_M5_noxref_d N_noxref_7_c_966_n ) capacitor c=0.00216577f \
 //x=9.795 //y=0.91 //x2=9.72 //y2=0.91
cc_606 ( N_noxref_6_c_786_n N_noxref_7_c_968_n ) capacitor c=0.0023507f \
 //x=9.905 //y=2.08 //x2=9.72 //y2=1.255
cc_607 ( N_noxref_6_M5_noxref_d N_noxref_7_c_968_n ) capacitor c=0.00599232f \
 //x=9.795 //y=0.91 //x2=9.72 //y2=1.255
cc_608 ( N_noxref_6_c_806_n N_noxref_7_c_1091_n ) capacitor c=0.00494191f \
 //x=9.9 //y=4.58 //x2=10.13 //y2=4.79
cc_609 ( N_noxref_6_M16_noxref_d N_noxref_7_c_1091_n ) capacitor c=0.0146106f \
 //x=9.84 //y=5.02 //x2=10.13 //y2=4.79
cc_610 ( N_noxref_6_c_807_n N_noxref_7_c_999_n ) capacitor c=0.00494191f \
 //x=9.705 //y=4.58 //x2=9.84 //y2=4.79
cc_611 ( N_noxref_6_M5_noxref_d N_noxref_7_c_969_n ) capacitor c=0.00220879f \
 //x=9.795 //y=0.91 //x2=10.095 //y2=0.755
cc_612 ( N_noxref_6_M5_noxref_d N_noxref_7_c_1095_n ) capacitor c=0.0138447f \
 //x=9.795 //y=0.91 //x2=10.095 //y2=1.41
cc_613 ( N_noxref_6_c_806_n N_noxref_7_c_1000_n ) capacitor c=0.00944945f \
 //x=9.9 //y=4.58 //x2=10.205 //y2=4.865
cc_614 ( N_noxref_6_M16_noxref_d N_noxref_7_c_1000_n ) capacitor c=0.00307344f \
 //x=9.84 //y=5.02 //x2=10.205 //y2=4.865
cc_615 ( N_noxref_6_M5_noxref_d N_noxref_7_c_970_n ) capacitor c=0.00220616f \
 //x=9.795 //y=0.91 //x2=10.25 //y2=0.91
cc_616 ( N_noxref_6_M5_noxref_d N_noxref_7_c_1099_n ) capacitor c=0.00347355f \
 //x=9.795 //y=0.91 //x2=10.25 //y2=1.255
cc_617 ( N_noxref_6_M5_noxref_d N_noxref_7_c_1100_n ) capacitor c=0.007449f \
 //x=9.795 //y=0.91 //x2=10.25 //y2=1.565
cc_618 ( N_noxref_6_M5_noxref_d N_noxref_7_c_972_n ) capacitor c=0.00957707f \
 //x=9.795 //y=0.91 //x2=10.25 //y2=1.92
cc_619 ( N_noxref_6_c_785_n N_noxref_7_c_973_n ) capacitor c=8.49451e-19 \
 //x=9.62 //y=2.96 //x2=10.25 //y2=2.085
cc_620 ( N_noxref_6_c_786_n N_noxref_7_c_973_n ) capacitor c=0.0167852f \
 //x=9.905 //y=2.08 //x2=10.25 //y2=2.085
cc_621 ( N_noxref_6_c_831_n N_noxref_9_c_1168_n ) capacitor c=0.00628626f \
 //x=4.105 //y=1.56 //x2=3.885 //y2=1.495
cc_622 ( N_noxref_6_c_826_n N_noxref_9_c_1169_n ) capacitor c=0.0197889f \
 //x=4.105 //y=0.905 //x2=4.77 //y2=0.53
cc_623 ( N_noxref_6_c_836_n N_noxref_9_c_1169_n ) capacitor c=0.00655813f \
 //x=4.635 //y=0.905 //x2=4.77 //y2=0.53
cc_624 ( N_noxref_6_c_826_n N_noxref_9_M1_noxref_s ) capacitor c=0.00628626f \
 //x=4.105 //y=0.905 //x2=2.78 //y2=0.365
cc_625 ( N_noxref_6_c_836_n N_noxref_9_M1_noxref_s ) capacitor c=0.0143002f \
 //x=4.635 //y=0.905 //x2=2.78 //y2=0.365
cc_626 ( N_noxref_6_c_837_n N_noxref_9_M1_noxref_s ) capacitor c=0.00290153f \
 //x=4.635 //y=1.25 //x2=2.78 //y2=0.365
cc_627 ( N_noxref_6_c_795_n N_noxref_10_c_1211_n ) capacitor c=0.0172642f \
 //x=9.505 //y=4.44 //x2=7.135 //y2=5.205
cc_628 ( N_noxref_6_c_801_n N_noxref_10_c_1211_n ) capacitor c=0.00485884f \
 //x=6.775 //y=4.44 //x2=7.135 //y2=5.205
cc_629 ( N_noxref_6_c_803_n N_noxref_10_c_1211_n ) capacitor c=0.0111238f \
 //x=6.66 //y=4.44 //x2=7.135 //y2=5.205
cc_630 ( N_noxref_6_M12_noxref_g N_noxref_10_c_1211_n ) capacitor c=0.018644f \
 //x=6.56 //y=6.02 //x2=7.135 //y2=5.205
cc_631 ( N_noxref_6_M13_noxref_g N_noxref_10_c_1211_n ) capacitor c=0.0169648f \
 //x=7 //y=6.02 //x2=7.135 //y2=5.205
cc_632 ( N_noxref_6_c_816_n N_noxref_10_c_1211_n ) capacitor c=0.00531676f \
 //x=6.66 //y=4.7 //x2=7.135 //y2=5.205
cc_633 ( N_noxref_6_c_795_n N_noxref_10_c_1217_n ) capacitor c=0.00389598f \
 //x=9.505 //y=4.44 //x2=8.015 //y2=6.905
cc_634 ( N_noxref_6_M12_noxref_g N_noxref_10_M12_noxref_s ) capacitor \
 c=0.0441361f //x=6.56 //y=6.02 //x2=6.205 //y2=5.02
cc_635 ( N_noxref_6_M13_noxref_g N_noxref_10_M13_noxref_d ) capacitor \
 c=0.0170604f //x=7 //y=6.02 //x2=7.075 //y2=5.02
cc_636 ( N_noxref_6_c_777_n N_noxref_11_M3_noxref_s ) capacitor c=6.20367e-19 \
 //x=9.505 //y=2.96 //x2=6.11 //y2=0.365
cc_637 ( N_noxref_7_M10_noxref_g N_noxref_8_c_1119_n ) capacitor c=0.0170604f \
 //x=4.11 //y=6.02 //x2=3.805 //y2=5.205
cc_638 ( N_noxref_7_M10_noxref_g N_noxref_8_c_1126_n ) capacitor c=0.0150677f \
 //x=4.11 //y=6.02 //x2=4.685 //y2=6.905
cc_639 ( N_noxref_7_M11_noxref_g N_noxref_8_c_1126_n ) capacitor c=0.016333f \
 //x=4.55 //y=6.02 //x2=4.685 //y2=6.905
cc_640 ( N_noxref_7_M11_noxref_g N_noxref_8_M11_noxref_d ) capacitor \
 c=0.0351101f //x=4.55 //y=6.02 //x2=4.625 //y2=5.02
cc_641 ( N_noxref_7_c_976_n N_noxref_10_c_1216_n ) capacitor c=0.0060417f \
 //x=10.245 //y=4.07 //x2=6.425 //y2=5.205
cc_642 ( N_noxref_7_c_960_n N_noxref_11_c_1278_n ) capacitor c=0.0034165f \
 //x=6.465 //y=1.915 //x2=6.245 //y2=1.495
cc_643 ( N_noxref_7_c_950_n N_noxref_11_c_1254_n ) capacitor c=0.0113474f \
 //x=6.66 //y=2.08 //x2=7.13 //y2=1.58
cc_644 ( N_noxref_7_c_959_n N_noxref_11_c_1254_n ) capacitor c=0.00703567f \
 //x=6.465 //y=1.52 //x2=7.13 //y2=1.58
cc_645 ( N_noxref_7_c_960_n N_noxref_11_c_1254_n ) capacitor c=0.018562f \
 //x=6.465 //y=1.915 //x2=7.13 //y2=1.58
cc_646 ( N_noxref_7_c_962_n N_noxref_11_c_1254_n ) capacitor c=0.00780629f \
 //x=6.84 //y=1.365 //x2=7.13 //y2=1.58
cc_647 ( N_noxref_7_c_965_n N_noxref_11_c_1254_n ) capacitor c=0.00339872f \
 //x=6.995 //y=1.21 //x2=7.13 //y2=1.58
cc_648 ( N_noxref_7_c_960_n N_noxref_11_c_1262_n ) capacitor c=6.71402e-19 \
 //x=6.465 //y=1.915 //x2=7.215 //y2=1.495
cc_649 ( N_noxref_7_c_956_n N_noxref_11_M3_noxref_s ) capacitor c=0.0326577f \
 //x=6.465 //y=0.865 //x2=6.11 //y2=0.365
cc_650 ( N_noxref_7_c_959_n N_noxref_11_M3_noxref_s ) capacitor c=3.48408e-19 \
 //x=6.465 //y=1.52 //x2=6.11 //y2=0.365
cc_651 ( N_noxref_7_c_963_n N_noxref_11_M3_noxref_s ) capacitor c=0.0120759f \
 //x=6.995 //y=0.865 //x2=6.11 //y2=0.365
cc_652 ( N_noxref_8_M11_noxref_d N_noxref_10_M12_noxref_s ) capacitor \
 c=0.00181587f //x=4.625 //y=5.02 //x2=6.205 //y2=5.02
cc_653 ( N_noxref_9_c_1172_n N_noxref_11_M3_noxref_s ) capacitor c=0.00174327f \
 //x=4.855 //y=0.615 //x2=6.11 //y2=0.365
