* SPICE3 file created from XOR2X1.ext - technology: sky130A

.subckt XOR2X1 Y A B VPB VNB
M1000 a_575_1004.t1 a_807_943.t3 Y pshort w=2u l=0.15u
+  ad=0p pd=0u as=1.16p ps=9.16u
M1001 VNB A a_556_74.t0 nshort w=-1.605u l=1.765u
+  ad=2.6398p pd=19.34u as=0p ps=0u
M1002 a_1241_1004.t1 B VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y a_807_943.t4 a_575_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1241_1004.t2 a_185_182.t4 Y pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y a_185_182.t3 a_1222_74.t0 nshort w=-1.605u l=1.765u
+  ad=0.3582p pd=3.14u as=0p ps=0u
M1006 VPB.t3 B a_807_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPB.t5 A a_575_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_807_943.t2 B VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B a_556_74.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPB.t6 A a_185_182.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPB.t1 B a_1241_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_575_1004.t3 A VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y a_185_182.t5 a_1241_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VNB a_807_943.t5 a_1222_74.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_185_182.t1 A VPB.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 B A 0.06fF
C1 VPB B 0.38fF
C2 VPB A 0.34fF
C3 Y B 0.81fF
C4 Y A 0.07fF
C5 Y VPB 0.53fF
R0 a_807_943.n2 a_807_943.t4 477.179
R1 a_807_943.n4 a_807_943.t5 420.747
R2 a_807_943.n2 a_807_943.t3 406.485
R3 a_807_943.n3 a_807_943.n2 211.151
R4 a_807_943.n6 a_807_943.n4 188.704
R5 a_807_943.n3 a_807_943.n1 114.038
R6 a_807_943.n4 a_807_943.n3 53.105
R7 a_807_943.n6 a_807_943.n5 30
R8 a_807_943.n7 a_807_943.n0 24.383
R9 a_807_943.n7 a_807_943.n6 23.684
R10 a_807_943.n1 a_807_943.t1 14.282
R11 a_807_943.n1 a_807_943.t2 14.282
R12 a_575_1004.t1 a_575_1004.n0 101.663
R13 a_575_1004.n0 a_575_1004.t2 101.661
R14 a_575_1004.n0 a_575_1004.t0 14.294
R15 a_575_1004.n0 a_575_1004.t3 14.282
R16 VPB VPB.n227 126.832
R17 VPB.n60 VPB.n58 94.117
R18 VPB.n202 VPB.n200 94.117
R19 VPB.n132 VPB.n130 94.117
R20 VPB.n184 VPB.n178 76.136
R21 VPB.n184 VPB.n183 76
R22 VPB.n198 VPB.n195 76
R23 VPB.n204 VPB.n203 76
R24 VPB.n208 VPB.n207 76
R25 VPB.n220 VPB.n219 76
R26 VPB.n181 VPB.n180 68.979
R27 VPB.n71 VPB.n70 68.979
R28 VPB.n46 VPB.n35 65.944
R29 VPB.n147 VPB.n96 65.944
R30 VPB.n122 VPB.n121 64.528
R31 VPB.n64 VPB.n63 64.528
R32 VPB.n20 VPB.n19 61.764
R33 VPB.n81 VPB.n80 61.764
R34 VPB.n103 VPB.n102 61.764
R35 VPB.n74 VPB.t7 55.106
R36 VPB.n62 VPB.t6 55.106
R37 VPB.n125 VPB.t2 55.106
R38 VPB.n179 VPB.t3 55.106
R39 VPB.n149 VPB.n148 44.502
R40 VPB.n48 VPB.n47 44.502
R41 VPB.n224 VPB.n220 20.452
R42 VPB.n178 VPB.n175 20.452
R43 VPB.n35 VPB.t4 14.282
R44 VPB.n35 VPB.t5 14.282
R45 VPB.n96 VPB.t0 14.282
R46 VPB.n96 VPB.t1 14.282
R47 VPB.n178 VPB.n177 13.653
R48 VPB.n177 VPB.n176 13.653
R49 VPB.n183 VPB.n182 13.653
R50 VPB.n182 VPB.n181 13.653
R51 VPB.n120 VPB.n119 13.653
R52 VPB.n119 VPB.n118 13.653
R53 VPB.n124 VPB.n123 13.653
R54 VPB.n123 VPB.n122 13.653
R55 VPB.n128 VPB.n127 13.653
R56 VPB.n127 VPB.n126 13.653
R57 VPB.n133 VPB.n132 13.653
R58 VPB.n132 VPB.n131 13.653
R59 VPB.n136 VPB.n135 13.653
R60 VPB.n135 VPB.n134 13.653
R61 VPB.n139 VPB.n138 13.653
R62 VPB.n138 VPB.n137 13.653
R63 VPB.n142 VPB.n141 13.653
R64 VPB.n141 VPB.n140 13.653
R65 VPB.n146 VPB.n145 13.653
R66 VPB.n145 VPB.n144 13.653
R67 VPB.n151 VPB.n150 13.653
R68 VPB.n150 VPB.n149 13.653
R69 VPB.n154 VPB.n153 13.653
R70 VPB.n153 VPB.n152 13.653
R71 VPB.n198 VPB.n197 13.653
R72 VPB.n197 VPB.n196 13.653
R73 VPB.n203 VPB.n202 13.653
R74 VPB.n202 VPB.n201 13.653
R75 VPB.n207 VPB.n206 13.653
R76 VPB.n206 VPB.n205 13.653
R77 VPB.n38 VPB.n37 13.653
R78 VPB.n37 VPB.n36 13.653
R79 VPB.n41 VPB.n40 13.653
R80 VPB.n40 VPB.n39 13.653
R81 VPB.n45 VPB.n44 13.653
R82 VPB.n44 VPB.n43 13.653
R83 VPB.n50 VPB.n49 13.653
R84 VPB.n49 VPB.n48 13.653
R85 VPB.n53 VPB.n52 13.653
R86 VPB.n52 VPB.n51 13.653
R87 VPB.n56 VPB.n55 13.653
R88 VPB.n55 VPB.n54 13.653
R89 VPB.n61 VPB.n60 13.653
R90 VPB.n60 VPB.n59 13.653
R91 VPB.n66 VPB.n65 13.653
R92 VPB.n65 VPB.n64 13.653
R93 VPB.n69 VPB.n68 13.653
R94 VPB.n68 VPB.n67 13.653
R95 VPB.n73 VPB.n72 13.653
R96 VPB.n72 VPB.n71 13.653
R97 VPB.n220 VPB.n0 13.653
R98 VPB VPB.n0 13.653
R99 VPB.n144 VPB.n143 13.35
R100 VPB.n43 VPB.n42 13.35
R101 VPB.n224 VPB.n223 13.276
R102 VPB.n223 VPB.n221 13.276
R103 VPB.n34 VPB.n16 13.276
R104 VPB.n16 VPB.n14 13.276
R105 VPB.n95 VPB.n77 13.276
R106 VPB.n77 VPB.n75 13.276
R107 VPB.n117 VPB.n99 13.276
R108 VPB.n99 VPB.n97 13.276
R109 VPB.n124 VPB.n120 13.276
R110 VPB.n129 VPB.n128 13.276
R111 VPB.n133 VPB.n129 13.276
R112 VPB.n136 VPB.n133 13.276
R113 VPB.n139 VPB.n136 13.276
R114 VPB.n142 VPB.n139 13.276
R115 VPB.n146 VPB.n142 13.276
R116 VPB.n154 VPB.n151 13.276
R117 VPB.n198 VPB.n154 13.276
R118 VPB.n199 VPB.n198 13.276
R119 VPB.n203 VPB.n199 13.276
R120 VPB.n41 VPB.n38 13.276
R121 VPB.n45 VPB.n41 13.276
R122 VPB.n53 VPB.n50 13.276
R123 VPB.n56 VPB.n53 13.276
R124 VPB.n57 VPB.n56 13.276
R125 VPB.n61 VPB.n57 13.276
R126 VPB.n69 VPB.n66 13.276
R127 VPB.n73 VPB.n69 13.276
R128 VPB.n175 VPB.n157 13.276
R129 VPB.n157 VPB.n155 13.276
R130 VPB.n162 VPB.n160 12.796
R131 VPB.n162 VPB.n161 12.564
R132 VPB.n171 VPB.n170 12.198
R133 VPB.n168 VPB.n167 12.198
R134 VPB.n165 VPB.n164 12.198
R135 VPB.n220 VPB.n74 10.944
R136 VPB.n128 VPB.n125 10.585
R137 VPB.n62 VPB.n61 10.585
R138 VPB.n147 VPB.n146 8.97
R139 VPB.n46 VPB.n45 8.97
R140 VPB.n175 VPB.n174 7.5
R141 VPB.n160 VPB.n159 7.5
R142 VPB.n164 VPB.n163 7.5
R143 VPB.n167 VPB.n166 7.5
R144 VPB.n157 VPB.n156 7.5
R145 VPB.n172 VPB.n158 7.5
R146 VPB.n99 VPB.n98 7.5
R147 VPB.n112 VPB.n111 7.5
R148 VPB.n106 VPB.n105 7.5
R149 VPB.n108 VPB.n107 7.5
R150 VPB.n101 VPB.n100 7.5
R151 VPB.n117 VPB.n116 7.5
R152 VPB.n77 VPB.n76 7.5
R153 VPB.n90 VPB.n89 7.5
R154 VPB.n84 VPB.n83 7.5
R155 VPB.n86 VPB.n85 7.5
R156 VPB.n79 VPB.n78 7.5
R157 VPB.n95 VPB.n94 7.5
R158 VPB.n16 VPB.n15 7.5
R159 VPB.n29 VPB.n28 7.5
R160 VPB.n23 VPB.n22 7.5
R161 VPB.n25 VPB.n24 7.5
R162 VPB.n18 VPB.n17 7.5
R163 VPB.n34 VPB.n33 7.5
R164 VPB.n223 VPB.n222 7.5
R165 VPB.n12 VPB.n11 7.5
R166 VPB.n6 VPB.n5 7.5
R167 VPB.n8 VPB.n7 7.5
R168 VPB.n2 VPB.n1 7.5
R169 VPB.n225 VPB.n224 7.5
R170 VPB.n57 VPB.n34 7.176
R171 VPB.n199 VPB.n95 7.176
R172 VPB.n129 VPB.n117 7.176
R173 VPB.n113 VPB.n110 6.729
R174 VPB.n109 VPB.n106 6.729
R175 VPB.n104 VPB.n101 6.729
R176 VPB.n91 VPB.n88 6.729
R177 VPB.n87 VPB.n84 6.729
R178 VPB.n82 VPB.n79 6.729
R179 VPB.n30 VPB.n27 6.729
R180 VPB.n26 VPB.n23 6.729
R181 VPB.n21 VPB.n18 6.729
R182 VPB.n13 VPB.n10 6.729
R183 VPB.n9 VPB.n6 6.729
R184 VPB.n4 VPB.n2 6.729
R185 VPB.n104 VPB.n103 6.728
R186 VPB.n109 VPB.n108 6.728
R187 VPB.n113 VPB.n112 6.728
R188 VPB.n116 VPB.n115 6.728
R189 VPB.n82 VPB.n81 6.728
R190 VPB.n87 VPB.n86 6.728
R191 VPB.n91 VPB.n90 6.728
R192 VPB.n94 VPB.n93 6.728
R193 VPB.n21 VPB.n20 6.728
R194 VPB.n26 VPB.n25 6.728
R195 VPB.n30 VPB.n29 6.728
R196 VPB.n33 VPB.n32 6.728
R197 VPB.n4 VPB.n3 6.728
R198 VPB.n9 VPB.n8 6.728
R199 VPB.n13 VPB.n12 6.728
R200 VPB.n226 VPB.n225 6.728
R201 VPB.n174 VPB.n173 6.398
R202 VPB.n151 VPB.n147 4.305
R203 VPB.n50 VPB.n46 4.305
R204 VPB.n125 VPB.n124 2.691
R205 VPB.n66 VPB.n62 2.691
R206 VPB.n183 VPB.n179 2.332
R207 VPB.n74 VPB.n73 2.332
R208 VPB.n172 VPB.n165 1.402
R209 VPB.n172 VPB.n168 1.402
R210 VPB.n172 VPB.n169 1.402
R211 VPB.n172 VPB.n171 1.402
R212 VPB.n173 VPB.n172 0.735
R213 VPB.n172 VPB.n162 0.735
R214 VPB.n114 VPB.n113 0.387
R215 VPB.n114 VPB.n109 0.387
R216 VPB.n114 VPB.n104 0.387
R217 VPB.n115 VPB.n114 0.387
R218 VPB.n92 VPB.n91 0.387
R219 VPB.n92 VPB.n87 0.387
R220 VPB.n92 VPB.n82 0.387
R221 VPB.n93 VPB.n92 0.387
R222 VPB.n31 VPB.n30 0.387
R223 VPB.n31 VPB.n26 0.387
R224 VPB.n31 VPB.n21 0.387
R225 VPB.n32 VPB.n31 0.387
R226 VPB.n227 VPB.n13 0.387
R227 VPB.n227 VPB.n9 0.387
R228 VPB.n227 VPB.n4 0.387
R229 VPB.n227 VPB.n226 0.387
R230 VPB.n188 VPB.n187 0.272
R231 VPB.n215 VPB.n214 0.272
R232 VPB.n219 VPB 0.198
R233 VPB.n185 VPB.n184 0.136
R234 VPB.n186 VPB.n185 0.136
R235 VPB.n187 VPB.n186 0.136
R236 VPB.n189 VPB.n188 0.136
R237 VPB.n190 VPB.n189 0.136
R238 VPB.n191 VPB.n190 0.136
R239 VPB.n192 VPB.n191 0.136
R240 VPB.n193 VPB.n192 0.136
R241 VPB.n194 VPB.n193 0.136
R242 VPB.n195 VPB.n194 0.136
R243 VPB.n195 VPB 0.136
R244 VPB.n204 VPB 0.136
R245 VPB.n208 VPB.n204 0.136
R246 VPB.n209 VPB.n208 0.136
R247 VPB.n210 VPB.n209 0.136
R248 VPB.n211 VPB.n210 0.136
R249 VPB.n212 VPB.n211 0.136
R250 VPB.n213 VPB.n212 0.136
R251 VPB.n214 VPB.n213 0.136
R252 VPB.n216 VPB.n215 0.136
R253 VPB.n217 VPB.n216 0.136
R254 VPB.n218 VPB.n217 0.136
R255 VPB.n219 VPB.n218 0.136
R256 a_1241_1004.n0 a_1241_1004.t2 101.66
R257 a_1241_1004.n0 a_1241_1004.t0 101.66
R258 a_1241_1004.n0 a_1241_1004.t3 14.294
R259 a_1241_1004.t1 a_1241_1004.n0 14.282
R260 a_185_182.n2 a_185_182.t5 477.179
R261 a_185_182.n2 a_185_182.t4 406.485
R262 a_185_182.n3 a_185_182.t3 225.731
R263 a_185_182.n4 a_185_182.n1 220.249
R264 a_185_182.n3 a_185_182.n2 161.6
R265 a_185_182.n4 a_185_182.n3 156.579
R266 a_185_182.n6 a_185_182.n4 135.599
R267 a_185_182.n6 a_185_182.n5 30
R268 a_185_182.n7 a_185_182.n0 24.383
R269 a_185_182.n7 a_185_182.n6 23.684
R270 a_185_182.n1 a_185_182.t2 14.282
R271 a_185_182.n1 a_185_182.t1 14.282
R272 a_1222_74.t0 a_1222_74.n1 93.333
R273 a_1222_74.n4 a_1222_74.n2 55.07
R274 a_1222_74.t0 a_1222_74.n0 8.137
R275 a_1222_74.n4 a_1222_74.n3 4.619
R276 a_1222_74.t0 a_1222_74.n4 0.071
R277 VNB VNB.n222 300.778
R278 VNB.n102 VNB.n101 199.897
R279 VNB.n85 VNB.n84 199.897
R280 VNB.n25 VNB.n24 199.897
R281 VNB.n191 VNB.n189 154.509
R282 VNB.n127 VNB.n125 154.509
R283 VNB.n61 VNB.n59 154.509
R284 VNB.n42 VNB.n41 121.366
R285 VNB.n141 VNB.n91 85.201
R286 VNB.n173 VNB.n165 76.136
R287 VNB.n173 VNB.n172 76
R288 VNB.n209 VNB.n208 76
R289 VNB.n197 VNB.n196 76
R290 VNB.n193 VNB.n192 76
R291 VNB.n187 VNB.n184 76
R292 VNB.n46 VNB.n34 64.194
R293 VNB.n69 VNB.n68 49.896
R294 VNB.n43 VNB.n42 36.937
R295 VNB.n143 VNB.n142 36.678
R296 VNB.n14 VNB.n13 35.01
R297 VNB.t2 VNB.n6 32.601
R298 VNB.n34 VNB.n33 28.421
R299 VNB.n49 VNB.n48 27.855
R300 VNB.n34 VNB.n32 25.263
R301 VNB.n32 VNB.n31 24.383
R302 VNB.n165 VNB.n162 20.452
R303 VNB.n210 VNB.n209 20.452
R304 VNB.n169 VNB.n168 20.094
R305 VNB.n116 VNB.n112 20.094
R306 VNB.n120 VNB.n110 20.094
R307 VNB.n63 VNB.n14 20.094
R308 VNB.n67 VNB.n11 20.094
R309 VNB.n74 VNB.n9 20.094
R310 VNB.n14 VNB.n12 19.017
R311 VNB.n114 VNB.n113 18.269
R312 VNB.n109 VNB.t0 17.595
R313 VNB.n8 VNB.t2 17.353
R314 VNB.n50 VNB.n49 16.721
R315 VNB.n172 VNB.n171 13.653
R316 VNB.n171 VNB.n170 13.653
R317 VNB.n115 VNB.n114 13.653
R318 VNB.n119 VNB.n118 13.653
R319 VNB.n118 VNB.n117 13.653
R320 VNB.n123 VNB.n122 13.653
R321 VNB.n122 VNB.n121 13.653
R322 VNB.n128 VNB.n127 13.653
R323 VNB.n127 VNB.n126 13.653
R324 VNB.n131 VNB.n130 13.653
R325 VNB.n130 VNB.n129 13.653
R326 VNB.n134 VNB.n133 13.653
R327 VNB.n133 VNB.n132 13.653
R328 VNB.n137 VNB.n136 13.653
R329 VNB.n136 VNB.n135 13.653
R330 VNB.n140 VNB.n139 13.653
R331 VNB.n139 VNB.n138 13.653
R332 VNB.n144 VNB.n143 13.653
R333 VNB.n147 VNB.n146 13.653
R334 VNB.n146 VNB.n145 13.653
R335 VNB.n187 VNB.n186 13.653
R336 VNB.n186 VNB.n185 13.653
R337 VNB.n192 VNB.n191 13.653
R338 VNB.n191 VNB.n190 13.653
R339 VNB.n196 VNB.n195 13.653
R340 VNB.n195 VNB.n194 13.653
R341 VNB.n37 VNB.n36 13.653
R342 VNB.n36 VNB.n35 13.653
R343 VNB.n40 VNB.n39 13.653
R344 VNB.n39 VNB.n38 13.653
R345 VNB.n45 VNB.n44 13.653
R346 VNB.n44 VNB.n43 13.653
R347 VNB.n51 VNB.n50 13.653
R348 VNB.n54 VNB.n53 13.653
R349 VNB.n53 VNB.n52 13.653
R350 VNB.n57 VNB.n56 13.653
R351 VNB.n56 VNB.n55 13.653
R352 VNB.n62 VNB.n61 13.653
R353 VNB.n61 VNB.n60 13.653
R354 VNB.n66 VNB.n65 13.653
R355 VNB.n65 VNB.n64 13.653
R356 VNB.n70 VNB.n69 13.653
R357 VNB.n73 VNB.n72 13.653
R358 VNB.n72 VNB.n71 13.653
R359 VNB.n209 VNB.n0 13.653
R360 VNB VNB.n0 13.653
R361 VNB.n165 VNB.n164 13.653
R362 VNB.n164 VNB.n163 13.653
R363 VNB.n110 VNB.n109 13.608
R364 VNB.n217 VNB.n214 13.577
R365 VNB.n150 VNB.n148 13.276
R366 VNB.n162 VNB.n150 13.276
R367 VNB.n94 VNB.n92 13.276
R368 VNB.n107 VNB.n94 13.276
R369 VNB.n77 VNB.n75 13.276
R370 VNB.n90 VNB.n77 13.276
R371 VNB.n17 VNB.n15 13.276
R372 VNB.n30 VNB.n17 13.276
R373 VNB.n124 VNB.n123 13.276
R374 VNB.n128 VNB.n124 13.276
R375 VNB.n131 VNB.n128 13.276
R376 VNB.n134 VNB.n131 13.276
R377 VNB.n137 VNB.n134 13.276
R378 VNB.n140 VNB.n137 13.276
R379 VNB.n147 VNB.n144 13.276
R380 VNB.n187 VNB.n147 13.276
R381 VNB.n188 VNB.n187 13.276
R382 VNB.n192 VNB.n188 13.276
R383 VNB.n40 VNB.n37 13.276
R384 VNB.n45 VNB.n40 13.276
R385 VNB.n54 VNB.n51 13.276
R386 VNB.n57 VNB.n54 13.276
R387 VNB.n58 VNB.n57 13.276
R388 VNB.n62 VNB.n58 13.276
R389 VNB.n73 VNB.n70 13.276
R390 VNB.n3 VNB.n1 13.276
R391 VNB.n210 VNB.n3 13.276
R392 VNB.n119 VNB.n116 13.097
R393 VNB.n67 VNB.n66 13.097
R394 VNB.n9 VNB.n8 12.837
R395 VNB.n168 VNB.n167 10.853
R396 VNB.n141 VNB.n140 10.764
R397 VNB.n46 VNB.n45 10.764
R398 VNB.n167 VNB.n166 10.417
R399 VNB.n209 VNB.n74 9.329
R400 VNB.n123 VNB.n120 8.97
R401 VNB.n63 VNB.n62 8.97
R402 VNB.n109 VNB.n108 7.858
R403 VNB.n8 VNB.n7 7.566
R404 VNB.n219 VNB.n218 7.5
R405 VNB.n100 VNB.n99 7.5
R406 VNB.n96 VNB.n95 7.5
R407 VNB.n94 VNB.n93 7.5
R408 VNB.n107 VNB.n106 7.5
R409 VNB.n83 VNB.n82 7.5
R410 VNB.n79 VNB.n78 7.5
R411 VNB.n77 VNB.n76 7.5
R412 VNB.n90 VNB.n89 7.5
R413 VNB.n23 VNB.n22 7.5
R414 VNB.n19 VNB.n18 7.5
R415 VNB.n17 VNB.n16 7.5
R416 VNB.n30 VNB.n29 7.5
R417 VNB.n211 VNB.n210 7.5
R418 VNB.n3 VNB.n2 7.5
R419 VNB.n216 VNB.n215 7.5
R420 VNB.n156 VNB.n155 7.5
R421 VNB.n152 VNB.n151 7.5
R422 VNB.n150 VNB.n149 7.5
R423 VNB.n162 VNB.n161 7.5
R424 VNB.n124 VNB.n107 7.176
R425 VNB.n188 VNB.n90 7.176
R426 VNB.n58 VNB.n30 7.176
R427 VNB.n221 VNB.n219 7.011
R428 VNB.n103 VNB.n100 7.011
R429 VNB.n98 VNB.n96 7.011
R430 VNB.n86 VNB.n83 7.011
R431 VNB.n81 VNB.n79 7.011
R432 VNB.n26 VNB.n23 7.011
R433 VNB.n21 VNB.n19 7.011
R434 VNB.n158 VNB.n156 7.011
R435 VNB.n154 VNB.n152 7.011
R436 VNB.n106 VNB.n105 7.01
R437 VNB.n98 VNB.n97 7.01
R438 VNB.n103 VNB.n102 7.01
R439 VNB.n89 VNB.n88 7.01
R440 VNB.n81 VNB.n80 7.01
R441 VNB.n86 VNB.n85 7.01
R442 VNB.n29 VNB.n28 7.01
R443 VNB.n21 VNB.n20 7.01
R444 VNB.n26 VNB.n25 7.01
R445 VNB.n161 VNB.n160 7.01
R446 VNB.n154 VNB.n153 7.01
R447 VNB.n158 VNB.n157 7.01
R448 VNB.n221 VNB.n220 7.01
R449 VNB.n217 VNB.n216 6.788
R450 VNB.n212 VNB.n211 6.788
R451 VNB.n5 VNB.n4 4.551
R452 VNB.n120 VNB.n119 4.305
R453 VNB.n66 VNB.n63 4.305
R454 VNB.n172 VNB.n169 3.947
R455 VNB.n74 VNB.n73 3.947
R456 VNB.n144 VNB.n141 2.511
R457 VNB.n51 VNB.n46 2.511
R458 VNB.t2 VNB.n5 2.238
R459 VNB.n49 VNB.n47 1.99
R460 VNB.n222 VNB.n213 0.921
R461 VNB.n222 VNB.n217 0.476
R462 VNB.n222 VNB.n212 0.475
R463 VNB.n112 VNB.n111 0.358
R464 VNB.n11 VNB.n10 0.358
R465 VNB.n177 VNB.n176 0.272
R466 VNB.n204 VNB.n203 0.272
R467 VNB.n104 VNB.n98 0.246
R468 VNB.n105 VNB.n104 0.246
R469 VNB.n104 VNB.n103 0.246
R470 VNB.n87 VNB.n81 0.246
R471 VNB.n88 VNB.n87 0.246
R472 VNB.n87 VNB.n86 0.246
R473 VNB.n27 VNB.n21 0.246
R474 VNB.n28 VNB.n27 0.246
R475 VNB.n27 VNB.n26 0.246
R476 VNB.n159 VNB.n154 0.246
R477 VNB.n160 VNB.n159 0.246
R478 VNB.n159 VNB.n158 0.246
R479 VNB.n222 VNB.n221 0.246
R480 VNB.n208 VNB 0.198
R481 VNB.n116 VNB.n115 0.179
R482 VNB.n70 VNB.n67 0.179
R483 VNB.n174 VNB.n173 0.136
R484 VNB.n175 VNB.n174 0.136
R485 VNB.n176 VNB.n175 0.136
R486 VNB.n178 VNB.n177 0.136
R487 VNB.n179 VNB.n178 0.136
R488 VNB.n180 VNB.n179 0.136
R489 VNB.n181 VNB.n180 0.136
R490 VNB.n182 VNB.n181 0.136
R491 VNB.n183 VNB.n182 0.136
R492 VNB.n184 VNB.n183 0.136
R493 VNB.n184 VNB 0.136
R494 VNB.n193 VNB 0.136
R495 VNB.n197 VNB.n193 0.136
R496 VNB.n198 VNB.n197 0.136
R497 VNB.n199 VNB.n198 0.136
R498 VNB.n200 VNB.n199 0.136
R499 VNB.n201 VNB.n200 0.136
R500 VNB.n202 VNB.n201 0.136
R501 VNB.n203 VNB.n202 0.136
R502 VNB.n205 VNB.n204 0.136
R503 VNB.n206 VNB.n205 0.136
R504 VNB.n207 VNB.n206 0.136
R505 VNB.n208 VNB.n207 0.136
R506 a_556_74.t0 a_556_74.n1 34.62
R507 a_556_74.t0 a_556_74.n0 8.137
R508 a_556_74.t0 a_556_74.n2 4.69
C6 VPB VNB 9.68fF
C7 a_556_74.n0 VNB 0.05fF
C8 a_556_74.n1 VNB 0.12fF
C9 a_556_74.n2 VNB 0.04fF
C10 a_1222_74.n0 VNB 0.05fF
C11 a_1222_74.n1 VNB 0.02fF
C12 a_1222_74.n2 VNB 0.12fF
C13 a_1222_74.n3 VNB 0.04fF
C14 a_1222_74.n4 VNB 0.17fF
C15 a_185_182.n0 VNB 0.05fF
C16 a_185_182.n1 VNB 0.99fF
C17 a_185_182.n2 VNB 0.56fF
C18 a_185_182.n3 VNB 1.14fF
C19 a_185_182.n4 VNB 1.21fF
C20 a_185_182.n5 VNB 0.04fF
C21 a_185_182.n6 VNB 0.25fF
C22 a_185_182.n7 VNB 0.07fF
C23 a_1241_1004.n0 VNB 0.52fF
C24 VPB.n0 VNB 0.03fF
C25 VPB.n1 VNB 0.04fF
C26 VPB.n2 VNB 0.02fF
C27 VPB.n3 VNB 0.10fF
C28 VPB.n5 VNB 0.02fF
C29 VPB.n6 VNB 0.02fF
C30 VPB.n7 VNB 0.02fF
C31 VPB.n8 VNB 0.02fF
C32 VPB.n10 VNB 0.02fF
C33 VPB.n11 VNB 0.02fF
C34 VPB.n12 VNB 0.02fF
C35 VPB.n14 VNB 0.02fF
C36 VPB.n15 VNB 0.02fF
C37 VPB.n16 VNB 0.02fF
C38 VPB.n17 VNB 0.04fF
C39 VPB.n18 VNB 0.02fF
C40 VPB.n19 VNB 0.17fF
C41 VPB.n20 VNB 0.04fF
C42 VPB.n22 VNB 0.02fF
C43 VPB.n23 VNB 0.02fF
C44 VPB.n24 VNB 0.02fF
C45 VPB.n25 VNB 0.02fF
C46 VPB.n27 VNB 0.02fF
C47 VPB.n28 VNB 0.02fF
C48 VPB.n29 VNB 0.02fF
C49 VPB.n31 VNB 0.27fF
C50 VPB.n33 VNB 0.03fF
C51 VPB.n34 VNB 0.02fF
C52 VPB.n35 VNB 0.09fF
C53 VPB.n36 VNB 0.27fF
C54 VPB.n37 VNB 0.02fF
C55 VPB.n38 VNB 0.02fF
C56 VPB.n39 VNB 0.27fF
C57 VPB.n40 VNB 0.02fF
C58 VPB.n41 VNB 0.02fF
C59 VPB.n42 VNB 0.13fF
C60 VPB.n43 VNB 0.15fF
C61 VPB.n44 VNB 0.02fF
C62 VPB.n45 VNB 0.02fF
C63 VPB.n46 VNB 0.03fF
C64 VPB.n47 VNB 0.13fF
C65 VPB.n48 VNB 0.16fF
C66 VPB.n49 VNB 0.02fF
C67 VPB.n50 VNB 0.02fF
C68 VPB.n51 VNB 0.23fF
C69 VPB.n52 VNB 0.02fF
C70 VPB.n53 VNB 0.02fF
C71 VPB.n54 VNB 0.27fF
C72 VPB.n55 VNB 0.01fF
C73 VPB.n56 VNB 0.02fF
C74 VPB.n57 VNB 0.03fF
C75 VPB.n58 VNB 0.03fF
C76 VPB.n59 VNB 0.27fF
C77 VPB.n60 VNB 0.01fF
C78 VPB.n61 VNB 0.02fF
C79 VPB.n62 VNB 0.06fF
C80 VPB.n63 VNB 0.13fF
C81 VPB.n64 VNB 0.19fF
C82 VPB.n65 VNB 0.02fF
C83 VPB.n66 VNB 0.01fF
C84 VPB.n67 VNB 0.16fF
C85 VPB.n68 VNB 0.02fF
C86 VPB.n69 VNB 0.02fF
C87 VPB.n70 VNB 0.13fF
C88 VPB.n71 VNB 0.19fF
C89 VPB.n72 VNB 0.02fF
C90 VPB.n73 VNB 0.01fF
C91 VPB.n74 VNB 0.06fF
C92 VPB.n75 VNB 0.02fF
C93 VPB.n76 VNB 0.02fF
C94 VPB.n77 VNB 0.02fF
C95 VPB.n78 VNB 0.04fF
C96 VPB.n79 VNB 0.02fF
C97 VPB.n80 VNB 0.19fF
C98 VPB.n81 VNB 0.04fF
C99 VPB.n83 VNB 0.02fF
C100 VPB.n84 VNB 0.02fF
C101 VPB.n85 VNB 0.02fF
C102 VPB.n86 VNB 0.02fF
C103 VPB.n88 VNB 0.02fF
C104 VPB.n89 VNB 0.02fF
C105 VPB.n90 VNB 0.02fF
C106 VPB.n92 VNB 0.27fF
C107 VPB.n94 VNB 0.03fF
C108 VPB.n95 VNB 0.02fF
C109 VPB.n96 VNB 0.09fF
C110 VPB.n97 VNB 0.02fF
C111 VPB.n98 VNB 0.02fF
C112 VPB.n99 VNB 0.02fF
C113 VPB.n100 VNB 0.04fF
C114 VPB.n101 VNB 0.02fF
C115 VPB.n102 VNB 0.17fF
C116 VPB.n103 VNB 0.04fF
C117 VPB.n105 VNB 0.02fF
C118 VPB.n106 VNB 0.02fF
C119 VPB.n107 VNB 0.02fF
C120 VPB.n108 VNB 0.02fF
C121 VPB.n110 VNB 0.02fF
C122 VPB.n111 VNB 0.02fF
C123 VPB.n112 VNB 0.02fF
C124 VPB.n114 VNB 0.27fF
C125 VPB.n116 VNB 0.03fF
C126 VPB.n117 VNB 0.02fF
C127 VPB.n118 VNB 0.16fF
C128 VPB.n119 VNB 0.02fF
C129 VPB.n120 VNB 0.02fF
C130 VPB.n121 VNB 0.13fF
C131 VPB.n122 VNB 0.19fF
C132 VPB.n123 VNB 0.02fF
C133 VPB.n124 VNB 0.01fF
C134 VPB.n125 VNB 0.06fF
C135 VPB.n126 VNB 0.27fF
C136 VPB.n127 VNB 0.01fF
C137 VPB.n128 VNB 0.02fF
C138 VPB.n129 VNB 0.03fF
C139 VPB.n130 VNB 0.03fF
C140 VPB.n131 VNB 0.27fF
C141 VPB.n132 VNB 0.01fF
C142 VPB.n133 VNB 0.02fF
C143 VPB.n134 VNB 0.27fF
C144 VPB.n135 VNB 0.02fF
C145 VPB.n136 VNB 0.02fF
C146 VPB.n137 VNB 0.27fF
C147 VPB.n138 VNB 0.02fF
C148 VPB.n139 VNB 0.02fF
C149 VPB.n140 VNB 0.27fF
C150 VPB.n141 VNB 0.02fF
C151 VPB.n142 VNB 0.02fF
C152 VPB.n143 VNB 0.13fF
C153 VPB.n144 VNB 0.15fF
C154 VPB.n145 VNB 0.02fF
C155 VPB.n146 VNB 0.02fF
C156 VPB.n147 VNB 0.03fF
C157 VPB.n148 VNB 0.13fF
C158 VPB.n149 VNB 0.16fF
C159 VPB.n150 VNB 0.02fF
C160 VPB.n151 VNB 0.02fF
C161 VPB.n152 VNB 0.23fF
C162 VPB.n153 VNB 0.02fF
C163 VPB.n154 VNB 0.02fF
C164 VPB.n155 VNB 0.02fF
C165 VPB.n156 VNB 0.02fF
C166 VPB.n157 VNB 0.02fF
C167 VPB.n158 VNB 0.10fF
C168 VPB.n159 VNB 0.03fF
C169 VPB.n160 VNB 0.02fF
C170 VPB.n161 VNB 0.05fF
C171 VPB.n162 VNB 0.01fF
C172 VPB.n163 VNB 0.02fF
C173 VPB.n164 VNB 0.02fF
C174 VPB.n166 VNB 0.02fF
C175 VPB.n167 VNB 0.02fF
C176 VPB.n170 VNB 0.02fF
C177 VPB.n172 VNB 0.45fF
C178 VPB.n174 VNB 0.04fF
C179 VPB.n175 VNB 0.04fF
C180 VPB.n176 VNB 0.27fF
C181 VPB.n177 VNB 0.03fF
C182 VPB.n178 VNB 0.03fF
C183 VPB.n179 VNB 0.06fF
C184 VPB.n180 VNB 0.13fF
C185 VPB.n181 VNB 0.19fF
C186 VPB.n182 VNB 0.02fF
C187 VPB.n183 VNB 0.01fF
C188 VPB.n184 VNB 0.07fF
C189 VPB.n185 VNB 0.02fF
C190 VPB.n186 VNB 0.02fF
C191 VPB.n187 VNB 0.04fF
C192 VPB.n188 VNB 0.04fF
C193 VPB.n189 VNB 0.02fF
C194 VPB.n190 VNB 0.02fF
C195 VPB.n191 VNB 0.02fF
C196 VPB.n192 VNB 0.02fF
C197 VPB.n193 VNB 0.02fF
C198 VPB.n194 VNB 0.02fF
C199 VPB.n195 VNB 0.02fF
C200 VPB.n196 VNB 0.27fF
C201 VPB.n197 VNB 0.01fF
C202 VPB.n198 VNB 0.02fF
C203 VPB.n199 VNB 0.03fF
C204 VPB.n200 VNB 0.03fF
C205 VPB.n201 VNB 0.27fF
C206 VPB.n202 VNB 0.01fF
C207 VPB.n203 VNB 0.02fF
C208 VPB.n204 VNB 0.02fF
C209 VPB.n205 VNB 0.27fF
C210 VPB.n206 VNB 0.02fF
C211 VPB.n207 VNB 0.02fF
C212 VPB.n208 VNB 0.02fF
C213 VPB.n209 VNB 0.02fF
C214 VPB.n210 VNB 0.02fF
C215 VPB.n211 VNB 0.02fF
C216 VPB.n212 VNB 0.02fF
C217 VPB.n213 VNB 0.02fF
C218 VPB.n214 VNB 0.04fF
C219 VPB.n215 VNB 0.04fF
C220 VPB.n216 VNB 0.02fF
C221 VPB.n217 VNB 0.02fF
C222 VPB.n218 VNB 0.02fF
C223 VPB.n219 VNB 0.03fF
C224 VPB.n220 VNB 0.03fF
C225 VPB.n221 VNB 0.02fF
C226 VPB.n222 VNB 0.02fF
C227 VPB.n223 VNB 0.02fF
C228 VPB.n224 VNB 0.04fF
C229 VPB.n225 VNB 0.04fF
C230 VPB.n227 VNB 0.42fF
C231 a_575_1004.n0 VNB 0.52fF
C232 a_807_943.n0 VNB 0.06fF
C233 a_807_943.n1 VNB 1.05fF
C234 a_807_943.n2 VNB 1.14fF
C235 a_807_943.n3 VNB 1.26fF
C236 a_807_943.n4 VNB 1.43fF
C237 a_807_943.n5 VNB 0.05fF
C238 a_807_943.n6 VNB 0.42fF
C239 a_807_943.n7 VNB 0.08fF
.ends
