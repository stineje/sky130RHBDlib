* SPICE3 file created from AND3X1.ext - technology: sky130A

.subckt AND3X1 Y A B C VDD GND
X0 Y and3x1_pcell_0/m1_867_649# GND GND nshort w=3 l=0.15
X1 VDD and3x1_pcell_0/m1_867_649# Y VDD pshort w=2 l=0.15
X2 GND A and3x1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X3 and3x1_pcell_0/m1_867_649# C and3x1_pcell_0/nand3x1_pcell_0/li_393_182# GND nshort w=3 l=0.15
X4 and3x1_pcell_0/nand3x1_pcell_0/li_393_182# B and3x1_pcell_0/nand3x1_pcell_0/nmos_bottom_0/a_0_0# GND nshort w=3 l=0.15
X5 VDD A and3x1_pcell_0/m1_867_649# VDD pshort w=2 l=0.15
X6 VDD B and3x1_pcell_0/m1_867_649# VDD pshort w=2 l=0.15
X7 VDD C and3x1_pcell_0/m1_867_649# VDD pshort w=2 l=0.15
C0 VDD GND 5.50fF
.ends
