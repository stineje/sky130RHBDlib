magic
tech sky130A
magscale 1 2
timestamp 1652323096
<< metal1 >>
rect 547 649 761 683
use nand2x1_pcell  nand2x1_pcell_0
timestamp 1652323009
transform 1 0 0 0 1 0
box -87 -34 753 1550
use invx1_pcell  invx1_pcell_0
timestamp 1652321374
transform 1 0 666 0 1 0
box -87 -34 531 1550
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 814 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 518 0 -1 666
box -53 -33 29 33
<< end >>
