// File: DFFRNX1.spi.pex
// Created: Tue Oct 15 15:46:41 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_DFFRNX1\%GND ( 1 47 51 54 59 69 77 87 95 103 109 119 125 135 146 150 \
 152 154 157 160 163 164 165 166 167 168 )
c292 ( 168 0 ) capacitor c=0.0208017f //x=23.56 //y=0.865
c293 ( 167 0 ) capacitor c=0.0225954f //x=18.645 //y=0.875
c294 ( 166 0 ) capacitor c=0.0226075f //x=13.835 //y=0.875
c295 ( 165 0 ) capacitor c=0.0207407f //x=10.61 //y=0.865
c296 ( 164 0 ) capacitor c=0.0226571f //x=5.695 //y=0.875
c297 ( 163 0 ) capacitor c=0.022675f //x=0.885 //y=0.875
c298 ( 162 0 ) capacitor c=0.00440095f //x=23.68 //y=0
c299 ( 160 0 ) capacitor c=0.109815f //x=22.57 //y=0
c300 ( 159 0 ) capacitor c=0.00440144f //x=18.87 //y=0
c301 ( 157 0 ) capacitor c=0.107954f //x=17.76 //y=0
c302 ( 156 0 ) capacitor c=0.00440144f //x=14.06 //y=0
c303 ( 154 0 ) capacitor c=0.10465f //x=12.95 //y=0
c304 ( 153 0 ) capacitor c=0.00440095f //x=10.8 //y=0
c305 ( 152 0 ) capacitor c=0.108705f //x=9.62 //y=0
c306 ( 151 0 ) capacitor c=0.00440144f //x=5.885 //y=0
c307 ( 150 0 ) capacitor c=0.10869f //x=4.81 //y=0
c308 ( 149 0 ) capacitor c=0.00440144f //x=1.075 //y=0
c309 ( 146 0 ) capacitor c=0.259877f //x=25.53 //y=0
c310 ( 135 0 ) capacitor c=0.0389288f //x=23.665 //y=0
c311 ( 125 0 ) capacitor c=0.131607f //x=22.4 //y=0
c312 ( 119 0 ) capacitor c=0.0339325f //x=18.75 //y=0
c313 ( 109 0 ) capacitor c=0.133561f //x=17.59 //y=0
c314 ( 103 0 ) capacitor c=0.0339325f //x=13.94 //y=0
c315 ( 95 0 ) capacitor c=0.0718026f //x=12.78 //y=0
c316 ( 87 0 ) capacitor c=0.0388888f //x=10.715 //y=0
c317 ( 77 0 ) capacitor c=0.133699f //x=9.45 //y=0
c318 ( 69 0 ) capacitor c=0.0339738f //x=5.8 //y=0
c319 ( 59 0 ) capacitor c=0.131745f //x=4.64 //y=0
c320 ( 54 0 ) capacitor c=0.178285f //x=0.74 //y=0
c321 ( 51 0 ) capacitor c=0.0367385f //x=0.99 //y=0
c322 ( 47 0 ) capacitor c=0.816614f //x=25.53 //y=0
r323 (  144 146 ) resistor r=26.5322 //w=0.357 //l=0.74 //layer=li \
 //thickness=0.1 //x=24.79 //y=0 //x2=25.53 //y2=0
r324 (  142 162 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.835 //y=0 //x2=23.75 //y2=0
r325 (  142 144 ) resistor r=34.2409 //w=0.357 //l=0.955 //layer=li \
 //thickness=0.1 //x=23.835 //y=0 //x2=24.79 //y2=0
r326 (  137 162 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.75 //y=0.17 //x2=23.75 //y2=0
r327 (  137 168 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=23.75 //y=0.17 //x2=23.75 //y2=0.955
r328 (  136 160 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.74 //y=0 //x2=22.57 //y2=0
r329 (  135 162 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.665 //y=0 //x2=23.75 //y2=0
r330 (  135 136 ) resistor r=33.1653 //w=0.357 //l=0.925 //layer=li \
 //thickness=0.1 //x=23.665 //y=0 //x2=22.74 //y2=0
r331 (  130 132 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=21.09 //y=0 //x2=22.2 //y2=0
r332 (  128 130 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=19.98 //y=0 //x2=21.09 //y2=0
r333 (  126 159 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.92 //y=0 //x2=18.835 //y2=0
r334 (  126 128 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=18.92 //y=0 //x2=19.98 //y2=0
r335 (  125 160 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.4 //y=0 //x2=22.57 //y2=0
r336 (  125 132 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=22.4 //y=0 //x2=22.2 //y2=0
r337 (  121 159 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.835 //y=0.17 //x2=18.835 //y2=0
r338 (  121 167 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=18.835 //y=0.17 //x2=18.835 //y2=0.965
r339 (  120 157 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.93 //y=0 //x2=17.76 //y2=0
r340 (  119 159 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.75 //y=0 //x2=18.835 //y2=0
r341 (  119 120 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=18.75 //y=0 //x2=17.93 //y2=0
r342 (  114 116 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=16.28 //y=0 //x2=17.39 //y2=0
r343 (  112 114 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=15.17 //y=0 //x2=16.28 //y2=0
r344 (  110 156 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.11 //y=0 //x2=14.025 //y2=0
r345 (  110 112 ) resistor r=38.0056 //w=0.357 //l=1.06 //layer=li \
 //thickness=0.1 //x=14.11 //y=0 //x2=15.17 //y2=0
r346 (  109 157 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.59 //y=0 //x2=17.76 //y2=0
r347 (  109 116 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=17.59 //y=0 //x2=17.39 //y2=0
r348 (  105 156 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.025 //y=0.17 //x2=14.025 //y2=0
r349 (  105 166 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=14.025 //y=0.17 //x2=14.025 //y2=0.965
r350 (  104 154 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.12 //y=0 //x2=12.95 //y2=0
r351 (  103 156 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.94 //y=0 //x2=14.025 //y2=0
r352 (  103 104 ) resistor r=29.4006 //w=0.357 //l=0.82 //layer=li \
 //thickness=0.1 //x=13.94 //y=0 //x2=13.12 //y2=0
r353 (  98 100 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=11.47 //y=0 //x2=12.58 //y2=0
r354 (  96 153 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.885 //y=0 //x2=10.8 //y2=0
r355 (  96 98 ) resistor r=20.9748 //w=0.357 //l=0.585 //layer=li \
 //thickness=0.1 //x=10.885 //y=0 //x2=11.47 //y2=0
r356 (  95 154 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.78 //y=0 //x2=12.95 //y2=0
r357 (  95 100 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.78 //y=0 //x2=12.58 //y2=0
r358 (  91 153 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.8 //y=0.17 //x2=10.8 //y2=0
r359 (  91 165 ) resistor r=53.7326 //w=0.187 //l=0.785 //layer=li \
 //thickness=0.1 //x=10.8 //y=0.17 //x2=10.8 //y2=0.955
r360 (  88 152 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.79 //y=0 //x2=9.62 //y2=0
r361 (  88 90 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.79 //y=0 //x2=10.36 //y2=0
r362 (  87 153 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.715 //y=0 //x2=10.8 //y2=0
r363 (  87 90 ) resistor r=12.7283 //w=0.357 //l=0.355 //layer=li \
 //thickness=0.1 //x=10.715 //y=0 //x2=10.36 //y2=0
r364 (  82 84 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=7.77 //y=0 //x2=8.88 //y2=0
r365 (  80 82 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=6.66 //y=0 //x2=7.77 //y2=0
r366 (  78 151 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.97 //y=0 //x2=5.885 //y2=0
r367 (  78 80 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=5.97 //y=0 //x2=6.66 //y2=0
r368 (  77 152 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.45 //y=0 //x2=9.62 //y2=0
r369 (  77 84 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.45 //y=0 //x2=8.88 //y2=0
r370 (  73 151 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.885 //y=0.17 //x2=5.885 //y2=0
r371 (  73 164 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=5.885 //y=0.17 //x2=5.885 //y2=0.965
r372 (  70 150 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=4.81 //y2=0
r373 (  70 72 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=0 //x2=5.55 //y2=0
r374 (  69 151 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.8 //y=0 //x2=5.885 //y2=0
r375 (  69 72 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=5.8 //y=0 //x2=5.55 //y2=0
r376 (  64 66 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=0 //x2=4.07 //y2=0
r377 (  62 64 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r378 (  60 149 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.075 //y2=0
r379 (  60 62 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.85 //y2=0
r380 (  59 150 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.81 //y2=0
r381 (  59 66 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.07 //y2=0
r382 (  55 149 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0
r383 (  55 163 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0.965
r384 (  51 149 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=1.075 //y2=0
r385 (  51 54 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=0.74 //y2=0
r386 (  47 146 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=25.53 //y=0 //x2=25.53 //y2=0
r387 (  45 144 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=0 //x2=24.79 //y2=0
r388 (  45 47 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=0 //x2=25.53 //y2=0
r389 (  43 162 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=0 //x2=23.68 //y2=0
r390 (  43 45 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=23.68 //y=0 //x2=24.79 //y2=0
r391 (  41 132 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.2 //y=0 //x2=22.2 //y2=0
r392 (  41 43 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=22.2 //y=0 //x2=23.68 //y2=0
r393 (  39 130 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=0 //x2=21.09 //y2=0
r394 (  39 41 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=0 //x2=22.2 //y2=0
r395 (  37 128 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=0 //x2=19.98 //y2=0
r396 (  37 39 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=0 //x2=21.09 //y2=0
r397 (  35 159 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.87 //y=0 //x2=18.87 //y2=0
r398 (  35 37 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=18.87 //y=0 //x2=19.98 //y2=0
r399 (  33 116 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=0 //x2=17.39 //y2=0
r400 (  33 35 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=0 //x2=18.87 //y2=0
r401 (  31 114 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=0 //x2=16.28 //y2=0
r402 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=0 //x2=17.39 //y2=0
r403 (  29 112 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=0 //x2=15.17 //y2=0
r404 (  29 31 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=0 //x2=16.28 //y2=0
r405 (  27 156 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=0 //x2=14.06 //y2=0
r406 (  27 29 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=0 //x2=15.17 //y2=0
r407 (  24 100 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=0 //x2=12.58 //y2=0
r408 (  22 98 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=0 //x2=11.47 //y2=0
r409 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=0 //x2=12.58 //y2=0
r410 (  20 90 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=0 //x2=10.36 //y2=0
r411 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=0 //x2=11.47 //y2=0
r412 (  18 84 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.88 //y=0 //x2=8.88 //y2=0
r413 (  18 20 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.88 //y=0 //x2=10.36 //y2=0
r414 (  16 82 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=0 //x2=7.77 //y2=0
r415 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=0 //x2=8.88 //y2=0
r416 (  14 80 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=0 //x2=6.66 //y2=0
r417 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=0 //x2=7.77 //y2=0
r418 (  12 72 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r419 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.66 //y2=0
r420 (  10 66 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r421 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=0 //x2=5.55 //y2=0
r422 (  8 64 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r423 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.07 //y2=0
r424 (  6 62 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r425 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r426 (  3 54 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r427 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r428 (  1 27 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.95 //y=0 //x2=14.06 //y2=0
r429 (  1 24 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=12.95 //y=0 //x2=12.58 //y2=0
ends PM_DFFRNX1\%GND

subckt PM_DFFRNX1\%VDD ( 1 47 54 61 71 79 89 95 105 115 123 133 139 147 155 \
 165 171 179 187 197 207 213 221 229 239 249 255 263 273 286 293 298 303 309 \
 315 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 \
 337 338 339 340 )
c323 ( 340 0 ) capacitor c=0.0382077f //x=24.975 //y=5.02
c324 ( 339 0 ) capacitor c=0.0240874f //x=24.095 //y=5.02
c325 ( 338 0 ) capacitor c=0.0495444f //x=23.225 //y=5.02
c326 ( 337 0 ) capacitor c=0.0453059f //x=21.345 //y=5.02
c327 ( 336 0 ) capacitor c=0.02424f //x=20.465 //y=5.02
c328 ( 335 0 ) capacitor c=0.02424f //x=19.585 //y=5.02
c329 ( 334 0 ) capacitor c=0.0531793f //x=18.715 //y=5.02
c330 ( 333 0 ) capacitor c=0.0453059f //x=16.535 //y=5.02
c331 ( 332 0 ) capacitor c=0.02424f //x=15.655 //y=5.02
c332 ( 331 0 ) capacitor c=0.024152f //x=14.775 //y=5.02
c333 ( 330 0 ) capacitor c=0.0531894f //x=13.905 //y=5.02
c334 ( 329 0 ) capacitor c=0.0380679f //x=12.025 //y=5.02
c335 ( 328 0 ) capacitor c=0.024008f //x=11.145 //y=5.02
c336 ( 327 0 ) capacitor c=0.049209f //x=10.275 //y=5.02
c337 ( 326 0 ) capacitor c=0.0452179f //x=8.395 //y=5.02
c338 ( 325 0 ) capacitor c=0.024152f //x=7.515 //y=5.02
c339 ( 324 0 ) capacitor c=0.024152f //x=6.635 //y=5.02
c340 ( 323 0 ) capacitor c=0.053132f //x=5.765 //y=5.02
c341 ( 322 0 ) capacitor c=0.0452179f //x=3.585 //y=5.02
c342 ( 321 0 ) capacitor c=0.024152f //x=2.705 //y=5.02
c343 ( 320 0 ) capacitor c=0.02424f //x=1.825 //y=5.02
c344 ( 319 0 ) capacitor c=0.0531407f //x=0.955 //y=5.02
c345 ( 318 0 ) capacitor c=0.00591168f //x=25.12 //y=7.4
c346 ( 317 0 ) capacitor c=0.00591168f //x=24.24 //y=7.4
c347 ( 316 0 ) capacitor c=0.00591168f //x=23.36 //y=7.4
c348 ( 315 0 ) capacitor c=0.136751f //x=22.57 //y=7.4
c349 ( 314 0 ) capacitor c=0.00591168f //x=21.49 //y=7.4
c350 ( 313 0 ) capacitor c=0.00591168f //x=20.61 //y=7.4
c351 ( 312 0 ) capacitor c=0.00591168f //x=19.73 //y=7.4
c352 ( 311 0 ) capacitor c=0.00591168f //x=18.87 //y=7.4
c353 ( 309 0 ) capacitor c=0.15714f //x=17.76 //y=7.4
c354 ( 308 0 ) capacitor c=0.00591168f //x=16.68 //y=7.4
c355 ( 307 0 ) capacitor c=0.00591168f //x=15.8 //y=7.4
c356 ( 306 0 ) capacitor c=0.00591168f //x=14.92 //y=7.4
c357 ( 305 0 ) capacitor c=0.00591168f //x=14.06 //y=7.4
c358 ( 303 0 ) capacitor c=0.135038f //x=12.95 //y=7.4
c359 ( 302 0 ) capacitor c=0.00591168f //x=12.17 //y=7.4
c360 ( 301 0 ) capacitor c=0.00591168f //x=11.29 //y=7.4
c361 ( 300 0 ) capacitor c=0.00591168f //x=10.36 //y=7.4
c362 ( 298 0 ) capacitor c=0.134558f //x=9.62 //y=7.4
c363 ( 297 0 ) capacitor c=0.00591168f //x=8.54 //y=7.4
c364 ( 296 0 ) capacitor c=0.00591168f //x=7.66 //y=7.4
c365 ( 295 0 ) capacitor c=0.00591168f //x=6.78 //y=7.4
c366 ( 294 0 ) capacitor c=0.00591168f //x=5.9 //y=7.4
c367 ( 293 0 ) capacitor c=0.15519f //x=4.81 //y=7.4
c368 ( 292 0 ) capacitor c=0.00591168f //x=3.73 //y=7.4
c369 ( 291 0 ) capacitor c=0.00591168f //x=2.85 //y=7.4
c370 ( 290 0 ) capacitor c=0.00591168f //x=1.97 //y=7.4
c371 ( 289 0 ) capacitor c=0.00591168f //x=1.09 //y=7.4
c372 ( 286 0 ) capacitor c=0.237727f //x=25.53 //y=7.4
c373 ( 273 0 ) capacitor c=0.0284327f //x=25.035 //y=7.4
c374 ( 263 0 ) capacitor c=0.0288633f //x=24.155 //y=7.4
c375 ( 255 0 ) capacitor c=0.0240981f //x=23.275 //y=7.4
c376 ( 249 0 ) capacitor c=0.0395236f //x=22.4 //y=7.4
c377 ( 239 0 ) capacitor c=0.0288769f //x=21.405 //y=7.4
c378 ( 229 0 ) capacitor c=0.0287757f //x=20.525 //y=7.4
c379 ( 221 0 ) capacitor c=0.028511f //x=19.645 //y=7.4
c380 ( 213 0 ) capacitor c=0.0383672f //x=18.765 //y=7.4
c381 ( 207 0 ) capacitor c=0.0395206f //x=17.59 //y=7.4
c382 ( 197 0 ) capacitor c=0.0288769f //x=16.595 //y=7.4
c383 ( 187 0 ) capacitor c=0.0287624f //x=15.715 //y=7.4
c384 ( 179 0 ) capacitor c=0.0284966f //x=14.835 //y=7.4
c385 ( 171 0 ) capacitor c=0.0383672f //x=13.955 //y=7.4
c386 ( 165 0 ) capacitor c=0.0236224f //x=12.78 //y=7.4
c387 ( 155 0 ) capacitor c=0.0288359f //x=12.085 //y=7.4
c388 ( 147 0 ) capacitor c=0.0288369f //x=11.205 //y=7.4
c389 ( 139 0 ) capacitor c=0.0240981f //x=10.325 //y=7.4
c390 ( 133 0 ) capacitor c=0.0394667f //x=9.45 //y=7.4
c391 ( 123 0 ) capacitor c=0.0288488f //x=8.455 //y=7.4
c392 ( 115 0 ) capacitor c=0.0287514f //x=7.575 //y=7.4
c393 ( 105 0 ) capacitor c=0.0284966f //x=6.695 //y=7.4
c394 ( 95 0 ) capacitor c=0.0383672f //x=5.815 //y=7.4
c395 ( 89 0 ) capacitor c=0.0394667f //x=4.64 //y=7.4
c396 ( 79 0 ) capacitor c=0.0288488f //x=3.645 //y=7.4
c397 ( 71 0 ) capacitor c=0.0287505f //x=2.765 //y=7.4
c398 ( 61 0 ) capacitor c=0.028511f //x=1.885 //y=7.4
c399 ( 54 0 ) capacitor c=0.234426f //x=0.74 //y=7.4
c400 ( 51 0 ) capacitor c=0.0452081f //x=1.005 //y=7.4
c401 ( 47 0 ) capacitor c=0.899931f //x=25.53 //y=7.4
r402 (  284 318 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.205 //y=7.4 //x2=25.12 //y2=7.4
r403 (  284 286 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=25.205 //y=7.4 //x2=25.53 //y2=7.4
r404 (  277 318 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=25.12 //y=7.23 //x2=25.12 //y2=7.4
r405 (  277 340 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=25.12 //y=7.23 //x2=25.12 //y2=6.745
r406 (  274 317 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.325 //y=7.4 //x2=24.24 //y2=7.4
r407 (  274 276 ) resistor r=16.6723 //w=0.357 //l=0.465 //layer=li \
 //thickness=0.1 //x=24.325 //y=7.4 //x2=24.79 //y2=7.4
r408 (  273 318 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=25.035 //y=7.4 //x2=25.12 //y2=7.4
r409 (  273 276 ) resistor r=8.78431 //w=0.357 //l=0.245 //layer=li \
 //thickness=0.1 //x=25.035 //y=7.4 //x2=24.79 //y2=7.4
r410 (  267 317 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=24.24 //y=7.23 //x2=24.24 //y2=7.4
r411 (  267 339 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=24.24 //y=7.23 //x2=24.24 //y2=6.745
r412 (  264 316 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.445 //y=7.4 //x2=23.36 //y2=7.4
r413 (  264 266 ) resistor r=8.42577 //w=0.357 //l=0.235 //layer=li \
 //thickness=0.1 //x=23.445 //y=7.4 //x2=23.68 //y2=7.4
r414 (  263 317 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.155 //y=7.4 //x2=24.24 //y2=7.4
r415 (  263 266 ) resistor r=17.0308 //w=0.357 //l=0.475 //layer=li \
 //thickness=0.1 //x=24.155 //y=7.4 //x2=23.68 //y2=7.4
r416 (  257 316 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=23.36 //y=7.23 //x2=23.36 //y2=7.4
r417 (  257 338 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=23.36 //y=7.23 //x2=23.36 //y2=6.405
r418 (  256 315 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.74 //y=7.4 //x2=22.57 //y2=7.4
r419 (  255 316 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=23.275 //y=7.4 //x2=23.36 //y2=7.4
r420 (  255 256 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=23.275 //y=7.4 //x2=22.74 //y2=7.4
r421 (  250 314 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.575 //y=7.4 //x2=21.49 //y2=7.4
r422 (  250 252 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=21.575 //y=7.4 //x2=22.2 //y2=7.4
r423 (  249 315 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=22.4 //y=7.4 //x2=22.57 //y2=7.4
r424 (  249 252 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=22.4 //y=7.4 //x2=22.2 //y2=7.4
r425 (  243 314 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=21.49 //y=7.23 //x2=21.49 //y2=7.4
r426 (  243 337 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.49 //y=7.23 //x2=21.49 //y2=6.745
r427 (  240 313 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.695 //y=7.4 //x2=20.61 //y2=7.4
r428 (  240 242 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=20.695 //y=7.4 //x2=21.09 //y2=7.4
r429 (  239 314 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.405 //y=7.4 //x2=21.49 //y2=7.4
r430 (  239 242 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=21.405 //y=7.4 //x2=21.09 //y2=7.4
r431 (  233 313 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=20.61 //y=7.23 //x2=20.61 //y2=7.4
r432 (  233 336 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.61 //y=7.23 //x2=20.61 //y2=6.745
r433 (  230 312 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.815 //y=7.4 //x2=19.73 //y2=7.4
r434 (  230 232 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=19.815 //y=7.4 //x2=19.98 //y2=7.4
r435 (  229 313 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.525 //y=7.4 //x2=20.61 //y2=7.4
r436 (  229 232 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=20.525 //y=7.4 //x2=19.98 //y2=7.4
r437 (  223 312 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=19.73 //y=7.23 //x2=19.73 //y2=7.4
r438 (  223 335 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=19.73 //y=7.23 //x2=19.73 //y2=6.745
r439 (  222 311 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.935 //y=7.4 //x2=18.85 //y2=7.4
r440 (  221 312 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.645 //y=7.4 //x2=19.73 //y2=7.4
r441 (  221 222 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=19.645 //y=7.4 //x2=18.935 //y2=7.4
r442 (  215 311 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=18.85 //y=7.23 //x2=18.85 //y2=7.4
r443 (  215 334 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=18.85 //y=7.23 //x2=18.85 //y2=6.405
r444 (  214 309 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.93 //y=7.4 //x2=17.76 //y2=7.4
r445 (  213 311 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=18.765 //y=7.4 //x2=18.85 //y2=7.4
r446 (  213 214 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=18.765 //y=7.4 //x2=17.93 //y2=7.4
r447 (  208 308 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.765 //y=7.4 //x2=16.68 //y2=7.4
r448 (  208 210 ) resistor r=22.409 //w=0.357 //l=0.625 //layer=li \
 //thickness=0.1 //x=16.765 //y=7.4 //x2=17.39 //y2=7.4
r449 (  207 309 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=17.59 //y=7.4 //x2=17.76 //y2=7.4
r450 (  207 210 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=17.59 //y=7.4 //x2=17.39 //y2=7.4
r451 (  201 308 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=16.68 //y=7.23 //x2=16.68 //y2=7.4
r452 (  201 333 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.68 //y=7.23 //x2=16.68 //y2=6.745
r453 (  198 307 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.885 //y=7.4 //x2=15.8 //y2=7.4
r454 (  198 200 ) resistor r=14.1625 //w=0.357 //l=0.395 //layer=li \
 //thickness=0.1 //x=15.885 //y=7.4 //x2=16.28 //y2=7.4
r455 (  197 308 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.595 //y=7.4 //x2=16.68 //y2=7.4
r456 (  197 200 ) resistor r=11.2941 //w=0.357 //l=0.315 //layer=li \
 //thickness=0.1 //x=16.595 //y=7.4 //x2=16.28 //y2=7.4
r457 (  191 307 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=15.8 //y=7.23 //x2=15.8 //y2=7.4
r458 (  191 332 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.8 //y=7.23 //x2=15.8 //y2=6.745
r459 (  188 306 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.005 //y=7.4 //x2=14.92 //y2=7.4
r460 (  188 190 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=15.005 //y=7.4 //x2=15.17 //y2=7.4
r461 (  187 307 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.715 //y=7.4 //x2=15.8 //y2=7.4
r462 (  187 190 ) resistor r=19.5406 //w=0.357 //l=0.545 //layer=li \
 //thickness=0.1 //x=15.715 //y=7.4 //x2=15.17 //y2=7.4
r463 (  181 306 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.92 //y=7.23 //x2=14.92 //y2=7.4
r464 (  181 331 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.92 //y=7.23 //x2=14.92 //y2=6.745
r465 (  180 305 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.125 //y=7.4 //x2=14.04 //y2=7.4
r466 (  179 306 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=14.835 //y=7.4 //x2=14.92 //y2=7.4
r467 (  179 180 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=14.835 //y=7.4 //x2=14.125 //y2=7.4
r468 (  173 305 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=14.04 //y=7.23 //x2=14.04 //y2=7.4
r469 (  173 330 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=14.04 //y=7.23 //x2=14.04 //y2=6.405
r470 (  172 303 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=13.12 //y=7.4 //x2=12.95 //y2=7.4
r471 (  171 305 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=13.955 //y=7.4 //x2=14.04 //y2=7.4
r472 (  171 172 ) resistor r=29.9384 //w=0.357 //l=0.835 //layer=li \
 //thickness=0.1 //x=13.955 //y=7.4 //x2=13.12 //y2=7.4
r473 (  166 302 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.255 //y=7.4 //x2=12.17 //y2=7.4
r474 (  166 168 ) resistor r=11.6527 //w=0.357 //l=0.325 //layer=li \
 //thickness=0.1 //x=12.255 //y=7.4 //x2=12.58 //y2=7.4
r475 (  165 303 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.78 //y=7.4 //x2=12.95 //y2=7.4
r476 (  165 168 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=12.78 //y=7.4 //x2=12.58 //y2=7.4
r477 (  159 302 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=12.17 //y=7.23 //x2=12.17 //y2=7.4
r478 (  159 329 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=12.17 //y=7.23 //x2=12.17 //y2=6.745
r479 (  156 301 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.375 //y=7.4 //x2=11.29 //y2=7.4
r480 (  156 158 ) resistor r=3.40616 //w=0.357 //l=0.095 //layer=li \
 //thickness=0.1 //x=11.375 //y=7.4 //x2=11.47 //y2=7.4
r481 (  155 302 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=12.085 //y=7.4 //x2=12.17 //y2=7.4
r482 (  155 158 ) resistor r=22.0504 //w=0.357 //l=0.615 //layer=li \
 //thickness=0.1 //x=12.085 //y=7.4 //x2=11.47 //y2=7.4
r483 (  149 301 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=11.29 //y=7.23 //x2=11.29 //y2=7.4
r484 (  149 328 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=11.29 //y=7.23 //x2=11.29 //y2=6.745
r485 (  148 300 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.495 //y=7.4 //x2=10.41 //y2=7.4
r486 (  147 301 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.205 //y=7.4 //x2=11.29 //y2=7.4
r487 (  147 148 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.205 //y=7.4 //x2=10.495 //y2=7.4
r488 (  141 300 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=10.41 //y=7.23 //x2=10.41 //y2=7.4
r489 (  141 327 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=10.41 //y=7.23 //x2=10.41 //y2=6.405
r490 (  140 298 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.79 //y=7.4 //x2=9.62 //y2=7.4
r491 (  139 300 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=10.325 //y=7.4 //x2=10.41 //y2=7.4
r492 (  139 140 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=10.325 //y=7.4 //x2=9.79 //y2=7.4
r493 (  134 297 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.625 //y=7.4 //x2=8.54 //y2=7.4
r494 (  134 136 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=8.625 //y=7.4 //x2=8.88 //y2=7.4
r495 (  133 298 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=9.45 //y=7.4 //x2=9.62 //y2=7.4
r496 (  133 136 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=9.45 //y=7.4 //x2=8.88 //y2=7.4
r497 (  127 297 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=8.54 //y=7.23 //x2=8.54 //y2=7.4
r498 (  127 326 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.54 //y=7.23 //x2=8.54 //y2=6.745
r499 (  124 296 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.745 //y=7.4 //x2=7.66 //y2=7.4
r500 (  124 126 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=7.745 //y=7.4 //x2=7.77 //y2=7.4
r501 (  123 297 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.455 //y=7.4 //x2=8.54 //y2=7.4
r502 (  123 126 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=8.455 //y=7.4 //x2=7.77 //y2=7.4
r503 (  117 296 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=7.66 //y=7.23 //x2=7.66 //y2=7.4
r504 (  117 325 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.66 //y=7.23 //x2=7.66 //y2=6.745
r505 (  116 295 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.865 //y=7.4 //x2=6.78 //y2=7.4
r506 (  115 296 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.575 //y=7.4 //x2=7.66 //y2=7.4
r507 (  115 116 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.575 //y=7.4 //x2=6.865 //y2=7.4
r508 (  109 295 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=7.4
r509 (  109 324 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.78 //y=7.23 //x2=6.78 //y2=6.745
r510 (  106 294 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.985 //y=7.4 //x2=5.9 //y2=7.4
r511 (  106 108 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=5.985 //y=7.4 //x2=6.66 //y2=7.4
r512 (  105 295 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.78 //y2=7.4
r513 (  105 108 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=6.695 //y=7.4 //x2=6.66 //y2=7.4
r514 (  99 294 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.9 //y=7.23 //x2=5.9 //y2=7.4
r515 (  99 323 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=5.9 //y=7.23 //x2=5.9 //y2=6.405
r516 (  96 293 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=4.81 //y2=7.4
r517 (  96 98 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.98 //y=7.4 //x2=5.55 //y2=7.4
r518 (  95 294 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.815 //y=7.4 //x2=5.9 //y2=7.4
r519 (  95 98 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=5.815 //y=7.4 //x2=5.55 //y2=7.4
r520 (  90 292 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=3.73 //y2=7.4
r521 (  90 92 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=4.07 //y2=7.4
r522 (  89 293 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.81 //y2=7.4
r523 (  89 92 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.07 //y2=7.4
r524 (  83 292 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=7.4
r525 (  83 322 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=6.745
r526 (  80 291 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.85 //y2=7.4
r527 (  80 82 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.96 //y2=7.4
r528 (  79 292 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=3.73 //y2=7.4
r529 (  79 82 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=2.96 //y2=7.4
r530 (  73 291 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=7.4
r531 (  73 321 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=6.745
r532 (  72 290 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.055 //y=7.4 //x2=1.97 //y2=7.4
r533 (  71 291 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.85 //y2=7.4
r534 (  71 72 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.055 //y2=7.4
r535 (  65 290 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=7.4
r536 (  65 320 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=6.745
r537 (  62 289 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.09 //y2=7.4
r538 (  62 64 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.85 //y2=7.4
r539 (  61 290 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.97 //y2=7.4
r540 (  61 64 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.85 //y2=7.4
r541 (  55 289 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=7.4
r542 (  55 319 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=6.405
r543 (  51 289 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=1.09 //y2=7.4
r544 (  51 54 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=0.74 //y2=7.4
r545 (  47 286 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=25.53 //y=7.4 //x2=25.53 //y2=7.4
r546 (  45 276 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=24.79 //y=7.4 //x2=24.79 //y2=7.4
r547 (  45 47 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=24.79 //y=7.4 //x2=25.53 //y2=7.4
r548 (  43 266 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=23.68 //y=7.4 //x2=23.68 //y2=7.4
r549 (  43 45 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=23.68 //y=7.4 //x2=24.79 //y2=7.4
r550 (  41 252 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=22.2 //y=7.4 //x2=22.2 //y2=7.4
r551 (  41 43 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=22.2 //y=7.4 //x2=23.68 //y2=7.4
r552 (  39 242 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=21.09 //y=7.4 //x2=21.09 //y2=7.4
r553 (  39 41 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=21.09 //y=7.4 //x2=22.2 //y2=7.4
r554 (  37 232 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=19.98 //y=7.4 //x2=19.98 //y2=7.4
r555 (  37 39 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=19.98 //y=7.4 //x2=21.09 //y2=7.4
r556 (  35 311 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=18.87 //y=7.4 //x2=18.87 //y2=7.4
r557 (  35 37 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=18.87 //y=7.4 //x2=19.98 //y2=7.4
r558 (  33 210 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=17.39 //y=7.4 //x2=17.39 //y2=7.4
r559 (  33 35 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=17.39 //y=7.4 //x2=18.87 //y2=7.4
r560 (  31 200 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=16.28 //y=7.4 //x2=16.28 //y2=7.4
r561 (  31 33 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=16.28 //y=7.4 //x2=17.39 //y2=7.4
r562 (  29 190 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=15.17 //y=7.4 //x2=15.17 //y2=7.4
r563 (  29 31 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=15.17 //y=7.4 //x2=16.28 //y2=7.4
r564 (  27 305 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=14.06 //y=7.4 //x2=14.06 //y2=7.4
r565 (  27 29 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=14.06 //y=7.4 //x2=15.17 //y2=7.4
r566 (  24 168 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=12.58 //y=7.4 //x2=12.58 //y2=7.4
r567 (  22 158 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=11.47 //y=7.4 //x2=11.47 //y2=7.4
r568 (  22 24 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=11.47 //y=7.4 //x2=12.58 //y2=7.4
r569 (  20 300 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=10.36 //y=7.4 //x2=10.36 //y2=7.4
r570 (  20 22 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=10.36 //y=7.4 //x2=11.47 //y2=7.4
r571 (  18 136 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=8.88 //y=7.4 //x2=8.88 //y2=7.4
r572 (  18 20 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=8.88 //y=7.4 //x2=10.36 //y2=7.4
r573 (  16 126 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=7.77 //y=7.4 //x2=7.77 //y2=7.4
r574 (  16 18 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=7.77 //y=7.4 //x2=8.88 //y2=7.4
r575 (  14 108 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=6.66 //y=7.4 //x2=6.66 //y2=7.4
r576 (  14 16 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=6.66 //y=7.4 //x2=7.77 //y2=7.4
r577 (  12 98 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r578 (  12 14 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.66 //y2=7.4
r579 (  10 92 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=7.4 //x2=4.07 //y2=7.4
r580 (  10 12 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=7.4 //x2=5.55 //y2=7.4
r581 (  8 82 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r582 (  8 10 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r583 (  6 64 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r584 (  6 8 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r585 (  3 54 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r586 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r587 (  1 27 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=12.95 //y=7.4 //x2=14.06 //y2=7.4
r588 (  1 24 ) resistor r=0.153654 //w=0.301 //l=0.37 //layer=m1 \
 //thickness=0.36 //x=12.95 //y=7.4 //x2=12.58 //y2=7.4
ends PM_DFFRNX1\%VDD

subckt PM_DFFRNX1\%noxref_3 ( 1 2 3 4 12 25 26 33 41 47 48 52 54 61 62 63 64 \
 65 66 67 68 72 73 74 79 81 84 85 86 87 88 89 93 95 98 99 104 105 110 119 122 \
 124 125 126 )
c246 ( 126 0 ) capacitor c=0.023087f //x=7.955 //y=5.02
c247 ( 125 0 ) capacitor c=0.023519f //x=7.075 //y=5.02
c248 ( 124 0 ) capacitor c=0.0224735f //x=6.195 //y=5.02
c249 ( 122 0 ) capacitor c=0.00872971f //x=8.205 //y=0.915
c250 ( 119 0 ) capacitor c=0.0588816f //x=10.73 //y=4.7
c251 ( 110 0 ) capacitor c=0.058931f //x=3.33 //y=4.7
c252 ( 105 0 ) capacitor c=0.0273931f //x=3.33 //y=1.915
c253 ( 104 0 ) capacitor c=0.0464411f //x=3.33 //y=2.08
c254 ( 99 0 ) capacitor c=0.0318948f //x=11.065 //y=1.21
c255 ( 98 0 ) capacitor c=0.0187384f //x=11.065 //y=0.865
c256 ( 95 0 ) capacitor c=0.0141798f //x=10.91 //y=1.365
c257 ( 93 0 ) capacitor c=0.0149844f //x=10.91 //y=0.71
c258 ( 89 0 ) capacitor c=0.0813322f //x=10.535 //y=1.915
c259 ( 88 0 ) capacitor c=0.0229267f //x=10.535 //y=1.52
c260 ( 87 0 ) capacitor c=0.0234352f //x=10.535 //y=1.21
c261 ( 86 0 ) capacitor c=0.0199343f //x=10.535 //y=0.865
c262 ( 85 0 ) capacitor c=0.0432517f //x=3.85 //y=1.26
c263 ( 84 0 ) capacitor c=0.0200379f //x=3.85 //y=0.915
c264 ( 81 0 ) capacitor c=0.0158629f //x=3.695 //y=1.415
c265 ( 79 0 ) capacitor c=0.0157803f //x=3.695 //y=0.76
c266 ( 74 0 ) capacitor c=0.0218028f //x=3.32 //y=1.57
c267 ( 73 0 ) capacitor c=0.0207459f //x=3.32 //y=1.26
c268 ( 72 0 ) capacitor c=0.0194308f //x=3.32 //y=0.915
c269 ( 68 0 ) capacitor c=0.110275f //x=11.07 //y=6.02
c270 ( 67 0 ) capacitor c=0.154305f //x=10.63 //y=6.02
c271 ( 66 0 ) capacitor c=0.158794f //x=3.51 //y=6.02
c272 ( 65 0 ) capacitor c=0.110114f //x=3.07 //y=6.02
c273 ( 62 0 ) capacitor c=0.00106608f //x=8.1 //y=5.155
c274 ( 61 0 ) capacitor c=0.00207319f //x=7.22 //y=5.155
c275 ( 54 0 ) capacitor c=0.0894789f //x=10.73 //y=2.08
c276 ( 52 0 ) capacitor c=0.108812f //x=8.88 //y=3.33
c277 ( 48 0 ) capacitor c=0.00398962f //x=8.48 //y=1.665
c278 ( 47 0 ) capacitor c=0.0137288f //x=8.795 //y=1.665
c279 ( 41 0 ) capacitor c=0.0284988f //x=8.795 //y=5.155
c280 ( 33 0 ) capacitor c=0.0176454f //x=8.015 //y=5.155
c281 ( 26 0 ) capacitor c=0.00332903f //x=6.425 //y=5.155
c282 ( 25 0 ) capacitor c=0.0148427f //x=7.135 //y=5.155
c283 ( 12 0 ) capacitor c=0.0883349f //x=3.33 //y=2.08
c284 ( 4 0 ) capacitor c=0.00479603f //x=8.995 //y=3.33
c285 ( 3 0 ) capacitor c=0.0449509f //x=10.615 //y=3.33
c286 ( 2 0 ) capacitor c=0.0164246f //x=3.445 //y=3.33
c287 ( 1 0 ) capacitor c=0.144217f //x=8.765 //y=3.33
r288 (  117 119 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=10.63 //y=4.7 //x2=10.73 //y2=4.7
r289 (  104 105 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.33 //y=2.08 //x2=3.33 //y2=1.915
r290 (  100 119 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=11.07 //y=4.865 //x2=10.73 //y2=4.7
r291 (  99 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.065 //y=1.21 //x2=11.025 //y2=1.365
r292 (  98 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.065 //y=0.865 //x2=11.025 //y2=0.71
r293 (  98 99 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.065 //y=0.865 //x2=11.065 //y2=1.21
r294 (  96 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.69 //y=1.365 //x2=10.575 //y2=1.365
r295 (  95 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.91 //y=1.365 //x2=11.025 //y2=1.365
r296 (  94 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.69 //y=0.71 //x2=10.575 //y2=0.71
r297 (  93 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=10.91 //y=0.71 //x2=11.025 //y2=0.71
r298 (  93 94 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=10.91 //y=0.71 //x2=10.69 //y2=0.71
r299 (  90 117 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=10.63 //y=4.865 //x2=10.63 //y2=4.7
r300 (  89 114 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=10.535 //y=1.915 //x2=10.73 //y2=2.08
r301 (  88 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.535 //y=1.52 //x2=10.575 //y2=1.365
r302 (  88 89 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=10.535 //y=1.52 //x2=10.535 //y2=1.915
r303 (  87 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.535 //y=1.21 //x2=10.575 //y2=1.365
r304 (  86 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=10.535 //y=0.865 //x2=10.575 //y2=0.71
r305 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=10.535 //y=0.865 //x2=10.535 //y2=1.21
r306 (  85 112 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=1.26 //x2=3.81 //y2=1.415
r307 (  84 111 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.81 //y2=0.76
r308 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.85 //y2=1.26
r309 (  82 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=1.415 //x2=3.36 //y2=1.415
r310 (  81 112 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=1.415 //x2=3.81 //y2=1.415
r311 (  80 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=0.76 //x2=3.36 //y2=0.76
r312 (  79 111 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.81 //y2=0.76
r313 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.475 //y2=0.76
r314 (  76 110 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=3.51 //y=4.865 //x2=3.33 //y2=4.7
r315 (  74 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.36 //y2=1.415
r316 (  74 105 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.32 //y2=1.915
r317 (  73 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.26 //x2=3.36 //y2=1.415
r318 (  72 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.36 //y2=0.76
r319 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.32 //y2=1.26
r320 (  69 110 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=3.07 //y=4.865 //x2=3.33 //y2=4.7
r321 (  68 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.07 //y=6.02 //x2=11.07 //y2=4.865
r322 (  67 90 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=10.63 //y=6.02 //x2=10.63 //y2=4.865
r323 (  66 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.51 //y=6.02 //x2=3.51 //y2=4.865
r324 (  65 69 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.07 //y=6.02 //x2=3.07 //y2=4.865
r325 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.8 //y=1.365 //x2=10.91 //y2=1.365
r326 (  64 96 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=10.8 //y=1.365 //x2=10.69 //y2=1.365
r327 (  63 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.695 //y2=1.415
r328 (  63 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.475 //y2=1.415
r329 (  59 119 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=4.7 //x2=10.73 //y2=4.7
r330 (  57 59 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=10.73 //y=3.33 //x2=10.73 //y2=4.7
r331 (  54 114 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=10.73 //y=2.08 //x2=10.73 //y2=2.08
r332 (  54 57 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=10.73 //y=2.08 //x2=10.73 //y2=3.33
r333 (  50 52 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=8.88 //y=5.07 //x2=8.88 //y2=3.33
r334 (  49 52 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=8.88 //y=1.75 //x2=8.88 //y2=3.33
r335 (  47 49 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.795 //y=1.665 //x2=8.88 //y2=1.75
r336 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=8.795 //y=1.665 //x2=8.48 //y2=1.665
r337 (  43 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.395 //y=1.58 //x2=8.48 //y2=1.665
r338 (  43 122 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=8.395 //y=1.58 //x2=8.395 //y2=1.01
r339 (  42 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.185 //y=5.155 //x2=8.1 //y2=5.155
r340 (  41 50 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=8.795 //y=5.155 //x2=8.88 //y2=5.07
r341 (  41 42 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=8.795 //y=5.155 //x2=8.185 //y2=5.155
r342 (  35 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.1 //y=5.24 //x2=8.1 //y2=5.155
r343 (  35 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=8.1 //y=5.24 //x2=8.1 //y2=5.725
r344 (  34 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.305 //y=5.155 //x2=7.22 //y2=5.155
r345 (  33 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=8.015 //y=5.155 //x2=8.1 //y2=5.155
r346 (  33 34 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=8.015 //y=5.155 //x2=7.305 //y2=5.155
r347 (  27 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.24 //x2=7.22 //y2=5.155
r348 (  27 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=7.22 //y=5.24 //x2=7.22 //y2=5.725
r349 (  25 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.155 //x2=7.22 //y2=5.155
r350 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=7.135 //y=5.155 //x2=6.425 //y2=5.155
r351 (  19 26 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.24 //x2=6.425 //y2=5.155
r352 (  19 124 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=6.34 //y=5.24 //x2=6.34 //y2=5.725
r353 (  17 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r354 (  15 17 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=3.33 //y=3.33 //x2=3.33 //y2=4.7
r355 (  12 104 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r356 (  12 15 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=3.33 //y=2.08 //x2=3.33 //y2=3.33
r357 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=10.73 //y=3.33 //x2=10.73 //y2=3.33
r358 (  8 52 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.88 //y=3.33 //x2=8.88 //y2=3.33
r359 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=3.33 //y=3.33 //x2=3.33 //y2=3.33
r360 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.995 //y=3.33 //x2=8.88 //y2=3.33
r361 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=10.615 //y=3.33 //x2=10.73 //y2=3.33
r362 (  3 4 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=10.615 //y=3.33 //x2=8.995 //y2=3.33
r363 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.445 //y=3.33 //x2=3.33 //y2=3.33
r364 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=3.33 //x2=8.88 //y2=3.33
r365 (  1 2 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=8.765 //y=3.33 //x2=3.445 //y2=3.33
ends PM_DFFRNX1\%noxref_3

subckt PM_DFFRNX1\%noxref_4 ( 1 2 13 14 25 27 28 32 34 41 42 43 44 45 46 47 48 \
 49 51 57 58 59 60 72 74 75 )
c147 ( 75 0 ) capacitor c=0.0220291f //x=11.585 //y=5.02
c148 ( 74 0 ) capacitor c=0.0217503f //x=10.705 //y=5.02
c149 ( 72 0 ) capacitor c=0.0084702f //x=11.58 //y=0.905
c150 ( 60 0 ) capacitor c=0.0556143f //x=14.335 //y=4.79
c151 ( 59 0 ) capacitor c=0.0293157f //x=14.625 //y=4.79
c152 ( 58 0 ) capacitor c=0.0347816f //x=14.29 //y=1.22
c153 ( 57 0 ) capacitor c=0.0187487f //x=14.29 //y=0.875
c154 ( 51 0 ) capacitor c=0.0137055f //x=14.135 //y=1.375
c155 ( 49 0 ) capacitor c=0.0149861f //x=14.135 //y=0.72
c156 ( 48 0 ) capacitor c=0.096037f //x=13.76 //y=1.915
c157 ( 47 0 ) capacitor c=0.0228993f //x=13.76 //y=1.53
c158 ( 46 0 ) capacitor c=0.0234352f //x=13.76 //y=1.22
c159 ( 45 0 ) capacitor c=0.0198724f //x=13.76 //y=0.875
c160 ( 44 0 ) capacitor c=0.110114f //x=14.7 //y=6.02
c161 ( 43 0 ) capacitor c=0.158956f //x=14.26 //y=6.02
c162 ( 41 0 ) capacitor c=0.00211606f //x=11.73 //y=5.2
c163 ( 34 0 ) capacitor c=0.0995893f //x=14.06 //y=2.08
c164 ( 32 0 ) capacitor c=0.10775f //x=12.21 //y=3.33
c165 ( 28 0 ) capacitor c=0.00404073f //x=11.855 //y=1.655
c166 ( 27 0 ) capacitor c=0.0122201f //x=12.125 //y=1.655
c167 ( 25 0 ) capacitor c=0.0137995f //x=12.125 //y=5.2
c168 ( 14 0 ) capacitor c=0.00251635f //x=10.935 //y=5.2
c169 ( 13 0 ) capacitor c=0.0143649f //x=11.645 //y=5.2
c170 ( 2 0 ) capacitor c=0.00733653f //x=12.325 //y=3.33
c171 ( 1 0 ) capacitor c=0.0503252f //x=13.945 //y=3.33
r172 (  59 61 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=14.625 //y=4.79 //x2=14.7 //y2=4.865
r173 (  59 60 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=14.625 //y=4.79 //x2=14.335 //y2=4.79
r174 (  58 71 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.29 //y=1.22 //x2=14.25 //y2=1.375
r175 (  57 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.29 //y=0.875 //x2=14.25 //y2=0.72
r176 (  57 58 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=14.29 //y=0.875 //x2=14.29 //y2=1.22
r177 (  54 60 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=14.26 //y=4.865 //x2=14.335 //y2=4.79
r178 (  54 69 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=14.26 //y=4.865 //x2=14.06 //y2=4.7
r179 (  52 65 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.915 //y=1.375 //x2=13.8 //y2=1.375
r180 (  51 71 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.135 //y=1.375 //x2=14.25 //y2=1.375
r181 (  50 64 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=13.915 //y=0.72 //x2=13.8 //y2=0.72
r182 (  49 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.135 //y=0.72 //x2=14.25 //y2=0.72
r183 (  49 50 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=14.135 //y=0.72 //x2=13.915 //y2=0.72
r184 (  48 67 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=13.76 //y=1.915 //x2=14.06 //y2=2.08
r185 (  47 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.76 //y=1.53 //x2=13.8 //y2=1.375
r186 (  47 48 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=13.76 //y=1.53 //x2=13.76 //y2=1.915
r187 (  46 65 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.76 //y=1.22 //x2=13.8 //y2=1.375
r188 (  45 64 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=13.76 //y=0.875 //x2=13.8 //y2=0.72
r189 (  45 46 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=13.76 //y=0.875 //x2=13.76 //y2=1.22
r190 (  44 61 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.7 //y=6.02 //x2=14.7 //y2=4.865
r191 (  43 54 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=14.26 //y=6.02 //x2=14.26 //y2=4.865
r192 (  42 51 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.025 //y=1.375 //x2=14.135 //y2=1.375
r193 (  42 52 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=14.025 //y=1.375 //x2=13.915 //y2=1.375
r194 (  39 69 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=4.7 //x2=14.06 //y2=4.7
r195 (  37 39 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=14.06 //y=3.33 //x2=14.06 //y2=4.7
r196 (  34 67 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=14.06 //y=2.08 //x2=14.06 //y2=2.08
r197 (  34 37 ) resistor r=85.5615 //w=0.187 //l=1.25 //layer=li \
 //thickness=0.1 //x=14.06 //y=2.08 //x2=14.06 //y2=3.33
r198 (  30 32 ) resistor r=122.182 //w=0.187 //l=1.785 //layer=li \
 //thickness=0.1 //x=12.21 //y=5.115 //x2=12.21 //y2=3.33
r199 (  29 32 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=12.21 //y=1.74 //x2=12.21 //y2=3.33
r200 (  27 29 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.125 //y=1.655 //x2=12.21 //y2=1.74
r201 (  27 28 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=12.125 //y=1.655 //x2=11.855 //y2=1.655
r202 (  26 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.815 //y=5.2 //x2=11.73 //y2=5.2
r203 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=12.125 //y=5.2 //x2=12.21 //y2=5.115
r204 (  25 26 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=12.125 //y=5.2 //x2=11.815 //y2=5.2
r205 (  21 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=11.77 //y=1.57 //x2=11.855 //y2=1.655
r206 (  21 72 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=11.77 //y=1.57 //x2=11.77 //y2=1
r207 (  15 41 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.73 //y=5.285 //x2=11.73 //y2=5.2
r208 (  15 75 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=11.73 //y=5.285 //x2=11.73 //y2=5.725
r209 (  13 41 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=11.645 //y=5.2 //x2=11.73 //y2=5.2
r210 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=11.645 //y=5.2 //x2=10.935 //y2=5.2
r211 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=10.85 //y=5.285 //x2=10.935 //y2=5.2
r212 (  7 74 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=10.85 //y=5.285 //x2=10.85 //y2=5.725
r213 (  6 37 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=14.06 //y=3.33 //x2=14.06 //y2=3.33
r214 (  4 32 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=12.21 //y=3.33 //x2=12.21 //y2=3.33
r215 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=12.325 //y=3.33 //x2=12.21 //y2=3.33
r216 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=13.945 //y=3.33 //x2=14.06 //y2=3.33
r217 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=13.945 //y=3.33 //x2=12.325 //y2=3.33
ends PM_DFFRNX1\%noxref_4

subckt PM_DFFRNX1\%CLK ( 1 2 7 8 9 10 11 12 13 14 15 16 17 19 32 43 44 45 46 \
 47 48 49 50 51 53 59 60 61 62 63 68 69 70 72 78 79 80 81 82 90 101 )
c215 ( 101 0 ) capacitor c=0.0334842f //x=15.17 //y=4.7
c216 ( 90 0 ) capacitor c=0.0334842f //x=2.22 //y=4.7
c217 ( 82 0 ) capacitor c=0.0249231f //x=15.505 //y=4.79
c218 ( 81 0 ) capacitor c=0.0825763f //x=15.26 //y=1.915
c219 ( 80 0 ) capacitor c=0.0170266f //x=15.26 //y=1.45
c220 ( 79 0 ) capacitor c=0.018609f //x=15.26 //y=1.22
c221 ( 78 0 ) capacitor c=0.0187309f //x=15.26 //y=0.91
c222 ( 72 0 ) capacitor c=0.014725f //x=15.105 //y=1.375
c223 ( 70 0 ) capacitor c=0.0146567f //x=15.105 //y=0.755
c224 ( 69 0 ) capacitor c=0.0335408f //x=14.735 //y=1.22
c225 ( 68 0 ) capacitor c=0.0173761f //x=14.735 //y=0.91
c226 ( 63 0 ) capacitor c=0.0245352f //x=2.555 //y=4.79
c227 ( 62 0 ) capacitor c=0.0850619f //x=2.31 //y=1.915
c228 ( 61 0 ) capacitor c=0.0170266f //x=2.31 //y=1.45
c229 ( 60 0 ) capacitor c=0.018609f //x=2.31 //y=1.22
c230 ( 59 0 ) capacitor c=0.0187309f //x=2.31 //y=0.91
c231 ( 53 0 ) capacitor c=0.014725f //x=2.155 //y=1.375
c232 ( 51 0 ) capacitor c=0.0146567f //x=2.155 //y=0.755
c233 ( 50 0 ) capacitor c=0.0335408f //x=1.785 //y=1.22
c234 ( 49 0 ) capacitor c=0.0173761f //x=1.785 //y=0.91
c235 ( 48 0 ) capacitor c=0.110114f //x=15.58 //y=6.02
c236 ( 47 0 ) capacitor c=0.11012f //x=15.14 //y=6.02
c237 ( 46 0 ) capacitor c=0.110114f //x=2.63 //y=6.02
c238 ( 45 0 ) capacitor c=0.11012f //x=2.19 //y=6.02
c239 ( 32 0 ) capacitor c=0.0952742f //x=15.17 //y=2.08
c240 ( 19 0 ) capacitor c=0.100158f //x=2.22 //y=2.08
c241 ( 2 0 ) capacitor c=0.0154455f //x=2.335 //y=4.44
c242 ( 1 0 ) capacitor c=0.301662f //x=15.055 //y=4.44
r243 (  103 104 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=15.17 //y=4.79 //x2=15.17 //y2=4.865
r244 (  101 103 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=15.17 //y=4.7 //x2=15.17 //y2=4.79
r245 (  92 93 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.79 //x2=2.22 //y2=4.865
r246 (  90 92 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.7 //x2=2.22 //y2=4.79
r247 (  83 103 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=15.305 //y=4.79 //x2=15.17 //y2=4.79
r248 (  82 84 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=15.505 //y=4.79 //x2=15.58 //y2=4.865
r249 (  82 83 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=15.505 //y=4.79 //x2=15.305 //y2=4.79
r250 (  81 108 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=15.26 //y=1.915 //x2=15.185 //y2=2.08
r251 (  80 106 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=15.26 //y=1.45 //x2=15.22 //y2=1.375
r252 (  80 81 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=15.26 //y=1.45 //x2=15.26 //y2=1.915
r253 (  79 106 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.26 //y=1.22 //x2=15.22 //y2=1.375
r254 (  78 105 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=15.26 //y=0.91 //x2=15.22 //y2=0.755
r255 (  78 79 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=15.26 //y=0.91 //x2=15.26 //y2=1.22
r256 (  73 99 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.89 //y=1.375 //x2=14.775 //y2=1.375
r257 (  72 106 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.105 //y=1.375 //x2=15.22 //y2=1.375
r258 (  71 98 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=14.89 //y=0.755 //x2=14.775 //y2=0.755
r259 (  70 105 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=15.105 //y=0.755 //x2=15.22 //y2=0.755
r260 (  70 71 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=15.105 //y=0.755 //x2=14.89 //y2=0.755
r261 (  69 99 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.735 //y=1.22 //x2=14.775 //y2=1.375
r262 (  68 98 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=14.735 //y=0.91 //x2=14.775 //y2=0.755
r263 (  68 69 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=14.735 //y=0.91 //x2=14.735 //y2=1.22
r264 (  64 92 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.355 //y=4.79 //x2=2.22 //y2=4.79
r265 (  63 65 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.63 //y2=4.865
r266 (  63 64 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.355 //y2=4.79
r267 (  62 97 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.915 //x2=2.235 //y2=2.08
r268 (  61 95 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.27 //y2=1.375
r269 (  61 62 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.31 //y2=1.915
r270 (  60 95 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.22 //x2=2.27 //y2=1.375
r271 (  59 94 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.27 //y2=0.755
r272 (  59 60 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.31 //y2=1.22
r273 (  54 88 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=1.375 //x2=1.825 //y2=1.375
r274 (  53 95 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=1.375 //x2=2.27 //y2=1.375
r275 (  52 87 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=0.755 //x2=1.825 //y2=0.755
r276 (  51 94 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=2.27 //y2=0.755
r277 (  51 52 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=1.94 //y2=0.755
r278 (  50 88 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=1.22 //x2=1.825 //y2=1.375
r279 (  49 87 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.825 //y2=0.755
r280 (  49 50 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.785 //y2=1.22
r281 (  48 84 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.58 //y=6.02 //x2=15.58 //y2=4.865
r282 (  47 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=15.14 //y=6.02 //x2=15.14 //y2=4.865
r283 (  46 65 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.63 //y=6.02 //x2=2.63 //y2=4.865
r284 (  45 93 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.19 //y=6.02 //x2=2.19 //y2=4.865
r285 (  44 72 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=14.997 //y=1.375 //x2=15.105 //y2=1.375
r286 (  44 73 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=14.997 //y=1.375 //x2=14.89 //y2=1.375
r287 (  43 53 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=2.155 //y2=1.375
r288 (  43 54 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=1.94 //y2=1.375
r289 (  41 101 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.17 //y=4.7 //x2=15.17 //y2=4.7
r290 (  32 108 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=15.17 //y=2.08 //x2=15.17 //y2=2.08
r291 (  29 90 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=4.7 //x2=2.22 //y2=4.7
r292 (  19 97 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=2.08
r293 (  17 41 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=15.17 //y=4.44 //x2=15.17 //y2=4.7
r294 (  16 17 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=15.17 //y=3.33 //x2=15.17 //y2=4.44
r295 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=15.17 //y=2.96 //x2=15.17 //y2=3.33
r296 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=15.17 //y=2.59 //x2=15.17 //y2=2.96
r297 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=15.17 //y=2.22 //x2=15.17 //y2=2.59
r298 (  13 32 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=15.17 //y=2.22 //x2=15.17 //y2=2.08
r299 (  12 29 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=2.22 //y=4.44 //x2=2.22 //y2=4.7
r300 (  11 12 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.7 //x2=2.22 //y2=4.44
r301 (  10 11 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=3.33 //x2=2.22 //y2=3.7
r302 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.96 //x2=2.22 //y2=3.33
r303 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=2.22 //y=2.59 //x2=2.22 //y2=2.96
r304 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=2.22 //y=2.22 //x2=2.22 //y2=2.59
r305 (  7 19 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=2.22 //y=2.22 //x2=2.22 //y2=2.08
r306 (  6 17 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=15.17 //y=4.44 //x2=15.17 //y2=4.44
r307 (  4 12 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.22 //y=4.44 //x2=2.22 //y2=4.44
r308 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.335 //y=4.44 //x2=2.22 //y2=4.44
r309 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=15.055 //y=4.44 //x2=15.17 //y2=4.44
r310 (  1 2 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=15.055 //y=4.44 //x2=2.335 //y2=4.44
ends PM_DFFRNX1\%CLK

subckt PM_DFFRNX1\%noxref_6 ( 1 2 3 4 17 18 25 33 39 40 44 46 54 61 62 63 64 \
 65 66 67 68 69 70 71 72 73 75 81 82 83 84 88 89 90 91 92 94 100 101 102 103 \
 123 125 126 127 )
c246 ( 127 0 ) capacitor c=0.023087f //x=3.145 //y=5.02
c247 ( 126 0 ) capacitor c=0.023519f //x=2.265 //y=5.02
c248 ( 125 0 ) capacitor c=0.0224735f //x=1.385 //y=5.02
c249 ( 123 0 ) capacitor c=0.00853354f //x=3.395 //y=0.915
c250 ( 103 0 ) capacitor c=0.0558396f //x=19.145 //y=4.79
c251 ( 102 0 ) capacitor c=0.0298189f //x=19.435 //y=4.79
c252 ( 101 0 ) capacitor c=0.0347816f //x=19.1 //y=1.22
c253 ( 100 0 ) capacitor c=0.0187487f //x=19.1 //y=0.875
c254 ( 94 0 ) capacitor c=0.0137055f //x=18.945 //y=1.375
c255 ( 92 0 ) capacitor c=0.0149861f //x=18.945 //y=0.72
c256 ( 91 0 ) capacitor c=0.096037f //x=18.57 //y=1.915
c257 ( 90 0 ) capacitor c=0.0228993f //x=18.57 //y=1.53
c258 ( 89 0 ) capacitor c=0.0234352f //x=18.57 //y=1.22
c259 ( 88 0 ) capacitor c=0.0198724f //x=18.57 //y=0.875
c260 ( 84 0 ) capacitor c=0.0556143f //x=6.195 //y=4.79
c261 ( 83 0 ) capacitor c=0.0293157f //x=6.485 //y=4.79
c262 ( 82 0 ) capacitor c=0.0347816f //x=6.15 //y=1.22
c263 ( 81 0 ) capacitor c=0.0187487f //x=6.15 //y=0.875
c264 ( 75 0 ) capacitor c=0.0137055f //x=5.995 //y=1.375
c265 ( 73 0 ) capacitor c=0.0149861f //x=5.995 //y=0.72
c266 ( 72 0 ) capacitor c=0.102158f //x=5.62 //y=1.915
c267 ( 71 0 ) capacitor c=0.0229444f //x=5.62 //y=1.53
c268 ( 70 0 ) capacitor c=0.0234352f //x=5.62 //y=1.22
c269 ( 69 0 ) capacitor c=0.0198724f //x=5.62 //y=0.875
c270 ( 68 0 ) capacitor c=0.110114f //x=19.51 //y=6.02
c271 ( 67 0 ) capacitor c=0.158956f //x=19.07 //y=6.02
c272 ( 66 0 ) capacitor c=0.110114f //x=6.56 //y=6.02
c273 ( 65 0 ) capacitor c=0.158956f //x=6.12 //y=6.02
c274 ( 62 0 ) capacitor c=0.00106608f //x=3.29 //y=5.155
c275 ( 61 0 ) capacitor c=0.00207162f //x=2.41 //y=5.155
c276 ( 54 0 ) capacitor c=0.106024f //x=18.87 //y=2.08
c277 ( 46 0 ) capacitor c=0.102261f //x=5.92 //y=2.08
c278 ( 44 0 ) capacitor c=0.109709f //x=4.07 //y=3.7
c279 ( 40 0 ) capacitor c=0.00493499f //x=3.67 //y=1.665
c280 ( 39 0 ) capacitor c=0.0154052f //x=3.985 //y=1.665
c281 ( 33 0 ) capacitor c=0.0283082f //x=3.985 //y=5.155
c282 ( 25 0 ) capacitor c=0.0176454f //x=3.205 //y=5.155
c283 ( 18 0 ) capacitor c=0.00351598f //x=1.615 //y=5.155
c284 ( 17 0 ) capacitor c=0.0154196f //x=2.325 //y=5.155
c285 ( 4 0 ) capacitor c=0.00424246f //x=6.035 //y=3.7
c286 ( 3 0 ) capacitor c=0.237637f //x=18.755 //y=3.7
c287 ( 2 0 ) capacitor c=0.0125346f //x=4.185 //y=3.7
c288 ( 1 0 ) capacitor c=0.0288301f //x=5.805 //y=3.7
r289 (  102 104 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=19.435 //y=4.79 //x2=19.51 //y2=4.865
r290 (  102 103 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=19.435 //y=4.79 //x2=19.145 //y2=4.79
r291 (  101 122 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.1 //y=1.22 //x2=19.06 //y2=1.375
r292 (  100 121 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.1 //y=0.875 //x2=19.06 //y2=0.72
r293 (  100 101 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=19.1 //y=0.875 //x2=19.1 //y2=1.22
r294 (  97 103 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=19.07 //y=4.865 //x2=19.145 //y2=4.79
r295 (  97 120 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=19.07 //y=4.865 //x2=18.87 //y2=4.7
r296 (  95 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.725 //y=1.375 //x2=18.61 //y2=1.375
r297 (  94 122 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.945 //y=1.375 //x2=19.06 //y2=1.375
r298 (  93 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.725 //y=0.72 //x2=18.61 //y2=0.72
r299 (  92 121 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=18.945 //y=0.72 //x2=19.06 //y2=0.72
r300 (  92 93 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=18.945 //y=0.72 //x2=18.725 //y2=0.72
r301 (  91 118 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=18.57 //y=1.915 //x2=18.87 //y2=2.08
r302 (  90 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.57 //y=1.53 //x2=18.61 //y2=1.375
r303 (  90 91 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=18.57 //y=1.53 //x2=18.57 //y2=1.915
r304 (  89 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.57 //y=1.22 //x2=18.61 //y2=1.375
r305 (  88 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=18.57 //y=0.875 //x2=18.61 //y2=0.72
r306 (  88 89 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=18.57 //y=0.875 //x2=18.57 //y2=1.22
r307 (  83 85 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.485 //y=4.79 //x2=6.56 //y2=4.865
r308 (  83 84 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=6.485 //y=4.79 //x2=6.195 //y2=4.79
r309 (  82 114 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.15 //y=1.22 //x2=6.11 //y2=1.375
r310 (  81 113 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.15 //y=0.875 //x2=6.11 //y2=0.72
r311 (  81 82 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.15 //y=0.875 //x2=6.15 //y2=1.22
r312 (  78 84 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.12 //y=4.865 //x2=6.195 //y2=4.79
r313 (  78 112 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=6.12 //y=4.865 //x2=5.92 //y2=4.7
r314 (  76 108 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.775 //y=1.375 //x2=5.66 //y2=1.375
r315 (  75 114 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.995 //y=1.375 //x2=6.11 //y2=1.375
r316 (  74 107 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.775 //y=0.72 //x2=5.66 //y2=0.72
r317 (  73 113 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.995 //y=0.72 //x2=6.11 //y2=0.72
r318 (  73 74 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=5.995 //y=0.72 //x2=5.775 //y2=0.72
r319 (  72 110 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.915 //x2=5.92 //y2=2.08
r320 (  71 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.53 //x2=5.66 //y2=1.375
r321 (  71 72 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.53 //x2=5.62 //y2=1.915
r322 (  70 108 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=1.22 //x2=5.66 //y2=1.375
r323 (  69 107 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.62 //y=0.875 //x2=5.66 //y2=0.72
r324 (  69 70 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.62 //y=0.875 //x2=5.62 //y2=1.22
r325 (  68 104 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.51 //y=6.02 //x2=19.51 //y2=4.865
r326 (  67 97 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.07 //y=6.02 //x2=19.07 //y2=4.865
r327 (  66 85 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.56 //y=6.02 //x2=6.56 //y2=4.865
r328 (  65 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.12 //y=6.02 //x2=6.12 //y2=4.865
r329 (  64 94 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.835 //y=1.375 //x2=18.945 //y2=1.375
r330 (  64 95 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=18.835 //y=1.375 //x2=18.725 //y2=1.375
r331 (  63 75 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.375 //x2=5.995 //y2=1.375
r332 (  63 76 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.885 //y=1.375 //x2=5.775 //y2=1.375
r333 (  59 120 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.87 //y=4.7 //x2=18.87 //y2=4.7
r334 (  57 59 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=18.87 //y=3.7 //x2=18.87 //y2=4.7
r335 (  54 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=18.87 //y=2.08 //x2=18.87 //y2=2.08
r336 (  54 57 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=18.87 //y=2.08 //x2=18.87 //y2=3.7
r337 (  51 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=4.7 //x2=5.92 //y2=4.7
r338 (  49 51 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=5.92 //y=3.7 //x2=5.92 //y2=4.7
r339 (  46 110 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.92 //y=2.08 //x2=5.92 //y2=2.08
r340 (  46 49 ) resistor r=110.888 //w=0.187 //l=1.62 //layer=li \
 //thickness=0.1 //x=5.92 //y=2.08 //x2=5.92 //y2=3.7
r341 (  42 44 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=4.07 //y=5.07 //x2=4.07 //y2=3.7
r342 (  41 44 ) resistor r=133.476 //w=0.187 //l=1.95 //layer=li \
 //thickness=0.1 //x=4.07 //y=1.75 //x2=4.07 //y2=3.7
r343 (  39 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=4.07 //y2=1.75
r344 (  39 40 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=3.67 //y2=1.665
r345 (  35 40 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.67 //y2=1.665
r346 (  35 123 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.585 //y2=1.01
r347 (  34 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.375 //y=5.155 //x2=3.29 //y2=5.155
r348 (  33 42 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=4.07 //y2=5.07
r349 (  33 34 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=3.375 //y2=5.155
r350 (  27 62 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.155
r351 (  27 127 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.725
r352 (  26 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.495 //y=5.155 //x2=2.41 //y2=5.155
r353 (  25 62 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=3.29 //y2=5.155
r354 (  25 26 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=2.495 //y2=5.155
r355 (  19 61 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.155
r356 (  19 126 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.725
r357 (  17 61 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=2.41 //y2=5.155
r358 (  17 18 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=1.615 //y2=5.155
r359 (  11 18 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.615 //y2=5.155
r360 (  11 125 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.53 //y2=5.725
r361 (  10 57 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=18.87 //y=3.7 //x2=18.87 //y2=3.7
r362 (  8 49 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.92 //y=3.7 //x2=5.92 //y2=3.7
r363 (  6 44 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=3.7 //x2=4.07 //y2=3.7
r364 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=6.035 //y=3.7 //x2=5.92 //y2=3.7
r365 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=18.755 //y=3.7 //x2=18.87 //y2=3.7
r366 (  3 4 ) resistor r=12.1374 //w=0.131 //l=12.72 //layer=m1 \
 //thickness=0.36 //x=18.755 //y=3.7 //x2=6.035 //y2=3.7
r367 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.185 //y=3.7 //x2=4.07 //y2=3.7
r368 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.805 //y=3.7 //x2=5.92 //y2=3.7
r369 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=5.805 //y=3.7 //x2=4.185 //y2=3.7
ends PM_DFFRNX1\%noxref_6

subckt PM_DFFRNX1\%RN ( 1 2 3 4 11 12 13 14 15 16 17 18 20 30 38 49 50 51 52 \
 53 54 55 56 57 61 62 63 68 70 73 74 78 79 80 85 87 90 91 92 93 94 96 102 103 \
 104 105 106 112 113 118 122 123 128 134 )
c269 ( 134 0 ) capacitor c=0.0336203f //x=19.98 //y=4.7
c270 ( 128 0 ) capacitor c=0.0593675f //x=16.28 //y=4.7
c271 ( 123 0 ) capacitor c=0.0273931f //x=16.28 //y=1.915
c272 ( 122 0 ) capacitor c=0.0461462f //x=16.28 //y=2.08
c273 ( 118 0 ) capacitor c=0.0587755f //x=8.14 //y=4.7
c274 ( 113 0 ) capacitor c=0.0273931f //x=8.14 //y=1.915
c275 ( 112 0 ) capacitor c=0.0463246f //x=8.14 //y=2.08
c276 ( 106 0 ) capacitor c=0.024933f //x=20.315 //y=4.79
c277 ( 105 0 ) capacitor c=0.0831166f //x=20.07 //y=1.915
c278 ( 104 0 ) capacitor c=0.0170266f //x=20.07 //y=1.45
c279 ( 103 0 ) capacitor c=0.018609f //x=20.07 //y=1.22
c280 ( 102 0 ) capacitor c=0.0187309f //x=20.07 //y=0.91
c281 ( 96 0 ) capacitor c=0.014725f //x=19.915 //y=1.375
c282 ( 94 0 ) capacitor c=0.0146567f //x=19.915 //y=0.755
c283 ( 93 0 ) capacitor c=0.0335408f //x=19.545 //y=1.22
c284 ( 92 0 ) capacitor c=0.0173761f //x=19.545 //y=0.91
c285 ( 91 0 ) capacitor c=0.0432517f //x=16.8 //y=1.26
c286 ( 90 0 ) capacitor c=0.0200379f //x=16.8 //y=0.915
c287 ( 87 0 ) capacitor c=0.0148873f //x=16.645 //y=1.415
c288 ( 85 0 ) capacitor c=0.0157803f //x=16.645 //y=0.76
c289 ( 80 0 ) capacitor c=0.0218028f //x=16.27 //y=1.57
c290 ( 79 0 ) capacitor c=0.0207459f //x=16.27 //y=1.26
c291 ( 78 0 ) capacitor c=0.0194308f //x=16.27 //y=0.915
c292 ( 74 0 ) capacitor c=0.0432517f //x=8.66 //y=1.26
c293 ( 73 0 ) capacitor c=0.0200379f //x=8.66 //y=0.915
c294 ( 70 0 ) capacitor c=0.0148873f //x=8.505 //y=1.415
c295 ( 68 0 ) capacitor c=0.0157803f //x=8.505 //y=0.76
c296 ( 63 0 ) capacitor c=0.0218028f //x=8.13 //y=1.57
c297 ( 62 0 ) capacitor c=0.0207459f //x=8.13 //y=1.26
c298 ( 61 0 ) capacitor c=0.0194308f //x=8.13 //y=0.915
c299 ( 57 0 ) capacitor c=0.110114f //x=20.39 //y=6.02
c300 ( 56 0 ) capacitor c=0.11012f //x=19.95 //y=6.02
c301 ( 55 0 ) capacitor c=0.158794f //x=16.46 //y=6.02
c302 ( 54 0 ) capacitor c=0.110114f //x=16.02 //y=6.02
c303 ( 53 0 ) capacitor c=0.158794f //x=8.32 //y=6.02
c304 ( 52 0 ) capacitor c=0.110114f //x=7.88 //y=6.02
c305 ( 38 0 ) capacitor c=0.0994642f //x=19.98 //y=2.08
c306 ( 30 0 ) capacitor c=0.0881589f //x=16.28 //y=2.08
c307 ( 20 0 ) capacitor c=0.0845523f //x=8.14 //y=2.08
c308 ( 4 0 ) capacitor c=0.00668196f //x=16.395 //y=2.22
c309 ( 3 0 ) capacitor c=0.115719f //x=19.865 //y=2.22
c310 ( 2 0 ) capacitor c=0.0160747f //x=8.255 //y=2.22
c311 ( 1 0 ) capacitor c=0.209784f //x=16.165 //y=2.22
r312 (  136 137 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=19.98 //y=4.79 //x2=19.98 //y2=4.865
r313 (  134 136 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=19.98 //y=4.7 //x2=19.98 //y2=4.79
r314 (  122 123 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=16.28 //y=2.08 //x2=16.28 //y2=1.915
r315 (  112 113 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=8.14 //y=2.08 //x2=8.14 //y2=1.915
r316 (  107 136 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=20.115 //y=4.79 //x2=19.98 //y2=4.79
r317 (  106 108 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=20.315 //y=4.79 //x2=20.39 //y2=4.865
r318 (  106 107 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=20.315 //y=4.79 //x2=20.115 //y2=4.79
r319 (  105 141 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=20.07 //y=1.915 //x2=19.995 //y2=2.08
r320 (  104 139 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=20.07 //y=1.45 //x2=20.03 //y2=1.375
r321 (  104 105 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=20.07 //y=1.45 //x2=20.07 //y2=1.915
r322 (  103 139 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.07 //y=1.22 //x2=20.03 //y2=1.375
r323 (  102 138 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=20.07 //y=0.91 //x2=20.03 //y2=0.755
r324 (  102 103 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=20.07 //y=0.91 //x2=20.07 //y2=1.22
r325 (  97 132 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.7 //y=1.375 //x2=19.585 //y2=1.375
r326 (  96 139 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.915 //y=1.375 //x2=20.03 //y2=1.375
r327 (  95 131 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.7 //y=0.755 //x2=19.585 //y2=0.755
r328 (  94 138 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=19.915 //y=0.755 //x2=20.03 //y2=0.755
r329 (  94 95 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=19.915 //y=0.755 //x2=19.7 //y2=0.755
r330 (  93 132 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.545 //y=1.22 //x2=19.585 //y2=1.375
r331 (  92 131 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=19.545 //y=0.91 //x2=19.585 //y2=0.755
r332 (  92 93 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=19.545 //y=0.91 //x2=19.545 //y2=1.22
r333 (  91 130 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.8 //y=1.26 //x2=16.76 //y2=1.415
r334 (  90 129 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.8 //y=0.915 //x2=16.76 //y2=0.76
r335 (  90 91 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.8 //y=0.915 //x2=16.8 //y2=1.26
r336 (  88 126 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.425 //y=1.415 //x2=16.31 //y2=1.415
r337 (  87 130 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.645 //y=1.415 //x2=16.76 //y2=1.415
r338 (  86 125 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.425 //y=0.76 //x2=16.31 //y2=0.76
r339 (  85 129 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=16.645 //y=0.76 //x2=16.76 //y2=0.76
r340 (  85 86 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=16.645 //y=0.76 //x2=16.425 //y2=0.76
r341 (  82 128 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=16.46 //y=4.865 //x2=16.28 //y2=4.7
r342 (  80 126 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.27 //y=1.57 //x2=16.31 //y2=1.415
r343 (  80 123 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.27 //y=1.57 //x2=16.27 //y2=1.915
r344 (  79 126 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.27 //y=1.26 //x2=16.31 //y2=1.415
r345 (  78 125 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=16.27 //y=0.915 //x2=16.31 //y2=0.76
r346 (  78 79 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=16.27 //y=0.915 //x2=16.27 //y2=1.26
r347 (  75 128 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=16.02 //y=4.865 //x2=16.28 //y2=4.7
r348 (  74 120 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.66 //y=1.26 //x2=8.62 //y2=1.415
r349 (  73 119 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.66 //y=0.915 //x2=8.62 //y2=0.76
r350 (  73 74 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.66 //y=0.915 //x2=8.66 //y2=1.26
r351 (  71 116 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.285 //y=1.415 //x2=8.17 //y2=1.415
r352 (  70 120 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.505 //y=1.415 //x2=8.62 //y2=1.415
r353 (  69 115 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.285 //y=0.76 //x2=8.17 //y2=0.76
r354 (  68 119 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=8.505 //y=0.76 //x2=8.62 //y2=0.76
r355 (  68 69 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=8.505 //y=0.76 //x2=8.285 //y2=0.76
r356 (  65 118 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=8.32 //y=4.865 //x2=8.14 //y2=4.7
r357 (  63 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.57 //x2=8.17 //y2=1.415
r358 (  63 113 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.57 //x2=8.13 //y2=1.915
r359 (  62 116 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=1.26 //x2=8.17 //y2=1.415
r360 (  61 115 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=8.13 //y=0.915 //x2=8.17 //y2=0.76
r361 (  61 62 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=8.13 //y=0.915 //x2=8.13 //y2=1.26
r362 (  58 118 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=7.88 //y=4.865 //x2=8.14 //y2=4.7
r363 (  57 108 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.39 //y=6.02 //x2=20.39 //y2=4.865
r364 (  56 137 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=19.95 //y=6.02 //x2=19.95 //y2=4.865
r365 (  55 82 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.46 //y=6.02 //x2=16.46 //y2=4.865
r366 (  54 75 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=16.02 //y=6.02 //x2=16.02 //y2=4.865
r367 (  53 65 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=8.32 //y=6.02 //x2=8.32 //y2=4.865
r368 (  52 58 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.88 //y=6.02 //x2=7.88 //y2=4.865
r369 (  51 96 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=19.807 //y=1.375 //x2=19.915 //y2=1.375
r370 (  51 97 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=19.807 //y=1.375 //x2=19.7 //y2=1.375
r371 (  50 87 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=16.535 //y=1.415 //x2=16.645 //y2=1.415
r372 (  50 88 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=16.535 //y=1.415 //x2=16.425 //y2=1.415
r373 (  49 70 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.395 //y=1.415 //x2=8.505 //y2=1.415
r374 (  49 71 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=8.395 //y=1.415 //x2=8.285 //y2=1.415
r375 (  47 134 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.98 //y=4.7 //x2=19.98 //y2=4.7
r376 (  38 141 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=19.98 //y=2.08 //x2=19.98 //y2=2.08
r377 (  35 128 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.28 //y=4.7 //x2=16.28 //y2=4.7
r378 (  33 35 ) resistor r=169.754 //w=0.187 //l=2.48 //layer=li \
 //thickness=0.1 //x=16.28 //y=2.22 //x2=16.28 //y2=4.7
r379 (  30 122 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=16.28 //y=2.08 //x2=16.28 //y2=2.08
r380 (  30 33 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=16.28 //y=2.08 //x2=16.28 //y2=2.22
r381 (  27 118 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.14 //y=4.7 //x2=8.14 //y2=4.7
r382 (  20 112 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=8.14 //y=2.08 //x2=8.14 //y2=2.08
r383 (  18 47 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=19.98 //y=3.7 //x2=19.98 //y2=4.7
r384 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=19.98 //y=3.33 //x2=19.98 //y2=3.7
r385 (  16 17 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.96 //x2=19.98 //y2=3.33
r386 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.59 //x2=19.98 //y2=2.96
r387 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.22 //x2=19.98 //y2=2.59
r388 (  14 38 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=19.98 //y=2.22 //x2=19.98 //y2=2.08
r389 (  13 27 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=8.14 //y=2.96 //x2=8.14 //y2=4.7
r390 (  12 13 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=8.14 //y=2.59 //x2=8.14 //y2=2.96
r391 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=8.14 //y=2.22 //x2=8.14 //y2=2.59
r392 (  11 20 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=8.14 //y=2.22 //x2=8.14 //y2=2.08
r393 (  10 14 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=19.98 //y=2.22 //x2=19.98 //y2=2.22
r394 (  8 33 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=16.28 //y=2.22 //x2=16.28 //y2=2.22
r395 (  6 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=8.14 //y=2.22 //x2=8.14 //y2=2.22
r396 (  4 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.395 //y=2.22 //x2=16.28 //y2=2.22
r397 (  3 10 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=19.865 //y=2.22 //x2=19.98 //y2=2.22
r398 (  3 4 ) resistor r=3.31107 //w=0.131 //l=3.47 //layer=m1 \
 //thickness=0.36 //x=19.865 //y=2.22 //x2=16.395 //y2=2.22
r399 (  2 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=8.255 //y=2.22 //x2=8.14 //y2=2.22
r400 (  1 8 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.165 //y=2.22 //x2=16.28 //y2=2.22
r401 (  1 2 ) resistor r=7.54771 //w=0.131 //l=7.91 //layer=m1 \
 //thickness=0.36 //x=16.165 //y=2.22 //x2=8.255 //y2=2.22
ends PM_DFFRNX1\%RN

subckt PM_DFFRNX1\%QN ( 1 2 7 8 9 10 11 12 13 14 15 16 23 24 31 39 45 46 57 67 \
 68 69 70 71 72 73 74 75 79 81 84 85 95 98 100 101 102 )
c156 ( 102 0 ) capacitor c=0.023087f //x=20.905 //y=5.02
c157 ( 101 0 ) capacitor c=0.023519f //x=20.025 //y=5.02
c158 ( 100 0 ) capacitor c=0.0224735f //x=19.145 //y=5.02
c159 ( 98 0 ) capacitor c=0.00872971f //x=21.155 //y=0.915
c160 ( 95 0 ) capacitor c=0.0593152f //x=23.68 //y=4.7
c161 ( 85 0 ) capacitor c=0.0318948f //x=24.015 //y=1.21
c162 ( 84 0 ) capacitor c=0.0187384f //x=24.015 //y=0.865
c163 ( 81 0 ) capacitor c=0.0141798f //x=23.86 //y=1.365
c164 ( 79 0 ) capacitor c=0.0149844f //x=23.86 //y=0.71
c165 ( 75 0 ) capacitor c=0.0853292f //x=23.485 //y=1.915
c166 ( 74 0 ) capacitor c=0.0229722f //x=23.485 //y=1.52
c167 ( 73 0 ) capacitor c=0.0234352f //x=23.485 //y=1.21
c168 ( 72 0 ) capacitor c=0.0199343f //x=23.485 //y=0.865
c169 ( 71 0 ) capacitor c=0.110275f //x=24.02 //y=6.02
c170 ( 70 0 ) capacitor c=0.154305f //x=23.58 //y=6.02
c171 ( 68 0 ) capacitor c=0.00116729f //x=21.05 //y=5.155
c172 ( 67 0 ) capacitor c=0.00226015f //x=20.17 //y=5.155
c173 ( 57 0 ) capacitor c=0.0933903f //x=23.68 //y=2.08
c174 ( 46 0 ) capacitor c=0.0052078f //x=21.43 //y=1.665
c175 ( 45 0 ) capacitor c=0.015794f //x=21.745 //y=1.665
c176 ( 39 0 ) capacitor c=0.0293025f //x=21.745 //y=5.155
c177 ( 31 0 ) capacitor c=0.0184197f //x=20.965 //y=5.155
c178 ( 24 0 ) capacitor c=0.00351598f //x=19.375 //y=5.155
c179 ( 23 0 ) capacitor c=0.0155255f //x=20.085 //y=5.155
c180 ( 7 0 ) capacitor c=0.111457f //x=21.83 //y=2.22
c181 ( 2 0 ) capacitor c=0.0140459f //x=21.945 //y=3.33
c182 ( 1 0 ) capacitor c=0.0669949f //x=23.565 //y=3.33
r183 (  93 95 ) resistor r=20.6867 //w=0.233 //l=0.1 //layer=ply \
 //thickness=0.18 //x=23.58 //y=4.7 //x2=23.68 //y2=4.7
r184 (  86 95 ) resistor r=70.3348 //w=0.233 //l=0.414367 //layer=ply \
 //thickness=0.18 //x=24.02 //y=4.865 //x2=23.68 //y2=4.7
r185 (  85 97 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.015 //y=1.21 //x2=23.975 //y2=1.365
r186 (  84 96 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.015 //y=0.865 //x2=23.975 //y2=0.71
r187 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.015 //y=0.865 //x2=24.015 //y2=1.21
r188 (  82 92 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.64 //y=1.365 //x2=23.525 //y2=1.365
r189 (  81 97 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.86 //y=1.365 //x2=23.975 //y2=1.365
r190 (  80 91 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.64 //y=0.71 //x2=23.525 //y2=0.71
r191 (  79 96 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=23.86 //y=0.71 //x2=23.975 //y2=0.71
r192 (  79 80 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=23.86 //y=0.71 //x2=23.64 //y2=0.71
r193 (  76 93 ) resistor r=13.0941 //w=0.233 //l=0.165 //layer=ply \
 //thickness=0.18 //x=23.58 //y=4.865 //x2=23.58 //y2=4.7
r194 (  75 90 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=23.485 //y=1.915 //x2=23.68 //y2=2.08
r195 (  74 92 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.485 //y=1.52 //x2=23.525 //y2=1.365
r196 (  74 75 ) resistor r=202.543 //w=0.094 //l=0.395 //layer=ply \
 //thickness=0.18 //x=23.485 //y=1.52 //x2=23.485 //y2=1.915
r197 (  73 92 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.485 //y=1.21 //x2=23.525 //y2=1.365
r198 (  72 91 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=23.485 //y=0.865 //x2=23.525 //y2=0.71
r199 (  72 73 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=23.485 //y=0.865 //x2=23.485 //y2=1.21
r200 (  71 86 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=24.02 //y=6.02 //x2=24.02 //y2=4.865
r201 (  70 76 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=23.58 //y=6.02 //x2=23.58 //y2=4.865
r202 (  69 81 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.75 //y=1.365 //x2=23.86 //y2=1.365
r203 (  69 82 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=23.75 //y=1.365 //x2=23.64 //y2=1.365
r204 (  65 95 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=23.68 //y=4.7 //x2=23.68 //y2=4.7
r205 (  57 90 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=23.68 //y=2.08 //x2=23.68 //y2=2.08
r206 (  45 47 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.745 //y=1.665 //x2=21.83 //y2=1.75
r207 (  45 46 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=21.745 //y=1.665 //x2=21.43 //y2=1.665
r208 (  41 46 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.345 //y=1.58 //x2=21.43 //y2=1.665
r209 (  41 98 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=21.345 //y=1.58 //x2=21.345 //y2=1.01
r210 (  40 68 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.135 //y=5.155 //x2=21.05 //y2=5.155
r211 (  39 48 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=21.745 //y=5.155 //x2=21.83 //y2=5.07
r212 (  39 40 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=21.745 //y=5.155 //x2=21.135 //y2=5.155
r213 (  33 68 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=21.05 //y=5.24 //x2=21.05 //y2=5.155
r214 (  33 102 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=21.05 //y=5.24 //x2=21.05 //y2=5.725
r215 (  32 67 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.255 //y=5.155 //x2=20.17 //y2=5.155
r216 (  31 68 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.965 //y=5.155 //x2=21.05 //y2=5.155
r217 (  31 32 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=20.965 //y=5.155 //x2=20.255 //y2=5.155
r218 (  25 67 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.17 //y=5.24 //x2=20.17 //y2=5.155
r219 (  25 101 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=20.17 //y=5.24 //x2=20.17 //y2=5.725
r220 (  23 67 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.085 //y=5.155 //x2=20.17 //y2=5.155
r221 (  23 24 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=20.085 //y=5.155 //x2=19.375 //y2=5.155
r222 (  17 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=19.29 //y=5.24 //x2=19.375 //y2=5.155
r223 (  17 100 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=19.29 //y=5.24 //x2=19.29 //y2=5.725
r224 (  16 65 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=23.68 //y=4.44 //x2=23.68 //y2=4.7
r225 (  15 16 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=23.68 //y=3.33 //x2=23.68 //y2=4.44
r226 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.68 //y=2.96 //x2=23.68 //y2=3.33
r227 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=23.68 //y=2.59 //x2=23.68 //y2=2.96
r228 (  13 57 ) resistor r=34.9091 //w=0.187 //l=0.51 //layer=li \
 //thickness=0.1 //x=23.68 //y=2.59 //x2=23.68 //y2=2.08
r229 (  12 48 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=21.83 //y=4.81 //x2=21.83 //y2=5.07
r230 (  11 12 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.83 //y=4.44 //x2=21.83 //y2=4.81
r231 (  10 11 ) resistor r=75.9786 //w=0.187 //l=1.11 //layer=li \
 //thickness=0.1 //x=21.83 //y=3.33 //x2=21.83 //y2=4.44
r232 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.96 //x2=21.83 //y2=3.33
r233 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=21.83 //y=2.59 //x2=21.83 //y2=2.96
r234 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=21.83 //y=2.22 //x2=21.83 //y2=2.59
r235 (  7 47 ) resistor r=32.1711 //w=0.187 //l=0.47 //layer=li \
 //thickness=0.1 //x=21.83 //y=2.22 //x2=21.83 //y2=1.75
r236 (  6 15 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=23.68 //y=3.33 //x2=23.68 //y2=3.33
r237 (  4 10 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.83 //y=3.33 //x2=21.83 //y2=3.33
r238 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.945 //y=3.33 //x2=21.83 //y2=3.33
r239 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=23.565 //y=3.33 //x2=23.68 //y2=3.33
r240 (  1 2 ) resistor r=1.5458 //w=0.131 //l=1.62 //layer=m1 //thickness=0.36 \
 //x=23.565 //y=3.33 //x2=21.945 //y2=3.33
ends PM_DFFRNX1\%QN

subckt PM_DFFRNX1\%noxref_9 ( 1 2 3 4 5 6 16 23 25 35 36 43 51 57 58 62 63 65 \
 71 72 75 76 77 78 79 80 81 82 83 84 85 86 87 88 90 96 97 98 99 103 104 105 \
 110 112 114 120 121 122 123 124 129 131 133 139 140 150 151 154 163 164 167 \
 175 177 178 179 )
c384 ( 179 0 ) capacitor c=0.023087f //x=16.095 //y=5.02
c385 ( 178 0 ) capacitor c=0.023519f //x=15.215 //y=5.02
c386 ( 177 0 ) capacitor c=0.0224735f //x=14.335 //y=5.02
c387 ( 175 0 ) capacitor c=0.00853354f //x=16.345 //y=0.915
c388 ( 167 0 ) capacitor c=0.0331844f //x=24.45 //y=4.7
c389 ( 164 0 ) capacitor c=0.0279499f //x=24.42 //y=1.915
c390 ( 163 0 ) capacitor c=0.0437302f //x=24.42 //y=2.08
c391 ( 154 0 ) capacitor c=0.0331095f //x=11.5 //y=4.7
c392 ( 151 0 ) capacitor c=0.0279499f //x=11.47 //y=1.915
c393 ( 150 0 ) capacitor c=0.0425269f //x=11.47 //y=2.08
c394 ( 140 0 ) capacitor c=0.0429696f //x=24.985 //y=1.25
c395 ( 139 0 ) capacitor c=0.0192208f //x=24.985 //y=0.905
c396 ( 133 0 ) capacitor c=0.0158629f //x=24.83 //y=1.405
c397 ( 131 0 ) capacitor c=0.0157803f //x=24.83 //y=0.75
c398 ( 129 0 ) capacitor c=0.0306375f //x=24.825 //y=4.79
c399 ( 124 0 ) capacitor c=0.0205163f //x=24.455 //y=1.56
c400 ( 123 0 ) capacitor c=0.0168481f //x=24.455 //y=1.25
c401 ( 122 0 ) capacitor c=0.0174783f //x=24.455 //y=0.905
c402 ( 121 0 ) capacitor c=0.0429696f //x=12.035 //y=1.25
c403 ( 120 0 ) capacitor c=0.0192208f //x=12.035 //y=0.905
c404 ( 114 0 ) capacitor c=0.0148884f //x=11.88 //y=1.405
c405 ( 112 0 ) capacitor c=0.0157803f //x=11.88 //y=0.75
c406 ( 110 0 ) capacitor c=0.0295235f //x=11.875 //y=4.79
c407 ( 105 0 ) capacitor c=0.0205163f //x=11.505 //y=1.56
c408 ( 104 0 ) capacitor c=0.0168481f //x=11.505 //y=1.25
c409 ( 103 0 ) capacitor c=0.0174783f //x=11.505 //y=0.905
c410 ( 99 0 ) capacitor c=0.0559896f //x=1.385 //y=4.79
c411 ( 98 0 ) capacitor c=0.0298189f //x=1.675 //y=4.79
c412 ( 97 0 ) capacitor c=0.0347816f //x=1.34 //y=1.22
c413 ( 96 0 ) capacitor c=0.0187487f //x=1.34 //y=0.875
c414 ( 90 0 ) capacitor c=0.0137055f //x=1.185 //y=1.375
c415 ( 88 0 ) capacitor c=0.0149861f //x=1.185 //y=0.72
c416 ( 87 0 ) capacitor c=0.102158f //x=0.81 //y=1.915
c417 ( 86 0 ) capacitor c=0.0229444f //x=0.81 //y=1.53
c418 ( 85 0 ) capacitor c=0.0234352f //x=0.81 //y=1.22
c419 ( 84 0 ) capacitor c=0.0198724f //x=0.81 //y=0.875
c420 ( 83 0 ) capacitor c=0.15358f //x=24.9 //y=6.02
c421 ( 82 0 ) capacitor c=0.110281f //x=24.46 //y=6.02
c422 ( 81 0 ) capacitor c=0.15358f //x=11.95 //y=6.02
c423 ( 80 0 ) capacitor c=0.110281f //x=11.51 //y=6.02
c424 ( 79 0 ) capacitor c=0.110114f //x=1.75 //y=6.02
c425 ( 78 0 ) capacitor c=0.158956f //x=1.31 //y=6.02
c426 ( 72 0 ) capacitor c=0.00116729f //x=16.24 //y=5.155
c427 ( 71 0 ) capacitor c=0.0021933f //x=15.36 //y=5.155
c428 ( 65 0 ) capacitor c=0.0765697f //x=24.42 //y=2.08
c429 ( 63 0 ) capacitor c=0.00453889f //x=24.42 //y=4.535
c430 ( 62 0 ) capacitor c=0.113069f //x=17.02 //y=4.07
c431 ( 58 0 ) capacitor c=0.00398962f //x=16.62 //y=1.665
c432 ( 57 0 ) capacitor c=0.0137288f //x=16.935 //y=1.665
c433 ( 51 0 ) capacitor c=0.0291076f //x=16.935 //y=5.155
c434 ( 43 0 ) capacitor c=0.0184197f //x=16.155 //y=5.155
c435 ( 36 0 ) capacitor c=0.00332903f //x=14.565 //y=5.155
c436 ( 35 0 ) capacitor c=0.014837f //x=15.275 //y=5.155
c437 ( 25 0 ) capacitor c=0.0719943f //x=11.47 //y=2.08
c438 ( 23 0 ) capacitor c=0.00453889f //x=11.47 //y=4.535
c439 ( 16 0 ) capacitor c=0.124161f //x=1.11 //y=2.08
c440 ( 6 0 ) capacitor c=0.00720076f //x=17.135 //y=4.07
c441 ( 5 0 ) capacitor c=0.228202f //x=24.305 //y=4.07
c442 ( 4 0 ) capacitor c=0.00557292f //x=11.585 //y=4.07
c443 ( 3 0 ) capacitor c=0.0897132f //x=16.905 //y=4.07
c444 ( 2 0 ) capacitor c=0.0160831f //x=1.225 //y=4.07
c445 ( 1 0 ) capacitor c=0.183938f //x=11.355 //y=4.07
r446 (  169 170 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=24.45 //y=4.79 //x2=24.45 //y2=4.865
r447 (  167 169 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=24.45 //y=4.7 //x2=24.45 //y2=4.79
r448 (  163 164 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=24.42 //y=2.08 //x2=24.42 //y2=1.915
r449 (  156 157 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=11.5 //y=4.79 //x2=11.5 //y2=4.865
r450 (  154 156 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=11.5 //y=4.7 //x2=11.5 //y2=4.79
r451 (  150 151 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=11.47 //y=2.08 //x2=11.47 //y2=1.915
r452 (  140 174 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.985 //y=1.25 //x2=24.945 //y2=1.405
r453 (  139 173 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.985 //y=0.905 //x2=24.945 //y2=0.75
r454 (  139 140 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.985 //y=0.905 //x2=24.985 //y2=1.25
r455 (  134 172 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.61 //y=1.405 //x2=24.495 //y2=1.405
r456 (  133 174 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.83 //y=1.405 //x2=24.945 //y2=1.405
r457 (  132 171 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.61 //y=0.75 //x2=24.495 //y2=0.75
r458 (  131 173 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=24.83 //y=0.75 //x2=24.945 //y2=0.75
r459 (  131 132 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=24.83 //y=0.75 //x2=24.61 //y2=0.75
r460 (  130 169 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=24.585 //y=4.79 //x2=24.45 //y2=4.79
r461 (  129 136 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=24.825 //y=4.79 //x2=24.9 //y2=4.865
r462 (  129 130 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=24.825 //y=4.79 //x2=24.585 //y2=4.79
r463 (  124 172 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.455 //y=1.56 //x2=24.495 //y2=1.405
r464 (  124 164 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=24.455 //y=1.56 //x2=24.455 //y2=1.915
r465 (  123 172 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.455 //y=1.25 //x2=24.495 //y2=1.405
r466 (  122 171 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=24.455 //y=0.905 //x2=24.495 //y2=0.75
r467 (  122 123 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=24.455 //y=0.905 //x2=24.455 //y2=1.25
r468 (  121 161 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.035 //y=1.25 //x2=11.995 //y2=1.405
r469 (  120 160 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=12.035 //y=0.905 //x2=11.995 //y2=0.75
r470 (  120 121 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=12.035 //y=0.905 //x2=12.035 //y2=1.25
r471 (  115 159 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.66 //y=1.405 //x2=11.545 //y2=1.405
r472 (  114 161 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.88 //y=1.405 //x2=11.995 //y2=1.405
r473 (  113 158 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.66 //y=0.75 //x2=11.545 //y2=0.75
r474 (  112 160 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=11.88 //y=0.75 //x2=11.995 //y2=0.75
r475 (  112 113 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=11.88 //y=0.75 //x2=11.66 //y2=0.75
r476 (  111 156 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=11.635 //y=4.79 //x2=11.5 //y2=4.79
r477 (  110 117 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=11.875 //y=4.79 //x2=11.95 //y2=4.865
r478 (  110 111 ) resistor r=123.064 //w=0.094 //l=0.24 //layer=ply \
 //thickness=0.18 //x=11.875 //y=4.79 //x2=11.635 //y2=4.79
r479 (  105 159 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.505 //y=1.56 //x2=11.545 //y2=1.405
r480 (  105 151 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=11.505 //y=1.56 //x2=11.505 //y2=1.915
r481 (  104 159 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.505 //y=1.25 //x2=11.545 //y2=1.405
r482 (  103 158 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=11.505 //y=0.905 //x2=11.545 //y2=0.75
r483 (  103 104 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=11.505 //y=0.905 //x2=11.505 //y2=1.25
r484 (  98 100 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.75 //y2=4.865
r485 (  98 99 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.385 //y2=4.79
r486 (  97 148 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=1.22 //x2=1.3 //y2=1.375
r487 (  96 147 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.3 //y2=0.72
r488 (  96 97 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.34 //y2=1.22
r489 (  93 99 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.385 //y2=4.79
r490 (  93 146 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.11 //y2=4.7
r491 (  91 142 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=1.375 //x2=0.85 //y2=1.375
r492 (  90 148 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=1.375 //x2=1.3 //y2=1.375
r493 (  89 141 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=0.72 //x2=0.85 //y2=0.72
r494 (  88 147 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=1.3 //y2=0.72
r495 (  88 89 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=0.965 //y2=0.72
r496 (  87 144 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.915 //x2=1.11 //y2=2.08
r497 (  86 142 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.85 //y2=1.375
r498 (  86 87 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.81 //y2=1.915
r499 (  85 142 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.22 //x2=0.85 //y2=1.375
r500 (  84 141 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.85 //y2=0.72
r501 (  84 85 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.81 //y2=1.22
r502 (  83 136 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=24.9 //y=6.02 //x2=24.9 //y2=4.865
r503 (  82 170 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=24.46 //y=6.02 //x2=24.46 //y2=4.865
r504 (  81 117 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.95 //y=6.02 //x2=11.95 //y2=4.865
r505 (  80 157 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=11.51 //y=6.02 //x2=11.51 //y2=4.865
r506 (  79 100 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.75 //y=6.02 //x2=1.75 //y2=4.865
r507 (  78 93 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.31 //y=6.02 //x2=1.31 //y2=4.865
r508 (  77 133 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=24.72 //y=1.405 //x2=24.83 //y2=1.405
r509 (  77 134 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=24.72 //y=1.405 //x2=24.61 //y2=1.405
r510 (  76 114 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.77 //y=1.405 //x2=11.88 //y2=1.405
r511 (  76 115 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=11.77 //y=1.405 //x2=11.66 //y2=1.405
r512 (  75 90 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=1.185 //y2=1.375
r513 (  75 91 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=0.965 //y2=1.375
r514 (  74 167 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=24.45 //y=4.7 //x2=24.45 //y2=4.7
r515 (  70 154 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.5 //y=4.7 //x2=11.5 //y2=4.7
r516 (  65 163 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=24.42 //y=2.08 //x2=24.42 //y2=2.08
r517 (  65 68 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=24.42 //y=2.08 //x2=24.42 //y2=4.07
r518 (  63 74 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=24.42 //y=4.535 //x2=24.435 //y2=4.7
r519 (  63 68 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=24.42 //y=4.535 //x2=24.42 //y2=4.07
r520 (  60 62 ) resistor r=68.4492 //w=0.187 //l=1 //layer=li //thickness=0.1 \
 //x=17.02 //y=5.07 //x2=17.02 //y2=4.07
r521 (  59 62 ) resistor r=158.802 //w=0.187 //l=2.32 //layer=li \
 //thickness=0.1 //x=17.02 //y=1.75 //x2=17.02 //y2=4.07
r522 (  57 59 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.935 //y=1.665 //x2=17.02 //y2=1.75
r523 (  57 58 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=16.935 //y=1.665 //x2=16.62 //y2=1.665
r524 (  53 58 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.535 //y=1.58 //x2=16.62 //y2=1.665
r525 (  53 175 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=16.535 //y=1.58 //x2=16.535 //y2=1.01
r526 (  52 72 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.325 //y=5.155 //x2=16.24 //y2=5.155
r527 (  51 60 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=16.935 //y=5.155 //x2=17.02 //y2=5.07
r528 (  51 52 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=16.935 //y=5.155 //x2=16.325 //y2=5.155
r529 (  45 72 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.24 //y=5.24 //x2=16.24 //y2=5.155
r530 (  45 179 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=16.24 //y=5.24 //x2=16.24 //y2=5.725
r531 (  44 71 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.445 //y=5.155 //x2=15.36 //y2=5.155
r532 (  43 72 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=16.155 //y=5.155 //x2=16.24 //y2=5.155
r533 (  43 44 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=16.155 //y=5.155 //x2=15.445 //y2=5.155
r534 (  37 71 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.36 //y=5.24 //x2=15.36 //y2=5.155
r535 (  37 178 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=15.36 //y=5.24 //x2=15.36 //y2=5.725
r536 (  35 71 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.275 //y=5.155 //x2=15.36 //y2=5.155
r537 (  35 36 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=15.275 //y=5.155 //x2=14.565 //y2=5.155
r538 (  29 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=14.48 //y=5.24 //x2=14.565 //y2=5.155
r539 (  29 177 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=14.48 //y=5.24 //x2=14.48 //y2=5.725
r540 (  25 150 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=11.47 //y=2.08 //x2=11.47 //y2=2.08
r541 (  25 28 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=11.47 //y=2.08 //x2=11.47 //y2=4.07
r542 (  23 70 ) resistor r=11.4737 //w=0.186 //l=0.172337 //layer=li \
 //thickness=0.1 //x=11.47 //y=4.535 //x2=11.485 //y2=4.7
r543 (  23 28 ) resistor r=31.8289 //w=0.187 //l=0.465 //layer=li \
 //thickness=0.1 //x=11.47 //y=4.535 //x2=11.47 //y2=4.07
r544 (  21 146 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r545 (  19 21 ) resistor r=43.123 //w=0.187 //l=0.63 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.07 //x2=1.11 //y2=4.7
r546 (  16 144 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r547 (  16 19 ) resistor r=136.214 //w=0.187 //l=1.99 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.08 //x2=1.11 //y2=4.07
r548 (  14 68 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=24.42 //y=4.07 //x2=24.42 //y2=4.07
r549 (  12 62 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=17.02 //y=4.07 //x2=17.02 //y2=4.07
r550 (  10 28 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=11.47 //y=4.07 //x2=11.47 //y2=4.07
r551 (  8 19 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.07
r552 (  6 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=17.135 //y=4.07 //x2=17.02 //y2=4.07
r553 (  5 14 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=24.305 //y=4.07 //x2=24.42 //y2=4.07
r554 (  5 6 ) resistor r=6.8416 //w=0.131 //l=7.17 //layer=m1 //thickness=0.36 \
 //x=24.305 //y=4.07 //x2=17.135 //y2=4.07
r555 (  4 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.585 //y=4.07 //x2=11.47 //y2=4.07
r556 (  3 12 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=16.905 //y=4.07 //x2=17.02 //y2=4.07
r557 (  3 4 ) resistor r=5.07634 //w=0.131 //l=5.32 //layer=m1 \
 //thickness=0.36 //x=16.905 //y=4.07 //x2=11.585 //y2=4.07
r558 (  2 8 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=1.225 //y=4.07 //x2=1.11 //y2=4.07
r559 (  1 10 ) resistor r=0.0880901 //w=0.191 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=11.355 //y=4.07 //x2=11.47 //y2=4.07
r560 (  1 2 ) resistor r=9.66603 //w=0.131 //l=10.13 //layer=m1 \
 //thickness=0.36 //x=11.355 //y=4.07 //x2=1.225 //y2=4.07
ends PM_DFFRNX1\%noxref_9

subckt PM_DFFRNX1\%Q ( 1 2 7 8 9 10 11 12 13 14 15 16 17 18 19 20 22 40 41 52 \
 54 55 67 68 69 70 74 75 76 81 83 86 87 89 90 95 98 100 101 )
c144 ( 101 0 ) capacitor c=0.0220291f //x=24.535 //y=5.02
c145 ( 100 0 ) capacitor c=0.0217503f //x=23.655 //y=5.02
c146 ( 98 0 ) capacitor c=0.0084702f //x=24.53 //y=0.905
c147 ( 95 0 ) capacitor c=0.059212f //x=21.09 //y=4.7
c148 ( 90 0 ) capacitor c=0.0273931f //x=21.09 //y=1.915
c149 ( 89 0 ) capacitor c=0.0471168f //x=21.09 //y=2.08
c150 ( 87 0 ) capacitor c=0.0432517f //x=21.61 //y=1.26
c151 ( 86 0 ) capacitor c=0.0200379f //x=21.61 //y=0.915
c152 ( 83 0 ) capacitor c=0.0158629f //x=21.455 //y=1.415
c153 ( 81 0 ) capacitor c=0.0157803f //x=21.455 //y=0.76
c154 ( 76 0 ) capacitor c=0.0218028f //x=21.08 //y=1.57
c155 ( 75 0 ) capacitor c=0.0207459f //x=21.08 //y=1.26
c156 ( 74 0 ) capacitor c=0.0194308f //x=21.08 //y=0.915
c157 ( 70 0 ) capacitor c=0.158794f //x=21.27 //y=6.02
c158 ( 69 0 ) capacitor c=0.110114f //x=20.83 //y=6.02
c159 ( 67 0 ) capacitor c=0.0024826f //x=24.68 //y=5.2
c160 ( 55 0 ) capacitor c=0.00525782f //x=24.805 //y=1.655
c161 ( 54 0 ) capacitor c=0.0140375f //x=25.075 //y=1.655
c162 ( 52 0 ) capacitor c=0.0142754f //x=25.075 //y=5.2
c163 ( 41 0 ) capacitor c=0.00265593f //x=23.885 //y=5.2
c164 ( 40 0 ) capacitor c=0.0150834f //x=24.595 //y=5.2
c165 ( 22 0 ) capacitor c=0.0910244f //x=21.09 //y=2.08
c166 ( 13 0 ) capacitor c=0.128349f //x=25.16 //y=2.22
c167 ( 2 0 ) capacitor c=0.0101384f //x=21.205 //y=3.7
c168 ( 1 0 ) capacitor c=0.102069f //x=25.045 //y=3.7
r169 (  89 90 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=21.09 //y=2.08 //x2=21.09 //y2=1.915
r170 (  87 97 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.61 //y=1.26 //x2=21.57 //y2=1.415
r171 (  86 96 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.61 //y=0.915 //x2=21.57 //y2=0.76
r172 (  86 87 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=21.61 //y=0.915 //x2=21.61 //y2=1.26
r173 (  84 93 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.235 //y=1.415 //x2=21.12 //y2=1.415
r174 (  83 97 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.455 //y=1.415 //x2=21.57 //y2=1.415
r175 (  82 92 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.235 //y=0.76 //x2=21.12 //y2=0.76
r176 (  81 96 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=21.455 //y=0.76 //x2=21.57 //y2=0.76
r177 (  81 82 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=21.455 //y=0.76 //x2=21.235 //y2=0.76
r178 (  78 95 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=21.27 //y=4.865 //x2=21.09 //y2=4.7
r179 (  76 93 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.08 //y=1.57 //x2=21.12 //y2=1.415
r180 (  76 90 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=21.08 //y=1.57 //x2=21.08 //y2=1.915
r181 (  75 93 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.08 //y=1.26 //x2=21.12 //y2=1.415
r182 (  74 92 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=21.08 //y=0.915 //x2=21.12 //y2=0.76
r183 (  74 75 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=21.08 //y=0.915 //x2=21.08 //y2=1.26
r184 (  71 95 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=20.83 //y=4.865 //x2=21.09 //y2=4.7
r185 (  70 78 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=21.27 //y=6.02 //x2=21.27 //y2=4.865
r186 (  69 71 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=20.83 //y=6.02 //x2=20.83 //y2=4.865
r187 (  68 83 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=21.345 //y=1.415 //x2=21.455 //y2=1.415
r188 (  68 84 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=21.345 //y=1.415 //x2=21.235 //y2=1.415
r189 (  54 56 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.075 //y=1.655 //x2=25.16 //y2=1.74
r190 (  54 55 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=25.075 //y=1.655 //x2=24.805 //y2=1.655
r191 (  53 67 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.765 //y=5.2 //x2=24.68 //y2=5.2
r192 (  52 57 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=25.075 //y=5.2 //x2=25.16 //y2=5.115
r193 (  52 53 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=25.075 //y=5.2 //x2=24.765 //y2=5.2
r194 (  48 55 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=24.72 //y=1.57 //x2=24.805 //y2=1.655
r195 (  48 98 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=24.72 //y=1.57 //x2=24.72 //y2=1
r196 (  42 67 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.68 //y=5.285 //x2=24.68 //y2=5.2
r197 (  42 101 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=24.68 //y=5.285 //x2=24.68 //y2=5.725
r198 (  40 67 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=24.595 //y=5.2 //x2=24.68 //y2=5.2
r199 (  40 41 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=24.595 //y=5.2 //x2=23.885 //y2=5.2
r200 (  34 41 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=23.8 //y=5.285 //x2=23.885 //y2=5.2
r201 (  34 100 ) resistor r=30.1176 //w=0.187 //l=0.44 //layer=li \
 //thickness=0.1 //x=23.8 //y=5.285 //x2=23.8 //y2=5.725
r202 (  32 95 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.09 //y=4.7 //x2=21.09 //y2=4.7
r203 (  22 89 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=21.09 //y=2.08 //x2=21.09 //y2=2.08
r204 (  20 57 ) resistor r=20.877 //w=0.187 //l=0.305 //layer=li \
 //thickness=0.1 //x=25.16 //y=4.81 //x2=25.16 //y2=5.115
r205 (  19 20 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=25.16 //y=4.44 //x2=25.16 //y2=4.81
r206 (  18 19 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=25.16 //y=4.07 //x2=25.16 //y2=4.44
r207 (  17 18 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=25.16 //y=3.7 //x2=25.16 //y2=4.07
r208 (  16 17 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=25.16 //y=3.33 //x2=25.16 //y2=3.7
r209 (  15 16 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=25.16 //y=2.96 //x2=25.16 //y2=3.33
r210 (  14 15 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=25.16 //y=2.59 //x2=25.16 //y2=2.96
r211 (  13 14 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=25.16 //y=2.22 //x2=25.16 //y2=2.59
r212 (  13 56 ) resistor r=32.8556 //w=0.187 //l=0.48 //layer=li \
 //thickness=0.1 //x=25.16 //y=2.22 //x2=25.16 //y2=1.74
r213 (  12 32 ) resistor r=17.7968 //w=0.187 //l=0.26 //layer=li \
 //thickness=0.1 //x=21.09 //y=4.44 //x2=21.09 //y2=4.7
r214 (  11 12 ) resistor r=50.6524 //w=0.187 //l=0.74 //layer=li \
 //thickness=0.1 //x=21.09 //y=3.7 //x2=21.09 //y2=4.44
r215 (  10 11 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.09 //y=3.33 //x2=21.09 //y2=3.7
r216 (  9 10 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li \
 //thickness=0.1 //x=21.09 //y=2.96 //x2=21.09 //y2=3.33
r217 (  8 9 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=21.09 //y=2.59 //x2=21.09 //y2=2.96
r218 (  7 8 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=21.09 //y=2.22 //x2=21.09 //y2=2.59
r219 (  7 22 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=21.09 //y=2.22 //x2=21.09 //y2=2.08
r220 (  6 17 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=25.16 //y=3.7 //x2=25.16 //y2=3.7
r221 (  4 11 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=21.09 //y=3.7 //x2=21.09 //y2=3.7
r222 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=21.205 //y=3.7 //x2=21.09 //y2=3.7
r223 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=25.045 //y=3.7 //x2=25.16 //y2=3.7
r224 (  1 2 ) resistor r=3.66412 //w=0.131 //l=3.84 //layer=m1 \
 //thickness=0.36 //x=25.045 //y=3.7 //x2=21.205 //y2=3.7
ends PM_DFFRNX1\%Q

subckt PM_DFFRNX1\%noxref_11 ( 1 5 9 13 17 35 )
c47 ( 35 0 ) capacitor c=0.0703709f //x=0.455 //y=0.375
c48 ( 17 0 ) capacitor c=0.0221229f //x=2.445 //y=1.59
c49 ( 13 0 ) capacitor c=0.0156939f //x=2.445 //y=0.54
c50 ( 9 0 ) capacitor c=0.00678203f //x=1.56 //y=0.625
c51 ( 5 0 ) capacitor c=0.0206412f //x=1.475 //y=1.59
c52 ( 1 0 ) capacitor c=0.0109947f //x=0.59 //y=1.505
r53 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=1.59 //x2=1.56 //y2=1.63
r54 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=1.59 //x2=2.045 //y2=1.59
r55 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=1.59 //x2=2.53 //y2=1.59
r56 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=1.59 //x2=2.045 //y2=1.59
r57 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=0.54 //x2=1.56 //y2=0.5
r58 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=0.54 //x2=2.045 //y2=0.54
r59 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=0.54 //x2=2.53 //y2=0.54
r60 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=0.54 //x2=2.045 //y2=0.54
r61 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=1.63
r62 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=0.89
r63 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.5
r64 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.89
r65 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.675 //y=1.59 //x2=0.59 //y2=1.63
r66 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.675 //y=1.59 //x2=1.075 //y2=1.59
r67 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.475 //y=1.59 //x2=1.56 //y2=1.63
r68 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.475 //y=1.59 //x2=1.075 //y2=1.59
r69 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.59 //y=1.505 //x2=0.59 //y2=1.63
r70 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.59 //y=1.505 //x2=0.59 //y2=0.89
ends PM_DFFRNX1\%noxref_11

subckt PM_DFFRNX1\%noxref_12 ( 1 3 11 15 25 28 29 )
c53 ( 29 0 ) capacitor c=0.043074f //x=2.965 //y=0.375
c54 ( 28 0 ) capacitor c=0.00465142f //x=1.86 //y=0.91
c55 ( 25 0 ) capacitor c=0.00156479f //x=3.1 //y=0.995
c56 ( 15 0 ) capacitor c=0.00737666f //x=4.07 //y=0.625
c57 ( 11 0 ) capacitor c=0.0149771f //x=3.985 //y=0.54
c58 ( 3 0 ) capacitor c=0.00718386f //x=3.1 //y=0.625
c59 ( 1 0 ) capacitor c=0.0253322f //x=3.015 //y=0.995
r60 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.5
r61 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.89
r62 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.185 //y=0.54 //x2=3.1 //y2=0.5
r63 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.185 //y=0.54 //x2=3.585 //y2=0.54
r64 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.985 //y=0.54 //x2=4.07 //y2=0.5
r65 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.985 //y=0.54 //x2=3.585 //y2=0.54
r66 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=0.995
r67 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=1.23
r68 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.995
r69 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.89
r70 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.5
r71 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.89
r72 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.135 //y=0.995 //x2=2.05 //y2=0.995
r73 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=3.1 //y2=0.995
r74 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=2.135 //y2=0.995
ends PM_DFFRNX1\%noxref_12

subckt PM_DFFRNX1\%D ( 1 2 3 5 13 14 15 16 17 18 20 26 27 28 29 30 38 )
c80 ( 38 0 ) capacitor c=0.0335551f //x=7.03 //y=4.7
c81 ( 30 0 ) capacitor c=0.0245352f //x=7.365 //y=4.79
c82 ( 29 0 ) capacitor c=0.0850619f //x=7.12 //y=1.915
c83 ( 28 0 ) capacitor c=0.0170266f //x=7.12 //y=1.45
c84 ( 27 0 ) capacitor c=0.018609f //x=7.12 //y=1.22
c85 ( 26 0 ) capacitor c=0.0187309f //x=7.12 //y=0.91
c86 ( 20 0 ) capacitor c=0.014725f //x=6.965 //y=1.375
c87 ( 18 0 ) capacitor c=0.0146567f //x=6.965 //y=0.755
c88 ( 17 0 ) capacitor c=0.0335408f //x=6.595 //y=1.22
c89 ( 16 0 ) capacitor c=0.0173761f //x=6.595 //y=0.91
c90 ( 15 0 ) capacitor c=0.110114f //x=7.44 //y=6.02
c91 ( 14 0 ) capacitor c=0.11012f //x=7 //y=6.02
c92 ( 5 0 ) capacitor c=0.0956955f //x=7.03 //y=2.08
r93 (  40 41 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=7.03 //y=4.79 //x2=7.03 //y2=4.865
r94 (  38 40 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=7.03 //y=4.7 //x2=7.03 //y2=4.79
r95 (  31 40 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=7.165 //y=4.79 //x2=7.03 //y2=4.79
r96 (  30 32 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=7.365 //y=4.79 //x2=7.44 //y2=4.865
r97 (  30 31 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=7.365 //y=4.79 //x2=7.165 //y2=4.79
r98 (  29 45 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.915 //x2=7.045 //y2=2.08
r99 (  28 43 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.45 //x2=7.08 //y2=1.375
r100 (  28 29 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.45 //x2=7.12 //y2=1.915
r101 (  27 43 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.12 //y=1.22 //x2=7.08 //y2=1.375
r102 (  26 42 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=7.12 //y=0.91 //x2=7.08 //y2=0.755
r103 (  26 27 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=7.12 //y=0.91 //x2=7.12 //y2=1.22
r104 (  21 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.75 //y=1.375 //x2=6.635 //y2=1.375
r105 (  20 43 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.965 //y=1.375 //x2=7.08 //y2=1.375
r106 (  19 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.75 //y=0.755 //x2=6.635 //y2=0.755
r107 (  18 42 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.965 //y=0.755 //x2=7.08 //y2=0.755
r108 (  18 19 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=6.965 //y=0.755 //x2=6.75 //y2=0.755
r109 (  17 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.595 //y=1.22 //x2=6.635 //y2=1.375
r110 (  16 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.595 //y=0.91 //x2=6.635 //y2=0.755
r111 (  16 17 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=6.595 //y=0.91 //x2=6.595 //y2=1.22
r112 (  15 32 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7.44 //y=6.02 //x2=7.44 //y2=4.865
r113 (  14 41 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=7 //y=6.02 //x2=7 //y2=4.865
r114 (  13 20 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=6.857 //y=1.375 //x2=6.965 //y2=1.375
r115 (  13 21 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=6.857 //y=1.375 //x2=6.75 //y2=1.375
r116 (  11 38 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.03 //y=4.7 //x2=7.03 //y2=4.7
r117 (  5 45 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=7.03 //y=2.08 //x2=7.03 //y2=2.08
r118 (  3 11 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=7.03 //y=2.96 //x2=7.03 //y2=4.7
r119 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=7.03 //y=2.59 //x2=7.03 //y2=2.96
r120 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=7.03 //y=2.22 //x2=7.03 //y2=2.59
r121 (  1 5 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li //thickness=0.1 \
 //x=7.03 //y=2.22 //x2=7.03 //y2=2.08
ends PM_DFFRNX1\%D

subckt PM_DFFRNX1\%noxref_14 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0693021f //x=5.265 //y=0.375
c51 ( 17 0 ) capacitor c=0.0206235f //x=7.255 //y=1.59
c52 ( 13 0 ) capacitor c=0.0156174f //x=7.255 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=6.37 //y=0.625
c54 ( 5 0 ) capacitor c=0.0183576f //x=6.285 //y=1.59
c55 ( 1 0 ) capacitor c=0.00791969f //x=5.4 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.455 //y=1.59 //x2=6.37 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.455 //y=1.59 //x2=6.855 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.255 //y=1.59 //x2=7.34 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.255 //y=1.59 //x2=6.855 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.455 //y=0.54 //x2=6.37 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.455 //y=0.54 //x2=6.855 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=7.255 //y=0.54 //x2=7.34 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.255 //y=0.54 //x2=6.855 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=6.37 //y=1.505 //x2=6.37 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=6.37 //y=1.505 //x2=6.37 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=6.37 //y=0.625 //x2=6.37 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=6.37 //y=0.625 //x2=6.37 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=5.485 //y=1.59 //x2=5.4 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=5.485 //y=1.59 //x2=5.885 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=6.285 //y=1.59 //x2=6.37 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=6.285 //y=1.59 //x2=5.885 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=5.4 //y=1.505 //x2=5.4 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=5.4 //y=1.505 //x2=5.4 //y2=0.89
ends PM_DFFRNX1\%noxref_14

subckt PM_DFFRNX1\%noxref_15 ( 1 3 11 15 25 28 29 )
c54 ( 29 0 ) capacitor c=0.0423432f //x=7.775 //y=0.375
c55 ( 28 0 ) capacitor c=0.00463374f //x=6.67 //y=0.91
c56 ( 25 0 ) capacitor c=0.00156479f //x=7.91 //y=0.995
c57 ( 15 0 ) capacitor c=0.00737666f //x=8.88 //y=0.625
c58 ( 11 0 ) capacitor c=0.0144218f //x=8.795 //y=0.54
c59 ( 3 0 ) capacitor c=0.00718386f //x=7.91 //y=0.625
c60 ( 1 0 ) capacitor c=0.0242666f //x=7.825 //y=0.995
r61 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=8.88 //y=0.625 //x2=8.88 //y2=0.5
r62 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=8.88 //y=0.625 //x2=8.88 //y2=0.89
r63 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=7.995 //y=0.54 //x2=7.91 //y2=0.5
r64 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=7.995 //y=0.54 //x2=8.395 //y2=0.54
r65 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=8.795 //y=0.54 //x2=8.88 //y2=0.5
r66 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=8.795 //y=0.54 //x2=8.395 //y2=0.54
r67 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.91 //y=1.08 //x2=7.91 //y2=0.995
r68 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=7.91 //y=1.08 //x2=7.91 //y2=1.23
r69 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.91 //x2=7.91 //y2=0.995
r70 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.91 //x2=7.91 //y2=0.89
r71 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.625 //x2=7.91 //y2=0.5
r72 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=7.91 //y=0.625 //x2=7.91 //y2=0.89
r73 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.945 //y=0.995 //x2=6.86 //y2=0.995
r74 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=7.825 //y=0.995 //x2=7.91 //y2=0.995
r75 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=7.825 //y=0.995 //x2=6.945 //y2=0.995
ends PM_DFFRNX1\%noxref_15

subckt PM_DFFRNX1\%noxref_16 ( 1 5 9 10 13 17 29 )
c52 ( 29 0 ) capacitor c=0.0632682f //x=10.18 //y=0.365
c53 ( 17 0 ) capacitor c=0.0072343f //x=12.255 //y=0.615
c54 ( 13 0 ) capacitor c=0.0145084f //x=12.17 //y=0.53
c55 ( 10 0 ) capacitor c=0.00582081f //x=11.285 //y=1.495
c56 ( 9 0 ) capacitor c=0.006761f //x=11.285 //y=0.615
c57 ( 5 0 ) capacitor c=0.0173046f //x=11.2 //y=1.58
c58 ( 1 0 ) capacitor c=0.00733328f //x=10.315 //y=1.495
r59 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=12.255 //y=0.615 //x2=12.255 //y2=0.49
r60 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=12.255 //y=0.615 //x2=12.255 //y2=0.88
r61 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.37 //y=0.53 //x2=11.285 //y2=0.49
r62 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.37 //y=0.53 //x2=11.77 //y2=0.53
r63 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=12.17 //y=0.53 //x2=12.255 //y2=0.49
r64 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=12.17 //y=0.53 //x2=11.77 //y2=0.53
r65 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=11.285 //y=1.495 //x2=11.285 //y2=1.62
r66 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=11.285 //y=1.495 //x2=11.285 //y2=0.88
r67 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=11.285 //y=0.615 //x2=11.285 //y2=0.49
r68 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=11.285 //y=0.615 //x2=11.285 //y2=0.88
r69 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=10.4 //y=1.58 //x2=10.315 //y2=1.62
r70 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=10.4 //y=1.58 //x2=10.8 //y2=1.58
r71 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=11.2 //y=1.58 //x2=11.285 //y2=1.62
r72 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=11.2 //y=1.58 //x2=10.8 //y2=1.58
r73 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=10.315 //y=1.495 //x2=10.315 //y2=1.62
r74 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=10.315 //y=1.495 //x2=10.315 //y2=0.88
ends PM_DFFRNX1\%noxref_16

subckt PM_DFFRNX1\%noxref_17 ( 1 5 9 13 17 35 )
c50 ( 35 0 ) capacitor c=0.0673029f //x=13.405 //y=0.375
c51 ( 17 0 ) capacitor c=0.0178317f //x=15.395 //y=1.59
c52 ( 13 0 ) capacitor c=0.0154936f //x=15.395 //y=0.54
c53 ( 9 0 ) capacitor c=0.00678203f //x=14.51 //y=0.625
c54 ( 5 0 ) capacitor c=0.0164013f //x=14.425 //y=1.59
c55 ( 1 0 ) capacitor c=0.00696517f //x=13.54 //y=1.505
r56 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.595 //y=1.59 //x2=14.51 //y2=1.63
r57 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.595 //y=1.59 //x2=14.995 //y2=1.59
r58 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.395 //y=1.59 //x2=15.48 //y2=1.59
r59 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.395 //y=1.59 //x2=14.995 //y2=1.59
r60 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.595 //y=0.54 //x2=14.51 //y2=0.5
r61 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.595 //y=0.54 //x2=14.995 //y2=0.54
r62 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.395 //y=0.54 //x2=15.48 //y2=0.54
r63 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=15.395 //y=0.54 //x2=14.995 //y2=0.54
r64 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=14.51 //y=1.505 //x2=14.51 //y2=1.63
r65 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=14.51 //y=1.505 //x2=14.51 //y2=0.89
r66 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=14.51 //y=0.625 //x2=14.51 //y2=0.5
r67 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=14.51 //y=0.625 //x2=14.51 //y2=0.89
r68 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=13.625 //y=1.59 //x2=13.54 //y2=1.63
r69 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=13.625 //y=1.59 //x2=14.025 //y2=1.59
r70 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=14.425 //y=1.59 //x2=14.51 //y2=1.63
r71 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=14.425 //y=1.59 //x2=14.025 //y2=1.59
r72 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=13.54 //y=1.505 //x2=13.54 //y2=1.63
r73 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=13.54 //y=1.505 //x2=13.54 //y2=0.89
ends PM_DFFRNX1\%noxref_17

subckt PM_DFFRNX1\%noxref_18 ( 1 3 11 15 25 28 29 )
c54 ( 29 0 ) capacitor c=0.0413887f //x=15.915 //y=0.375
c55 ( 28 0 ) capacitor c=0.0045748f //x=14.81 //y=0.91
c56 ( 25 0 ) capacitor c=0.00156479f //x=16.05 //y=0.995
c57 ( 15 0 ) capacitor c=0.00737666f //x=17.02 //y=0.625
c58 ( 11 0 ) capacitor c=0.0144218f //x=16.935 //y=0.54
c59 ( 3 0 ) capacitor c=0.00718386f //x=16.05 //y=0.625
c60 ( 1 0 ) capacitor c=0.0220678f //x=15.965 //y=0.995
r61 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=17.02 //y=0.625 //x2=17.02 //y2=0.5
r62 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=17.02 //y=0.625 //x2=17.02 //y2=0.89
r63 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.135 //y=0.54 //x2=16.05 //y2=0.5
r64 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.135 //y=0.54 //x2=16.535 //y2=0.54
r65 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=16.935 //y=0.54 //x2=17.02 //y2=0.5
r66 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=16.935 //y=0.54 //x2=16.535 //y2=0.54
r67 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=16.05 //y=1.08 //x2=16.05 //y2=0.995
r68 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=16.05 //y=1.08 //x2=16.05 //y2=1.23
r69 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=16.05 //y=0.91 //x2=16.05 //y2=0.995
r70 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=16.05 //y=0.91 //x2=16.05 //y2=0.89
r71 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=16.05 //y=0.625 //x2=16.05 //y2=0.5
r72 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=16.05 //y=0.625 //x2=16.05 //y2=0.89
r73 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=15.085 //y=0.995 //x2=15 //y2=0.995
r74 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=15.965 //y=0.995 //x2=16.05 //y2=0.995
r75 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=15.965 //y=0.995 //x2=15.085 //y2=0.995
ends PM_DFFRNX1\%noxref_18

subckt PM_DFFRNX1\%noxref_19 ( 1 5 9 13 17 35 )
c52 ( 35 0 ) capacitor c=0.0688914f //x=18.215 //y=0.375
c53 ( 17 0 ) capacitor c=0.018313f //x=20.205 //y=1.59
c54 ( 13 0 ) capacitor c=0.0155692f //x=20.205 //y=0.54
c55 ( 9 0 ) capacitor c=0.00678203f //x=19.32 //y=0.625
c56 ( 5 0 ) capacitor c=0.0164013f //x=19.235 //y=1.59
c57 ( 1 0 ) capacitor c=0.00696517f //x=18.35 //y=1.505
r58 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.405 //y=1.59 //x2=19.32 //y2=1.63
r59 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.405 //y=1.59 //x2=19.805 //y2=1.59
r60 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.205 //y=1.59 //x2=20.29 //y2=1.59
r61 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.205 //y=1.59 //x2=19.805 //y2=1.59
r62 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.405 //y=0.54 //x2=19.32 //y2=0.5
r63 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.405 //y=0.54 //x2=19.805 //y2=0.54
r64 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=20.205 //y=0.54 //x2=20.29 //y2=0.54
r65 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.205 //y=0.54 //x2=19.805 //y2=0.54
r66 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=19.32 //y=1.505 //x2=19.32 //y2=1.63
r67 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=19.32 //y=1.505 //x2=19.32 //y2=0.89
r68 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=19.32 //y=0.625 //x2=19.32 //y2=0.5
r69 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=19.32 //y=0.625 //x2=19.32 //y2=0.89
r70 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=18.435 //y=1.59 //x2=18.35 //y2=1.63
r71 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=18.435 //y=1.59 //x2=18.835 //y2=1.59
r72 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=19.235 //y=1.59 //x2=19.32 //y2=1.63
r73 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=19.235 //y=1.59 //x2=18.835 //y2=1.59
r74 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=18.35 //y=1.505 //x2=18.35 //y2=1.63
r75 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=18.35 //y=1.505 //x2=18.35 //y2=0.89
ends PM_DFFRNX1\%noxref_19

subckt PM_DFFRNX1\%noxref_20 ( 1 3 11 15 25 28 29 )
c52 ( 29 0 ) capacitor c=0.0430705f //x=20.725 //y=0.375
c53 ( 28 0 ) capacitor c=0.00457437f //x=19.62 //y=0.91
c54 ( 25 0 ) capacitor c=0.00156479f //x=20.86 //y=0.995
c55 ( 15 0 ) capacitor c=0.00737666f //x=21.83 //y=0.625
c56 ( 11 0 ) capacitor c=0.0152164f //x=21.745 //y=0.54
c57 ( 3 0 ) capacitor c=0.00718386f //x=20.86 //y=0.625
c58 ( 1 0 ) capacitor c=0.0252837f //x=20.775 //y=0.995
r59 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=21.83 //y=0.625 //x2=21.83 //y2=0.5
r60 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=21.83 //y=0.625 //x2=21.83 //y2=0.89
r61 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=20.945 //y=0.54 //x2=20.86 //y2=0.5
r62 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=20.945 //y=0.54 //x2=21.345 //y2=0.54
r63 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=21.745 //y=0.54 //x2=21.83 //y2=0.5
r64 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=21.745 //y=0.54 //x2=21.345 //y2=0.54
r65 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.86 //y=1.08 //x2=20.86 //y2=0.995
r66 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=20.86 //y=1.08 //x2=20.86 //y2=1.23
r67 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.86 //y=0.91 //x2=20.86 //y2=0.995
r68 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=20.86 //y=0.91 //x2=20.86 //y2=0.89
r69 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=20.86 //y=0.625 //x2=20.86 //y2=0.5
r70 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=20.86 //y=0.625 //x2=20.86 //y2=0.89
r71 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=19.895 //y=0.995 //x2=19.81 //y2=0.995
r72 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=20.775 //y=0.995 //x2=20.86 //y2=0.995
r73 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=20.775 //y=0.995 //x2=19.895 //y2=0.995
ends PM_DFFRNX1\%noxref_20

subckt PM_DFFRNX1\%noxref_21 ( 1 5 9 10 13 17 29 )
c50 ( 29 0 ) capacitor c=0.0637432f //x=23.13 //y=0.365
c51 ( 17 0 ) capacitor c=0.00722223f //x=25.205 //y=0.615
c52 ( 13 0 ) capacitor c=0.0149664f //x=25.12 //y=0.53
c53 ( 10 0 ) capacitor c=0.00687696f //x=24.235 //y=1.495
c54 ( 9 0 ) capacitor c=0.006761f //x=24.235 //y=0.615
c55 ( 5 0 ) capacitor c=0.0201208f //x=24.15 //y=1.58
c56 ( 1 0 ) capacitor c=0.00828748f //x=23.265 //y=1.495
r57 (  17 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=25.205 //y=0.615 //x2=25.205 //y2=0.49
r58 (  17 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=25.205 //y=0.615 //x2=25.205 //y2=0.88
r59 (  14 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=24.32 //y=0.53 //x2=24.235 //y2=0.49
r60 (  14 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=24.32 //y=0.53 //x2=24.72 //y2=0.53
r61 (  13 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=25.12 //y=0.53 //x2=25.205 //y2=0.49
r62 (  13 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=25.12 //y=0.53 //x2=24.72 //y2=0.53
r63 (  10 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=24.235 //y=1.495 //x2=24.235 //y2=1.62
r64 (  10 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=24.235 //y=1.495 //x2=24.235 //y2=0.88
r65 (  9 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=24.235 //y=0.615 //x2=24.235 //y2=0.49
r66 (  9 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=24.235 //y=0.615 //x2=24.235 //y2=0.88
r67 (  6 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=23.35 //y=1.58 //x2=23.265 //y2=1.62
r68 (  6 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=23.35 //y=1.58 //x2=23.75 //y2=1.58
r69 (  5 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=24.15 //y=1.58 //x2=24.235 //y2=1.62
r70 (  5 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=24.15 //y=1.58 //x2=23.75 //y2=1.58
r71 (  1 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=23.265 //y=1.495 //x2=23.265 //y2=1.62
r72 (  1 29 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=23.265 //y=1.495 //x2=23.265 //y2=0.88
ends PM_DFFRNX1\%noxref_21

