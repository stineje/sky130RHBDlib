// File: OR2X1.spi.pex
// Created: Tue Oct 15 15:50:42 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_OR2X1\%GND ( 1 13 25 29 37 41 49 55 63 67 78 81 100 112 113 )
c74 ( 113 0 ) capacitor c=0.0600324f //x=3.825 //y=0.37
c75 ( 112 0 ) capacitor c=0.0737024f //x=0.56 //y=0.365
c76 ( 100 0 ) capacitor c=0.0992376f //x=3.33 //y=0
c77 ( 81 0 ) capacitor c=0.202778f //x=0.695 //y=0
c78 ( 78 0 ) capacitor c=0.198211f //x=5.18 //y=0
c79 ( 76 0 ) capacitor c=0.0360689f //x=5.015 //y=0
c80 ( 70 0 ) capacitor c=0.00587411f //x=4.93 //y=0.45
c81 ( 67 0 ) capacitor c=0.00542558f //x=4.845 //y=0.535
c82 ( 66 0 ) capacitor c=0.00479856f //x=4.445 //y=0.45
c83 ( 63 0 ) capacitor c=0.0068422f //x=4.36 //y=0.535
c84 ( 58 0 ) capacitor c=0.00592191f //x=3.96 //y=0.45
c85 ( 55 0 ) capacitor c=0.0164879f //x=3.875 //y=0
c86 ( 50 0 ) capacitor c=0.0659516f //x=2.72 //y=0
c87 ( 49 0 ) capacitor c=0.0195795f //x=3.16 //y=0
c88 ( 44 0 ) capacitor c=0.00609805f //x=2.635 //y=0.445
c89 ( 41 0 ) capacitor c=0.00508468f //x=2.55 //y=0.53
c90 ( 40 0 ) capacitor c=0.00468234f //x=2.15 //y=0.445
c91 ( 37 0 ) capacitor c=0.00556167f //x=2.065 //y=0.53
c92 ( 32 0 ) capacitor c=0.00468234f //x=1.665 //y=0.445
c93 ( 29 0 ) capacitor c=0.00556167f //x=1.58 //y=0.53
c94 ( 28 0 ) capacitor c=0.00468234f //x=1.18 //y=0.445
c95 ( 25 0 ) capacitor c=0.00709092f //x=1.095 //y=0.53
c96 ( 20 0 ) capacitor c=0.00609805f //x=0.695 //y=0.445
c97 ( 13 0 ) capacitor c=0.224767f //x=5.18 //y=0
r98 (  104 105 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=4.445 //y=0 //x2=4.93 //y2=0
r99 (  103 104 ) resistor r=0.179272 //w=0.357 //l=0.005 //layer=li \
 //thickness=0.1 //x=4.44 //y=0 //x2=4.445 //y2=0
r100 (  101 103 ) resistor r=17.2101 //w=0.357 //l=0.48 //layer=li \
 //thickness=0.1 //x=3.96 //y=0 //x2=4.44 //y2=0
r101 (  88 89 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.15 //y=0 //x2=2.635 //y2=0
r102 (  87 88 ) resistor r=10.7563 //w=0.357 //l=0.3 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.15 //y2=0
r103 (  85 87 ) resistor r=6.63305 //w=0.357 //l=0.185 //layer=li \
 //thickness=0.1 //x=1.665 //y=0 //x2=1.85 //y2=0
r104 (  84 85 ) resistor r=17.3894 //w=0.357 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.18 //y=0 //x2=1.665 //y2=0
r105 (  83 84 ) resistor r=15.7759 //w=0.357 //l=0.44 //layer=li \
 //thickness=0.1 //x=0.74 //y=0 //x2=1.18 //y2=0
r106 (  81 83 ) resistor r=1.61345 //w=0.357 //l=0.045 //layer=li \
 //thickness=0.1 //x=0.695 //y=0 //x2=0.74 //y2=0
r107 (  76 105 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.015 //y=0 //x2=4.93 //y2=0
r108 (  76 78 ) resistor r=5.91597 //w=0.357 //l=0.165 //layer=li \
 //thickness=0.1 //x=5.015 //y=0 //x2=5.18 //y2=0
r109 (  71 113 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.62 //x2=4.93 //y2=0.535
r110 (  71 113 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.62 //x2=4.93 //y2=1.225
r111 (  70 113 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.45 //x2=4.93 //y2=0.535
r112 (  69 105 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.17 //x2=4.93 //y2=0
r113 (  69 70 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=4.93 //y=0.17 //x2=4.93 //y2=0.45
r114 (  68 113 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.53 //y=0.535 //x2=4.445 //y2=0.535
r115 (  67 113 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.845 //y=0.535 //x2=4.93 //y2=0.535
r116 (  67 68 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=4.845 //y=0.535 //x2=4.53 //y2=0.535
r117 (  66 113 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.445 //y=0.45 //x2=4.445 //y2=0.535
r118 (  65 104 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=4.445 //y=0.17 //x2=4.445 //y2=0
r119 (  65 66 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=4.445 //y=0.17 //x2=4.445 //y2=0.45
r120 (  64 113 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.045 //y=0.535 //x2=3.96 //y2=0.535
r121 (  63 113 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.36 //y=0.535 //x2=4.445 //y2=0.535
r122 (  63 64 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=4.36 //y=0.535 //x2=4.045 //y2=0.535
r123 (  59 113 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.62 //x2=3.96 //y2=0.535
r124 (  59 113 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.62 //x2=3.96 //y2=1.225
r125 (  58 113 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.45 //x2=3.96 //y2=0.535
r126 (  57 101 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.17 //x2=3.96 //y2=0
r127 (  57 58 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=3.96 //y=0.17 //x2=3.96 //y2=0.45
r128 (  56 100 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.5 //y=0 //x2=3.33 //y2=0
r129 (  55 101 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.875 //y=0 //x2=3.96 //y2=0
r130 (  55 56 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=3.875 //y=0 //x2=3.5 //y2=0
r131 (  50 89 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.72 //y=0 //x2=2.635 //y2=0
r132 (  50 52 ) resistor r=8.60504 //w=0.357 //l=0.24 //layer=li \
 //thickness=0.1 //x=2.72 //y=0 //x2=2.96 //y2=0
r133 (  49 100 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=3.33 //y2=0
r134 (  49 52 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=0 //x2=2.96 //y2=0
r135 (  45 112 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.53
r136 (  45 112 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.615 //x2=2.635 //y2=0.88
r137 (  44 112 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.445 //x2=2.635 //y2=0.53
r138 (  43 89 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.17 //x2=2.635 //y2=0
r139 (  43 44 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=2.635 //y=0.17 //x2=2.635 //y2=0.445
r140 (  42 112 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.235 //y=0.53 //x2=2.15 //y2=0.53
r141 (  41 112 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.635 //y2=0.53
r142 (  41 42 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=2.55 //y=0.53 //x2=2.235 //y2=0.53
r143 (  40 112 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.445 //x2=2.15 //y2=0.53
r144 (  39 88 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.17 //x2=2.15 //y2=0
r145 (  39 40 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=2.15 //y=0.17 //x2=2.15 //y2=0.445
r146 (  38 112 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.75 //y=0.53 //x2=1.665 //y2=0.53
r147 (  37 112 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.065 //y=0.53 //x2=2.15 //y2=0.53
r148 (  37 38 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=2.065 //y=0.53 //x2=1.75 //y2=0.53
r149 (  33 112 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.615 //x2=1.665 //y2=0.53
r150 (  33 112 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.615 //x2=1.665 //y2=0.88
r151 (  32 112 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.665 //y=0.445 //x2=1.665 //y2=0.53
r152 (  31 85 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.17 //x2=1.665 //y2=0
r153 (  31 32 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=1.665 //y=0.17 //x2=1.665 //y2=0.445
r154 (  30 112 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.265 //y=0.53 //x2=1.18 //y2=0.53
r155 (  29 112 ) resistor r=6.4 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=1.58 //y=0.53 //x2=1.665 //y2=0.53
r156 (  29 30 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.58 //y=0.53 //x2=1.265 //y2=0.53
r157 (  28 112 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.445 //x2=1.18 //y2=0.53
r158 (  27 84 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0
r159 (  27 28 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=1.18 //y=0.17 //x2=1.18 //y2=0.445
r160 (  26 112 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.78 //y=0.53 //x2=0.695 //y2=0.53
r161 (  25 112 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.095 //y=0.53 //x2=1.18 //y2=0.53
r162 (  25 26 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=1.095 //y=0.53 //x2=0.78 //y2=0.53
r163 (  21 112 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.615 //x2=0.695 //y2=0.53
r164 (  21 112 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.615 //x2=0.695 //y2=1.22
r165 (  20 112 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.445 //x2=0.695 //y2=0.53
r166 (  19 81 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.17 //x2=0.695 //y2=0
r167 (  19 20 ) resistor r=18.8235 //w=0.187 //l=0.275 //layer=li \
 //thickness=0.1 //x=0.695 //y=0.17 //x2=0.695 //y2=0.445
r168 (  13 78 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.18 //y=0 //x2=5.18 //y2=0
r169 (  11 103 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=0 //x2=4.44 //y2=0
r170 (  11 13 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=0 //x2=5.18 //y2=0
r171 (  9 52 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r172 (  9 11 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.44 //y2=0
r173 (  6 87 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r174 (  3 83 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r175 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
r176 (  1 9 ) resistor r=0.0768272 //w=0.301 //l=0.185 //layer=m1 \
 //thickness=0.36 //x=2.775 //y=0 //x2=2.96 //y2=0
r177 (  1 6 ) resistor r=0.384136 //w=0.301 //l=0.925 //layer=m1 \
 //thickness=0.36 //x=2.775 //y=0 //x2=1.85 //y2=0
ends PM_OR2X1\%GND

subckt PM_OR2X1\%VDD ( 1 13 17 20 27 43 56 60 63 64 65 )
c72 ( 65 0 ) capacitor c=0.0451925f //x=4.74 //y=5.02
c73 ( 64 0 ) capacitor c=0.0423715f //x=3.87 //y=5.02
c74 ( 63 0 ) capacitor c=0.0256796f //x=1.085 //y=5.025
c75 ( 62 0 ) capacitor c=0.00591168f //x=4.885 //y=7.4
c76 ( 61 0 ) capacitor c=0.00591168f //x=4.005 //y=7.4
c77 ( 60 0 ) capacitor c=0.109776f //x=3.33 //y=7.4
c78 ( 59 0 ) capacitor c=0.00591168f //x=1.23 //y=7.4
c79 ( 56 0 ) capacitor c=0.228884f //x=5.18 //y=7.4
c80 ( 43 0 ) capacitor c=0.0287207f //x=4.8 //y=7.4
c81 ( 35 0 ) capacitor c=0.0216067f //x=3.92 //y=7.4
c82 ( 27 0 ) capacitor c=0.0778183f //x=3.16 //y=7.4
c83 ( 20 0 ) capacitor c=0.210107f //x=0.74 //y=7.4
c84 ( 17 0 ) capacitor c=0.0465804f //x=1.145 //y=7.4
c85 ( 13 0 ) capacitor c=0.22902f //x=5.18 //y=7.4
r86 (  54 62 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.97 //y=7.4 //x2=4.885 //y2=7.4
r87 (  54 56 ) resistor r=7.52941 //w=0.357 //l=0.21 //layer=li \
 //thickness=0.1 //x=4.97 //y=7.4 //x2=5.18 //y2=7.4
r88 (  47 62 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=4.885 //y=7.23 //x2=4.885 //y2=7.4
r89 (  47 65 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=4.885 //y=7.23 //x2=4.885 //y2=6.405
r90 (  44 61 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.09 //y=7.4 //x2=4.005 //y2=7.4
r91 (  44 46 ) resistor r=12.549 //w=0.357 //l=0.35 //layer=li //thickness=0.1 \
 //x=4.09 //y=7.4 //x2=4.44 //y2=7.4
r92 (  43 62 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=4.8 //y=7.4 //x2=4.885 //y2=7.4
r93 (  43 46 ) resistor r=12.9076 //w=0.357 //l=0.36 //layer=li \
 //thickness=0.1 //x=4.8 //y=7.4 //x2=4.44 //y2=7.4
r94 (  37 61 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=4.005 //y=7.23 //x2=4.005 //y2=7.4
r95 (  37 64 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=4.005 //y=7.23 //x2=4.005 //y2=6.405
r96 (  36 60 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.5 //y=7.4 //x2=3.33 //y2=7.4
r97 (  35 61 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.92 //y=7.4 //x2=4.005 //y2=7.4
r98 (  35 36 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=3.92 //y=7.4 //x2=3.5 //y2=7.4
r99 (  30 32 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r100 (  28 59 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.315 //y=7.4 //x2=1.23 //y2=7.4
r101 (  28 30 ) resistor r=19.1821 //w=0.357 //l=0.535 //layer=li \
 //thickness=0.1 //x=1.315 //y=7.4 //x2=1.85 //y2=7.4
r102 (  27 60 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.16 //y=7.4 //x2=3.33 //y2=7.4
r103 (  27 32 ) resistor r=7.17087 //w=0.357 //l=0.2 //layer=li \
 //thickness=0.1 //x=3.16 //y=7.4 //x2=2.96 //y2=7.4
r104 (  21 59 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.23 //y=7.23 //x2=1.23 //y2=7.4
r105 (  21 63 ) resistor r=33.5401 //w=0.187 //l=0.49 //layer=li \
 //thickness=0.1 //x=1.23 //y=7.23 //x2=1.23 //y2=6.74
r106 (  17 59 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.145 //y=7.4 //x2=1.23 //y2=7.4
r107 (  17 20 ) resistor r=14.521 //w=0.357 //l=0.405 //layer=li \
 //thickness=0.1 //x=1.145 //y=7.4 //x2=0.74 //y2=7.4
r108 (  13 56 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.18 //y=7.4 //x2=5.18 //y2=7.4
r109 (  11 46 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.44 //y=7.4 //x2=4.44 //y2=7.4
r110 (  11 13 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=4.44 //y=7.4 //x2=5.18 //y2=7.4
r111 (  9 32 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r112 (  9 11 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.44 //y2=7.4
r113 (  6 30 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r114 (  3 20 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r115 (  3 6 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
r116 (  1 9 ) resistor r=0.0768272 //w=0.301 //l=0.185 //layer=m1 \
 //thickness=0.36 //x=2.775 //y=7.4 //x2=2.96 //y2=7.4
r117 (  1 6 ) resistor r=0.384136 //w=0.301 //l=0.925 //layer=m1 \
 //thickness=0.36 //x=2.775 //y=7.4 //x2=1.85 //y2=7.4
ends PM_OR2X1\%VDD

subckt PM_OR2X1\%noxref_3 ( 1 2 11 12 23 24 25 30 32 40 41 42 43 44 45 46 50 \
 51 52 54 60 61 63 71 72 75 )
c136 ( 75 0 ) capacitor c=0.0159573f //x=1.965 //y=5.025
c137 ( 72 0 ) capacitor c=0.00905936f //x=1.96 //y=0.905
c138 ( 71 0 ) capacitor c=0.007684f //x=0.99 //y=0.905
c139 ( 63 0 ) capacitor c=0.0528806f //x=4.07 //y=2.085
c140 ( 61 0 ) capacitor c=0.0435629f //x=4.71 //y=1.255
c141 ( 60 0 ) capacitor c=0.0200386f //x=4.71 //y=0.91
c142 ( 54 0 ) capacitor c=0.0152946f //x=4.555 //y=1.41
c143 ( 52 0 ) capacitor c=0.0157804f //x=4.555 //y=0.755
c144 ( 51 0 ) capacitor c=0.0524991f //x=4.3 //y=4.79
c145 ( 50 0 ) capacitor c=0.0322983f //x=4.59 //y=4.79
c146 ( 46 0 ) capacitor c=0.0290017f //x=4.18 //y=1.92
c147 ( 45 0 ) capacitor c=0.0250027f //x=4.18 //y=1.565
c148 ( 44 0 ) capacitor c=0.0234316f //x=4.18 //y=1.255
c149 ( 43 0 ) capacitor c=0.0200596f //x=4.18 //y=0.91
c150 ( 42 0 ) capacitor c=0.154218f //x=4.665 //y=6.02
c151 ( 41 0 ) capacitor c=0.154243f //x=4.225 //y=6.02
c152 ( 39 0 ) capacitor c=0.00710337f //x=2.15 //y=1.655
c153 ( 32 0 ) capacitor c=0.0944546f //x=4.07 //y=2.085
c154 ( 30 0 ) capacitor c=0.112871f //x=2.59 //y=3.33
c155 ( 25 0 ) capacitor c=0.0162468f //x=2.505 //y=1.655
c156 ( 24 0 ) capacitor c=0.00499395f //x=2.195 //y=5.21
c157 ( 23 0 ) capacitor c=0.0155365f //x=2.505 //y=5.21
c158 ( 12 0 ) capacitor c=0.00277607f //x=1.265 //y=1.655
c159 ( 11 0 ) capacitor c=0.0280953f //x=2.065 //y=1.655
c160 ( 2 0 ) capacitor c=0.0155913f //x=2.705 //y=3.33
c161 ( 1 0 ) capacitor c=0.0801529f //x=3.955 //y=3.33
r162 (  63 64 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.07 //y=2.085 //x2=4.18 //y2=2.085
r163 (  61 70 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.71 //y=1.255 //x2=4.67 //y2=1.41
r164 (  60 69 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.71 //y=0.91 //x2=4.67 //y2=0.755
r165 (  60 61 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.71 //y=0.91 //x2=4.71 //y2=1.255
r166 (  55 68 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.335 //y=1.41 //x2=4.22 //y2=1.41
r167 (  54 70 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.555 //y=1.41 //x2=4.67 //y2=1.41
r168 (  53 67 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.335 //y=0.755 //x2=4.22 //y2=0.755
r169 (  52 69 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=4.555 //y=0.755 //x2=4.67 //y2=0.755
r170 (  52 53 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=4.555 //y=0.755 //x2=4.335 //y2=0.755
r171 (  50 57 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.59 //y=4.79 //x2=4.665 //y2=4.865
r172 (  50 51 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=4.59 //y=4.79 //x2=4.3 //y2=4.79
r173 (  47 51 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=4.225 //y=4.865 //x2=4.3 //y2=4.79
r174 (  47 66 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=4.225 //y=4.865 //x2=4.07 //y2=4.7
r175 (  46 64 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.92 //x2=4.18 //y2=2.085
r176 (  45 68 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.565 //x2=4.22 //y2=1.41
r177 (  45 46 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.565 //x2=4.18 //y2=1.92
r178 (  44 68 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.18 //y=1.255 //x2=4.22 //y2=1.41
r179 (  43 67 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=4.18 //y=0.91 //x2=4.22 //y2=0.755
r180 (  43 44 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=4.18 //y=0.91 //x2=4.18 //y2=1.255
r181 (  42 57 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.665 //y=6.02 //x2=4.665 //y2=4.865
r182 (  41 47 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=4.225 //y=6.02 //x2=4.225 //y2=4.865
r183 (  40 54 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.445 //y=1.41 //x2=4.555 //y2=1.41
r184 (  40 55 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=4.445 //y=1.41 //x2=4.335 //y2=1.41
r185 (  37 66 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.07 //y=4.7 //x2=4.07 //y2=4.7
r186 (  35 37 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=4.07 //y=3.33 //x2=4.07 //y2=4.7
r187 (  32 63 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=4.07 //y=2.085 //x2=4.07 //y2=2.085
r188 (  32 35 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=4.07 //y=2.085 //x2=4.07 //y2=3.33
r189 (  28 30 ) resistor r=122.866 //w=0.187 //l=1.795 //layer=li \
 //thickness=0.1 //x=2.59 //y=5.125 //x2=2.59 //y2=3.33
r190 (  27 30 ) resistor r=108.834 //w=0.187 //l=1.59 //layer=li \
 //thickness=0.1 //x=2.59 //y=1.74 //x2=2.59 //y2=3.33
r191 (  26 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.235 //y=1.655 //x2=2.15 //y2=1.655
r192 (  25 27 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.59 //y2=1.74
r193 (  25 26 ) resistor r=18.4813 //w=0.187 //l=0.27 //layer=li \
 //thickness=0.1 //x=2.505 //y=1.655 //x2=2.235 //y2=1.655
r194 (  23 28 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.21 //x2=2.59 //y2=5.125
r195 (  23 24 ) resistor r=21.2193 //w=0.187 //l=0.31 //layer=li \
 //thickness=0.1 //x=2.505 //y=5.21 //x2=2.195 //y2=5.21
r196 (  19 39 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1.655
r197 (  19 72 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=2.15 //y=1.57 //x2=2.15 //y2=1
r198 (  13 24 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.295 //x2=2.195 //y2=5.21
r199 (  13 75 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=2.11 //y=5.295 //x2=2.11 //y2=5.72
r200 (  11 39 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.065 //y=1.655 //x2=2.15 //y2=1.655
r201 (  11 12 ) resistor r=54.7594 //w=0.187 //l=0.8 //layer=li \
 //thickness=0.1 //x=2.065 //y=1.655 //x2=1.265 //y2=1.655
r202 (  7 12 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.18 //y=1.57 //x2=1.265 //y2=1.655
r203 (  7 71 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=1.18 //y=1.57 //x2=1.18 //y2=1
r204 (  6 35 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=3.33 //x2=4.07 //y2=3.33
r205 (  4 30 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=2.59 //y=3.33 //x2=2.59 //y2=3.33
r206 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=2.705 //y=3.33 //x2=2.59 //y2=3.33
r207 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=3.955 //y=3.33 //x2=4.07 //y2=3.33
r208 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=3.955 //y=3.33 //x2=2.705 //y2=3.33
ends PM_OR2X1\%noxref_3

subckt PM_OR2X1\%A ( 1 2 3 4 5 6 7 10 20 22 23 24 25 26 27 28 32 34 37 39 40 \
 45 )
c66 ( 45 0 ) capacitor c=0.04214f //x=0.955 //y=4.705
c67 ( 40 0 ) capacitor c=0.0321911f //x=1.445 //y=1.25
c68 ( 39 0 ) capacitor c=0.0185201f //x=1.445 //y=0.905
c69 ( 37 0 ) capacitor c=0.0344254f //x=1.375 //y=4.795
c70 ( 34 0 ) capacitor c=0.0133656f //x=1.29 //y=1.405
c71 ( 32 0 ) capacitor c=0.0157804f //x=1.29 //y=0.75
c72 ( 28 0 ) capacitor c=0.0828832f //x=0.915 //y=1.915
c73 ( 27 0 ) capacitor c=0.022867f //x=0.915 //y=1.56
c74 ( 26 0 ) capacitor c=0.0234318f //x=0.915 //y=1.25
c75 ( 25 0 ) capacitor c=0.0192004f //x=0.915 //y=0.905
c76 ( 24 0 ) capacitor c=0.110795f //x=1.45 //y=6.025
c77 ( 23 0 ) capacitor c=0.153847f //x=1.01 //y=6.025
c78 ( 20 0 ) capacitor c=0.00993392f //x=0.955 //y=4.705
c79 ( 10 0 ) capacitor c=0.112424f //x=1.11 //y=2.08
r80 (  47 48 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=0.955 //y=4.795 //x2=0.955 //y2=4.87
r81 (  45 47 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=0.955 //y=4.705 //x2=0.955 //y2=4.795
r82 (  40 54 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=1.25 //x2=1.405 //y2=1.405
r83 (  39 53 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.905 //x2=1.405 //y2=0.75
r84 (  39 40 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.445 //y=0.905 //x2=1.445 //y2=1.25
r85 (  38 47 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=1.09 //y=4.795 //x2=0.955 //y2=4.795
r86 (  37 41 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.375 //y=4.795 //x2=1.45 //y2=4.87
r87 (  37 38 ) resistor r=146.138 //w=0.094 //l=0.285 //layer=ply \
 //thickness=0.18 //x=1.375 //y=4.795 //x2=1.09 //y2=4.795
r88 (  35 52 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=1.405 //x2=0.955 //y2=1.405
r89 (  34 54 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=1.405 //x2=1.405 //y2=1.405
r90 (  33 51 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.07 //y=0.75 //x2=0.955 //y2=0.75
r91 (  32 53 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.75 //x2=1.405 //y2=0.75
r92 (  32 33 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.29 //y=0.75 //x2=1.07 //y2=0.75
r93 (  28 50 ) resistor r=34.8111 //w=0.27 //l=0.264953 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.915 //x2=1.11 //y2=2.08
r94 (  27 52 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.56 //x2=0.955 //y2=1.405
r95 (  27 28 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.56 //x2=0.915 //y2=1.915
r96 (  26 52 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=1.25 //x2=0.955 //y2=1.405
r97 (  25 51 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.905 //x2=0.955 //y2=0.75
r98 (  25 26 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.915 //y=0.905 //x2=0.915 //y2=1.25
r99 (  24 41 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.45 //y=6.025 //x2=1.45 //y2=4.87
r100 (  23 48 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.01 //y=6.025 //x2=1.01 //y2=4.87
r101 (  22 34 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.405 //x2=1.29 //y2=1.405
r102 (  22 35 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.18 //y=1.405 //x2=1.07 //y2=1.405
r103 (  20 45 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=0.955 //y=4.705 //x2=0.955 //y2=4.705
r104 (  20 21 ) resistor r=7.81102 //w=0.254 //l=0.155 //layer=li \
 //thickness=0.1 //x=0.955 //y=4.705 //x2=1.11 //y2=4.705
r105 (  10 50 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r106 (  8 21 ) resistor r=3.23951 //w=0.254 //l=0.165 //layer=li \
 //thickness=0.1 //x=1.11 //y=4.54 //x2=1.11 //y2=4.705
r107 (  7 8 ) resistor r=6.84492 //w=0.187 //l=0.1 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.44 //x2=1.11 //y2=4.54
r108 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=4.07 //x2=1.11 //y2=4.44
r109 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=3.7 //x2=1.11 //y2=4.07
r110 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=3.33 //x2=1.11 //y2=3.7
r111 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.96 //x2=1.11 //y2=3.33
r112 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.59 //x2=1.11 //y2=2.96
r113 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.22 //x2=1.11 //y2=2.59
r114 (  1 10 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=1.11 //y=2.22 //x2=1.11 //y2=2.08
ends PM_OR2X1\%A

subckt PM_OR2X1\%B ( 1 2 3 4 5 6 7 8 10 21 22 23 24 25 26 31 33 35 41 42 44 45 \
 48 )
c69 ( 48 0 ) capacitor c=0.0369822f //x=1.885 //y=4.705
c70 ( 45 0 ) capacitor c=0.0279572f //x=1.85 //y=1.915
c71 ( 44 0 ) capacitor c=0.0422144f //x=1.85 //y=2.08
c72 ( 42 0 ) capacitor c=0.0237734f //x=2.415 //y=1.255
c73 ( 41 0 ) capacitor c=0.0191782f //x=2.415 //y=0.905
c74 ( 35 0 ) capacitor c=0.0346941f //x=2.26 //y=1.405
c75 ( 33 0 ) capacitor c=0.0157803f //x=2.26 //y=0.75
c76 ( 31 0 ) capacitor c=0.0360787f //x=2.255 //y=4.795
c77 ( 26 0 ) capacitor c=0.0199921f //x=1.885 //y=1.56
c78 ( 25 0 ) capacitor c=0.0169608f //x=1.885 //y=1.255
c79 ( 24 0 ) capacitor c=0.0185462f //x=1.885 //y=0.905
c80 ( 23 0 ) capacitor c=0.15325f //x=2.33 //y=6.025
c81 ( 22 0 ) capacitor c=0.110232f //x=1.89 //y=6.025
c82 ( 10 0 ) capacitor c=0.0809838f //x=1.85 //y=2.08
c83 ( 8 0 ) capacitor c=0.00521267f //x=1.85 //y=4.54
r84 (  50 51 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=1.885 //y=4.795 //x2=1.885 //y2=4.87
r85 (  48 50 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=1.885 //y=4.705 //x2=1.885 //y2=4.795
r86 (  44 45 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=1.85 //y=2.08 //x2=1.85 //y2=1.915
r87 (  42 55 ) resistor r=4.95774 //w=0.164 //l=0.112 //layer=ply \
 //thickness=0.18 //x=2.415 //y=1.255 //x2=2.415 //y2=1.367
r88 (  41 54 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.375 //y2=0.75
r89 (  41 42 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=2.415 //y=0.905 //x2=2.415 //y2=1.255
r90 (  36 53 ) resistor r=10.8103 //w=0.211 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=1.405 //x2=1.925 //y2=1.405
r91 (  35 55 ) resistor r=45.9962 //w=0.164 //l=0.17296 //layer=ply \
 //thickness=0.18 //x=2.26 //y=1.405 //x2=2.415 //y2=1.367
r92 (  34 52 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.04 //y=0.75 //x2=1.925 //y2=0.75
r93 (  33 54 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.375 //y2=0.75
r94 (  33 34 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=2.26 //y=0.75 //x2=2.04 //y2=0.75
r95 (  32 50 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.02 //y=4.795 //x2=1.885 //y2=4.795
r96 (  31 38 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.795 //x2=2.33 //y2=4.87
r97 (  31 32 ) resistor r=120.5 //w=0.094 //l=0.235 //layer=ply \
 //thickness=0.18 //x=2.255 //y=4.795 //x2=2.02 //y2=4.795
r98 (  26 53 ) resistor r=39.5036 //w=0.211 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.925 //y2=1.405
r99 (  26 45 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.56 //x2=1.885 //y2=1.915
r100 (  25 53 ) resistor r=38.3614 //w=0.211 //l=0.168819 //layer=ply \
 //thickness=0.18 //x=1.885 //y=1.255 //x2=1.925 //y2=1.405
r101 (  24 52 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.925 //y2=0.75
r102 (  24 25 ) resistor r=179.468 //w=0.094 //l=0.35 //layer=ply \
 //thickness=0.18 //x=1.885 //y=0.905 //x2=1.885 //y2=1.255
r103 (  23 38 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.33 //y=6.025 //x2=2.33 //y2=4.87
r104 (  22 51 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.89 //y=6.025 //x2=1.89 //y2=4.87
r105 (  21 35 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.26 //y2=1.405
r106 (  21 36 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=2.15 //y=1.405 //x2=2.04 //y2=1.405
r107 (  20 48 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.885 //y=4.705 //x2=1.885 //y2=4.705
r108 (  10 44 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.85 //y=2.08 //x2=1.85 //y2=2.08
r109 (  8 20 ) resistor r=11.332 //w=0.189 //l=0.173292 //layer=li \
 //thickness=0.1 //x=1.85 //y=4.54 //x2=1.867 //y2=4.705
r110 (  7 8 ) resistor r=6.84492 //w=0.187 //l=0.1 //layer=li //thickness=0.1 \
 //x=1.85 //y=4.44 //x2=1.85 //y2=4.54
r111 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=4.07 //x2=1.85 //y2=4.44
r112 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=3.7 //x2=1.85 //y2=4.07
r113 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=3.33 //x2=1.85 //y2=3.7
r114 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=2.96 //x2=1.85 //y2=3.33
r115 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=2.59 //x2=1.85 //y2=2.96
r116 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=1.85 //y=2.22 //x2=1.85 //y2=2.59
r117 (  1 10 ) resistor r=9.58289 //w=0.187 //l=0.14 //layer=li \
 //thickness=0.1 //x=1.85 //y=2.22 //x2=1.85 //y2=2.08
ends PM_OR2X1\%B

subckt PM_OR2X1\%noxref_6 ( 7 8 15 16 23 24 25 )
c41 ( 25 0 ) capacitor c=0.030764f //x=2.405 //y=5.025
c42 ( 24 0 ) capacitor c=0.0185379f //x=1.525 //y=5.025
c43 ( 23 0 ) capacitor c=0.0409962f //x=0.655 //y=5.025
c44 ( 16 0 ) capacitor c=0.00193672f //x=1.755 //y=6.91
c45 ( 15 0 ) capacitor c=0.01354f //x=2.465 //y=6.91
c46 ( 8 0 ) capacitor c=0.00844339f //x=0.875 //y=5.21
c47 ( 7 0 ) capacitor c=0.0240359f //x=1.585 //y=5.21
r48 (  17 25 ) resistor r=5.81818 //w=0.187 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.55 //y=6.825 //x2=2.55 //y2=6.74
r49 (  15 17 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=2.465 //y=6.91 //x2=2.55 //y2=6.825
r50 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.465 //y=6.91 //x2=1.755 //y2=6.91
r51 (  10 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.67 //y=6.825 //x2=1.755 //y2=6.91
r52 (  10 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.67 //y=6.825 //x2=1.67 //y2=6.4
r53 (  9 24 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=1.67 //y=5.295 //x2=1.67 //y2=5.72
r54 (  7 9 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.585 //y=5.21 //x2=1.67 //y2=5.295
r55 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=1.585 //y=5.21 //x2=0.875 //y2=5.21
r56 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=0.79 //y=5.295 //x2=0.875 //y2=5.21
r57 (  1 23 ) resistor r=29.0909 //w=0.187 //l=0.425 //layer=li \
 //thickness=0.1 //x=0.79 //y=5.295 //x2=0.79 //y2=5.72
ends PM_OR2X1\%noxref_6

subckt PM_OR2X1\%Y ( 1 2 3 4 5 6 7 18 19 20 21 31 33 )
c44 ( 33 0 ) capacitor c=0.028734f //x=4.3 //y=5.02
c45 ( 31 0 ) capacitor c=0.0173218f //x=4.255 //y=0.91
c46 ( 21 0 ) capacitor c=0.00575887f //x=4.53 //y=4.58
c47 ( 20 0 ) capacitor c=0.0136889f //x=4.725 //y=4.58
c48 ( 19 0 ) capacitor c=0.00636159f //x=4.525 //y=2.08
c49 ( 18 0 ) capacitor c=0.0140707f //x=4.725 //y=2.08
c50 ( 1 0 ) capacitor c=0.105613f //x=4.81 //y=2.22
r51 (  20 23 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=4.58 //x2=4.81 //y2=4.495
r52 (  20 21 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=4.725 //y=4.58 //x2=4.53 //y2=4.58
r53 (  18 22 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.725 //y=2.08 //x2=4.81 //y2=2.165
r54 (  18 19 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=4.725 //y=2.08 //x2=4.525 //y2=2.08
r55 (  12 21 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.445 //y=4.665 //x2=4.53 //y2=4.58
r56 (  12 33 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li \
 //thickness=0.1 //x=4.445 //y=4.665 //x2=4.445 //y2=5.725
r57 (  8 19 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=4.44 //y=1.995 //x2=4.525 //y2=2.08
r58 (  8 31 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=4.44 //y=1.995 //x2=4.44 //y2=1.005
r59 (  7 23 ) resistor r=3.76471 //w=0.187 //l=0.055 //layer=li \
 //thickness=0.1 //x=4.81 //y=4.44 //x2=4.81 //y2=4.495
r60 (  6 7 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.81 //y=4.07 //x2=4.81 //y2=4.44
r61 (  5 6 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.81 //y=3.7 //x2=4.81 //y2=4.07
r62 (  4 5 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.81 //y=3.33 //x2=4.81 //y2=3.7
r63 (  3 4 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.81 //y=2.96 //x2=4.81 //y2=3.33
r64 (  2 3 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.81 //y=2.59 //x2=4.81 //y2=2.96
r65 (  1 2 ) resistor r=25.3262 //w=0.187 //l=0.37 //layer=li //thickness=0.1 \
 //x=4.81 //y=2.22 //x2=4.81 //y2=2.59
r66 (  1 22 ) resistor r=3.76471 //w=0.187 //l=0.055 //layer=li \
 //thickness=0.1 //x=4.81 //y=2.22 //x2=4.81 //y2=2.165
ends PM_OR2X1\%Y

