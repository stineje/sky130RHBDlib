VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO VOTERN3X1
  CLASS CORE ;
  FOREIGN VOTERN3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.990 BY 7.400 ;
  SYMMETRY X Y R90 ;
  SITE unitrh ;
  PIN YN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.734950 ;
    PORT
      LAYER li1 ;
        RECT 7.805 5.295 7.975 6.565 ;
        RECT 8.685 5.295 8.855 6.565 ;
        RECT 7.805 5.125 9.335 5.295 ;
        RECT 9.165 1.730 9.335 5.125 ;
        RECT 8.725 1.560 9.335 1.730 ;
        RECT 2.065 1.170 2.235 1.345 ;
        RECT 2.060 1.015 2.235 1.170 ;
        RECT 2.060 0.835 2.230 1.015 ;
        RECT 5.395 0.835 5.565 1.345 ;
        RECT 8.725 0.835 8.895 1.560 ;
      LAYER mcon ;
        RECT 2.065 1.095 2.235 1.265 ;
        RECT 5.395 1.095 5.565 1.265 ;
        RECT 8.725 1.095 8.895 1.265 ;
      LAYER met1 ;
        RECT 2.035 1.265 2.265 1.295 ;
        RECT 5.365 1.265 5.595 1.295 ;
        RECT 8.695 1.265 8.925 1.295 ;
        RECT 2.005 1.095 8.955 1.265 ;
        RECT 2.035 1.065 2.265 1.095 ;
        RECT 5.365 1.065 5.595 1.095 ;
        RECT 8.695 1.065 8.925 1.095 ;
    END
  END YN
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.053700 ;
    PORT
      LAYER li1 ;
        RECT 1.805 4.710 1.975 4.870 ;
        RECT 1.765 4.540 1.975 4.710 ;
        RECT 8.425 4.540 8.615 4.870 ;
        RECT 1.765 1.915 1.935 4.540 ;
        RECT 8.425 1.915 8.595 4.540 ;
      LAYER mcon ;
        RECT 1.765 3.985 1.935 4.155 ;
        RECT 8.425 3.985 8.595 4.155 ;
      LAYER met1 ;
        RECT 1.735 4.155 1.965 4.185 ;
        RECT 8.395 4.155 8.625 4.185 ;
        RECT 1.705 3.985 8.655 4.155 ;
        RECT 1.735 3.955 1.965 3.985 ;
        RECT 8.395 3.955 8.625 3.985 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.066500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.915 0.825 4.870 ;
        RECT 4.355 1.915 4.525 4.870 ;
      LAYER mcon ;
        RECT 0.655 4.355 0.825 4.525 ;
        RECT 4.355 4.355 4.525 4.525 ;
      LAYER met1 ;
        RECT 0.625 4.525 0.855 4.555 ;
        RECT 4.325 4.525 4.555 4.555 ;
        RECT 0.595 4.355 4.585 4.525 ;
        RECT 0.625 4.325 0.855 4.355 ;
        RECT 4.325 4.325 4.555 4.355 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.060500 ;
    PORT
      LAYER li1 ;
        RECT 5.835 1.915 6.005 4.870 ;
        RECT 7.315 1.915 7.485 4.870 ;
      LAYER mcon ;
        RECT 5.835 1.995 6.005 2.165 ;
        RECT 7.315 1.995 7.485 2.165 ;
      LAYER met1 ;
        RECT 5.805 2.165 6.035 2.195 ;
        RECT 7.285 2.165 7.515 2.195 ;
        RECT 5.775 1.995 7.545 2.165 ;
        RECT 5.805 1.965 6.035 1.995 ;
        RECT 7.285 1.965 7.515 1.995 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.435 3.930 10.425 7.750 ;
      LAYER li1 ;
        RECT -0.170 7.230 10.160 7.570 ;
        RECT -0.170 4.110 0.170 7.230 ;
        RECT 0.705 5.125 0.875 7.230 ;
        RECT 1.585 5.555 1.755 7.230 ;
        RECT 2.465 5.125 2.635 7.230 ;
        RECT 3.160 4.110 3.500 7.230 ;
        RECT 6.490 4.110 6.830 7.230 ;
        RECT 9.820 4.110 10.160 7.230 ;
      LAYER mcon ;
        RECT 0.285 7.315 0.455 7.485 ;
        RECT 0.655 7.315 0.825 7.485 ;
        RECT 1.025 7.315 1.195 7.485 ;
        RECT 1.395 7.315 1.565 7.485 ;
        RECT 1.765 7.315 1.935 7.485 ;
        RECT 2.135 7.315 2.305 7.485 ;
        RECT 2.505 7.315 2.675 7.485 ;
        RECT 2.875 7.315 3.045 7.485 ;
        RECT 3.615 7.315 3.785 7.485 ;
        RECT 3.985 7.315 4.155 7.485 ;
        RECT 4.355 7.315 4.525 7.485 ;
        RECT 4.725 7.315 4.895 7.485 ;
        RECT 5.095 7.315 5.265 7.485 ;
        RECT 5.465 7.315 5.635 7.485 ;
        RECT 5.835 7.315 6.005 7.485 ;
        RECT 6.205 7.315 6.375 7.485 ;
        RECT 6.945 7.315 7.115 7.485 ;
        RECT 7.315 7.315 7.485 7.485 ;
        RECT 7.685 7.315 7.855 7.485 ;
        RECT 8.055 7.315 8.225 7.485 ;
        RECT 8.425 7.315 8.595 7.485 ;
        RECT 8.795 7.315 8.965 7.485 ;
        RECT 9.165 7.315 9.335 7.485 ;
        RECT 9.535 7.315 9.705 7.485 ;
      LAYER met1 ;
        RECT -0.170 7.230 10.160 7.570 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT -0.170 -0.170 10.160 2.720 ;
      LAYER li1 ;
        RECT -0.170 0.170 0.170 2.720 ;
        RECT 1.095 0.170 1.265 1.120 ;
        RECT 3.160 0.170 3.500 2.720 ;
        RECT 4.425 0.170 4.595 1.120 ;
        RECT 6.490 0.170 6.830 2.720 ;
        RECT 7.755 0.170 7.925 1.120 ;
        RECT 9.820 0.170 10.160 2.720 ;
        RECT -0.170 -0.170 10.160 0.170 ;
      LAYER mcon ;
        RECT 0.285 -0.085 0.455 0.085 ;
        RECT 0.655 -0.085 0.825 0.085 ;
        RECT 1.025 -0.085 1.195 0.085 ;
        RECT 1.395 -0.085 1.565 0.085 ;
        RECT 1.765 -0.085 1.935 0.085 ;
        RECT 2.135 -0.085 2.305 0.085 ;
        RECT 2.505 -0.085 2.675 0.085 ;
        RECT 2.875 -0.085 3.045 0.085 ;
        RECT 3.615 -0.085 3.785 0.085 ;
        RECT 3.985 -0.085 4.155 0.085 ;
        RECT 4.355 -0.085 4.525 0.085 ;
        RECT 4.725 -0.085 4.895 0.085 ;
        RECT 5.095 -0.085 5.265 0.085 ;
        RECT 5.465 -0.085 5.635 0.085 ;
        RECT 5.835 -0.085 6.005 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.945 -0.085 7.115 0.085 ;
        RECT 7.315 -0.085 7.485 0.085 ;
        RECT 7.685 -0.085 7.855 0.085 ;
        RECT 8.055 -0.085 8.225 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.795 -0.085 8.965 0.085 ;
        RECT 9.165 -0.085 9.335 0.085 ;
        RECT 9.535 -0.085 9.705 0.085 ;
      LAYER met1 ;
        RECT -0.170 -0.170 10.160 0.170 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 1.145 6.825 1.325 6.995 ;
        RECT 1.145 5.295 1.315 6.825 ;
        RECT 2.025 5.295 2.195 6.995 ;
        RECT 1.145 5.125 2.195 5.295 ;
        RECT 2.025 5.045 2.195 5.125 ;
        RECT 4.025 6.825 5.955 6.995 ;
        RECT 4.025 5.045 4.195 6.825 ;
        RECT 4.465 5.295 4.635 6.565 ;
        RECT 4.905 5.555 5.075 6.825 ;
        RECT 5.345 5.295 5.515 6.565 ;
        RECT 5.785 5.375 5.955 6.825 ;
        RECT 7.365 6.825 9.295 6.995 ;
        RECT 4.465 5.125 5.515 5.295 ;
        RECT 5.345 5.045 5.515 5.125 ;
        RECT 7.365 5.045 7.535 6.825 ;
        RECT 8.245 5.555 8.415 6.825 ;
        RECT 9.125 5.555 9.295 6.825 ;
        RECT 0.610 1.665 0.780 1.745 ;
        RECT 1.580 1.665 1.750 1.745 ;
        RECT 0.610 1.495 1.750 1.665 ;
        RECT 0.610 0.365 0.780 1.495 ;
        RECT 1.580 0.615 1.750 1.495 ;
        RECT 2.550 0.615 2.720 1.745 ;
        RECT 1.580 0.445 2.720 0.615 ;
        RECT 1.580 0.365 1.750 0.445 ;
        RECT 2.550 0.365 2.720 0.445 ;
        RECT 3.940 1.665 4.110 1.745 ;
        RECT 4.910 1.665 5.080 1.745 ;
        RECT 3.940 1.495 5.080 1.665 ;
        RECT 3.940 0.365 4.110 1.495 ;
        RECT 4.910 0.615 5.080 1.495 ;
        RECT 5.880 0.615 6.050 1.745 ;
        RECT 4.910 0.445 6.050 0.615 ;
        RECT 4.910 0.365 5.080 0.445 ;
        RECT 5.880 0.365 6.050 0.445 ;
        RECT 7.270 1.665 7.440 1.745 ;
        RECT 8.240 1.665 8.410 1.745 ;
        RECT 7.270 1.495 8.410 1.665 ;
        RECT 7.270 0.365 7.440 1.495 ;
        RECT 8.240 0.615 8.410 1.495 ;
        RECT 9.210 0.615 9.380 1.390 ;
        RECT 8.240 0.445 9.380 0.615 ;
        RECT 8.240 0.365 8.410 0.445 ;
        RECT 9.210 0.365 9.380 0.445 ;
      LAYER mcon ;
        RECT 2.025 5.125 2.195 5.295 ;
        RECT 4.025 5.125 4.195 5.295 ;
        RECT 5.345 5.125 5.515 5.295 ;
        RECT 7.365 5.125 7.535 5.295 ;
      LAYER met1 ;
        RECT 1.995 5.295 2.225 5.325 ;
        RECT 3.995 5.295 4.225 5.325 ;
        RECT 5.315 5.295 5.545 5.325 ;
        RECT 7.335 5.295 7.565 5.325 ;
        RECT 1.965 5.125 4.255 5.295 ;
        RECT 5.285 5.125 7.595 5.295 ;
        RECT 1.995 5.095 2.225 5.125 ;
        RECT 3.995 5.095 4.225 5.125 ;
        RECT 5.315 5.095 5.545 5.125 ;
        RECT 7.335 5.095 7.565 5.125 ;
  END
END VOTERN3X1
END LIBRARY

