// File: and3x1_pcell.spi.pex
// Created: Tue Oct 15 15:54:33 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_AND3X1_PCELL\%noxref_1 ( 13 17 20 25 35 38 43 47 60 67 74 75 )
c88 ( 75 0 ) capacitor c=0.0598672f //x=5.305 //y=0.37
c89 ( 74 0 ) capacitor c=0.0226959f //x=0.885 //y=0.875
c90 ( 67 0 ) capacitor c=0.23428f //x=6.41 //y=0
c91 ( 60 0 ) capacitor c=0.104423f //x=4.81 //y=0
c92 ( 59 0 ) capacitor c=0.00440144f //x=1.075 //y=0
c93 ( 50 0 ) capacitor c=0.00587411f //x=6.41 //y=0.45
c94 ( 47 0 ) capacitor c=0.00542558f //x=6.325 //y=0.535
c95 ( 46 0 ) capacitor c=0.00479856f //x=5.925 //y=0.45
c96 ( 43 0 ) capacitor c=0.0068422f //x=5.84 //y=0.535
c97 ( 38 0 ) capacitor c=0.00592191f //x=5.44 //y=0.45
c98 ( 35 0 ) capacitor c=0.0164879f //x=5.355 //y=0
c99 ( 25 0 ) capacitor c=0.131647f //x=4.64 //y=0
c100 ( 20 0 ) capacitor c=0.178285f //x=0.74 //y=0
c101 ( 17 0 ) capacitor c=0.0367385f //x=0.99 //y=0
c102 ( 13 0 ) capacitor c=0.259992f //x=6.29 //y=0
r103 (  66 67 ) resistor r=4.30252 //w=0.357 //l=0.12 //layer=li \
 //thickness=0.1 //x=6.29 //y=0 //x2=6.41 //y2=0
r104 (  64 66 ) resistor r=13.0868 //w=0.357 //l=0.365 //layer=li \
 //thickness=0.1 //x=5.925 //y=0 //x2=6.29 //y2=0
r105 (  63 64 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=5.55 //y=0 //x2=5.925 //y2=0
r106 (  61 63 ) resistor r=3.94398 //w=0.357 //l=0.11 //layer=li \
 //thickness=0.1 //x=5.44 //y=0 //x2=5.55 //y2=0
r107 (  51 75 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.41 //y=0.62 //x2=6.41 //y2=0.535
r108 (  51 75 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=6.41 //y=0.62 //x2=6.41 //y2=1.225
r109 (  50 75 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.41 //y=0.45 //x2=6.41 //y2=0.535
r110 (  49 67 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.41 //y=0.17 //x2=6.41 //y2=0
r111 (  49 50 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=6.41 //y=0.17 //x2=6.41 //y2=0.45
r112 (  48 75 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.01 //y=0.535 //x2=5.925 //y2=0.535
r113 (  47 75 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.325 //y=0.535 //x2=6.41 //y2=0.535
r114 (  47 48 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=6.325 //y=0.535 //x2=6.01 //y2=0.535
r115 (  46 75 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.925 //y=0.45 //x2=5.925 //y2=0.535
r116 (  45 64 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.925 //y=0.17 //x2=5.925 //y2=0
r117 (  45 46 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=5.925 //y=0.17 //x2=5.925 //y2=0.45
r118 (  44 75 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.525 //y=0.535 //x2=5.44 //y2=0.535
r119 (  43 75 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.84 //y=0.535 //x2=5.925 //y2=0.535
r120 (  43 44 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=5.84 //y=0.535 //x2=5.525 //y2=0.535
r121 (  39 75 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.44 //y=0.62 //x2=5.44 //y2=0.535
r122 (  39 75 ) resistor r=41.4118 //w=0.187 //l=0.605 //layer=li \
 //thickness=0.1 //x=5.44 //y=0.62 //x2=5.44 //y2=1.225
r123 (  38 75 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.44 //y=0.45 //x2=5.44 //y2=0.535
r124 (  37 61 ) resistor r=5.03728 //w=0.34 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.44 //y=0.17 //x2=5.44 //y2=0
r125 (  37 38 ) resistor r=19.1658 //w=0.187 //l=0.28 //layer=li \
 //thickness=0.1 //x=5.44 //y=0.17 //x2=5.44 //y2=0.45
r126 (  36 60 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=4.98 //y=0 //x2=4.81 //y2=0
r127 (  35 61 ) resistor r=3.04762 //w=0.357 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.355 //y=0 //x2=5.44 //y2=0
r128 (  35 36 ) resistor r=13.4454 //w=0.357 //l=0.375 //layer=li \
 //thickness=0.1 //x=5.355 //y=0 //x2=4.98 //y2=0
r129 (  30 32 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=2.96 //y=0 //x2=4.07 //y2=0
r130 (  28 30 ) resistor r=39.7983 //w=0.357 //l=1.11 //layer=li \
 //thickness=0.1 //x=1.85 //y=0 //x2=2.96 //y2=0
r131 (  26 59 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.075 //y2=0
r132 (  26 28 ) resistor r=24.7395 //w=0.357 //l=0.69 //layer=li \
 //thickness=0.1 //x=1.16 //y=0 //x2=1.85 //y2=0
r133 (  25 60 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=4.64 //y=0 //x2=4.81 //y2=0
r134 (  25 32 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=0 //x2=4.07 //y2=0
r135 (  21 59 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0
r136 (  21 74 ) resistor r=54.4171 //w=0.187 //l=0.795 //layer=li \
 //thickness=0.1 //x=1.075 //y=0.17 //x2=1.075 //y2=0.965
r137 (  17 59 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=1.075 //y2=0
r138 (  17 20 ) resistor r=8.96359 //w=0.357 //l=0.25 //layer=li \
 //thickness=0.1 //x=0.99 //y=0 //x2=0.74 //y2=0
r139 (  13 66 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=6.29 //y=0 //x2=6.29 //y2=0
r140 (  11 63 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=0 //x2=5.55 //y2=0
r141 (  11 13 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=0 //x2=6.29 //y2=0
r142 (  9 32 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=0 //x2=4.07 //y2=0
r143 (  9 11 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=0 //x2=5.55 //y2=0
r144 (  7 30 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=0 //x2=2.96 //y2=0
r145 (  7 9 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=0 //x2=4.07 //y2=0
r146 (  5 28 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=0 //x2=1.85 //y2=0
r147 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=0 //x2=2.96 //y2=0
r148 (  2 20 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=0 //x2=0.74 //y2=0
r149 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=0 //x2=1.85 //y2=0
ends PM_AND3X1_PCELL\%noxref_1

subckt PM_AND3X1_PCELL\%noxref_2 ( 13 20 27 37 45 55 69 85 89 90 91 92 93 94 \
 95 )
c83 ( 95 0 ) capacitor c=0.0451925f //x=6.22 //y=5.02
c84 ( 94 0 ) capacitor c=0.0422823f //x=5.35 //y=5.02
c85 ( 93 0 ) capacitor c=0.0455453f //x=3.585 //y=5.02
c86 ( 92 0 ) capacitor c=0.0244794f //x=2.705 //y=5.02
c87 ( 91 0 ) capacitor c=0.0244794f //x=1.825 //y=5.02
c88 ( 90 0 ) capacitor c=0.0533644f //x=0.955 //y=5.02
c89 ( 89 0 ) capacitor c=0.234796f //x=6.29 //y=7.4
c90 ( 87 0 ) capacitor c=0.00591168f //x=5.55 //y=7.4
c91 ( 85 0 ) capacitor c=0.130858f //x=4.81 //y=7.4
c92 ( 84 0 ) capacitor c=0.00591168f //x=3.73 //y=7.4
c93 ( 83 0 ) capacitor c=0.00591168f //x=2.85 //y=7.4
c94 ( 82 0 ) capacitor c=0.00591168f //x=1.97 //y=7.4
c95 ( 81 0 ) capacitor c=0.00591168f //x=1.09 //y=7.4
c96 ( 69 0 ) capacitor c=0.0287207f //x=6.28 //y=7.4
c97 ( 61 0 ) capacitor c=0.0216067f //x=5.4 //y=7.4
c98 ( 55 0 ) capacitor c=0.0418861f //x=4.64 //y=7.4
c99 ( 45 0 ) capacitor c=0.028513f //x=3.645 //y=7.4
c100 ( 37 0 ) capacitor c=0.0287069f //x=2.765 //y=7.4
c101 ( 27 0 ) capacitor c=0.0292055f //x=1.885 //y=7.4
c102 ( 20 0 ) capacitor c=0.235022f //x=0.74 //y=7.4
c103 ( 17 0 ) capacitor c=0.0452081f //x=1.005 //y=7.4
c104 ( 13 0 ) capacitor c=0.291287f //x=6.29 //y=7.4
r105 (  71 89 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=6.365 //y=7.23 //x2=6.365 //y2=7.4
r106 (  71 95 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=6.365 //y=7.23 //x2=6.365 //y2=6.405
r107 (  70 87 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.57 //y=7.4 //x2=5.485 //y2=7.4
r108 (  69 89 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=6.28 //y=7.4 //x2=6.365 //y2=7.4
r109 (  69 70 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=6.28 //y=7.4 //x2=5.57 //y2=7.4
r110 (  63 87 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=5.485 //y=7.23 //x2=5.485 //y2=7.4
r111 (  63 94 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=5.485 //y=7.23 //x2=5.485 //y2=6.405
r112 (  62 85 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=4.98 //y=7.4 //x2=4.81 //y2=7.4
r113 (  61 87 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=5.4 //y=7.4 //x2=5.485 //y2=7.4
r114 (  61 62 ) resistor r=15.0588 //w=0.357 //l=0.42 //layer=li \
 //thickness=0.1 //x=5.4 //y=7.4 //x2=4.98 //y2=7.4
r115 (  56 84 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=3.73 //y2=7.4
r116 (  56 58 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=4.07 //y2=7.4
r117 (  55 85 ) resistor r=5.4201 //w=0.34 //l=0.17 //layer=li //thickness=0.1 \
 //x=4.64 //y=7.4 //x2=4.81 //y2=7.4
r118 (  55 58 ) resistor r=20.437 //w=0.357 //l=0.57 //layer=li \
 //thickness=0.1 //x=4.64 //y=7.4 //x2=4.07 //y2=7.4
r119 (  49 84 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=7.4
r120 (  49 93 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=6.745
r121 (  46 83 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.85 //y2=7.4
r122 (  46 48 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.96 //y2=7.4
r123 (  45 84 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=3.73 //y2=7.4
r124 (  45 48 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=2.96 //y2=7.4
r125 (  39 83 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=7.4
r126 (  39 92 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=6.745
r127 (  38 82 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.055 //y=7.4 //x2=1.97 //y2=7.4
r128 (  37 83 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.85 //y2=7.4
r129 (  37 38 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.055 //y2=7.4
r130 (  31 82 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=7.4
r131 (  31 91 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=6.745
r132 (  28 81 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.09 //y2=7.4
r133 (  28 30 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.85 //y2=7.4
r134 (  27 82 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.97 //y2=7.4
r135 (  27 30 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.85 //y2=7.4
r136 (  21 81 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=7.4
r137 (  21 90 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=6.405
r138 (  17 81 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=1.09 //y2=7.4
r139 (  17 20 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=0.74 //y2=7.4
r140 (  13 89 ) resistor r=4.65 //w=0.17 //l=0.34 //layer=mcon //count=2 \
 //x=6.29 //y=7.4 //x2=6.29 //y2=7.4
r141 (  11 87 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=5.55 //y=7.4 //x2=5.55 //y2=7.4
r142 (  11 13 ) resistor r=0.307309 //w=0.301 //l=0.74 //layer=m1 \
 //thickness=0.36 //x=5.55 //y=7.4 //x2=6.29 //y2=7.4
r143 (  9 58 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=4.07 //y=7.4 //x2=4.07 //y2=7.4
r144 (  9 11 ) resistor r=0.614618 //w=0.301 //l=1.48 //layer=m1 \
 //thickness=0.36 //x=4.07 //y=7.4 //x2=5.55 //y2=7.4
r145 (  7 48 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=2.96 //y=7.4 //x2=2.96 //y2=7.4
r146 (  7 9 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r147 (  5 30 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=1.85 //y=7.4 //x2=1.85 //y2=7.4
r148 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r149 (  2 20 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 \
 //x=0.74 //y=7.4 //x2=0.74 //y2=7.4
r150 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_AND3X1_PCELL\%noxref_2

subckt PM_AND3X1_PCELL\%noxref_3 ( 1 2 13 14 21 29 35 36 40 42 49 50 51 52 53 \
 54 55 56 57 61 62 63 65 71 72 74 82 84 85 86 )
c141 ( 86 0 ) capacitor c=0.023087f //x=3.145 //y=5.02
c142 ( 85 0 ) capacitor c=0.023519f //x=2.265 //y=5.02
c143 ( 84 0 ) capacitor c=0.0224735f //x=1.385 //y=5.02
c144 ( 82 0 ) capacitor c=0.00853354f //x=3.395 //y=0.915
c145 ( 74 0 ) capacitor c=0.0528806f //x=5.55 //y=2.085
c146 ( 72 0 ) capacitor c=0.0435629f //x=6.19 //y=1.255
c147 ( 71 0 ) capacitor c=0.0200386f //x=6.19 //y=0.91
c148 ( 65 0 ) capacitor c=0.0152946f //x=6.035 //y=1.41
c149 ( 63 0 ) capacitor c=0.0157804f //x=6.035 //y=0.755
c150 ( 62 0 ) capacitor c=0.0524167f //x=5.78 //y=4.79
c151 ( 61 0 ) capacitor c=0.0322983f //x=6.07 //y=4.79
c152 ( 57 0 ) capacitor c=0.0290017f //x=5.66 //y=1.92
c153 ( 56 0 ) capacitor c=0.0250027f //x=5.66 //y=1.565
c154 ( 55 0 ) capacitor c=0.0234316f //x=5.66 //y=1.255
c155 ( 54 0 ) capacitor c=0.0200596f //x=5.66 //y=0.91
c156 ( 53 0 ) capacitor c=0.154218f //x=6.145 //y=6.02
c157 ( 52 0 ) capacitor c=0.154243f //x=5.705 //y=6.02
c158 ( 50 0 ) capacitor c=0.0019954f //x=3.29 //y=5.155
c159 ( 49 0 ) capacitor c=0.00424403f //x=2.41 //y=5.155
c160 ( 42 0 ) capacitor c=0.0944546f //x=5.55 //y=2.085
c161 ( 40 0 ) capacitor c=0.114111f //x=4.07 //y=3.33
c162 ( 36 0 ) capacitor c=0.00777616f //x=3.67 //y=1.665
c163 ( 35 0 ) capacitor c=0.018423f //x=3.985 //y=1.665
c164 ( 29 0 ) capacitor c=0.0347121f //x=3.985 //y=5.155
c165 ( 21 0 ) capacitor c=0.0254521f //x=3.205 //y=5.155
c166 ( 14 0 ) capacitor c=0.00549987f //x=1.615 //y=5.155
c167 ( 13 0 ) capacitor c=0.0214591f //x=2.325 //y=5.155
c168 ( 2 0 ) capacitor c=0.0158372f //x=4.185 //y=3.33
c169 ( 1 0 ) capacitor c=0.0799791f //x=5.435 //y=3.33
r170 (  74 75 ) resistor r=17.5563 //w=0.302 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.55 //y=2.085 //x2=5.66 //y2=2.085
r171 (  72 81 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.19 //y=1.255 //x2=6.15 //y2=1.41
r172 (  71 80 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=6.19 //y=0.91 //x2=6.15 //y2=0.755
r173 (  71 72 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=6.19 //y=0.91 //x2=6.19 //y2=1.255
r174 (  66 79 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.815 //y=1.41 //x2=5.7 //y2=1.41
r175 (  65 81 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.035 //y=1.41 //x2=6.15 //y2=1.41
r176 (  64 78 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=5.815 //y=0.755 //x2=5.7 //y2=0.755
r177 (  63 80 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=6.035 //y=0.755 //x2=6.15 //y2=0.755
r178 (  63 64 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=6.035 //y=0.755 //x2=5.815 //y2=0.755
r179 (  61 68 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=6.07 //y=4.79 //x2=6.145 //y2=4.865
r180 (  61 62 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=6.07 //y=4.79 //x2=5.78 //y2=4.79
r181 (  58 62 ) resistor r=23.403 //w=0.284 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=5.705 //y=4.865 //x2=5.78 //y2=4.79
r182 (  58 77 ) resistor r=26.3063 //w=0.284 //l=0.229783 //layer=ply \
 //thickness=0.18 //x=5.705 //y=4.865 //x2=5.55 //y2=4.7
r183 (  57 75 ) resistor r=19.1248 //w=0.302 //l=0.165 //layer=ply \
 //thickness=0.18 //x=5.66 //y=1.92 //x2=5.66 //y2=2.085
r184 (  56 79 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.66 //y=1.565 //x2=5.7 //y2=1.41
r185 (  56 57 ) resistor r=182.032 //w=0.094 //l=0.355 //layer=ply \
 //thickness=0.18 //x=5.66 //y=1.565 //x2=5.66 //y2=1.92
r186 (  55 79 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.66 //y=1.255 //x2=5.7 //y2=1.41
r187 (  54 78 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=5.66 //y=0.91 //x2=5.7 //y2=0.755
r188 (  54 55 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=5.66 //y=0.91 //x2=5.66 //y2=1.255
r189 (  53 68 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=6.145 //y=6.02 //x2=6.145 //y2=4.865
r190 (  52 58 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=5.705 //y=6.02 //x2=5.705 //y2=4.865
r191 (  51 65 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.925 //y=1.41 //x2=6.035 //y2=1.41
r192 (  51 66 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=5.925 //y=1.41 //x2=5.815 //y2=1.41
r193 (  47 77 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.55 //y=4.7 //x2=5.55 //y2=4.7
r194 (  45 47 ) resistor r=93.7754 //w=0.187 //l=1.37 //layer=li \
 //thickness=0.1 //x=5.55 //y=3.33 //x2=5.55 //y2=4.7
r195 (  42 74 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=5.55 //y=2.085 //x2=5.55 //y2=2.085
r196 (  42 45 ) resistor r=85.2193 //w=0.187 //l=1.245 //layer=li \
 //thickness=0.1 //x=5.55 //y=2.085 //x2=5.55 //y2=3.33
r197 (  38 40 ) resistor r=119.102 //w=0.187 //l=1.74 //layer=li \
 //thickness=0.1 //x=4.07 //y=5.07 //x2=4.07 //y2=3.33
r198 (  37 40 ) resistor r=108.15 //w=0.187 //l=1.58 //layer=li \
 //thickness=0.1 //x=4.07 //y=1.75 //x2=4.07 //y2=3.33
r199 (  35 37 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=4.07 //y2=1.75
r200 (  35 36 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=3.67 //y2=1.665
r201 (  31 36 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.67 //y2=1.665
r202 (  31 82 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.585 //y2=1.01
r203 (  30 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.375 //y=5.155 //x2=3.29 //y2=5.155
r204 (  29 38 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=4.07 //y2=5.07
r205 (  29 30 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=3.375 //y2=5.155
r206 (  23 50 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.155
r207 (  23 86 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.725
r208 (  22 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.495 //y=5.155 //x2=2.41 //y2=5.155
r209 (  21 50 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=3.29 //y2=5.155
r210 (  21 22 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=2.495 //y2=5.155
r211 (  15 49 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.155
r212 (  15 85 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.725
r213 (  13 49 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=2.41 //y2=5.155
r214 (  13 14 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.325 //y=5.155 //x2=1.615 //y2=5.155
r215 (  7 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.615 //y2=5.155
r216 (  7 84 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.53 //y2=5.725
r217 (  6 45 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=5.55 //y=3.33 //x2=5.55 //y2=3.33
r218 (  4 40 ) resistor r=9.3 //w=0.17 //l=0.17 //layer=mcon //count=1 \
 //x=4.07 //y=3.33 //x2=4.07 //y2=3.33
r219 (  2 4 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=4.185 //y=3.33 //x2=4.07 //y2=3.33
r220 (  1 6 ) resistor r=0.0717383 //w=0.224 //l=0.115 //layer=m1 \
 //thickness=0.36 //x=5.435 //y=3.33 //x2=5.55 //y2=3.33
r221 (  1 2 ) resistor r=1.19275 //w=0.131 //l=1.25 //layer=m1 \
 //thickness=0.36 //x=5.435 //y=3.33 //x2=4.185 //y2=3.33
ends PM_AND3X1_PCELL\%noxref_3

subckt PM_AND3X1_PCELL\%noxref_4 ( 2 7 8 9 10 11 12 13 14 16 22 23 24 25 )
c55 ( 25 0 ) capacitor c=0.0598646f //x=1.385 //y=4.79
c56 ( 24 0 ) capacitor c=0.0375015f //x=1.675 //y=4.79
c57 ( 23 0 ) capacitor c=0.0347816f //x=1.34 //y=1.22
c58 ( 22 0 ) capacitor c=0.0187487f //x=1.34 //y=0.875
c59 ( 16 0 ) capacitor c=0.0137055f //x=1.185 //y=1.375
c60 ( 14 0 ) capacitor c=0.0149861f //x=1.185 //y=0.72
c61 ( 13 0 ) capacitor c=0.102158f //x=0.81 //y=1.915
c62 ( 12 0 ) capacitor c=0.0229444f //x=0.81 //y=1.53
c63 ( 11 0 ) capacitor c=0.0234352f //x=0.81 //y=1.22
c64 ( 10 0 ) capacitor c=0.0198724f //x=0.81 //y=0.875
c65 ( 9 0 ) capacitor c=0.110114f //x=1.75 //y=6.02
c66 ( 8 0 ) capacitor c=0.158956f //x=1.31 //y=6.02
c67 ( 2 0 ) capacitor c=0.128679f //x=1.11 //y=2.08
r68 (  24 26 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.75 //y2=4.865
r69 (  24 25 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.385 //y2=4.79
r70 (  23 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=1.22 //x2=1.3 //y2=1.375
r71 (  22 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.3 //y2=0.72
r72 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.34 //y2=1.22
r73 (  19 25 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.385 //y2=4.79
r74 (  19 34 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.11 //y2=4.7
r75 (  17 30 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=1.375 //x2=0.85 //y2=1.375
r76 (  16 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=1.375 //x2=1.3 //y2=1.375
r77 (  15 29 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=0.72 //x2=0.85 //y2=0.72
r78 (  14 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=1.3 //y2=0.72
r79 (  14 15 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=0.965 //y2=0.72
r80 (  13 32 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.915 //x2=1.11 //y2=2.08
r81 (  12 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.85 //y2=1.375
r82 (  12 13 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.81 //y2=1.915
r83 (  11 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.22 //x2=0.85 //y2=1.375
r84 (  10 29 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.85 //y2=0.72
r85 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.81 //y2=1.22
r86 (  9 26 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.75 //y=6.02 //x2=1.75 //y2=4.865
r87 (  8 19 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.31 //y=6.02 //x2=1.31 //y2=4.865
r88 (  7 16 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=1.185 //y2=1.375
r89 (  7 17 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=0.965 //y2=1.375
r90 (  5 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r91 (  2 32 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r92 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=4.7
ends PM_AND3X1_PCELL\%noxref_4

subckt PM_AND3X1_PCELL\%noxref_5 ( 2 7 8 9 10 11 12 14 20 21 22 23 24 32 )
c70 ( 32 0 ) capacitor c=0.0354872f //x=2.22 //y=4.7
c71 ( 24 0 ) capacitor c=0.0307682f //x=2.555 //y=4.79
c72 ( 23 0 ) capacitor c=0.0850619f //x=2.31 //y=1.915
c73 ( 22 0 ) capacitor c=0.0170266f //x=2.31 //y=1.45
c74 ( 21 0 ) capacitor c=0.018609f //x=2.31 //y=1.22
c75 ( 20 0 ) capacitor c=0.0187309f //x=2.31 //y=0.91
c76 ( 14 0 ) capacitor c=0.014725f //x=2.155 //y=1.375
c77 ( 12 0 ) capacitor c=0.0146567f //x=2.155 //y=0.755
c78 ( 11 0 ) capacitor c=0.0335408f //x=1.785 //y=1.22
c79 ( 10 0 ) capacitor c=0.0173761f //x=1.785 //y=0.91
c80 ( 9 0 ) capacitor c=0.110114f //x=2.63 //y=6.02
c81 ( 8 0 ) capacitor c=0.11012f //x=2.19 //y=6.02
c82 ( 2 0 ) capacitor c=0.106476f //x=2.22 //y=2.08
r83 (  34 35 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.79 //x2=2.22 //y2=4.865
r84 (  32 34 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.7 //x2=2.22 //y2=4.79
r85 (  25 34 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.355 //y=4.79 //x2=2.22 //y2=4.79
r86 (  24 26 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.63 //y2=4.865
r87 (  24 25 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.355 //y2=4.79
r88 (  23 39 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.915 //x2=2.235 //y2=2.08
r89 (  22 37 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.27 //y2=1.375
r90 (  22 23 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.31 //y2=1.915
r91 (  21 37 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.22 //x2=2.27 //y2=1.375
r92 (  20 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.27 //y2=0.755
r93 (  20 21 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.31 //y2=1.22
r94 (  15 30 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=1.375 //x2=1.825 //y2=1.375
r95 (  14 37 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=1.375 //x2=2.27 //y2=1.375
r96 (  13 29 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=0.755 //x2=1.825 //y2=0.755
r97 (  12 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=2.27 //y2=0.755
r98 (  12 13 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=1.94 //y2=0.755
r99 (  11 30 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=1.22 //x2=1.825 //y2=1.375
r100 (  10 29 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.825 //y2=0.755
r101 (  10 11 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.785 //y2=1.22
r102 (  9 26 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.63 //y=6.02 //x2=2.63 //y2=4.865
r103 (  8 35 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.19 //y=6.02 //x2=2.19 //y2=4.865
r104 (  7 14 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=2.155 //y2=1.375
r105 (  7 15 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=1.94 //y2=1.375
r106 (  5 32 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=4.7 //x2=2.22 //y2=4.7
r107 (  2 39 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=2.08
r108 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=4.7
ends PM_AND3X1_PCELL\%noxref_5

subckt PM_AND3X1_PCELL\%noxref_6 ( 1 5 9 13 17 35 )
c45 ( 35 0 ) capacitor c=0.0747858f //x=0.455 //y=0.375
c46 ( 17 0 ) capacitor c=0.0266691f //x=2.445 //y=1.59
c47 ( 13 0 ) capacitor c=0.0156939f //x=2.445 //y=0.54
c48 ( 9 0 ) capacitor c=0.00678203f //x=1.56 //y=0.625
c49 ( 5 0 ) capacitor c=0.0236189f //x=1.475 //y=1.59
c50 ( 1 0 ) capacitor c=0.0109947f //x=0.59 //y=1.505
r51 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=1.59 //x2=1.56 //y2=1.63
r52 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=1.59 //x2=2.045 //y2=1.59
r53 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=1.59 //x2=2.53 //y2=1.59
r54 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=1.59 //x2=2.045 //y2=1.59
r55 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=0.54 //x2=1.56 //y2=0.5
r56 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=0.54 //x2=2.045 //y2=0.54
r57 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=0.54 //x2=2.53 //y2=0.54
r58 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=0.54 //x2=2.045 //y2=0.54
r59 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=1.63
r60 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=0.89
r61 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.5
r62 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.89
r63 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.675 //y=1.59 //x2=0.59 //y2=1.63
r64 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.675 //y=1.59 //x2=1.075 //y2=1.59
r65 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.475 //y=1.59 //x2=1.56 //y2=1.63
r66 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.475 //y=1.59 //x2=1.075 //y2=1.59
r67 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.59 //y=1.505 //x2=0.59 //y2=1.63
r68 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.59 //y=1.505 //x2=0.59 //y2=0.89
ends PM_AND3X1_PCELL\%noxref_6

subckt PM_AND3X1_PCELL\%noxref_7 ( 2 7 8 9 13 14 15 20 22 25 26 28 29 34 )
c54 ( 34 0 ) capacitor c=0.0672371f //x=3.33 //y=4.7
c55 ( 29 0 ) capacitor c=0.0273931f //x=3.33 //y=1.915
c56 ( 28 0 ) capacitor c=0.0471168f //x=3.33 //y=2.08
c57 ( 26 0 ) capacitor c=0.0432517f //x=3.85 //y=1.26
c58 ( 25 0 ) capacitor c=0.0200379f //x=3.85 //y=0.915
c59 ( 22 0 ) capacitor c=0.0158629f //x=3.695 //y=1.415
c60 ( 20 0 ) capacitor c=0.0157803f //x=3.695 //y=0.76
c61 ( 15 0 ) capacitor c=0.0218028f //x=3.32 //y=1.57
c62 ( 14 0 ) capacitor c=0.0207459f //x=3.32 //y=1.26
c63 ( 13 0 ) capacitor c=0.0194308f //x=3.32 //y=0.915
c64 ( 9 0 ) capacitor c=0.158794f //x=3.51 //y=6.02
c65 ( 8 0 ) capacitor c=0.110114f //x=3.07 //y=6.02
c66 ( 2 0 ) capacitor c=0.095837f //x=3.33 //y=2.08
r67 (  28 29 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.33 //y=2.08 //x2=3.33 //y2=1.915
r68 (  26 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=1.26 //x2=3.81 //y2=1.415
r69 (  25 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.81 //y2=0.76
r70 (  25 26 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.85 //y2=1.26
r71 (  23 32 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=1.415 //x2=3.36 //y2=1.415
r72 (  22 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=1.415 //x2=3.81 //y2=1.415
r73 (  21 31 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=0.76 //x2=3.36 //y2=0.76
r74 (  20 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.81 //y2=0.76
r75 (  20 21 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.475 //y2=0.76
r76 (  17 34 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=3.51 //y=4.865 //x2=3.33 //y2=4.7
r77 (  15 32 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.36 //y2=1.415
r78 (  15 29 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.32 //y2=1.915
r79 (  14 32 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.26 //x2=3.36 //y2=1.415
r80 (  13 31 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.36 //y2=0.76
r81 (  13 14 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.32 //y2=1.26
r82 (  10 34 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=3.07 //y=4.865 //x2=3.33 //y2=4.7
r83 (  9 17 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.51 //y=6.02 //x2=3.51 //y2=4.865
r84 (  8 10 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.07 //y=6.02 //x2=3.07 //y2=4.865
r85 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.695 //y2=1.415
r86 (  7 23 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.475 //y2=1.415
r87 (  5 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r88 (  2 28 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r89 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=4.7
ends PM_AND3X1_PCELL\%noxref_7

subckt PM_AND3X1_PCELL\%noxref_8 ( 1 3 11 15 25 28 29 )
c54 ( 29 0 ) capacitor c=0.0456206f //x=2.965 //y=0.375
c55 ( 28 0 ) capacitor c=0.00467097f //x=1.86 //y=0.91
c56 ( 25 0 ) capacitor c=0.00156479f //x=3.1 //y=0.995
c57 ( 15 0 ) capacitor c=0.00737666f //x=4.07 //y=0.625
c58 ( 11 0 ) capacitor c=0.0152819f //x=3.985 //y=0.54
c59 ( 3 0 ) capacitor c=0.00718386f //x=3.1 //y=0.625
c60 ( 1 0 ) capacitor c=0.0279585f //x=3.015 //y=0.995
r61 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.5
r62 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.89
r63 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.185 //y=0.54 //x2=3.1 //y2=0.5
r64 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.185 //y=0.54 //x2=3.585 //y2=0.54
r65 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.985 //y=0.54 //x2=4.07 //y2=0.5
r66 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.985 //y=0.54 //x2=3.585 //y2=0.54
r67 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=0.995
r68 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=1.23
r69 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.995
r70 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.89
r71 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.5
r72 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.89
r73 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.135 //y=0.995 //x2=2.05 //y2=0.995
r74 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=3.1 //y2=0.995
r75 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=2.135 //y2=0.995
ends PM_AND3X1_PCELL\%noxref_8

subckt PM_AND3X1_PCELL\%noxref_9 ( 11 12 13 14 16 17 19 )
c44 ( 19 0 ) capacitor c=0.028734f //x=5.78 //y=5.02
c45 ( 17 0 ) capacitor c=0.0173218f //x=5.735 //y=0.91
c46 ( 16 0 ) capacitor c=0.105613f //x=6.29 //y=4.495
c47 ( 14 0 ) capacitor c=0.00575887f //x=6.01 //y=4.58
c48 ( 13 0 ) capacitor c=0.0136889f //x=6.205 //y=4.58
c49 ( 12 0 ) capacitor c=0.00636159f //x=6.005 //y=2.08
c50 ( 11 0 ) capacitor c=0.0140707f //x=6.205 //y=2.08
r51 (  15 16 ) resistor r=159.487 //w=0.187 //l=2.33 //layer=li \
 //thickness=0.1 //x=6.29 //y=2.165 //x2=6.29 //y2=4.495
r52 (  13 16 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.205 //y=4.58 //x2=6.29 //y2=4.495
r53 (  13 14 ) resistor r=13.3476 //w=0.187 //l=0.195 //layer=li \
 //thickness=0.1 //x=6.205 //y=4.58 //x2=6.01 //y2=4.58
r54 (  11 15 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=6.205 //y=2.08 //x2=6.29 //y2=2.165
r55 (  11 12 ) resistor r=13.6898 //w=0.187 //l=0.2 //layer=li //thickness=0.1 \
 //x=6.205 //y=2.08 //x2=6.005 //y2=2.08
r56 (  5 14 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5.925 //y=4.665 //x2=6.01 //y2=4.58
r57 (  5 19 ) resistor r=72.5562 //w=0.187 //l=1.06 //layer=li //thickness=0.1 \
 //x=5.925 //y=4.665 //x2=5.925 //y2=5.725
r58 (  1 12 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=5.92 //y=1.995 //x2=6.005 //y2=2.08
r59 (  1 17 ) resistor r=67.7647 //w=0.187 //l=0.99 //layer=li //thickness=0.1 \
 //x=5.92 //y=1.995 //x2=5.92 //y2=1.005
ends PM_AND3X1_PCELL\%noxref_9

