magic
tech sky130A
magscale 1 2
timestamp 1652455925
<< nwell >>
rect 57 1463 91 1497
rect 31 822 117 884
<< pwell >>
rect -34 -34 182 544
<< psubdiff >>
rect 34 482 114 544
rect 34 -17 57 17
rect 91 -17 114 17
rect 34 -34 114 -17
<< nsubdiff >>
rect 34 1497 114 1514
rect 34 1463 57 1497
rect 91 1463 114 1497
rect 34 822 114 884
<< psubdiffcont >>
rect 57 -17 91 17
<< nsubdiffcont >>
rect 57 1463 91 1497
<< locali >>
rect 34 1497 114 1514
rect 34 1463 57 1497
rect 91 1463 114 1497
rect 34 1446 114 1463
rect 34 17 114 34
rect 34 -17 57 17
rect 91 -17 114 17
rect 34 -34 114 -17
<< metal1 >>
rect -34 1446 182 1514
rect -34 -34 182 34
use diff_ring_side  diff_ring_side_0 pcells
timestamp 1652319726
transform 1 0 0 0 1 0
box -87 -34 87 1550
use diff_ring_side  diff_ring_side_1
timestamp 1652319726
transform 1 0 148 0 1 0
box -87 -34 87 1550
<< labels >>
rlabel metal1 -34 1446 182 1514 1 VPWR
port 1 nsew power bidirectional abutment
rlabel metal1 -34 -34 182 34 1 VGND
port 2 nsew ground bidirectional abutment
rlabel nwell 57 1463 91 1497 1 VPB
port 3 nsew power bidirectional
rlabel pwell 57 -17 91 17 1 VNB
port 4 nsew ground bidirectional
<< properties >>
string LEFclass CORE SPACER
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
