* SPICE3 file created from TMRDFFSNRNQX1.ext - technology: sky130A

.subckt TMRDFFSNRNQX1 Q D CLK SN RN VDD GND
X0 VDD RN a_277_1004 VDD pshort w=2 l=0.15 M=2
X1 GND a_7973_1004 a_8749_75 GND nshort w=3 l=0.15
X2 a_6371_943 a_6049_1004 VDD VDD pshort w=2 l=0.15 M=2
X3 VDD a_7973_1004 a_7333_943 VDD pshort w=2 l=0.15 M=2
X4 VDD a_9897_1004 a_10219_943 VDD pshort w=2 l=0.15 M=2
X5 a_17533_1005 a_4447_943 VDD VDD pshort w=2 l=0.15 M=2
X6 a_12143_943 CLK VDD VDD pshort w=2 l=0.15 M=2
X7 GND D a_91_75 GND nshort w=3 l=0.15
X8 a_15991_943 a_15669_1004 VDD VDD pshort w=2 l=0.15 M=2
X9 a_599_943 a_1561_943 VDD VDD pshort w=2 l=0.15 M=2
X10 VDD RN a_1561_943 VDD pshort w=2 l=0.15 M=2
X11 a_11916_182 RN a_11635_75 GND nshort w=3 l=0.15
X12 a_9897_1004 a_6371_943 VDD VDD pshort w=2 l=0.15 M=2
X13 a_4125_1004 a_599_943 VDD VDD pshort w=2 l=0.15 M=2
X14 a_9992_182 RN a_9711_75 GND nshort w=3 l=0.15
X15 VDD SN a_2201_1004 VDD pshort w=2 l=0.15 M=2
X16 a_4125_1004 a_4447_943 VDD VDD pshort w=2 l=0.15 M=2
X17 GND a_4447_943 a_17428_73 GND nshort w=3 l=0.15
X18 VDD a_6371_943 a_6049_1004 VDD pshort w=2 l=0.15 M=2
X19 a_18197_1005 a_4447_943 a_17533_1005 VDD pshort w=2 l=0.15 M=2
X20 a_1561_943 CLK VDD VDD pshort w=2 l=0.15 M=2
X21 GND a_11821_1004 a_13559_75 GND nshort w=3 l=0.15
X22 GND a_12143_943 a_15483_75 GND nshort w=3 l=0.15
X23 VDD a_599_943 a_277_1004 VDD pshort w=2 l=0.15 M=2
X24 a_13745_1004 SN VDD VDD pshort w=2 l=0.15 M=2
X25 a_17533_1005 a_10219_943 VDD VDD pshort w=2 l=0.15 M=2
X26 a_12143_943 a_11821_1004 VDD VDD pshort w=2 l=0.15 M=2
X27 a_14802_182 CLK a_14521_75 GND nshort w=3 l=0.15
X28 VDD a_13745_1004 a_13105_943 VDD pshort w=2 l=0.15 M=2
X29 a_17708_181 a_15991_943 a_18094_73 GND nshort w=3 l=0.15
X30 a_10954_182 SN a_10673_75 GND nshort w=3 l=0.15
X31 a_15991_943 SN VDD VDD pshort w=2 l=0.15 M=2
X32 a_16726_182 SN a_16445_75 GND nshort w=3 l=0.15
X33 a_12878_182 CLK a_12597_75 GND nshort w=3 l=0.15
X34 a_15669_1004 a_12143_943 VDD VDD pshort w=2 l=0.15 M=2
X35 VDD a_1561_943 a_2201_1004 VDD pshort w=2 l=0.15 M=2
X36 a_4125_1004 RN VDD VDD pshort w=2 l=0.15 M=2
X37 VDD RN a_6049_1004 VDD pshort w=2 l=0.15 M=2
X38 a_7973_1004 a_7333_943 VDD VDD pshort w=2 l=0.15 M=2
X39 a_9897_1004 a_10219_943 VDD VDD pshort w=2 l=0.15 M=2
X40 GND a_15669_1004 a_16445_75 GND nshort w=3 l=0.15
X41 VDD a_13105_943 a_15991_943 VDD pshort w=2 l=0.15 M=2
X42 a_1561_943 a_2201_1004 VDD VDD pshort w=2 l=0.15 M=2
X43 a_2201_1004 a_1561_943 a_2296_182 GND nshort w=3 l=0.15
X44 a_372_182 RN a_91_75 GND nshort w=3 l=0.15
X45 a_18197_1005 a_15991_943 a_17533_1005 VDD pshort w=2 l=0.15 M=2
X46 VDD a_4125_1004 a_4447_943 VDD pshort w=2 l=0.15 M=2
X47 a_6371_943 CLK VDD VDD pshort w=2 l=0.15 M=2
X48 a_4125_1004 a_4447_943 a_4220_182 GND nshort w=3 l=0.15
X49 VDD CLK a_7333_943 VDD pshort w=2 l=0.15 M=2
X50 a_6049_1004 D VDD VDD pshort w=2 l=0.15 M=2
X51 a_17708_181 a_10219_943 a_18197_1005 VDD pshort w=2 l=0.15 M=2
X52 a_13840_182 SN a_13559_75 GND nshort w=3 l=0.15
X53 a_277_1004 D VDD VDD pshort w=2 l=0.15 M=2
X54 a_15764_182 RN a_15483_75 GND nshort w=3 l=0.15
X55 VDD CLK a_13105_943 VDD pshort w=2 l=0.15 M=2
X56 a_10219_943 a_7333_943 VDD VDD pshort w=2 l=0.15 M=2
X57 VDD a_11821_1004 a_13745_1004 VDD pshort w=2 l=0.15 M=2
X58 VDD a_13105_943 a_12143_943 VDD pshort w=2 l=0.15 M=2
X59 a_15669_1004 RN VDD VDD pshort w=2 l=0.15 M=2
X60 VDD a_277_1004 a_599_943 VDD pshort w=2 l=0.15 M=2
X61 a_9897_1004 RN VDD VDD pshort w=2 l=0.15 M=2
X62 VDD RN a_11821_1004 VDD pshort w=2 l=0.15 M=2
X63 GND a_277_1004 a_2015_75 GND nshort w=3 l=0.15
X64 a_599_943 a_1561_943 a_1334_182 GND nshort w=3 l=0.15
X65 Q a_17708_181 GND GND nshort w=3 l=0.15
X66 a_6371_943 a_7333_943 a_7106_182 GND nshort w=3 l=0.15
X67 a_13745_1004 a_13105_943 VDD VDD pshort w=2 l=0.15 M=2
X68 VDD SN a_4447_943 VDD pshort w=2 l=0.15 M=2
X69 a_1561_943 RN a_3258_182 GND nshort w=3 l=0.15
X70 a_18197_1005 a_15991_943 a_17708_181 VDD pshort w=2 l=0.15 M=2
X71 VDD a_15991_943 a_15669_1004 VDD pshort w=2 l=0.15 M=2
X72 a_6371_943 a_7333_943 VDD VDD pshort w=2 l=0.15 M=2
X73 Q a_17708_181 VDD VDD pshort w=2 l=0.15 M=2
X74 VDD RN a_7333_943 VDD pshort w=2 l=0.15 M=2
X75 a_4447_943 a_1561_943 a_5182_182 GND nshort w=3 l=0.15
X76 VDD SN a_7973_1004 VDD pshort w=2 l=0.15 M=2
X77 a_11821_1004 a_12143_943 a_11916_182 GND nshort w=3 l=0.15
X78 a_17708_181 a_10219_943 a_17428_73 GND nshort w=3 l=0.15
X79 a_6049_1004 a_6371_943 a_6144_182 GND nshort w=3 l=0.15
X80 VDD CLK a_599_943 VDD pshort w=2 l=0.15 M=2
X81 a_9897_1004 a_10219_943 a_9992_182 GND nshort w=3 l=0.15
X82 VDD a_12143_943 a_11821_1004 VDD pshort w=2 l=0.15 M=2
X83 a_7973_1004 a_7333_943 a_8068_182 GND nshort w=3 l=0.15
X84 GND a_2201_1004 a_2977_75 GND nshort w=3 l=0.15
X85 VDD a_1561_943 a_4447_943 VDD pshort w=2 l=0.15 M=2
X86 GND a_277_1004 a_1053_75 GND nshort w=3 l=0.15
X87 VDD a_6049_1004 a_7973_1004 VDD pshort w=2 l=0.15 M=2
X88 VDD RN a_13105_943 VDD pshort w=2 l=0.15 M=2
X89 a_4220_182 RN a_3939_75 GND nshort w=3 l=0.15
X90 a_11821_1004 D VDD VDD pshort w=2 l=0.15 M=2
X91 a_10219_943 a_7333_943 a_10954_182 GND nshort w=3 l=0.15
X92 a_2296_182 SN a_2015_75 GND nshort w=3 l=0.15
X93 a_12143_943 a_13105_943 a_12878_182 GND nshort w=3 l=0.15
X94 a_13105_943 RN a_14802_182 GND nshort w=3 l=0.15
X95 GND a_599_943 a_3939_75 GND nshort w=3 l=0.15
X96 a_2201_1004 a_277_1004 VDD VDD pshort w=2 l=0.15 M=2
X97 a_7333_943 RN a_9030_182 GND nshort w=3 l=0.15
X98 a_5182_182 SN a_4901_75 GND nshort w=3 l=0.15
X99 a_15669_1004 a_15991_943 a_15764_182 GND nshort w=3 l=0.15
X100 a_7106_182 CLK a_6825_75 GND nshort w=3 l=0.15
X101 a_1334_182 CLK a_1053_75 GND nshort w=3 l=0.15
X102 a_3258_182 CLK a_2977_75 GND nshort w=3 l=0.15
X103 a_13745_1004 a_13105_943 a_13840_182 GND nshort w=3 l=0.15
X104 GND a_6049_1004 a_6825_75 GND nshort w=3 l=0.15
X105 VDD SN a_10219_943 VDD pshort w=2 l=0.15 M=2
X106 GND a_4125_1004 a_4901_75 GND nshort w=3 l=0.15
X107 GND a_15991_943 a_18760_73 GND nshort w=3 l=0.15
X108 GND a_4447_943 a_18094_73 GND nshort w=3 l=0.15
X109 a_6144_182 RN a_5863_75 GND nshort w=3 l=0.15
X110 GND D a_11635_75 GND nshort w=3 l=0.15
X111 a_15991_943 a_13105_943 a_16726_182 GND nshort w=3 l=0.15
X112 a_8068_182 SN a_7787_75 GND nshort w=3 l=0.15
X113 GND a_6049_1004 a_7787_75 GND nshort w=3 l=0.15
X114 GND a_6371_943 a_9711_75 GND nshort w=3 l=0.15
X115 a_17708_181 a_10219_943 a_18760_73 GND nshort w=3 l=0.15
X116 GND D a_5863_75 GND nshort w=3 l=0.15
X117 a_277_1004 a_599_943 a_372_182 GND nshort w=3 l=0.15
X118 a_9030_182 CLK a_8749_75 GND nshort w=3 l=0.15
X119 GND a_11821_1004 a_12597_75 GND nshort w=3 l=0.15
X120 GND a_13745_1004 a_14521_75 GND nshort w=3 l=0.15
X121 GND a_9897_1004 a_10673_75 GND nshort w=3 l=0.15
C0 SN a_12143_943 3.98fF
C1 VDD a_277_1004 2.25fF
C2 VDD a_6049_1004 2.38fF
C3 VDD a_10219_943 4.07fF
C4 VDD CLK 5.12fF
C5 VDD D 3.63fF
C6 VDD a_7333_943 2.66fF
C7 VDD a_1561_943 2.66fF
C8 a_6371_943 a_7333_943 3.19fF
C9 VDD a_15991_943 2.64fF
C10 a_6371_943 SN 3.98fF
C11 VDD a_599_943 2.45fF
C12 VDD RN 2.54fF
C13 VDD a_2201_1004 2.07fF
C14 a_13105_943 a_12143_943 3.19fF
C15 VDD a_4447_943 6.41fF
C16 VDD a_4125_1004 2.07fF
C17 VDD a_13745_1004 2.07fF
C18 VDD a_12143_943 2.46fF
C19 a_10219_943 CLK 3.10fF
C20 VDD a_7973_1004 2.07fF
C21 VDD a_13105_943 2.67fF
C22 VDD a_11821_1004 2.38fF
C23 D CLK 11.68fF
C24 a_10219_943 SN 3.07fF
C25 D a_7333_943 4.46fF
C26 D a_1561_943 4.46fF
C27 CLK SN 2.43fF
C28 D SN 2.38fF
C29 RN CLK 2.23fF
C30 a_10219_943 a_4447_943 5.28fF
C31 RN D 2.04fF
C32 a_599_943 a_1561_943 3.19fF
C33 VDD a_6371_943 2.46fF
C34 CLK a_4447_943 10.85fF
C35 a_599_943 SN 2.03fF
C36 D a_4447_943 3.08fF
C37 RN SN 5.64fF
C38 a_10219_943 a_12143_943 2.04fF
C39 SN a_4447_943 3.24fF
C40 VDD a_15669_1004 2.09fF
C41 a_9897_1004 VDD 2.07fF
C42 a_10219_943 a_13105_943 4.45fF
C43 SN GND 4.14fF
C44 RN GND 5.23fF
C45 VDD GND 46.80fF
.ends
