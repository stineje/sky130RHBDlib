magic
tech sky130A
magscale 1 2
timestamp 1651250934
<< nwell >>
rect -84 832 4376 1575
<< nmos >>
rect 147 318 177 379
tri 177 318 193 334 sw
rect 447 318 477 379
rect 147 288 253 318
tri 253 288 283 318 sw
rect 147 187 177 288
tri 177 272 193 288 nw
tri 237 272 253 288 ne
tri 177 187 193 203 sw
tri 237 187 253 203 se
rect 253 187 283 288
tri 342 288 372 318 se
rect 372 288 477 318
rect 342 194 372 288
tri 372 272 388 288 nw
tri 431 272 447 288 ne
tri 372 194 388 210 sw
tri 431 194 447 210 se
rect 447 194 477 288
tri 147 157 177 187 ne
rect 177 157 253 187
tri 253 157 283 187 nw
tri 342 164 372 194 ne
rect 372 164 447 194
tri 447 164 477 194 nw
rect 649 326 679 379
tri 679 326 695 342 sw
rect 649 296 755 326
tri 755 296 785 326 sw
rect 649 195 679 296
tri 679 280 695 296 nw
tri 739 280 755 296 ne
tri 679 195 695 211 sw
tri 739 195 755 211 se
rect 755 195 785 296
tri 649 165 679 195 ne
rect 679 165 755 195
tri 755 165 785 195 nw
rect 1130 316 1160 377
tri 1160 316 1176 332 sw
rect 1324 324 1354 377
tri 1354 324 1370 340 sw
rect 1130 286 1236 316
tri 1236 286 1266 316 sw
rect 1324 294 1430 324
tri 1430 294 1460 324 sw
rect 1130 185 1160 286
tri 1160 270 1176 286 nw
tri 1220 270 1236 286 ne
tri 1160 185 1176 201 sw
tri 1220 185 1236 201 se
rect 1236 185 1266 286
rect 1324 193 1354 294
tri 1354 278 1370 294 nw
tri 1414 278 1430 294 ne
tri 1354 193 1370 209 sw
tri 1414 193 1430 209 se
rect 1430 193 1460 294
tri 1130 155 1160 185 ne
rect 1160 155 1236 185
tri 1236 155 1266 185 nw
tri 1324 163 1354 193 ne
rect 1354 163 1430 193
tri 1430 163 1460 193 nw
rect 1796 316 1826 377
tri 1826 316 1842 332 sw
rect 1990 324 2020 377
tri 2020 324 2036 340 sw
rect 1796 286 1902 316
tri 1902 286 1932 316 sw
rect 1990 294 2096 324
tri 2096 294 2126 324 sw
rect 1796 185 1826 286
tri 1826 270 1842 286 nw
tri 1886 270 1902 286 ne
tri 1826 185 1842 201 sw
tri 1886 185 1902 201 se
rect 1902 185 1932 286
rect 1990 193 2020 294
tri 2020 278 2036 294 nw
tri 2080 278 2096 294 ne
tri 2020 193 2036 209 sw
tri 2080 193 2096 209 se
rect 2096 193 2126 294
tri 1796 155 1826 185 ne
rect 1826 155 1902 185
tri 1902 155 1932 185 nw
tri 1990 163 2020 193 ne
rect 2020 163 2096 193
tri 2096 163 2126 193 nw
rect 2462 316 2492 377
tri 2492 316 2508 332 sw
rect 2656 324 2686 377
tri 2686 324 2702 340 sw
rect 2462 286 2568 316
tri 2568 286 2598 316 sw
rect 2656 294 2762 324
tri 2762 294 2792 324 sw
rect 2462 185 2492 286
tri 2492 270 2508 286 nw
tri 2552 270 2568 286 ne
tri 2492 185 2508 201 sw
tri 2552 185 2568 201 se
rect 2568 185 2598 286
rect 2656 193 2686 294
tri 2686 278 2702 294 nw
tri 2746 278 2762 294 ne
tri 2686 193 2702 209 sw
tri 2746 193 2762 209 se
rect 2762 193 2792 294
tri 2462 155 2492 185 ne
rect 2492 155 2568 185
tri 2568 155 2598 185 nw
tri 2656 163 2686 193 ne
rect 2686 163 2762 193
tri 2762 163 2792 193 nw
rect 3128 316 3158 377
tri 3158 316 3174 332 sw
rect 3322 324 3352 377
tri 3352 324 3368 340 sw
rect 3128 286 3234 316
tri 3234 286 3264 316 sw
rect 3322 294 3428 324
tri 3428 294 3458 324 sw
rect 3128 185 3158 286
tri 3158 270 3174 286 nw
tri 3218 270 3234 286 ne
tri 3158 185 3174 201 sw
tri 3218 185 3234 201 se
rect 3234 185 3264 286
rect 3322 193 3352 294
tri 3352 278 3368 294 nw
tri 3412 278 3428 294 ne
tri 3352 193 3368 209 sw
tri 3412 193 3428 209 se
rect 3428 193 3458 294
tri 3128 155 3158 185 ne
rect 3158 155 3234 185
tri 3234 155 3264 185 nw
tri 3322 163 3352 193 ne
rect 3352 163 3428 193
tri 3428 163 3458 193 nw
rect 3794 316 3824 377
tri 3824 316 3840 332 sw
rect 3988 324 4018 377
tri 4018 324 4034 340 sw
rect 3794 286 3900 316
tri 3900 286 3930 316 sw
rect 3988 294 4094 324
tri 4094 294 4124 324 sw
rect 3794 185 3824 286
tri 3824 270 3840 286 nw
tri 3884 270 3900 286 ne
tri 3824 185 3840 201 sw
tri 3884 185 3900 201 se
rect 3900 185 3930 286
rect 3988 193 4018 294
tri 4018 278 4034 294 nw
tri 4078 278 4094 294 ne
tri 4018 193 4034 209 sw
tri 4078 193 4094 209 se
rect 4094 193 4124 294
tri 3794 155 3824 185 ne
rect 3824 155 3900 185
tri 3900 155 3930 185 nw
tri 3988 163 4018 193 ne
rect 4018 163 4094 193
tri 4094 163 4124 193 nw
<< pmos >>
rect 247 1050 277 1450
rect 335 1050 365 1450
rect 423 1050 453 1450
rect 511 1050 541 1450
rect 599 1050 629 1450
rect 687 1050 717 1450
rect 1149 1050 1179 1450
rect 1237 1050 1267 1450
rect 1325 1050 1355 1450
rect 1413 1050 1443 1450
rect 1815 1050 1845 1450
rect 1903 1050 1933 1450
rect 1991 1050 2021 1450
rect 2079 1050 2109 1450
rect 2481 1050 2511 1450
rect 2569 1050 2599 1450
rect 2657 1050 2687 1450
rect 2745 1050 2775 1450
rect 3147 1050 3177 1450
rect 3235 1050 3265 1450
rect 3323 1050 3353 1450
rect 3411 1050 3441 1450
rect 3813 1050 3843 1450
rect 3901 1050 3931 1450
rect 3989 1050 4019 1450
rect 4077 1050 4107 1450
<< ndiff >>
rect 91 363 147 379
rect 91 329 101 363
rect 135 329 147 363
rect 91 291 147 329
rect 177 363 447 379
rect 177 334 198 363
tri 177 318 193 334 ne
rect 193 329 198 334
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 447 363
rect 193 318 447 329
rect 477 363 533 379
rect 477 329 489 363
rect 523 329 533 363
rect 91 257 101 291
rect 135 257 147 291
tri 253 288 283 318 ne
rect 283 291 342 318
rect 91 223 147 257
rect 91 189 101 223
rect 135 189 147 223
rect 91 157 147 189
tri 177 272 193 288 se
rect 193 272 237 288
tri 237 272 253 288 sw
rect 177 238 253 272
rect 177 204 198 238
rect 232 204 253 238
rect 177 203 253 204
tri 177 187 193 203 ne
rect 193 187 237 203
tri 237 187 253 203 nw
rect 283 257 295 291
rect 329 257 342 291
tri 342 288 372 318 nw
rect 283 223 342 257
rect 283 189 295 223
rect 329 189 342 223
tri 372 272 388 288 se
rect 388 272 431 288
tri 431 272 447 288 sw
rect 372 244 447 272
rect 372 210 393 244
rect 427 210 447 244
tri 372 194 388 210 ne
rect 388 194 431 210
tri 431 194 447 210 nw
tri 147 157 177 187 sw
tri 253 157 283 187 se
rect 283 164 342 189
tri 342 164 372 194 sw
tri 447 164 477 194 se
rect 477 164 533 329
rect 283 157 533 164
rect 91 153 533 157
rect 91 119 101 153
rect 135 119 295 153
rect 329 119 392 153
rect 426 119 489 153
rect 523 119 533 153
rect 91 103 533 119
rect 593 363 649 379
rect 593 329 603 363
rect 637 329 649 363
rect 593 291 649 329
rect 679 342 841 379
tri 679 326 695 342 ne
rect 695 326 841 342
tri 755 296 785 326 ne
rect 593 257 603 291
rect 637 257 649 291
rect 593 223 649 257
rect 593 189 603 223
rect 637 189 649 223
tri 679 280 695 296 se
rect 695 280 739 296
tri 739 280 755 296 sw
rect 679 247 755 280
rect 679 213 700 247
rect 734 213 755 247
rect 679 211 755 213
tri 679 195 695 211 ne
rect 695 195 739 211
tri 739 195 755 211 nw
rect 785 291 841 326
rect 785 257 797 291
rect 831 257 841 291
rect 785 223 841 257
rect 593 165 649 189
tri 649 165 679 195 sw
tri 755 165 785 195 se
rect 785 189 797 223
rect 831 189 841 223
rect 785 165 841 189
rect 593 153 841 165
rect 593 119 603 153
rect 637 119 700 153
rect 734 119 797 153
rect 831 119 841 153
rect 593 103 841 119
rect 1074 361 1130 377
rect 1074 327 1084 361
rect 1118 327 1130 361
rect 1074 289 1130 327
rect 1160 361 1324 377
rect 1160 332 1181 361
tri 1160 316 1176 332 ne
rect 1176 327 1181 332
rect 1215 327 1278 361
rect 1312 327 1324 361
rect 1176 316 1324 327
rect 1354 340 1516 377
tri 1354 324 1370 340 ne
rect 1370 324 1516 340
rect 1074 255 1084 289
rect 1118 255 1130 289
tri 1236 286 1266 316 ne
rect 1266 289 1324 316
tri 1430 294 1460 324 ne
rect 1074 221 1130 255
rect 1074 187 1084 221
rect 1118 187 1130 221
rect 1074 155 1130 187
tri 1160 270 1176 286 se
rect 1176 270 1220 286
tri 1220 270 1236 286 sw
rect 1160 236 1236 270
rect 1160 202 1181 236
rect 1215 202 1236 236
rect 1160 201 1236 202
tri 1160 185 1176 201 ne
rect 1176 185 1220 201
tri 1220 185 1236 201 nw
rect 1266 255 1278 289
rect 1312 255 1324 289
rect 1266 221 1324 255
rect 1266 187 1278 221
rect 1312 187 1324 221
tri 1354 278 1370 294 se
rect 1370 278 1414 294
tri 1414 278 1430 294 sw
rect 1354 245 1430 278
rect 1354 211 1375 245
rect 1409 211 1430 245
rect 1354 209 1430 211
tri 1354 193 1370 209 ne
rect 1370 193 1414 209
tri 1414 193 1430 209 nw
rect 1460 289 1516 324
rect 1460 255 1472 289
rect 1506 255 1516 289
rect 1460 221 1516 255
tri 1130 155 1160 185 sw
tri 1236 155 1266 185 se
rect 1266 163 1324 187
tri 1324 163 1354 193 sw
tri 1430 163 1460 193 se
rect 1460 187 1472 221
rect 1506 187 1516 221
rect 1460 163 1516 187
rect 1266 155 1516 163
rect 1074 151 1516 155
rect 1074 117 1084 151
rect 1118 117 1278 151
rect 1312 117 1375 151
rect 1409 117 1472 151
rect 1506 117 1516 151
rect 1074 101 1516 117
rect 1740 361 1796 377
rect 1740 327 1750 361
rect 1784 327 1796 361
rect 1740 289 1796 327
rect 1826 361 1990 377
rect 1826 332 1847 361
tri 1826 316 1842 332 ne
rect 1842 327 1847 332
rect 1881 327 1944 361
rect 1978 327 1990 361
rect 1842 316 1990 327
rect 2020 340 2182 377
tri 2020 324 2036 340 ne
rect 2036 324 2182 340
rect 1740 255 1750 289
rect 1784 255 1796 289
tri 1902 286 1932 316 ne
rect 1932 289 1990 316
tri 2096 294 2126 324 ne
rect 1740 221 1796 255
rect 1740 187 1750 221
rect 1784 187 1796 221
rect 1740 155 1796 187
tri 1826 270 1842 286 se
rect 1842 270 1886 286
tri 1886 270 1902 286 sw
rect 1826 236 1902 270
rect 1826 202 1847 236
rect 1881 202 1902 236
rect 1826 201 1902 202
tri 1826 185 1842 201 ne
rect 1842 185 1886 201
tri 1886 185 1902 201 nw
rect 1932 255 1944 289
rect 1978 255 1990 289
rect 1932 221 1990 255
rect 1932 187 1944 221
rect 1978 187 1990 221
tri 2020 278 2036 294 se
rect 2036 278 2080 294
tri 2080 278 2096 294 sw
rect 2020 245 2096 278
rect 2020 211 2041 245
rect 2075 211 2096 245
rect 2020 209 2096 211
tri 2020 193 2036 209 ne
rect 2036 193 2080 209
tri 2080 193 2096 209 nw
rect 2126 289 2182 324
rect 2126 255 2138 289
rect 2172 255 2182 289
rect 2126 221 2182 255
tri 1796 155 1826 185 sw
tri 1902 155 1932 185 se
rect 1932 163 1990 187
tri 1990 163 2020 193 sw
tri 2096 163 2126 193 se
rect 2126 187 2138 221
rect 2172 187 2182 221
rect 2126 163 2182 187
rect 1932 155 2182 163
rect 1740 151 2182 155
rect 1740 117 1750 151
rect 1784 117 1944 151
rect 1978 117 2041 151
rect 2075 117 2138 151
rect 2172 117 2182 151
rect 1740 101 2182 117
rect 2406 361 2462 377
rect 2406 327 2416 361
rect 2450 327 2462 361
rect 2406 289 2462 327
rect 2492 361 2656 377
rect 2492 332 2513 361
tri 2492 316 2508 332 ne
rect 2508 327 2513 332
rect 2547 327 2610 361
rect 2644 327 2656 361
rect 2508 316 2656 327
rect 2686 340 2848 377
tri 2686 324 2702 340 ne
rect 2702 324 2848 340
rect 2406 255 2416 289
rect 2450 255 2462 289
tri 2568 286 2598 316 ne
rect 2598 289 2656 316
tri 2762 294 2792 324 ne
rect 2406 221 2462 255
rect 2406 187 2416 221
rect 2450 187 2462 221
rect 2406 155 2462 187
tri 2492 270 2508 286 se
rect 2508 270 2552 286
tri 2552 270 2568 286 sw
rect 2492 236 2568 270
rect 2492 202 2513 236
rect 2547 202 2568 236
rect 2492 201 2568 202
tri 2492 185 2508 201 ne
rect 2508 185 2552 201
tri 2552 185 2568 201 nw
rect 2598 255 2610 289
rect 2644 255 2656 289
rect 2598 221 2656 255
rect 2598 187 2610 221
rect 2644 187 2656 221
tri 2686 278 2702 294 se
rect 2702 278 2746 294
tri 2746 278 2762 294 sw
rect 2686 245 2762 278
rect 2686 211 2707 245
rect 2741 211 2762 245
rect 2686 209 2762 211
tri 2686 193 2702 209 ne
rect 2702 193 2746 209
tri 2746 193 2762 209 nw
rect 2792 289 2848 324
rect 2792 255 2804 289
rect 2838 255 2848 289
rect 2792 221 2848 255
tri 2462 155 2492 185 sw
tri 2568 155 2598 185 se
rect 2598 163 2656 187
tri 2656 163 2686 193 sw
tri 2762 163 2792 193 se
rect 2792 187 2804 221
rect 2838 187 2848 221
rect 2792 163 2848 187
rect 2598 155 2848 163
rect 2406 151 2848 155
rect 2406 117 2416 151
rect 2450 117 2610 151
rect 2644 117 2707 151
rect 2741 117 2804 151
rect 2838 117 2848 151
rect 2406 101 2848 117
rect 3072 361 3128 377
rect 3072 327 3082 361
rect 3116 327 3128 361
rect 3072 289 3128 327
rect 3158 361 3322 377
rect 3158 332 3179 361
tri 3158 316 3174 332 ne
rect 3174 327 3179 332
rect 3213 327 3276 361
rect 3310 327 3322 361
rect 3174 316 3322 327
rect 3352 340 3514 377
tri 3352 324 3368 340 ne
rect 3368 324 3514 340
rect 3072 255 3082 289
rect 3116 255 3128 289
tri 3234 286 3264 316 ne
rect 3264 289 3322 316
tri 3428 294 3458 324 ne
rect 3072 221 3128 255
rect 3072 187 3082 221
rect 3116 187 3128 221
rect 3072 155 3128 187
tri 3158 270 3174 286 se
rect 3174 270 3218 286
tri 3218 270 3234 286 sw
rect 3158 236 3234 270
rect 3158 202 3179 236
rect 3213 202 3234 236
rect 3158 201 3234 202
tri 3158 185 3174 201 ne
rect 3174 185 3218 201
tri 3218 185 3234 201 nw
rect 3264 255 3276 289
rect 3310 255 3322 289
rect 3264 221 3322 255
rect 3264 187 3276 221
rect 3310 187 3322 221
tri 3352 278 3368 294 se
rect 3368 278 3412 294
tri 3412 278 3428 294 sw
rect 3352 245 3428 278
rect 3352 211 3373 245
rect 3407 211 3428 245
rect 3352 209 3428 211
tri 3352 193 3368 209 ne
rect 3368 193 3412 209
tri 3412 193 3428 209 nw
rect 3458 289 3514 324
rect 3458 255 3470 289
rect 3504 255 3514 289
rect 3458 221 3514 255
tri 3128 155 3158 185 sw
tri 3234 155 3264 185 se
rect 3264 163 3322 187
tri 3322 163 3352 193 sw
tri 3428 163 3458 193 se
rect 3458 187 3470 221
rect 3504 187 3514 221
rect 3458 163 3514 187
rect 3264 155 3514 163
rect 3072 151 3514 155
rect 3072 117 3082 151
rect 3116 117 3276 151
rect 3310 117 3373 151
rect 3407 117 3470 151
rect 3504 117 3514 151
rect 3072 101 3514 117
rect 3738 361 3794 377
rect 3738 327 3748 361
rect 3782 327 3794 361
rect 3738 289 3794 327
rect 3824 361 3988 377
rect 3824 332 3845 361
tri 3824 316 3840 332 ne
rect 3840 327 3845 332
rect 3879 327 3942 361
rect 3976 327 3988 361
rect 3840 316 3988 327
rect 4018 340 4180 377
tri 4018 324 4034 340 ne
rect 4034 324 4180 340
rect 3738 255 3748 289
rect 3782 255 3794 289
tri 3900 286 3930 316 ne
rect 3930 289 3988 316
tri 4094 294 4124 324 ne
rect 3738 221 3794 255
rect 3738 187 3748 221
rect 3782 187 3794 221
rect 3738 155 3794 187
tri 3824 270 3840 286 se
rect 3840 270 3884 286
tri 3884 270 3900 286 sw
rect 3824 236 3900 270
rect 3824 202 3845 236
rect 3879 202 3900 236
rect 3824 201 3900 202
tri 3824 185 3840 201 ne
rect 3840 185 3884 201
tri 3884 185 3900 201 nw
rect 3930 255 3942 289
rect 3976 255 3988 289
rect 3930 221 3988 255
rect 3930 187 3942 221
rect 3976 187 3988 221
tri 4018 278 4034 294 se
rect 4034 278 4078 294
tri 4078 278 4094 294 sw
rect 4018 245 4094 278
rect 4018 211 4039 245
rect 4073 211 4094 245
rect 4018 209 4094 211
tri 4018 193 4034 209 ne
rect 4034 193 4078 209
tri 4078 193 4094 209 nw
rect 4124 289 4180 324
rect 4124 255 4136 289
rect 4170 255 4180 289
rect 4124 221 4180 255
tri 3794 155 3824 185 sw
tri 3900 155 3930 185 se
rect 3930 163 3988 187
tri 3988 163 4018 193 sw
tri 4094 163 4124 193 se
rect 4124 187 4136 221
rect 4170 187 4180 221
rect 4124 163 4180 187
rect 3930 155 4180 163
rect 3738 151 4180 155
rect 3738 117 3748 151
rect 3782 117 3942 151
rect 3976 117 4039 151
rect 4073 117 4136 151
rect 4170 117 4180 151
rect 3738 101 4180 117
<< pdiff >>
rect 191 1412 247 1450
rect 191 1378 201 1412
rect 235 1378 247 1412
rect 191 1344 247 1378
rect 191 1310 201 1344
rect 235 1310 247 1344
rect 191 1276 247 1310
rect 191 1242 201 1276
rect 235 1242 247 1276
rect 191 1208 247 1242
rect 191 1174 201 1208
rect 235 1174 247 1208
rect 191 1139 247 1174
rect 191 1105 201 1139
rect 235 1105 247 1139
rect 191 1050 247 1105
rect 277 1412 335 1450
rect 277 1378 289 1412
rect 323 1378 335 1412
rect 277 1344 335 1378
rect 277 1310 289 1344
rect 323 1310 335 1344
rect 277 1276 335 1310
rect 277 1242 289 1276
rect 323 1242 335 1276
rect 277 1208 335 1242
rect 277 1174 289 1208
rect 323 1174 335 1208
rect 277 1139 335 1174
rect 277 1105 289 1139
rect 323 1105 335 1139
rect 277 1050 335 1105
rect 365 1412 423 1450
rect 365 1378 377 1412
rect 411 1378 423 1412
rect 365 1344 423 1378
rect 365 1310 377 1344
rect 411 1310 423 1344
rect 365 1276 423 1310
rect 365 1242 377 1276
rect 411 1242 423 1276
rect 365 1208 423 1242
rect 365 1174 377 1208
rect 411 1174 423 1208
rect 365 1050 423 1174
rect 453 1412 511 1450
rect 453 1378 465 1412
rect 499 1378 511 1412
rect 453 1344 511 1378
rect 453 1310 465 1344
rect 499 1310 511 1344
rect 453 1276 511 1310
rect 453 1242 465 1276
rect 499 1242 511 1276
rect 453 1208 511 1242
rect 453 1174 465 1208
rect 499 1174 511 1208
rect 453 1139 511 1174
rect 453 1105 465 1139
rect 499 1105 511 1139
rect 453 1050 511 1105
rect 541 1412 599 1450
rect 541 1378 553 1412
rect 587 1378 599 1412
rect 541 1344 599 1378
rect 541 1310 553 1344
rect 587 1310 599 1344
rect 541 1276 599 1310
rect 541 1242 553 1276
rect 587 1242 599 1276
rect 541 1208 599 1242
rect 541 1174 553 1208
rect 587 1174 599 1208
rect 541 1050 599 1174
rect 629 1412 687 1450
rect 629 1378 641 1412
rect 675 1378 687 1412
rect 629 1344 687 1378
rect 629 1310 641 1344
rect 675 1310 687 1344
rect 629 1276 687 1310
rect 629 1242 641 1276
rect 675 1242 687 1276
rect 629 1208 687 1242
rect 629 1174 641 1208
rect 675 1174 687 1208
rect 629 1139 687 1174
rect 629 1105 641 1139
rect 675 1105 687 1139
rect 629 1050 687 1105
rect 717 1412 771 1450
rect 717 1378 729 1412
rect 763 1378 771 1412
rect 717 1344 771 1378
rect 717 1310 729 1344
rect 763 1310 771 1344
rect 717 1276 771 1310
rect 717 1242 729 1276
rect 763 1242 771 1276
rect 717 1208 771 1242
rect 717 1174 729 1208
rect 763 1174 771 1208
rect 717 1050 771 1174
rect 1093 1412 1149 1450
rect 1093 1378 1103 1412
rect 1137 1378 1149 1412
rect 1093 1344 1149 1378
rect 1093 1310 1103 1344
rect 1137 1310 1149 1344
rect 1093 1276 1149 1310
rect 1093 1242 1103 1276
rect 1137 1242 1149 1276
rect 1093 1208 1149 1242
rect 1093 1174 1103 1208
rect 1137 1174 1149 1208
rect 1093 1139 1149 1174
rect 1093 1105 1103 1139
rect 1137 1105 1149 1139
rect 1093 1050 1149 1105
rect 1179 1412 1237 1450
rect 1179 1378 1191 1412
rect 1225 1378 1237 1412
rect 1179 1344 1237 1378
rect 1179 1310 1191 1344
rect 1225 1310 1237 1344
rect 1179 1276 1237 1310
rect 1179 1242 1191 1276
rect 1225 1242 1237 1276
rect 1179 1208 1237 1242
rect 1179 1174 1191 1208
rect 1225 1174 1237 1208
rect 1179 1139 1237 1174
rect 1179 1105 1191 1139
rect 1225 1105 1237 1139
rect 1179 1050 1237 1105
rect 1267 1412 1325 1450
rect 1267 1378 1279 1412
rect 1313 1378 1325 1412
rect 1267 1344 1325 1378
rect 1267 1310 1279 1344
rect 1313 1310 1325 1344
rect 1267 1276 1325 1310
rect 1267 1242 1279 1276
rect 1313 1242 1325 1276
rect 1267 1208 1325 1242
rect 1267 1174 1279 1208
rect 1313 1174 1325 1208
rect 1267 1050 1325 1174
rect 1355 1412 1413 1450
rect 1355 1378 1367 1412
rect 1401 1378 1413 1412
rect 1355 1344 1413 1378
rect 1355 1310 1367 1344
rect 1401 1310 1413 1344
rect 1355 1276 1413 1310
rect 1355 1242 1367 1276
rect 1401 1242 1413 1276
rect 1355 1208 1413 1242
rect 1355 1174 1367 1208
rect 1401 1174 1413 1208
rect 1355 1139 1413 1174
rect 1355 1105 1367 1139
rect 1401 1105 1413 1139
rect 1355 1050 1413 1105
rect 1443 1412 1497 1450
rect 1443 1378 1455 1412
rect 1489 1378 1497 1412
rect 1443 1344 1497 1378
rect 1443 1310 1455 1344
rect 1489 1310 1497 1344
rect 1443 1276 1497 1310
rect 1443 1242 1455 1276
rect 1489 1242 1497 1276
rect 1443 1208 1497 1242
rect 1443 1174 1455 1208
rect 1489 1174 1497 1208
rect 1443 1050 1497 1174
rect 1759 1412 1815 1450
rect 1759 1378 1769 1412
rect 1803 1378 1815 1412
rect 1759 1344 1815 1378
rect 1759 1310 1769 1344
rect 1803 1310 1815 1344
rect 1759 1276 1815 1310
rect 1759 1242 1769 1276
rect 1803 1242 1815 1276
rect 1759 1208 1815 1242
rect 1759 1174 1769 1208
rect 1803 1174 1815 1208
rect 1759 1139 1815 1174
rect 1759 1105 1769 1139
rect 1803 1105 1815 1139
rect 1759 1050 1815 1105
rect 1845 1412 1903 1450
rect 1845 1378 1857 1412
rect 1891 1378 1903 1412
rect 1845 1344 1903 1378
rect 1845 1310 1857 1344
rect 1891 1310 1903 1344
rect 1845 1276 1903 1310
rect 1845 1242 1857 1276
rect 1891 1242 1903 1276
rect 1845 1208 1903 1242
rect 1845 1174 1857 1208
rect 1891 1174 1903 1208
rect 1845 1139 1903 1174
rect 1845 1105 1857 1139
rect 1891 1105 1903 1139
rect 1845 1050 1903 1105
rect 1933 1412 1991 1450
rect 1933 1378 1945 1412
rect 1979 1378 1991 1412
rect 1933 1344 1991 1378
rect 1933 1310 1945 1344
rect 1979 1310 1991 1344
rect 1933 1276 1991 1310
rect 1933 1242 1945 1276
rect 1979 1242 1991 1276
rect 1933 1208 1991 1242
rect 1933 1174 1945 1208
rect 1979 1174 1991 1208
rect 1933 1050 1991 1174
rect 2021 1412 2079 1450
rect 2021 1378 2033 1412
rect 2067 1378 2079 1412
rect 2021 1344 2079 1378
rect 2021 1310 2033 1344
rect 2067 1310 2079 1344
rect 2021 1276 2079 1310
rect 2021 1242 2033 1276
rect 2067 1242 2079 1276
rect 2021 1208 2079 1242
rect 2021 1174 2033 1208
rect 2067 1174 2079 1208
rect 2021 1139 2079 1174
rect 2021 1105 2033 1139
rect 2067 1105 2079 1139
rect 2021 1050 2079 1105
rect 2109 1412 2163 1450
rect 2109 1378 2121 1412
rect 2155 1378 2163 1412
rect 2109 1344 2163 1378
rect 2109 1310 2121 1344
rect 2155 1310 2163 1344
rect 2109 1276 2163 1310
rect 2109 1242 2121 1276
rect 2155 1242 2163 1276
rect 2109 1208 2163 1242
rect 2109 1174 2121 1208
rect 2155 1174 2163 1208
rect 2109 1050 2163 1174
rect 2425 1412 2481 1450
rect 2425 1378 2435 1412
rect 2469 1378 2481 1412
rect 2425 1344 2481 1378
rect 2425 1310 2435 1344
rect 2469 1310 2481 1344
rect 2425 1276 2481 1310
rect 2425 1242 2435 1276
rect 2469 1242 2481 1276
rect 2425 1208 2481 1242
rect 2425 1174 2435 1208
rect 2469 1174 2481 1208
rect 2425 1139 2481 1174
rect 2425 1105 2435 1139
rect 2469 1105 2481 1139
rect 2425 1050 2481 1105
rect 2511 1412 2569 1450
rect 2511 1378 2523 1412
rect 2557 1378 2569 1412
rect 2511 1344 2569 1378
rect 2511 1310 2523 1344
rect 2557 1310 2569 1344
rect 2511 1276 2569 1310
rect 2511 1242 2523 1276
rect 2557 1242 2569 1276
rect 2511 1208 2569 1242
rect 2511 1174 2523 1208
rect 2557 1174 2569 1208
rect 2511 1139 2569 1174
rect 2511 1105 2523 1139
rect 2557 1105 2569 1139
rect 2511 1050 2569 1105
rect 2599 1412 2657 1450
rect 2599 1378 2611 1412
rect 2645 1378 2657 1412
rect 2599 1344 2657 1378
rect 2599 1310 2611 1344
rect 2645 1310 2657 1344
rect 2599 1276 2657 1310
rect 2599 1242 2611 1276
rect 2645 1242 2657 1276
rect 2599 1208 2657 1242
rect 2599 1174 2611 1208
rect 2645 1174 2657 1208
rect 2599 1050 2657 1174
rect 2687 1412 2745 1450
rect 2687 1378 2699 1412
rect 2733 1378 2745 1412
rect 2687 1344 2745 1378
rect 2687 1310 2699 1344
rect 2733 1310 2745 1344
rect 2687 1276 2745 1310
rect 2687 1242 2699 1276
rect 2733 1242 2745 1276
rect 2687 1208 2745 1242
rect 2687 1174 2699 1208
rect 2733 1174 2745 1208
rect 2687 1139 2745 1174
rect 2687 1105 2699 1139
rect 2733 1105 2745 1139
rect 2687 1050 2745 1105
rect 2775 1412 2829 1450
rect 2775 1378 2787 1412
rect 2821 1378 2829 1412
rect 2775 1344 2829 1378
rect 2775 1310 2787 1344
rect 2821 1310 2829 1344
rect 2775 1276 2829 1310
rect 2775 1242 2787 1276
rect 2821 1242 2829 1276
rect 2775 1208 2829 1242
rect 2775 1174 2787 1208
rect 2821 1174 2829 1208
rect 2775 1050 2829 1174
rect 3091 1412 3147 1450
rect 3091 1378 3101 1412
rect 3135 1378 3147 1412
rect 3091 1344 3147 1378
rect 3091 1310 3101 1344
rect 3135 1310 3147 1344
rect 3091 1276 3147 1310
rect 3091 1242 3101 1276
rect 3135 1242 3147 1276
rect 3091 1208 3147 1242
rect 3091 1174 3101 1208
rect 3135 1174 3147 1208
rect 3091 1139 3147 1174
rect 3091 1105 3101 1139
rect 3135 1105 3147 1139
rect 3091 1050 3147 1105
rect 3177 1412 3235 1450
rect 3177 1378 3189 1412
rect 3223 1378 3235 1412
rect 3177 1344 3235 1378
rect 3177 1310 3189 1344
rect 3223 1310 3235 1344
rect 3177 1276 3235 1310
rect 3177 1242 3189 1276
rect 3223 1242 3235 1276
rect 3177 1208 3235 1242
rect 3177 1174 3189 1208
rect 3223 1174 3235 1208
rect 3177 1139 3235 1174
rect 3177 1105 3189 1139
rect 3223 1105 3235 1139
rect 3177 1050 3235 1105
rect 3265 1412 3323 1450
rect 3265 1378 3277 1412
rect 3311 1378 3323 1412
rect 3265 1344 3323 1378
rect 3265 1310 3277 1344
rect 3311 1310 3323 1344
rect 3265 1276 3323 1310
rect 3265 1242 3277 1276
rect 3311 1242 3323 1276
rect 3265 1208 3323 1242
rect 3265 1174 3277 1208
rect 3311 1174 3323 1208
rect 3265 1050 3323 1174
rect 3353 1412 3411 1450
rect 3353 1378 3365 1412
rect 3399 1378 3411 1412
rect 3353 1344 3411 1378
rect 3353 1310 3365 1344
rect 3399 1310 3411 1344
rect 3353 1276 3411 1310
rect 3353 1242 3365 1276
rect 3399 1242 3411 1276
rect 3353 1208 3411 1242
rect 3353 1174 3365 1208
rect 3399 1174 3411 1208
rect 3353 1139 3411 1174
rect 3353 1105 3365 1139
rect 3399 1105 3411 1139
rect 3353 1050 3411 1105
rect 3441 1412 3495 1450
rect 3441 1378 3453 1412
rect 3487 1378 3495 1412
rect 3441 1344 3495 1378
rect 3441 1310 3453 1344
rect 3487 1310 3495 1344
rect 3441 1276 3495 1310
rect 3441 1242 3453 1276
rect 3487 1242 3495 1276
rect 3441 1208 3495 1242
rect 3441 1174 3453 1208
rect 3487 1174 3495 1208
rect 3441 1050 3495 1174
rect 3757 1412 3813 1450
rect 3757 1378 3767 1412
rect 3801 1378 3813 1412
rect 3757 1344 3813 1378
rect 3757 1310 3767 1344
rect 3801 1310 3813 1344
rect 3757 1276 3813 1310
rect 3757 1242 3767 1276
rect 3801 1242 3813 1276
rect 3757 1208 3813 1242
rect 3757 1174 3767 1208
rect 3801 1174 3813 1208
rect 3757 1139 3813 1174
rect 3757 1105 3767 1139
rect 3801 1105 3813 1139
rect 3757 1050 3813 1105
rect 3843 1412 3901 1450
rect 3843 1378 3855 1412
rect 3889 1378 3901 1412
rect 3843 1344 3901 1378
rect 3843 1310 3855 1344
rect 3889 1310 3901 1344
rect 3843 1276 3901 1310
rect 3843 1242 3855 1276
rect 3889 1242 3901 1276
rect 3843 1208 3901 1242
rect 3843 1174 3855 1208
rect 3889 1174 3901 1208
rect 3843 1139 3901 1174
rect 3843 1105 3855 1139
rect 3889 1105 3901 1139
rect 3843 1050 3901 1105
rect 3931 1412 3989 1450
rect 3931 1378 3943 1412
rect 3977 1378 3989 1412
rect 3931 1344 3989 1378
rect 3931 1310 3943 1344
rect 3977 1310 3989 1344
rect 3931 1276 3989 1310
rect 3931 1242 3943 1276
rect 3977 1242 3989 1276
rect 3931 1208 3989 1242
rect 3931 1174 3943 1208
rect 3977 1174 3989 1208
rect 3931 1050 3989 1174
rect 4019 1412 4077 1450
rect 4019 1378 4031 1412
rect 4065 1378 4077 1412
rect 4019 1344 4077 1378
rect 4019 1310 4031 1344
rect 4065 1310 4077 1344
rect 4019 1276 4077 1310
rect 4019 1242 4031 1276
rect 4065 1242 4077 1276
rect 4019 1208 4077 1242
rect 4019 1174 4031 1208
rect 4065 1174 4077 1208
rect 4019 1139 4077 1174
rect 4019 1105 4031 1139
rect 4065 1105 4077 1139
rect 4019 1050 4077 1105
rect 4107 1412 4161 1450
rect 4107 1378 4119 1412
rect 4153 1378 4161 1412
rect 4107 1344 4161 1378
rect 4107 1310 4119 1344
rect 4153 1310 4161 1344
rect 4107 1276 4161 1310
rect 4107 1242 4119 1276
rect 4153 1242 4161 1276
rect 4107 1208 4161 1242
rect 4107 1174 4119 1208
rect 4153 1174 4161 1208
rect 4107 1050 4161 1174
<< ndiffc >>
rect 101 329 135 363
rect 198 329 232 363
rect 295 329 329 363
rect 392 329 426 363
rect 489 329 523 363
rect 101 257 135 291
rect 101 189 135 223
rect 198 204 232 238
rect 295 257 329 291
rect 295 189 329 223
rect 393 210 427 244
rect 101 119 135 153
rect 295 119 329 153
rect 392 119 426 153
rect 489 119 523 153
rect 603 329 637 363
rect 603 257 637 291
rect 603 189 637 223
rect 700 213 734 247
rect 797 257 831 291
rect 797 189 831 223
rect 603 119 637 153
rect 700 119 734 153
rect 797 119 831 153
rect 1084 327 1118 361
rect 1181 327 1215 361
rect 1278 327 1312 361
rect 1084 255 1118 289
rect 1084 187 1118 221
rect 1181 202 1215 236
rect 1278 255 1312 289
rect 1278 187 1312 221
rect 1375 211 1409 245
rect 1472 255 1506 289
rect 1472 187 1506 221
rect 1084 117 1118 151
rect 1278 117 1312 151
rect 1375 117 1409 151
rect 1472 117 1506 151
rect 1750 327 1784 361
rect 1847 327 1881 361
rect 1944 327 1978 361
rect 1750 255 1784 289
rect 1750 187 1784 221
rect 1847 202 1881 236
rect 1944 255 1978 289
rect 1944 187 1978 221
rect 2041 211 2075 245
rect 2138 255 2172 289
rect 2138 187 2172 221
rect 1750 117 1784 151
rect 1944 117 1978 151
rect 2041 117 2075 151
rect 2138 117 2172 151
rect 2416 327 2450 361
rect 2513 327 2547 361
rect 2610 327 2644 361
rect 2416 255 2450 289
rect 2416 187 2450 221
rect 2513 202 2547 236
rect 2610 255 2644 289
rect 2610 187 2644 221
rect 2707 211 2741 245
rect 2804 255 2838 289
rect 2804 187 2838 221
rect 2416 117 2450 151
rect 2610 117 2644 151
rect 2707 117 2741 151
rect 2804 117 2838 151
rect 3082 327 3116 361
rect 3179 327 3213 361
rect 3276 327 3310 361
rect 3082 255 3116 289
rect 3082 187 3116 221
rect 3179 202 3213 236
rect 3276 255 3310 289
rect 3276 187 3310 221
rect 3373 211 3407 245
rect 3470 255 3504 289
rect 3470 187 3504 221
rect 3082 117 3116 151
rect 3276 117 3310 151
rect 3373 117 3407 151
rect 3470 117 3504 151
rect 3748 327 3782 361
rect 3845 327 3879 361
rect 3942 327 3976 361
rect 3748 255 3782 289
rect 3748 187 3782 221
rect 3845 202 3879 236
rect 3942 255 3976 289
rect 3942 187 3976 221
rect 4039 211 4073 245
rect 4136 255 4170 289
rect 4136 187 4170 221
rect 3748 117 3782 151
rect 3942 117 3976 151
rect 4039 117 4073 151
rect 4136 117 4170 151
<< pdiffc >>
rect 201 1378 235 1412
rect 201 1310 235 1344
rect 201 1242 235 1276
rect 201 1174 235 1208
rect 201 1105 235 1139
rect 289 1378 323 1412
rect 289 1310 323 1344
rect 289 1242 323 1276
rect 289 1174 323 1208
rect 289 1105 323 1139
rect 377 1378 411 1412
rect 377 1310 411 1344
rect 377 1242 411 1276
rect 377 1174 411 1208
rect 465 1378 499 1412
rect 465 1310 499 1344
rect 465 1242 499 1276
rect 465 1174 499 1208
rect 465 1105 499 1139
rect 553 1378 587 1412
rect 553 1310 587 1344
rect 553 1242 587 1276
rect 553 1174 587 1208
rect 641 1378 675 1412
rect 641 1310 675 1344
rect 641 1242 675 1276
rect 641 1174 675 1208
rect 641 1105 675 1139
rect 729 1378 763 1412
rect 729 1310 763 1344
rect 729 1242 763 1276
rect 729 1174 763 1208
rect 1103 1378 1137 1412
rect 1103 1310 1137 1344
rect 1103 1242 1137 1276
rect 1103 1174 1137 1208
rect 1103 1105 1137 1139
rect 1191 1378 1225 1412
rect 1191 1310 1225 1344
rect 1191 1242 1225 1276
rect 1191 1174 1225 1208
rect 1191 1105 1225 1139
rect 1279 1378 1313 1412
rect 1279 1310 1313 1344
rect 1279 1242 1313 1276
rect 1279 1174 1313 1208
rect 1367 1378 1401 1412
rect 1367 1310 1401 1344
rect 1367 1242 1401 1276
rect 1367 1174 1401 1208
rect 1367 1105 1401 1139
rect 1455 1378 1489 1412
rect 1455 1310 1489 1344
rect 1455 1242 1489 1276
rect 1455 1174 1489 1208
rect 1769 1378 1803 1412
rect 1769 1310 1803 1344
rect 1769 1242 1803 1276
rect 1769 1174 1803 1208
rect 1769 1105 1803 1139
rect 1857 1378 1891 1412
rect 1857 1310 1891 1344
rect 1857 1242 1891 1276
rect 1857 1174 1891 1208
rect 1857 1105 1891 1139
rect 1945 1378 1979 1412
rect 1945 1310 1979 1344
rect 1945 1242 1979 1276
rect 1945 1174 1979 1208
rect 2033 1378 2067 1412
rect 2033 1310 2067 1344
rect 2033 1242 2067 1276
rect 2033 1174 2067 1208
rect 2033 1105 2067 1139
rect 2121 1378 2155 1412
rect 2121 1310 2155 1344
rect 2121 1242 2155 1276
rect 2121 1174 2155 1208
rect 2435 1378 2469 1412
rect 2435 1310 2469 1344
rect 2435 1242 2469 1276
rect 2435 1174 2469 1208
rect 2435 1105 2469 1139
rect 2523 1378 2557 1412
rect 2523 1310 2557 1344
rect 2523 1242 2557 1276
rect 2523 1174 2557 1208
rect 2523 1105 2557 1139
rect 2611 1378 2645 1412
rect 2611 1310 2645 1344
rect 2611 1242 2645 1276
rect 2611 1174 2645 1208
rect 2699 1378 2733 1412
rect 2699 1310 2733 1344
rect 2699 1242 2733 1276
rect 2699 1174 2733 1208
rect 2699 1105 2733 1139
rect 2787 1378 2821 1412
rect 2787 1310 2821 1344
rect 2787 1242 2821 1276
rect 2787 1174 2821 1208
rect 3101 1378 3135 1412
rect 3101 1310 3135 1344
rect 3101 1242 3135 1276
rect 3101 1174 3135 1208
rect 3101 1105 3135 1139
rect 3189 1378 3223 1412
rect 3189 1310 3223 1344
rect 3189 1242 3223 1276
rect 3189 1174 3223 1208
rect 3189 1105 3223 1139
rect 3277 1378 3311 1412
rect 3277 1310 3311 1344
rect 3277 1242 3311 1276
rect 3277 1174 3311 1208
rect 3365 1378 3399 1412
rect 3365 1310 3399 1344
rect 3365 1242 3399 1276
rect 3365 1174 3399 1208
rect 3365 1105 3399 1139
rect 3453 1378 3487 1412
rect 3453 1310 3487 1344
rect 3453 1242 3487 1276
rect 3453 1174 3487 1208
rect 3767 1378 3801 1412
rect 3767 1310 3801 1344
rect 3767 1242 3801 1276
rect 3767 1174 3801 1208
rect 3767 1105 3801 1139
rect 3855 1378 3889 1412
rect 3855 1310 3889 1344
rect 3855 1242 3889 1276
rect 3855 1174 3889 1208
rect 3855 1105 3889 1139
rect 3943 1378 3977 1412
rect 3943 1310 3977 1344
rect 3943 1242 3977 1276
rect 3943 1174 3977 1208
rect 4031 1378 4065 1412
rect 4031 1310 4065 1344
rect 4031 1242 4065 1276
rect 4031 1174 4065 1208
rect 4031 1105 4065 1139
rect 4119 1378 4153 1412
rect 4119 1310 4153 1344
rect 4119 1242 4153 1276
rect 4119 1174 4153 1208
<< psubdiff >>
rect -31 546 4323 572
rect -31 512 -17 546
rect 17 512 945 546
rect 979 512 1611 546
rect 1645 512 2277 546
rect 2311 512 2943 546
rect 2977 512 3609 546
rect 3643 512 4275 546
rect 4309 512 4323 546
rect -31 510 4323 512
rect -31 474 31 510
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect -31 368 -17 402
rect 17 368 31 402
rect 931 474 993 510
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 931 368 945 402
rect 979 368 993 402
rect 1597 474 1659 510
rect 1597 440 1611 474
rect 1645 440 1659 474
rect 1597 402 1659 440
rect 931 330 993 368
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect -31 47 31 80
rect 931 80 945 114
rect 979 80 993 114
rect 1597 368 1611 402
rect 1645 368 1659 402
rect 2263 474 2325 510
rect 2263 440 2277 474
rect 2311 440 2325 474
rect 2263 402 2325 440
rect 1597 330 1659 368
rect 1597 296 1611 330
rect 1645 296 1659 330
rect 1597 258 1659 296
rect 1597 224 1611 258
rect 1645 224 1659 258
rect 1597 186 1659 224
rect 1597 152 1611 186
rect 1645 152 1659 186
rect 1597 114 1659 152
rect 931 47 993 80
rect 1597 80 1611 114
rect 1645 80 1659 114
rect 2263 368 2277 402
rect 2311 368 2325 402
rect 2929 474 2991 510
rect 2929 440 2943 474
rect 2977 440 2991 474
rect 2929 402 2991 440
rect 2263 330 2325 368
rect 2263 296 2277 330
rect 2311 296 2325 330
rect 2263 258 2325 296
rect 2263 224 2277 258
rect 2311 224 2325 258
rect 2263 186 2325 224
rect 2263 152 2277 186
rect 2311 152 2325 186
rect 2263 114 2325 152
rect 1597 47 1659 80
rect 2263 80 2277 114
rect 2311 80 2325 114
rect 2929 368 2943 402
rect 2977 368 2991 402
rect 3595 474 3657 510
rect 3595 440 3609 474
rect 3643 440 3657 474
rect 3595 402 3657 440
rect 2929 330 2991 368
rect 2929 296 2943 330
rect 2977 296 2991 330
rect 2929 258 2991 296
rect 2929 224 2943 258
rect 2977 224 2991 258
rect 2929 186 2991 224
rect 2929 152 2943 186
rect 2977 152 2991 186
rect 2929 114 2991 152
rect 2263 47 2325 80
rect 2929 80 2943 114
rect 2977 80 2991 114
rect 3595 368 3609 402
rect 3643 368 3657 402
rect 4261 474 4323 510
rect 4261 440 4275 474
rect 4309 440 4323 474
rect 4261 402 4323 440
rect 3595 330 3657 368
rect 3595 296 3609 330
rect 3643 296 3657 330
rect 3595 258 3657 296
rect 3595 224 3609 258
rect 3643 224 3657 258
rect 3595 186 3657 224
rect 3595 152 3609 186
rect 3643 152 3657 186
rect 3595 114 3657 152
rect 2929 47 2991 80
rect 3595 80 3609 114
rect 3643 80 3657 114
rect 4261 368 4275 402
rect 4309 368 4323 402
rect 4261 330 4323 368
rect 4261 296 4275 330
rect 4309 296 4323 330
rect 4261 258 4323 296
rect 4261 224 4275 258
rect 4309 224 4323 258
rect 4261 186 4323 224
rect 4261 152 4275 186
rect 4309 152 4323 186
rect 4261 114 4323 152
rect 3595 47 3657 80
rect 4261 80 4275 114
rect 4309 80 4323 114
rect 4261 47 4323 80
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1323 47
rect 1357 13 1395 47
rect 1429 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1683 47
rect 1717 13 1755 47
rect 1789 13 1827 47
rect 1861 13 1899 47
rect 1933 13 1989 47
rect 2023 13 2061 47
rect 2095 13 2133 47
rect 2167 13 2205 47
rect 2239 13 2349 47
rect 2383 13 2421 47
rect 2455 13 2493 47
rect 2527 13 2565 47
rect 2599 13 2655 47
rect 2689 13 2727 47
rect 2761 13 2799 47
rect 2833 13 2871 47
rect 2905 13 3015 47
rect 3049 13 3087 47
rect 3121 13 3159 47
rect 3193 13 3231 47
rect 3265 13 3321 47
rect 3355 13 3393 47
rect 3427 13 3465 47
rect 3499 13 3537 47
rect 3571 13 3681 47
rect 3715 13 3753 47
rect 3787 13 3825 47
rect 3859 13 3897 47
rect 3931 13 3987 47
rect 4021 13 4059 47
rect 4093 13 4131 47
rect 4165 13 4203 47
rect 4237 13 4323 47
rect -31 11 31 13
rect 931 11 993 13
rect 1597 11 1659 13
rect 2263 11 2325 13
rect 2929 11 2991 13
rect 3595 11 3657 13
rect 4261 11 4323 13
<< nsubdiff >>
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1323 1539
rect 1357 1505 1395 1539
rect 1429 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1683 1539
rect 1717 1505 1755 1539
rect 1789 1505 1827 1539
rect 1861 1505 1899 1539
rect 1933 1505 1989 1539
rect 2023 1505 2061 1539
rect 2095 1505 2133 1539
rect 2167 1505 2205 1539
rect 2239 1505 2349 1539
rect 2383 1505 2421 1539
rect 2455 1505 2493 1539
rect 2527 1505 2565 1539
rect 2599 1505 2655 1539
rect 2689 1505 2727 1539
rect 2761 1505 2799 1539
rect 2833 1505 2871 1539
rect 2905 1505 3015 1539
rect 3049 1505 3087 1539
rect 3121 1505 3159 1539
rect 3193 1505 3231 1539
rect 3265 1505 3321 1539
rect 3355 1505 3393 1539
rect 3427 1505 3465 1539
rect 3499 1505 3537 1539
rect 3571 1505 3681 1539
rect 3715 1505 3753 1539
rect 3787 1505 3825 1539
rect 3859 1505 3897 1539
rect 3931 1505 3987 1539
rect 4021 1505 4059 1539
rect 4093 1505 4131 1539
rect 4165 1505 4203 1539
rect 4237 1505 4323 1539
rect -31 1470 31 1505
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect 931 1470 993 1505
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect -31 1038 31 1076
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 1597 1470 1659 1505
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect 931 1076 945 1110
rect 979 1076 993 1110
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect 931 1038 993 1076
rect 1597 1436 1611 1470
rect 1645 1436 1659 1470
rect 2263 1470 2325 1505
rect 1597 1398 1659 1436
rect 1597 1364 1611 1398
rect 1645 1364 1659 1398
rect 1597 1326 1659 1364
rect 1597 1292 1611 1326
rect 1645 1292 1659 1326
rect 1597 1254 1659 1292
rect 1597 1220 1611 1254
rect 1645 1220 1659 1254
rect 1597 1182 1659 1220
rect 1597 1148 1611 1182
rect 1645 1148 1659 1182
rect 1597 1110 1659 1148
rect 1597 1076 1611 1110
rect 1645 1076 1659 1110
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect -31 930 31 932
rect 931 932 945 966
rect 979 932 993 966
rect 1597 1038 1659 1076
rect 2263 1436 2277 1470
rect 2311 1436 2325 1470
rect 2929 1470 2991 1505
rect 2263 1398 2325 1436
rect 2263 1364 2277 1398
rect 2311 1364 2325 1398
rect 2263 1326 2325 1364
rect 2263 1292 2277 1326
rect 2311 1292 2325 1326
rect 2263 1254 2325 1292
rect 2263 1220 2277 1254
rect 2311 1220 2325 1254
rect 2263 1182 2325 1220
rect 2263 1148 2277 1182
rect 2311 1148 2325 1182
rect 2263 1110 2325 1148
rect 2263 1076 2277 1110
rect 2311 1076 2325 1110
rect 1597 1004 1611 1038
rect 1645 1004 1659 1038
rect 1597 966 1659 1004
rect 931 930 993 932
rect 1597 932 1611 966
rect 1645 932 1659 966
rect 2263 1038 2325 1076
rect 2929 1436 2943 1470
rect 2977 1436 2991 1470
rect 3595 1470 3657 1505
rect 2929 1398 2991 1436
rect 2929 1364 2943 1398
rect 2977 1364 2991 1398
rect 2929 1326 2991 1364
rect 2929 1292 2943 1326
rect 2977 1292 2991 1326
rect 2929 1254 2991 1292
rect 2929 1220 2943 1254
rect 2977 1220 2991 1254
rect 2929 1182 2991 1220
rect 2929 1148 2943 1182
rect 2977 1148 2991 1182
rect 2929 1110 2991 1148
rect 2929 1076 2943 1110
rect 2977 1076 2991 1110
rect 2263 1004 2277 1038
rect 2311 1004 2325 1038
rect 2263 966 2325 1004
rect 1597 930 1659 932
rect 2263 932 2277 966
rect 2311 932 2325 966
rect 2929 1038 2991 1076
rect 3595 1436 3609 1470
rect 3643 1436 3657 1470
rect 4261 1470 4323 1505
rect 3595 1398 3657 1436
rect 3595 1364 3609 1398
rect 3643 1364 3657 1398
rect 3595 1326 3657 1364
rect 3595 1292 3609 1326
rect 3643 1292 3657 1326
rect 3595 1254 3657 1292
rect 3595 1220 3609 1254
rect 3643 1220 3657 1254
rect 3595 1182 3657 1220
rect 3595 1148 3609 1182
rect 3643 1148 3657 1182
rect 3595 1110 3657 1148
rect 3595 1076 3609 1110
rect 3643 1076 3657 1110
rect 2929 1004 2943 1038
rect 2977 1004 2991 1038
rect 2929 966 2991 1004
rect 2263 930 2325 932
rect 2929 932 2943 966
rect 2977 932 2991 966
rect 3595 1038 3657 1076
rect 4261 1436 4275 1470
rect 4309 1436 4323 1470
rect 4261 1398 4323 1436
rect 4261 1364 4275 1398
rect 4309 1364 4323 1398
rect 4261 1326 4323 1364
rect 4261 1292 4275 1326
rect 4309 1292 4323 1326
rect 4261 1254 4323 1292
rect 4261 1220 4275 1254
rect 4309 1220 4323 1254
rect 4261 1182 4323 1220
rect 4261 1148 4275 1182
rect 4309 1148 4323 1182
rect 4261 1110 4323 1148
rect 4261 1076 4275 1110
rect 4309 1076 4323 1110
rect 3595 1004 3609 1038
rect 3643 1004 3657 1038
rect 3595 966 3657 1004
rect 2929 930 2991 932
rect 3595 932 3609 966
rect 3643 932 3657 966
rect 4261 1038 4323 1076
rect 4261 1004 4275 1038
rect 4309 1004 4323 1038
rect 4261 966 4323 1004
rect 3595 930 3657 932
rect 4261 932 4275 966
rect 4309 932 4323 966
rect 4261 930 4323 932
rect -31 868 4323 930
<< psubdiffcont >>
rect -17 512 17 546
rect 945 512 979 546
rect 1611 512 1645 546
rect 2277 512 2311 546
rect 2943 512 2977 546
rect 3609 512 3643 546
rect 4275 512 4309 546
rect -17 440 17 474
rect -17 368 17 402
rect 945 440 979 474
rect -17 296 17 330
rect -17 224 17 258
rect -17 152 17 186
rect -17 80 17 114
rect 945 368 979 402
rect 1611 440 1645 474
rect 945 296 979 330
rect 945 224 979 258
rect 945 152 979 186
rect 945 80 979 114
rect 1611 368 1645 402
rect 2277 440 2311 474
rect 1611 296 1645 330
rect 1611 224 1645 258
rect 1611 152 1645 186
rect 1611 80 1645 114
rect 2277 368 2311 402
rect 2943 440 2977 474
rect 2277 296 2311 330
rect 2277 224 2311 258
rect 2277 152 2311 186
rect 2277 80 2311 114
rect 2943 368 2977 402
rect 3609 440 3643 474
rect 2943 296 2977 330
rect 2943 224 2977 258
rect 2943 152 2977 186
rect 2943 80 2977 114
rect 3609 368 3643 402
rect 4275 440 4309 474
rect 3609 296 3643 330
rect 3609 224 3643 258
rect 3609 152 3643 186
rect 3609 80 3643 114
rect 4275 368 4309 402
rect 4275 296 4309 330
rect 4275 224 4309 258
rect 4275 152 4309 186
rect 4275 80 4309 114
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1161 13 1195 47
rect 1233 13 1267 47
rect 1323 13 1357 47
rect 1395 13 1429 47
rect 1467 13 1501 47
rect 1539 13 1573 47
rect 1683 13 1717 47
rect 1755 13 1789 47
rect 1827 13 1861 47
rect 1899 13 1933 47
rect 1989 13 2023 47
rect 2061 13 2095 47
rect 2133 13 2167 47
rect 2205 13 2239 47
rect 2349 13 2383 47
rect 2421 13 2455 47
rect 2493 13 2527 47
rect 2565 13 2599 47
rect 2655 13 2689 47
rect 2727 13 2761 47
rect 2799 13 2833 47
rect 2871 13 2905 47
rect 3015 13 3049 47
rect 3087 13 3121 47
rect 3159 13 3193 47
rect 3231 13 3265 47
rect 3321 13 3355 47
rect 3393 13 3427 47
rect 3465 13 3499 47
rect 3537 13 3571 47
rect 3681 13 3715 47
rect 3753 13 3787 47
rect 3825 13 3859 47
rect 3897 13 3931 47
rect 3987 13 4021 47
rect 4059 13 4093 47
rect 4131 13 4165 47
rect 4203 13 4237 47
<< nsubdiffcont >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1161 1505 1195 1539
rect 1233 1505 1267 1539
rect 1323 1505 1357 1539
rect 1395 1505 1429 1539
rect 1467 1505 1501 1539
rect 1539 1505 1573 1539
rect 1683 1505 1717 1539
rect 1755 1505 1789 1539
rect 1827 1505 1861 1539
rect 1899 1505 1933 1539
rect 1989 1505 2023 1539
rect 2061 1505 2095 1539
rect 2133 1505 2167 1539
rect 2205 1505 2239 1539
rect 2349 1505 2383 1539
rect 2421 1505 2455 1539
rect 2493 1505 2527 1539
rect 2565 1505 2599 1539
rect 2655 1505 2689 1539
rect 2727 1505 2761 1539
rect 2799 1505 2833 1539
rect 2871 1505 2905 1539
rect 3015 1505 3049 1539
rect 3087 1505 3121 1539
rect 3159 1505 3193 1539
rect 3231 1505 3265 1539
rect 3321 1505 3355 1539
rect 3393 1505 3427 1539
rect 3465 1505 3499 1539
rect 3537 1505 3571 1539
rect 3681 1505 3715 1539
rect 3753 1505 3787 1539
rect 3825 1505 3859 1539
rect 3897 1505 3931 1539
rect 3987 1505 4021 1539
rect 4059 1505 4093 1539
rect 4131 1505 4165 1539
rect 4203 1505 4237 1539
rect -17 1436 17 1470
rect -17 1364 17 1398
rect -17 1292 17 1326
rect -17 1220 17 1254
rect -17 1148 17 1182
rect -17 1076 17 1110
rect 945 1436 979 1470
rect 945 1364 979 1398
rect 945 1292 979 1326
rect 945 1220 979 1254
rect 945 1148 979 1182
rect 945 1076 979 1110
rect -17 1004 17 1038
rect -17 932 17 966
rect 1611 1436 1645 1470
rect 1611 1364 1645 1398
rect 1611 1292 1645 1326
rect 1611 1220 1645 1254
rect 1611 1148 1645 1182
rect 1611 1076 1645 1110
rect 945 1004 979 1038
rect 945 932 979 966
rect 2277 1436 2311 1470
rect 2277 1364 2311 1398
rect 2277 1292 2311 1326
rect 2277 1220 2311 1254
rect 2277 1148 2311 1182
rect 2277 1076 2311 1110
rect 1611 1004 1645 1038
rect 1611 932 1645 966
rect 2943 1436 2977 1470
rect 2943 1364 2977 1398
rect 2943 1292 2977 1326
rect 2943 1220 2977 1254
rect 2943 1148 2977 1182
rect 2943 1076 2977 1110
rect 2277 1004 2311 1038
rect 2277 932 2311 966
rect 3609 1436 3643 1470
rect 3609 1364 3643 1398
rect 3609 1292 3643 1326
rect 3609 1220 3643 1254
rect 3609 1148 3643 1182
rect 3609 1076 3643 1110
rect 2943 1004 2977 1038
rect 2943 932 2977 966
rect 4275 1436 4309 1470
rect 4275 1364 4309 1398
rect 4275 1292 4309 1326
rect 4275 1220 4309 1254
rect 4275 1148 4309 1182
rect 4275 1076 4309 1110
rect 3609 1004 3643 1038
rect 3609 932 3643 966
rect 4275 1004 4309 1038
rect 4275 932 4309 966
<< poly >>
rect 247 1450 277 1476
rect 335 1450 365 1476
rect 423 1450 453 1476
rect 511 1450 541 1476
rect 599 1450 629 1476
rect 687 1450 717 1476
rect 1149 1450 1179 1476
rect 1237 1450 1267 1476
rect 1325 1450 1355 1476
rect 1413 1450 1443 1476
rect 247 1019 277 1050
rect 335 1019 365 1050
rect 423 1019 453 1050
rect 511 1019 541 1050
rect 195 1003 365 1019
rect 195 969 205 1003
rect 239 989 365 1003
rect 417 1003 541 1019
rect 239 969 249 989
rect 195 953 249 969
rect 417 969 427 1003
rect 461 989 541 1003
rect 599 1019 629 1050
rect 687 1019 717 1050
rect 599 1003 717 1019
rect 599 989 649 1003
rect 461 969 471 989
rect 417 953 471 969
rect 639 969 649 989
rect 683 989 717 1003
rect 1815 1450 1845 1476
rect 1903 1450 1933 1476
rect 1991 1450 2021 1476
rect 2079 1450 2109 1476
rect 683 969 693 989
rect 639 953 693 969
rect 1149 1019 1179 1050
rect 1237 1019 1267 1050
rect 1325 1019 1355 1050
rect 1413 1019 1443 1050
rect 1149 1003 1267 1019
rect 1149 989 1167 1003
rect 1157 969 1167 989
rect 1201 989 1267 1003
rect 1311 1003 1443 1019
rect 1201 969 1211 989
rect 1157 953 1211 969
rect 1311 969 1321 1003
rect 1355 989 1443 1003
rect 2481 1450 2511 1476
rect 2569 1450 2599 1476
rect 2657 1450 2687 1476
rect 2745 1450 2775 1476
rect 1355 969 1365 989
rect 1311 953 1365 969
rect 1815 1019 1845 1050
rect 1903 1019 1933 1050
rect 1991 1019 2021 1050
rect 2079 1019 2109 1050
rect 1815 1003 1933 1019
rect 1815 989 1833 1003
rect 1823 969 1833 989
rect 1867 989 1933 1003
rect 1977 1003 2109 1019
rect 1867 969 1877 989
rect 1823 953 1877 969
rect 1977 969 1987 1003
rect 2021 989 2109 1003
rect 3147 1450 3177 1476
rect 3235 1450 3265 1476
rect 3323 1450 3353 1476
rect 3411 1450 3441 1476
rect 2021 969 2031 989
rect 1977 953 2031 969
rect 2481 1019 2511 1050
rect 2569 1019 2599 1050
rect 2657 1019 2687 1050
rect 2745 1019 2775 1050
rect 2481 1003 2599 1019
rect 2481 989 2499 1003
rect 2489 969 2499 989
rect 2533 989 2599 1003
rect 2643 1003 2775 1019
rect 2533 969 2543 989
rect 2489 953 2543 969
rect 2643 969 2653 1003
rect 2687 989 2775 1003
rect 3813 1450 3843 1476
rect 3901 1450 3931 1476
rect 3989 1450 4019 1476
rect 4077 1450 4107 1476
rect 2687 969 2697 989
rect 2643 953 2697 969
rect 3147 1019 3177 1050
rect 3235 1019 3265 1050
rect 3323 1019 3353 1050
rect 3411 1019 3441 1050
rect 3147 1003 3265 1019
rect 3147 989 3165 1003
rect 3155 969 3165 989
rect 3199 989 3265 1003
rect 3309 1003 3441 1019
rect 3199 969 3209 989
rect 3155 953 3209 969
rect 3309 969 3319 1003
rect 3353 989 3441 1003
rect 3353 969 3363 989
rect 3309 953 3363 969
rect 3813 1019 3843 1050
rect 3901 1019 3931 1050
rect 3989 1019 4019 1050
rect 4077 1019 4107 1050
rect 3813 1003 3931 1019
rect 3813 989 3831 1003
rect 3821 969 3831 989
rect 3865 989 3931 1003
rect 3975 1003 4107 1019
rect 3865 969 3875 989
rect 3821 953 3875 969
rect 3975 969 3985 1003
rect 4019 989 4107 1003
rect 4019 969 4029 989
rect 3975 953 4029 969
rect 195 461 249 477
rect 195 441 205 461
rect 147 427 205 441
rect 239 427 249 461
rect 147 411 249 427
rect 417 461 471 477
rect 417 427 427 461
rect 461 441 471 461
rect 639 461 693 477
rect 461 427 477 441
rect 417 411 477 427
rect 639 427 649 461
rect 683 427 693 461
rect 639 411 693 427
rect 1157 461 1211 477
rect 1157 441 1167 461
rect 147 379 177 411
rect 447 379 477 411
rect 649 379 679 411
rect 1130 427 1167 441
rect 1201 427 1211 461
rect 1130 411 1211 427
rect 1305 461 1359 477
rect 1305 427 1315 461
rect 1349 427 1359 461
rect 1305 411 1359 427
rect 1823 461 1877 477
rect 1823 441 1833 461
rect 1130 377 1160 411
rect 1324 377 1354 411
rect 1796 427 1833 441
rect 1867 427 1877 461
rect 1796 411 1877 427
rect 1971 461 2025 477
rect 1971 427 1981 461
rect 2015 427 2025 461
rect 1971 411 2025 427
rect 2489 461 2543 477
rect 2489 441 2499 461
rect 1796 377 1826 411
rect 1990 377 2020 411
rect 2462 427 2499 441
rect 2533 427 2543 461
rect 2462 411 2543 427
rect 2637 461 2691 477
rect 2637 427 2647 461
rect 2681 427 2691 461
rect 2637 411 2691 427
rect 3155 461 3209 477
rect 3155 441 3165 461
rect 2462 377 2492 411
rect 2656 377 2686 411
rect 3128 427 3165 441
rect 3199 427 3209 461
rect 3128 411 3209 427
rect 3303 461 3357 477
rect 3303 427 3313 461
rect 3347 427 3357 461
rect 3303 411 3357 427
rect 3821 461 3875 477
rect 3821 441 3831 461
rect 3128 377 3158 411
rect 3322 377 3352 411
rect 3794 427 3831 441
rect 3865 427 3875 461
rect 3794 411 3875 427
rect 3969 461 4023 477
rect 3969 427 3979 461
rect 4013 427 4023 461
rect 3969 411 4023 427
rect 3794 377 3824 411
rect 3988 377 4018 411
<< polycont >>
rect 205 969 239 1003
rect 427 969 461 1003
rect 649 969 683 1003
rect 1167 969 1201 1003
rect 1321 969 1355 1003
rect 1833 969 1867 1003
rect 1987 969 2021 1003
rect 2499 969 2533 1003
rect 2653 969 2687 1003
rect 3165 969 3199 1003
rect 3319 969 3353 1003
rect 3831 969 3865 1003
rect 3985 969 4019 1003
rect 205 427 239 461
rect 427 427 461 461
rect 649 427 683 461
rect 1167 427 1201 461
rect 1315 427 1349 461
rect 1833 427 1867 461
rect 1981 427 2015 461
rect 2499 427 2533 461
rect 2647 427 2681 461
rect 3165 427 3199 461
rect 3313 427 3347 461
rect 3831 427 3865 461
rect 3979 427 4013 461
<< locali >>
rect -31 1539 4323 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1323 1539
rect 1357 1505 1395 1539
rect 1429 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1683 1539
rect 1717 1505 1755 1539
rect 1789 1505 1827 1539
rect 1861 1505 1899 1539
rect 1933 1505 1989 1539
rect 2023 1505 2061 1539
rect 2095 1505 2133 1539
rect 2167 1505 2205 1539
rect 2239 1505 2349 1539
rect 2383 1505 2421 1539
rect 2455 1505 2493 1539
rect 2527 1505 2565 1539
rect 2599 1505 2655 1539
rect 2689 1505 2727 1539
rect 2761 1505 2799 1539
rect 2833 1505 2871 1539
rect 2905 1505 3015 1539
rect 3049 1505 3087 1539
rect 3121 1505 3159 1539
rect 3193 1505 3231 1539
rect 3265 1505 3321 1539
rect 3355 1505 3393 1539
rect 3427 1505 3465 1539
rect 3499 1505 3537 1539
rect 3571 1505 3681 1539
rect 3715 1505 3753 1539
rect 3787 1505 3825 1539
rect 3859 1505 3897 1539
rect 3931 1505 3987 1539
rect 4021 1505 4059 1539
rect 4093 1505 4131 1539
rect 4165 1505 4203 1539
rect 4237 1505 4323 1539
rect -31 1492 4323 1505
rect -31 1470 31 1492
rect -31 1436 -17 1470
rect 17 1436 31 1470
rect -31 1398 31 1436
rect -31 1364 -17 1398
rect 17 1364 31 1398
rect -31 1326 31 1364
rect -31 1292 -17 1326
rect 17 1292 31 1326
rect -31 1254 31 1292
rect -31 1220 -17 1254
rect 17 1220 31 1254
rect -31 1182 31 1220
rect -31 1148 -17 1182
rect 17 1148 31 1182
rect -31 1110 31 1148
rect -31 1076 -17 1110
rect 17 1076 31 1110
rect 201 1412 235 1492
rect 201 1344 235 1378
rect 201 1276 235 1310
rect 201 1208 235 1242
rect 201 1139 235 1174
rect 201 1089 235 1105
rect 289 1412 323 1450
rect 289 1344 323 1378
rect 289 1276 323 1310
rect 289 1208 323 1242
rect 289 1139 323 1174
rect 377 1412 411 1492
rect 377 1344 411 1378
rect 377 1276 411 1310
rect 377 1208 411 1242
rect 377 1157 411 1174
rect 465 1412 499 1450
rect 465 1344 499 1378
rect 465 1276 499 1310
rect 465 1208 499 1242
rect 289 1094 323 1105
rect 465 1139 499 1174
rect 553 1412 587 1492
rect 553 1344 587 1378
rect 553 1276 587 1310
rect 553 1208 587 1242
rect 553 1157 587 1174
rect 641 1412 675 1450
rect 641 1344 675 1378
rect 641 1276 675 1310
rect 641 1208 675 1242
rect 465 1094 499 1105
rect 641 1139 675 1174
rect 729 1412 763 1492
rect 729 1344 763 1378
rect 729 1276 763 1310
rect 729 1208 763 1242
rect 729 1157 763 1174
rect 931 1470 993 1492
rect 931 1436 945 1470
rect 979 1436 993 1470
rect 931 1398 993 1436
rect 931 1364 945 1398
rect 979 1364 993 1398
rect 931 1326 993 1364
rect 931 1292 945 1326
rect 979 1292 993 1326
rect 931 1254 993 1292
rect 931 1220 945 1254
rect 979 1220 993 1254
rect 931 1182 993 1220
rect 641 1094 675 1105
rect 931 1148 945 1182
rect 979 1148 993 1182
rect 931 1110 993 1148
rect -31 1038 31 1076
rect 289 1060 831 1094
rect -31 1004 -17 1038
rect 17 1004 31 1038
rect -31 966 31 1004
rect -31 932 -17 966
rect 17 932 31 966
rect -31 868 31 932
rect 205 1003 239 1019
rect 205 905 239 969
rect -31 546 31 572
rect -31 512 -17 546
rect 17 512 31 546
rect -31 474 31 512
rect -31 440 -17 474
rect 17 440 31 474
rect -31 402 31 440
rect 205 461 239 871
rect 205 411 239 427
rect 427 1003 461 1019
rect 427 461 461 945
rect 427 411 461 427
rect 649 1003 683 1019
rect 649 757 683 969
rect 649 461 683 723
rect 649 411 683 427
rect 797 831 831 1060
rect 931 1076 945 1110
rect 979 1076 993 1110
rect 931 1038 993 1076
rect 1103 1412 1137 1492
rect 1103 1344 1137 1378
rect 1103 1276 1137 1310
rect 1103 1208 1137 1242
rect 1103 1139 1137 1174
rect 1103 1073 1137 1105
rect 1191 1412 1225 1450
rect 1191 1344 1225 1378
rect 1191 1276 1225 1310
rect 1191 1208 1225 1242
rect 1191 1139 1225 1174
rect 1279 1412 1313 1492
rect 1279 1344 1313 1378
rect 1279 1276 1313 1310
rect 1279 1208 1313 1242
rect 1279 1157 1313 1174
rect 1367 1412 1401 1450
rect 1367 1344 1401 1378
rect 1367 1276 1401 1310
rect 1367 1208 1401 1242
rect 1191 1103 1225 1105
rect 1367 1139 1401 1174
rect 1455 1412 1489 1492
rect 1455 1344 1489 1378
rect 1455 1276 1489 1310
rect 1455 1208 1489 1242
rect 1455 1157 1489 1174
rect 1597 1470 1659 1492
rect 1597 1436 1611 1470
rect 1645 1436 1659 1470
rect 1597 1398 1659 1436
rect 1597 1364 1611 1398
rect 1645 1364 1659 1398
rect 1597 1326 1659 1364
rect 1597 1292 1611 1326
rect 1645 1292 1659 1326
rect 1597 1254 1659 1292
rect 1597 1220 1611 1254
rect 1645 1220 1659 1254
rect 1597 1182 1659 1220
rect 1367 1103 1401 1105
rect 1597 1148 1611 1182
rect 1645 1148 1659 1182
rect 1597 1110 1659 1148
rect 1191 1069 1497 1103
rect 931 1004 945 1038
rect 979 1004 993 1038
rect 931 966 993 1004
rect 931 932 945 966
rect 979 932 993 966
rect 931 868 993 932
rect 1167 1003 1201 1019
rect 1321 1003 1355 1019
rect -31 368 -17 402
rect 17 368 31 402
rect -31 330 31 368
rect -31 296 -17 330
rect 17 296 31 330
rect -31 258 31 296
rect -31 224 -17 258
rect 17 224 31 258
rect -31 186 31 224
rect -31 152 -17 186
rect 17 152 31 186
rect -31 114 31 152
rect -31 80 -17 114
rect 17 80 31 114
rect 101 363 135 379
rect 295 363 329 379
rect 489 363 523 379
rect 135 329 198 363
rect 232 329 295 363
rect 329 329 392 363
rect 426 329 489 363
rect 101 291 135 329
rect 101 223 135 257
rect 295 291 329 329
rect 489 313 523 329
rect 603 363 637 379
rect 797 378 831 797
rect 1167 831 1201 969
rect 603 291 637 329
rect 101 153 135 189
rect 101 103 135 119
rect 198 238 232 254
rect -31 62 31 80
rect 198 62 232 204
rect 295 223 329 257
rect 393 244 427 260
rect 603 244 637 257
rect 427 223 637 244
rect 427 210 603 223
rect 393 194 427 210
rect 295 153 329 189
rect 700 344 831 378
rect 931 546 993 572
rect 931 512 945 546
rect 979 512 993 546
rect 931 474 993 512
rect 931 440 945 474
rect 979 440 993 474
rect 931 402 993 440
rect 1167 461 1201 797
rect 1167 411 1201 427
rect 1315 969 1321 988
rect 1315 953 1355 969
rect 1315 683 1349 953
rect 1315 461 1349 649
rect 1315 411 1349 427
rect 1463 757 1497 1069
rect 1597 1076 1611 1110
rect 1645 1076 1659 1110
rect 1597 1038 1659 1076
rect 1769 1412 1803 1492
rect 1769 1344 1803 1378
rect 1769 1276 1803 1310
rect 1769 1208 1803 1242
rect 1769 1139 1803 1174
rect 1769 1073 1803 1105
rect 1857 1412 1891 1450
rect 1857 1344 1891 1378
rect 1857 1276 1891 1310
rect 1857 1208 1891 1242
rect 1857 1139 1891 1174
rect 1945 1412 1979 1492
rect 1945 1344 1979 1378
rect 1945 1276 1979 1310
rect 1945 1208 1979 1242
rect 1945 1157 1979 1174
rect 2033 1412 2067 1450
rect 2033 1344 2067 1378
rect 2033 1276 2067 1310
rect 2033 1208 2067 1242
rect 1857 1103 1891 1105
rect 2033 1139 2067 1174
rect 2121 1412 2155 1492
rect 2121 1344 2155 1378
rect 2121 1276 2155 1310
rect 2121 1208 2155 1242
rect 2121 1157 2155 1174
rect 2263 1470 2325 1492
rect 2263 1436 2277 1470
rect 2311 1436 2325 1470
rect 2263 1398 2325 1436
rect 2263 1364 2277 1398
rect 2311 1364 2325 1398
rect 2263 1326 2325 1364
rect 2263 1292 2277 1326
rect 2311 1292 2325 1326
rect 2263 1254 2325 1292
rect 2263 1220 2277 1254
rect 2311 1220 2325 1254
rect 2263 1182 2325 1220
rect 2033 1103 2067 1105
rect 2263 1148 2277 1182
rect 2311 1148 2325 1182
rect 2263 1110 2325 1148
rect 1857 1069 2163 1103
rect 1597 1004 1611 1038
rect 1645 1004 1659 1038
rect 1597 966 1659 1004
rect 1597 932 1611 966
rect 1645 932 1659 966
rect 1597 868 1659 932
rect 1833 1003 1867 1019
rect 1987 1003 2021 1019
rect 931 368 945 402
rect 979 368 993 402
rect 700 247 734 344
rect 931 330 993 368
rect 700 197 734 213
rect 797 291 831 307
rect 797 223 831 257
rect 489 153 523 169
rect 329 119 392 153
rect 426 119 489 153
rect 295 103 329 119
rect 489 103 523 119
rect 603 153 637 189
rect 797 153 831 189
rect 637 119 700 153
rect 734 119 797 153
rect 603 103 637 119
rect 797 103 831 119
rect 931 296 945 330
rect 979 296 993 330
rect 931 258 993 296
rect 931 224 945 258
rect 979 224 993 258
rect 931 186 993 224
rect 931 152 945 186
rect 979 152 993 186
rect 931 114 993 152
rect 931 80 945 114
rect 979 80 993 114
rect 1084 361 1118 377
rect 1278 361 1312 377
rect 1463 376 1497 723
rect 1833 757 1867 969
rect 1118 327 1181 361
rect 1215 327 1278 361
rect 1084 289 1118 327
rect 1084 221 1118 255
rect 1278 289 1312 327
rect 1084 151 1118 187
rect 1084 101 1118 117
rect 1181 236 1215 252
rect 931 62 993 80
rect 1181 62 1215 202
rect 1278 221 1312 255
rect 1375 342 1497 376
rect 1597 546 1659 572
rect 1597 512 1611 546
rect 1645 512 1659 546
rect 1597 474 1659 512
rect 1597 440 1611 474
rect 1645 440 1659 474
rect 1597 402 1659 440
rect 1833 461 1867 723
rect 1833 411 1867 427
rect 1981 969 1987 988
rect 1981 953 2021 969
rect 1981 905 2015 953
rect 1981 461 2015 871
rect 1981 411 2015 427
rect 2129 757 2163 1069
rect 2263 1076 2277 1110
rect 2311 1076 2325 1110
rect 2263 1038 2325 1076
rect 2435 1412 2469 1492
rect 2435 1344 2469 1378
rect 2435 1276 2469 1310
rect 2435 1208 2469 1242
rect 2435 1139 2469 1174
rect 2435 1073 2469 1105
rect 2523 1412 2557 1450
rect 2523 1344 2557 1378
rect 2523 1276 2557 1310
rect 2523 1208 2557 1242
rect 2523 1139 2557 1174
rect 2611 1412 2645 1492
rect 2611 1344 2645 1378
rect 2611 1276 2645 1310
rect 2611 1208 2645 1242
rect 2611 1157 2645 1174
rect 2699 1412 2733 1450
rect 2699 1344 2733 1378
rect 2699 1276 2733 1310
rect 2699 1208 2733 1242
rect 2523 1103 2557 1105
rect 2699 1139 2733 1174
rect 2787 1412 2821 1492
rect 2787 1344 2821 1378
rect 2787 1276 2821 1310
rect 2787 1208 2821 1242
rect 2787 1157 2821 1174
rect 2929 1470 2991 1492
rect 2929 1436 2943 1470
rect 2977 1436 2991 1470
rect 2929 1398 2991 1436
rect 2929 1364 2943 1398
rect 2977 1364 2991 1398
rect 2929 1326 2991 1364
rect 2929 1292 2943 1326
rect 2977 1292 2991 1326
rect 2929 1254 2991 1292
rect 2929 1220 2943 1254
rect 2977 1220 2991 1254
rect 2929 1182 2991 1220
rect 2699 1103 2733 1105
rect 2929 1148 2943 1182
rect 2977 1148 2991 1182
rect 2929 1110 2991 1148
rect 2523 1069 2829 1103
rect 2263 1004 2277 1038
rect 2311 1004 2325 1038
rect 2263 966 2325 1004
rect 2263 932 2277 966
rect 2311 932 2325 966
rect 2263 868 2325 932
rect 2499 1003 2533 1019
rect 2653 1003 2687 1019
rect 1597 368 1611 402
rect 1645 368 1659 402
rect 1375 245 1409 342
rect 1597 330 1659 368
rect 1375 195 1409 211
rect 1472 289 1506 305
rect 1472 221 1506 255
rect 1278 151 1312 187
rect 1472 151 1506 187
rect 1312 117 1375 151
rect 1409 117 1472 151
rect 1278 101 1312 117
rect 1472 101 1506 117
rect 1597 296 1611 330
rect 1645 296 1659 330
rect 1597 258 1659 296
rect 1597 224 1611 258
rect 1645 224 1659 258
rect 1597 186 1659 224
rect 1597 152 1611 186
rect 1645 152 1659 186
rect 1597 114 1659 152
rect 1597 80 1611 114
rect 1645 80 1659 114
rect 1750 361 1784 377
rect 1944 361 1978 377
rect 2129 376 2163 723
rect 2499 757 2533 969
rect 1784 327 1847 361
rect 1881 327 1944 361
rect 1750 289 1784 327
rect 1750 221 1784 255
rect 1944 289 1978 327
rect 1750 151 1784 187
rect 1750 101 1784 117
rect 1847 236 1881 252
rect 1597 62 1659 80
rect 1847 62 1881 202
rect 1944 221 1978 255
rect 2041 342 2163 376
rect 2263 546 2325 572
rect 2263 512 2277 546
rect 2311 512 2325 546
rect 2263 474 2325 512
rect 2263 440 2277 474
rect 2311 440 2325 474
rect 2263 402 2325 440
rect 2499 461 2533 723
rect 2499 411 2533 427
rect 2647 979 2653 995
rect 2681 953 2687 969
rect 2647 461 2681 945
rect 2647 411 2681 427
rect 2795 905 2829 1069
rect 2263 368 2277 402
rect 2311 368 2325 402
rect 2041 245 2075 342
rect 2263 330 2325 368
rect 2041 195 2075 211
rect 2138 289 2172 305
rect 2138 221 2172 255
rect 1944 151 1978 187
rect 2138 151 2172 187
rect 1978 117 2041 151
rect 2075 117 2138 151
rect 1944 101 1978 117
rect 2138 101 2172 117
rect 2263 296 2277 330
rect 2311 296 2325 330
rect 2263 258 2325 296
rect 2263 224 2277 258
rect 2311 224 2325 258
rect 2263 186 2325 224
rect 2263 152 2277 186
rect 2311 152 2325 186
rect 2263 114 2325 152
rect 2263 80 2277 114
rect 2311 80 2325 114
rect 2416 361 2450 377
rect 2610 361 2644 377
rect 2795 376 2829 871
rect 2929 1076 2943 1110
rect 2977 1076 2991 1110
rect 2929 1038 2991 1076
rect 3101 1412 3135 1492
rect 3101 1344 3135 1378
rect 3101 1276 3135 1310
rect 3101 1208 3135 1242
rect 3101 1139 3135 1174
rect 3101 1073 3135 1105
rect 3189 1412 3223 1450
rect 3189 1344 3223 1378
rect 3189 1276 3223 1310
rect 3189 1208 3223 1242
rect 3189 1139 3223 1174
rect 3277 1412 3311 1492
rect 3277 1344 3311 1378
rect 3277 1276 3311 1310
rect 3277 1208 3311 1242
rect 3277 1157 3311 1174
rect 3365 1412 3399 1450
rect 3365 1344 3399 1378
rect 3365 1276 3399 1310
rect 3365 1208 3399 1242
rect 3189 1103 3223 1105
rect 3365 1139 3399 1174
rect 3453 1412 3487 1492
rect 3453 1344 3487 1378
rect 3453 1276 3487 1310
rect 3453 1208 3487 1242
rect 3453 1157 3487 1174
rect 3595 1470 3657 1492
rect 3595 1436 3609 1470
rect 3643 1436 3657 1470
rect 3595 1398 3657 1436
rect 3595 1364 3609 1398
rect 3643 1364 3657 1398
rect 3595 1326 3657 1364
rect 3595 1292 3609 1326
rect 3643 1292 3657 1326
rect 3595 1254 3657 1292
rect 3595 1220 3609 1254
rect 3643 1220 3657 1254
rect 3595 1182 3657 1220
rect 3365 1103 3399 1105
rect 3595 1148 3609 1182
rect 3643 1148 3657 1182
rect 3595 1110 3657 1148
rect 3189 1069 3495 1103
rect 2929 1004 2943 1038
rect 2977 1004 2991 1038
rect 2929 966 2991 1004
rect 2929 932 2943 966
rect 2977 932 2991 966
rect 2929 868 2991 932
rect 3165 1003 3199 1019
rect 3319 1003 3353 1019
rect 3165 831 3199 969
rect 2450 327 2513 361
rect 2547 327 2610 361
rect 2416 289 2450 327
rect 2416 221 2450 255
rect 2610 289 2644 327
rect 2416 151 2450 187
rect 2416 101 2450 117
rect 2513 236 2547 252
rect 2263 62 2325 80
rect 2513 62 2547 202
rect 2610 221 2644 255
rect 2707 342 2829 376
rect 2929 546 2991 572
rect 2929 512 2943 546
rect 2977 512 2991 546
rect 2929 474 2991 512
rect 2929 440 2943 474
rect 2977 440 2991 474
rect 2929 402 2991 440
rect 3165 461 3199 797
rect 3165 411 3199 427
rect 3313 969 3319 988
rect 3313 953 3353 969
rect 3313 831 3347 953
rect 3313 461 3347 797
rect 3313 411 3347 427
rect 3461 757 3495 1069
rect 3595 1076 3609 1110
rect 3643 1076 3657 1110
rect 3595 1038 3657 1076
rect 3767 1412 3801 1492
rect 3767 1344 3801 1378
rect 3767 1276 3801 1310
rect 3767 1208 3801 1242
rect 3767 1139 3801 1174
rect 3767 1073 3801 1105
rect 3855 1412 3889 1450
rect 3855 1344 3889 1378
rect 3855 1276 3889 1310
rect 3855 1208 3889 1242
rect 3855 1139 3889 1174
rect 3943 1412 3977 1492
rect 3943 1344 3977 1378
rect 3943 1276 3977 1310
rect 3943 1208 3977 1242
rect 3943 1157 3977 1174
rect 4031 1412 4065 1450
rect 4031 1344 4065 1378
rect 4031 1276 4065 1310
rect 4031 1208 4065 1242
rect 3855 1103 3889 1105
rect 4031 1139 4065 1174
rect 4119 1412 4153 1492
rect 4119 1344 4153 1378
rect 4119 1276 4153 1310
rect 4119 1208 4153 1242
rect 4119 1157 4153 1174
rect 4261 1470 4323 1492
rect 4261 1436 4275 1470
rect 4309 1436 4323 1470
rect 4261 1398 4323 1436
rect 4261 1364 4275 1398
rect 4309 1364 4323 1398
rect 4261 1326 4323 1364
rect 4261 1292 4275 1326
rect 4309 1292 4323 1326
rect 4261 1254 4323 1292
rect 4261 1220 4275 1254
rect 4309 1220 4323 1254
rect 4261 1182 4323 1220
rect 4031 1103 4065 1105
rect 4261 1148 4275 1182
rect 4309 1148 4323 1182
rect 4261 1110 4323 1148
rect 3855 1069 4161 1103
rect 3595 1004 3609 1038
rect 3643 1004 3657 1038
rect 3595 966 3657 1004
rect 3595 932 3609 966
rect 3643 932 3657 966
rect 3595 868 3657 932
rect 3831 1003 3865 1019
rect 3985 1003 4019 1019
rect 2929 368 2943 402
rect 2977 368 2991 402
rect 2707 245 2741 342
rect 2929 330 2991 368
rect 2707 195 2741 211
rect 2804 289 2838 305
rect 2804 221 2838 255
rect 2610 151 2644 187
rect 2804 151 2838 187
rect 2644 117 2707 151
rect 2741 117 2804 151
rect 2610 101 2644 117
rect 2804 101 2838 117
rect 2929 296 2943 330
rect 2977 296 2991 330
rect 2929 258 2991 296
rect 2929 224 2943 258
rect 2977 224 2991 258
rect 2929 186 2991 224
rect 2929 152 2943 186
rect 2977 152 2991 186
rect 2929 114 2991 152
rect 2929 80 2943 114
rect 2977 80 2991 114
rect 3082 361 3116 377
rect 3276 361 3310 377
rect 3461 376 3495 723
rect 3831 757 3865 969
rect 3116 327 3179 361
rect 3213 327 3276 361
rect 3082 289 3116 327
rect 3082 221 3116 255
rect 3276 289 3310 327
rect 3082 151 3116 187
rect 3082 101 3116 117
rect 3179 236 3213 252
rect 2929 62 2991 80
rect 3179 62 3213 202
rect 3276 221 3310 255
rect 3373 342 3495 376
rect 3595 546 3657 572
rect 3595 512 3609 546
rect 3643 512 3657 546
rect 3595 474 3657 512
rect 3595 440 3609 474
rect 3643 440 3657 474
rect 3595 402 3657 440
rect 3831 461 3865 723
rect 3831 411 3865 427
rect 3979 969 3985 988
rect 3979 953 4019 969
rect 3979 905 4013 953
rect 3979 461 4013 871
rect 3979 411 4013 427
rect 4127 831 4161 1069
rect 4261 1076 4275 1110
rect 4309 1076 4323 1110
rect 4261 1038 4323 1076
rect 4261 1004 4275 1038
rect 4309 1004 4323 1038
rect 4261 966 4323 1004
rect 4261 932 4275 966
rect 4309 932 4323 966
rect 4261 868 4323 932
rect 3595 368 3609 402
rect 3643 368 3657 402
rect 3373 245 3407 342
rect 3595 330 3657 368
rect 3373 195 3407 211
rect 3470 289 3504 305
rect 3470 221 3504 255
rect 3276 151 3310 187
rect 3470 151 3504 187
rect 3310 117 3373 151
rect 3407 117 3470 151
rect 3276 101 3310 117
rect 3470 101 3504 117
rect 3595 296 3609 330
rect 3643 296 3657 330
rect 3595 258 3657 296
rect 3595 224 3609 258
rect 3643 224 3657 258
rect 3595 186 3657 224
rect 3595 152 3609 186
rect 3643 152 3657 186
rect 3595 114 3657 152
rect 3595 80 3609 114
rect 3643 80 3657 114
rect 3748 361 3782 377
rect 3942 361 3976 377
rect 4127 376 4161 797
rect 3782 327 3845 361
rect 3879 327 3942 361
rect 3748 289 3782 327
rect 3748 221 3782 255
rect 3942 289 3976 327
rect 3748 151 3782 187
rect 3748 101 3782 117
rect 3845 236 3879 252
rect 3595 62 3657 80
rect 3845 62 3879 202
rect 3942 221 3976 255
rect 4039 342 4161 376
rect 4261 546 4323 572
rect 4261 512 4275 546
rect 4309 512 4323 546
rect 4261 474 4323 512
rect 4261 440 4275 474
rect 4309 440 4323 474
rect 4261 402 4323 440
rect 4261 368 4275 402
rect 4309 368 4323 402
rect 4039 245 4073 342
rect 4261 330 4323 368
rect 4039 195 4073 211
rect 4136 289 4170 305
rect 4136 221 4170 255
rect 3942 151 3976 187
rect 4136 151 4170 187
rect 3976 117 4039 151
rect 4073 117 4136 151
rect 3942 101 3976 117
rect 4136 101 4170 117
rect 4261 296 4275 330
rect 4309 296 4323 330
rect 4261 258 4323 296
rect 4261 224 4275 258
rect 4309 224 4323 258
rect 4261 186 4323 224
rect 4261 152 4275 186
rect 4309 152 4323 186
rect 4261 114 4323 152
rect 4261 80 4275 114
rect 4309 80 4323 114
rect 4261 62 4323 80
rect -31 47 4323 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1323 47
rect 1357 13 1395 47
rect 1429 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1683 47
rect 1717 13 1755 47
rect 1789 13 1827 47
rect 1861 13 1899 47
rect 1933 13 1989 47
rect 2023 13 2061 47
rect 2095 13 2133 47
rect 2167 13 2205 47
rect 2239 13 2349 47
rect 2383 13 2421 47
rect 2455 13 2493 47
rect 2527 13 2565 47
rect 2599 13 2655 47
rect 2689 13 2727 47
rect 2761 13 2799 47
rect 2833 13 2871 47
rect 2905 13 3015 47
rect 3049 13 3087 47
rect 3121 13 3159 47
rect 3193 13 3231 47
rect 3265 13 3321 47
rect 3355 13 3393 47
rect 3427 13 3465 47
rect 3499 13 3537 47
rect 3571 13 3681 47
rect 3715 13 3753 47
rect 3787 13 3825 47
rect 3859 13 3897 47
rect 3931 13 3987 47
rect 4021 13 4059 47
rect 4093 13 4131 47
rect 4165 13 4203 47
rect 4237 13 4323 47
rect -31 0 4323 13
<< viali >>
rect 55 1505 89 1539
rect 127 1505 161 1539
rect 199 1505 233 1539
rect 271 1505 305 1539
rect 343 1505 377 1539
rect 415 1505 449 1539
rect 513 1505 547 1539
rect 585 1505 619 1539
rect 657 1505 691 1539
rect 729 1505 763 1539
rect 801 1505 835 1539
rect 873 1505 907 1539
rect 1017 1505 1051 1539
rect 1089 1505 1123 1539
rect 1161 1505 1195 1539
rect 1233 1505 1267 1539
rect 1323 1505 1357 1539
rect 1395 1505 1429 1539
rect 1467 1505 1501 1539
rect 1539 1505 1573 1539
rect 1683 1505 1717 1539
rect 1755 1505 1789 1539
rect 1827 1505 1861 1539
rect 1899 1505 1933 1539
rect 1989 1505 2023 1539
rect 2061 1505 2095 1539
rect 2133 1505 2167 1539
rect 2205 1505 2239 1539
rect 2349 1505 2383 1539
rect 2421 1505 2455 1539
rect 2493 1505 2527 1539
rect 2565 1505 2599 1539
rect 2655 1505 2689 1539
rect 2727 1505 2761 1539
rect 2799 1505 2833 1539
rect 2871 1505 2905 1539
rect 3015 1505 3049 1539
rect 3087 1505 3121 1539
rect 3159 1505 3193 1539
rect 3231 1505 3265 1539
rect 3321 1505 3355 1539
rect 3393 1505 3427 1539
rect 3465 1505 3499 1539
rect 3537 1505 3571 1539
rect 3681 1505 3715 1539
rect 3753 1505 3787 1539
rect 3825 1505 3859 1539
rect 3897 1505 3931 1539
rect 3987 1505 4021 1539
rect 4059 1505 4093 1539
rect 4131 1505 4165 1539
rect 4203 1505 4237 1539
rect 205 871 239 905
rect 427 969 461 979
rect 427 945 461 969
rect 649 723 683 757
rect 797 797 831 831
rect 1167 797 1201 831
rect 1315 649 1349 683
rect 1315 427 1349 461
rect 1463 723 1497 757
rect 1833 723 1867 757
rect 1981 871 2015 905
rect 2129 723 2163 757
rect 2499 723 2533 757
rect 2647 969 2653 979
rect 2653 969 2681 979
rect 2647 945 2681 969
rect 2795 871 2829 905
rect 3165 797 3199 831
rect 3313 797 3347 831
rect 3461 723 3495 757
rect 3831 723 3865 757
rect 3979 871 4013 905
rect 4127 797 4161 831
rect 55 13 89 47
rect 127 13 161 47
rect 199 13 233 47
rect 271 13 305 47
rect 343 13 377 47
rect 415 13 449 47
rect 513 13 547 47
rect 585 13 619 47
rect 657 13 691 47
rect 729 13 763 47
rect 801 13 835 47
rect 873 13 907 47
rect 1017 13 1051 47
rect 1089 13 1123 47
rect 1161 13 1195 47
rect 1233 13 1267 47
rect 1323 13 1357 47
rect 1395 13 1429 47
rect 1467 13 1501 47
rect 1539 13 1573 47
rect 1683 13 1717 47
rect 1755 13 1789 47
rect 1827 13 1861 47
rect 1899 13 1933 47
rect 1989 13 2023 47
rect 2061 13 2095 47
rect 2133 13 2167 47
rect 2205 13 2239 47
rect 2349 13 2383 47
rect 2421 13 2455 47
rect 2493 13 2527 47
rect 2565 13 2599 47
rect 2655 13 2689 47
rect 2727 13 2761 47
rect 2799 13 2833 47
rect 2871 13 2905 47
rect 3015 13 3049 47
rect 3087 13 3121 47
rect 3159 13 3193 47
rect 3231 13 3265 47
rect 3321 13 3355 47
rect 3393 13 3427 47
rect 3465 13 3499 47
rect 3537 13 3571 47
rect 3681 13 3715 47
rect 3753 13 3787 47
rect 3825 13 3859 47
rect 3897 13 3931 47
rect 3987 13 4021 47
rect 4059 13 4093 47
rect 4131 13 4165 47
rect 4203 13 4237 47
<< metal1 >>
rect -31 1539 4323 1554
rect -31 1505 55 1539
rect 89 1505 127 1539
rect 161 1505 199 1539
rect 233 1505 271 1539
rect 305 1505 343 1539
rect 377 1505 415 1539
rect 449 1505 513 1539
rect 547 1505 585 1539
rect 619 1505 657 1539
rect 691 1505 729 1539
rect 763 1505 801 1539
rect 835 1505 873 1539
rect 907 1505 1017 1539
rect 1051 1505 1089 1539
rect 1123 1505 1161 1539
rect 1195 1505 1233 1539
rect 1267 1505 1323 1539
rect 1357 1505 1395 1539
rect 1429 1505 1467 1539
rect 1501 1505 1539 1539
rect 1573 1505 1683 1539
rect 1717 1505 1755 1539
rect 1789 1505 1827 1539
rect 1861 1505 1899 1539
rect 1933 1505 1989 1539
rect 2023 1505 2061 1539
rect 2095 1505 2133 1539
rect 2167 1505 2205 1539
rect 2239 1505 2349 1539
rect 2383 1505 2421 1539
rect 2455 1505 2493 1539
rect 2527 1505 2565 1539
rect 2599 1505 2655 1539
rect 2689 1505 2727 1539
rect 2761 1505 2799 1539
rect 2833 1505 2871 1539
rect 2905 1505 3015 1539
rect 3049 1505 3087 1539
rect 3121 1505 3159 1539
rect 3193 1505 3231 1539
rect 3265 1505 3321 1539
rect 3355 1505 3393 1539
rect 3427 1505 3465 1539
rect 3499 1505 3537 1539
rect 3571 1505 3681 1539
rect 3715 1505 3753 1539
rect 3787 1505 3825 1539
rect 3859 1505 3897 1539
rect 3931 1505 3987 1539
rect 4021 1505 4059 1539
rect 4093 1505 4131 1539
rect 4165 1505 4203 1539
rect 4237 1505 4323 1539
rect -31 1492 4323 1505
rect 421 979 467 985
rect 2641 979 2687 985
rect 415 945 427 979
rect 461 945 2647 979
rect 2681 945 2693 979
rect 421 939 467 945
rect 2641 939 2687 945
rect 199 905 245 911
rect 1975 905 2021 911
rect 2789 905 2835 911
rect 3973 905 4019 911
rect 193 871 205 905
rect 239 871 1981 905
rect 2015 871 2795 905
rect 2829 871 3979 905
rect 4013 871 4025 905
rect 199 865 245 871
rect 1975 865 2021 871
rect 2789 865 2835 871
rect 3973 865 4019 871
rect 791 831 837 837
rect 1161 831 1207 837
rect 3159 831 3205 837
rect 3307 831 3353 837
rect 4121 831 4167 837
rect 785 797 797 831
rect 831 797 1167 831
rect 1201 797 3165 831
rect 3199 797 3211 831
rect 3301 797 3313 831
rect 3347 797 4127 831
rect 4161 797 4173 831
rect 791 791 837 797
rect 1161 791 1207 797
rect 3159 791 3205 797
rect 3307 791 3353 797
rect 4121 791 4167 797
rect 643 757 689 763
rect 1457 757 1503 763
rect 1827 757 1873 763
rect 2123 757 2169 763
rect 2493 757 2539 763
rect 3455 757 3501 763
rect 3825 757 3871 763
rect 637 723 649 757
rect 683 723 1463 757
rect 1497 723 1833 757
rect 1867 723 1879 757
rect 2117 723 2129 757
rect 2163 723 2499 757
rect 2533 723 2545 757
rect 3449 723 3461 757
rect 3495 723 3831 757
rect 3865 723 3877 757
rect 643 717 689 723
rect 1457 717 1503 723
rect 1827 717 1873 723
rect 2123 717 2169 723
rect 2493 717 2539 723
rect 3455 717 3501 723
rect 3825 717 3871 723
rect 1309 683 1355 689
rect 1279 649 1315 683
rect 1349 649 1361 683
rect 1309 643 1355 649
rect 1309 461 1355 467
rect 1279 427 1315 461
rect 1349 427 1361 461
rect 1309 421 1355 427
rect -31 47 4323 62
rect -31 13 55 47
rect 89 13 127 47
rect 161 13 199 47
rect 233 13 271 47
rect 305 13 343 47
rect 377 13 415 47
rect 449 13 513 47
rect 547 13 585 47
rect 619 13 657 47
rect 691 13 729 47
rect 763 13 801 47
rect 835 13 873 47
rect 907 13 1017 47
rect 1051 13 1089 47
rect 1123 13 1161 47
rect 1195 13 1233 47
rect 1267 13 1323 47
rect 1357 13 1395 47
rect 1429 13 1467 47
rect 1501 13 1539 47
rect 1573 13 1683 47
rect 1717 13 1755 47
rect 1789 13 1827 47
rect 1861 13 1899 47
rect 1933 13 1989 47
rect 2023 13 2061 47
rect 2095 13 2133 47
rect 2167 13 2205 47
rect 2239 13 2349 47
rect 2383 13 2421 47
rect 2455 13 2493 47
rect 2527 13 2565 47
rect 2599 13 2655 47
rect 2689 13 2727 47
rect 2761 13 2799 47
rect 2833 13 2871 47
rect 2905 13 3015 47
rect 3049 13 3087 47
rect 3121 13 3159 47
rect 3193 13 3231 47
rect 3265 13 3321 47
rect 3355 13 3393 47
rect 3427 13 3465 47
rect 3499 13 3537 47
rect 3571 13 3681 47
rect 3715 13 3753 47
rect 3787 13 3825 47
rect 3859 13 3897 47
rect 3931 13 3987 47
rect 4021 13 4059 47
rect 4093 13 4131 47
rect 4165 13 4203 47
rect 4237 13 4323 47
rect -31 0 4323 13
<< labels >>
rlabel metal1 4127 797 4161 831 1 Q
port 1 n
rlabel metal1 1315 649 1349 683 1 D
port 2 n
rlabel metal1 427 945 461 979 1 CLK
port 3 n
rlabel metal1 -31 1492 4323 1554 1 VDD
port 4 n
rlabel metal1 -31 0 4323 62 1 GND
port 5 n
<< end >>
