* SPICE3 file created from TMRDFFQNX1.ext - technology: sky130A

.subckt TMRDFFQNX1 QN D CLK VPB VNB
M1000 a_13093_1005.t2 a_11887_383.t5 VPB.t53 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 VPB.t33 a_147_159.t5 a_1845_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_6137_1004.t4 a_4891_943.t5 VPB.t16 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPB.t7 a_4569_1004.t7 a_4891_943.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_13093_1005.t3 a_11887_383.t6 a_13757_1005.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPB.t26 a_4439_159.t6 a_7595_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPB.t21 a_147_159.t6 a_277_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPB.t5 a_6137_1004.t5 a_4439_159.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VNB a_8861_1004.t11 a_11656_73.t0 nshort w=-1.605u l=1.765u
+  ad=3.7611p pd=32.97u as=0p ps=0u
M1009 VPB.t81 a_8731_159.t5 a_8861_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_3177_1004.t3 a_277_1004.t7 VPB.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPB.t6 a_1845_1004.t5 a_147_159.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_11887_383.t1 a_11761_1004.t5 VPB.t40 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPB.t48 D a_9183_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VNB a_10429_1004.t5 a_10990_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1015 VNB a_8731_159.t9 a_8675_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPB.t43 D a_4891_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPB.t49 a_7469_1004.t5 a_7595_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPB.t70 CLK a_277_1004.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VNB a_4569_1004.t8 a_5366_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1020 VNB a_599_943.t5 a_1740_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_13757_1005.t1 a_7595_383.t5 a_13268_181.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VNB a_11887_383.t7 a_13654_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_3177_1004.t0 a_3303_383.t5 VPB.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPB.t65 CLK a_147_159.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_11887_383.t4 a_8731_159.t6 VPB.t79 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPB.t56 a_11887_383.t9 a_11761_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 VNB a_11887_383.t8 a_12988_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPB.t72 CLK a_4439_159.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_9183_943.t1 D VPB.t44 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_3303_383.t1 a_3177_1004.t6 VPB.t41 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPB.t29 a_599_943.t6 a_277_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 VNB a_147_159.t13 a_91_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPB.t10 a_277_1004.t8 a_599_943.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_8731_159.t1 a_10429_1004.t6 VPB.t37 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_4569_1004.t3 a_4891_943.t6 VPB.t61 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_13757_1005.t3 a_3303_383.t6 a_13268_181.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPB.t31 a_9183_943.t7 a_10429_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPB.t8 a_147_159.t7 a_3303_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_7595_383.t4 a_7469_1004.t6 VPB.t50 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 VNB a_4569_1004.t9 a_7364_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1041 VNB a_3177_1004.t5 a_3738_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPB.t3 a_4569_1004.t10 a_7469_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1043 VNB a_9183_943.t5 a_10324_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_4439_159.t2 CLK VPB.t71 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_1845_1004.t1 a_147_159.t8 VPB.t60 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_8861_1004.t4 a_9183_943.t8 VPB.t52 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPB.t24 a_4439_159.t8 a_4569_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_6137_1004.t1 a_4439_159.t9 VPB.t22 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_9183_943.t4 a_8861_1004.t7 VPB.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 VNB a_4439_159.t5 a_4383_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_13093_1005.t0 a_3303_383.t7 a_13757_1005.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 a_11761_1004.t0 a_11887_383.t11 VPB.t55 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 a_3303_383.t2 a_147_159.t10 VPB.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1054 VPB.t63 a_7595_383.t6 a_13093_1005.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 VNB a_277_1004.t9 a_1074_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1056 VPB.t46 D a_599_943.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_13757_1005.t5 a_11887_383.t12 a_13093_1005.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 a_8731_159.t4 CLK VPB.t76 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1059 VPB.t38 a_8731_159.t7 a_10429_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1060 a_277_1004.t2 a_147_159.t11 VPB.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 a_4439_159.t0 a_6137_1004.t6 VPB.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 VPB.t64 a_7595_383.t7 a_7469_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 VPB.t68 CLK a_4569_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1064 VPB.t58 a_599_943.t7 a_1845_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 a_11761_1004.t4 a_8861_1004.t8 VPB.t51 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 VNB a_11761_1004.t6 a_12322_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1067 VPB.t54 a_11887_383.t13 a_13093_1005.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_4891_943.t2 D VPB.t47 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 a_13757_1005.t7 a_3303_383.t10 a_13093_1005.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 a_277_1004.t4 CLK VPB.t69 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 VNB a_6137_1004.t7 a_6698_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1072 VNB a_277_1004.t10 a_3072_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1073 VPB.t13 a_4891_943.t8 a_4569_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1074 VPB.t14 a_277_1004.t11 a_3177_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 a_147_159.t3 CLK VPB.t66 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1076 VPB.t78 a_11761_1004.t7 a_11887_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 VNB a_4891_943.t7 a_6032_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1078 VNB a_3303_383.t9 a_14320_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1079 a_4891_943.t0 a_4569_1004.t11 VPB.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 a_7595_383.t0 a_4439_159.t10 VPB.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 a_277_1004.t1 a_599_943.t8 VPB.t30 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1082 a_599_943.t3 a_277_1004.t12 VPB.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_8861_1004.t0 a_8731_159.t10 VPB.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 a_13268_181.t1 a_3303_383.t11 a_13757_1005.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 VPB.t74 CLK a_8731_159.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_10429_1004.t1 a_9183_943.t9 VPB.t34 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 a_147_159.t1 a_1845_1004.t6 VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 a_7469_1004.t0 a_4569_1004.t12 VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 VPB.t80 a_3303_383.t12 a_3177_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 VPB.t32 a_8731_159.t12 a_11887_383.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 VPB.t75 CLK a_8861_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1092 a_4569_1004.t0 a_4439_159.t11 VPB.t25 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1093 VPB.t15 a_4891_943.t9 a_6137_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 VNB a_7469_1004.t7 a_8030_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1095 VPB.t59 a_8861_1004.t10 a_11761_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1096 VPB.t57 a_3177_1004.t7 a_3303_383.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 a_13093_1005.t6 a_7595_383.t10 VPB.t62 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 a_599_943.t1 D VPB.t45 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1099 VPB.t36 a_10429_1004.t7 a_8731_159.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 VNB a_1845_1004.t7 a_2406_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1101 a_13268_181.t4 a_7595_383.t11 a_13757_1005.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1102 a_10429_1004.t3 a_8731_159.t13 VPB.t42 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_7469_1004.t3 a_7595_383.t12 VPB.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 VNB a_8861_1004.t9 a_9658_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1105 VPB.t39 a_9183_943.t10 a_8861_1004.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 a_4569_1004.t5 CLK VPB.t67 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 VPB.t23 a_4439_159.t13 a_6137_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 VPB.t35 a_8861_1004.t12 a_9183_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 a_1845_1004.t4 a_599_943.t10 VPB.t77 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 a_8861_1004.t5 CLK VPB.t73 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 D CLK 1.40fF
C1 VPB D 0.22fF
C2 VPB CLK 3.13fF
R0 a_10429_1004.n3 a_10429_1004.t7 480.392
R1 a_10429_1004.n3 a_10429_1004.t6 403.272
R2 a_10429_1004.n4 a_10429_1004.t5 266.974
R3 a_10429_1004.n7 a_10429_1004.n5 200.608
R4 a_10429_1004.n5 a_10429_1004.n2 162.547
R5 a_10429_1004.n5 a_10429_1004.n4 153.315
R6 a_10429_1004.n4 a_10429_1004.n3 108.494
R7 a_10429_1004.n2 a_10429_1004.n1 76.002
R8 a_10429_1004.n7 a_10429_1004.n6 15.218
R9 a_10429_1004.n0 a_10429_1004.t2 14.282
R10 a_10429_1004.n0 a_10429_1004.t3 14.282
R11 a_10429_1004.n1 a_10429_1004.t0 14.282
R12 a_10429_1004.n1 a_10429_1004.t1 14.282
R13 a_10429_1004.n2 a_10429_1004.n0 12.85
R14 a_10429_1004.n8 a_10429_1004.n7 12.014
R15 a_10990_73.t0 a_10990_73.n6 93.333
R16 a_10990_73.n4 a_10990_73.n3 41.622
R17 a_10990_73.t0 a_10990_73.n4 21.209
R18 a_10990_73.t0 a_10990_73.n5 11.595
R19 a_10990_73.t0 a_10990_73.n7 8.137
R20 a_10990_73.n2 a_10990_73.n0 4.031
R21 a_10990_73.n2 a_10990_73.n1 3.644
R22 a_10990_73.t0 a_10990_73.n2 1.093
R23 VNB VNB.n1157 300.778
R24 VNB.n174 VNB.n173 199.897
R25 VNB.n226 VNB.n225 199.897
R26 VNB.n278 VNB.n277 199.897
R27 VNB.n330 VNB.n329 199.897
R28 VNB.n382 VNB.n381 199.897
R29 VNB.n434 VNB.n433 199.897
R30 VNB.n486 VNB.n485 199.897
R31 VNB.n538 VNB.n537 199.897
R32 VNB.n606 VNB.n605 199.897
R33 VNB.n68 VNB.n67 199.897
R34 VNB.n658 VNB.n657 199.897
R35 VNB.n710 VNB.n709 199.897
R36 VNB.n762 VNB.n761 199.897
R37 VNB.n814 VNB.n813 199.897
R38 VNB.n882 VNB.n881 199.897
R39 VNB.n934 VNB.n933 199.897
R40 VNB.n986 VNB.n985 199.897
R41 VNB.n1038 VNB.n1037 199.897
R42 VNB.n1090 VNB.n1089 199.897
R43 VNB.n15 VNB.n14 199.897
R44 VNB.n183 VNB.n181 154.509
R45 VNB.n287 VNB.n285 154.509
R46 VNB.n235 VNB.n233 154.509
R47 VNB.n391 VNB.n389 154.509
R48 VNB.n339 VNB.n337 154.509
R49 VNB.n495 VNB.n493 154.509
R50 VNB.n443 VNB.n441 154.509
R51 VNB.n615 VNB.n613 154.509
R52 VNB.n547 VNB.n545 154.509
R53 VNB.n667 VNB.n665 154.509
R54 VNB.n101 VNB.n99 154.509
R55 VNB.n771 VNB.n769 154.509
R56 VNB.n719 VNB.n717 154.509
R57 VNB.n891 VNB.n889 154.509
R58 VNB.n823 VNB.n821 154.509
R59 VNB.n995 VNB.n993 154.509
R60 VNB.n943 VNB.n941 154.509
R61 VNB.n1099 VNB.n1097 154.509
R62 VNB.n1047 VNB.n1045 154.509
R63 VNB.n24 VNB.n22 154.509
R64 VNB.n82 VNB.n81 121.366
R65 VNB.n583 VNB.n582 85.559
R66 VNB.n859 VNB.n858 85.559
R67 VNB.n53 VNB.n4 85.559
R68 VNB.n151 VNB.n150 84.842
R69 VNB.n203 VNB.n202 84.842
R70 VNB.n255 VNB.n254 84.842
R71 VNB.n307 VNB.n306 84.842
R72 VNB.n359 VNB.n358 84.842
R73 VNB.n411 VNB.n410 84.842
R74 VNB.n463 VNB.n462 84.842
R75 VNB.n515 VNB.n514 84.842
R76 VNB.n115 VNB.n57 84.842
R77 VNB.n687 VNB.n686 84.842
R78 VNB.n739 VNB.n738 84.842
R79 VNB.n791 VNB.n790 84.842
R80 VNB.n911 VNB.n910 84.842
R81 VNB.n963 VNB.n962 84.842
R82 VNB.n1015 VNB.n1014 84.842
R83 VNB.n1067 VNB.n1066 84.842
R84 VNB.n1119 VNB.n1118 84.842
R85 VNB.n1144 VNB.n1143 76
R86 VNB.n1131 VNB.n1130 76
R87 VNB.n1127 VNB.n1126 76
R88 VNB.n1123 VNB.n1122 76
R89 VNB.n1117 VNB.n1116 76
R90 VNB.n1113 VNB.n1112 76
R91 VNB.n1109 VNB.n1108 76
R92 VNB.n1105 VNB.n1104 76
R93 VNB.n1101 VNB.n1100 76
R94 VNB.n1079 VNB.n1078 76
R95 VNB.n1075 VNB.n1074 76
R96 VNB.n1071 VNB.n1070 76
R97 VNB.n1065 VNB.n1064 76
R98 VNB.n1061 VNB.n1060 76
R99 VNB.n1057 VNB.n1056 76
R100 VNB.n1053 VNB.n1052 76
R101 VNB.n1049 VNB.n1048 76
R102 VNB.n1027 VNB.n1026 76
R103 VNB.n1023 VNB.n1022 76
R104 VNB.n1019 VNB.n1018 76
R105 VNB.n1013 VNB.n1012 76
R106 VNB.n1009 VNB.n1008 76
R107 VNB.n1005 VNB.n1004 76
R108 VNB.n1001 VNB.n1000 76
R109 VNB.n997 VNB.n996 76
R110 VNB.n975 VNB.n974 76
R111 VNB.n971 VNB.n970 76
R112 VNB.n967 VNB.n966 76
R113 VNB.n961 VNB.n960 76
R114 VNB.n957 VNB.n956 76
R115 VNB.n953 VNB.n952 76
R116 VNB.n949 VNB.n948 76
R117 VNB.n945 VNB.n944 76
R118 VNB.n923 VNB.n922 76
R119 VNB.n919 VNB.n918 76
R120 VNB.n915 VNB.n914 76
R121 VNB.n909 VNB.n908 76
R122 VNB.n905 VNB.n904 76
R123 VNB.n901 VNB.n900 76
R124 VNB.n897 VNB.n896 76
R125 VNB.n893 VNB.n892 76
R126 VNB.n871 VNB.n870 76
R127 VNB.n867 VNB.n866 76
R128 VNB.n863 VNB.n862 76
R129 VNB.n857 VNB.n856 76
R130 VNB.n853 VNB.n852 76
R131 VNB.n849 VNB.n848 76
R132 VNB.n845 VNB.n844 76
R133 VNB.n841 VNB.n840 76
R134 VNB.n837 VNB.n836 76
R135 VNB.n833 VNB.n832 76
R136 VNB.n829 VNB.n828 76
R137 VNB.n825 VNB.n824 76
R138 VNB.n803 VNB.n802 76
R139 VNB.n799 VNB.n798 76
R140 VNB.n795 VNB.n794 76
R141 VNB.n789 VNB.n788 76
R142 VNB.n785 VNB.n784 76
R143 VNB.n781 VNB.n780 76
R144 VNB.n777 VNB.n776 76
R145 VNB.n773 VNB.n772 76
R146 VNB.n751 VNB.n750 76
R147 VNB.n747 VNB.n746 76
R148 VNB.n743 VNB.n742 76
R149 VNB.n737 VNB.n736 76
R150 VNB.n733 VNB.n732 76
R151 VNB.n729 VNB.n728 76
R152 VNB.n725 VNB.n724 76
R153 VNB.n721 VNB.n720 76
R154 VNB.n699 VNB.n698 76
R155 VNB.n695 VNB.n694 76
R156 VNB.n691 VNB.n690 76
R157 VNB.n685 VNB.n684 76
R158 VNB.n681 VNB.n680 76
R159 VNB.n677 VNB.n676 76
R160 VNB.n673 VNB.n672 76
R161 VNB.n669 VNB.n668 76
R162 VNB.n647 VNB.n646 76
R163 VNB.n643 VNB.n642 76
R164 VNB.n639 VNB.n636 76
R165 VNB.n625 VNB.n624 76
R166 VNB.n621 VNB.n620 76
R167 VNB.n617 VNB.n616 76
R168 VNB.n595 VNB.n594 76
R169 VNB.n591 VNB.n590 76
R170 VNB.n587 VNB.n586 76
R171 VNB.n581 VNB.n580 76
R172 VNB.n577 VNB.n576 76
R173 VNB.n573 VNB.n572 76
R174 VNB.n569 VNB.n568 76
R175 VNB.n565 VNB.n564 76
R176 VNB.n561 VNB.n560 76
R177 VNB.n557 VNB.n556 76
R178 VNB.n553 VNB.n552 76
R179 VNB.n549 VNB.n548 76
R180 VNB.n527 VNB.n526 76
R181 VNB.n523 VNB.n522 76
R182 VNB.n519 VNB.n518 76
R183 VNB.n513 VNB.n512 76
R184 VNB.n509 VNB.n508 76
R185 VNB.n505 VNB.n504 76
R186 VNB.n501 VNB.n500 76
R187 VNB.n497 VNB.n496 76
R188 VNB.n475 VNB.n474 76
R189 VNB.n471 VNB.n470 76
R190 VNB.n467 VNB.n466 76
R191 VNB.n461 VNB.n460 76
R192 VNB.n457 VNB.n456 76
R193 VNB.n453 VNB.n452 76
R194 VNB.n449 VNB.n448 76
R195 VNB.n445 VNB.n444 76
R196 VNB.n423 VNB.n422 76
R197 VNB.n419 VNB.n418 76
R198 VNB.n415 VNB.n414 76
R199 VNB.n409 VNB.n408 76
R200 VNB.n405 VNB.n404 76
R201 VNB.n401 VNB.n400 76
R202 VNB.n397 VNB.n396 76
R203 VNB.n393 VNB.n392 76
R204 VNB.n371 VNB.n370 76
R205 VNB.n367 VNB.n366 76
R206 VNB.n363 VNB.n362 76
R207 VNB.n357 VNB.n356 76
R208 VNB.n353 VNB.n352 76
R209 VNB.n349 VNB.n348 76
R210 VNB.n345 VNB.n344 76
R211 VNB.n341 VNB.n340 76
R212 VNB.n319 VNB.n318 76
R213 VNB.n315 VNB.n314 76
R214 VNB.n311 VNB.n310 76
R215 VNB.n305 VNB.n304 76
R216 VNB.n301 VNB.n300 76
R217 VNB.n297 VNB.n296 76
R218 VNB.n293 VNB.n292 76
R219 VNB.n289 VNB.n288 76
R220 VNB.n267 VNB.n266 76
R221 VNB.n263 VNB.n262 76
R222 VNB.n259 VNB.n258 76
R223 VNB.n253 VNB.n252 76
R224 VNB.n249 VNB.n248 76
R225 VNB.n245 VNB.n244 76
R226 VNB.n241 VNB.n240 76
R227 VNB.n237 VNB.n236 76
R228 VNB.n215 VNB.n214 76
R229 VNB.n211 VNB.n210 76
R230 VNB.n207 VNB.n206 76
R231 VNB.n201 VNB.n200 76
R232 VNB.n197 VNB.n196 76
R233 VNB.n193 VNB.n192 76
R234 VNB.n189 VNB.n188 76
R235 VNB.n185 VNB.n184 76
R236 VNB.n163 VNB.n162 76
R237 VNB.n159 VNB.n158 76
R238 VNB.n155 VNB.n154 76
R239 VNB.n149 VNB.n148 76
R240 VNB.n86 VNB.n77 63.835
R241 VNB.n585 VNB.n584 41.971
R242 VNB.n861 VNB.n860 41.971
R243 VNB.n51 VNB.n50 41.971
R244 VNB.n83 VNB.n82 36.937
R245 VNB.n153 VNB.n152 36.678
R246 VNB.n205 VNB.n204 36.678
R247 VNB.n257 VNB.n256 36.678
R248 VNB.n309 VNB.n308 36.678
R249 VNB.n361 VNB.n360 36.678
R250 VNB.n413 VNB.n412 36.678
R251 VNB.n465 VNB.n464 36.678
R252 VNB.n517 VNB.n516 36.678
R253 VNB.n638 VNB.n637 36.678
R254 VNB.n689 VNB.n688 36.678
R255 VNB.n741 VNB.n740 36.678
R256 VNB.n793 VNB.n792 36.678
R257 VNB.n913 VNB.n912 36.678
R258 VNB.n965 VNB.n964 36.678
R259 VNB.n1017 VNB.n1016 36.678
R260 VNB.n1069 VNB.n1068 36.678
R261 VNB.n1121 VNB.n1120 36.678
R262 VNB.n144 VNB.n143 35.118
R263 VNB.n77 VNB.n76 28.421
R264 VNB.n89 VNB.n88 27.855
R265 VNB.n77 VNB.n75 25.263
R266 VNB.n75 VNB.n74 24.383
R267 VNB.n133 VNB.n130 20.452
R268 VNB.n1145 VNB.n1144 20.452
R269 VNB.n90 VNB.n89 16.721
R270 VNB.n142 VNB.n141 13.653
R271 VNB.n141 VNB.n140 13.653
R272 VNB.n139 VNB.n138 13.653
R273 VNB.n138 VNB.n137 13.653
R274 VNB.n136 VNB.n135 13.653
R275 VNB.n135 VNB.n134 13.653
R276 VNB.n148 VNB.n147 13.653
R277 VNB.n147 VNB.n146 13.653
R278 VNB.n154 VNB.n153 13.653
R279 VNB.n158 VNB.n157 13.653
R280 VNB.n157 VNB.n156 13.653
R281 VNB.n162 VNB.n161 13.653
R282 VNB.n161 VNB.n160 13.653
R283 VNB.n184 VNB.n183 13.653
R284 VNB.n183 VNB.n182 13.653
R285 VNB.n188 VNB.n187 13.653
R286 VNB.n187 VNB.n186 13.653
R287 VNB.n192 VNB.n191 13.653
R288 VNB.n191 VNB.n190 13.653
R289 VNB.n196 VNB.n195 13.653
R290 VNB.n195 VNB.n194 13.653
R291 VNB.n200 VNB.n199 13.653
R292 VNB.n199 VNB.n198 13.653
R293 VNB.n206 VNB.n205 13.653
R294 VNB.n210 VNB.n209 13.653
R295 VNB.n209 VNB.n208 13.653
R296 VNB.n214 VNB.n213 13.653
R297 VNB.n213 VNB.n212 13.653
R298 VNB.n236 VNB.n235 13.653
R299 VNB.n235 VNB.n234 13.653
R300 VNB.n240 VNB.n239 13.653
R301 VNB.n239 VNB.n238 13.653
R302 VNB.n244 VNB.n243 13.653
R303 VNB.n243 VNB.n242 13.653
R304 VNB.n248 VNB.n247 13.653
R305 VNB.n247 VNB.n246 13.653
R306 VNB.n252 VNB.n251 13.653
R307 VNB.n251 VNB.n250 13.653
R308 VNB.n258 VNB.n257 13.653
R309 VNB.n262 VNB.n261 13.653
R310 VNB.n261 VNB.n260 13.653
R311 VNB.n266 VNB.n265 13.653
R312 VNB.n265 VNB.n264 13.653
R313 VNB.n288 VNB.n287 13.653
R314 VNB.n287 VNB.n286 13.653
R315 VNB.n292 VNB.n291 13.653
R316 VNB.n291 VNB.n290 13.653
R317 VNB.n296 VNB.n295 13.653
R318 VNB.n295 VNB.n294 13.653
R319 VNB.n300 VNB.n299 13.653
R320 VNB.n299 VNB.n298 13.653
R321 VNB.n304 VNB.n303 13.653
R322 VNB.n303 VNB.n302 13.653
R323 VNB.n310 VNB.n309 13.653
R324 VNB.n314 VNB.n313 13.653
R325 VNB.n313 VNB.n312 13.653
R326 VNB.n318 VNB.n317 13.653
R327 VNB.n317 VNB.n316 13.653
R328 VNB.n340 VNB.n339 13.653
R329 VNB.n339 VNB.n338 13.653
R330 VNB.n344 VNB.n343 13.653
R331 VNB.n343 VNB.n342 13.653
R332 VNB.n348 VNB.n347 13.653
R333 VNB.n347 VNB.n346 13.653
R334 VNB.n352 VNB.n351 13.653
R335 VNB.n351 VNB.n350 13.653
R336 VNB.n356 VNB.n355 13.653
R337 VNB.n355 VNB.n354 13.653
R338 VNB.n362 VNB.n361 13.653
R339 VNB.n366 VNB.n365 13.653
R340 VNB.n365 VNB.n364 13.653
R341 VNB.n370 VNB.n369 13.653
R342 VNB.n369 VNB.n368 13.653
R343 VNB.n392 VNB.n391 13.653
R344 VNB.n391 VNB.n390 13.653
R345 VNB.n396 VNB.n395 13.653
R346 VNB.n395 VNB.n394 13.653
R347 VNB.n400 VNB.n399 13.653
R348 VNB.n399 VNB.n398 13.653
R349 VNB.n404 VNB.n403 13.653
R350 VNB.n403 VNB.n402 13.653
R351 VNB.n408 VNB.n407 13.653
R352 VNB.n407 VNB.n406 13.653
R353 VNB.n414 VNB.n413 13.653
R354 VNB.n418 VNB.n417 13.653
R355 VNB.n417 VNB.n416 13.653
R356 VNB.n422 VNB.n421 13.653
R357 VNB.n421 VNB.n420 13.653
R358 VNB.n444 VNB.n443 13.653
R359 VNB.n443 VNB.n442 13.653
R360 VNB.n448 VNB.n447 13.653
R361 VNB.n447 VNB.n446 13.653
R362 VNB.n452 VNB.n451 13.653
R363 VNB.n451 VNB.n450 13.653
R364 VNB.n456 VNB.n455 13.653
R365 VNB.n455 VNB.n454 13.653
R366 VNB.n460 VNB.n459 13.653
R367 VNB.n459 VNB.n458 13.653
R368 VNB.n466 VNB.n465 13.653
R369 VNB.n470 VNB.n469 13.653
R370 VNB.n469 VNB.n468 13.653
R371 VNB.n474 VNB.n473 13.653
R372 VNB.n473 VNB.n472 13.653
R373 VNB.n496 VNB.n495 13.653
R374 VNB.n495 VNB.n494 13.653
R375 VNB.n500 VNB.n499 13.653
R376 VNB.n499 VNB.n498 13.653
R377 VNB.n504 VNB.n503 13.653
R378 VNB.n503 VNB.n502 13.653
R379 VNB.n508 VNB.n507 13.653
R380 VNB.n507 VNB.n506 13.653
R381 VNB.n512 VNB.n511 13.653
R382 VNB.n511 VNB.n510 13.653
R383 VNB.n518 VNB.n517 13.653
R384 VNB.n522 VNB.n521 13.653
R385 VNB.n521 VNB.n520 13.653
R386 VNB.n526 VNB.n525 13.653
R387 VNB.n525 VNB.n524 13.653
R388 VNB.n548 VNB.n547 13.653
R389 VNB.n547 VNB.n546 13.653
R390 VNB.n552 VNB.n551 13.653
R391 VNB.n551 VNB.n550 13.653
R392 VNB.n556 VNB.n555 13.653
R393 VNB.n555 VNB.n554 13.653
R394 VNB.n560 VNB.n559 13.653
R395 VNB.n559 VNB.n558 13.653
R396 VNB.n564 VNB.n563 13.653
R397 VNB.n563 VNB.n562 13.653
R398 VNB.n568 VNB.n567 13.653
R399 VNB.n567 VNB.n566 13.653
R400 VNB.n572 VNB.n571 13.653
R401 VNB.n571 VNB.n570 13.653
R402 VNB.n576 VNB.n575 13.653
R403 VNB.n575 VNB.n574 13.653
R404 VNB.n580 VNB.n579 13.653
R405 VNB.n579 VNB.n578 13.653
R406 VNB.n586 VNB.n585 13.653
R407 VNB.n590 VNB.n589 13.653
R408 VNB.n589 VNB.n588 13.653
R409 VNB.n594 VNB.n593 13.653
R410 VNB.n593 VNB.n592 13.653
R411 VNB.n616 VNB.n615 13.653
R412 VNB.n615 VNB.n614 13.653
R413 VNB.n620 VNB.n619 13.653
R414 VNB.n619 VNB.n618 13.653
R415 VNB.n624 VNB.n623 13.653
R416 VNB.n623 VNB.n622 13.653
R417 VNB.n80 VNB.n79 13.653
R418 VNB.n79 VNB.n78 13.653
R419 VNB.n85 VNB.n84 13.653
R420 VNB.n84 VNB.n83 13.653
R421 VNB.n91 VNB.n90 13.653
R422 VNB.n94 VNB.n93 13.653
R423 VNB.n93 VNB.n92 13.653
R424 VNB.n97 VNB.n96 13.653
R425 VNB.n96 VNB.n95 13.653
R426 VNB.n102 VNB.n101 13.653
R427 VNB.n101 VNB.n100 13.653
R428 VNB.n105 VNB.n104 13.653
R429 VNB.n104 VNB.n103 13.653
R430 VNB.n108 VNB.n107 13.653
R431 VNB.n107 VNB.n106 13.653
R432 VNB.n111 VNB.n110 13.653
R433 VNB.n110 VNB.n109 13.653
R434 VNB.n114 VNB.n113 13.653
R435 VNB.n113 VNB.n112 13.653
R436 VNB.n639 VNB.n638 13.653
R437 VNB.n642 VNB.n641 13.653
R438 VNB.n641 VNB.n640 13.653
R439 VNB.n646 VNB.n645 13.653
R440 VNB.n645 VNB.n644 13.653
R441 VNB.n668 VNB.n667 13.653
R442 VNB.n667 VNB.n666 13.653
R443 VNB.n672 VNB.n671 13.653
R444 VNB.n671 VNB.n670 13.653
R445 VNB.n676 VNB.n675 13.653
R446 VNB.n675 VNB.n674 13.653
R447 VNB.n680 VNB.n679 13.653
R448 VNB.n679 VNB.n678 13.653
R449 VNB.n684 VNB.n683 13.653
R450 VNB.n683 VNB.n682 13.653
R451 VNB.n690 VNB.n689 13.653
R452 VNB.n694 VNB.n693 13.653
R453 VNB.n693 VNB.n692 13.653
R454 VNB.n698 VNB.n697 13.653
R455 VNB.n697 VNB.n696 13.653
R456 VNB.n720 VNB.n719 13.653
R457 VNB.n719 VNB.n718 13.653
R458 VNB.n724 VNB.n723 13.653
R459 VNB.n723 VNB.n722 13.653
R460 VNB.n728 VNB.n727 13.653
R461 VNB.n727 VNB.n726 13.653
R462 VNB.n732 VNB.n731 13.653
R463 VNB.n731 VNB.n730 13.653
R464 VNB.n736 VNB.n735 13.653
R465 VNB.n735 VNB.n734 13.653
R466 VNB.n742 VNB.n741 13.653
R467 VNB.n746 VNB.n745 13.653
R468 VNB.n745 VNB.n744 13.653
R469 VNB.n750 VNB.n749 13.653
R470 VNB.n749 VNB.n748 13.653
R471 VNB.n772 VNB.n771 13.653
R472 VNB.n771 VNB.n770 13.653
R473 VNB.n776 VNB.n775 13.653
R474 VNB.n775 VNB.n774 13.653
R475 VNB.n780 VNB.n779 13.653
R476 VNB.n779 VNB.n778 13.653
R477 VNB.n784 VNB.n783 13.653
R478 VNB.n783 VNB.n782 13.653
R479 VNB.n788 VNB.n787 13.653
R480 VNB.n787 VNB.n786 13.653
R481 VNB.n794 VNB.n793 13.653
R482 VNB.n798 VNB.n797 13.653
R483 VNB.n797 VNB.n796 13.653
R484 VNB.n802 VNB.n801 13.653
R485 VNB.n801 VNB.n800 13.653
R486 VNB.n824 VNB.n823 13.653
R487 VNB.n823 VNB.n822 13.653
R488 VNB.n828 VNB.n827 13.653
R489 VNB.n827 VNB.n826 13.653
R490 VNB.n832 VNB.n831 13.653
R491 VNB.n831 VNB.n830 13.653
R492 VNB.n836 VNB.n835 13.653
R493 VNB.n835 VNB.n834 13.653
R494 VNB.n840 VNB.n839 13.653
R495 VNB.n839 VNB.n838 13.653
R496 VNB.n844 VNB.n843 13.653
R497 VNB.n843 VNB.n842 13.653
R498 VNB.n848 VNB.n847 13.653
R499 VNB.n847 VNB.n846 13.653
R500 VNB.n852 VNB.n851 13.653
R501 VNB.n851 VNB.n850 13.653
R502 VNB.n856 VNB.n855 13.653
R503 VNB.n855 VNB.n854 13.653
R504 VNB.n862 VNB.n861 13.653
R505 VNB.n866 VNB.n865 13.653
R506 VNB.n865 VNB.n864 13.653
R507 VNB.n870 VNB.n869 13.653
R508 VNB.n869 VNB.n868 13.653
R509 VNB.n892 VNB.n891 13.653
R510 VNB.n891 VNB.n890 13.653
R511 VNB.n896 VNB.n895 13.653
R512 VNB.n895 VNB.n894 13.653
R513 VNB.n900 VNB.n899 13.653
R514 VNB.n899 VNB.n898 13.653
R515 VNB.n904 VNB.n903 13.653
R516 VNB.n903 VNB.n902 13.653
R517 VNB.n908 VNB.n907 13.653
R518 VNB.n907 VNB.n906 13.653
R519 VNB.n914 VNB.n913 13.653
R520 VNB.n918 VNB.n917 13.653
R521 VNB.n917 VNB.n916 13.653
R522 VNB.n922 VNB.n921 13.653
R523 VNB.n921 VNB.n920 13.653
R524 VNB.n944 VNB.n943 13.653
R525 VNB.n943 VNB.n942 13.653
R526 VNB.n948 VNB.n947 13.653
R527 VNB.n947 VNB.n946 13.653
R528 VNB.n952 VNB.n951 13.653
R529 VNB.n951 VNB.n950 13.653
R530 VNB.n956 VNB.n955 13.653
R531 VNB.n955 VNB.n954 13.653
R532 VNB.n960 VNB.n959 13.653
R533 VNB.n959 VNB.n958 13.653
R534 VNB.n966 VNB.n965 13.653
R535 VNB.n970 VNB.n969 13.653
R536 VNB.n969 VNB.n968 13.653
R537 VNB.n974 VNB.n973 13.653
R538 VNB.n973 VNB.n972 13.653
R539 VNB.n996 VNB.n995 13.653
R540 VNB.n995 VNB.n994 13.653
R541 VNB.n1000 VNB.n999 13.653
R542 VNB.n999 VNB.n998 13.653
R543 VNB.n1004 VNB.n1003 13.653
R544 VNB.n1003 VNB.n1002 13.653
R545 VNB.n1008 VNB.n1007 13.653
R546 VNB.n1007 VNB.n1006 13.653
R547 VNB.n1012 VNB.n1011 13.653
R548 VNB.n1011 VNB.n1010 13.653
R549 VNB.n1018 VNB.n1017 13.653
R550 VNB.n1022 VNB.n1021 13.653
R551 VNB.n1021 VNB.n1020 13.653
R552 VNB.n1026 VNB.n1025 13.653
R553 VNB.n1025 VNB.n1024 13.653
R554 VNB.n1048 VNB.n1047 13.653
R555 VNB.n1047 VNB.n1046 13.653
R556 VNB.n1052 VNB.n1051 13.653
R557 VNB.n1051 VNB.n1050 13.653
R558 VNB.n1056 VNB.n1055 13.653
R559 VNB.n1055 VNB.n1054 13.653
R560 VNB.n1060 VNB.n1059 13.653
R561 VNB.n1059 VNB.n1058 13.653
R562 VNB.n1064 VNB.n1063 13.653
R563 VNB.n1063 VNB.n1062 13.653
R564 VNB.n1070 VNB.n1069 13.653
R565 VNB.n1074 VNB.n1073 13.653
R566 VNB.n1073 VNB.n1072 13.653
R567 VNB.n1078 VNB.n1077 13.653
R568 VNB.n1077 VNB.n1076 13.653
R569 VNB.n1100 VNB.n1099 13.653
R570 VNB.n1099 VNB.n1098 13.653
R571 VNB.n1104 VNB.n1103 13.653
R572 VNB.n1103 VNB.n1102 13.653
R573 VNB.n1108 VNB.n1107 13.653
R574 VNB.n1107 VNB.n1106 13.653
R575 VNB.n1112 VNB.n1111 13.653
R576 VNB.n1111 VNB.n1110 13.653
R577 VNB.n1116 VNB.n1115 13.653
R578 VNB.n1115 VNB.n1114 13.653
R579 VNB.n1122 VNB.n1121 13.653
R580 VNB.n1126 VNB.n1125 13.653
R581 VNB.n1125 VNB.n1124 13.653
R582 VNB.n1130 VNB.n1129 13.653
R583 VNB.n1129 VNB.n1128 13.653
R584 VNB.n25 VNB.n24 13.653
R585 VNB.n24 VNB.n23 13.653
R586 VNB.n28 VNB.n27 13.653
R587 VNB.n27 VNB.n26 13.653
R588 VNB.n31 VNB.n30 13.653
R589 VNB.n30 VNB.n29 13.653
R590 VNB.n34 VNB.n33 13.653
R591 VNB.n33 VNB.n32 13.653
R592 VNB.n37 VNB.n36 13.653
R593 VNB.n36 VNB.n35 13.653
R594 VNB.n40 VNB.n39 13.653
R595 VNB.n39 VNB.n38 13.653
R596 VNB.n43 VNB.n42 13.653
R597 VNB.n42 VNB.n41 13.653
R598 VNB.n46 VNB.n45 13.653
R599 VNB.n45 VNB.n44 13.653
R600 VNB.n49 VNB.n48 13.653
R601 VNB.n48 VNB.n47 13.653
R602 VNB.n52 VNB.n51 13.653
R603 VNB.n56 VNB.n55 13.653
R604 VNB.n55 VNB.n54 13.653
R605 VNB.n1144 VNB.n0 13.653
R606 VNB VNB.n0 13.653
R607 VNB.n133 VNB.n132 13.653
R608 VNB.n132 VNB.n131 13.653
R609 VNB.n1152 VNB.n1149 13.577
R610 VNB.n118 VNB.n116 13.276
R611 VNB.n130 VNB.n118 13.276
R612 VNB.n166 VNB.n164 13.276
R613 VNB.n179 VNB.n166 13.276
R614 VNB.n218 VNB.n216 13.276
R615 VNB.n231 VNB.n218 13.276
R616 VNB.n270 VNB.n268 13.276
R617 VNB.n283 VNB.n270 13.276
R618 VNB.n322 VNB.n320 13.276
R619 VNB.n335 VNB.n322 13.276
R620 VNB.n374 VNB.n372 13.276
R621 VNB.n387 VNB.n374 13.276
R622 VNB.n426 VNB.n424 13.276
R623 VNB.n439 VNB.n426 13.276
R624 VNB.n478 VNB.n476 13.276
R625 VNB.n491 VNB.n478 13.276
R626 VNB.n530 VNB.n528 13.276
R627 VNB.n543 VNB.n530 13.276
R628 VNB.n598 VNB.n596 13.276
R629 VNB.n611 VNB.n598 13.276
R630 VNB.n60 VNB.n58 13.276
R631 VNB.n73 VNB.n60 13.276
R632 VNB.n650 VNB.n648 13.276
R633 VNB.n663 VNB.n650 13.276
R634 VNB.n702 VNB.n700 13.276
R635 VNB.n715 VNB.n702 13.276
R636 VNB.n754 VNB.n752 13.276
R637 VNB.n767 VNB.n754 13.276
R638 VNB.n806 VNB.n804 13.276
R639 VNB.n819 VNB.n806 13.276
R640 VNB.n874 VNB.n872 13.276
R641 VNB.n887 VNB.n874 13.276
R642 VNB.n926 VNB.n924 13.276
R643 VNB.n939 VNB.n926 13.276
R644 VNB.n978 VNB.n976 13.276
R645 VNB.n991 VNB.n978 13.276
R646 VNB.n1030 VNB.n1028 13.276
R647 VNB.n1043 VNB.n1030 13.276
R648 VNB.n1082 VNB.n1080 13.276
R649 VNB.n1095 VNB.n1082 13.276
R650 VNB.n7 VNB.n5 13.276
R651 VNB.n20 VNB.n7 13.276
R652 VNB.n142 VNB.n139 13.276
R653 VNB.n139 VNB.n136 13.276
R654 VNB.n184 VNB.n180 13.276
R655 VNB.n236 VNB.n232 13.276
R656 VNB.n288 VNB.n284 13.276
R657 VNB.n340 VNB.n336 13.276
R658 VNB.n392 VNB.n388 13.276
R659 VNB.n444 VNB.n440 13.276
R660 VNB.n496 VNB.n492 13.276
R661 VNB.n548 VNB.n544 13.276
R662 VNB.n616 VNB.n612 13.276
R663 VNB.n85 VNB.n80 13.276
R664 VNB.n94 VNB.n91 13.276
R665 VNB.n97 VNB.n94 13.276
R666 VNB.n98 VNB.n97 13.276
R667 VNB.n102 VNB.n98 13.276
R668 VNB.n105 VNB.n102 13.276
R669 VNB.n108 VNB.n105 13.276
R670 VNB.n111 VNB.n108 13.276
R671 VNB.n114 VNB.n111 13.276
R672 VNB.n642 VNB.n639 13.276
R673 VNB.n668 VNB.n664 13.276
R674 VNB.n720 VNB.n716 13.276
R675 VNB.n772 VNB.n768 13.276
R676 VNB.n824 VNB.n820 13.276
R677 VNB.n892 VNB.n888 13.276
R678 VNB.n944 VNB.n940 13.276
R679 VNB.n996 VNB.n992 13.276
R680 VNB.n1048 VNB.n1044 13.276
R681 VNB.n1100 VNB.n1096 13.276
R682 VNB.n25 VNB.n21 13.276
R683 VNB.n28 VNB.n25 13.276
R684 VNB.n31 VNB.n28 13.276
R685 VNB.n34 VNB.n31 13.276
R686 VNB.n37 VNB.n34 13.276
R687 VNB.n40 VNB.n37 13.276
R688 VNB.n43 VNB.n40 13.276
R689 VNB.n46 VNB.n43 13.276
R690 VNB.n49 VNB.n46 13.276
R691 VNB.n52 VNB.n49 13.276
R692 VNB.n1144 VNB.n56 13.276
R693 VNB.n3 VNB.n1 13.276
R694 VNB.n1145 VNB.n3 13.276
R695 VNB.n56 VNB.n53 12.02
R696 VNB.n86 VNB.n85 10.764
R697 VNB.n115 VNB.n114 10.764
R698 VNB.n1154 VNB.n1153 7.5
R699 VNB.n172 VNB.n171 7.5
R700 VNB.n168 VNB.n167 7.5
R701 VNB.n166 VNB.n165 7.5
R702 VNB.n179 VNB.n178 7.5
R703 VNB.n224 VNB.n223 7.5
R704 VNB.n220 VNB.n219 7.5
R705 VNB.n218 VNB.n217 7.5
R706 VNB.n231 VNB.n230 7.5
R707 VNB.n276 VNB.n275 7.5
R708 VNB.n272 VNB.n271 7.5
R709 VNB.n270 VNB.n269 7.5
R710 VNB.n283 VNB.n282 7.5
R711 VNB.n328 VNB.n327 7.5
R712 VNB.n324 VNB.n323 7.5
R713 VNB.n322 VNB.n321 7.5
R714 VNB.n335 VNB.n334 7.5
R715 VNB.n380 VNB.n379 7.5
R716 VNB.n376 VNB.n375 7.5
R717 VNB.n374 VNB.n373 7.5
R718 VNB.n387 VNB.n386 7.5
R719 VNB.n432 VNB.n431 7.5
R720 VNB.n428 VNB.n427 7.5
R721 VNB.n426 VNB.n425 7.5
R722 VNB.n439 VNB.n438 7.5
R723 VNB.n484 VNB.n483 7.5
R724 VNB.n480 VNB.n479 7.5
R725 VNB.n478 VNB.n477 7.5
R726 VNB.n491 VNB.n490 7.5
R727 VNB.n536 VNB.n535 7.5
R728 VNB.n532 VNB.n531 7.5
R729 VNB.n530 VNB.n529 7.5
R730 VNB.n543 VNB.n542 7.5
R731 VNB.n604 VNB.n603 7.5
R732 VNB.n600 VNB.n599 7.5
R733 VNB.n598 VNB.n597 7.5
R734 VNB.n611 VNB.n610 7.5
R735 VNB.n66 VNB.n65 7.5
R736 VNB.n62 VNB.n61 7.5
R737 VNB.n60 VNB.n59 7.5
R738 VNB.n73 VNB.n72 7.5
R739 VNB.n656 VNB.n655 7.5
R740 VNB.n652 VNB.n651 7.5
R741 VNB.n650 VNB.n649 7.5
R742 VNB.n663 VNB.n662 7.5
R743 VNB.n708 VNB.n707 7.5
R744 VNB.n704 VNB.n703 7.5
R745 VNB.n702 VNB.n701 7.5
R746 VNB.n715 VNB.n714 7.5
R747 VNB.n760 VNB.n759 7.5
R748 VNB.n756 VNB.n755 7.5
R749 VNB.n754 VNB.n753 7.5
R750 VNB.n767 VNB.n766 7.5
R751 VNB.n812 VNB.n811 7.5
R752 VNB.n808 VNB.n807 7.5
R753 VNB.n806 VNB.n805 7.5
R754 VNB.n819 VNB.n818 7.5
R755 VNB.n880 VNB.n879 7.5
R756 VNB.n876 VNB.n875 7.5
R757 VNB.n874 VNB.n873 7.5
R758 VNB.n887 VNB.n886 7.5
R759 VNB.n932 VNB.n931 7.5
R760 VNB.n928 VNB.n927 7.5
R761 VNB.n926 VNB.n925 7.5
R762 VNB.n939 VNB.n938 7.5
R763 VNB.n984 VNB.n983 7.5
R764 VNB.n980 VNB.n979 7.5
R765 VNB.n978 VNB.n977 7.5
R766 VNB.n991 VNB.n990 7.5
R767 VNB.n1036 VNB.n1035 7.5
R768 VNB.n1032 VNB.n1031 7.5
R769 VNB.n1030 VNB.n1029 7.5
R770 VNB.n1043 VNB.n1042 7.5
R771 VNB.n1088 VNB.n1087 7.5
R772 VNB.n1084 VNB.n1083 7.5
R773 VNB.n1082 VNB.n1081 7.5
R774 VNB.n1095 VNB.n1094 7.5
R775 VNB.n13 VNB.n12 7.5
R776 VNB.n9 VNB.n8 7.5
R777 VNB.n7 VNB.n6 7.5
R778 VNB.n20 VNB.n19 7.5
R779 VNB.n1146 VNB.n1145 7.5
R780 VNB.n3 VNB.n2 7.5
R781 VNB.n1151 VNB.n1150 7.5
R782 VNB.n124 VNB.n123 7.5
R783 VNB.n120 VNB.n119 7.5
R784 VNB.n118 VNB.n117 7.5
R785 VNB.n130 VNB.n129 7.5
R786 VNB.n180 VNB.n179 7.176
R787 VNB.n232 VNB.n231 7.176
R788 VNB.n284 VNB.n283 7.176
R789 VNB.n336 VNB.n335 7.176
R790 VNB.n388 VNB.n387 7.176
R791 VNB.n440 VNB.n439 7.176
R792 VNB.n492 VNB.n491 7.176
R793 VNB.n544 VNB.n543 7.176
R794 VNB.n612 VNB.n611 7.176
R795 VNB.n98 VNB.n73 7.176
R796 VNB.n664 VNB.n663 7.176
R797 VNB.n716 VNB.n715 7.176
R798 VNB.n768 VNB.n767 7.176
R799 VNB.n820 VNB.n819 7.176
R800 VNB.n888 VNB.n887 7.176
R801 VNB.n940 VNB.n939 7.176
R802 VNB.n992 VNB.n991 7.176
R803 VNB.n1044 VNB.n1043 7.176
R804 VNB.n1096 VNB.n1095 7.176
R805 VNB.n21 VNB.n20 7.176
R806 VNB.n1156 VNB.n1154 7.011
R807 VNB.n175 VNB.n172 7.011
R808 VNB.n170 VNB.n168 7.011
R809 VNB.n227 VNB.n224 7.011
R810 VNB.n222 VNB.n220 7.011
R811 VNB.n279 VNB.n276 7.011
R812 VNB.n274 VNB.n272 7.011
R813 VNB.n331 VNB.n328 7.011
R814 VNB.n326 VNB.n324 7.011
R815 VNB.n383 VNB.n380 7.011
R816 VNB.n378 VNB.n376 7.011
R817 VNB.n435 VNB.n432 7.011
R818 VNB.n430 VNB.n428 7.011
R819 VNB.n487 VNB.n484 7.011
R820 VNB.n482 VNB.n480 7.011
R821 VNB.n539 VNB.n536 7.011
R822 VNB.n534 VNB.n532 7.011
R823 VNB.n607 VNB.n604 7.011
R824 VNB.n602 VNB.n600 7.011
R825 VNB.n69 VNB.n66 7.011
R826 VNB.n64 VNB.n62 7.011
R827 VNB.n659 VNB.n656 7.011
R828 VNB.n654 VNB.n652 7.011
R829 VNB.n711 VNB.n708 7.011
R830 VNB.n706 VNB.n704 7.011
R831 VNB.n763 VNB.n760 7.011
R832 VNB.n758 VNB.n756 7.011
R833 VNB.n815 VNB.n812 7.011
R834 VNB.n810 VNB.n808 7.011
R835 VNB.n883 VNB.n880 7.011
R836 VNB.n878 VNB.n876 7.011
R837 VNB.n935 VNB.n932 7.011
R838 VNB.n930 VNB.n928 7.011
R839 VNB.n987 VNB.n984 7.011
R840 VNB.n982 VNB.n980 7.011
R841 VNB.n1039 VNB.n1036 7.011
R842 VNB.n1034 VNB.n1032 7.011
R843 VNB.n1091 VNB.n1088 7.011
R844 VNB.n1086 VNB.n1084 7.011
R845 VNB.n16 VNB.n13 7.011
R846 VNB.n11 VNB.n9 7.011
R847 VNB.n126 VNB.n124 7.011
R848 VNB.n122 VNB.n120 7.011
R849 VNB.n178 VNB.n177 7.01
R850 VNB.n170 VNB.n169 7.01
R851 VNB.n175 VNB.n174 7.01
R852 VNB.n230 VNB.n229 7.01
R853 VNB.n222 VNB.n221 7.01
R854 VNB.n227 VNB.n226 7.01
R855 VNB.n282 VNB.n281 7.01
R856 VNB.n274 VNB.n273 7.01
R857 VNB.n279 VNB.n278 7.01
R858 VNB.n334 VNB.n333 7.01
R859 VNB.n326 VNB.n325 7.01
R860 VNB.n331 VNB.n330 7.01
R861 VNB.n386 VNB.n385 7.01
R862 VNB.n378 VNB.n377 7.01
R863 VNB.n383 VNB.n382 7.01
R864 VNB.n438 VNB.n437 7.01
R865 VNB.n430 VNB.n429 7.01
R866 VNB.n435 VNB.n434 7.01
R867 VNB.n490 VNB.n489 7.01
R868 VNB.n482 VNB.n481 7.01
R869 VNB.n487 VNB.n486 7.01
R870 VNB.n542 VNB.n541 7.01
R871 VNB.n534 VNB.n533 7.01
R872 VNB.n539 VNB.n538 7.01
R873 VNB.n610 VNB.n609 7.01
R874 VNB.n602 VNB.n601 7.01
R875 VNB.n607 VNB.n606 7.01
R876 VNB.n72 VNB.n71 7.01
R877 VNB.n64 VNB.n63 7.01
R878 VNB.n69 VNB.n68 7.01
R879 VNB.n662 VNB.n661 7.01
R880 VNB.n654 VNB.n653 7.01
R881 VNB.n659 VNB.n658 7.01
R882 VNB.n714 VNB.n713 7.01
R883 VNB.n706 VNB.n705 7.01
R884 VNB.n711 VNB.n710 7.01
R885 VNB.n766 VNB.n765 7.01
R886 VNB.n758 VNB.n757 7.01
R887 VNB.n763 VNB.n762 7.01
R888 VNB.n818 VNB.n817 7.01
R889 VNB.n810 VNB.n809 7.01
R890 VNB.n815 VNB.n814 7.01
R891 VNB.n886 VNB.n885 7.01
R892 VNB.n878 VNB.n877 7.01
R893 VNB.n883 VNB.n882 7.01
R894 VNB.n938 VNB.n937 7.01
R895 VNB.n930 VNB.n929 7.01
R896 VNB.n935 VNB.n934 7.01
R897 VNB.n990 VNB.n989 7.01
R898 VNB.n982 VNB.n981 7.01
R899 VNB.n987 VNB.n986 7.01
R900 VNB.n1042 VNB.n1041 7.01
R901 VNB.n1034 VNB.n1033 7.01
R902 VNB.n1039 VNB.n1038 7.01
R903 VNB.n1094 VNB.n1093 7.01
R904 VNB.n1086 VNB.n1085 7.01
R905 VNB.n1091 VNB.n1090 7.01
R906 VNB.n19 VNB.n18 7.01
R907 VNB.n11 VNB.n10 7.01
R908 VNB.n16 VNB.n15 7.01
R909 VNB.n129 VNB.n128 7.01
R910 VNB.n122 VNB.n121 7.01
R911 VNB.n126 VNB.n125 7.01
R912 VNB.n1156 VNB.n1155 7.01
R913 VNB.n1152 VNB.n1151 6.788
R914 VNB.n1147 VNB.n1146 6.788
R915 VNB.n143 VNB.n133 6.111
R916 VNB.n143 VNB.n142 6.1
R917 VNB.n154 VNB.n151 2.511
R918 VNB.n206 VNB.n203 2.511
R919 VNB.n258 VNB.n255 2.511
R920 VNB.n310 VNB.n307 2.511
R921 VNB.n362 VNB.n359 2.511
R922 VNB.n414 VNB.n411 2.511
R923 VNB.n466 VNB.n463 2.511
R924 VNB.n518 VNB.n515 2.511
R925 VNB.n91 VNB.n86 2.511
R926 VNB.n639 VNB.n115 2.511
R927 VNB.n690 VNB.n687 2.511
R928 VNB.n742 VNB.n739 2.511
R929 VNB.n794 VNB.n791 2.511
R930 VNB.n914 VNB.n911 2.511
R931 VNB.n966 VNB.n963 2.511
R932 VNB.n1018 VNB.n1015 2.511
R933 VNB.n1070 VNB.n1067 2.511
R934 VNB.n1122 VNB.n1119 2.511
R935 VNB.n89 VNB.n87 1.99
R936 VNB.n586 VNB.n583 1.255
R937 VNB.n862 VNB.n859 1.255
R938 VNB.n53 VNB.n52 1.255
R939 VNB.n1157 VNB.n1148 0.921
R940 VNB.n1157 VNB.n1152 0.476
R941 VNB.n1157 VNB.n1147 0.475
R942 VNB.n185 VNB.n163 0.272
R943 VNB.n237 VNB.n215 0.272
R944 VNB.n289 VNB.n267 0.272
R945 VNB.n341 VNB.n319 0.272
R946 VNB.n393 VNB.n371 0.272
R947 VNB.n445 VNB.n423 0.272
R948 VNB.n497 VNB.n475 0.272
R949 VNB.n549 VNB.n527 0.272
R950 VNB.n617 VNB.n595 0.272
R951 VNB.n631 VNB.n630 0.272
R952 VNB.n669 VNB.n647 0.272
R953 VNB.n721 VNB.n699 0.272
R954 VNB.n773 VNB.n751 0.272
R955 VNB.n825 VNB.n803 0.272
R956 VNB.n893 VNB.n871 0.272
R957 VNB.n945 VNB.n923 0.272
R958 VNB.n997 VNB.n975 0.272
R959 VNB.n1049 VNB.n1027 0.272
R960 VNB.n1101 VNB.n1079 0.272
R961 VNB.n1132 VNB.n1131 0.272
R962 VNB.n176 VNB.n170 0.246
R963 VNB.n177 VNB.n176 0.246
R964 VNB.n176 VNB.n175 0.246
R965 VNB.n228 VNB.n222 0.246
R966 VNB.n229 VNB.n228 0.246
R967 VNB.n228 VNB.n227 0.246
R968 VNB.n280 VNB.n274 0.246
R969 VNB.n281 VNB.n280 0.246
R970 VNB.n280 VNB.n279 0.246
R971 VNB.n332 VNB.n326 0.246
R972 VNB.n333 VNB.n332 0.246
R973 VNB.n332 VNB.n331 0.246
R974 VNB.n384 VNB.n378 0.246
R975 VNB.n385 VNB.n384 0.246
R976 VNB.n384 VNB.n383 0.246
R977 VNB.n436 VNB.n430 0.246
R978 VNB.n437 VNB.n436 0.246
R979 VNB.n436 VNB.n435 0.246
R980 VNB.n488 VNB.n482 0.246
R981 VNB.n489 VNB.n488 0.246
R982 VNB.n488 VNB.n487 0.246
R983 VNB.n540 VNB.n534 0.246
R984 VNB.n541 VNB.n540 0.246
R985 VNB.n540 VNB.n539 0.246
R986 VNB.n608 VNB.n602 0.246
R987 VNB.n609 VNB.n608 0.246
R988 VNB.n608 VNB.n607 0.246
R989 VNB.n70 VNB.n64 0.246
R990 VNB.n71 VNB.n70 0.246
R991 VNB.n70 VNB.n69 0.246
R992 VNB.n660 VNB.n654 0.246
R993 VNB.n661 VNB.n660 0.246
R994 VNB.n660 VNB.n659 0.246
R995 VNB.n712 VNB.n706 0.246
R996 VNB.n713 VNB.n712 0.246
R997 VNB.n712 VNB.n711 0.246
R998 VNB.n764 VNB.n758 0.246
R999 VNB.n765 VNB.n764 0.246
R1000 VNB.n764 VNB.n763 0.246
R1001 VNB.n816 VNB.n810 0.246
R1002 VNB.n817 VNB.n816 0.246
R1003 VNB.n816 VNB.n815 0.246
R1004 VNB.n884 VNB.n878 0.246
R1005 VNB.n885 VNB.n884 0.246
R1006 VNB.n884 VNB.n883 0.246
R1007 VNB.n936 VNB.n930 0.246
R1008 VNB.n937 VNB.n936 0.246
R1009 VNB.n936 VNB.n935 0.246
R1010 VNB.n988 VNB.n982 0.246
R1011 VNB.n989 VNB.n988 0.246
R1012 VNB.n988 VNB.n987 0.246
R1013 VNB.n1040 VNB.n1034 0.246
R1014 VNB.n1041 VNB.n1040 0.246
R1015 VNB.n1040 VNB.n1039 0.246
R1016 VNB.n1092 VNB.n1086 0.246
R1017 VNB.n1093 VNB.n1092 0.246
R1018 VNB.n1092 VNB.n1091 0.246
R1019 VNB.n17 VNB.n11 0.246
R1020 VNB.n18 VNB.n17 0.246
R1021 VNB.n17 VNB.n16 0.246
R1022 VNB.n127 VNB.n122 0.246
R1023 VNB.n128 VNB.n127 0.246
R1024 VNB.n127 VNB.n126 0.246
R1025 VNB.n1157 VNB.n1156 0.246
R1026 VNB.n1143 VNB 0.198
R1027 VNB.n145 VNB.n144 0.136
R1028 VNB.n149 VNB.n145 0.136
R1029 VNB.n155 VNB.n149 0.136
R1030 VNB.n159 VNB.n155 0.136
R1031 VNB.n163 VNB.n159 0.136
R1032 VNB.n189 VNB.n185 0.136
R1033 VNB.n193 VNB.n189 0.136
R1034 VNB.n197 VNB.n193 0.136
R1035 VNB.n201 VNB.n197 0.136
R1036 VNB.n207 VNB.n201 0.136
R1037 VNB.n211 VNB.n207 0.136
R1038 VNB.n215 VNB.n211 0.136
R1039 VNB.n241 VNB.n237 0.136
R1040 VNB.n245 VNB.n241 0.136
R1041 VNB.n249 VNB.n245 0.136
R1042 VNB.n253 VNB.n249 0.136
R1043 VNB.n259 VNB.n253 0.136
R1044 VNB.n263 VNB.n259 0.136
R1045 VNB.n267 VNB.n263 0.136
R1046 VNB.n293 VNB.n289 0.136
R1047 VNB.n297 VNB.n293 0.136
R1048 VNB.n301 VNB.n297 0.136
R1049 VNB.n305 VNB.n301 0.136
R1050 VNB.n311 VNB.n305 0.136
R1051 VNB.n315 VNB.n311 0.136
R1052 VNB.n319 VNB.n315 0.136
R1053 VNB.n345 VNB.n341 0.136
R1054 VNB.n349 VNB.n345 0.136
R1055 VNB.n353 VNB.n349 0.136
R1056 VNB.n357 VNB.n353 0.136
R1057 VNB.n363 VNB.n357 0.136
R1058 VNB.n367 VNB.n363 0.136
R1059 VNB.n371 VNB.n367 0.136
R1060 VNB.n397 VNB.n393 0.136
R1061 VNB.n401 VNB.n397 0.136
R1062 VNB.n405 VNB.n401 0.136
R1063 VNB.n409 VNB.n405 0.136
R1064 VNB.n415 VNB.n409 0.136
R1065 VNB.n419 VNB.n415 0.136
R1066 VNB.n423 VNB.n419 0.136
R1067 VNB.n449 VNB.n445 0.136
R1068 VNB.n453 VNB.n449 0.136
R1069 VNB.n457 VNB.n453 0.136
R1070 VNB.n461 VNB.n457 0.136
R1071 VNB.n467 VNB.n461 0.136
R1072 VNB.n471 VNB.n467 0.136
R1073 VNB.n475 VNB.n471 0.136
R1074 VNB.n501 VNB.n497 0.136
R1075 VNB.n505 VNB.n501 0.136
R1076 VNB.n509 VNB.n505 0.136
R1077 VNB.n513 VNB.n509 0.136
R1078 VNB.n519 VNB.n513 0.136
R1079 VNB.n523 VNB.n519 0.136
R1080 VNB.n527 VNB.n523 0.136
R1081 VNB.n553 VNB.n549 0.136
R1082 VNB.n557 VNB.n553 0.136
R1083 VNB.n561 VNB.n557 0.136
R1084 VNB.n565 VNB.n561 0.136
R1085 VNB.n569 VNB.n565 0.136
R1086 VNB.n573 VNB.n569 0.136
R1087 VNB.n577 VNB.n573 0.136
R1088 VNB.n581 VNB.n577 0.136
R1089 VNB.n587 VNB.n581 0.136
R1090 VNB.n591 VNB.n587 0.136
R1091 VNB.n595 VNB.n591 0.136
R1092 VNB.n621 VNB.n617 0.136
R1093 VNB.n625 VNB.n621 0.136
R1094 VNB.n626 VNB.n625 0.136
R1095 VNB.n627 VNB.n626 0.136
R1096 VNB.n628 VNB.n627 0.136
R1097 VNB.n629 VNB.n628 0.136
R1098 VNB.n630 VNB.n629 0.136
R1099 VNB.n632 VNB.n631 0.136
R1100 VNB.n633 VNB.n632 0.136
R1101 VNB.n634 VNB.n633 0.136
R1102 VNB.n635 VNB.n634 0.136
R1103 VNB.n636 VNB.n635 0.136
R1104 VNB.n647 VNB.n643 0.136
R1105 VNB.n673 VNB.n669 0.136
R1106 VNB.n677 VNB.n673 0.136
R1107 VNB.n681 VNB.n677 0.136
R1108 VNB.n685 VNB.n681 0.136
R1109 VNB.n691 VNB.n685 0.136
R1110 VNB.n695 VNB.n691 0.136
R1111 VNB.n699 VNB.n695 0.136
R1112 VNB.n725 VNB.n721 0.136
R1113 VNB.n729 VNB.n725 0.136
R1114 VNB.n733 VNB.n729 0.136
R1115 VNB.n737 VNB.n733 0.136
R1116 VNB.n743 VNB.n737 0.136
R1117 VNB.n747 VNB.n743 0.136
R1118 VNB.n751 VNB.n747 0.136
R1119 VNB.n777 VNB.n773 0.136
R1120 VNB.n781 VNB.n777 0.136
R1121 VNB.n785 VNB.n781 0.136
R1122 VNB.n789 VNB.n785 0.136
R1123 VNB.n795 VNB.n789 0.136
R1124 VNB.n799 VNB.n795 0.136
R1125 VNB.n803 VNB.n799 0.136
R1126 VNB.n829 VNB.n825 0.136
R1127 VNB.n833 VNB.n829 0.136
R1128 VNB.n837 VNB.n833 0.136
R1129 VNB.n841 VNB.n837 0.136
R1130 VNB.n845 VNB.n841 0.136
R1131 VNB.n849 VNB.n845 0.136
R1132 VNB.n853 VNB.n849 0.136
R1133 VNB.n857 VNB.n853 0.136
R1134 VNB.n863 VNB.n857 0.136
R1135 VNB.n867 VNB.n863 0.136
R1136 VNB.n871 VNB.n867 0.136
R1137 VNB.n897 VNB.n893 0.136
R1138 VNB.n901 VNB.n897 0.136
R1139 VNB.n905 VNB.n901 0.136
R1140 VNB.n909 VNB.n905 0.136
R1141 VNB.n915 VNB.n909 0.136
R1142 VNB.n919 VNB.n915 0.136
R1143 VNB.n923 VNB.n919 0.136
R1144 VNB.n949 VNB.n945 0.136
R1145 VNB.n953 VNB.n949 0.136
R1146 VNB.n957 VNB.n953 0.136
R1147 VNB.n961 VNB.n957 0.136
R1148 VNB.n967 VNB.n961 0.136
R1149 VNB.n971 VNB.n967 0.136
R1150 VNB.n975 VNB.n971 0.136
R1151 VNB.n1001 VNB.n997 0.136
R1152 VNB.n1005 VNB.n1001 0.136
R1153 VNB.n1009 VNB.n1005 0.136
R1154 VNB.n1013 VNB.n1009 0.136
R1155 VNB.n1019 VNB.n1013 0.136
R1156 VNB.n1023 VNB.n1019 0.136
R1157 VNB.n1027 VNB.n1023 0.136
R1158 VNB.n1053 VNB.n1049 0.136
R1159 VNB.n1057 VNB.n1053 0.136
R1160 VNB.n1061 VNB.n1057 0.136
R1161 VNB.n1065 VNB.n1061 0.136
R1162 VNB.n1071 VNB.n1065 0.136
R1163 VNB.n1075 VNB.n1071 0.136
R1164 VNB.n1079 VNB.n1075 0.136
R1165 VNB.n1105 VNB.n1101 0.136
R1166 VNB.n1109 VNB.n1105 0.136
R1167 VNB.n1113 VNB.n1109 0.136
R1168 VNB.n1117 VNB.n1113 0.136
R1169 VNB.n1123 VNB.n1117 0.136
R1170 VNB.n1127 VNB.n1123 0.136
R1171 VNB.n1131 VNB.n1127 0.136
R1172 VNB.n1133 VNB.n1132 0.136
R1173 VNB.n1134 VNB.n1133 0.136
R1174 VNB.n1135 VNB.n1134 0.136
R1175 VNB.n1136 VNB.n1135 0.136
R1176 VNB.n1137 VNB.n1136 0.136
R1177 VNB.n1138 VNB.n1137 0.136
R1178 VNB.n1139 VNB.n1138 0.136
R1179 VNB.n1140 VNB.n1139 0.136
R1180 VNB.n1141 VNB.n1140 0.136
R1181 VNB.n1142 VNB.n1141 0.136
R1182 VNB.n1143 VNB.n1142 0.136
R1183 VNB.n636 VNB 0.068
R1184 VNB.n643 VNB 0.068
R1185 a_4439_159.n8 a_4439_159.t8 512.525
R1186 a_4439_159.n6 a_4439_159.t13 472.359
R1187 a_4439_159.n4 a_4439_159.t6 472.359
R1188 a_4439_159.n6 a_4439_159.t9 384.527
R1189 a_4439_159.n4 a_4439_159.t10 384.527
R1190 a_4439_159.n8 a_4439_159.t11 371.139
R1191 a_4439_159.n9 a_4439_159.t5 324.268
R1192 a_4439_159.n7 a_4439_159.t12 277.772
R1193 a_4439_159.n5 a_4439_159.t7 277.772
R1194 a_4439_159.n14 a_4439_159.n12 247.192
R1195 a_4439_159.n9 a_4439_159.n8 119.654
R1196 a_4439_159.n12 a_4439_159.n3 109.441
R1197 a_4439_159.n10 a_4439_159.n9 82.484
R1198 a_4439_159.n11 a_4439_159.n5 80.307
R1199 a_4439_159.n3 a_4439_159.n2 76.002
R1200 a_4439_159.n10 a_4439_159.n7 76
R1201 a_4439_159.n12 a_4439_159.n11 76
R1202 a_4439_159.n7 a_4439_159.n6 67.001
R1203 a_4439_159.n5 a_4439_159.n4 67.001
R1204 a_4439_159.n14 a_4439_159.n13 30
R1205 a_4439_159.n15 a_4439_159.n0 24.383
R1206 a_4439_159.n15 a_4439_159.n14 23.684
R1207 a_4439_159.n1 a_4439_159.t3 14.282
R1208 a_4439_159.n1 a_4439_159.t2 14.282
R1209 a_4439_159.n2 a_4439_159.t1 14.282
R1210 a_4439_159.n2 a_4439_159.t0 14.282
R1211 a_4439_159.n3 a_4439_159.n1 12.85
R1212 a_4439_159.n11 a_4439_159.n10 2.947
R1213 a_4383_75.n4 a_4383_75.n3 19.724
R1214 a_4383_75.t0 a_4383_75.n5 11.595
R1215 a_4383_75.t0 a_4383_75.n4 9.207
R1216 a_4383_75.n2 a_4383_75.n0 8.543
R1217 a_4383_75.t0 a_4383_75.n2 3.034
R1218 a_4383_75.n2 a_4383_75.n1 0.443
R1219 a_11887_383.n3 a_11887_383.t13 512.525
R1220 a_11887_383.n4 a_11887_383.t6 477.179
R1221 a_11887_383.n8 a_11887_383.t9 472.359
R1222 a_11887_383.n4 a_11887_383.t12 406.485
R1223 a_11887_383.n8 a_11887_383.t11 384.527
R1224 a_11887_383.n3 a_11887_383.t5 371.139
R1225 a_11887_383.n5 a_11887_383.t7 346.633
R1226 a_11887_383.n7 a_11887_383.t8 287.1
R1227 a_11887_383.n9 a_11887_383.t10 251.219
R1228 a_11887_383.n13 a_11887_383.n11 227.161
R1229 a_11887_383.n6 a_11887_383.n5 154.675
R1230 a_11887_383.n11 a_11887_383.n2 135.994
R1231 a_11887_383.n9 a_11887_383.n8 93.554
R1232 a_11887_383.n6 a_11887_383.n3 89.615
R1233 a_11887_383.n10 a_11887_383.n9 78.947
R1234 a_11887_383.n10 a_11887_383.n7 77.043
R1235 a_11887_383.n2 a_11887_383.n1 76.002
R1236 a_11887_383.n11 a_11887_383.n10 76
R1237 a_11887_383.n7 a_11887_383.n6 53.105
R1238 a_11887_383.n5 a_11887_383.n4 29.194
R1239 a_11887_383.n13 a_11887_383.n12 15.218
R1240 a_11887_383.n0 a_11887_383.t0 14.282
R1241 a_11887_383.n0 a_11887_383.t4 14.282
R1242 a_11887_383.n1 a_11887_383.t3 14.282
R1243 a_11887_383.n1 a_11887_383.t1 14.282
R1244 a_11887_383.n2 a_11887_383.n0 12.85
R1245 a_11887_383.n14 a_11887_383.n13 12.014
R1246 VPB VPB.n1382 126.832
R1247 VPB.n40 VPB.n38 94.117
R1248 VPB.n1324 VPB.n1322 94.117
R1249 VPB.n1261 VPB.n1259 94.117
R1250 VPB.n1198 VPB.n1196 94.117
R1251 VPB.n1135 VPB.n1133 94.117
R1252 VPB.n1072 VPB.n1070 94.117
R1253 VPB.n989 VPB.n987 94.117
R1254 VPB.n926 VPB.n924 94.117
R1255 VPB.n863 VPB.n861 94.117
R1256 VPB.n800 VPB.n798 94.117
R1257 VPB.n128 VPB.n126 94.117
R1258 VPB.n739 VPB.n737 94.117
R1259 VPB.n656 VPB.n654 94.117
R1260 VPB.n593 VPB.n591 94.117
R1261 VPB.n530 VPB.n528 94.117
R1262 VPB.n467 VPB.n465 94.117
R1263 VPB.n404 VPB.n402 94.117
R1264 VPB.n341 VPB.n339 94.117
R1265 VPB.n278 VPB.n276 94.117
R1266 VPB.n223 VPB.n221 94.117
R1267 VPB.n669 VPB.n668 80.104
R1268 VPB.n1002 VPB.n1001 80.104
R1269 VPB.n50 VPB.n49 80.104
R1270 VPB.n186 VPB.n185 76
R1271 VPB.n190 VPB.n189 76
R1272 VPB.n194 VPB.n193 76
R1273 VPB.n198 VPB.n197 76
R1274 VPB.n225 VPB.n224 76
R1275 VPB.n229 VPB.n228 76
R1276 VPB.n233 VPB.n232 76
R1277 VPB.n237 VPB.n236 76
R1278 VPB.n241 VPB.n240 76
R1279 VPB.n245 VPB.n244 76
R1280 VPB.n249 VPB.n248 76
R1281 VPB.n253 VPB.n252 76
R1282 VPB.n280 VPB.n279 76
R1283 VPB.n285 VPB.n284 76
R1284 VPB.n290 VPB.n289 76
R1285 VPB.n297 VPB.n296 76
R1286 VPB.n302 VPB.n301 76
R1287 VPB.n307 VPB.n306 76
R1288 VPB.n312 VPB.n311 76
R1289 VPB.n316 VPB.n315 76
R1290 VPB.n343 VPB.n342 76
R1291 VPB.n348 VPB.n347 76
R1292 VPB.n353 VPB.n352 76
R1293 VPB.n360 VPB.n359 76
R1294 VPB.n365 VPB.n364 76
R1295 VPB.n370 VPB.n369 76
R1296 VPB.n375 VPB.n374 76
R1297 VPB.n379 VPB.n378 76
R1298 VPB.n406 VPB.n405 76
R1299 VPB.n411 VPB.n410 76
R1300 VPB.n416 VPB.n415 76
R1301 VPB.n423 VPB.n422 76
R1302 VPB.n428 VPB.n427 76
R1303 VPB.n433 VPB.n432 76
R1304 VPB.n438 VPB.n437 76
R1305 VPB.n442 VPB.n441 76
R1306 VPB.n469 VPB.n468 76
R1307 VPB.n474 VPB.n473 76
R1308 VPB.n479 VPB.n478 76
R1309 VPB.n486 VPB.n485 76
R1310 VPB.n491 VPB.n490 76
R1311 VPB.n496 VPB.n495 76
R1312 VPB.n501 VPB.n500 76
R1313 VPB.n505 VPB.n504 76
R1314 VPB.n532 VPB.n531 76
R1315 VPB.n537 VPB.n536 76
R1316 VPB.n542 VPB.n541 76
R1317 VPB.n549 VPB.n548 76
R1318 VPB.n554 VPB.n553 76
R1319 VPB.n559 VPB.n558 76
R1320 VPB.n564 VPB.n563 76
R1321 VPB.n568 VPB.n567 76
R1322 VPB.n595 VPB.n594 76
R1323 VPB.n600 VPB.n599 76
R1324 VPB.n605 VPB.n604 76
R1325 VPB.n612 VPB.n611 76
R1326 VPB.n617 VPB.n616 76
R1327 VPB.n622 VPB.n621 76
R1328 VPB.n627 VPB.n626 76
R1329 VPB.n631 VPB.n630 76
R1330 VPB.n658 VPB.n657 76
R1331 VPB.n662 VPB.n661 76
R1332 VPB.n667 VPB.n666 76
R1333 VPB.n672 VPB.n671 76
R1334 VPB.n679 VPB.n678 76
R1335 VPB.n684 VPB.n683 76
R1336 VPB.n689 VPB.n688 76
R1337 VPB.n696 VPB.n695 76
R1338 VPB.n701 VPB.n700 76
R1339 VPB.n706 VPB.n705 76
R1340 VPB.n710 VPB.n709 76
R1341 VPB.n714 VPB.n713 76
R1342 VPB.n741 VPB.n740 76
R1343 VPB.n746 VPB.n745 76
R1344 VPB.n751 VPB.n750 76
R1345 VPB.n766 VPB.n762 76
R1346 VPB.n771 VPB.n770 76
R1347 VPB.n775 VPB.n774 76
R1348 VPB.n802 VPB.n801 76
R1349 VPB.n807 VPB.n806 76
R1350 VPB.n812 VPB.n811 76
R1351 VPB.n819 VPB.n818 76
R1352 VPB.n824 VPB.n823 76
R1353 VPB.n829 VPB.n828 76
R1354 VPB.n834 VPB.n833 76
R1355 VPB.n838 VPB.n837 76
R1356 VPB.n865 VPB.n864 76
R1357 VPB.n870 VPB.n869 76
R1358 VPB.n875 VPB.n874 76
R1359 VPB.n882 VPB.n881 76
R1360 VPB.n887 VPB.n886 76
R1361 VPB.n892 VPB.n891 76
R1362 VPB.n897 VPB.n896 76
R1363 VPB.n901 VPB.n900 76
R1364 VPB.n928 VPB.n927 76
R1365 VPB.n933 VPB.n932 76
R1366 VPB.n938 VPB.n937 76
R1367 VPB.n945 VPB.n944 76
R1368 VPB.n950 VPB.n949 76
R1369 VPB.n955 VPB.n954 76
R1370 VPB.n960 VPB.n959 76
R1371 VPB.n964 VPB.n963 76
R1372 VPB.n991 VPB.n990 76
R1373 VPB.n995 VPB.n994 76
R1374 VPB.n1000 VPB.n999 76
R1375 VPB.n1005 VPB.n1004 76
R1376 VPB.n1012 VPB.n1011 76
R1377 VPB.n1017 VPB.n1016 76
R1378 VPB.n1022 VPB.n1021 76
R1379 VPB.n1029 VPB.n1028 76
R1380 VPB.n1034 VPB.n1033 76
R1381 VPB.n1039 VPB.n1038 76
R1382 VPB.n1043 VPB.n1042 76
R1383 VPB.n1047 VPB.n1046 76
R1384 VPB.n1074 VPB.n1073 76
R1385 VPB.n1079 VPB.n1078 76
R1386 VPB.n1084 VPB.n1083 76
R1387 VPB.n1091 VPB.n1090 76
R1388 VPB.n1096 VPB.n1095 76
R1389 VPB.n1101 VPB.n1100 76
R1390 VPB.n1106 VPB.n1105 76
R1391 VPB.n1110 VPB.n1109 76
R1392 VPB.n1137 VPB.n1136 76
R1393 VPB.n1142 VPB.n1141 76
R1394 VPB.n1147 VPB.n1146 76
R1395 VPB.n1154 VPB.n1153 76
R1396 VPB.n1159 VPB.n1158 76
R1397 VPB.n1164 VPB.n1163 76
R1398 VPB.n1169 VPB.n1168 76
R1399 VPB.n1173 VPB.n1172 76
R1400 VPB.n1200 VPB.n1199 76
R1401 VPB.n1205 VPB.n1204 76
R1402 VPB.n1210 VPB.n1209 76
R1403 VPB.n1217 VPB.n1216 76
R1404 VPB.n1222 VPB.n1221 76
R1405 VPB.n1227 VPB.n1226 76
R1406 VPB.n1232 VPB.n1231 76
R1407 VPB.n1236 VPB.n1235 76
R1408 VPB.n1263 VPB.n1262 76
R1409 VPB.n1268 VPB.n1267 76
R1410 VPB.n1273 VPB.n1272 76
R1411 VPB.n1280 VPB.n1279 76
R1412 VPB.n1285 VPB.n1284 76
R1413 VPB.n1290 VPB.n1289 76
R1414 VPB.n1295 VPB.n1294 76
R1415 VPB.n1299 VPB.n1298 76
R1416 VPB.n1326 VPB.n1325 76
R1417 VPB.n1331 VPB.n1330 76
R1418 VPB.n1336 VPB.n1335 76
R1419 VPB.n1343 VPB.n1342 76
R1420 VPB.n1348 VPB.n1347 76
R1421 VPB.n1353 VPB.n1352 76
R1422 VPB.n1358 VPB.n1357 76
R1423 VPB.n1362 VPB.n1361 76
R1424 VPB.n1375 VPB.n1374 76
R1425 VPB.n698 VPB.n697 75.654
R1426 VPB.n1031 VPB.n1030 75.654
R1427 VPB.n72 VPB.n71 75.654
R1428 VPB.n22 VPB.n21 61.764
R1429 VPB.n1306 VPB.n1305 61.764
R1430 VPB.n1243 VPB.n1242 61.764
R1431 VPB.n1180 VPB.n1179 61.764
R1432 VPB.n1117 VPB.n1116 61.764
R1433 VPB.n1054 VPB.n1053 61.764
R1434 VPB.n971 VPB.n970 61.764
R1435 VPB.n908 VPB.n907 61.764
R1436 VPB.n845 VPB.n844 61.764
R1437 VPB.n782 VPB.n781 61.764
R1438 VPB.n89 VPB.n88 61.764
R1439 VPB.n721 VPB.n720 61.764
R1440 VPB.n638 VPB.n637 61.764
R1441 VPB.n575 VPB.n574 61.764
R1442 VPB.n512 VPB.n511 61.764
R1443 VPB.n449 VPB.n448 61.764
R1444 VPB.n386 VPB.n385 61.764
R1445 VPB.n323 VPB.n322 61.764
R1446 VPB.n260 VPB.n259 61.764
R1447 VPB.n205 VPB.n204 61.764
R1448 VPB.n308 VPB.t53 55.465
R1449 VPB.n281 VPB.t63 55.465
R1450 VPB.n78 VPB.t9 55.106
R1451 VPB.n1354 VPB.t17 55.106
R1452 VPB.n1291 VPB.t77 55.106
R1453 VPB.n1228 VPB.t12 55.106
R1454 VPB.n1165 VPB.t18 55.106
R1455 VPB.n1102 VPB.t41 55.106
R1456 VPB.n1035 VPB.t25 55.106
R1457 VPB.n956 VPB.t2 55.106
R1458 VPB.n893 VPB.t16 55.106
R1459 VPB.n830 VPB.t4 55.106
R1460 VPB.n767 VPB.t1 55.106
R1461 VPB.n118 VPB.t50 55.106
R1462 VPB.n702 VPB.t28 55.106
R1463 VPB.n623 VPB.t19 55.106
R1464 VPB.n560 VPB.t34 55.106
R1465 VPB.n497 VPB.t37 55.106
R1466 VPB.n434 VPB.t51 55.106
R1467 VPB.n371 VPB.t40 55.106
R1468 VPB.n45 VPB.t29 55.106
R1469 VPB.n1327 VPB.t46 55.106
R1470 VPB.n1264 VPB.t33 55.106
R1471 VPB.n1201 VPB.t65 55.106
R1472 VPB.n1138 VPB.t80 55.106
R1473 VPB.n1075 VPB.t8 55.106
R1474 VPB.n996 VPB.t13 55.106
R1475 VPB.n929 VPB.t43 55.106
R1476 VPB.n866 VPB.t23 55.106
R1477 VPB.n803 VPB.t72 55.106
R1478 VPB.n133 VPB.t64 55.106
R1479 VPB.n742 VPB.t26 55.106
R1480 VPB.n663 VPB.t39 55.106
R1481 VPB.n596 VPB.t48 55.106
R1482 VPB.n533 VPB.t38 55.106
R1483 VPB.n470 VPB.t74 55.106
R1484 VPB.n407 VPB.t56 55.106
R1485 VPB.n344 VPB.t32 55.106
R1486 VPB.n287 VPB.n286 48.952
R1487 VPB.n350 VPB.n349 48.952
R1488 VPB.n413 VPB.n412 48.952
R1489 VPB.n476 VPB.n475 48.952
R1490 VPB.n539 VPB.n538 48.952
R1491 VPB.n602 VPB.n601 48.952
R1492 VPB.n676 VPB.n675 48.952
R1493 VPB.n748 VPB.n747 48.952
R1494 VPB.n135 VPB.n134 48.952
R1495 VPB.n809 VPB.n808 48.952
R1496 VPB.n872 VPB.n871 48.952
R1497 VPB.n935 VPB.n934 48.952
R1498 VPB.n1009 VPB.n1008 48.952
R1499 VPB.n1081 VPB.n1080 48.952
R1500 VPB.n1144 VPB.n1143 48.952
R1501 VPB.n1207 VPB.n1206 48.952
R1502 VPB.n1270 VPB.n1269 48.952
R1503 VPB.n1333 VPB.n1332 48.952
R1504 VPB.n54 VPB.n53 48.952
R1505 VPB.n304 VPB.n303 44.502
R1506 VPB.n367 VPB.n366 44.502
R1507 VPB.n430 VPB.n429 44.502
R1508 VPB.n493 VPB.n492 44.502
R1509 VPB.n556 VPB.n555 44.502
R1510 VPB.n619 VPB.n618 44.502
R1511 VPB.n693 VPB.n692 44.502
R1512 VPB.n115 VPB.n114 44.502
R1513 VPB.n764 VPB.n763 44.502
R1514 VPB.n826 VPB.n825 44.502
R1515 VPB.n889 VPB.n888 44.502
R1516 VPB.n952 VPB.n951 44.502
R1517 VPB.n1026 VPB.n1025 44.502
R1518 VPB.n1098 VPB.n1097 44.502
R1519 VPB.n1161 VPB.n1160 44.502
R1520 VPB.n1224 VPB.n1223 44.502
R1521 VPB.n1287 VPB.n1286 44.502
R1522 VPB.n1350 VPB.n1349 44.502
R1523 VPB.n68 VPB.n67 44.502
R1524 VPB.n292 VPB.n291 41.183
R1525 VPB.n66 VPB.n14 40.824
R1526 VPB.n57 VPB.n15 40.824
R1527 VPB.n1338 VPB.n1337 40.824
R1528 VPB.n1275 VPB.n1274 40.824
R1529 VPB.n1212 VPB.n1211 40.824
R1530 VPB.n1149 VPB.n1148 40.824
R1531 VPB.n1086 VPB.n1085 40.824
R1532 VPB.n1024 VPB.n1023 40.824
R1533 VPB.n1007 VPB.n1006 40.824
R1534 VPB.n940 VPB.n939 40.824
R1535 VPB.n877 VPB.n876 40.824
R1536 VPB.n814 VPB.n813 40.824
R1537 VPB.n142 VPB.n82 40.824
R1538 VPB.n109 VPB.n104 40.824
R1539 VPB.n691 VPB.n690 40.824
R1540 VPB.n674 VPB.n673 40.824
R1541 VPB.n607 VPB.n606 40.824
R1542 VPB.n544 VPB.n543 40.824
R1543 VPB.n481 VPB.n480 40.824
R1544 VPB.n418 VPB.n417 40.824
R1545 VPB.n355 VPB.n354 40.824
R1546 VPB.n181 VPB.n180 35.118
R1547 VPB.n1379 VPB.n1375 20.452
R1548 VPB.n170 VPB.n167 20.452
R1549 VPB.n294 VPB.n293 17.801
R1550 VPB.n357 VPB.n356 17.801
R1551 VPB.n420 VPB.n419 17.801
R1552 VPB.n483 VPB.n482 17.801
R1553 VPB.n546 VPB.n545 17.801
R1554 VPB.n609 VPB.n608 17.801
R1555 VPB.n681 VPB.n680 17.801
R1556 VPB.n106 VPB.n105 17.801
R1557 VPB.n139 VPB.n138 17.801
R1558 VPB.n816 VPB.n815 17.801
R1559 VPB.n879 VPB.n878 17.801
R1560 VPB.n942 VPB.n941 17.801
R1561 VPB.n1014 VPB.n1013 17.801
R1562 VPB.n1088 VPB.n1087 17.801
R1563 VPB.n1151 VPB.n1150 17.801
R1564 VPB.n1214 VPB.n1213 17.801
R1565 VPB.n1277 VPB.n1276 17.801
R1566 VPB.n1340 VPB.n1339 17.801
R1567 VPB.n59 VPB.n58 17.801
R1568 VPB.n14 VPB.t69 14.282
R1569 VPB.n14 VPB.t21 14.282
R1570 VPB.n15 VPB.t30 14.282
R1571 VPB.n15 VPB.t70 14.282
R1572 VPB.n1337 VPB.t45 14.282
R1573 VPB.n1337 VPB.t10 14.282
R1574 VPB.n1274 VPB.t60 14.282
R1575 VPB.n1274 VPB.t58 14.282
R1576 VPB.n1211 VPB.t66 14.282
R1577 VPB.n1211 VPB.t6 14.282
R1578 VPB.n1148 VPB.t20 14.282
R1579 VPB.n1148 VPB.t14 14.282
R1580 VPB.n1085 VPB.t11 14.282
R1581 VPB.n1085 VPB.t57 14.282
R1582 VPB.n1023 VPB.t67 14.282
R1583 VPB.n1023 VPB.t24 14.282
R1584 VPB.n1006 VPB.t61 14.282
R1585 VPB.n1006 VPB.t68 14.282
R1586 VPB.n939 VPB.t47 14.282
R1587 VPB.n939 VPB.t7 14.282
R1588 VPB.n876 VPB.t22 14.282
R1589 VPB.n876 VPB.t15 14.282
R1590 VPB.n813 VPB.t71 14.282
R1591 VPB.n813 VPB.t5 14.282
R1592 VPB.n82 VPB.t0 14.282
R1593 VPB.n82 VPB.t3 14.282
R1594 VPB.n104 VPB.t27 14.282
R1595 VPB.n104 VPB.t49 14.282
R1596 VPB.n690 VPB.t73 14.282
R1597 VPB.n690 VPB.t81 14.282
R1598 VPB.n673 VPB.t52 14.282
R1599 VPB.n673 VPB.t75 14.282
R1600 VPB.n606 VPB.t44 14.282
R1601 VPB.n606 VPB.t35 14.282
R1602 VPB.n543 VPB.t42 14.282
R1603 VPB.n543 VPB.t31 14.282
R1604 VPB.n480 VPB.t76 14.282
R1605 VPB.n480 VPB.t36 14.282
R1606 VPB.n417 VPB.t55 14.282
R1607 VPB.n417 VPB.t59 14.282
R1608 VPB.n354 VPB.t79 14.282
R1609 VPB.n354 VPB.t78 14.282
R1610 VPB.n291 VPB.t62 14.282
R1611 VPB.n291 VPB.t54 14.282
R1612 VPB.n170 VPB.n169 13.653
R1613 VPB.n169 VPB.n168 13.653
R1614 VPB.n179 VPB.n178 13.653
R1615 VPB.n178 VPB.n177 13.653
R1616 VPB.n176 VPB.n175 13.653
R1617 VPB.n175 VPB.n174 13.653
R1618 VPB.n173 VPB.n172 13.653
R1619 VPB.n172 VPB.n171 13.653
R1620 VPB.n185 VPB.n184 13.653
R1621 VPB.n184 VPB.n183 13.653
R1622 VPB.n189 VPB.n188 13.653
R1623 VPB.n188 VPB.n187 13.653
R1624 VPB.n193 VPB.n192 13.653
R1625 VPB.n192 VPB.n191 13.653
R1626 VPB.n197 VPB.n196 13.653
R1627 VPB.n196 VPB.n195 13.653
R1628 VPB.n224 VPB.n223 13.653
R1629 VPB.n223 VPB.n222 13.653
R1630 VPB.n228 VPB.n227 13.653
R1631 VPB.n227 VPB.n226 13.653
R1632 VPB.n232 VPB.n231 13.653
R1633 VPB.n231 VPB.n230 13.653
R1634 VPB.n236 VPB.n235 13.653
R1635 VPB.n235 VPB.n234 13.653
R1636 VPB.n240 VPB.n239 13.653
R1637 VPB.n239 VPB.n238 13.653
R1638 VPB.n244 VPB.n243 13.653
R1639 VPB.n243 VPB.n242 13.653
R1640 VPB.n248 VPB.n247 13.653
R1641 VPB.n247 VPB.n246 13.653
R1642 VPB.n252 VPB.n251 13.653
R1643 VPB.n251 VPB.n250 13.653
R1644 VPB.n279 VPB.n278 13.653
R1645 VPB.n278 VPB.n277 13.653
R1646 VPB.n284 VPB.n283 13.653
R1647 VPB.n283 VPB.n282 13.653
R1648 VPB.n289 VPB.n288 13.653
R1649 VPB.n288 VPB.n287 13.653
R1650 VPB.n296 VPB.n295 13.653
R1651 VPB.n295 VPB.n294 13.653
R1652 VPB.n301 VPB.n300 13.653
R1653 VPB.n300 VPB.n299 13.653
R1654 VPB.n306 VPB.n305 13.653
R1655 VPB.n305 VPB.n304 13.653
R1656 VPB.n311 VPB.n310 13.653
R1657 VPB.n310 VPB.n309 13.653
R1658 VPB.n315 VPB.n314 13.653
R1659 VPB.n314 VPB.n313 13.653
R1660 VPB.n342 VPB.n341 13.653
R1661 VPB.n341 VPB.n340 13.653
R1662 VPB.n347 VPB.n346 13.653
R1663 VPB.n346 VPB.n345 13.653
R1664 VPB.n352 VPB.n351 13.653
R1665 VPB.n351 VPB.n350 13.653
R1666 VPB.n359 VPB.n358 13.653
R1667 VPB.n358 VPB.n357 13.653
R1668 VPB.n364 VPB.n363 13.653
R1669 VPB.n363 VPB.n362 13.653
R1670 VPB.n369 VPB.n368 13.653
R1671 VPB.n368 VPB.n367 13.653
R1672 VPB.n374 VPB.n373 13.653
R1673 VPB.n373 VPB.n372 13.653
R1674 VPB.n378 VPB.n377 13.653
R1675 VPB.n377 VPB.n376 13.653
R1676 VPB.n405 VPB.n404 13.653
R1677 VPB.n404 VPB.n403 13.653
R1678 VPB.n410 VPB.n409 13.653
R1679 VPB.n409 VPB.n408 13.653
R1680 VPB.n415 VPB.n414 13.653
R1681 VPB.n414 VPB.n413 13.653
R1682 VPB.n422 VPB.n421 13.653
R1683 VPB.n421 VPB.n420 13.653
R1684 VPB.n427 VPB.n426 13.653
R1685 VPB.n426 VPB.n425 13.653
R1686 VPB.n432 VPB.n431 13.653
R1687 VPB.n431 VPB.n430 13.653
R1688 VPB.n437 VPB.n436 13.653
R1689 VPB.n436 VPB.n435 13.653
R1690 VPB.n441 VPB.n440 13.653
R1691 VPB.n440 VPB.n439 13.653
R1692 VPB.n468 VPB.n467 13.653
R1693 VPB.n467 VPB.n466 13.653
R1694 VPB.n473 VPB.n472 13.653
R1695 VPB.n472 VPB.n471 13.653
R1696 VPB.n478 VPB.n477 13.653
R1697 VPB.n477 VPB.n476 13.653
R1698 VPB.n485 VPB.n484 13.653
R1699 VPB.n484 VPB.n483 13.653
R1700 VPB.n490 VPB.n489 13.653
R1701 VPB.n489 VPB.n488 13.653
R1702 VPB.n495 VPB.n494 13.653
R1703 VPB.n494 VPB.n493 13.653
R1704 VPB.n500 VPB.n499 13.653
R1705 VPB.n499 VPB.n498 13.653
R1706 VPB.n504 VPB.n503 13.653
R1707 VPB.n503 VPB.n502 13.653
R1708 VPB.n531 VPB.n530 13.653
R1709 VPB.n530 VPB.n529 13.653
R1710 VPB.n536 VPB.n535 13.653
R1711 VPB.n535 VPB.n534 13.653
R1712 VPB.n541 VPB.n540 13.653
R1713 VPB.n540 VPB.n539 13.653
R1714 VPB.n548 VPB.n547 13.653
R1715 VPB.n547 VPB.n546 13.653
R1716 VPB.n553 VPB.n552 13.653
R1717 VPB.n552 VPB.n551 13.653
R1718 VPB.n558 VPB.n557 13.653
R1719 VPB.n557 VPB.n556 13.653
R1720 VPB.n563 VPB.n562 13.653
R1721 VPB.n562 VPB.n561 13.653
R1722 VPB.n567 VPB.n566 13.653
R1723 VPB.n566 VPB.n565 13.653
R1724 VPB.n594 VPB.n593 13.653
R1725 VPB.n593 VPB.n592 13.653
R1726 VPB.n599 VPB.n598 13.653
R1727 VPB.n598 VPB.n597 13.653
R1728 VPB.n604 VPB.n603 13.653
R1729 VPB.n603 VPB.n602 13.653
R1730 VPB.n611 VPB.n610 13.653
R1731 VPB.n610 VPB.n609 13.653
R1732 VPB.n616 VPB.n615 13.653
R1733 VPB.n615 VPB.n614 13.653
R1734 VPB.n621 VPB.n620 13.653
R1735 VPB.n620 VPB.n619 13.653
R1736 VPB.n626 VPB.n625 13.653
R1737 VPB.n625 VPB.n624 13.653
R1738 VPB.n630 VPB.n629 13.653
R1739 VPB.n629 VPB.n628 13.653
R1740 VPB.n657 VPB.n656 13.653
R1741 VPB.n656 VPB.n655 13.653
R1742 VPB.n661 VPB.n660 13.653
R1743 VPB.n660 VPB.n659 13.653
R1744 VPB.n666 VPB.n665 13.653
R1745 VPB.n665 VPB.n664 13.653
R1746 VPB.n671 VPB.n670 13.653
R1747 VPB.n670 VPB.n669 13.653
R1748 VPB.n678 VPB.n677 13.653
R1749 VPB.n677 VPB.n676 13.653
R1750 VPB.n683 VPB.n682 13.653
R1751 VPB.n682 VPB.n681 13.653
R1752 VPB.n688 VPB.n687 13.653
R1753 VPB.n687 VPB.n686 13.653
R1754 VPB.n695 VPB.n694 13.653
R1755 VPB.n694 VPB.n693 13.653
R1756 VPB.n700 VPB.n699 13.653
R1757 VPB.n699 VPB.n698 13.653
R1758 VPB.n705 VPB.n704 13.653
R1759 VPB.n704 VPB.n703 13.653
R1760 VPB.n709 VPB.n708 13.653
R1761 VPB.n708 VPB.n707 13.653
R1762 VPB.n713 VPB.n712 13.653
R1763 VPB.n712 VPB.n711 13.653
R1764 VPB.n740 VPB.n739 13.653
R1765 VPB.n739 VPB.n738 13.653
R1766 VPB.n745 VPB.n744 13.653
R1767 VPB.n744 VPB.n743 13.653
R1768 VPB.n750 VPB.n749 13.653
R1769 VPB.n749 VPB.n748 13.653
R1770 VPB.n108 VPB.n107 13.653
R1771 VPB.n107 VPB.n106 13.653
R1772 VPB.n113 VPB.n112 13.653
R1773 VPB.n112 VPB.n111 13.653
R1774 VPB.n117 VPB.n116 13.653
R1775 VPB.n116 VPB.n115 13.653
R1776 VPB.n121 VPB.n120 13.653
R1777 VPB.n120 VPB.n119 13.653
R1778 VPB.n124 VPB.n123 13.653
R1779 VPB.n123 VPB.n122 13.653
R1780 VPB.n129 VPB.n128 13.653
R1781 VPB.n128 VPB.n127 13.653
R1782 VPB.n132 VPB.n131 13.653
R1783 VPB.n131 VPB.n130 13.653
R1784 VPB.n137 VPB.n136 13.653
R1785 VPB.n136 VPB.n135 13.653
R1786 VPB.n141 VPB.n140 13.653
R1787 VPB.n140 VPB.n139 13.653
R1788 VPB.n146 VPB.n145 13.653
R1789 VPB.n145 VPB.n144 13.653
R1790 VPB.n766 VPB.n765 13.653
R1791 VPB.n765 VPB.n764 13.653
R1792 VPB.n770 VPB.n769 13.653
R1793 VPB.n769 VPB.n768 13.653
R1794 VPB.n774 VPB.n773 13.653
R1795 VPB.n773 VPB.n772 13.653
R1796 VPB.n801 VPB.n800 13.653
R1797 VPB.n800 VPB.n799 13.653
R1798 VPB.n806 VPB.n805 13.653
R1799 VPB.n805 VPB.n804 13.653
R1800 VPB.n811 VPB.n810 13.653
R1801 VPB.n810 VPB.n809 13.653
R1802 VPB.n818 VPB.n817 13.653
R1803 VPB.n817 VPB.n816 13.653
R1804 VPB.n823 VPB.n822 13.653
R1805 VPB.n822 VPB.n821 13.653
R1806 VPB.n828 VPB.n827 13.653
R1807 VPB.n827 VPB.n826 13.653
R1808 VPB.n833 VPB.n832 13.653
R1809 VPB.n832 VPB.n831 13.653
R1810 VPB.n837 VPB.n836 13.653
R1811 VPB.n836 VPB.n835 13.653
R1812 VPB.n864 VPB.n863 13.653
R1813 VPB.n863 VPB.n862 13.653
R1814 VPB.n869 VPB.n868 13.653
R1815 VPB.n868 VPB.n867 13.653
R1816 VPB.n874 VPB.n873 13.653
R1817 VPB.n873 VPB.n872 13.653
R1818 VPB.n881 VPB.n880 13.653
R1819 VPB.n880 VPB.n879 13.653
R1820 VPB.n886 VPB.n885 13.653
R1821 VPB.n885 VPB.n884 13.653
R1822 VPB.n891 VPB.n890 13.653
R1823 VPB.n890 VPB.n889 13.653
R1824 VPB.n896 VPB.n895 13.653
R1825 VPB.n895 VPB.n894 13.653
R1826 VPB.n900 VPB.n899 13.653
R1827 VPB.n899 VPB.n898 13.653
R1828 VPB.n927 VPB.n926 13.653
R1829 VPB.n926 VPB.n925 13.653
R1830 VPB.n932 VPB.n931 13.653
R1831 VPB.n931 VPB.n930 13.653
R1832 VPB.n937 VPB.n936 13.653
R1833 VPB.n936 VPB.n935 13.653
R1834 VPB.n944 VPB.n943 13.653
R1835 VPB.n943 VPB.n942 13.653
R1836 VPB.n949 VPB.n948 13.653
R1837 VPB.n948 VPB.n947 13.653
R1838 VPB.n954 VPB.n953 13.653
R1839 VPB.n953 VPB.n952 13.653
R1840 VPB.n959 VPB.n958 13.653
R1841 VPB.n958 VPB.n957 13.653
R1842 VPB.n963 VPB.n962 13.653
R1843 VPB.n962 VPB.n961 13.653
R1844 VPB.n990 VPB.n989 13.653
R1845 VPB.n989 VPB.n988 13.653
R1846 VPB.n994 VPB.n993 13.653
R1847 VPB.n993 VPB.n992 13.653
R1848 VPB.n999 VPB.n998 13.653
R1849 VPB.n998 VPB.n997 13.653
R1850 VPB.n1004 VPB.n1003 13.653
R1851 VPB.n1003 VPB.n1002 13.653
R1852 VPB.n1011 VPB.n1010 13.653
R1853 VPB.n1010 VPB.n1009 13.653
R1854 VPB.n1016 VPB.n1015 13.653
R1855 VPB.n1015 VPB.n1014 13.653
R1856 VPB.n1021 VPB.n1020 13.653
R1857 VPB.n1020 VPB.n1019 13.653
R1858 VPB.n1028 VPB.n1027 13.653
R1859 VPB.n1027 VPB.n1026 13.653
R1860 VPB.n1033 VPB.n1032 13.653
R1861 VPB.n1032 VPB.n1031 13.653
R1862 VPB.n1038 VPB.n1037 13.653
R1863 VPB.n1037 VPB.n1036 13.653
R1864 VPB.n1042 VPB.n1041 13.653
R1865 VPB.n1041 VPB.n1040 13.653
R1866 VPB.n1046 VPB.n1045 13.653
R1867 VPB.n1045 VPB.n1044 13.653
R1868 VPB.n1073 VPB.n1072 13.653
R1869 VPB.n1072 VPB.n1071 13.653
R1870 VPB.n1078 VPB.n1077 13.653
R1871 VPB.n1077 VPB.n1076 13.653
R1872 VPB.n1083 VPB.n1082 13.653
R1873 VPB.n1082 VPB.n1081 13.653
R1874 VPB.n1090 VPB.n1089 13.653
R1875 VPB.n1089 VPB.n1088 13.653
R1876 VPB.n1095 VPB.n1094 13.653
R1877 VPB.n1094 VPB.n1093 13.653
R1878 VPB.n1100 VPB.n1099 13.653
R1879 VPB.n1099 VPB.n1098 13.653
R1880 VPB.n1105 VPB.n1104 13.653
R1881 VPB.n1104 VPB.n1103 13.653
R1882 VPB.n1109 VPB.n1108 13.653
R1883 VPB.n1108 VPB.n1107 13.653
R1884 VPB.n1136 VPB.n1135 13.653
R1885 VPB.n1135 VPB.n1134 13.653
R1886 VPB.n1141 VPB.n1140 13.653
R1887 VPB.n1140 VPB.n1139 13.653
R1888 VPB.n1146 VPB.n1145 13.653
R1889 VPB.n1145 VPB.n1144 13.653
R1890 VPB.n1153 VPB.n1152 13.653
R1891 VPB.n1152 VPB.n1151 13.653
R1892 VPB.n1158 VPB.n1157 13.653
R1893 VPB.n1157 VPB.n1156 13.653
R1894 VPB.n1163 VPB.n1162 13.653
R1895 VPB.n1162 VPB.n1161 13.653
R1896 VPB.n1168 VPB.n1167 13.653
R1897 VPB.n1167 VPB.n1166 13.653
R1898 VPB.n1172 VPB.n1171 13.653
R1899 VPB.n1171 VPB.n1170 13.653
R1900 VPB.n1199 VPB.n1198 13.653
R1901 VPB.n1198 VPB.n1197 13.653
R1902 VPB.n1204 VPB.n1203 13.653
R1903 VPB.n1203 VPB.n1202 13.653
R1904 VPB.n1209 VPB.n1208 13.653
R1905 VPB.n1208 VPB.n1207 13.653
R1906 VPB.n1216 VPB.n1215 13.653
R1907 VPB.n1215 VPB.n1214 13.653
R1908 VPB.n1221 VPB.n1220 13.653
R1909 VPB.n1220 VPB.n1219 13.653
R1910 VPB.n1226 VPB.n1225 13.653
R1911 VPB.n1225 VPB.n1224 13.653
R1912 VPB.n1231 VPB.n1230 13.653
R1913 VPB.n1230 VPB.n1229 13.653
R1914 VPB.n1235 VPB.n1234 13.653
R1915 VPB.n1234 VPB.n1233 13.653
R1916 VPB.n1262 VPB.n1261 13.653
R1917 VPB.n1261 VPB.n1260 13.653
R1918 VPB.n1267 VPB.n1266 13.653
R1919 VPB.n1266 VPB.n1265 13.653
R1920 VPB.n1272 VPB.n1271 13.653
R1921 VPB.n1271 VPB.n1270 13.653
R1922 VPB.n1279 VPB.n1278 13.653
R1923 VPB.n1278 VPB.n1277 13.653
R1924 VPB.n1284 VPB.n1283 13.653
R1925 VPB.n1283 VPB.n1282 13.653
R1926 VPB.n1289 VPB.n1288 13.653
R1927 VPB.n1288 VPB.n1287 13.653
R1928 VPB.n1294 VPB.n1293 13.653
R1929 VPB.n1293 VPB.n1292 13.653
R1930 VPB.n1298 VPB.n1297 13.653
R1931 VPB.n1297 VPB.n1296 13.653
R1932 VPB.n1325 VPB.n1324 13.653
R1933 VPB.n1324 VPB.n1323 13.653
R1934 VPB.n1330 VPB.n1329 13.653
R1935 VPB.n1329 VPB.n1328 13.653
R1936 VPB.n1335 VPB.n1334 13.653
R1937 VPB.n1334 VPB.n1333 13.653
R1938 VPB.n1342 VPB.n1341 13.653
R1939 VPB.n1341 VPB.n1340 13.653
R1940 VPB.n1347 VPB.n1346 13.653
R1941 VPB.n1346 VPB.n1345 13.653
R1942 VPB.n1352 VPB.n1351 13.653
R1943 VPB.n1351 VPB.n1350 13.653
R1944 VPB.n1357 VPB.n1356 13.653
R1945 VPB.n1356 VPB.n1355 13.653
R1946 VPB.n1361 VPB.n1360 13.653
R1947 VPB.n1360 VPB.n1359 13.653
R1948 VPB.n41 VPB.n40 13.653
R1949 VPB.n40 VPB.n39 13.653
R1950 VPB.n44 VPB.n43 13.653
R1951 VPB.n43 VPB.n42 13.653
R1952 VPB.n48 VPB.n47 13.653
R1953 VPB.n47 VPB.n46 13.653
R1954 VPB.n52 VPB.n51 13.653
R1955 VPB.n51 VPB.n50 13.653
R1956 VPB.n56 VPB.n55 13.653
R1957 VPB.n55 VPB.n54 13.653
R1958 VPB.n61 VPB.n60 13.653
R1959 VPB.n60 VPB.n59 13.653
R1960 VPB.n65 VPB.n64 13.653
R1961 VPB.n64 VPB.n63 13.653
R1962 VPB.n70 VPB.n69 13.653
R1963 VPB.n69 VPB.n68 13.653
R1964 VPB.n74 VPB.n73 13.653
R1965 VPB.n73 VPB.n72 13.653
R1966 VPB.n77 VPB.n76 13.653
R1967 VPB.n76 VPB.n75 13.653
R1968 VPB.n81 VPB.n80 13.653
R1969 VPB.n80 VPB.n79 13.653
R1970 VPB.n1375 VPB.n0 13.653
R1971 VPB VPB.n0 13.653
R1972 VPB.n299 VPB.n298 13.35
R1973 VPB.n362 VPB.n361 13.35
R1974 VPB.n425 VPB.n424 13.35
R1975 VPB.n488 VPB.n487 13.35
R1976 VPB.n551 VPB.n550 13.35
R1977 VPB.n614 VPB.n613 13.35
R1978 VPB.n686 VPB.n685 13.35
R1979 VPB.n111 VPB.n110 13.35
R1980 VPB.n144 VPB.n143 13.35
R1981 VPB.n821 VPB.n820 13.35
R1982 VPB.n884 VPB.n883 13.35
R1983 VPB.n947 VPB.n946 13.35
R1984 VPB.n1019 VPB.n1018 13.35
R1985 VPB.n1093 VPB.n1092 13.35
R1986 VPB.n1156 VPB.n1155 13.35
R1987 VPB.n1219 VPB.n1218 13.35
R1988 VPB.n1282 VPB.n1281 13.35
R1989 VPB.n1345 VPB.n1344 13.35
R1990 VPB.n63 VPB.n62 13.35
R1991 VPB.n1379 VPB.n1378 13.276
R1992 VPB.n1378 VPB.n1376 13.276
R1993 VPB.n36 VPB.n18 13.276
R1994 VPB.n18 VPB.n16 13.276
R1995 VPB.n1320 VPB.n1302 13.276
R1996 VPB.n1302 VPB.n1300 13.276
R1997 VPB.n1257 VPB.n1239 13.276
R1998 VPB.n1239 VPB.n1237 13.276
R1999 VPB.n1194 VPB.n1176 13.276
R2000 VPB.n1176 VPB.n1174 13.276
R2001 VPB.n1131 VPB.n1113 13.276
R2002 VPB.n1113 VPB.n1111 13.276
R2003 VPB.n1068 VPB.n1050 13.276
R2004 VPB.n1050 VPB.n1048 13.276
R2005 VPB.n985 VPB.n967 13.276
R2006 VPB.n967 VPB.n965 13.276
R2007 VPB.n922 VPB.n904 13.276
R2008 VPB.n904 VPB.n902 13.276
R2009 VPB.n859 VPB.n841 13.276
R2010 VPB.n841 VPB.n839 13.276
R2011 VPB.n796 VPB.n778 13.276
R2012 VPB.n778 VPB.n776 13.276
R2013 VPB.n103 VPB.n85 13.276
R2014 VPB.n85 VPB.n83 13.276
R2015 VPB.n735 VPB.n717 13.276
R2016 VPB.n717 VPB.n715 13.276
R2017 VPB.n652 VPB.n634 13.276
R2018 VPB.n634 VPB.n632 13.276
R2019 VPB.n589 VPB.n571 13.276
R2020 VPB.n571 VPB.n569 13.276
R2021 VPB.n526 VPB.n508 13.276
R2022 VPB.n508 VPB.n506 13.276
R2023 VPB.n463 VPB.n445 13.276
R2024 VPB.n445 VPB.n443 13.276
R2025 VPB.n400 VPB.n382 13.276
R2026 VPB.n382 VPB.n380 13.276
R2027 VPB.n337 VPB.n319 13.276
R2028 VPB.n319 VPB.n317 13.276
R2029 VPB.n274 VPB.n256 13.276
R2030 VPB.n256 VPB.n254 13.276
R2031 VPB.n219 VPB.n201 13.276
R2032 VPB.n201 VPB.n199 13.276
R2033 VPB.n179 VPB.n176 13.276
R2034 VPB.n176 VPB.n173 13.276
R2035 VPB.n224 VPB.n220 13.276
R2036 VPB.n279 VPB.n275 13.276
R2037 VPB.n342 VPB.n338 13.276
R2038 VPB.n405 VPB.n401 13.276
R2039 VPB.n468 VPB.n464 13.276
R2040 VPB.n531 VPB.n527 13.276
R2041 VPB.n594 VPB.n590 13.276
R2042 VPB.n657 VPB.n653 13.276
R2043 VPB.n740 VPB.n736 13.276
R2044 VPB.n117 VPB.n113 13.276
R2045 VPB.n124 VPB.n121 13.276
R2046 VPB.n125 VPB.n124 13.276
R2047 VPB.n129 VPB.n125 13.276
R2048 VPB.n132 VPB.n129 13.276
R2049 VPB.n141 VPB.n137 13.276
R2050 VPB.n766 VPB.n146 13.276
R2051 VPB.n801 VPB.n797 13.276
R2052 VPB.n864 VPB.n860 13.276
R2053 VPB.n927 VPB.n923 13.276
R2054 VPB.n990 VPB.n986 13.276
R2055 VPB.n1073 VPB.n1069 13.276
R2056 VPB.n1136 VPB.n1132 13.276
R2057 VPB.n1199 VPB.n1195 13.276
R2058 VPB.n1262 VPB.n1258 13.276
R2059 VPB.n1325 VPB.n1321 13.276
R2060 VPB.n41 VPB.n37 13.276
R2061 VPB.n44 VPB.n41 13.276
R2062 VPB.n52 VPB.n48 13.276
R2063 VPB.n56 VPB.n52 13.276
R2064 VPB.n65 VPB.n61 13.276
R2065 VPB.n74 VPB.n70 13.276
R2066 VPB.n77 VPB.n74 13.276
R2067 VPB.n1375 VPB.n81 13.276
R2068 VPB.n167 VPB.n149 13.276
R2069 VPB.n149 VPB.n147 13.276
R2070 VPB.n154 VPB.n152 12.796
R2071 VPB.n154 VPB.n153 12.564
R2072 VPB.n81 VPB.n78 12.558
R2073 VPB.n45 VPB.n44 12.2
R2074 VPB.n162 VPB.n161 12.198
R2075 VPB.n158 VPB.n157 12.198
R2076 VPB.n162 VPB.n159 12.198
R2077 VPB.n137 VPB.n133 11.841
R2078 VPB.n118 VPB.n117 11.482
R2079 VPB.n767 VPB.n766 11.482
R2080 VPB.n61 VPB.n57 9.329
R2081 VPB.n66 VPB.n65 8.97
R2082 VPB.n167 VPB.n166 7.5
R2083 VPB.n152 VPB.n151 7.5
R2084 VPB.n157 VPB.n156 7.5
R2085 VPB.n161 VPB.n160 7.5
R2086 VPB.n149 VPB.n148 7.5
R2087 VPB.n164 VPB.n150 7.5
R2088 VPB.n201 VPB.n200 7.5
R2089 VPB.n214 VPB.n213 7.5
R2090 VPB.n208 VPB.n207 7.5
R2091 VPB.n210 VPB.n209 7.5
R2092 VPB.n203 VPB.n202 7.5
R2093 VPB.n219 VPB.n218 7.5
R2094 VPB.n256 VPB.n255 7.5
R2095 VPB.n269 VPB.n268 7.5
R2096 VPB.n263 VPB.n262 7.5
R2097 VPB.n265 VPB.n264 7.5
R2098 VPB.n258 VPB.n257 7.5
R2099 VPB.n274 VPB.n273 7.5
R2100 VPB.n319 VPB.n318 7.5
R2101 VPB.n332 VPB.n331 7.5
R2102 VPB.n326 VPB.n325 7.5
R2103 VPB.n328 VPB.n327 7.5
R2104 VPB.n321 VPB.n320 7.5
R2105 VPB.n337 VPB.n336 7.5
R2106 VPB.n382 VPB.n381 7.5
R2107 VPB.n395 VPB.n394 7.5
R2108 VPB.n389 VPB.n388 7.5
R2109 VPB.n391 VPB.n390 7.5
R2110 VPB.n384 VPB.n383 7.5
R2111 VPB.n400 VPB.n399 7.5
R2112 VPB.n445 VPB.n444 7.5
R2113 VPB.n458 VPB.n457 7.5
R2114 VPB.n452 VPB.n451 7.5
R2115 VPB.n454 VPB.n453 7.5
R2116 VPB.n447 VPB.n446 7.5
R2117 VPB.n463 VPB.n462 7.5
R2118 VPB.n508 VPB.n507 7.5
R2119 VPB.n521 VPB.n520 7.5
R2120 VPB.n515 VPB.n514 7.5
R2121 VPB.n517 VPB.n516 7.5
R2122 VPB.n510 VPB.n509 7.5
R2123 VPB.n526 VPB.n525 7.5
R2124 VPB.n571 VPB.n570 7.5
R2125 VPB.n584 VPB.n583 7.5
R2126 VPB.n578 VPB.n577 7.5
R2127 VPB.n580 VPB.n579 7.5
R2128 VPB.n573 VPB.n572 7.5
R2129 VPB.n589 VPB.n588 7.5
R2130 VPB.n634 VPB.n633 7.5
R2131 VPB.n647 VPB.n646 7.5
R2132 VPB.n641 VPB.n640 7.5
R2133 VPB.n643 VPB.n642 7.5
R2134 VPB.n636 VPB.n635 7.5
R2135 VPB.n652 VPB.n651 7.5
R2136 VPB.n717 VPB.n716 7.5
R2137 VPB.n730 VPB.n729 7.5
R2138 VPB.n724 VPB.n723 7.5
R2139 VPB.n726 VPB.n725 7.5
R2140 VPB.n719 VPB.n718 7.5
R2141 VPB.n735 VPB.n734 7.5
R2142 VPB.n85 VPB.n84 7.5
R2143 VPB.n98 VPB.n97 7.5
R2144 VPB.n92 VPB.n91 7.5
R2145 VPB.n94 VPB.n93 7.5
R2146 VPB.n87 VPB.n86 7.5
R2147 VPB.n103 VPB.n102 7.5
R2148 VPB.n778 VPB.n777 7.5
R2149 VPB.n791 VPB.n790 7.5
R2150 VPB.n785 VPB.n784 7.5
R2151 VPB.n787 VPB.n786 7.5
R2152 VPB.n780 VPB.n779 7.5
R2153 VPB.n796 VPB.n795 7.5
R2154 VPB.n841 VPB.n840 7.5
R2155 VPB.n854 VPB.n853 7.5
R2156 VPB.n848 VPB.n847 7.5
R2157 VPB.n850 VPB.n849 7.5
R2158 VPB.n843 VPB.n842 7.5
R2159 VPB.n859 VPB.n858 7.5
R2160 VPB.n904 VPB.n903 7.5
R2161 VPB.n917 VPB.n916 7.5
R2162 VPB.n911 VPB.n910 7.5
R2163 VPB.n913 VPB.n912 7.5
R2164 VPB.n906 VPB.n905 7.5
R2165 VPB.n922 VPB.n921 7.5
R2166 VPB.n967 VPB.n966 7.5
R2167 VPB.n980 VPB.n979 7.5
R2168 VPB.n974 VPB.n973 7.5
R2169 VPB.n976 VPB.n975 7.5
R2170 VPB.n969 VPB.n968 7.5
R2171 VPB.n985 VPB.n984 7.5
R2172 VPB.n1050 VPB.n1049 7.5
R2173 VPB.n1063 VPB.n1062 7.5
R2174 VPB.n1057 VPB.n1056 7.5
R2175 VPB.n1059 VPB.n1058 7.5
R2176 VPB.n1052 VPB.n1051 7.5
R2177 VPB.n1068 VPB.n1067 7.5
R2178 VPB.n1113 VPB.n1112 7.5
R2179 VPB.n1126 VPB.n1125 7.5
R2180 VPB.n1120 VPB.n1119 7.5
R2181 VPB.n1122 VPB.n1121 7.5
R2182 VPB.n1115 VPB.n1114 7.5
R2183 VPB.n1131 VPB.n1130 7.5
R2184 VPB.n1176 VPB.n1175 7.5
R2185 VPB.n1189 VPB.n1188 7.5
R2186 VPB.n1183 VPB.n1182 7.5
R2187 VPB.n1185 VPB.n1184 7.5
R2188 VPB.n1178 VPB.n1177 7.5
R2189 VPB.n1194 VPB.n1193 7.5
R2190 VPB.n1239 VPB.n1238 7.5
R2191 VPB.n1252 VPB.n1251 7.5
R2192 VPB.n1246 VPB.n1245 7.5
R2193 VPB.n1248 VPB.n1247 7.5
R2194 VPB.n1241 VPB.n1240 7.5
R2195 VPB.n1257 VPB.n1256 7.5
R2196 VPB.n1302 VPB.n1301 7.5
R2197 VPB.n1315 VPB.n1314 7.5
R2198 VPB.n1309 VPB.n1308 7.5
R2199 VPB.n1311 VPB.n1310 7.5
R2200 VPB.n1304 VPB.n1303 7.5
R2201 VPB.n1320 VPB.n1319 7.5
R2202 VPB.n18 VPB.n17 7.5
R2203 VPB.n31 VPB.n30 7.5
R2204 VPB.n25 VPB.n24 7.5
R2205 VPB.n27 VPB.n26 7.5
R2206 VPB.n20 VPB.n19 7.5
R2207 VPB.n36 VPB.n35 7.5
R2208 VPB.n1378 VPB.n1377 7.5
R2209 VPB.n12 VPB.n11 7.5
R2210 VPB.n6 VPB.n5 7.5
R2211 VPB.n8 VPB.n7 7.5
R2212 VPB.n2 VPB.n1 7.5
R2213 VPB.n1380 VPB.n1379 7.5
R2214 VPB.n37 VPB.n36 7.176
R2215 VPB.n1321 VPB.n1320 7.176
R2216 VPB.n1258 VPB.n1257 7.176
R2217 VPB.n1195 VPB.n1194 7.176
R2218 VPB.n1132 VPB.n1131 7.176
R2219 VPB.n1069 VPB.n1068 7.176
R2220 VPB.n986 VPB.n985 7.176
R2221 VPB.n923 VPB.n922 7.176
R2222 VPB.n860 VPB.n859 7.176
R2223 VPB.n797 VPB.n796 7.176
R2224 VPB.n125 VPB.n103 7.176
R2225 VPB.n736 VPB.n735 7.176
R2226 VPB.n653 VPB.n652 7.176
R2227 VPB.n590 VPB.n589 7.176
R2228 VPB.n527 VPB.n526 7.176
R2229 VPB.n464 VPB.n463 7.176
R2230 VPB.n401 VPB.n400 7.176
R2231 VPB.n338 VPB.n337 7.176
R2232 VPB.n275 VPB.n274 7.176
R2233 VPB.n220 VPB.n219 7.176
R2234 VPB.n113 VPB.n109 6.817
R2235 VPB.n146 VPB.n142 6.817
R2236 VPB.n215 VPB.n212 6.729
R2237 VPB.n211 VPB.n208 6.729
R2238 VPB.n206 VPB.n203 6.729
R2239 VPB.n270 VPB.n267 6.729
R2240 VPB.n266 VPB.n263 6.729
R2241 VPB.n261 VPB.n258 6.729
R2242 VPB.n333 VPB.n330 6.729
R2243 VPB.n329 VPB.n326 6.729
R2244 VPB.n324 VPB.n321 6.729
R2245 VPB.n396 VPB.n393 6.729
R2246 VPB.n392 VPB.n389 6.729
R2247 VPB.n387 VPB.n384 6.729
R2248 VPB.n459 VPB.n456 6.729
R2249 VPB.n455 VPB.n452 6.729
R2250 VPB.n450 VPB.n447 6.729
R2251 VPB.n522 VPB.n519 6.729
R2252 VPB.n518 VPB.n515 6.729
R2253 VPB.n513 VPB.n510 6.729
R2254 VPB.n585 VPB.n582 6.729
R2255 VPB.n581 VPB.n578 6.729
R2256 VPB.n576 VPB.n573 6.729
R2257 VPB.n648 VPB.n645 6.729
R2258 VPB.n644 VPB.n641 6.729
R2259 VPB.n639 VPB.n636 6.729
R2260 VPB.n731 VPB.n728 6.729
R2261 VPB.n727 VPB.n724 6.729
R2262 VPB.n722 VPB.n719 6.729
R2263 VPB.n99 VPB.n96 6.729
R2264 VPB.n95 VPB.n92 6.729
R2265 VPB.n90 VPB.n87 6.729
R2266 VPB.n792 VPB.n789 6.729
R2267 VPB.n788 VPB.n785 6.729
R2268 VPB.n783 VPB.n780 6.729
R2269 VPB.n855 VPB.n852 6.729
R2270 VPB.n851 VPB.n848 6.729
R2271 VPB.n846 VPB.n843 6.729
R2272 VPB.n918 VPB.n915 6.729
R2273 VPB.n914 VPB.n911 6.729
R2274 VPB.n909 VPB.n906 6.729
R2275 VPB.n981 VPB.n978 6.729
R2276 VPB.n977 VPB.n974 6.729
R2277 VPB.n972 VPB.n969 6.729
R2278 VPB.n1064 VPB.n1061 6.729
R2279 VPB.n1060 VPB.n1057 6.729
R2280 VPB.n1055 VPB.n1052 6.729
R2281 VPB.n1127 VPB.n1124 6.729
R2282 VPB.n1123 VPB.n1120 6.729
R2283 VPB.n1118 VPB.n1115 6.729
R2284 VPB.n1190 VPB.n1187 6.729
R2285 VPB.n1186 VPB.n1183 6.729
R2286 VPB.n1181 VPB.n1178 6.729
R2287 VPB.n1253 VPB.n1250 6.729
R2288 VPB.n1249 VPB.n1246 6.729
R2289 VPB.n1244 VPB.n1241 6.729
R2290 VPB.n1316 VPB.n1313 6.729
R2291 VPB.n1312 VPB.n1309 6.729
R2292 VPB.n1307 VPB.n1304 6.729
R2293 VPB.n32 VPB.n29 6.729
R2294 VPB.n28 VPB.n25 6.729
R2295 VPB.n23 VPB.n20 6.729
R2296 VPB.n13 VPB.n10 6.729
R2297 VPB.n9 VPB.n6 6.729
R2298 VPB.n4 VPB.n2 6.729
R2299 VPB.n206 VPB.n205 6.728
R2300 VPB.n211 VPB.n210 6.728
R2301 VPB.n215 VPB.n214 6.728
R2302 VPB.n218 VPB.n217 6.728
R2303 VPB.n261 VPB.n260 6.728
R2304 VPB.n266 VPB.n265 6.728
R2305 VPB.n270 VPB.n269 6.728
R2306 VPB.n273 VPB.n272 6.728
R2307 VPB.n324 VPB.n323 6.728
R2308 VPB.n329 VPB.n328 6.728
R2309 VPB.n333 VPB.n332 6.728
R2310 VPB.n336 VPB.n335 6.728
R2311 VPB.n387 VPB.n386 6.728
R2312 VPB.n392 VPB.n391 6.728
R2313 VPB.n396 VPB.n395 6.728
R2314 VPB.n399 VPB.n398 6.728
R2315 VPB.n450 VPB.n449 6.728
R2316 VPB.n455 VPB.n454 6.728
R2317 VPB.n459 VPB.n458 6.728
R2318 VPB.n462 VPB.n461 6.728
R2319 VPB.n513 VPB.n512 6.728
R2320 VPB.n518 VPB.n517 6.728
R2321 VPB.n522 VPB.n521 6.728
R2322 VPB.n525 VPB.n524 6.728
R2323 VPB.n576 VPB.n575 6.728
R2324 VPB.n581 VPB.n580 6.728
R2325 VPB.n585 VPB.n584 6.728
R2326 VPB.n588 VPB.n587 6.728
R2327 VPB.n639 VPB.n638 6.728
R2328 VPB.n644 VPB.n643 6.728
R2329 VPB.n648 VPB.n647 6.728
R2330 VPB.n651 VPB.n650 6.728
R2331 VPB.n722 VPB.n721 6.728
R2332 VPB.n727 VPB.n726 6.728
R2333 VPB.n731 VPB.n730 6.728
R2334 VPB.n734 VPB.n733 6.728
R2335 VPB.n90 VPB.n89 6.728
R2336 VPB.n95 VPB.n94 6.728
R2337 VPB.n99 VPB.n98 6.728
R2338 VPB.n102 VPB.n101 6.728
R2339 VPB.n783 VPB.n782 6.728
R2340 VPB.n788 VPB.n787 6.728
R2341 VPB.n792 VPB.n791 6.728
R2342 VPB.n795 VPB.n794 6.728
R2343 VPB.n846 VPB.n845 6.728
R2344 VPB.n851 VPB.n850 6.728
R2345 VPB.n855 VPB.n854 6.728
R2346 VPB.n858 VPB.n857 6.728
R2347 VPB.n909 VPB.n908 6.728
R2348 VPB.n914 VPB.n913 6.728
R2349 VPB.n918 VPB.n917 6.728
R2350 VPB.n921 VPB.n920 6.728
R2351 VPB.n972 VPB.n971 6.728
R2352 VPB.n977 VPB.n976 6.728
R2353 VPB.n981 VPB.n980 6.728
R2354 VPB.n984 VPB.n983 6.728
R2355 VPB.n1055 VPB.n1054 6.728
R2356 VPB.n1060 VPB.n1059 6.728
R2357 VPB.n1064 VPB.n1063 6.728
R2358 VPB.n1067 VPB.n1066 6.728
R2359 VPB.n1118 VPB.n1117 6.728
R2360 VPB.n1123 VPB.n1122 6.728
R2361 VPB.n1127 VPB.n1126 6.728
R2362 VPB.n1130 VPB.n1129 6.728
R2363 VPB.n1181 VPB.n1180 6.728
R2364 VPB.n1186 VPB.n1185 6.728
R2365 VPB.n1190 VPB.n1189 6.728
R2366 VPB.n1193 VPB.n1192 6.728
R2367 VPB.n1244 VPB.n1243 6.728
R2368 VPB.n1249 VPB.n1248 6.728
R2369 VPB.n1253 VPB.n1252 6.728
R2370 VPB.n1256 VPB.n1255 6.728
R2371 VPB.n1307 VPB.n1306 6.728
R2372 VPB.n1312 VPB.n1311 6.728
R2373 VPB.n1316 VPB.n1315 6.728
R2374 VPB.n1319 VPB.n1318 6.728
R2375 VPB.n23 VPB.n22 6.728
R2376 VPB.n28 VPB.n27 6.728
R2377 VPB.n32 VPB.n31 6.728
R2378 VPB.n35 VPB.n34 6.728
R2379 VPB.n4 VPB.n3 6.728
R2380 VPB.n9 VPB.n8 6.728
R2381 VPB.n13 VPB.n12 6.728
R2382 VPB.n1381 VPB.n1380 6.728
R2383 VPB.n296 VPB.n292 6.458
R2384 VPB.n359 VPB.n355 6.458
R2385 VPB.n422 VPB.n418 6.458
R2386 VPB.n485 VPB.n481 6.458
R2387 VPB.n548 VPB.n544 6.458
R2388 VPB.n611 VPB.n607 6.458
R2389 VPB.n109 VPB.n108 6.458
R2390 VPB.n142 VPB.n141 6.458
R2391 VPB.n818 VPB.n814 6.458
R2392 VPB.n881 VPB.n877 6.458
R2393 VPB.n944 VPB.n940 6.458
R2394 VPB.n1090 VPB.n1086 6.458
R2395 VPB.n1153 VPB.n1149 6.458
R2396 VPB.n1216 VPB.n1212 6.458
R2397 VPB.n1279 VPB.n1275 6.458
R2398 VPB.n1342 VPB.n1338 6.458
R2399 VPB.n166 VPB.n165 6.398
R2400 VPB.n180 VPB.n170 6.112
R2401 VPB.n180 VPB.n179 6.101
R2402 VPB.n695 VPB.n691 4.305
R2403 VPB.n1028 VPB.n1024 4.305
R2404 VPB.n70 VPB.n66 4.305
R2405 VPB.n678 VPB.n674 3.947
R2406 VPB.n1011 VPB.n1007 3.947
R2407 VPB.n57 VPB.n56 3.947
R2408 VPB.n311 VPB.n308 1.794
R2409 VPB.n374 VPB.n371 1.794
R2410 VPB.n437 VPB.n434 1.794
R2411 VPB.n500 VPB.n497 1.794
R2412 VPB.n563 VPB.n560 1.794
R2413 VPB.n626 VPB.n623 1.794
R2414 VPB.n121 VPB.n118 1.794
R2415 VPB.n770 VPB.n767 1.794
R2416 VPB.n833 VPB.n830 1.794
R2417 VPB.n896 VPB.n893 1.794
R2418 VPB.n959 VPB.n956 1.794
R2419 VPB.n1105 VPB.n1102 1.794
R2420 VPB.n1168 VPB.n1165 1.794
R2421 VPB.n1231 VPB.n1228 1.794
R2422 VPB.n1294 VPB.n1291 1.794
R2423 VPB.n1357 VPB.n1354 1.794
R2424 VPB.n284 VPB.n281 1.435
R2425 VPB.n347 VPB.n344 1.435
R2426 VPB.n410 VPB.n407 1.435
R2427 VPB.n473 VPB.n470 1.435
R2428 VPB.n536 VPB.n533 1.435
R2429 VPB.n599 VPB.n596 1.435
R2430 VPB.n745 VPB.n742 1.435
R2431 VPB.n133 VPB.n132 1.435
R2432 VPB.n806 VPB.n803 1.435
R2433 VPB.n869 VPB.n866 1.435
R2434 VPB.n932 VPB.n929 1.435
R2435 VPB.n1078 VPB.n1075 1.435
R2436 VPB.n1141 VPB.n1138 1.435
R2437 VPB.n1204 VPB.n1201 1.435
R2438 VPB.n1267 VPB.n1264 1.435
R2439 VPB.n1330 VPB.n1327 1.435
R2440 VPB.n164 VPB.n155 1.402
R2441 VPB.n164 VPB.n158 1.402
R2442 VPB.n164 VPB.n162 1.402
R2443 VPB.n164 VPB.n163 1.402
R2444 VPB.n666 VPB.n663 1.076
R2445 VPB.n999 VPB.n996 1.076
R2446 VPB.n48 VPB.n45 1.076
R2447 VPB.n165 VPB.n164 0.735
R2448 VPB.n164 VPB.n154 0.735
R2449 VPB.n705 VPB.n702 0.717
R2450 VPB.n1038 VPB.n1035 0.717
R2451 VPB.n78 VPB.n77 0.717
R2452 VPB.n216 VPB.n215 0.387
R2453 VPB.n216 VPB.n211 0.387
R2454 VPB.n216 VPB.n206 0.387
R2455 VPB.n217 VPB.n216 0.387
R2456 VPB.n271 VPB.n270 0.387
R2457 VPB.n271 VPB.n266 0.387
R2458 VPB.n271 VPB.n261 0.387
R2459 VPB.n272 VPB.n271 0.387
R2460 VPB.n334 VPB.n333 0.387
R2461 VPB.n334 VPB.n329 0.387
R2462 VPB.n334 VPB.n324 0.387
R2463 VPB.n335 VPB.n334 0.387
R2464 VPB.n397 VPB.n396 0.387
R2465 VPB.n397 VPB.n392 0.387
R2466 VPB.n397 VPB.n387 0.387
R2467 VPB.n398 VPB.n397 0.387
R2468 VPB.n460 VPB.n459 0.387
R2469 VPB.n460 VPB.n455 0.387
R2470 VPB.n460 VPB.n450 0.387
R2471 VPB.n461 VPB.n460 0.387
R2472 VPB.n523 VPB.n522 0.387
R2473 VPB.n523 VPB.n518 0.387
R2474 VPB.n523 VPB.n513 0.387
R2475 VPB.n524 VPB.n523 0.387
R2476 VPB.n586 VPB.n585 0.387
R2477 VPB.n586 VPB.n581 0.387
R2478 VPB.n586 VPB.n576 0.387
R2479 VPB.n587 VPB.n586 0.387
R2480 VPB.n649 VPB.n648 0.387
R2481 VPB.n649 VPB.n644 0.387
R2482 VPB.n649 VPB.n639 0.387
R2483 VPB.n650 VPB.n649 0.387
R2484 VPB.n732 VPB.n731 0.387
R2485 VPB.n732 VPB.n727 0.387
R2486 VPB.n732 VPB.n722 0.387
R2487 VPB.n733 VPB.n732 0.387
R2488 VPB.n100 VPB.n99 0.387
R2489 VPB.n100 VPB.n95 0.387
R2490 VPB.n100 VPB.n90 0.387
R2491 VPB.n101 VPB.n100 0.387
R2492 VPB.n793 VPB.n792 0.387
R2493 VPB.n793 VPB.n788 0.387
R2494 VPB.n793 VPB.n783 0.387
R2495 VPB.n794 VPB.n793 0.387
R2496 VPB.n856 VPB.n855 0.387
R2497 VPB.n856 VPB.n851 0.387
R2498 VPB.n856 VPB.n846 0.387
R2499 VPB.n857 VPB.n856 0.387
R2500 VPB.n919 VPB.n918 0.387
R2501 VPB.n919 VPB.n914 0.387
R2502 VPB.n919 VPB.n909 0.387
R2503 VPB.n920 VPB.n919 0.387
R2504 VPB.n982 VPB.n981 0.387
R2505 VPB.n982 VPB.n977 0.387
R2506 VPB.n982 VPB.n972 0.387
R2507 VPB.n983 VPB.n982 0.387
R2508 VPB.n1065 VPB.n1064 0.387
R2509 VPB.n1065 VPB.n1060 0.387
R2510 VPB.n1065 VPB.n1055 0.387
R2511 VPB.n1066 VPB.n1065 0.387
R2512 VPB.n1128 VPB.n1127 0.387
R2513 VPB.n1128 VPB.n1123 0.387
R2514 VPB.n1128 VPB.n1118 0.387
R2515 VPB.n1129 VPB.n1128 0.387
R2516 VPB.n1191 VPB.n1190 0.387
R2517 VPB.n1191 VPB.n1186 0.387
R2518 VPB.n1191 VPB.n1181 0.387
R2519 VPB.n1192 VPB.n1191 0.387
R2520 VPB.n1254 VPB.n1253 0.387
R2521 VPB.n1254 VPB.n1249 0.387
R2522 VPB.n1254 VPB.n1244 0.387
R2523 VPB.n1255 VPB.n1254 0.387
R2524 VPB.n1317 VPB.n1316 0.387
R2525 VPB.n1317 VPB.n1312 0.387
R2526 VPB.n1317 VPB.n1307 0.387
R2527 VPB.n1318 VPB.n1317 0.387
R2528 VPB.n33 VPB.n32 0.387
R2529 VPB.n33 VPB.n28 0.387
R2530 VPB.n33 VPB.n23 0.387
R2531 VPB.n34 VPB.n33 0.387
R2532 VPB.n1382 VPB.n13 0.387
R2533 VPB.n1382 VPB.n9 0.387
R2534 VPB.n1382 VPB.n4 0.387
R2535 VPB.n1382 VPB.n1381 0.387
R2536 VPB.n225 VPB.n198 0.272
R2537 VPB.n280 VPB.n253 0.272
R2538 VPB.n343 VPB.n316 0.272
R2539 VPB.n406 VPB.n379 0.272
R2540 VPB.n469 VPB.n442 0.272
R2541 VPB.n532 VPB.n505 0.272
R2542 VPB.n595 VPB.n568 0.272
R2543 VPB.n658 VPB.n631 0.272
R2544 VPB.n741 VPB.n714 0.272
R2545 VPB.n757 VPB.n756 0.272
R2546 VPB.n802 VPB.n775 0.272
R2547 VPB.n865 VPB.n838 0.272
R2548 VPB.n928 VPB.n901 0.272
R2549 VPB.n991 VPB.n964 0.272
R2550 VPB.n1074 VPB.n1047 0.272
R2551 VPB.n1137 VPB.n1110 0.272
R2552 VPB.n1200 VPB.n1173 0.272
R2553 VPB.n1263 VPB.n1236 0.272
R2554 VPB.n1326 VPB.n1299 0.272
R2555 VPB.n1363 VPB.n1362 0.272
R2556 VPB.n1374 VPB 0.198
R2557 VPB.n182 VPB.n181 0.136
R2558 VPB.n186 VPB.n182 0.136
R2559 VPB.n190 VPB.n186 0.136
R2560 VPB.n194 VPB.n190 0.136
R2561 VPB.n198 VPB.n194 0.136
R2562 VPB.n229 VPB.n225 0.136
R2563 VPB.n233 VPB.n229 0.136
R2564 VPB.n237 VPB.n233 0.136
R2565 VPB.n241 VPB.n237 0.136
R2566 VPB.n245 VPB.n241 0.136
R2567 VPB.n249 VPB.n245 0.136
R2568 VPB.n253 VPB.n249 0.136
R2569 VPB.n285 VPB.n280 0.136
R2570 VPB.n290 VPB.n285 0.136
R2571 VPB.n297 VPB.n290 0.136
R2572 VPB.n302 VPB.n297 0.136
R2573 VPB.n307 VPB.n302 0.136
R2574 VPB.n312 VPB.n307 0.136
R2575 VPB.n316 VPB.n312 0.136
R2576 VPB.n348 VPB.n343 0.136
R2577 VPB.n353 VPB.n348 0.136
R2578 VPB.n360 VPB.n353 0.136
R2579 VPB.n365 VPB.n360 0.136
R2580 VPB.n370 VPB.n365 0.136
R2581 VPB.n375 VPB.n370 0.136
R2582 VPB.n379 VPB.n375 0.136
R2583 VPB.n411 VPB.n406 0.136
R2584 VPB.n416 VPB.n411 0.136
R2585 VPB.n423 VPB.n416 0.136
R2586 VPB.n428 VPB.n423 0.136
R2587 VPB.n433 VPB.n428 0.136
R2588 VPB.n438 VPB.n433 0.136
R2589 VPB.n442 VPB.n438 0.136
R2590 VPB.n474 VPB.n469 0.136
R2591 VPB.n479 VPB.n474 0.136
R2592 VPB.n486 VPB.n479 0.136
R2593 VPB.n491 VPB.n486 0.136
R2594 VPB.n496 VPB.n491 0.136
R2595 VPB.n501 VPB.n496 0.136
R2596 VPB.n505 VPB.n501 0.136
R2597 VPB.n537 VPB.n532 0.136
R2598 VPB.n542 VPB.n537 0.136
R2599 VPB.n549 VPB.n542 0.136
R2600 VPB.n554 VPB.n549 0.136
R2601 VPB.n559 VPB.n554 0.136
R2602 VPB.n564 VPB.n559 0.136
R2603 VPB.n568 VPB.n564 0.136
R2604 VPB.n600 VPB.n595 0.136
R2605 VPB.n605 VPB.n600 0.136
R2606 VPB.n612 VPB.n605 0.136
R2607 VPB.n617 VPB.n612 0.136
R2608 VPB.n622 VPB.n617 0.136
R2609 VPB.n627 VPB.n622 0.136
R2610 VPB.n631 VPB.n627 0.136
R2611 VPB.n662 VPB.n658 0.136
R2612 VPB.n667 VPB.n662 0.136
R2613 VPB.n672 VPB.n667 0.136
R2614 VPB.n679 VPB.n672 0.136
R2615 VPB.n684 VPB.n679 0.136
R2616 VPB.n689 VPB.n684 0.136
R2617 VPB.n696 VPB.n689 0.136
R2618 VPB.n701 VPB.n696 0.136
R2619 VPB.n706 VPB.n701 0.136
R2620 VPB.n710 VPB.n706 0.136
R2621 VPB.n714 VPB.n710 0.136
R2622 VPB.n746 VPB.n741 0.136
R2623 VPB.n751 VPB.n746 0.136
R2624 VPB.n752 VPB.n751 0.136
R2625 VPB.n753 VPB.n752 0.136
R2626 VPB.n754 VPB.n753 0.136
R2627 VPB.n755 VPB.n754 0.136
R2628 VPB.n756 VPB.n755 0.136
R2629 VPB.n758 VPB.n757 0.136
R2630 VPB.n759 VPB.n758 0.136
R2631 VPB.n760 VPB.n759 0.136
R2632 VPB.n761 VPB.n760 0.136
R2633 VPB.n762 VPB.n761 0.136
R2634 VPB.n775 VPB.n771 0.136
R2635 VPB.n807 VPB.n802 0.136
R2636 VPB.n812 VPB.n807 0.136
R2637 VPB.n819 VPB.n812 0.136
R2638 VPB.n824 VPB.n819 0.136
R2639 VPB.n829 VPB.n824 0.136
R2640 VPB.n834 VPB.n829 0.136
R2641 VPB.n838 VPB.n834 0.136
R2642 VPB.n870 VPB.n865 0.136
R2643 VPB.n875 VPB.n870 0.136
R2644 VPB.n882 VPB.n875 0.136
R2645 VPB.n887 VPB.n882 0.136
R2646 VPB.n892 VPB.n887 0.136
R2647 VPB.n897 VPB.n892 0.136
R2648 VPB.n901 VPB.n897 0.136
R2649 VPB.n933 VPB.n928 0.136
R2650 VPB.n938 VPB.n933 0.136
R2651 VPB.n945 VPB.n938 0.136
R2652 VPB.n950 VPB.n945 0.136
R2653 VPB.n955 VPB.n950 0.136
R2654 VPB.n960 VPB.n955 0.136
R2655 VPB.n964 VPB.n960 0.136
R2656 VPB.n995 VPB.n991 0.136
R2657 VPB.n1000 VPB.n995 0.136
R2658 VPB.n1005 VPB.n1000 0.136
R2659 VPB.n1012 VPB.n1005 0.136
R2660 VPB.n1017 VPB.n1012 0.136
R2661 VPB.n1022 VPB.n1017 0.136
R2662 VPB.n1029 VPB.n1022 0.136
R2663 VPB.n1034 VPB.n1029 0.136
R2664 VPB.n1039 VPB.n1034 0.136
R2665 VPB.n1043 VPB.n1039 0.136
R2666 VPB.n1047 VPB.n1043 0.136
R2667 VPB.n1079 VPB.n1074 0.136
R2668 VPB.n1084 VPB.n1079 0.136
R2669 VPB.n1091 VPB.n1084 0.136
R2670 VPB.n1096 VPB.n1091 0.136
R2671 VPB.n1101 VPB.n1096 0.136
R2672 VPB.n1106 VPB.n1101 0.136
R2673 VPB.n1110 VPB.n1106 0.136
R2674 VPB.n1142 VPB.n1137 0.136
R2675 VPB.n1147 VPB.n1142 0.136
R2676 VPB.n1154 VPB.n1147 0.136
R2677 VPB.n1159 VPB.n1154 0.136
R2678 VPB.n1164 VPB.n1159 0.136
R2679 VPB.n1169 VPB.n1164 0.136
R2680 VPB.n1173 VPB.n1169 0.136
R2681 VPB.n1205 VPB.n1200 0.136
R2682 VPB.n1210 VPB.n1205 0.136
R2683 VPB.n1217 VPB.n1210 0.136
R2684 VPB.n1222 VPB.n1217 0.136
R2685 VPB.n1227 VPB.n1222 0.136
R2686 VPB.n1232 VPB.n1227 0.136
R2687 VPB.n1236 VPB.n1232 0.136
R2688 VPB.n1268 VPB.n1263 0.136
R2689 VPB.n1273 VPB.n1268 0.136
R2690 VPB.n1280 VPB.n1273 0.136
R2691 VPB.n1285 VPB.n1280 0.136
R2692 VPB.n1290 VPB.n1285 0.136
R2693 VPB.n1295 VPB.n1290 0.136
R2694 VPB.n1299 VPB.n1295 0.136
R2695 VPB.n1331 VPB.n1326 0.136
R2696 VPB.n1336 VPB.n1331 0.136
R2697 VPB.n1343 VPB.n1336 0.136
R2698 VPB.n1348 VPB.n1343 0.136
R2699 VPB.n1353 VPB.n1348 0.136
R2700 VPB.n1358 VPB.n1353 0.136
R2701 VPB.n1362 VPB.n1358 0.136
R2702 VPB.n1364 VPB.n1363 0.136
R2703 VPB.n1365 VPB.n1364 0.136
R2704 VPB.n1366 VPB.n1365 0.136
R2705 VPB.n1367 VPB.n1366 0.136
R2706 VPB.n1368 VPB.n1367 0.136
R2707 VPB.n1369 VPB.n1368 0.136
R2708 VPB.n1370 VPB.n1369 0.136
R2709 VPB.n1371 VPB.n1370 0.136
R2710 VPB.n1372 VPB.n1371 0.136
R2711 VPB.n1373 VPB.n1372 0.136
R2712 VPB.n1374 VPB.n1373 0.136
R2713 VPB.n762 VPB 0.068
R2714 VPB.n771 VPB 0.068
R2715 a_13093_1005.n4 a_13093_1005.n3 195.987
R2716 a_13093_1005.n2 a_13093_1005.t0 89.553
R2717 a_13093_1005.n5 a_13093_1005.n4 75.27
R2718 a_13093_1005.n3 a_13093_1005.n2 75.214
R2719 a_13093_1005.n4 a_13093_1005.n0 36.519
R2720 a_13093_1005.n3 a_13093_1005.t4 14.338
R2721 a_13093_1005.n0 a_13093_1005.t7 14.282
R2722 a_13093_1005.n0 a_13093_1005.t6 14.282
R2723 a_13093_1005.n1 a_13093_1005.t5 14.282
R2724 a_13093_1005.n1 a_13093_1005.t3 14.282
R2725 a_13093_1005.n5 a_13093_1005.t1 14.282
R2726 a_13093_1005.t2 a_13093_1005.n5 14.282
R2727 a_13093_1005.n2 a_13093_1005.n1 12.119
R2728 a_147_159.n8 a_147_159.t6 512.525
R2729 a_147_159.n6 a_147_159.t5 472.359
R2730 a_147_159.n4 a_147_159.t7 472.359
R2731 a_147_159.n6 a_147_159.t8 384.527
R2732 a_147_159.n4 a_147_159.t10 384.527
R2733 a_147_159.n8 a_147_159.t11 371.139
R2734 a_147_159.n9 a_147_159.t13 324.268
R2735 a_147_159.n7 a_147_159.t9 277.772
R2736 a_147_159.n5 a_147_159.t12 277.772
R2737 a_147_159.n14 a_147_159.n12 247.192
R2738 a_147_159.n9 a_147_159.n8 119.654
R2739 a_147_159.n12 a_147_159.n3 109.441
R2740 a_147_159.n10 a_147_159.n9 82.484
R2741 a_147_159.n11 a_147_159.n5 80.307
R2742 a_147_159.n3 a_147_159.n2 76.002
R2743 a_147_159.n10 a_147_159.n7 76
R2744 a_147_159.n12 a_147_159.n11 76
R2745 a_147_159.n7 a_147_159.n6 67.001
R2746 a_147_159.n5 a_147_159.n4 67.001
R2747 a_147_159.n14 a_147_159.n13 30
R2748 a_147_159.n15 a_147_159.n0 24.383
R2749 a_147_159.n15 a_147_159.n14 23.684
R2750 a_147_159.n1 a_147_159.t4 14.282
R2751 a_147_159.n1 a_147_159.t3 14.282
R2752 a_147_159.n2 a_147_159.t0 14.282
R2753 a_147_159.n2 a_147_159.t1 14.282
R2754 a_147_159.n3 a_147_159.n1 12.85
R2755 a_147_159.n11 a_147_159.n10 2.947
R2756 a_1845_1004.n4 a_1845_1004.t5 480.392
R2757 a_1845_1004.n4 a_1845_1004.t6 403.272
R2758 a_1845_1004.n5 a_1845_1004.t7 266.974
R2759 a_1845_1004.n8 a_1845_1004.n6 194.086
R2760 a_1845_1004.n6 a_1845_1004.n3 162.547
R2761 a_1845_1004.n6 a_1845_1004.n5 153.315
R2762 a_1845_1004.n5 a_1845_1004.n4 108.494
R2763 a_1845_1004.n3 a_1845_1004.n2 76.002
R2764 a_1845_1004.n8 a_1845_1004.n7 30
R2765 a_1845_1004.n9 a_1845_1004.n0 24.383
R2766 a_1845_1004.n9 a_1845_1004.n8 23.684
R2767 a_1845_1004.n1 a_1845_1004.t2 14.282
R2768 a_1845_1004.n1 a_1845_1004.t1 14.282
R2769 a_1845_1004.n2 a_1845_1004.t3 14.282
R2770 a_1845_1004.n2 a_1845_1004.t4 14.282
R2771 a_1845_1004.n3 a_1845_1004.n1 12.85
R2772 a_4891_943.n4 a_4891_943.t9 480.392
R2773 a_4891_943.n6 a_4891_943.t6 454.685
R2774 a_4891_943.n6 a_4891_943.t8 428.979
R2775 a_4891_943.n4 a_4891_943.t5 403.272
R2776 a_4891_943.n5 a_4891_943.t7 266.974
R2777 a_4891_943.n7 a_4891_943.t10 221.453
R2778 a_4891_943.n11 a_4891_943.n9 194.086
R2779 a_4891_943.n9 a_4891_943.n3 162.547
R2780 a_4891_943.n7 a_4891_943.n6 108.494
R2781 a_4891_943.n5 a_4891_943.n4 108.494
R2782 a_4891_943.n8 a_4891_943.n7 78.947
R2783 a_4891_943.n8 a_4891_943.n5 77.315
R2784 a_4891_943.n3 a_4891_943.n2 76.002
R2785 a_4891_943.n9 a_4891_943.n8 76
R2786 a_4891_943.n11 a_4891_943.n10 30
R2787 a_4891_943.n12 a_4891_943.n0 24.383
R2788 a_4891_943.n12 a_4891_943.n11 23.684
R2789 a_4891_943.n1 a_4891_943.t3 14.282
R2790 a_4891_943.n1 a_4891_943.t2 14.282
R2791 a_4891_943.n2 a_4891_943.t1 14.282
R2792 a_4891_943.n2 a_4891_943.t0 14.282
R2793 a_4891_943.n3 a_4891_943.n1 12.85
R2794 a_6137_1004.n4 a_6137_1004.t5 480.392
R2795 a_6137_1004.n4 a_6137_1004.t6 403.272
R2796 a_6137_1004.n5 a_6137_1004.t7 266.974
R2797 a_6137_1004.n8 a_6137_1004.n6 194.086
R2798 a_6137_1004.n6 a_6137_1004.n3 162.547
R2799 a_6137_1004.n6 a_6137_1004.n5 153.315
R2800 a_6137_1004.n5 a_6137_1004.n4 108.494
R2801 a_6137_1004.n3 a_6137_1004.n2 76.002
R2802 a_6137_1004.n8 a_6137_1004.n7 30
R2803 a_6137_1004.n9 a_6137_1004.n0 24.383
R2804 a_6137_1004.n9 a_6137_1004.n8 23.684
R2805 a_6137_1004.n1 a_6137_1004.t0 14.282
R2806 a_6137_1004.n1 a_6137_1004.t1 14.282
R2807 a_6137_1004.n2 a_6137_1004.t3 14.282
R2808 a_6137_1004.n2 a_6137_1004.t4 14.282
R2809 a_6137_1004.n3 a_6137_1004.n1 12.85
R2810 a_4569_1004.n8 a_4569_1004.t7 480.392
R2811 a_4569_1004.n6 a_4569_1004.t10 480.392
R2812 a_4569_1004.n8 a_4569_1004.t11 403.272
R2813 a_4569_1004.n6 a_4569_1004.t12 403.272
R2814 a_4569_1004.n9 a_4569_1004.t8 293.527
R2815 a_4569_1004.n7 a_4569_1004.t9 293.527
R2816 a_4569_1004.n13 a_4569_1004.n11 223.151
R2817 a_4569_1004.n11 a_4569_1004.n5 154.293
R2818 a_4569_1004.n10 a_4569_1004.n7 83.3
R2819 a_4569_1004.n9 a_4569_1004.n8 81.941
R2820 a_4569_1004.n7 a_4569_1004.n6 81.941
R2821 a_4569_1004.n4 a_4569_1004.n3 79.232
R2822 a_4569_1004.n11 a_4569_1004.n10 77.315
R2823 a_4569_1004.n10 a_4569_1004.n9 76
R2824 a_4569_1004.n5 a_4569_1004.n4 63.152
R2825 a_4569_1004.n13 a_4569_1004.n12 30
R2826 a_4569_1004.n14 a_4569_1004.n0 24.383
R2827 a_4569_1004.n14 a_4569_1004.n13 23.684
R2828 a_4569_1004.n5 a_4569_1004.n1 16.08
R2829 a_4569_1004.n4 a_4569_1004.n2 16.08
R2830 a_4569_1004.n1 a_4569_1004.t2 14.282
R2831 a_4569_1004.n1 a_4569_1004.t3 14.282
R2832 a_4569_1004.n2 a_4569_1004.t6 14.282
R2833 a_4569_1004.n2 a_4569_1004.t5 14.282
R2834 a_4569_1004.n3 a_4569_1004.t1 14.282
R2835 a_4569_1004.n3 a_4569_1004.t0 14.282
R2836 a_13757_1005.n4 a_13757_1005.n3 196.002
R2837 a_13757_1005.n2 a_13757_1005.t1 89.553
R2838 a_13757_1005.n5 a_13757_1005.n4 75.27
R2839 a_13757_1005.n3 a_13757_1005.n2 75.214
R2840 a_13757_1005.n4 a_13757_1005.n0 36.52
R2841 a_13757_1005.n3 a_13757_1005.t4 14.338
R2842 a_13757_1005.n0 a_13757_1005.t2 14.282
R2843 a_13757_1005.n0 a_13757_1005.t7 14.282
R2844 a_13757_1005.n1 a_13757_1005.t0 14.282
R2845 a_13757_1005.n1 a_13757_1005.t3 14.282
R2846 a_13757_1005.t6 a_13757_1005.n5 14.282
R2847 a_13757_1005.n5 a_13757_1005.t5 14.282
R2848 a_13757_1005.n2 a_13757_1005.n1 12.119
R2849 a_7595_383.n5 a_7595_383.t5 475.572
R2850 a_7595_383.n9 a_7595_383.t7 472.359
R2851 a_7595_383.n4 a_7595_383.t6 469.145
R2852 a_7595_383.n9 a_7595_383.t12 384.527
R2853 a_7595_383.n5 a_7595_383.t11 384.527
R2854 a_7595_383.n4 a_7595_383.t10 384.527
R2855 a_7595_383.n6 a_7595_383.t13 277.772
R2856 a_7595_383.n12 a_7595_383.n3 242.205
R2857 a_7595_383.n10 a_7595_383.n9 201.031
R2858 a_7595_383.n7 a_7595_383.n6 156.851
R2859 a_7595_383.n10 a_7595_383.t9 141.018
R2860 a_7595_383.n8 a_7595_383.t8 141.018
R2861 a_7595_383.n8 a_7595_383.n7 134.03
R2862 a_7595_383.n14 a_7595_383.n12 114.428
R2863 a_7595_383.n3 a_7595_383.n2 76.002
R2864 a_7595_383.n12 a_7595_383.n11 76
R2865 a_7595_383.n6 a_7595_383.n5 67.889
R2866 a_7595_383.n11 a_7595_383.n8 66.982
R2867 a_7595_383.n7 a_7595_383.n4 66.88
R2868 a_7595_383.n11 a_7595_383.n10 52.291
R2869 a_7595_383.n14 a_7595_383.n13 30
R2870 a_7595_383.n15 a_7595_383.n0 24.383
R2871 a_7595_383.n15 a_7595_383.n14 23.684
R2872 a_7595_383.n1 a_7595_383.t1 14.282
R2873 a_7595_383.n1 a_7595_383.t0 14.282
R2874 a_7595_383.n2 a_7595_383.t3 14.282
R2875 a_7595_383.n2 a_7595_383.t4 14.282
R2876 a_7595_383.n3 a_7595_383.n1 12.85
R2877 a_277_1004.n7 a_277_1004.t8 480.392
R2878 a_277_1004.n5 a_277_1004.t11 480.392
R2879 a_277_1004.n7 a_277_1004.t12 403.272
R2880 a_277_1004.n5 a_277_1004.t7 403.272
R2881 a_277_1004.n8 a_277_1004.t9 293.527
R2882 a_277_1004.n6 a_277_1004.t10 293.527
R2883 a_277_1004.n12 a_277_1004.n10 229.673
R2884 a_277_1004.n10 a_277_1004.n4 154.293
R2885 a_277_1004.n9 a_277_1004.n6 83.3
R2886 a_277_1004.n8 a_277_1004.n7 81.941
R2887 a_277_1004.n6 a_277_1004.n5 81.941
R2888 a_277_1004.n3 a_277_1004.n2 79.232
R2889 a_277_1004.n10 a_277_1004.n9 77.315
R2890 a_277_1004.n9 a_277_1004.n8 76
R2891 a_277_1004.n4 a_277_1004.n3 63.152
R2892 a_277_1004.n4 a_277_1004.n0 16.08
R2893 a_277_1004.n3 a_277_1004.n1 16.08
R2894 a_277_1004.n12 a_277_1004.n11 15.218
R2895 a_277_1004.n0 a_277_1004.t0 14.282
R2896 a_277_1004.n0 a_277_1004.t1 14.282
R2897 a_277_1004.n1 a_277_1004.t5 14.282
R2898 a_277_1004.n1 a_277_1004.t4 14.282
R2899 a_277_1004.n2 a_277_1004.t3 14.282
R2900 a_277_1004.n2 a_277_1004.t2 14.282
R2901 a_277_1004.n13 a_277_1004.n12 12.014
R2902 a_8030_73.n12 a_8030_73.n11 26.811
R2903 a_8030_73.n6 a_8030_73.n5 24.977
R2904 a_8030_73.n2 a_8030_73.n1 24.877
R2905 a_8030_73.t0 a_8030_73.n2 12.677
R2906 a_8030_73.t0 a_8030_73.n3 11.595
R2907 a_8030_73.t1 a_8030_73.n8 8.137
R2908 a_8030_73.t0 a_8030_73.n4 7.273
R2909 a_8030_73.t0 a_8030_73.n0 6.109
R2910 a_8030_73.t1 a_8030_73.n7 4.864
R2911 a_8030_73.t0 a_8030_73.n12 2.074
R2912 a_8030_73.n7 a_8030_73.n6 1.13
R2913 a_8030_73.n12 a_8030_73.t1 0.937
R2914 a_8030_73.t1 a_8030_73.n10 0.804
R2915 a_8030_73.n10 a_8030_73.n9 0.136
R2916 a_8731_159.n7 a_8731_159.t5 512.525
R2917 a_8731_159.n5 a_8731_159.t7 472.359
R2918 a_8731_159.n3 a_8731_159.t12 472.359
R2919 a_8731_159.n5 a_8731_159.t13 384.527
R2920 a_8731_159.n3 a_8731_159.t6 384.527
R2921 a_8731_159.n7 a_8731_159.t10 371.139
R2922 a_8731_159.n8 a_8731_159.t9 324.268
R2923 a_8731_159.n6 a_8731_159.t8 277.772
R2924 a_8731_159.n4 a_8731_159.t11 277.772
R2925 a_8731_159.n13 a_8731_159.n11 253.714
R2926 a_8731_159.n8 a_8731_159.n7 119.654
R2927 a_8731_159.n11 a_8731_159.n2 109.441
R2928 a_8731_159.n9 a_8731_159.n8 82.484
R2929 a_8731_159.n10 a_8731_159.n4 80.307
R2930 a_8731_159.n2 a_8731_159.n1 76.002
R2931 a_8731_159.n9 a_8731_159.n6 76
R2932 a_8731_159.n11 a_8731_159.n10 76
R2933 a_8731_159.n6 a_8731_159.n5 67.001
R2934 a_8731_159.n4 a_8731_159.n3 67.001
R2935 a_8731_159.n13 a_8731_159.n12 15.218
R2936 a_8731_159.n0 a_8731_159.t3 14.282
R2937 a_8731_159.n0 a_8731_159.t4 14.282
R2938 a_8731_159.n1 a_8731_159.t0 14.282
R2939 a_8731_159.n1 a_8731_159.t1 14.282
R2940 a_8731_159.n2 a_8731_159.n0 12.85
R2941 a_8731_159.n14 a_8731_159.n13 12.014
R2942 a_8731_159.n10 a_8731_159.n9 2.947
R2943 a_8861_1004.n7 a_8861_1004.t12 480.392
R2944 a_8861_1004.n5 a_8861_1004.t10 480.392
R2945 a_8861_1004.n7 a_8861_1004.t7 403.272
R2946 a_8861_1004.n5 a_8861_1004.t8 403.272
R2947 a_8861_1004.n8 a_8861_1004.t9 293.527
R2948 a_8861_1004.n6 a_8861_1004.t11 293.527
R2949 a_8861_1004.n12 a_8861_1004.n10 229.673
R2950 a_8861_1004.n10 a_8861_1004.n4 154.293
R2951 a_8861_1004.n9 a_8861_1004.n6 83.3
R2952 a_8861_1004.n8 a_8861_1004.n7 81.941
R2953 a_8861_1004.n6 a_8861_1004.n5 81.941
R2954 a_8861_1004.n3 a_8861_1004.n2 79.232
R2955 a_8861_1004.n10 a_8861_1004.n9 77.315
R2956 a_8861_1004.n9 a_8861_1004.n8 76
R2957 a_8861_1004.n4 a_8861_1004.n3 63.152
R2958 a_8861_1004.n4 a_8861_1004.n0 16.08
R2959 a_8861_1004.n3 a_8861_1004.n1 16.08
R2960 a_8861_1004.n12 a_8861_1004.n11 15.218
R2961 a_8861_1004.n0 a_8861_1004.t3 14.282
R2962 a_8861_1004.n0 a_8861_1004.t4 14.282
R2963 a_8861_1004.n1 a_8861_1004.t6 14.282
R2964 a_8861_1004.n1 a_8861_1004.t5 14.282
R2965 a_8861_1004.n2 a_8861_1004.t1 14.282
R2966 a_8861_1004.n2 a_8861_1004.t0 14.282
R2967 a_8861_1004.n13 a_8861_1004.n12 12.014
R2968 a_5366_73.n12 a_5366_73.n11 26.811
R2969 a_5366_73.n6 a_5366_73.n5 24.977
R2970 a_5366_73.n2 a_5366_73.n1 24.877
R2971 a_5366_73.t0 a_5366_73.n2 12.677
R2972 a_5366_73.t0 a_5366_73.n3 11.595
R2973 a_5366_73.t1 a_5366_73.n8 8.137
R2974 a_5366_73.t0 a_5366_73.n4 7.273
R2975 a_5366_73.t0 a_5366_73.n0 6.109
R2976 a_5366_73.t1 a_5366_73.n7 4.864
R2977 a_5366_73.t0 a_5366_73.n12 2.074
R2978 a_5366_73.n7 a_5366_73.n6 1.13
R2979 a_5366_73.n12 a_5366_73.t1 0.937
R2980 a_5366_73.t1 a_5366_73.n10 0.804
R2981 a_5366_73.n10 a_5366_73.n9 0.136
R2982 a_599_943.n4 a_599_943.t7 480.392
R2983 a_599_943.n6 a_599_943.t8 454.685
R2984 a_599_943.n6 a_599_943.t6 428.979
R2985 a_599_943.n4 a_599_943.t10 403.272
R2986 a_599_943.n5 a_599_943.t5 266.974
R2987 a_599_943.n7 a_599_943.t9 221.453
R2988 a_599_943.n11 a_599_943.n9 194.086
R2989 a_599_943.n9 a_599_943.n3 162.547
R2990 a_599_943.n7 a_599_943.n6 108.494
R2991 a_599_943.n5 a_599_943.n4 108.494
R2992 a_599_943.n8 a_599_943.n7 78.947
R2993 a_599_943.n8 a_599_943.n5 77.315
R2994 a_599_943.n3 a_599_943.n2 76.002
R2995 a_599_943.n9 a_599_943.n8 76
R2996 a_599_943.n11 a_599_943.n10 30
R2997 a_599_943.n12 a_599_943.n0 24.383
R2998 a_599_943.n12 a_599_943.n11 23.684
R2999 a_599_943.n1 a_599_943.t2 14.282
R3000 a_599_943.n1 a_599_943.t1 14.282
R3001 a_599_943.n2 a_599_943.t4 14.282
R3002 a_599_943.n2 a_599_943.t3 14.282
R3003 a_599_943.n3 a_599_943.n1 12.85
R3004 a_1740_73.n12 a_1740_73.n11 26.811
R3005 a_1740_73.n6 a_1740_73.n5 24.977
R3006 a_1740_73.n2 a_1740_73.n1 24.877
R3007 a_1740_73.t0 a_1740_73.n2 12.677
R3008 a_1740_73.t0 a_1740_73.n3 11.595
R3009 a_1740_73.t1 a_1740_73.n8 8.137
R3010 a_1740_73.t0 a_1740_73.n4 7.273
R3011 a_1740_73.t0 a_1740_73.n0 6.109
R3012 a_1740_73.t1 a_1740_73.n7 4.864
R3013 a_1740_73.t0 a_1740_73.n12 2.074
R3014 a_1740_73.n7 a_1740_73.n6 1.13
R3015 a_1740_73.n12 a_1740_73.t1 0.937
R3016 a_1740_73.t1 a_1740_73.n10 0.804
R3017 a_1740_73.n10 a_1740_73.n9 0.136
R3018 a_3177_1004.n3 a_3177_1004.t7 480.392
R3019 a_3177_1004.n3 a_3177_1004.t6 403.272
R3020 a_3177_1004.n4 a_3177_1004.t5 293.527
R3021 a_3177_1004.n7 a_3177_1004.n5 227.161
R3022 a_3177_1004.n5 a_3177_1004.n4 153.315
R3023 a_3177_1004.n5 a_3177_1004.n2 135.994
R3024 a_3177_1004.n4 a_3177_1004.n3 81.941
R3025 a_3177_1004.n2 a_3177_1004.n1 76.002
R3026 a_3177_1004.n7 a_3177_1004.n6 15.218
R3027 a_3177_1004.n0 a_3177_1004.t4 14.282
R3028 a_3177_1004.n0 a_3177_1004.t0 14.282
R3029 a_3177_1004.n1 a_3177_1004.t2 14.282
R3030 a_3177_1004.n1 a_3177_1004.t3 14.282
R3031 a_3177_1004.n2 a_3177_1004.n0 12.85
R3032 a_3177_1004.n8 a_3177_1004.n7 12.014
R3033 a_11761_1004.n4 a_11761_1004.t7 480.392
R3034 a_11761_1004.n4 a_11761_1004.t5 403.272
R3035 a_11761_1004.n5 a_11761_1004.t6 346.633
R3036 a_11761_1004.n8 a_11761_1004.n6 273.745
R3037 a_11761_1004.n6 a_11761_1004.n5 153.315
R3038 a_11761_1004.n6 a_11761_1004.n3 82.888
R3039 a_11761_1004.n3 a_11761_1004.n2 76.002
R3040 a_11761_1004.n8 a_11761_1004.n7 30
R3041 a_11761_1004.n5 a_11761_1004.n4 28.835
R3042 a_11761_1004.n9 a_11761_1004.n0 24.383
R3043 a_11761_1004.n9 a_11761_1004.n8 23.684
R3044 a_11761_1004.n1 a_11761_1004.t1 14.282
R3045 a_11761_1004.n1 a_11761_1004.t0 14.282
R3046 a_11761_1004.n2 a_11761_1004.t3 14.282
R3047 a_11761_1004.n2 a_11761_1004.t4 14.282
R3048 a_11761_1004.n3 a_11761_1004.n1 12.85
R3049 a_9183_943.n4 a_9183_943.t7 480.392
R3050 a_9183_943.n6 a_9183_943.t8 454.685
R3051 a_9183_943.n6 a_9183_943.t10 428.979
R3052 a_9183_943.n4 a_9183_943.t9 403.272
R3053 a_9183_943.n5 a_9183_943.t5 266.974
R3054 a_9183_943.n7 a_9183_943.t6 221.453
R3055 a_9183_943.n11 a_9183_943.n9 194.086
R3056 a_9183_943.n9 a_9183_943.n3 162.547
R3057 a_9183_943.n7 a_9183_943.n6 108.494
R3058 a_9183_943.n5 a_9183_943.n4 108.494
R3059 a_9183_943.n8 a_9183_943.n7 78.947
R3060 a_9183_943.n8 a_9183_943.n5 77.315
R3061 a_9183_943.n3 a_9183_943.n2 76.002
R3062 a_9183_943.n9 a_9183_943.n8 76
R3063 a_9183_943.n11 a_9183_943.n10 30
R3064 a_9183_943.n12 a_9183_943.n0 24.383
R3065 a_9183_943.n12 a_9183_943.n11 23.684
R3066 a_9183_943.n1 a_9183_943.t2 14.282
R3067 a_9183_943.n1 a_9183_943.t1 14.282
R3068 a_9183_943.n2 a_9183_943.t3 14.282
R3069 a_9183_943.n2 a_9183_943.t4 14.282
R3070 a_9183_943.n3 a_9183_943.n1 12.85
R3071 a_91_75.n4 a_91_75.n3 19.724
R3072 a_91_75.t0 a_91_75.n5 11.595
R3073 a_91_75.t0 a_91_75.n4 9.207
R3074 a_91_75.n2 a_91_75.n0 8.543
R3075 a_91_75.t0 a_91_75.n2 3.034
R3076 a_91_75.n2 a_91_75.n1 0.443
R3077 a_372_182.n8 a_372_182.n6 96.467
R3078 a_372_182.n3 a_372_182.n1 44.628
R3079 a_372_182.t0 a_372_182.n8 32.417
R3080 a_372_182.n3 a_372_182.n2 23.284
R3081 a_372_182.n6 a_372_182.n5 22.349
R3082 a_372_182.t0 a_372_182.n10 20.241
R3083 a_372_182.n10 a_372_182.n9 13.494
R3084 a_372_182.n6 a_372_182.n4 8.443
R3085 a_372_182.t0 a_372_182.n0 8.137
R3086 a_372_182.t0 a_372_182.n3 5.727
R3087 a_372_182.n8 a_372_182.n7 1.435
R3088 a_13654_73.n2 a_13654_73.n0 34.606
R3089 a_13654_73.n2 a_13654_73.n1 2.115
R3090 a_13654_73.t0 a_13654_73.n2 0.065
R3091 a_12988_73.n1 a_12988_73.n0 32.249
R3092 a_12988_73.t0 a_12988_73.n5 7.911
R3093 a_12988_73.n4 a_12988_73.n2 4.032
R3094 a_12988_73.n4 a_12988_73.n3 3.644
R3095 a_12988_73.t0 a_12988_73.n1 2.534
R3096 a_12988_73.t0 a_12988_73.n4 1.099
R3097 a_7469_1004.n4 a_7469_1004.t5 480.392
R3098 a_7469_1004.n4 a_7469_1004.t6 403.272
R3099 a_7469_1004.n5 a_7469_1004.t7 293.527
R3100 a_7469_1004.n8 a_7469_1004.n6 220.639
R3101 a_7469_1004.n6 a_7469_1004.n5 153.315
R3102 a_7469_1004.n6 a_7469_1004.n3 135.994
R3103 a_7469_1004.n5 a_7469_1004.n4 81.941
R3104 a_7469_1004.n3 a_7469_1004.n2 76.002
R3105 a_7469_1004.n8 a_7469_1004.n7 30
R3106 a_7469_1004.n9 a_7469_1004.n0 24.383
R3107 a_7469_1004.n9 a_7469_1004.n8 23.684
R3108 a_7469_1004.n1 a_7469_1004.t4 14.282
R3109 a_7469_1004.n1 a_7469_1004.t3 14.282
R3110 a_7469_1004.n2 a_7469_1004.t1 14.282
R3111 a_7469_1004.n2 a_7469_1004.t0 14.282
R3112 a_7469_1004.n3 a_7469_1004.n1 12.85
R3113 a_2406_73.n12 a_2406_73.n11 26.811
R3114 a_2406_73.n6 a_2406_73.n5 24.977
R3115 a_2406_73.n2 a_2406_73.n1 24.877
R3116 a_2406_73.t0 a_2406_73.n2 12.677
R3117 a_2406_73.t0 a_2406_73.n3 11.595
R3118 a_2406_73.t1 a_2406_73.n8 8.137
R3119 a_2406_73.t0 a_2406_73.n4 7.273
R3120 a_2406_73.t0 a_2406_73.n0 6.109
R3121 a_2406_73.t1 a_2406_73.n7 4.864
R3122 a_2406_73.t0 a_2406_73.n12 2.074
R3123 a_2406_73.n7 a_2406_73.n6 1.13
R3124 a_2406_73.n12 a_2406_73.t1 0.937
R3125 a_2406_73.t1 a_2406_73.n10 0.804
R3126 a_2406_73.n10 a_2406_73.n9 0.136
R3127 a_4664_182.n8 a_4664_182.n6 96.467
R3128 a_4664_182.n3 a_4664_182.n1 44.628
R3129 a_4664_182.t0 a_4664_182.n8 32.417
R3130 a_4664_182.n3 a_4664_182.n2 23.284
R3131 a_4664_182.n6 a_4664_182.n5 22.349
R3132 a_4664_182.t0 a_4664_182.n10 20.241
R3133 a_4664_182.n10 a_4664_182.n9 13.494
R3134 a_4664_182.n6 a_4664_182.n4 8.443
R3135 a_4664_182.t0 a_4664_182.n0 8.137
R3136 a_4664_182.t0 a_4664_182.n3 5.727
R3137 a_4664_182.n8 a_4664_182.n7 1.435
R3138 a_9658_73.t0 a_9658_73.n1 34.62
R3139 a_9658_73.t0 a_9658_73.n0 8.137
R3140 a_9658_73.t0 a_9658_73.n2 4.69
R3141 a_13268_181.n11 a_13268_181.n3 336.934
R3142 a_13268_181.n10 a_13268_181.n9 114.024
R3143 a_13268_181.n10 a_13268_181.n6 111.94
R3144 a_13268_181.n11 a_13268_181.n10 78.403
R3145 a_13268_181.n3 a_13268_181.n2 75.271
R3146 a_13268_181.n14 a_13268_181.n0 55.263
R3147 a_13268_181.n13 a_13268_181.n12 30
R3148 a_13268_181.n14 a_13268_181.n13 25.263
R3149 a_13268_181.n6 a_13268_181.n5 22.578
R3150 a_13268_181.n9 a_13268_181.n8 22.578
R3151 a_13268_181.n13 a_13268_181.n11 20.417
R3152 a_13268_181.n1 a_13268_181.t5 14.282
R3153 a_13268_181.n1 a_13268_181.t4 14.282
R3154 a_13268_181.n2 a_13268_181.t0 14.282
R3155 a_13268_181.n2 a_13268_181.t1 14.282
R3156 a_13268_181.n3 a_13268_181.n1 12.119
R3157 a_13268_181.n6 a_13268_181.n4 8.58
R3158 a_13268_181.n9 a_13268_181.n7 8.58
R3159 a_3303_383.n5 a_3303_383.t6 512.525
R3160 a_3303_383.n4 a_3303_383.t10 512.525
R3161 a_3303_383.n9 a_3303_383.t12 472.359
R3162 a_3303_383.n9 a_3303_383.t5 384.527
R3163 a_3303_383.n5 a_3303_383.t11 371.139
R3164 a_3303_383.n4 a_3303_383.t7 371.139
R3165 a_3303_383.n6 a_3303_383.n5 258.98
R3166 a_3303_383.n10 a_3303_383.t13 198.113
R3167 a_3303_383.n8 a_3303_383.n4 195.827
R3168 a_3303_383.n12 a_3303_383.n3 189.099
R3169 a_3303_383.n6 a_3303_383.t9 176.995
R3170 a_3303_383.n7 a_3303_383.t8 170.569
R3171 a_3303_383.n14 a_3303_383.n12 167.533
R3172 a_3303_383.n7 a_3303_383.n6 153.043
R3173 a_3303_383.n10 a_3303_383.n9 146.66
R3174 a_3303_383.n11 a_3303_383.n8 112.41
R3175 a_3303_383.n11 a_3303_383.n10 78.947
R3176 a_3303_383.n3 a_3303_383.n2 76.002
R3177 a_3303_383.n12 a_3303_383.n11 76
R3178 a_3303_383.n8 a_3303_383.n7 63.152
R3179 a_3303_383.n14 a_3303_383.n13 30
R3180 a_3303_383.n15 a_3303_383.n0 24.383
R3181 a_3303_383.n15 a_3303_383.n14 23.684
R3182 a_3303_383.n1 a_3303_383.t3 14.282
R3183 a_3303_383.n1 a_3303_383.t2 14.282
R3184 a_3303_383.n2 a_3303_383.t0 14.282
R3185 a_3303_383.n2 a_3303_383.t1 14.282
R3186 a_3303_383.n3 a_3303_383.n1 12.85
R3187 a_7364_73.n12 a_7364_73.n11 26.811
R3188 a_7364_73.n6 a_7364_73.n5 24.977
R3189 a_7364_73.n2 a_7364_73.n1 24.877
R3190 a_7364_73.t0 a_7364_73.n2 12.677
R3191 a_7364_73.t0 a_7364_73.n3 11.595
R3192 a_7364_73.t1 a_7364_73.n8 8.137
R3193 a_7364_73.t0 a_7364_73.n4 7.273
R3194 a_7364_73.t0 a_7364_73.n0 6.109
R3195 a_7364_73.t1 a_7364_73.n7 4.864
R3196 a_7364_73.t0 a_7364_73.n12 2.074
R3197 a_7364_73.n7 a_7364_73.n6 1.13
R3198 a_7364_73.n12 a_7364_73.t1 0.937
R3199 a_7364_73.t1 a_7364_73.n10 0.804
R3200 a_7364_73.n10 a_7364_73.n9 0.136
R3201 a_3738_73.n12 a_3738_73.n11 26.811
R3202 a_3738_73.n6 a_3738_73.n5 24.977
R3203 a_3738_73.n2 a_3738_73.n1 24.877
R3204 a_3738_73.t0 a_3738_73.n2 12.677
R3205 a_3738_73.t0 a_3738_73.n3 11.595
R3206 a_3738_73.t1 a_3738_73.n8 8.137
R3207 a_3738_73.t0 a_3738_73.n4 7.273
R3208 a_3738_73.t0 a_3738_73.n0 6.109
R3209 a_3738_73.t1 a_3738_73.n7 4.864
R3210 a_3738_73.t0 a_3738_73.n12 2.074
R3211 a_3738_73.n7 a_3738_73.n6 1.13
R3212 a_3738_73.n12 a_3738_73.t1 0.937
R3213 a_3738_73.t1 a_3738_73.n10 0.804
R3214 a_3738_73.n10 a_3738_73.n9 0.136
R3215 a_10324_73.t0 a_10324_73.n1 34.62
R3216 a_10324_73.t0 a_10324_73.n0 8.137
R3217 a_10324_73.t0 a_10324_73.n2 4.69
R3218 a_8956_182.n9 a_8956_182.n7 82.852
R3219 a_8956_182.n3 a_8956_182.n1 44.628
R3220 a_8956_182.t0 a_8956_182.n9 32.417
R3221 a_8956_182.n7 a_8956_182.n6 27.2
R3222 a_8956_182.n5 a_8956_182.n4 23.498
R3223 a_8956_182.n3 a_8956_182.n2 23.284
R3224 a_8956_182.n7 a_8956_182.n5 22.4
R3225 a_8956_182.t0 a_8956_182.n11 20.241
R3226 a_8956_182.n11 a_8956_182.n10 13.494
R3227 a_8956_182.t0 a_8956_182.n0 8.137
R3228 a_8956_182.t0 a_8956_182.n3 5.727
R3229 a_8956_182.n9 a_8956_182.n8 1.435
R3230 a_11656_73.t0 a_11656_73.n1 34.62
R3231 a_11656_73.t0 a_11656_73.n0 8.137
R3232 a_11656_73.t0 a_11656_73.n2 4.69
R3233 a_1074_73.t0 a_1074_73.n1 34.62
R3234 a_1074_73.t0 a_1074_73.n0 8.137
R3235 a_1074_73.t0 a_1074_73.n2 4.69
R3236 a_12322_73.t0 a_12322_73.n1 34.62
R3237 a_12322_73.t0 a_12322_73.n0 8.137
R3238 a_12322_73.t0 a_12322_73.n2 4.69
R3239 a_6698_73.n12 a_6698_73.n11 26.811
R3240 a_6698_73.n6 a_6698_73.n5 24.977
R3241 a_6698_73.n2 a_6698_73.n1 24.877
R3242 a_6698_73.t0 a_6698_73.n2 12.677
R3243 a_6698_73.t0 a_6698_73.n3 11.595
R3244 a_6698_73.t1 a_6698_73.n8 8.137
R3245 a_6698_73.t0 a_6698_73.n4 7.273
R3246 a_6698_73.t0 a_6698_73.n0 6.109
R3247 a_6698_73.t1 a_6698_73.n7 4.864
R3248 a_6698_73.t0 a_6698_73.n12 2.074
R3249 a_6698_73.n7 a_6698_73.n6 1.13
R3250 a_6698_73.n12 a_6698_73.t1 0.937
R3251 a_6698_73.t1 a_6698_73.n10 0.804
R3252 a_6698_73.n10 a_6698_73.n9 0.136
R3253 a_3072_73.t0 a_3072_73.n1 34.62
R3254 a_3072_73.t0 a_3072_73.n0 8.137
R3255 a_3072_73.t0 a_3072_73.n2 4.69
R3256 a_6032_73.t0 a_6032_73.n1 34.62
R3257 a_6032_73.t0 a_6032_73.n0 8.137
R3258 a_6032_73.t0 a_6032_73.n2 4.69
R3259 a_14320_73.t0 a_14320_73.n1 34.62
R3260 a_14320_73.t0 a_14320_73.n0 8.137
R3261 a_14320_73.t0 a_14320_73.n2 4.69
R3262 a_8675_75.n5 a_8675_75.n4 19.724
R3263 a_8675_75.t0 a_8675_75.n3 11.595
R3264 a_8675_75.t0 a_8675_75.n5 9.207
R3265 a_8675_75.n2 a_8675_75.n1 2.455
R3266 a_8675_75.n2 a_8675_75.n0 1.32
R3267 a_8675_75.t0 a_8675_75.n2 0.246
C3 VPB VNB 56.35fF
C4 a_8675_75.n0 VNB 0.10fF
C5 a_8675_75.n1 VNB 0.04fF
C6 a_8675_75.n2 VNB 0.03fF
C7 a_8675_75.n3 VNB 0.07fF
C8 a_8675_75.n4 VNB 0.08fF
C9 a_8675_75.n5 VNB 0.06fF
C10 a_14320_73.n0 VNB 0.06fF
C11 a_14320_73.n1 VNB 0.13fF
C12 a_14320_73.n2 VNB 0.04fF
C13 a_6032_73.n0 VNB 0.05fF
C14 a_6032_73.n1 VNB 0.12fF
C15 a_6032_73.n2 VNB 0.04fF
C16 a_3072_73.n0 VNB 0.05fF
C17 a_3072_73.n1 VNB 0.12fF
C18 a_3072_73.n2 VNB 0.04fF
C19 a_6698_73.n0 VNB 0.02fF
C20 a_6698_73.n1 VNB 0.10fF
C21 a_6698_73.n2 VNB 0.06fF
C22 a_6698_73.n3 VNB 0.06fF
C23 a_6698_73.n4 VNB 0.00fF
C24 a_6698_73.n5 VNB 0.04fF
C25 a_6698_73.n6 VNB 0.05fF
C26 a_6698_73.n7 VNB 0.02fF
C27 a_6698_73.n8 VNB 0.05fF
C28 a_6698_73.n9 VNB 0.08fF
C29 a_6698_73.n10 VNB 0.17fF
C30 a_6698_73.t1 VNB 0.23fF
C31 a_6698_73.n11 VNB 0.09fF
C32 a_6698_73.n12 VNB 0.00fF
C33 a_12322_73.n0 VNB 0.05fF
C34 a_12322_73.n1 VNB 0.12fF
C35 a_12322_73.n2 VNB 0.04fF
C36 a_1074_73.n0 VNB 0.05fF
C37 a_1074_73.n1 VNB 0.12fF
C38 a_1074_73.n2 VNB 0.04fF
C39 a_11656_73.n0 VNB 0.05fF
C40 a_11656_73.n1 VNB 0.12fF
C41 a_11656_73.n2 VNB 0.04fF
C42 a_8956_182.n0 VNB 0.07fF
C43 a_8956_182.n1 VNB 0.09fF
C44 a_8956_182.n2 VNB 0.13fF
C45 a_8956_182.n3 VNB 0.11fF
C46 a_8956_182.n4 VNB 0.02fF
C47 a_8956_182.n5 VNB 0.03fF
C48 a_8956_182.n6 VNB 0.02fF
C49 a_8956_182.n7 VNB 0.05fF
C50 a_8956_182.n8 VNB 0.03fF
C51 a_8956_182.n9 VNB 0.11fF
C52 a_8956_182.n10 VNB 0.06fF
C53 a_8956_182.n11 VNB 0.01fF
C54 a_8956_182.t0 VNB 0.33fF
C55 a_10324_73.n0 VNB 0.05fF
C56 a_10324_73.n1 VNB 0.12fF
C57 a_10324_73.n2 VNB 0.04fF
C58 a_3738_73.n0 VNB 0.02fF
C59 a_3738_73.n1 VNB 0.10fF
C60 a_3738_73.n2 VNB 0.06fF
C61 a_3738_73.n3 VNB 0.06fF
C62 a_3738_73.n4 VNB 0.00fF
C63 a_3738_73.n5 VNB 0.04fF
C64 a_3738_73.n6 VNB 0.05fF
C65 a_3738_73.n7 VNB 0.02fF
C66 a_3738_73.n8 VNB 0.05fF
C67 a_3738_73.n9 VNB 0.08fF
C68 a_3738_73.n10 VNB 0.17fF
C69 a_3738_73.t1 VNB 0.23fF
C70 a_3738_73.n11 VNB 0.09fF
C71 a_3738_73.n12 VNB 0.00fF
C72 a_7364_73.n0 VNB 0.02fF
C73 a_7364_73.n1 VNB 0.10fF
C74 a_7364_73.n2 VNB 0.06fF
C75 a_7364_73.n3 VNB 0.06fF
C76 a_7364_73.n4 VNB 0.00fF
C77 a_7364_73.n5 VNB 0.04fF
C78 a_7364_73.n6 VNB 0.05fF
C79 a_7364_73.n7 VNB 0.02fF
C80 a_7364_73.n8 VNB 0.05fF
C81 a_7364_73.n9 VNB 0.08fF
C82 a_7364_73.n10 VNB 0.17fF
C83 a_7364_73.t1 VNB 0.23fF
C84 a_7364_73.n11 VNB 0.09fF
C85 a_7364_73.n12 VNB 0.00fF
C86 a_3303_383.n0 VNB 0.08fF
C87 a_3303_383.n1 VNB 1.00fF
C88 a_3303_383.n2 VNB 1.18fF
C89 a_3303_383.n3 VNB 0.66fF
C90 a_3303_383.n4 VNB 0.74fF
C91 a_3303_383.n5 VNB 0.88fF
C92 a_3303_383.n6 VNB 1.08fF
C93 a_3303_383.t8 VNB 0.83fF
C94 a_3303_383.n7 VNB 0.65fF
C95 a_3303_383.n8 VNB 3.06fF
C96 a_3303_383.n9 VNB 0.71fF
C97 a_3303_383.t13 VNB 0.92fF
C98 a_3303_383.n10 VNB 0.72fF
C99 a_3303_383.n11 VNB 14.13fF
C100 a_3303_383.n12 VNB 0.79fF
C101 a_3303_383.n13 VNB 0.06fF
C102 a_3303_383.n14 VNB 0.47fF
C103 a_3303_383.n15 VNB 0.10fF
C104 a_13268_181.n0 VNB 0.04fF
C105 a_13268_181.n1 VNB 0.42fF
C106 a_13268_181.n2 VNB 0.51fF
C107 a_13268_181.n3 VNB 0.48fF
C108 a_13268_181.n4 VNB 0.04fF
C109 a_13268_181.n5 VNB 0.05fF
C110 a_13268_181.n6 VNB 0.11fF
C111 a_13268_181.n7 VNB 0.04fF
C112 a_13268_181.n8 VNB 0.05fF
C113 a_13268_181.n9 VNB 0.11fF
C114 a_13268_181.n10 VNB 1.11fF
C115 a_13268_181.n11 VNB 0.41fF
C116 a_13268_181.n12 VNB 0.03fF
C117 a_13268_181.n13 VNB 0.05fF
C118 a_13268_181.n14 VNB 0.04fF
C119 a_9658_73.n0 VNB 0.05fF
C120 a_9658_73.n1 VNB 0.12fF
C121 a_9658_73.n2 VNB 0.04fF
C122 a_4664_182.n0 VNB 0.07fF
C123 a_4664_182.n1 VNB 0.09fF
C124 a_4664_182.n2 VNB 0.13fF
C125 a_4664_182.n3 VNB 0.11fF
C126 a_4664_182.n4 VNB 0.02fF
C127 a_4664_182.n5 VNB 0.03fF
C128 a_4664_182.n6 VNB 0.06fF
C129 a_4664_182.n7 VNB 0.03fF
C130 a_4664_182.n8 VNB 0.12fF
C131 a_4664_182.n9 VNB 0.06fF
C132 a_4664_182.n10 VNB 0.01fF
C133 a_4664_182.t0 VNB 0.33fF
C134 a_2406_73.n0 VNB 0.02fF
C135 a_2406_73.n1 VNB 0.10fF
C136 a_2406_73.n2 VNB 0.06fF
C137 a_2406_73.n3 VNB 0.06fF
C138 a_2406_73.n4 VNB 0.00fF
C139 a_2406_73.n5 VNB 0.04fF
C140 a_2406_73.n6 VNB 0.05fF
C141 a_2406_73.n7 VNB 0.02fF
C142 a_2406_73.n8 VNB 0.05fF
C143 a_2406_73.n9 VNB 0.08fF
C144 a_2406_73.n10 VNB 0.17fF
C145 a_2406_73.t1 VNB 0.23fF
C146 a_2406_73.n11 VNB 0.09fF
C147 a_2406_73.n12 VNB 0.00fF
C148 a_7469_1004.n0 VNB 0.04fF
C149 a_7469_1004.n1 VNB 0.57fF
C150 a_7469_1004.n2 VNB 0.67fF
C151 a_7469_1004.n3 VNB 0.31fF
C152 a_7469_1004.n4 VNB 0.38fF
C153 a_7469_1004.n5 VNB 0.61fF
C154 a_7469_1004.n6 VNB 0.64fF
C155 a_7469_1004.n7 VNB 0.04fF
C156 a_7469_1004.n8 VNB 0.33fF
C157 a_7469_1004.n9 VNB 0.06fF
C158 a_12988_73.n0 VNB 0.11fF
C159 a_12988_73.n1 VNB 0.09fF
C160 a_12988_73.n2 VNB 0.08fF
C161 a_12988_73.n3 VNB 0.02fF
C162 a_12988_73.n4 VNB 0.01fF
C163 a_12988_73.n5 VNB 0.06fF
C164 a_13654_73.n0 VNB 0.13fF
C165 a_13654_73.n1 VNB 0.14fF
C166 a_13654_73.n2 VNB 0.16fF
C167 a_372_182.n0 VNB 0.07fF
C168 a_372_182.n1 VNB 0.09fF
C169 a_372_182.n2 VNB 0.13fF
C170 a_372_182.n3 VNB 0.11fF
C171 a_372_182.n4 VNB 0.02fF
C172 a_372_182.n5 VNB 0.03fF
C173 a_372_182.n6 VNB 0.06fF
C174 a_372_182.n7 VNB 0.03fF
C175 a_372_182.n8 VNB 0.12fF
C176 a_372_182.n9 VNB 0.06fF
C177 a_372_182.n10 VNB 0.01fF
C178 a_372_182.t0 VNB 0.33fF
C179 a_91_75.n0 VNB 0.19fF
C180 a_91_75.n1 VNB 0.04fF
C181 a_91_75.n2 VNB 0.01fF
C182 a_91_75.n3 VNB 0.08fF
C183 a_91_75.n4 VNB 0.06fF
C184 a_91_75.n5 VNB 0.06fF
C185 a_9183_943.n0 VNB 0.05fF
C186 a_9183_943.n1 VNB 0.72fF
C187 a_9183_943.n2 VNB 0.85fF
C188 a_9183_943.n3 VNB 0.43fF
C189 a_9183_943.n4 VNB 0.53fF
C190 a_9183_943.n5 VNB 0.53fF
C191 a_9183_943.n6 VNB 0.53fF
C192 a_9183_943.t6 VNB 0.70fF
C193 a_9183_943.n7 VNB 0.51fF
C194 a_9183_943.n8 VNB 1.39fF
C195 a_9183_943.n9 VNB 0.57fF
C196 a_9183_943.n10 VNB 0.05fF
C197 a_9183_943.n11 VNB 0.38fF
C198 a_9183_943.n12 VNB 0.07fF
C199 a_11761_1004.n0 VNB 0.04fF
C200 a_11761_1004.n1 VNB 0.53fF
C201 a_11761_1004.n2 VNB 0.63fF
C202 a_11761_1004.n3 VNB 0.23fF
C203 a_11761_1004.n4 VNB 0.29fF
C204 a_11761_1004.n5 VNB 0.58fF
C205 a_11761_1004.n6 VNB 0.60fF
C206 a_11761_1004.n7 VNB 0.03fF
C207 a_11761_1004.n8 VNB 0.37fF
C208 a_11761_1004.n9 VNB 0.05fF
C209 a_3177_1004.n0 VNB 0.55fF
C210 a_3177_1004.n1 VNB 0.65fF
C211 a_3177_1004.n2 VNB 0.30fF
C212 a_3177_1004.n3 VNB 0.37fF
C213 a_3177_1004.n4 VNB 0.59fF
C214 a_3177_1004.n5 VNB 0.63fF
C215 a_3177_1004.n6 VNB 0.09fF
C216 a_3177_1004.n7 VNB 0.31fF
C217 a_3177_1004.n8 VNB 0.05fF
C218 a_1740_73.n0 VNB 0.02fF
C219 a_1740_73.n1 VNB 0.10fF
C220 a_1740_73.n2 VNB 0.06fF
C221 a_1740_73.n3 VNB 0.06fF
C222 a_1740_73.n4 VNB 0.00fF
C223 a_1740_73.n5 VNB 0.04fF
C224 a_1740_73.n6 VNB 0.05fF
C225 a_1740_73.n7 VNB 0.02fF
C226 a_1740_73.n8 VNB 0.05fF
C227 a_1740_73.n9 VNB 0.08fF
C228 a_1740_73.n10 VNB 0.17fF
C229 a_1740_73.t1 VNB 0.23fF
C230 a_1740_73.n11 VNB 0.09fF
C231 a_1740_73.n12 VNB 0.00fF
C232 a_599_943.n0 VNB 0.04fF
C233 a_599_943.n1 VNB 0.58fF
C234 a_599_943.n2 VNB 0.69fF
C235 a_599_943.n3 VNB 0.35fF
C236 a_599_943.n4 VNB 0.42fF
C237 a_599_943.n5 VNB 0.42fF
C238 a_599_943.n6 VNB 0.42fF
C239 a_599_943.t9 VNB 0.56fF
C240 a_599_943.n7 VNB 0.41fF
C241 a_599_943.n8 VNB 1.11fF
C242 a_599_943.n9 VNB 0.46fF
C243 a_599_943.n10 VNB 0.04fF
C244 a_599_943.n11 VNB 0.31fF
C245 a_599_943.n12 VNB 0.06fF
C246 a_5366_73.n0 VNB 0.02fF
C247 a_5366_73.n1 VNB 0.10fF
C248 a_5366_73.n2 VNB 0.06fF
C249 a_5366_73.n3 VNB 0.06fF
C250 a_5366_73.n4 VNB 0.00fF
C251 a_5366_73.n5 VNB 0.04fF
C252 a_5366_73.n6 VNB 0.05fF
C253 a_5366_73.n7 VNB 0.02fF
C254 a_5366_73.n8 VNB 0.05fF
C255 a_5366_73.n9 VNB 0.08fF
C256 a_5366_73.n10 VNB 0.17fF
C257 a_5366_73.t1 VNB 0.23fF
C258 a_5366_73.n11 VNB 0.09fF
C259 a_5366_73.n12 VNB 0.00fF
C260 a_8861_1004.n0 VNB 0.80fF
C261 a_8861_1004.n1 VNB 0.80fF
C262 a_8861_1004.n2 VNB 0.94fF
C263 a_8861_1004.n3 VNB 0.30fF
C264 a_8861_1004.n4 VNB 0.43fF
C265 a_8861_1004.n5 VNB 0.53fF
C266 a_8861_1004.n6 VNB 0.69fF
C267 a_8861_1004.n7 VNB 0.53fF
C268 a_8861_1004.n8 VNB 0.58fF
C269 a_8861_1004.n9 VNB 2.86fF
C270 a_8861_1004.n10 VNB 0.68fF
C271 a_8861_1004.n11 VNB 0.12fF
C272 a_8861_1004.n12 VNB 0.45fF
C273 a_8861_1004.n13 VNB 0.07fF
C274 a_8731_159.n0 VNB 0.85fF
C275 a_8731_159.n1 VNB 1.01fF
C276 a_8731_159.n2 VNB 0.41fF
C277 a_8731_159.n3 VNB 0.46fF
C278 a_8731_159.t11 VNB 0.92fF
C279 a_8731_159.n4 VNB 0.65fF
C280 a_8731_159.n5 VNB 0.46fF
C281 a_8731_159.t8 VNB 0.92fF
C282 a_8731_159.n6 VNB 0.60fF
C283 a_8731_159.n7 VNB 0.46fF
C284 a_8731_159.n8 VNB 0.86fF
C285 a_8731_159.n9 VNB 2.83fF
C286 a_8731_159.n10 VNB 2.11fF
C287 a_8731_159.n11 VNB 0.68fF
C288 a_8731_159.n12 VNB 0.13fF
C289 a_8731_159.n13 VNB 0.54fF
C290 a_8731_159.n14 VNB 0.07fF
C291 a_8030_73.n0 VNB 0.02fF
C292 a_8030_73.n1 VNB 0.10fF
C293 a_8030_73.n2 VNB 0.06fF
C294 a_8030_73.n3 VNB 0.06fF
C295 a_8030_73.n4 VNB 0.00fF
C296 a_8030_73.n5 VNB 0.04fF
C297 a_8030_73.n6 VNB 0.05fF
C298 a_8030_73.n7 VNB 0.02fF
C299 a_8030_73.n8 VNB 0.05fF
C300 a_8030_73.n9 VNB 0.08fF
C301 a_8030_73.n10 VNB 0.17fF
C302 a_8030_73.t1 VNB 0.23fF
C303 a_8030_73.n11 VNB 0.09fF
C304 a_8030_73.n12 VNB 0.00fF
C305 a_277_1004.n0 VNB 0.74fF
C306 a_277_1004.n1 VNB 0.74fF
C307 a_277_1004.n2 VNB 0.86fF
C308 a_277_1004.n3 VNB 0.27fF
C309 a_277_1004.n4 VNB 0.39fF
C310 a_277_1004.n5 VNB 0.49fF
C311 a_277_1004.n6 VNB 0.63fF
C312 a_277_1004.n7 VNB 0.49fF
C313 a_277_1004.n8 VNB 0.53fF
C314 a_277_1004.n9 VNB 2.63fF
C315 a_277_1004.n10 VNB 0.62fF
C316 a_277_1004.n11 VNB 0.11fF
C317 a_277_1004.n12 VNB 0.42fF
C318 a_277_1004.n13 VNB 0.06fF
C319 a_7595_383.n0 VNB 0.05fF
C320 a_7595_383.n1 VNB 0.72fF
C321 a_7595_383.n2 VNB 0.85fF
C322 a_7595_383.n3 VNB 0.55fF
C323 a_7595_383.n4 VNB 0.39fF
C324 a_7595_383.n5 VNB 0.44fF
C325 a_7595_383.t13 VNB 0.77fF
C326 a_7595_383.n6 VNB 1.30fF
C327 a_7595_383.n7 VNB 1.08fF
C328 a_7595_383.t8 VNB 0.59fF
C329 a_7595_383.n8 VNB 1.09fF
C330 a_7595_383.n9 VNB 0.60fF
C331 a_7595_383.t9 VNB 0.59fF
C332 a_7595_383.n10 VNB 0.51fF
C333 a_7595_383.n11 VNB 5.56fF
C334 a_7595_383.n12 VNB 0.57fF
C335 a_7595_383.n13 VNB 0.05fF
C336 a_7595_383.n14 VNB 0.25fF
C337 a_7595_383.n15 VNB 0.07fF
C338 a_13757_1005.n0 VNB 0.28fF
C339 a_13757_1005.n1 VNB 0.29fF
C340 a_13757_1005.n2 VNB 0.20fF
C341 a_13757_1005.n3 VNB 0.56fF
C342 a_13757_1005.n4 VNB 0.25fF
C343 a_13757_1005.n5 VNB 0.35fF
C344 a_4569_1004.n0 VNB 0.06fF
C345 a_4569_1004.n1 VNB 0.81fF
C346 a_4569_1004.n2 VNB 0.81fF
C347 a_4569_1004.n3 VNB 0.95fF
C348 a_4569_1004.n4 VNB 0.30fF
C349 a_4569_1004.n5 VNB 0.43fF
C350 a_4569_1004.n6 VNB 0.54fF
C351 a_4569_1004.n7 VNB 0.69fF
C352 a_4569_1004.n8 VNB 0.54fF
C353 a_4569_1004.n9 VNB 0.58fF
C354 a_4569_1004.n10 VNB 2.89fF
C355 a_4569_1004.n11 VNB 0.67fF
C356 a_4569_1004.n12 VNB 0.05fF
C357 a_4569_1004.n13 VNB 0.47fF
C358 a_4569_1004.n14 VNB 0.08fF
C359 a_6137_1004.n0 VNB 0.05fF
C360 a_6137_1004.n1 VNB 0.61fF
C361 a_6137_1004.n2 VNB 0.73fF
C362 a_6137_1004.n3 VNB 0.37fF
C363 a_6137_1004.n4 VNB 0.45fF
C364 a_6137_1004.n5 VNB 0.65fF
C365 a_6137_1004.n6 VNB 0.69fF
C366 a_6137_1004.n7 VNB 0.04fF
C367 a_6137_1004.n8 VNB 0.32fF
C368 a_6137_1004.n9 VNB 0.06fF
C369 a_4891_943.n0 VNB 0.05fF
C370 a_4891_943.n1 VNB 0.71fF
C371 a_4891_943.n2 VNB 0.84fF
C372 a_4891_943.n3 VNB 0.43fF
C373 a_4891_943.n4 VNB 0.52fF
C374 a_4891_943.n5 VNB 0.52fF
C375 a_4891_943.n6 VNB 0.52fF
C376 a_4891_943.t10 VNB 0.69fF
C377 a_4891_943.n7 VNB 0.50fF
C378 a_4891_943.n8 VNB 1.37fF
C379 a_4891_943.n9 VNB 0.56fF
C380 a_4891_943.n10 VNB 0.05fF
C381 a_4891_943.n11 VNB 0.37fF
C382 a_4891_943.n12 VNB 0.07fF
C383 a_1845_1004.n0 VNB 0.04fF
C384 a_1845_1004.n1 VNB 0.55fF
C385 a_1845_1004.n2 VNB 0.65fF
C386 a_1845_1004.n3 VNB 0.33fF
C387 a_1845_1004.n4 VNB 0.40fF
C388 a_1845_1004.n5 VNB 0.58fF
C389 a_1845_1004.n6 VNB 0.62fF
C390 a_1845_1004.n7 VNB 0.04fF
C391 a_1845_1004.n8 VNB 0.29fF
C392 a_1845_1004.n9 VNB 0.06fF
C393 a_147_159.n0 VNB 0.06fF
C394 a_147_159.n1 VNB 0.81fF
C395 a_147_159.n2 VNB 0.96fF
C396 a_147_159.n3 VNB 0.39fF
C397 a_147_159.n4 VNB 0.44fF
C398 a_147_159.t12 VNB 0.88fF
C399 a_147_159.n5 VNB 0.61fF
C400 a_147_159.n6 VNB 0.44fF
C401 a_147_159.t9 VNB 0.88fF
C402 a_147_159.n7 VNB 0.57fF
C403 a_147_159.n8 VNB 0.44fF
C404 a_147_159.n9 VNB 0.82fF
C405 a_147_159.n10 VNB 2.69fF
C406 a_147_159.n11 VNB 2.00fF
C407 a_147_159.n12 VNB 0.64fF
C408 a_147_159.n13 VNB 0.05fF
C409 a_147_159.n14 VNB 0.52fF
C410 a_147_159.n15 VNB 0.08fF
C411 a_13093_1005.n0 VNB 0.36fF
C412 a_13093_1005.n1 VNB 0.32fF
C413 a_13093_1005.n2 VNB 0.23fF
C414 a_13093_1005.n3 VNB 0.62fF
C415 a_13093_1005.n4 VNB 0.28fF
C416 a_13093_1005.n5 VNB 0.40fF
C417 VPB.n0 VNB 0.03fF
C418 VPB.n1 VNB 0.04fF
C419 VPB.n2 VNB 0.02fF
C420 VPB.n3 VNB 0.19fF
C421 VPB.n5 VNB 0.02fF
C422 VPB.n6 VNB 0.02fF
C423 VPB.n7 VNB 0.02fF
C424 VPB.n8 VNB 0.02fF
C425 VPB.n10 VNB 0.02fF
C426 VPB.n11 VNB 0.02fF
C427 VPB.n12 VNB 0.02fF
C428 VPB.n14 VNB 0.10fF
C429 VPB.n15 VNB 0.10fF
C430 VPB.n16 VNB 0.02fF
C431 VPB.n17 VNB 0.02fF
C432 VPB.n18 VNB 0.02fF
C433 VPB.n19 VNB 0.04fF
C434 VPB.n20 VNB 0.02fF
C435 VPB.n21 VNB 0.25fF
C436 VPB.n22 VNB 0.04fF
C437 VPB.n24 VNB 0.02fF
C438 VPB.n25 VNB 0.02fF
C439 VPB.n26 VNB 0.02fF
C440 VPB.n27 VNB 0.02fF
C441 VPB.n29 VNB 0.02fF
C442 VPB.n30 VNB 0.02fF
C443 VPB.n31 VNB 0.02fF
C444 VPB.n33 VNB 0.28fF
C445 VPB.n35 VNB 0.03fF
C446 VPB.n36 VNB 0.02fF
C447 VPB.n37 VNB 0.03fF
C448 VPB.n38 VNB 0.03fF
C449 VPB.n39 VNB 0.28fF
C450 VPB.n40 VNB 0.01fF
C451 VPB.n41 VNB 0.02fF
C452 VPB.n42 VNB 0.28fF
C453 VPB.n43 VNB 0.02fF
C454 VPB.n44 VNB 0.02fF
C455 VPB.n45 VNB 0.06fF
C456 VPB.n46 VNB 0.21fF
C457 VPB.n47 VNB 0.02fF
C458 VPB.n48 VNB 0.01fF
C459 VPB.n49 VNB 0.14fF
C460 VPB.n50 VNB 0.17fF
C461 VPB.n51 VNB 0.02fF
C462 VPB.n52 VNB 0.02fF
C463 VPB.n53 VNB 0.14fF
C464 VPB.n54 VNB 0.17fF
C465 VPB.n55 VNB 0.02fF
C466 VPB.n56 VNB 0.02fF
C467 VPB.n57 VNB 0.02fF
C468 VPB.n58 VNB 0.14fF
C469 VPB.n59 VNB 0.16fF
C470 VPB.n60 VNB 0.02fF
C471 VPB.n61 VNB 0.02fF
C472 VPB.n62 VNB 0.14fF
C473 VPB.n63 VNB 0.15fF
C474 VPB.n64 VNB 0.02fF
C475 VPB.n65 VNB 0.02fF
C476 VPB.n66 VNB 0.02fF
C477 VPB.n67 VNB 0.14fF
C478 VPB.n68 VNB 0.17fF
C479 VPB.n69 VNB 0.02fF
C480 VPB.n70 VNB 0.02fF
C481 VPB.n71 VNB 0.14fF
C482 VPB.n72 VNB 0.17fF
C483 VPB.n73 VNB 0.02fF
C484 VPB.n74 VNB 0.02fF
C485 VPB.n75 VNB 0.22fF
C486 VPB.n76 VNB 0.02fF
C487 VPB.n77 VNB 0.01fF
C488 VPB.n78 VNB 0.06fF
C489 VPB.n79 VNB 0.28fF
C490 VPB.n80 VNB 0.02fF
C491 VPB.n81 VNB 0.02fF
C492 VPB.n82 VNB 0.10fF
C493 VPB.n83 VNB 0.02fF
C494 VPB.n84 VNB 0.02fF
C495 VPB.n85 VNB 0.02fF
C496 VPB.n86 VNB 0.04fF
C497 VPB.n87 VNB 0.02fF
C498 VPB.n88 VNB 0.20fF
C499 VPB.n89 VNB 0.04fF
C500 VPB.n91 VNB 0.02fF
C501 VPB.n92 VNB 0.02fF
C502 VPB.n93 VNB 0.02fF
C503 VPB.n94 VNB 0.02fF
C504 VPB.n96 VNB 0.02fF
C505 VPB.n97 VNB 0.02fF
C506 VPB.n98 VNB 0.02fF
C507 VPB.n100 VNB 0.28fF
C508 VPB.n102 VNB 0.03fF
C509 VPB.n103 VNB 0.02fF
C510 VPB.n104 VNB 0.10fF
C511 VPB.n105 VNB 0.14fF
C512 VPB.n106 VNB 0.16fF
C513 VPB.n107 VNB 0.02fF
C514 VPB.n108 VNB 0.02fF
C515 VPB.n109 VNB 0.02fF
C516 VPB.n110 VNB 0.14fF
C517 VPB.n111 VNB 0.15fF
C518 VPB.n112 VNB 0.02fF
C519 VPB.n113 VNB 0.02fF
C520 VPB.n114 VNB 0.14fF
C521 VPB.n115 VNB 0.17fF
C522 VPB.n116 VNB 0.02fF
C523 VPB.n117 VNB 0.02fF
C524 VPB.n118 VNB 0.06fF
C525 VPB.n119 VNB 0.24fF
C526 VPB.n120 VNB 0.02fF
C527 VPB.n121 VNB 0.01fF
C528 VPB.n122 VNB 0.28fF
C529 VPB.n123 VNB 0.01fF
C530 VPB.n124 VNB 0.02fF
C531 VPB.n125 VNB 0.03fF
C532 VPB.n126 VNB 0.03fF
C533 VPB.n127 VNB 0.28fF
C534 VPB.n128 VNB 0.01fF
C535 VPB.n129 VNB 0.02fF
C536 VPB.n130 VNB 0.24fF
C537 VPB.n131 VNB 0.02fF
C538 VPB.n132 VNB 0.01fF
C539 VPB.n133 VNB 0.06fF
C540 VPB.n134 VNB 0.14fF
C541 VPB.n135 VNB 0.17fF
C542 VPB.n136 VNB 0.02fF
C543 VPB.n137 VNB 0.02fF
C544 VPB.n138 VNB 0.14fF
C545 VPB.n139 VNB 0.16fF
C546 VPB.n140 VNB 0.02fF
C547 VPB.n141 VNB 0.02fF
C548 VPB.n142 VNB 0.02fF
C549 VPB.n143 VNB 0.14fF
C550 VPB.n144 VNB 0.15fF
C551 VPB.n145 VNB 0.02fF
C552 VPB.n146 VNB 0.02fF
C553 VPB.n147 VNB 0.02fF
C554 VPB.n148 VNB 0.02fF
C555 VPB.n149 VNB 0.02fF
C556 VPB.n150 VNB 0.14fF
C557 VPB.n151 VNB 0.03fF
C558 VPB.n152 VNB 0.02fF
C559 VPB.n153 VNB 0.05fF
C560 VPB.n154 VNB 0.01fF
C561 VPB.n156 VNB 0.02fF
C562 VPB.n157 VNB 0.02fF
C563 VPB.n159 VNB 0.02fF
C564 VPB.n160 VNB 0.02fF
C565 VPB.n161 VNB 0.02fF
C566 VPB.n164 VNB 0.47fF
C567 VPB.n166 VNB 0.04fF
C568 VPB.n167 VNB 0.04fF
C569 VPB.n168 VNB 0.28fF
C570 VPB.n169 VNB 0.03fF
C571 VPB.n170 VNB 0.04fF
C572 VPB.n171 VNB 0.28fF
C573 VPB.n172 VNB 0.02fF
C574 VPB.n173 VNB 0.02fF
C575 VPB.n174 VNB 0.28fF
C576 VPB.n175 VNB 0.02fF
C577 VPB.n176 VNB 0.02fF
C578 VPB.n177 VNB 0.28fF
C579 VPB.n178 VNB 0.02fF
C580 VPB.n179 VNB 0.02fF
C581 VPB.n180 VNB 0.00fF
C582 VPB.n181 VNB 0.10fF
C583 VPB.n182 VNB 0.02fF
C584 VPB.n183 VNB 0.28fF
C585 VPB.n184 VNB 0.02fF
C586 VPB.n185 VNB 0.02fF
C587 VPB.n186 VNB 0.02fF
C588 VPB.n187 VNB 0.28fF
C589 VPB.n188 VNB 0.02fF
C590 VPB.n189 VNB 0.02fF
C591 VPB.n190 VNB 0.02fF
C592 VPB.n191 VNB 0.28fF
C593 VPB.n192 VNB 0.02fF
C594 VPB.n193 VNB 0.02fF
C595 VPB.n194 VNB 0.02fF
C596 VPB.n195 VNB 0.28fF
C597 VPB.n196 VNB 0.01fF
C598 VPB.n197 VNB 0.02fF
C599 VPB.n198 VNB 0.04fF
C600 VPB.n199 VNB 0.02fF
C601 VPB.n200 VNB 0.02fF
C602 VPB.n201 VNB 0.02fF
C603 VPB.n202 VNB 0.04fF
C604 VPB.n203 VNB 0.02fF
C605 VPB.n204 VNB 0.21fF
C606 VPB.n205 VNB 0.04fF
C607 VPB.n207 VNB 0.02fF
C608 VPB.n208 VNB 0.02fF
C609 VPB.n209 VNB 0.02fF
C610 VPB.n210 VNB 0.02fF
C611 VPB.n212 VNB 0.02fF
C612 VPB.n213 VNB 0.02fF
C613 VPB.n214 VNB 0.02fF
C614 VPB.n216 VNB 0.28fF
C615 VPB.n218 VNB 0.03fF
C616 VPB.n219 VNB 0.02fF
C617 VPB.n220 VNB 0.03fF
C618 VPB.n221 VNB 0.03fF
C619 VPB.n222 VNB 0.28fF
C620 VPB.n223 VNB 0.01fF
C621 VPB.n224 VNB 0.02fF
C622 VPB.n225 VNB 0.04fF
C623 VPB.n226 VNB 0.28fF
C624 VPB.n227 VNB 0.02fF
C625 VPB.n228 VNB 0.02fF
C626 VPB.n229 VNB 0.02fF
C627 VPB.n230 VNB 0.28fF
C628 VPB.n231 VNB 0.02fF
C629 VPB.n232 VNB 0.02fF
C630 VPB.n233 VNB 0.02fF
C631 VPB.n234 VNB 0.28fF
C632 VPB.n235 VNB 0.02fF
C633 VPB.n236 VNB 0.02fF
C634 VPB.n237 VNB 0.02fF
C635 VPB.n238 VNB 0.28fF
C636 VPB.n239 VNB 0.02fF
C637 VPB.n240 VNB 0.02fF
C638 VPB.n241 VNB 0.02fF
C639 VPB.n242 VNB 0.28fF
C640 VPB.n243 VNB 0.02fF
C641 VPB.n244 VNB 0.02fF
C642 VPB.n245 VNB 0.02fF
C643 VPB.n246 VNB 0.28fF
C644 VPB.n247 VNB 0.02fF
C645 VPB.n248 VNB 0.02fF
C646 VPB.n249 VNB 0.02fF
C647 VPB.n250 VNB 0.28fF
C648 VPB.n251 VNB 0.01fF
C649 VPB.n252 VNB 0.02fF
C650 VPB.n253 VNB 0.04fF
C651 VPB.n254 VNB 0.02fF
C652 VPB.n255 VNB 0.02fF
C653 VPB.n256 VNB 0.02fF
C654 VPB.n257 VNB 0.04fF
C655 VPB.n258 VNB 0.02fF
C656 VPB.n259 VNB 0.20fF
C657 VPB.n260 VNB 0.04fF
C658 VPB.n262 VNB 0.02fF
C659 VPB.n263 VNB 0.02fF
C660 VPB.n264 VNB 0.02fF
C661 VPB.n265 VNB 0.02fF
C662 VPB.n267 VNB 0.02fF
C663 VPB.n268 VNB 0.02fF
C664 VPB.n269 VNB 0.02fF
C665 VPB.n271 VNB 0.28fF
C666 VPB.n273 VNB 0.03fF
C667 VPB.n274 VNB 0.02fF
C668 VPB.n275 VNB 0.03fF
C669 VPB.n276 VNB 0.03fF
C670 VPB.n277 VNB 0.28fF
C671 VPB.n278 VNB 0.01fF
C672 VPB.n279 VNB 0.02fF
C673 VPB.n280 VNB 0.04fF
C674 VPB.n281 VNB 0.06fF
C675 VPB.n282 VNB 0.24fF
C676 VPB.n283 VNB 0.02fF
C677 VPB.n284 VNB 0.01fF
C678 VPB.n285 VNB 0.02fF
C679 VPB.n286 VNB 0.14fF
C680 VPB.n287 VNB 0.17fF
C681 VPB.n288 VNB 0.02fF
C682 VPB.n289 VNB 0.02fF
C683 VPB.n290 VNB 0.02fF
C684 VPB.n291 VNB 0.10fF
C685 VPB.n292 VNB 0.02fF
C686 VPB.n293 VNB 0.14fF
C687 VPB.n294 VNB 0.16fF
C688 VPB.n295 VNB 0.02fF
C689 VPB.n296 VNB 0.02fF
C690 VPB.n297 VNB 0.02fF
C691 VPB.n298 VNB 0.14fF
C692 VPB.n299 VNB 0.15fF
C693 VPB.n300 VNB 0.02fF
C694 VPB.n301 VNB 0.02fF
C695 VPB.n302 VNB 0.02fF
C696 VPB.n303 VNB 0.14fF
C697 VPB.n304 VNB 0.17fF
C698 VPB.n305 VNB 0.02fF
C699 VPB.n306 VNB 0.02fF
C700 VPB.n307 VNB 0.02fF
C701 VPB.n308 VNB 0.06fF
C702 VPB.n309 VNB 0.24fF
C703 VPB.n310 VNB 0.02fF
C704 VPB.n311 VNB 0.01fF
C705 VPB.n312 VNB 0.02fF
C706 VPB.n313 VNB 0.28fF
C707 VPB.n314 VNB 0.01fF
C708 VPB.n315 VNB 0.02fF
C709 VPB.n316 VNB 0.04fF
C710 VPB.n317 VNB 0.02fF
C711 VPB.n318 VNB 0.02fF
C712 VPB.n319 VNB 0.02fF
C713 VPB.n320 VNB 0.04fF
C714 VPB.n321 VNB 0.02fF
C715 VPB.n322 VNB 0.20fF
C716 VPB.n323 VNB 0.04fF
C717 VPB.n325 VNB 0.02fF
C718 VPB.n326 VNB 0.02fF
C719 VPB.n327 VNB 0.02fF
C720 VPB.n328 VNB 0.02fF
C721 VPB.n330 VNB 0.02fF
C722 VPB.n331 VNB 0.02fF
C723 VPB.n332 VNB 0.02fF
C724 VPB.n334 VNB 0.28fF
C725 VPB.n336 VNB 0.03fF
C726 VPB.n337 VNB 0.02fF
C727 VPB.n338 VNB 0.03fF
C728 VPB.n339 VNB 0.03fF
C729 VPB.n340 VNB 0.28fF
C730 VPB.n341 VNB 0.01fF
C731 VPB.n342 VNB 0.02fF
C732 VPB.n343 VNB 0.04fF
C733 VPB.n344 VNB 0.06fF
C734 VPB.n345 VNB 0.24fF
C735 VPB.n346 VNB 0.02fF
C736 VPB.n347 VNB 0.01fF
C737 VPB.n348 VNB 0.02fF
C738 VPB.n349 VNB 0.14fF
C739 VPB.n350 VNB 0.17fF
C740 VPB.n351 VNB 0.02fF
C741 VPB.n352 VNB 0.02fF
C742 VPB.n353 VNB 0.02fF
C743 VPB.n354 VNB 0.10fF
C744 VPB.n355 VNB 0.02fF
C745 VPB.n356 VNB 0.14fF
C746 VPB.n357 VNB 0.16fF
C747 VPB.n358 VNB 0.02fF
C748 VPB.n359 VNB 0.02fF
C749 VPB.n360 VNB 0.02fF
C750 VPB.n361 VNB 0.14fF
C751 VPB.n362 VNB 0.15fF
C752 VPB.n363 VNB 0.02fF
C753 VPB.n364 VNB 0.02fF
C754 VPB.n365 VNB 0.02fF
C755 VPB.n366 VNB 0.14fF
C756 VPB.n367 VNB 0.17fF
C757 VPB.n368 VNB 0.02fF
C758 VPB.n369 VNB 0.02fF
C759 VPB.n370 VNB 0.02fF
C760 VPB.n371 VNB 0.06fF
C761 VPB.n372 VNB 0.24fF
C762 VPB.n373 VNB 0.02fF
C763 VPB.n374 VNB 0.01fF
C764 VPB.n375 VNB 0.02fF
C765 VPB.n376 VNB 0.28fF
C766 VPB.n377 VNB 0.01fF
C767 VPB.n378 VNB 0.02fF
C768 VPB.n379 VNB 0.04fF
C769 VPB.n380 VNB 0.02fF
C770 VPB.n381 VNB 0.02fF
C771 VPB.n382 VNB 0.02fF
C772 VPB.n383 VNB 0.04fF
C773 VPB.n384 VNB 0.02fF
C774 VPB.n385 VNB 0.20fF
C775 VPB.n386 VNB 0.04fF
C776 VPB.n388 VNB 0.02fF
C777 VPB.n389 VNB 0.02fF
C778 VPB.n390 VNB 0.02fF
C779 VPB.n391 VNB 0.02fF
C780 VPB.n393 VNB 0.02fF
C781 VPB.n394 VNB 0.02fF
C782 VPB.n395 VNB 0.02fF
C783 VPB.n397 VNB 0.28fF
C784 VPB.n399 VNB 0.03fF
C785 VPB.n400 VNB 0.02fF
C786 VPB.n401 VNB 0.03fF
C787 VPB.n402 VNB 0.03fF
C788 VPB.n403 VNB 0.28fF
C789 VPB.n404 VNB 0.01fF
C790 VPB.n405 VNB 0.02fF
C791 VPB.n406 VNB 0.04fF
C792 VPB.n407 VNB 0.06fF
C793 VPB.n408 VNB 0.24fF
C794 VPB.n409 VNB 0.02fF
C795 VPB.n410 VNB 0.01fF
C796 VPB.n411 VNB 0.02fF
C797 VPB.n412 VNB 0.14fF
C798 VPB.n413 VNB 0.17fF
C799 VPB.n414 VNB 0.02fF
C800 VPB.n415 VNB 0.02fF
C801 VPB.n416 VNB 0.02fF
C802 VPB.n417 VNB 0.10fF
C803 VPB.n418 VNB 0.02fF
C804 VPB.n419 VNB 0.14fF
C805 VPB.n420 VNB 0.16fF
C806 VPB.n421 VNB 0.02fF
C807 VPB.n422 VNB 0.02fF
C808 VPB.n423 VNB 0.02fF
C809 VPB.n424 VNB 0.14fF
C810 VPB.n425 VNB 0.15fF
C811 VPB.n426 VNB 0.02fF
C812 VPB.n427 VNB 0.02fF
C813 VPB.n428 VNB 0.02fF
C814 VPB.n429 VNB 0.14fF
C815 VPB.n430 VNB 0.17fF
C816 VPB.n431 VNB 0.02fF
C817 VPB.n432 VNB 0.02fF
C818 VPB.n433 VNB 0.02fF
C819 VPB.n434 VNB 0.06fF
C820 VPB.n435 VNB 0.24fF
C821 VPB.n436 VNB 0.02fF
C822 VPB.n437 VNB 0.01fF
C823 VPB.n438 VNB 0.02fF
C824 VPB.n439 VNB 0.28fF
C825 VPB.n440 VNB 0.01fF
C826 VPB.n441 VNB 0.02fF
C827 VPB.n442 VNB 0.04fF
C828 VPB.n443 VNB 0.02fF
C829 VPB.n444 VNB 0.02fF
C830 VPB.n445 VNB 0.02fF
C831 VPB.n446 VNB 0.04fF
C832 VPB.n447 VNB 0.02fF
C833 VPB.n448 VNB 0.20fF
C834 VPB.n449 VNB 0.04fF
C835 VPB.n451 VNB 0.02fF
C836 VPB.n452 VNB 0.02fF
C837 VPB.n453 VNB 0.02fF
C838 VPB.n454 VNB 0.02fF
C839 VPB.n456 VNB 0.02fF
C840 VPB.n457 VNB 0.02fF
C841 VPB.n458 VNB 0.02fF
C842 VPB.n460 VNB 0.28fF
C843 VPB.n462 VNB 0.03fF
C844 VPB.n463 VNB 0.02fF
C845 VPB.n464 VNB 0.03fF
C846 VPB.n465 VNB 0.03fF
C847 VPB.n466 VNB 0.28fF
C848 VPB.n467 VNB 0.01fF
C849 VPB.n468 VNB 0.02fF
C850 VPB.n469 VNB 0.04fF
C851 VPB.n470 VNB 0.06fF
C852 VPB.n471 VNB 0.24fF
C853 VPB.n472 VNB 0.02fF
C854 VPB.n473 VNB 0.01fF
C855 VPB.n474 VNB 0.02fF
C856 VPB.n475 VNB 0.14fF
C857 VPB.n476 VNB 0.17fF
C858 VPB.n477 VNB 0.02fF
C859 VPB.n478 VNB 0.02fF
C860 VPB.n479 VNB 0.02fF
C861 VPB.n480 VNB 0.10fF
C862 VPB.n481 VNB 0.02fF
C863 VPB.n482 VNB 0.14fF
C864 VPB.n483 VNB 0.16fF
C865 VPB.n484 VNB 0.02fF
C866 VPB.n485 VNB 0.02fF
C867 VPB.n486 VNB 0.02fF
C868 VPB.n487 VNB 0.14fF
C869 VPB.n488 VNB 0.15fF
C870 VPB.n489 VNB 0.02fF
C871 VPB.n490 VNB 0.02fF
C872 VPB.n491 VNB 0.02fF
C873 VPB.n492 VNB 0.14fF
C874 VPB.n493 VNB 0.17fF
C875 VPB.n494 VNB 0.02fF
C876 VPB.n495 VNB 0.02fF
C877 VPB.n496 VNB 0.02fF
C878 VPB.n497 VNB 0.06fF
C879 VPB.n498 VNB 0.24fF
C880 VPB.n499 VNB 0.02fF
C881 VPB.n500 VNB 0.01fF
C882 VPB.n501 VNB 0.02fF
C883 VPB.n502 VNB 0.28fF
C884 VPB.n503 VNB 0.01fF
C885 VPB.n504 VNB 0.02fF
C886 VPB.n505 VNB 0.04fF
C887 VPB.n506 VNB 0.02fF
C888 VPB.n507 VNB 0.02fF
C889 VPB.n508 VNB 0.02fF
C890 VPB.n509 VNB 0.04fF
C891 VPB.n510 VNB 0.02fF
C892 VPB.n511 VNB 0.20fF
C893 VPB.n512 VNB 0.04fF
C894 VPB.n514 VNB 0.02fF
C895 VPB.n515 VNB 0.02fF
C896 VPB.n516 VNB 0.02fF
C897 VPB.n517 VNB 0.02fF
C898 VPB.n519 VNB 0.02fF
C899 VPB.n520 VNB 0.02fF
C900 VPB.n521 VNB 0.02fF
C901 VPB.n523 VNB 0.28fF
C902 VPB.n525 VNB 0.03fF
C903 VPB.n526 VNB 0.02fF
C904 VPB.n527 VNB 0.03fF
C905 VPB.n528 VNB 0.03fF
C906 VPB.n529 VNB 0.28fF
C907 VPB.n530 VNB 0.01fF
C908 VPB.n531 VNB 0.02fF
C909 VPB.n532 VNB 0.04fF
C910 VPB.n533 VNB 0.06fF
C911 VPB.n534 VNB 0.24fF
C912 VPB.n535 VNB 0.02fF
C913 VPB.n536 VNB 0.01fF
C914 VPB.n537 VNB 0.02fF
C915 VPB.n538 VNB 0.14fF
C916 VPB.n539 VNB 0.17fF
C917 VPB.n540 VNB 0.02fF
C918 VPB.n541 VNB 0.02fF
C919 VPB.n542 VNB 0.02fF
C920 VPB.n543 VNB 0.10fF
C921 VPB.n544 VNB 0.02fF
C922 VPB.n545 VNB 0.14fF
C923 VPB.n546 VNB 0.16fF
C924 VPB.n547 VNB 0.02fF
C925 VPB.n548 VNB 0.02fF
C926 VPB.n549 VNB 0.02fF
C927 VPB.n550 VNB 0.14fF
C928 VPB.n551 VNB 0.15fF
C929 VPB.n552 VNB 0.02fF
C930 VPB.n553 VNB 0.02fF
C931 VPB.n554 VNB 0.02fF
C932 VPB.n555 VNB 0.14fF
C933 VPB.n556 VNB 0.17fF
C934 VPB.n557 VNB 0.02fF
C935 VPB.n558 VNB 0.02fF
C936 VPB.n559 VNB 0.02fF
C937 VPB.n560 VNB 0.06fF
C938 VPB.n561 VNB 0.24fF
C939 VPB.n562 VNB 0.02fF
C940 VPB.n563 VNB 0.01fF
C941 VPB.n564 VNB 0.02fF
C942 VPB.n565 VNB 0.28fF
C943 VPB.n566 VNB 0.01fF
C944 VPB.n567 VNB 0.02fF
C945 VPB.n568 VNB 0.04fF
C946 VPB.n569 VNB 0.02fF
C947 VPB.n570 VNB 0.02fF
C948 VPB.n571 VNB 0.02fF
C949 VPB.n572 VNB 0.04fF
C950 VPB.n573 VNB 0.02fF
C951 VPB.n574 VNB 0.20fF
C952 VPB.n575 VNB 0.04fF
C953 VPB.n577 VNB 0.02fF
C954 VPB.n578 VNB 0.02fF
C955 VPB.n579 VNB 0.02fF
C956 VPB.n580 VNB 0.02fF
C957 VPB.n582 VNB 0.02fF
C958 VPB.n583 VNB 0.02fF
C959 VPB.n584 VNB 0.02fF
C960 VPB.n586 VNB 0.28fF
C961 VPB.n588 VNB 0.03fF
C962 VPB.n589 VNB 0.02fF
C963 VPB.n590 VNB 0.03fF
C964 VPB.n591 VNB 0.03fF
C965 VPB.n592 VNB 0.28fF
C966 VPB.n593 VNB 0.01fF
C967 VPB.n594 VNB 0.02fF
C968 VPB.n595 VNB 0.04fF
C969 VPB.n596 VNB 0.06fF
C970 VPB.n597 VNB 0.24fF
C971 VPB.n598 VNB 0.02fF
C972 VPB.n599 VNB 0.01fF
C973 VPB.n600 VNB 0.02fF
C974 VPB.n601 VNB 0.14fF
C975 VPB.n602 VNB 0.17fF
C976 VPB.n603 VNB 0.02fF
C977 VPB.n604 VNB 0.02fF
C978 VPB.n605 VNB 0.02fF
C979 VPB.n606 VNB 0.10fF
C980 VPB.n607 VNB 0.02fF
C981 VPB.n608 VNB 0.14fF
C982 VPB.n609 VNB 0.16fF
C983 VPB.n610 VNB 0.02fF
C984 VPB.n611 VNB 0.02fF
C985 VPB.n612 VNB 0.02fF
C986 VPB.n613 VNB 0.14fF
C987 VPB.n614 VNB 0.15fF
C988 VPB.n615 VNB 0.02fF
C989 VPB.n616 VNB 0.02fF
C990 VPB.n617 VNB 0.02fF
C991 VPB.n618 VNB 0.14fF
C992 VPB.n619 VNB 0.17fF
C993 VPB.n620 VNB 0.02fF
C994 VPB.n621 VNB 0.02fF
C995 VPB.n622 VNB 0.02fF
C996 VPB.n623 VNB 0.06fF
C997 VPB.n624 VNB 0.24fF
C998 VPB.n625 VNB 0.02fF
C999 VPB.n626 VNB 0.01fF
C1000 VPB.n627 VNB 0.02fF
C1001 VPB.n628 VNB 0.28fF
C1002 VPB.n629 VNB 0.01fF
C1003 VPB.n630 VNB 0.02fF
C1004 VPB.n631 VNB 0.04fF
C1005 VPB.n632 VNB 0.02fF
C1006 VPB.n633 VNB 0.02fF
C1007 VPB.n634 VNB 0.02fF
C1008 VPB.n635 VNB 0.04fF
C1009 VPB.n636 VNB 0.02fF
C1010 VPB.n637 VNB 0.25fF
C1011 VPB.n638 VNB 0.04fF
C1012 VPB.n640 VNB 0.02fF
C1013 VPB.n641 VNB 0.02fF
C1014 VPB.n642 VNB 0.02fF
C1015 VPB.n643 VNB 0.02fF
C1016 VPB.n645 VNB 0.02fF
C1017 VPB.n646 VNB 0.02fF
C1018 VPB.n647 VNB 0.02fF
C1019 VPB.n649 VNB 0.28fF
C1020 VPB.n651 VNB 0.03fF
C1021 VPB.n652 VNB 0.02fF
C1022 VPB.n653 VNB 0.03fF
C1023 VPB.n654 VNB 0.03fF
C1024 VPB.n655 VNB 0.28fF
C1025 VPB.n656 VNB 0.01fF
C1026 VPB.n657 VNB 0.02fF
C1027 VPB.n658 VNB 0.04fF
C1028 VPB.n659 VNB 0.28fF
C1029 VPB.n660 VNB 0.02fF
C1030 VPB.n661 VNB 0.02fF
C1031 VPB.n662 VNB 0.02fF
C1032 VPB.n663 VNB 0.06fF
C1033 VPB.n664 VNB 0.21fF
C1034 VPB.n665 VNB 0.02fF
C1035 VPB.n666 VNB 0.01fF
C1036 VPB.n667 VNB 0.02fF
C1037 VPB.n668 VNB 0.14fF
C1038 VPB.n669 VNB 0.17fF
C1039 VPB.n670 VNB 0.02fF
C1040 VPB.n671 VNB 0.02fF
C1041 VPB.n672 VNB 0.02fF
C1042 VPB.n673 VNB 0.10fF
C1043 VPB.n674 VNB 0.02fF
C1044 VPB.n675 VNB 0.14fF
C1045 VPB.n676 VNB 0.17fF
C1046 VPB.n677 VNB 0.02fF
C1047 VPB.n678 VNB 0.02fF
C1048 VPB.n679 VNB 0.02fF
C1049 VPB.n680 VNB 0.14fF
C1050 VPB.n681 VNB 0.16fF
C1051 VPB.n682 VNB 0.02fF
C1052 VPB.n683 VNB 0.02fF
C1053 VPB.n684 VNB 0.02fF
C1054 VPB.n685 VNB 0.14fF
C1055 VPB.n686 VNB 0.15fF
C1056 VPB.n687 VNB 0.02fF
C1057 VPB.n688 VNB 0.02fF
C1058 VPB.n689 VNB 0.02fF
C1059 VPB.n690 VNB 0.10fF
C1060 VPB.n691 VNB 0.02fF
C1061 VPB.n692 VNB 0.14fF
C1062 VPB.n693 VNB 0.17fF
C1063 VPB.n694 VNB 0.02fF
C1064 VPB.n695 VNB 0.02fF
C1065 VPB.n696 VNB 0.02fF
C1066 VPB.n697 VNB 0.14fF
C1067 VPB.n698 VNB 0.17fF
C1068 VPB.n699 VNB 0.02fF
C1069 VPB.n700 VNB 0.02fF
C1070 VPB.n701 VNB 0.02fF
C1071 VPB.n702 VNB 0.06fF
C1072 VPB.n703 VNB 0.22fF
C1073 VPB.n704 VNB 0.02fF
C1074 VPB.n705 VNB 0.01fF
C1075 VPB.n706 VNB 0.02fF
C1076 VPB.n707 VNB 0.28fF
C1077 VPB.n708 VNB 0.02fF
C1078 VPB.n709 VNB 0.02fF
C1079 VPB.n710 VNB 0.02fF
C1080 VPB.n711 VNB 0.28fF
C1081 VPB.n712 VNB 0.01fF
C1082 VPB.n713 VNB 0.02fF
C1083 VPB.n714 VNB 0.04fF
C1084 VPB.n715 VNB 0.02fF
C1085 VPB.n716 VNB 0.02fF
C1086 VPB.n717 VNB 0.02fF
C1087 VPB.n718 VNB 0.04fF
C1088 VPB.n719 VNB 0.02fF
C1089 VPB.n720 VNB 0.25fF
C1090 VPB.n721 VNB 0.04fF
C1091 VPB.n723 VNB 0.02fF
C1092 VPB.n724 VNB 0.02fF
C1093 VPB.n725 VNB 0.02fF
C1094 VPB.n726 VNB 0.02fF
C1095 VPB.n728 VNB 0.02fF
C1096 VPB.n729 VNB 0.02fF
C1097 VPB.n730 VNB 0.02fF
C1098 VPB.n732 VNB 0.28fF
C1099 VPB.n734 VNB 0.03fF
C1100 VPB.n735 VNB 0.02fF
C1101 VPB.n736 VNB 0.03fF
C1102 VPB.n737 VNB 0.03fF
C1103 VPB.n738 VNB 0.28fF
C1104 VPB.n739 VNB 0.01fF
C1105 VPB.n740 VNB 0.02fF
C1106 VPB.n741 VNB 0.04fF
C1107 VPB.n742 VNB 0.06fF
C1108 VPB.n743 VNB 0.24fF
C1109 VPB.n744 VNB 0.02fF
C1110 VPB.n745 VNB 0.01fF
C1111 VPB.n746 VNB 0.02fF
C1112 VPB.n747 VNB 0.14fF
C1113 VPB.n748 VNB 0.17fF
C1114 VPB.n749 VNB 0.02fF
C1115 VPB.n750 VNB 0.02fF
C1116 VPB.n751 VNB 0.02fF
C1117 VPB.n752 VNB 0.02fF
C1118 VPB.n753 VNB 0.02fF
C1119 VPB.n754 VNB 0.02fF
C1120 VPB.n755 VNB 0.02fF
C1121 VPB.n756 VNB 0.04fF
C1122 VPB.n757 VNB 0.04fF
C1123 VPB.n758 VNB 0.02fF
C1124 VPB.n759 VNB 0.02fF
C1125 VPB.n760 VNB 0.02fF
C1126 VPB.n761 VNB 0.02fF
C1127 VPB.n762 VNB 0.02fF
C1128 VPB.n763 VNB 0.14fF
C1129 VPB.n764 VNB 0.17fF
C1130 VPB.n765 VNB 0.02fF
C1131 VPB.n766 VNB 0.02fF
C1132 VPB.n767 VNB 0.06fF
C1133 VPB.n768 VNB 0.24fF
C1134 VPB.n769 VNB 0.02fF
C1135 VPB.n770 VNB 0.01fF
C1136 VPB.n771 VNB 0.02fF
C1137 VPB.n772 VNB 0.28fF
C1138 VPB.n773 VNB 0.01fF
C1139 VPB.n774 VNB 0.02fF
C1140 VPB.n775 VNB 0.04fF
C1141 VPB.n776 VNB 0.02fF
C1142 VPB.n777 VNB 0.02fF
C1143 VPB.n778 VNB 0.02fF
C1144 VPB.n779 VNB 0.04fF
C1145 VPB.n780 VNB 0.02fF
C1146 VPB.n781 VNB 0.20fF
C1147 VPB.n782 VNB 0.04fF
C1148 VPB.n784 VNB 0.02fF
C1149 VPB.n785 VNB 0.02fF
C1150 VPB.n786 VNB 0.02fF
C1151 VPB.n787 VNB 0.02fF
C1152 VPB.n789 VNB 0.02fF
C1153 VPB.n790 VNB 0.02fF
C1154 VPB.n791 VNB 0.02fF
C1155 VPB.n793 VNB 0.28fF
C1156 VPB.n795 VNB 0.03fF
C1157 VPB.n796 VNB 0.02fF
C1158 VPB.n797 VNB 0.03fF
C1159 VPB.n798 VNB 0.03fF
C1160 VPB.n799 VNB 0.28fF
C1161 VPB.n800 VNB 0.01fF
C1162 VPB.n801 VNB 0.02fF
C1163 VPB.n802 VNB 0.04fF
C1164 VPB.n803 VNB 0.06fF
C1165 VPB.n804 VNB 0.24fF
C1166 VPB.n805 VNB 0.02fF
C1167 VPB.n806 VNB 0.01fF
C1168 VPB.n807 VNB 0.02fF
C1169 VPB.n808 VNB 0.14fF
C1170 VPB.n809 VNB 0.17fF
C1171 VPB.n810 VNB 0.02fF
C1172 VPB.n811 VNB 0.02fF
C1173 VPB.n812 VNB 0.02fF
C1174 VPB.n813 VNB 0.10fF
C1175 VPB.n814 VNB 0.02fF
C1176 VPB.n815 VNB 0.14fF
C1177 VPB.n816 VNB 0.16fF
C1178 VPB.n817 VNB 0.02fF
C1179 VPB.n818 VNB 0.02fF
C1180 VPB.n819 VNB 0.02fF
C1181 VPB.n820 VNB 0.14fF
C1182 VPB.n821 VNB 0.15fF
C1183 VPB.n822 VNB 0.02fF
C1184 VPB.n823 VNB 0.02fF
C1185 VPB.n824 VNB 0.02fF
C1186 VPB.n825 VNB 0.14fF
C1187 VPB.n826 VNB 0.17fF
C1188 VPB.n827 VNB 0.02fF
C1189 VPB.n828 VNB 0.02fF
C1190 VPB.n829 VNB 0.02fF
C1191 VPB.n830 VNB 0.06fF
C1192 VPB.n831 VNB 0.24fF
C1193 VPB.n832 VNB 0.02fF
C1194 VPB.n833 VNB 0.01fF
C1195 VPB.n834 VNB 0.02fF
C1196 VPB.n835 VNB 0.28fF
C1197 VPB.n836 VNB 0.01fF
C1198 VPB.n837 VNB 0.02fF
C1199 VPB.n838 VNB 0.04fF
C1200 VPB.n839 VNB 0.02fF
C1201 VPB.n840 VNB 0.02fF
C1202 VPB.n841 VNB 0.02fF
C1203 VPB.n842 VNB 0.04fF
C1204 VPB.n843 VNB 0.02fF
C1205 VPB.n844 VNB 0.20fF
C1206 VPB.n845 VNB 0.04fF
C1207 VPB.n847 VNB 0.02fF
C1208 VPB.n848 VNB 0.02fF
C1209 VPB.n849 VNB 0.02fF
C1210 VPB.n850 VNB 0.02fF
C1211 VPB.n852 VNB 0.02fF
C1212 VPB.n853 VNB 0.02fF
C1213 VPB.n854 VNB 0.02fF
C1214 VPB.n856 VNB 0.28fF
C1215 VPB.n858 VNB 0.03fF
C1216 VPB.n859 VNB 0.02fF
C1217 VPB.n860 VNB 0.03fF
C1218 VPB.n861 VNB 0.03fF
C1219 VPB.n862 VNB 0.28fF
C1220 VPB.n863 VNB 0.01fF
C1221 VPB.n864 VNB 0.02fF
C1222 VPB.n865 VNB 0.04fF
C1223 VPB.n866 VNB 0.06fF
C1224 VPB.n867 VNB 0.24fF
C1225 VPB.n868 VNB 0.02fF
C1226 VPB.n869 VNB 0.01fF
C1227 VPB.n870 VNB 0.02fF
C1228 VPB.n871 VNB 0.14fF
C1229 VPB.n872 VNB 0.17fF
C1230 VPB.n873 VNB 0.02fF
C1231 VPB.n874 VNB 0.02fF
C1232 VPB.n875 VNB 0.02fF
C1233 VPB.n876 VNB 0.10fF
C1234 VPB.n877 VNB 0.02fF
C1235 VPB.n878 VNB 0.14fF
C1236 VPB.n879 VNB 0.16fF
C1237 VPB.n880 VNB 0.02fF
C1238 VPB.n881 VNB 0.02fF
C1239 VPB.n882 VNB 0.02fF
C1240 VPB.n883 VNB 0.14fF
C1241 VPB.n884 VNB 0.15fF
C1242 VPB.n885 VNB 0.02fF
C1243 VPB.n886 VNB 0.02fF
C1244 VPB.n887 VNB 0.02fF
C1245 VPB.n888 VNB 0.14fF
C1246 VPB.n889 VNB 0.17fF
C1247 VPB.n890 VNB 0.02fF
C1248 VPB.n891 VNB 0.02fF
C1249 VPB.n892 VNB 0.02fF
C1250 VPB.n893 VNB 0.06fF
C1251 VPB.n894 VNB 0.24fF
C1252 VPB.n895 VNB 0.02fF
C1253 VPB.n896 VNB 0.01fF
C1254 VPB.n897 VNB 0.02fF
C1255 VPB.n898 VNB 0.28fF
C1256 VPB.n899 VNB 0.01fF
C1257 VPB.n900 VNB 0.02fF
C1258 VPB.n901 VNB 0.04fF
C1259 VPB.n902 VNB 0.02fF
C1260 VPB.n903 VNB 0.02fF
C1261 VPB.n904 VNB 0.02fF
C1262 VPB.n905 VNB 0.04fF
C1263 VPB.n906 VNB 0.02fF
C1264 VPB.n907 VNB 0.20fF
C1265 VPB.n908 VNB 0.04fF
C1266 VPB.n910 VNB 0.02fF
C1267 VPB.n911 VNB 0.02fF
C1268 VPB.n912 VNB 0.02fF
C1269 VPB.n913 VNB 0.02fF
C1270 VPB.n915 VNB 0.02fF
C1271 VPB.n916 VNB 0.02fF
C1272 VPB.n917 VNB 0.02fF
C1273 VPB.n919 VNB 0.28fF
C1274 VPB.n921 VNB 0.03fF
C1275 VPB.n922 VNB 0.02fF
C1276 VPB.n923 VNB 0.03fF
C1277 VPB.n924 VNB 0.03fF
C1278 VPB.n925 VNB 0.28fF
C1279 VPB.n926 VNB 0.01fF
C1280 VPB.n927 VNB 0.02fF
C1281 VPB.n928 VNB 0.04fF
C1282 VPB.n929 VNB 0.06fF
C1283 VPB.n930 VNB 0.24fF
C1284 VPB.n931 VNB 0.02fF
C1285 VPB.n932 VNB 0.01fF
C1286 VPB.n933 VNB 0.02fF
C1287 VPB.n934 VNB 0.14fF
C1288 VPB.n935 VNB 0.17fF
C1289 VPB.n936 VNB 0.02fF
C1290 VPB.n937 VNB 0.02fF
C1291 VPB.n938 VNB 0.02fF
C1292 VPB.n939 VNB 0.10fF
C1293 VPB.n940 VNB 0.02fF
C1294 VPB.n941 VNB 0.14fF
C1295 VPB.n942 VNB 0.16fF
C1296 VPB.n943 VNB 0.02fF
C1297 VPB.n944 VNB 0.02fF
C1298 VPB.n945 VNB 0.02fF
C1299 VPB.n946 VNB 0.14fF
C1300 VPB.n947 VNB 0.15fF
C1301 VPB.n948 VNB 0.02fF
C1302 VPB.n949 VNB 0.02fF
C1303 VPB.n950 VNB 0.02fF
C1304 VPB.n951 VNB 0.14fF
C1305 VPB.n952 VNB 0.17fF
C1306 VPB.n953 VNB 0.02fF
C1307 VPB.n954 VNB 0.02fF
C1308 VPB.n955 VNB 0.02fF
C1309 VPB.n956 VNB 0.06fF
C1310 VPB.n957 VNB 0.24fF
C1311 VPB.n958 VNB 0.02fF
C1312 VPB.n959 VNB 0.01fF
C1313 VPB.n960 VNB 0.02fF
C1314 VPB.n961 VNB 0.28fF
C1315 VPB.n962 VNB 0.01fF
C1316 VPB.n963 VNB 0.02fF
C1317 VPB.n964 VNB 0.04fF
C1318 VPB.n965 VNB 0.02fF
C1319 VPB.n966 VNB 0.02fF
C1320 VPB.n967 VNB 0.02fF
C1321 VPB.n968 VNB 0.04fF
C1322 VPB.n969 VNB 0.02fF
C1323 VPB.n970 VNB 0.25fF
C1324 VPB.n971 VNB 0.04fF
C1325 VPB.n973 VNB 0.02fF
C1326 VPB.n974 VNB 0.02fF
C1327 VPB.n975 VNB 0.02fF
C1328 VPB.n976 VNB 0.02fF
C1329 VPB.n978 VNB 0.02fF
C1330 VPB.n979 VNB 0.02fF
C1331 VPB.n980 VNB 0.02fF
C1332 VPB.n982 VNB 0.28fF
C1333 VPB.n984 VNB 0.03fF
C1334 VPB.n985 VNB 0.02fF
C1335 VPB.n986 VNB 0.03fF
C1336 VPB.n987 VNB 0.03fF
C1337 VPB.n988 VNB 0.28fF
C1338 VPB.n989 VNB 0.01fF
C1339 VPB.n990 VNB 0.02fF
C1340 VPB.n991 VNB 0.04fF
C1341 VPB.n992 VNB 0.28fF
C1342 VPB.n993 VNB 0.02fF
C1343 VPB.n994 VNB 0.02fF
C1344 VPB.n995 VNB 0.02fF
C1345 VPB.n996 VNB 0.06fF
C1346 VPB.n997 VNB 0.21fF
C1347 VPB.n998 VNB 0.02fF
C1348 VPB.n999 VNB 0.01fF
C1349 VPB.n1000 VNB 0.02fF
C1350 VPB.n1001 VNB 0.14fF
C1351 VPB.n1002 VNB 0.17fF
C1352 VPB.n1003 VNB 0.02fF
C1353 VPB.n1004 VNB 0.02fF
C1354 VPB.n1005 VNB 0.02fF
C1355 VPB.n1006 VNB 0.10fF
C1356 VPB.n1007 VNB 0.02fF
C1357 VPB.n1008 VNB 0.14fF
C1358 VPB.n1009 VNB 0.17fF
C1359 VPB.n1010 VNB 0.02fF
C1360 VPB.n1011 VNB 0.02fF
C1361 VPB.n1012 VNB 0.02fF
C1362 VPB.n1013 VNB 0.14fF
C1363 VPB.n1014 VNB 0.16fF
C1364 VPB.n1015 VNB 0.02fF
C1365 VPB.n1016 VNB 0.02fF
C1366 VPB.n1017 VNB 0.02fF
C1367 VPB.n1018 VNB 0.14fF
C1368 VPB.n1019 VNB 0.15fF
C1369 VPB.n1020 VNB 0.02fF
C1370 VPB.n1021 VNB 0.02fF
C1371 VPB.n1022 VNB 0.02fF
C1372 VPB.n1023 VNB 0.10fF
C1373 VPB.n1024 VNB 0.02fF
C1374 VPB.n1025 VNB 0.14fF
C1375 VPB.n1026 VNB 0.17fF
C1376 VPB.n1027 VNB 0.02fF
C1377 VPB.n1028 VNB 0.02fF
C1378 VPB.n1029 VNB 0.02fF
C1379 VPB.n1030 VNB 0.14fF
C1380 VPB.n1031 VNB 0.17fF
C1381 VPB.n1032 VNB 0.02fF
C1382 VPB.n1033 VNB 0.02fF
C1383 VPB.n1034 VNB 0.02fF
C1384 VPB.n1035 VNB 0.06fF
C1385 VPB.n1036 VNB 0.22fF
C1386 VPB.n1037 VNB 0.02fF
C1387 VPB.n1038 VNB 0.01fF
C1388 VPB.n1039 VNB 0.02fF
C1389 VPB.n1040 VNB 0.28fF
C1390 VPB.n1041 VNB 0.02fF
C1391 VPB.n1042 VNB 0.02fF
C1392 VPB.n1043 VNB 0.02fF
C1393 VPB.n1044 VNB 0.28fF
C1394 VPB.n1045 VNB 0.01fF
C1395 VPB.n1046 VNB 0.02fF
C1396 VPB.n1047 VNB 0.04fF
C1397 VPB.n1048 VNB 0.02fF
C1398 VPB.n1049 VNB 0.02fF
C1399 VPB.n1050 VNB 0.02fF
C1400 VPB.n1051 VNB 0.04fF
C1401 VPB.n1052 VNB 0.02fF
C1402 VPB.n1053 VNB 0.25fF
C1403 VPB.n1054 VNB 0.04fF
C1404 VPB.n1056 VNB 0.02fF
C1405 VPB.n1057 VNB 0.02fF
C1406 VPB.n1058 VNB 0.02fF
C1407 VPB.n1059 VNB 0.02fF
C1408 VPB.n1061 VNB 0.02fF
C1409 VPB.n1062 VNB 0.02fF
C1410 VPB.n1063 VNB 0.02fF
C1411 VPB.n1065 VNB 0.28fF
C1412 VPB.n1067 VNB 0.03fF
C1413 VPB.n1068 VNB 0.02fF
C1414 VPB.n1069 VNB 0.03fF
C1415 VPB.n1070 VNB 0.03fF
C1416 VPB.n1071 VNB 0.28fF
C1417 VPB.n1072 VNB 0.01fF
C1418 VPB.n1073 VNB 0.02fF
C1419 VPB.n1074 VNB 0.04fF
C1420 VPB.n1075 VNB 0.06fF
C1421 VPB.n1076 VNB 0.24fF
C1422 VPB.n1077 VNB 0.02fF
C1423 VPB.n1078 VNB 0.01fF
C1424 VPB.n1079 VNB 0.02fF
C1425 VPB.n1080 VNB 0.14fF
C1426 VPB.n1081 VNB 0.17fF
C1427 VPB.n1082 VNB 0.02fF
C1428 VPB.n1083 VNB 0.02fF
C1429 VPB.n1084 VNB 0.02fF
C1430 VPB.n1085 VNB 0.10fF
C1431 VPB.n1086 VNB 0.02fF
C1432 VPB.n1087 VNB 0.14fF
C1433 VPB.n1088 VNB 0.16fF
C1434 VPB.n1089 VNB 0.02fF
C1435 VPB.n1090 VNB 0.02fF
C1436 VPB.n1091 VNB 0.02fF
C1437 VPB.n1092 VNB 0.14fF
C1438 VPB.n1093 VNB 0.15fF
C1439 VPB.n1094 VNB 0.02fF
C1440 VPB.n1095 VNB 0.02fF
C1441 VPB.n1096 VNB 0.02fF
C1442 VPB.n1097 VNB 0.14fF
C1443 VPB.n1098 VNB 0.17fF
C1444 VPB.n1099 VNB 0.02fF
C1445 VPB.n1100 VNB 0.02fF
C1446 VPB.n1101 VNB 0.02fF
C1447 VPB.n1102 VNB 0.06fF
C1448 VPB.n1103 VNB 0.24fF
C1449 VPB.n1104 VNB 0.02fF
C1450 VPB.n1105 VNB 0.01fF
C1451 VPB.n1106 VNB 0.02fF
C1452 VPB.n1107 VNB 0.28fF
C1453 VPB.n1108 VNB 0.01fF
C1454 VPB.n1109 VNB 0.02fF
C1455 VPB.n1110 VNB 0.04fF
C1456 VPB.n1111 VNB 0.02fF
C1457 VPB.n1112 VNB 0.02fF
C1458 VPB.n1113 VNB 0.02fF
C1459 VPB.n1114 VNB 0.04fF
C1460 VPB.n1115 VNB 0.02fF
C1461 VPB.n1116 VNB 0.20fF
C1462 VPB.n1117 VNB 0.04fF
C1463 VPB.n1119 VNB 0.02fF
C1464 VPB.n1120 VNB 0.02fF
C1465 VPB.n1121 VNB 0.02fF
C1466 VPB.n1122 VNB 0.02fF
C1467 VPB.n1124 VNB 0.02fF
C1468 VPB.n1125 VNB 0.02fF
C1469 VPB.n1126 VNB 0.02fF
C1470 VPB.n1128 VNB 0.28fF
C1471 VPB.n1130 VNB 0.03fF
C1472 VPB.n1131 VNB 0.02fF
C1473 VPB.n1132 VNB 0.03fF
C1474 VPB.n1133 VNB 0.03fF
C1475 VPB.n1134 VNB 0.28fF
C1476 VPB.n1135 VNB 0.01fF
C1477 VPB.n1136 VNB 0.02fF
C1478 VPB.n1137 VNB 0.04fF
C1479 VPB.n1138 VNB 0.06fF
C1480 VPB.n1139 VNB 0.24fF
C1481 VPB.n1140 VNB 0.02fF
C1482 VPB.n1141 VNB 0.01fF
C1483 VPB.n1142 VNB 0.02fF
C1484 VPB.n1143 VNB 0.14fF
C1485 VPB.n1144 VNB 0.17fF
C1486 VPB.n1145 VNB 0.02fF
C1487 VPB.n1146 VNB 0.02fF
C1488 VPB.n1147 VNB 0.02fF
C1489 VPB.n1148 VNB 0.10fF
C1490 VPB.n1149 VNB 0.02fF
C1491 VPB.n1150 VNB 0.14fF
C1492 VPB.n1151 VNB 0.16fF
C1493 VPB.n1152 VNB 0.02fF
C1494 VPB.n1153 VNB 0.02fF
C1495 VPB.n1154 VNB 0.02fF
C1496 VPB.n1155 VNB 0.14fF
C1497 VPB.n1156 VNB 0.15fF
C1498 VPB.n1157 VNB 0.02fF
C1499 VPB.n1158 VNB 0.02fF
C1500 VPB.n1159 VNB 0.02fF
C1501 VPB.n1160 VNB 0.14fF
C1502 VPB.n1161 VNB 0.17fF
C1503 VPB.n1162 VNB 0.02fF
C1504 VPB.n1163 VNB 0.02fF
C1505 VPB.n1164 VNB 0.02fF
C1506 VPB.n1165 VNB 0.06fF
C1507 VPB.n1166 VNB 0.24fF
C1508 VPB.n1167 VNB 0.02fF
C1509 VPB.n1168 VNB 0.01fF
C1510 VPB.n1169 VNB 0.02fF
C1511 VPB.n1170 VNB 0.28fF
C1512 VPB.n1171 VNB 0.01fF
C1513 VPB.n1172 VNB 0.02fF
C1514 VPB.n1173 VNB 0.04fF
C1515 VPB.n1174 VNB 0.02fF
C1516 VPB.n1175 VNB 0.02fF
C1517 VPB.n1176 VNB 0.02fF
C1518 VPB.n1177 VNB 0.04fF
C1519 VPB.n1178 VNB 0.02fF
C1520 VPB.n1179 VNB 0.20fF
C1521 VPB.n1180 VNB 0.04fF
C1522 VPB.n1182 VNB 0.02fF
C1523 VPB.n1183 VNB 0.02fF
C1524 VPB.n1184 VNB 0.02fF
C1525 VPB.n1185 VNB 0.02fF
C1526 VPB.n1187 VNB 0.02fF
C1527 VPB.n1188 VNB 0.02fF
C1528 VPB.n1189 VNB 0.02fF
C1529 VPB.n1191 VNB 0.28fF
C1530 VPB.n1193 VNB 0.03fF
C1531 VPB.n1194 VNB 0.02fF
C1532 VPB.n1195 VNB 0.03fF
C1533 VPB.n1196 VNB 0.03fF
C1534 VPB.n1197 VNB 0.28fF
C1535 VPB.n1198 VNB 0.01fF
C1536 VPB.n1199 VNB 0.02fF
C1537 VPB.n1200 VNB 0.04fF
C1538 VPB.n1201 VNB 0.06fF
C1539 VPB.n1202 VNB 0.24fF
C1540 VPB.n1203 VNB 0.02fF
C1541 VPB.n1204 VNB 0.01fF
C1542 VPB.n1205 VNB 0.02fF
C1543 VPB.n1206 VNB 0.14fF
C1544 VPB.n1207 VNB 0.17fF
C1545 VPB.n1208 VNB 0.02fF
C1546 VPB.n1209 VNB 0.02fF
C1547 VPB.n1210 VNB 0.02fF
C1548 VPB.n1211 VNB 0.10fF
C1549 VPB.n1212 VNB 0.02fF
C1550 VPB.n1213 VNB 0.14fF
C1551 VPB.n1214 VNB 0.16fF
C1552 VPB.n1215 VNB 0.02fF
C1553 VPB.n1216 VNB 0.02fF
C1554 VPB.n1217 VNB 0.02fF
C1555 VPB.n1218 VNB 0.14fF
C1556 VPB.n1219 VNB 0.15fF
C1557 VPB.n1220 VNB 0.02fF
C1558 VPB.n1221 VNB 0.02fF
C1559 VPB.n1222 VNB 0.02fF
C1560 VPB.n1223 VNB 0.14fF
C1561 VPB.n1224 VNB 0.17fF
C1562 VPB.n1225 VNB 0.02fF
C1563 VPB.n1226 VNB 0.02fF
C1564 VPB.n1227 VNB 0.02fF
C1565 VPB.n1228 VNB 0.06fF
C1566 VPB.n1229 VNB 0.24fF
C1567 VPB.n1230 VNB 0.02fF
C1568 VPB.n1231 VNB 0.01fF
C1569 VPB.n1232 VNB 0.02fF
C1570 VPB.n1233 VNB 0.28fF
C1571 VPB.n1234 VNB 0.01fF
C1572 VPB.n1235 VNB 0.02fF
C1573 VPB.n1236 VNB 0.04fF
C1574 VPB.n1237 VNB 0.02fF
C1575 VPB.n1238 VNB 0.02fF
C1576 VPB.n1239 VNB 0.02fF
C1577 VPB.n1240 VNB 0.04fF
C1578 VPB.n1241 VNB 0.02fF
C1579 VPB.n1242 VNB 0.20fF
C1580 VPB.n1243 VNB 0.04fF
C1581 VPB.n1245 VNB 0.02fF
C1582 VPB.n1246 VNB 0.02fF
C1583 VPB.n1247 VNB 0.02fF
C1584 VPB.n1248 VNB 0.02fF
C1585 VPB.n1250 VNB 0.02fF
C1586 VPB.n1251 VNB 0.02fF
C1587 VPB.n1252 VNB 0.02fF
C1588 VPB.n1254 VNB 0.28fF
C1589 VPB.n1256 VNB 0.03fF
C1590 VPB.n1257 VNB 0.02fF
C1591 VPB.n1258 VNB 0.03fF
C1592 VPB.n1259 VNB 0.03fF
C1593 VPB.n1260 VNB 0.28fF
C1594 VPB.n1261 VNB 0.01fF
C1595 VPB.n1262 VNB 0.02fF
C1596 VPB.n1263 VNB 0.04fF
C1597 VPB.n1264 VNB 0.06fF
C1598 VPB.n1265 VNB 0.24fF
C1599 VPB.n1266 VNB 0.02fF
C1600 VPB.n1267 VNB 0.01fF
C1601 VPB.n1268 VNB 0.02fF
C1602 VPB.n1269 VNB 0.14fF
C1603 VPB.n1270 VNB 0.17fF
C1604 VPB.n1271 VNB 0.02fF
C1605 VPB.n1272 VNB 0.02fF
C1606 VPB.n1273 VNB 0.02fF
C1607 VPB.n1274 VNB 0.10fF
C1608 VPB.n1275 VNB 0.02fF
C1609 VPB.n1276 VNB 0.14fF
C1610 VPB.n1277 VNB 0.16fF
C1611 VPB.n1278 VNB 0.02fF
C1612 VPB.n1279 VNB 0.02fF
C1613 VPB.n1280 VNB 0.02fF
C1614 VPB.n1281 VNB 0.14fF
C1615 VPB.n1282 VNB 0.15fF
C1616 VPB.n1283 VNB 0.02fF
C1617 VPB.n1284 VNB 0.02fF
C1618 VPB.n1285 VNB 0.02fF
C1619 VPB.n1286 VNB 0.14fF
C1620 VPB.n1287 VNB 0.17fF
C1621 VPB.n1288 VNB 0.02fF
C1622 VPB.n1289 VNB 0.02fF
C1623 VPB.n1290 VNB 0.02fF
C1624 VPB.n1291 VNB 0.06fF
C1625 VPB.n1292 VNB 0.24fF
C1626 VPB.n1293 VNB 0.02fF
C1627 VPB.n1294 VNB 0.01fF
C1628 VPB.n1295 VNB 0.02fF
C1629 VPB.n1296 VNB 0.28fF
C1630 VPB.n1297 VNB 0.01fF
C1631 VPB.n1298 VNB 0.02fF
C1632 VPB.n1299 VNB 0.04fF
C1633 VPB.n1300 VNB 0.02fF
C1634 VPB.n1301 VNB 0.02fF
C1635 VPB.n1302 VNB 0.02fF
C1636 VPB.n1303 VNB 0.04fF
C1637 VPB.n1304 VNB 0.02fF
C1638 VPB.n1305 VNB 0.20fF
C1639 VPB.n1306 VNB 0.04fF
C1640 VPB.n1308 VNB 0.02fF
C1641 VPB.n1309 VNB 0.02fF
C1642 VPB.n1310 VNB 0.02fF
C1643 VPB.n1311 VNB 0.02fF
C1644 VPB.n1313 VNB 0.02fF
C1645 VPB.n1314 VNB 0.02fF
C1646 VPB.n1315 VNB 0.02fF
C1647 VPB.n1317 VNB 0.28fF
C1648 VPB.n1319 VNB 0.03fF
C1649 VPB.n1320 VNB 0.02fF
C1650 VPB.n1321 VNB 0.03fF
C1651 VPB.n1322 VNB 0.03fF
C1652 VPB.n1323 VNB 0.28fF
C1653 VPB.n1324 VNB 0.01fF
C1654 VPB.n1325 VNB 0.02fF
C1655 VPB.n1326 VNB 0.04fF
C1656 VPB.n1327 VNB 0.06fF
C1657 VPB.n1328 VNB 0.24fF
C1658 VPB.n1329 VNB 0.02fF
C1659 VPB.n1330 VNB 0.01fF
C1660 VPB.n1331 VNB 0.02fF
C1661 VPB.n1332 VNB 0.14fF
C1662 VPB.n1333 VNB 0.17fF
C1663 VPB.n1334 VNB 0.02fF
C1664 VPB.n1335 VNB 0.02fF
C1665 VPB.n1336 VNB 0.02fF
C1666 VPB.n1337 VNB 0.10fF
C1667 VPB.n1338 VNB 0.02fF
C1668 VPB.n1339 VNB 0.14fF
C1669 VPB.n1340 VNB 0.16fF
C1670 VPB.n1341 VNB 0.02fF
C1671 VPB.n1342 VNB 0.02fF
C1672 VPB.n1343 VNB 0.02fF
C1673 VPB.n1344 VNB 0.14fF
C1674 VPB.n1345 VNB 0.15fF
C1675 VPB.n1346 VNB 0.02fF
C1676 VPB.n1347 VNB 0.02fF
C1677 VPB.n1348 VNB 0.02fF
C1678 VPB.n1349 VNB 0.14fF
C1679 VPB.n1350 VNB 0.17fF
C1680 VPB.n1351 VNB 0.02fF
C1681 VPB.n1352 VNB 0.02fF
C1682 VPB.n1353 VNB 0.02fF
C1683 VPB.n1354 VNB 0.06fF
C1684 VPB.n1355 VNB 0.24fF
C1685 VPB.n1356 VNB 0.02fF
C1686 VPB.n1357 VNB 0.01fF
C1687 VPB.n1358 VNB 0.02fF
C1688 VPB.n1359 VNB 0.28fF
C1689 VPB.n1360 VNB 0.01fF
C1690 VPB.n1361 VNB 0.02fF
C1691 VPB.n1362 VNB 0.04fF
C1692 VPB.n1363 VNB 0.04fF
C1693 VPB.n1364 VNB 0.02fF
C1694 VPB.n1365 VNB 0.02fF
C1695 VPB.n1366 VNB 0.02fF
C1696 VPB.n1367 VNB 0.02fF
C1697 VPB.n1368 VNB 0.02fF
C1698 VPB.n1369 VNB 0.02fF
C1699 VPB.n1370 VNB 0.02fF
C1700 VPB.n1371 VNB 0.02fF
C1701 VPB.n1372 VNB 0.02fF
C1702 VPB.n1373 VNB 0.02fF
C1703 VPB.n1374 VNB 0.03fF
C1704 VPB.n1375 VNB 0.04fF
C1705 VPB.n1376 VNB 0.02fF
C1706 VPB.n1377 VNB 0.02fF
C1707 VPB.n1378 VNB 0.02fF
C1708 VPB.n1379 VNB 0.04fF
C1709 VPB.n1380 VNB 0.04fF
C1710 VPB.n1382 VNB 0.44fF
C1711 a_11887_383.n0 VNB 0.54fF
C1712 a_11887_383.n1 VNB 0.64fF
C1713 a_11887_383.n2 VNB 0.29fF
C1714 a_11887_383.n3 VNB 0.26fF
C1715 a_11887_383.n4 VNB 0.29fF
C1716 a_11887_383.n5 VNB 0.74fF
C1717 a_11887_383.n6 VNB 0.52fF
C1718 a_11887_383.n7 VNB 0.36fF
C1719 a_11887_383.n8 VNB 0.32fF
C1720 a_11887_383.t10 VNB 0.55fF
C1721 a_11887_383.n9 VNB 0.39fF
C1722 a_11887_383.n10 VNB 0.97fF
C1723 a_11887_383.n11 VNB 0.43fF
C1724 a_11887_383.n12 VNB 0.08fF
C1725 a_11887_383.n13 VNB 0.31fF
C1726 a_11887_383.n14 VNB 0.05fF
C1727 a_4383_75.n0 VNB 0.20fF
C1728 a_4383_75.n1 VNB 0.04fF
C1729 a_4383_75.n2 VNB 0.01fF
C1730 a_4383_75.n3 VNB 0.08fF
C1731 a_4383_75.n4 VNB 0.06fF
C1732 a_4383_75.n5 VNB 0.07fF
C1733 a_4439_159.n0 VNB 0.07fF
C1734 a_4439_159.n1 VNB 0.89fF
C1735 a_4439_159.n2 VNB 1.05fF
C1736 a_4439_159.n3 VNB 0.43fF
C1737 a_4439_159.n4 VNB 0.48fF
C1738 a_4439_159.t7 VNB 0.96fF
C1739 a_4439_159.n5 VNB 0.67fF
C1740 a_4439_159.n6 VNB 0.48fF
C1741 a_4439_159.t12 VNB 0.96fF
C1742 a_4439_159.n7 VNB 0.63fF
C1743 a_4439_159.n8 VNB 0.48fF
C1744 a_4439_159.n9 VNB 0.90fF
C1745 a_4439_159.n10 VNB 2.95fF
C1746 a_4439_159.n11 VNB 2.19fF
C1747 a_4439_159.n12 VNB 0.70fF
C1748 a_4439_159.n13 VNB 0.06fF
C1749 a_4439_159.n14 VNB 0.57fF
C1750 a_4439_159.n15 VNB 0.09fF
C1751 a_10990_73.n0 VNB 0.08fF
C1752 a_10990_73.n1 VNB 0.02fF
C1753 a_10990_73.n2 VNB 0.01fF
C1754 a_10990_73.n3 VNB 0.10fF
C1755 a_10990_73.n4 VNB 0.07fF
C1756 a_10990_73.n5 VNB 0.05fF
C1757 a_10990_73.n6 VNB 0.02fF
C1758 a_10990_73.n7 VNB 0.05fF
C1759 a_10429_1004.n0 VNB 0.61fF
C1760 a_10429_1004.n1 VNB 0.72fF
C1761 a_10429_1004.n2 VNB 0.36fF
C1762 a_10429_1004.n3 VNB 0.44fF
C1763 a_10429_1004.n4 VNB 0.64fF
C1764 a_10429_1004.n5 VNB 0.69fF
C1765 a_10429_1004.n6 VNB 0.09fF
C1766 a_10429_1004.n7 VNB 0.31fF
C1767 a_10429_1004.n8 VNB 0.05fF
.ends
