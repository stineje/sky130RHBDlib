* SPICE3 file created from AND2X1.ext - technology: sky130A

.subckt AND2X1 Y A B VDD GND
M1000 GND A.t1 a_112_101.t0 nshort w=-1.605u l=1.765u
+  ad=1.3199p pd=9.67u as=0p ps=0u
M1001 VDD.t3 A.t0 a_217_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y.t0 a_217_1050.t6 VDD.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1003 VDD.t0 B.t0 a_217_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_217_1050.t3 A.t2 VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_217_1050.t2 B.t2 VDD.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 VDD.t4 a_217_1050.t7 Y.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y a_217_1050.t5 GND.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
C0 A VDD 0.08fF
C1 B VDD 0.07fF
C2 A B 0.27fF
C3 Y VDD 0.78fF
R0 a_217_1050.n4 a_217_1050.t7 512.525
R1 a_217_1050.n4 a_217_1050.t6 371.139
R2 a_217_1050.n5 a_217_1050.t5 210.434
R3 a_217_1050.n8 a_217_1050.n6 184.039
R4 a_217_1050.n6 a_217_1050.n3 179.052
R5 a_217_1050.n5 a_217_1050.n4 173.2
R6 a_217_1050.n6 a_217_1050.n5 153.043
R7 a_217_1050.n3 a_217_1050.n2 76.002
R8 a_217_1050.n8 a_217_1050.n7 30
R9 a_217_1050.n9 a_217_1050.n0 24.383
R10 a_217_1050.n9 a_217_1050.n8 23.684
R11 a_217_1050.n1 a_217_1050.t0 14.282
R12 a_217_1050.n1 a_217_1050.t2 14.282
R13 a_217_1050.n2 a_217_1050.t4 14.282
R14 a_217_1050.n2 a_217_1050.t3 14.282
R15 a_217_1050.n3 a_217_1050.n1 12.85
R16 GND.n32 GND.n31 219.745
R17 GND.n32 GND.n30 85.529
R18 GND.n44 GND.n43 84.842
R19 GND.n9 GND.n1 76.145
R20 GND.n39 GND.n38 76
R21 GND.n9 GND.n8 76
R22 GND.n17 GND.n16 76
R23 GND.n26 GND.n25 76
R24 GND.n29 GND.n28 76
R25 GND.n36 GND.n35 76
R26 GND.n59 GND.n58 76
R27 GND.n56 GND.n55 76
R28 GND.n53 GND.n52 76
R29 GND.n50 GND.n49 76
R30 GND.n47 GND.n46 76
R31 GND.n42 GND.n41 76
R32 GND.n22 GND.t1 39.412
R33 GND.n5 GND.n4 35.01
R34 GND.n6 GND.n5 19.735
R35 GND.n14 GND.n13 19.735
R36 GND.n24 GND.n23 19.735
R37 GND.n5 GND.n3 19.017
R38 GND.n22 GND.n21 17.185
R39 GND.n35 GND.n33 14.167
R40 GND.n41 GND.n40 13.653
R41 GND.n46 GND.n45 13.653
R42 GND.n49 GND.n48 13.653
R43 GND.n52 GND.n51 13.653
R44 GND.n55 GND.n54 13.653
R45 GND.n58 GND.n57 13.653
R46 GND.n35 GND.n34 13.653
R47 GND.n28 GND.n27 13.653
R48 GND.n25 GND.n18 13.653
R49 GND.n16 GND.n15 13.653
R50 GND.n8 GND.n7 13.653
R51 GND.n3 GND.n2 7.5
R52 GND.n12 GND.n11 7.5
R53 GND.n33 GND.n32 7.312
R54 GND.n23 GND.n22 6.139
R55 GND.n20 GND.n19 4.551
R56 GND.n8 GND.n6 3.935
R57 GND.n46 GND.n44 3.935
R58 GND.n25 GND.n24 3.541
R59 GND.t1 GND.n20 2.238
R60 GND.n11 GND.n10 1.935
R61 GND.n1 GND.n0 0.596
R62 GND.n38 GND.n37 0.596
R63 GND.n13 GND.n12 0.358
R64 GND.n36 GND.n29 0.29
R65 GND.n39 GND 0.207
R66 GND.n16 GND.n14 0.196
R67 GND.n53 GND.n50 0.181
R68 GND.n17 GND.n9 0.157
R69 GND.n26 GND.n17 0.157
R70 GND.n29 GND.n26 0.145
R71 GND.n59 GND.n56 0.145
R72 GND.n56 GND.n53 0.145
R73 GND.n50 GND.n47 0.145
R74 GND.n47 GND.n42 0.145
R75 GND.n42 GND.n39 0.145
R76 GND GND.n36 0.078
R77 GND GND.n59 0.066
R78 Y.n2 Y.n1 200.754
R79 Y.n2 Y.n0 184.007
R80 Y Y.n2 76
R81 Y.n0 Y.t1 14.282
R82 Y.n0 Y.t0 14.282
R83 A.n0 A.t0 480.392
R84 A.n0 A.t2 403.272
R85 A.n1 A.t1 310.033
R86 A A.n1 76
R87 A.n1 A.n0 71.894
R88 VDD.n68 VDD.n66 144.705
R89 VDD.n26 VDD.n25 77.792
R90 VDD.n35 VDD.n34 77.792
R91 VDD.n29 VDD.n23 76.145
R92 VDD.n29 VDD.n28 76
R93 VDD.n33 VDD.n32 76
R94 VDD.n39 VDD.n38 76
R95 VDD.n43 VDD.n42 76
R96 VDD.n70 VDD.n69 76
R97 VDD.n124 VDD.n123 76
R98 VDD.n119 VDD.n118 76
R99 VDD.n114 VDD.n113 76
R100 VDD.n108 VDD.n107 76
R101 VDD.n103 VDD.n102 76
R102 VDD.n98 VDD.n97 76
R103 VDD.n93 VDD.n92 76
R104 VDD.n94 VDD.t2 55.106
R105 VDD.n37 VDD.t5 55.106
R106 VDD.n24 VDD.t4 55.106
R107 VDD.n120 VDD.t0 55.106
R108 VDD.n110 VDD.n109 40.824
R109 VDD.n59 VDD.n58 36.774
R110 VDD.n116 VDD.n115 36.608
R111 VDD.n100 VDD.n99 32.032
R112 VDD.n92 VDD.n89 21.841
R113 VDD.n23 VDD.n20 21.841
R114 VDD.n109 VDD.t1 14.282
R115 VDD.n109 VDD.t3 14.282
R116 VDD.n89 VDD.n72 14.167
R117 VDD.n72 VDD.n71 14.167
R118 VDD.n64 VDD.n45 14.167
R119 VDD.n45 VDD.n44 14.167
R120 VDD.n20 VDD.n19 14.167
R121 VDD.n19 VDD.n17 14.167
R122 VDD.n69 VDD.n65 14.167
R123 VDD.n23 VDD.n22 13.653
R124 VDD.n22 VDD.n21 13.653
R125 VDD.n28 VDD.n27 13.653
R126 VDD.n27 VDD.n26 13.653
R127 VDD.n32 VDD.n31 13.653
R128 VDD.n31 VDD.n30 13.653
R129 VDD.n38 VDD.n36 13.653
R130 VDD.n36 VDD.n35 13.653
R131 VDD.n42 VDD.n41 13.653
R132 VDD.n41 VDD.n40 13.653
R133 VDD.n69 VDD.n68 13.653
R134 VDD.n68 VDD.n67 13.653
R135 VDD.n123 VDD.n122 13.653
R136 VDD.n122 VDD.n121 13.653
R137 VDD.n118 VDD.n117 13.653
R138 VDD.n117 VDD.n116 13.653
R139 VDD.n113 VDD.n112 13.653
R140 VDD.n112 VDD.n111 13.653
R141 VDD.n107 VDD.n106 13.653
R142 VDD.n106 VDD.n105 13.653
R143 VDD.n102 VDD.n101 13.653
R144 VDD.n101 VDD.n100 13.653
R145 VDD.n97 VDD.n96 13.653
R146 VDD.n96 VDD.n95 13.653
R147 VDD.n92 VDD.n91 13.653
R148 VDD.n91 VDD.n90 13.653
R149 VDD.n4 VDD.n2 12.915
R150 VDD.n4 VDD.n3 12.66
R151 VDD.n12 VDD.n11 12.343
R152 VDD.n10 VDD.n9 12.343
R153 VDD.n7 VDD.n6 12.343
R154 VDD.n113 VDD.n110 8.658
R155 VDD.n65 VDD.n64 7.674
R156 VDD.n49 VDD.n48 7.5
R157 VDD.n52 VDD.n51 7.5
R158 VDD.n54 VDD.n53 7.5
R159 VDD.n57 VDD.n56 7.5
R160 VDD.n64 VDD.n63 7.5
R161 VDD.n84 VDD.n83 7.5
R162 VDD.n78 VDD.n77 7.5
R163 VDD.n80 VDD.n79 7.5
R164 VDD.n86 VDD.n76 7.5
R165 VDD.n86 VDD.n74 7.5
R166 VDD.n89 VDD.n88 7.5
R167 VDD.n20 VDD.n16 7.5
R168 VDD.n2 VDD.n1 7.5
R169 VDD.n6 VDD.n5 7.5
R170 VDD.n9 VDD.n8 7.5
R171 VDD.n19 VDD.n18 7.5
R172 VDD.n14 VDD.n0 7.5
R173 VDD.n87 VDD.n73 6.772
R174 VDD.n85 VDD.n82 6.772
R175 VDD.n81 VDD.n78 6.772
R176 VDD.n81 VDD.n80 6.772
R177 VDD.n85 VDD.n84 6.772
R178 VDD.n88 VDD.n87 6.772
R179 VDD.n63 VDD.n62 6.772
R180 VDD.n50 VDD.n47 6.772
R181 VDD.n55 VDD.n52 6.772
R182 VDD.n60 VDD.n57 6.772
R183 VDD.n60 VDD.n59 6.772
R184 VDD.n55 VDD.n54 6.772
R185 VDD.n50 VDD.n49 6.772
R186 VDD.n62 VDD.n46 6.772
R187 VDD.n16 VDD.n15 6.458
R188 VDD.n76 VDD.n75 6.202
R189 VDD.n105 VDD.n104 4.576
R190 VDD.n97 VDD.n94 2.754
R191 VDD.n123 VDD.n120 2.361
R192 VDD.n28 VDD.n24 1.967
R193 VDD.n38 VDD.n37 1.967
R194 VDD.n14 VDD.n7 1.329
R195 VDD.n14 VDD.n10 1.329
R196 VDD.n14 VDD.n12 1.329
R197 VDD.n14 VDD.n13 1.329
R198 VDD.n15 VDD.n14 0.696
R199 VDD.n14 VDD.n4 0.696
R200 VDD.n86 VDD.n85 0.365
R201 VDD.n86 VDD.n81 0.365
R202 VDD.n87 VDD.n86 0.365
R203 VDD.n61 VDD.n60 0.365
R204 VDD.n61 VDD.n55 0.365
R205 VDD.n61 VDD.n50 0.365
R206 VDD.n62 VDD.n61 0.365
R207 VDD.n70 VDD.n43 0.29
R208 VDD.n93 VDD 0.207
R209 VDD.n114 VDD.n108 0.181
R210 VDD.n33 VDD.n29 0.157
R211 VDD.n39 VDD.n33 0.157
R212 VDD.n43 VDD.n39 0.145
R213 VDD.n124 VDD.n119 0.145
R214 VDD.n119 VDD.n114 0.145
R215 VDD.n108 VDD.n103 0.145
R216 VDD.n103 VDD.n98 0.145
R217 VDD.n98 VDD.n93 0.145
R218 VDD VDD.n70 0.078
R219 VDD VDD.n124 0.066
R220 a_112_101.t0 a_112_101.n1 34.62
R221 a_112_101.t0 a_112_101.n0 8.137
R222 a_112_101.t0 a_112_101.n2 4.69
R223 B.n0 B.t0 472.359
R224 B.n0 B.t2 384.527
R225 B.n1 B.t1 241.172
R226 B.n1 B.n0 110.06
R227 B B.n1 76
C4 VDD GND 5.00fF
C5 a_112_101.n0 GND 0.05fF
C6 a_112_101.n1 GND 0.12fF
C7 a_112_101.n2 GND 0.04fF
C8 VDD.n0 GND 0.11fF
C9 VDD.n1 GND 0.02fF
C10 VDD.n2 GND 0.02fF
C11 VDD.n3 GND 0.04fF
C12 VDD.n4 GND 0.01fF
C13 VDD.n5 GND 0.02fF
C14 VDD.n6 GND 0.02fF
C15 VDD.n8 GND 0.02fF
C16 VDD.n9 GND 0.02fF
C17 VDD.n11 GND 0.02fF
C18 VDD.n14 GND 0.41fF
C19 VDD.n16 GND 0.03fF
C20 VDD.n17 GND 0.02fF
C21 VDD.n18 GND 0.02fF
C22 VDD.n19 GND 0.02fF
C23 VDD.n20 GND 0.03fF
C24 VDD.n21 GND 0.25fF
C25 VDD.n22 GND 0.02fF
C26 VDD.n23 GND 0.03fF
C27 VDD.n24 GND 0.05fF
C28 VDD.n25 GND 0.13fF
C29 VDD.n26 GND 0.18fF
C30 VDD.n27 GND 0.01fF
C31 VDD.n28 GND 0.01fF
C32 VDD.n29 GND 0.06fF
C33 VDD.n30 GND 0.15fF
C34 VDD.n31 GND 0.01fF
C35 VDD.n32 GND 0.02fF
C36 VDD.n33 GND 0.02fF
C37 VDD.n34 GND 0.13fF
C38 VDD.n35 GND 0.18fF
C39 VDD.n36 GND 0.01fF
C40 VDD.n37 GND 0.05fF
C41 VDD.n38 GND 0.01fF
C42 VDD.n39 GND 0.02fF
C43 VDD.n40 GND 0.25fF
C44 VDD.n41 GND 0.01fF
C45 VDD.n42 GND 0.02fF
C46 VDD.n43 GND 0.03fF
C47 VDD.n44 GND 0.02fF
C48 VDD.n45 GND 0.02fF
C49 VDD.n46 GND 0.02fF
C50 VDD.n47 GND 0.02fF
C51 VDD.n48 GND 0.02fF
C52 VDD.n49 GND 0.02fF
C53 VDD.n51 GND 0.02fF
C54 VDD.n52 GND 0.02fF
C55 VDD.n53 GND 0.02fF
C56 VDD.n54 GND 0.02fF
C57 VDD.n56 GND 0.03fF
C58 VDD.n57 GND 0.02fF
C59 VDD.n58 GND 0.17fF
C60 VDD.n59 GND 0.03fF
C61 VDD.n61 GND 0.25fF
C62 VDD.n63 GND 0.02fF
C63 VDD.n64 GND 0.02fF
C64 VDD.n65 GND 0.03fF
C65 VDD.n66 GND 0.02fF
C66 VDD.n67 GND 0.25fF
C67 VDD.n68 GND 0.01fF
C68 VDD.n69 GND 0.02fF
C69 VDD.n70 GND 0.03fF
C70 VDD.n71 GND 0.02fF
C71 VDD.n72 GND 0.02fF
C72 VDD.n73 GND 0.02fF
C73 VDD.n74 GND 0.14fF
C74 VDD.n75 GND 0.03fF
C75 VDD.n76 GND 0.02fF
C76 VDD.n77 GND 0.02fF
C77 VDD.n78 GND 0.02fF
C78 VDD.n79 GND 0.02fF
C79 VDD.n80 GND 0.02fF
C80 VDD.n82 GND 0.02fF
C81 VDD.n83 GND 0.02fF
C82 VDD.n84 GND 0.02fF
C83 VDD.n86 GND 0.41fF
C84 VDD.n88 GND 0.03fF
C85 VDD.n89 GND 0.03fF
C86 VDD.n90 GND 0.25fF
C87 VDD.n91 GND 0.02fF
C88 VDD.n92 GND 0.03fF
C89 VDD.n93 GND 0.02fF
C90 VDD.n94 GND 0.05fF
C91 VDD.n95 GND 0.22fF
C92 VDD.n96 GND 0.01fF
C93 VDD.n97 GND 0.01fF
C94 VDD.n98 GND 0.02fF
C95 VDD.n99 GND 0.12fF
C96 VDD.n100 GND 0.15fF
C97 VDD.n101 GND 0.01fF
C98 VDD.n102 GND 0.02fF
C99 VDD.n103 GND 0.02fF
C100 VDD.n104 GND 0.15fF
C101 VDD.n105 GND 0.13fF
C102 VDD.n106 GND 0.01fF
C103 VDD.n107 GND 0.02fF
C104 VDD.n108 GND 0.02fF
C105 VDD.n109 GND 0.10fF
C106 VDD.n110 GND 0.02fF
C107 VDD.n111 GND 0.27fF
C108 VDD.n112 GND 0.01fF
C109 VDD.n113 GND 0.02fF
C110 VDD.n114 GND 0.02fF
C111 VDD.n115 GND 0.12fF
C112 VDD.n116 GND 0.15fF
C113 VDD.n117 GND 0.01fF
C114 VDD.n118 GND 0.02fF
C115 VDD.n119 GND 0.02fF
C116 VDD.n120 GND 0.05fF
C117 VDD.n121 GND 0.22fF
C118 VDD.n122 GND 0.01fF
C119 VDD.n123 GND 0.01fF
C120 VDD.n124 GND 0.01fF
C121 Y.n0 GND 0.81fF
C122 Y.n1 GND 0.38fF
C123 Y.n2 GND 0.51fF
C124 a_217_1050.n0 GND 0.03fF
C125 a_217_1050.n1 GND 0.41fF
C126 a_217_1050.n2 GND 0.49fF
C127 a_217_1050.n3 GND 0.26fF
C128 a_217_1050.n4 GND 0.29fF
C129 a_217_1050.n5 GND 0.45fF
C130 a_217_1050.n6 GND 0.45fF
C131 a_217_1050.n7 GND 0.03fF
C132 a_217_1050.n8 GND 0.21fF
C133 a_217_1050.n9 GND 0.04fF
.ends
