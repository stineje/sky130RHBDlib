magic
tech sky130A
magscale 1 2
timestamp 1648156629
<< metal1 >>
rect 315 649 1297 683
rect 1647 649 2103 683
rect 95 575 636 609
rect 981 575 1967 609
use li1_M1_contact  li1_M1_contact_3
timestamp 1648061256
transform -1 0 962 0 -1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform -1 0 296 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform 1 0 666 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_6
timestamp 1648061256
transform 1 0 148 0 1 592
box -53 -33 29 33
use nand2x1_pcell  nand2x1_pcell_0
timestamp 1648064633
transform 1 0 444 0 1 0
box -84 0 750 1575
use nand2x1_pcell  nand2x1_pcell_1
timestamp 1648064633
transform 1 0 1110 0 1 0
box -84 0 750 1575
use invx1_pcell  invx1_pcell_0
timestamp 1648064504
transform 1 0 0 0 1 0
box -84 0 528 1575
use li1_M1_contact  li1_M1_contact_5
timestamp 1648061256
transform 1 0 1998 0 1 592
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_7
timestamp 1648061256
transform 1 0 2146 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_4
timestamp 1648061256
transform -1 0 1628 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_2
timestamp 1648061256
transform 1 0 1332 0 1 666
box -53 -33 29 33
use nand2x1_pcell  nand2x1_pcell_2
timestamp 1648064633
transform 1 0 1776 0 1 0
box -84 0 750 1575
<< end >>
