* SPICE3 file created from DFFSNQX1.ext - technology: sky130A

.subckt DFFSNQX1 Q D CLK SN VPB VNB
M1000 VNB a_168_157# a_112_73.t0 nshort w=-1.605u l=1.765u
+  ad=1.0746p pd=9.42u as=0p ps=0u
M1001 VNB a_343_383.t12 a_3368_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1002 Q SN VPB.t16 pshort w=2u l=0.15u
+  ad=1.74p pd=13.74u as=0p ps=0u
M1003 VPB.t22 a_168_157# a_217_1004.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPB.t2 a_1265_943.t5 a_1905_1004.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 Q a_1265_943.t6 VPB.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_1905_1004.t1 a_217_1004.t6 VPB.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPB.t19 a_343_383.t7 a_217_1004.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPB.t0 a_217_1004.t7 a_343_383.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_3473_1004.t3 Q VPB.t28 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VNB a_217_1004.t10 a_757_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1011 VNB a_1905_1004.t7 a_2702_73.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1012 Q a_1265_943.t7 a_4294_182.t1 nshort w=-1.605u l=1.765u
+  ad=0.1791p pd=1.57u as=0p ps=0u
M1013 VPB.t25 CLK a_343_383.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPB.t10 a_1905_1004.t8 a_1265_943.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_3473_1004.t1 a_343_383.t9 VPB.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPB.t11 a_3473_1004.t6 Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPB.t23 a_1265_943.t8 Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 VNB a_217_1004.t5 a_1719_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPB.t18 a_1265_943.t9 a_343_383.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_217_1004.t3 a_168_157# VPB.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1905_1004.t5 a_1265_943.t10 VPB.t17 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPB.t15 SN Q pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_217_1004.t2 a_343_383.t10 VPB.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1905_1004.t3 SN VPB.t14 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_343_383.t0 a_217_1004.t8 VPB.t7 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPB.t8 a_217_1004.t9 a_1905_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_343_383.t5 CLK VPB.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1265_943.t1 a_1905_1004.t9 VPB.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPB.t29 Q a_3473_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 VNB a_3473_1004.t5 a_4013_75.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPB.t26 CLK a_1265_943.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1032 Q a_3473_1004.t7 VPB.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_343_383.t2 a_1265_943.t13 VPB.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPB.t4 a_343_383.t11 a_3473_1004.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPB.t13 SN a_1905_1004.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1265_943.t2 CLK VPB.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
C0 VPB CLK 0.59fF
C1 VPB Q 1.84fF
C2 VPB a_168_157# 0.08fF
C3 VPB SN 0.10fF
C4 CLK SN 0.08fF
C5 Q SN 0.39fF
R0 VPB.n313 VPB.n311 94.117
R1 VPB.n227 VPB.n225 94.117
R2 VPB.n395 VPB.n393 94.117
R3 VPB.n165 VPB.n163 94.117
R4 VPB.n103 VPB.n101 94.117
R5 VPB.n25 VPB.n24 84.554
R6 VPB.n437 VPB.n436 80.104
R7 VPB.n355 VPB.n354 80.104
R8 VPB.n44 VPB.n43 76
R9 VPB.n49 VPB.n48 76
R10 VPB.n54 VPB.n53 76
R11 VPB.n61 VPB.n60 76
R12 VPB.n66 VPB.n65 76
R13 VPB.n71 VPB.n70 76
R14 VPB.n75 VPB.n74 76
R15 VPB.n79 VPB.n78 76
R16 VPB.n105 VPB.n104 76
R17 VPB.n110 VPB.n109 76
R18 VPB.n115 VPB.n114 76
R19 VPB.n122 VPB.n121 76
R20 VPB.n127 VPB.n126 76
R21 VPB.n132 VPB.n131 76
R22 VPB.n137 VPB.n136 76
R23 VPB.n141 VPB.n140 76
R24 VPB.n167 VPB.n166 76
R25 VPB.n172 VPB.n171 76
R26 VPB.n177 VPB.n176 76
R27 VPB.n184 VPB.n183 76
R28 VPB.n189 VPB.n188 76
R29 VPB.n194 VPB.n193 76
R30 VPB.n199 VPB.n198 76
R31 VPB.n203 VPB.n202 76
R32 VPB.n229 VPB.n228 76
R33 VPB.n449 VPB.n448 76
R34 VPB.n445 VPB.n444 76
R35 VPB.n440 VPB.n439 76
R36 VPB.n435 VPB.n434 76
R37 VPB.n428 VPB.n427 76
R38 VPB.n423 VPB.n422 76
R39 VPB.n418 VPB.n417 76
R40 VPB.n411 VPB.n410 76
R41 VPB.n406 VPB.n405 76
R42 VPB.n401 VPB.n400 76
R43 VPB.n397 VPB.n396 76
R44 VPB.n371 VPB.n370 76
R45 VPB.n367 VPB.n366 76
R46 VPB.n363 VPB.n362 76
R47 VPB.n358 VPB.n357 76
R48 VPB.n353 VPB.n352 76
R49 VPB.n346 VPB.n345 76
R50 VPB.n341 VPB.n340 76
R51 VPB.n336 VPB.n335 76
R52 VPB.n329 VPB.n328 76
R53 VPB.n324 VPB.n323 76
R54 VPB.n319 VPB.n318 76
R55 VPB.n315 VPB.n314 76
R56 VPB.n289 VPB.n288 76
R57 VPB.n285 VPB.n284 76
R58 VPB.n280 VPB.n279 76
R59 VPB.n275 VPB.n274 76
R60 VPB.n268 VPB.n267 76
R61 VPB.n263 VPB.n262 76
R62 VPB.n258 VPB.n257 76
R63 VPB.n256 VPB.n230 76
R64 VPB.n63 VPB.n62 75.654
R65 VPB.n408 VPB.n407 75.654
R66 VPB.n326 VPB.n325 75.654
R67 VPB.n294 VPB.n293 61.764
R68 VPB.n376 VPB.n375 61.764
R69 VPB.n208 VPB.n207 61.764
R70 VPB.n146 VPB.n145 61.764
R71 VPB.n84 VPB.n83 61.764
R72 VPB.n231 VPB.t21 55.106
R73 VPB.n320 VPB.t7 55.106
R74 VPB.n402 VPB.t9 55.106
R75 VPB.n195 VPB.t12 55.106
R76 VPB.n133 VPB.t5 55.106
R77 VPB.n67 VPB.t3 55.106
R78 VPB.n281 VPB.t19 55.106
R79 VPB.n359 VPB.t18 55.106
R80 VPB.n441 VPB.t2 55.106
R81 VPB.n168 VPB.t26 55.106
R82 VPB.n106 VPB.t29 55.106
R83 VPB.n31 VPB.t23 55.106
R84 VPB.n39 VPB.n38 48.952
R85 VPB.n112 VPB.n111 48.952
R86 VPB.n174 VPB.n173 48.952
R87 VPB.n430 VPB.n429 48.952
R88 VPB.n348 VPB.n347 48.952
R89 VPB.n277 VPB.n276 48.952
R90 VPB.n58 VPB.n57 44.502
R91 VPB.n129 VPB.n128 44.502
R92 VPB.n191 VPB.n190 44.502
R93 VPB.n415 VPB.n414 44.502
R94 VPB.n333 VPB.n332 44.502
R95 VPB.n260 VPB.n259 44.502
R96 VPB.n270 VPB.n269 40.824
R97 VPB.n331 VPB.n330 40.824
R98 VPB.n351 VPB.n350 40.824
R99 VPB.n413 VPB.n412 40.824
R100 VPB.n433 VPB.n432 40.824
R101 VPB.n179 VPB.n178 40.824
R102 VPB.n117 VPB.n116 40.824
R103 VPB.n56 VPB.n55 40.824
R104 VPB.n42 VPB.n41 40.824
R105 VPB.n36 VPB.n35 35.118
R106 VPB.n256 VPB.n253 20.452
R107 VPB.n23 VPB.n20 20.452
R108 VPB.n46 VPB.n45 17.801
R109 VPB.n119 VPB.n118 17.801
R110 VPB.n181 VPB.n180 17.801
R111 VPB.n425 VPB.n424 17.801
R112 VPB.n343 VPB.n342 17.801
R113 VPB.n272 VPB.n271 17.801
R114 VPB.n269 VPB.t20 14.282
R115 VPB.n269 VPB.t22 14.282
R116 VPB.n330 VPB.t27 14.282
R117 VPB.n330 VPB.t0 14.282
R118 VPB.n350 VPB.t6 14.282
R119 VPB.n350 VPB.t25 14.282
R120 VPB.n412 VPB.t14 14.282
R121 VPB.n412 VPB.t8 14.282
R122 VPB.n432 VPB.t17 14.282
R123 VPB.n432 VPB.t13 14.282
R124 VPB.n178 VPB.t24 14.282
R125 VPB.n178 VPB.t10 14.282
R126 VPB.n116 VPB.t28 14.282
R127 VPB.n116 VPB.t4 14.282
R128 VPB.n55 VPB.t16 14.282
R129 VPB.n55 VPB.t11 14.282
R130 VPB.n41 VPB.t1 14.282
R131 VPB.n41 VPB.t15 14.282
R132 VPB.n23 VPB.n22 13.653
R133 VPB.n22 VPB.n21 13.653
R134 VPB.n34 VPB.n33 13.653
R135 VPB.n33 VPB.n32 13.653
R136 VPB.n30 VPB.n26 13.653
R137 VPB.n26 VPB.n25 13.653
R138 VPB.n29 VPB.n28 13.653
R139 VPB.n28 VPB.n27 13.653
R140 VPB.n43 VPB.n40 13.653
R141 VPB.n40 VPB.n39 13.653
R142 VPB.n48 VPB.n47 13.653
R143 VPB.n47 VPB.n46 13.653
R144 VPB.n53 VPB.n52 13.653
R145 VPB.n52 VPB.n51 13.653
R146 VPB.n60 VPB.n59 13.653
R147 VPB.n59 VPB.n58 13.653
R148 VPB.n65 VPB.n64 13.653
R149 VPB.n64 VPB.n63 13.653
R150 VPB.n70 VPB.n69 13.653
R151 VPB.n69 VPB.n68 13.653
R152 VPB.n74 VPB.n73 13.653
R153 VPB.n73 VPB.n72 13.653
R154 VPB.n78 VPB.n77 13.653
R155 VPB.n77 VPB.n76 13.653
R156 VPB.n104 VPB.n103 13.653
R157 VPB.n103 VPB.n102 13.653
R158 VPB.n109 VPB.n108 13.653
R159 VPB.n108 VPB.n107 13.653
R160 VPB.n114 VPB.n113 13.653
R161 VPB.n113 VPB.n112 13.653
R162 VPB.n121 VPB.n120 13.653
R163 VPB.n120 VPB.n119 13.653
R164 VPB.n126 VPB.n125 13.653
R165 VPB.n125 VPB.n124 13.653
R166 VPB.n131 VPB.n130 13.653
R167 VPB.n130 VPB.n129 13.653
R168 VPB.n136 VPB.n135 13.653
R169 VPB.n135 VPB.n134 13.653
R170 VPB.n140 VPB.n139 13.653
R171 VPB.n139 VPB.n138 13.653
R172 VPB.n166 VPB.n165 13.653
R173 VPB.n165 VPB.n164 13.653
R174 VPB.n171 VPB.n170 13.653
R175 VPB.n170 VPB.n169 13.653
R176 VPB.n176 VPB.n175 13.653
R177 VPB.n175 VPB.n174 13.653
R178 VPB.n183 VPB.n182 13.653
R179 VPB.n182 VPB.n181 13.653
R180 VPB.n188 VPB.n187 13.653
R181 VPB.n187 VPB.n186 13.653
R182 VPB.n193 VPB.n192 13.653
R183 VPB.n192 VPB.n191 13.653
R184 VPB.n198 VPB.n197 13.653
R185 VPB.n197 VPB.n196 13.653
R186 VPB.n202 VPB.n201 13.653
R187 VPB.n201 VPB.n200 13.653
R188 VPB.n228 VPB.n227 13.653
R189 VPB.n227 VPB.n226 13.653
R190 VPB.n448 VPB.n447 13.653
R191 VPB.n447 VPB.n446 13.653
R192 VPB.n444 VPB.n443 13.653
R193 VPB.n443 VPB.n442 13.653
R194 VPB.n439 VPB.n438 13.653
R195 VPB.n438 VPB.n437 13.653
R196 VPB.n434 VPB.n431 13.653
R197 VPB.n431 VPB.n430 13.653
R198 VPB.n427 VPB.n426 13.653
R199 VPB.n426 VPB.n425 13.653
R200 VPB.n422 VPB.n421 13.653
R201 VPB.n421 VPB.n420 13.653
R202 VPB.n417 VPB.n416 13.653
R203 VPB.n416 VPB.n415 13.653
R204 VPB.n410 VPB.n409 13.653
R205 VPB.n409 VPB.n408 13.653
R206 VPB.n405 VPB.n404 13.653
R207 VPB.n404 VPB.n403 13.653
R208 VPB.n400 VPB.n399 13.653
R209 VPB.n399 VPB.n398 13.653
R210 VPB.n396 VPB.n395 13.653
R211 VPB.n395 VPB.n394 13.653
R212 VPB.n370 VPB.n369 13.653
R213 VPB.n369 VPB.n368 13.653
R214 VPB.n366 VPB.n365 13.653
R215 VPB.n365 VPB.n364 13.653
R216 VPB.n362 VPB.n361 13.653
R217 VPB.n361 VPB.n360 13.653
R218 VPB.n357 VPB.n356 13.653
R219 VPB.n356 VPB.n355 13.653
R220 VPB.n352 VPB.n349 13.653
R221 VPB.n349 VPB.n348 13.653
R222 VPB.n345 VPB.n344 13.653
R223 VPB.n344 VPB.n343 13.653
R224 VPB.n340 VPB.n339 13.653
R225 VPB.n339 VPB.n338 13.653
R226 VPB.n335 VPB.n334 13.653
R227 VPB.n334 VPB.n333 13.653
R228 VPB.n328 VPB.n327 13.653
R229 VPB.n327 VPB.n326 13.653
R230 VPB.n323 VPB.n322 13.653
R231 VPB.n322 VPB.n321 13.653
R232 VPB.n318 VPB.n317 13.653
R233 VPB.n317 VPB.n316 13.653
R234 VPB.n314 VPB.n313 13.653
R235 VPB.n313 VPB.n312 13.653
R236 VPB.n288 VPB.n287 13.653
R237 VPB.n287 VPB.n286 13.653
R238 VPB.n284 VPB.n283 13.653
R239 VPB.n283 VPB.n282 13.653
R240 VPB.n279 VPB.n278 13.653
R241 VPB.n278 VPB.n277 13.653
R242 VPB.n274 VPB.n273 13.653
R243 VPB.n273 VPB.n272 13.653
R244 VPB.n267 VPB.n266 13.653
R245 VPB.n266 VPB.n265 13.653
R246 VPB.n262 VPB.n261 13.653
R247 VPB.n261 VPB.n260 13.653
R248 VPB.n257 VPB.n233 13.653
R249 VPB.n233 VPB.n232 13.653
R250 VPB.n256 VPB.n255 13.653
R251 VPB.n255 VPB.n254 13.653
R252 VPB.n51 VPB.n50 13.35
R253 VPB.n124 VPB.n123 13.35
R254 VPB.n186 VPB.n185 13.35
R255 VPB.n420 VPB.n419 13.35
R256 VPB.n338 VPB.n337 13.35
R257 VPB.n265 VPB.n264 13.35
R258 VPB.n99 VPB.n82 13.276
R259 VPB.n82 VPB.n80 13.276
R260 VPB.n161 VPB.n144 13.276
R261 VPB.n144 VPB.n142 13.276
R262 VPB.n223 VPB.n206 13.276
R263 VPB.n206 VPB.n204 13.276
R264 VPB.n391 VPB.n374 13.276
R265 VPB.n374 VPB.n372 13.276
R266 VPB.n309 VPB.n292 13.276
R267 VPB.n292 VPB.n290 13.276
R268 VPB.n253 VPB.n236 13.276
R269 VPB.n236 VPB.n234 13.276
R270 VPB.n20 VPB.n19 13.276
R271 VPB.n19 VPB.n17 13.276
R272 VPB.n30 VPB.n29 13.276
R273 VPB.n104 VPB.n100 13.276
R274 VPB.n166 VPB.n162 13.276
R275 VPB.n228 VPB.n224 13.276
R276 VPB.n396 VPB.n392 13.276
R277 VPB.n314 VPB.n310 13.276
R278 VPB.n257 VPB.n256 13.276
R279 VPB.n4 VPB.n2 12.796
R280 VPB.n4 VPB.n3 12.564
R281 VPB.n34 VPB.n31 12.2
R282 VPB.n10 VPB.n9 12.198
R283 VPB.n12 VPB.n11 12.198
R284 VPB.n10 VPB.n7 12.198
R285 VPB.n236 VPB.n235 7.5
R286 VPB.n239 VPB.n238 7.5
R287 VPB.n242 VPB.n241 7.5
R288 VPB.n244 VPB.n243 7.5
R289 VPB.n247 VPB.n246 7.5
R290 VPB.n253 VPB.n252 7.5
R291 VPB.n292 VPB.n291 7.5
R292 VPB.n304 VPB.n303 7.5
R293 VPB.n298 VPB.n297 7.5
R294 VPB.n300 VPB.n299 7.5
R295 VPB.n306 VPB.n296 7.5
R296 VPB.n306 VPB.n294 7.5
R297 VPB.n309 VPB.n308 7.5
R298 VPB.n374 VPB.n373 7.5
R299 VPB.n386 VPB.n385 7.5
R300 VPB.n380 VPB.n379 7.5
R301 VPB.n382 VPB.n381 7.5
R302 VPB.n388 VPB.n378 7.5
R303 VPB.n388 VPB.n376 7.5
R304 VPB.n391 VPB.n390 7.5
R305 VPB.n206 VPB.n205 7.5
R306 VPB.n218 VPB.n217 7.5
R307 VPB.n212 VPB.n211 7.5
R308 VPB.n214 VPB.n213 7.5
R309 VPB.n220 VPB.n210 7.5
R310 VPB.n220 VPB.n208 7.5
R311 VPB.n223 VPB.n222 7.5
R312 VPB.n144 VPB.n143 7.5
R313 VPB.n156 VPB.n155 7.5
R314 VPB.n150 VPB.n149 7.5
R315 VPB.n152 VPB.n151 7.5
R316 VPB.n158 VPB.n148 7.5
R317 VPB.n158 VPB.n146 7.5
R318 VPB.n161 VPB.n160 7.5
R319 VPB.n82 VPB.n81 7.5
R320 VPB.n94 VPB.n93 7.5
R321 VPB.n88 VPB.n87 7.5
R322 VPB.n90 VPB.n89 7.5
R323 VPB.n96 VPB.n86 7.5
R324 VPB.n96 VPB.n84 7.5
R325 VPB.n99 VPB.n98 7.5
R326 VPB.n20 VPB.n16 7.5
R327 VPB.n2 VPB.n1 7.5
R328 VPB.n9 VPB.n8 7.5
R329 VPB.n7 VPB.n6 7.5
R330 VPB.n19 VPB.n18 7.5
R331 VPB.n14 VPB.n0 7.5
R332 VPB.n100 VPB.n99 7.176
R333 VPB.n162 VPB.n161 7.176
R334 VPB.n224 VPB.n223 7.176
R335 VPB.n392 VPB.n391 7.176
R336 VPB.n310 VPB.n309 7.176
R337 VPB.n305 VPB.n302 6.729
R338 VPB.n301 VPB.n298 6.729
R339 VPB.n387 VPB.n384 6.729
R340 VPB.n383 VPB.n380 6.729
R341 VPB.n219 VPB.n216 6.729
R342 VPB.n215 VPB.n212 6.729
R343 VPB.n157 VPB.n154 6.729
R344 VPB.n153 VPB.n150 6.729
R345 VPB.n95 VPB.n92 6.729
R346 VPB.n91 VPB.n88 6.729
R347 VPB.n301 VPB.n300 6.728
R348 VPB.n305 VPB.n304 6.728
R349 VPB.n308 VPB.n307 6.728
R350 VPB.n383 VPB.n382 6.728
R351 VPB.n387 VPB.n386 6.728
R352 VPB.n390 VPB.n389 6.728
R353 VPB.n215 VPB.n214 6.728
R354 VPB.n219 VPB.n218 6.728
R355 VPB.n222 VPB.n221 6.728
R356 VPB.n153 VPB.n152 6.728
R357 VPB.n157 VPB.n156 6.728
R358 VPB.n160 VPB.n159 6.728
R359 VPB.n91 VPB.n90 6.728
R360 VPB.n95 VPB.n94 6.728
R361 VPB.n98 VPB.n97 6.728
R362 VPB.n252 VPB.n251 6.728
R363 VPB.n240 VPB.n237 6.728
R364 VPB.n245 VPB.n242 6.728
R365 VPB.n249 VPB.n247 6.728
R366 VPB.n249 VPB.n248 6.728
R367 VPB.n245 VPB.n244 6.728
R368 VPB.n240 VPB.n239 6.728
R369 VPB.n121 VPB.n117 6.458
R370 VPB.n183 VPB.n179 6.458
R371 VPB.n274 VPB.n270 6.458
R372 VPB.n16 VPB.n15 6.398
R373 VPB.n296 VPB.n295 6.166
R374 VPB.n378 VPB.n377 6.166
R375 VPB.n210 VPB.n209 6.166
R376 VPB.n148 VPB.n147 6.166
R377 VPB.n86 VPB.n85 6.166
R378 VPB.n35 VPB.n23 6.112
R379 VPB.n35 VPB.n34 6.101
R380 VPB.n60 VPB.n56 4.305
R381 VPB.n417 VPB.n413 4.305
R382 VPB.n335 VPB.n331 4.305
R383 VPB.n43 VPB.n42 3.947
R384 VPB.n434 VPB.n433 3.947
R385 VPB.n352 VPB.n351 3.947
R386 VPB.n136 VPB.n133 1.794
R387 VPB.n198 VPB.n195 1.794
R388 VPB.n257 VPB.n231 1.794
R389 VPB.n109 VPB.n106 1.435
R390 VPB.n171 VPB.n168 1.435
R391 VPB.n284 VPB.n281 1.435
R392 VPB.n14 VPB.n5 1.402
R393 VPB.n14 VPB.n10 1.402
R394 VPB.n14 VPB.n12 1.402
R395 VPB.n14 VPB.n13 1.402
R396 VPB.n31 VPB.n30 1.076
R397 VPB.n444 VPB.n441 1.076
R398 VPB.n362 VPB.n359 1.076
R399 VPB.n15 VPB.n14 0.735
R400 VPB.n14 VPB.n4 0.735
R401 VPB.n70 VPB.n67 0.717
R402 VPB.n405 VPB.n402 0.717
R403 VPB.n323 VPB.n320 0.717
R404 VPB.n306 VPB.n305 0.387
R405 VPB.n306 VPB.n301 0.387
R406 VPB.n307 VPB.n306 0.387
R407 VPB.n388 VPB.n387 0.387
R408 VPB.n388 VPB.n383 0.387
R409 VPB.n389 VPB.n388 0.387
R410 VPB.n220 VPB.n219 0.387
R411 VPB.n220 VPB.n215 0.387
R412 VPB.n221 VPB.n220 0.387
R413 VPB.n158 VPB.n157 0.387
R414 VPB.n158 VPB.n153 0.387
R415 VPB.n159 VPB.n158 0.387
R416 VPB.n96 VPB.n95 0.387
R417 VPB.n96 VPB.n91 0.387
R418 VPB.n97 VPB.n96 0.387
R419 VPB.n250 VPB.n249 0.387
R420 VPB.n250 VPB.n245 0.387
R421 VPB.n250 VPB.n240 0.387
R422 VPB.n251 VPB.n250 0.387
R423 VPB.n105 VPB.n79 0.272
R424 VPB.n167 VPB.n141 0.272
R425 VPB.n229 VPB.n203 0.272
R426 VPB.n397 VPB.n371 0.272
R427 VPB.n315 VPB.n289 0.272
R428 VPB.n37 VPB.n36 0.136
R429 VPB.n44 VPB.n37 0.136
R430 VPB.n49 VPB.n44 0.136
R431 VPB.n54 VPB.n49 0.136
R432 VPB.n61 VPB.n54 0.136
R433 VPB.n66 VPB.n61 0.136
R434 VPB.n71 VPB.n66 0.136
R435 VPB.n75 VPB.n71 0.136
R436 VPB.n79 VPB.n75 0.136
R437 VPB.n110 VPB.n105 0.136
R438 VPB.n115 VPB.n110 0.136
R439 VPB.n122 VPB.n115 0.136
R440 VPB.n127 VPB.n122 0.136
R441 VPB.n132 VPB.n127 0.136
R442 VPB.n137 VPB.n132 0.136
R443 VPB.n141 VPB.n137 0.136
R444 VPB.n172 VPB.n167 0.136
R445 VPB.n177 VPB.n172 0.136
R446 VPB.n184 VPB.n177 0.136
R447 VPB.n189 VPB.n184 0.136
R448 VPB.n194 VPB.n189 0.136
R449 VPB.n199 VPB.n194 0.136
R450 VPB.n203 VPB.n199 0.136
R451 VPB.n449 VPB.n229 0.136
R452 VPB.n449 VPB.n445 0.136
R453 VPB.n445 VPB.n440 0.136
R454 VPB.n440 VPB.n435 0.136
R455 VPB.n435 VPB.n428 0.136
R456 VPB.n428 VPB.n423 0.136
R457 VPB.n423 VPB.n418 0.136
R458 VPB.n418 VPB.n411 0.136
R459 VPB.n411 VPB.n406 0.136
R460 VPB.n406 VPB.n401 0.136
R461 VPB.n401 VPB.n397 0.136
R462 VPB.n371 VPB.n367 0.136
R463 VPB.n367 VPB.n363 0.136
R464 VPB.n363 VPB.n358 0.136
R465 VPB.n358 VPB.n353 0.136
R466 VPB.n353 VPB.n346 0.136
R467 VPB.n346 VPB.n341 0.136
R468 VPB.n341 VPB.n336 0.136
R469 VPB.n336 VPB.n329 0.136
R470 VPB.n329 VPB.n324 0.136
R471 VPB.n324 VPB.n319 0.136
R472 VPB.n319 VPB.n315 0.136
R473 VPB.n289 VPB.n285 0.136
R474 VPB.n285 VPB.n280 0.136
R475 VPB.n280 VPB.n275 0.136
R476 VPB.n275 VPB.n268 0.136
R477 VPB.n268 VPB.n263 0.136
R478 VPB.n263 VPB.n258 0.136
R479 VPB.n258 VPB.n230 0.136
R480 VPB.n230 VPB 0.031
R481 a_217_1004.n5 a_217_1004.t7 512.525
R482 a_217_1004.n3 a_217_1004.t9 512.525
R483 a_217_1004.n5 a_217_1004.t8 371.139
R484 a_217_1004.n3 a_217_1004.t6 371.139
R485 a_217_1004.n6 a_217_1004.n5 226.225
R486 a_217_1004.n4 a_217_1004.n3 225.866
R487 a_217_1004.n4 a_217_1004.t5 218.057
R488 a_217_1004.n6 a_217_1004.t10 217.698
R489 a_217_1004.n8 a_217_1004.n2 215.652
R490 a_217_1004.n10 a_217_1004.n8 147.503
R491 a_217_1004.n7 a_217_1004.n4 79.488
R492 a_217_1004.n8 a_217_1004.n7 77.314
R493 a_217_1004.n2 a_217_1004.n1 76.002
R494 a_217_1004.n7 a_217_1004.n6 76
R495 a_217_1004.n10 a_217_1004.n9 15.218
R496 a_217_1004.n0 a_217_1004.t1 14.282
R497 a_217_1004.n0 a_217_1004.t2 14.282
R498 a_217_1004.n1 a_217_1004.t4 14.282
R499 a_217_1004.n1 a_217_1004.t3 14.282
R500 a_217_1004.n2 a_217_1004.n0 12.85
R501 a_217_1004.n11 a_217_1004.n10 12.014
R502 a_1265_943.n6 a_1265_943.t10 454.685
R503 a_1265_943.n8 a_1265_943.t13 454.685
R504 a_1265_943.n4 a_1265_943.t6 454.685
R505 a_1265_943.n6 a_1265_943.t5 428.979
R506 a_1265_943.n8 a_1265_943.t9 428.979
R507 a_1265_943.n4 a_1265_943.t8 428.979
R508 a_1265_943.n7 a_1265_943.t11 248.006
R509 a_1265_943.n9 a_1265_943.t12 248.006
R510 a_1265_943.n5 a_1265_943.t7 248.006
R511 a_1265_943.n14 a_1265_943.n12 220.639
R512 a_1265_943.n12 a_1265_943.n3 135.994
R513 a_1265_943.n7 a_1265_943.n6 81.941
R514 a_1265_943.n9 a_1265_943.n8 81.941
R515 a_1265_943.n5 a_1265_943.n4 81.941
R516 a_1265_943.n11 a_1265_943.n5 81.396
R517 a_1265_943.n10 a_1265_943.n9 79.491
R518 a_1265_943.n3 a_1265_943.n2 76.002
R519 a_1265_943.n10 a_1265_943.n7 76
R520 a_1265_943.n12 a_1265_943.n11 76
R521 a_1265_943.n14 a_1265_943.n13 30
R522 a_1265_943.n15 a_1265_943.n0 24.383
R523 a_1265_943.n15 a_1265_943.n14 23.684
R524 a_1265_943.n1 a_1265_943.t3 14.282
R525 a_1265_943.n1 a_1265_943.t2 14.282
R526 a_1265_943.n2 a_1265_943.t0 14.282
R527 a_1265_943.n2 a_1265_943.t1 14.282
R528 a_1265_943.n3 a_1265_943.n1 12.85
R529 a_1265_943.n11 a_1265_943.n10 2.947
R530 a_1905_1004.n6 a_1905_1004.t8 480.392
R531 a_1905_1004.n6 a_1905_1004.t9 403.272
R532 a_1905_1004.n8 a_1905_1004.n5 233.952
R533 a_1905_1004.n7 a_1905_1004.t7 213.869
R534 a_1905_1004.n7 a_1905_1004.n6 161.6
R535 a_1905_1004.n8 a_1905_1004.n7 153.315
R536 a_1905_1004.n10 a_1905_1004.n8 143.492
R537 a_1905_1004.n4 a_1905_1004.n3 79.232
R538 a_1905_1004.n5 a_1905_1004.n4 63.152
R539 a_1905_1004.n10 a_1905_1004.n9 30
R540 a_1905_1004.n11 a_1905_1004.n0 24.383
R541 a_1905_1004.n11 a_1905_1004.n10 23.684
R542 a_1905_1004.n5 a_1905_1004.n1 16.08
R543 a_1905_1004.n4 a_1905_1004.n2 16.08
R544 a_1905_1004.n1 a_1905_1004.t6 14.282
R545 a_1905_1004.n1 a_1905_1004.t5 14.282
R546 a_1905_1004.n2 a_1905_1004.t2 14.282
R547 a_1905_1004.n2 a_1905_1004.t3 14.282
R548 a_1905_1004.n3 a_1905_1004.t0 14.282
R549 a_1905_1004.n3 a_1905_1004.t1 14.282
R550 a_1719_75.t0 a_1719_75.n3 117.777
R551 a_1719_75.n6 a_1719_75.n5 45.444
R552 a_1719_75.t0 a_1719_75.n6 21.213
R553 a_1719_75.t0 a_1719_75.n4 11.595
R554 a_1719_75.n2 a_1719_75.n0 8.543
R555 a_1719_75.t0 a_1719_75.n2 3.034
R556 a_1719_75.n2 a_1719_75.n1 0.443
R557 VNB VNB.n391 300.778
R558 VNB.n215 VNB.n214 199.897
R559 VNB.n100 VNB.n99 199.897
R560 VNB.n80 VNB.n79 199.897
R561 VNB.n322 VNB.n321 199.897
R562 VNB.n18 VNB.n17 199.897
R563 VNB.n112 VNB.n110 154.509
R564 VNB.n224 VNB.n222 154.509
R565 VNB.n331 VNB.n329 154.509
R566 VNB.n265 VNB.n263 154.509
R567 VNB.n44 VNB.n42 154.509
R568 VNB.n363 VNB.n362 147.75
R569 VNB.n124 VNB.n123 121.366
R570 VNB.n30 VNB.n28 121.366
R571 VNB.n56 VNB.n55 121.366
R572 VNB.n192 VNB.n191 85.559
R573 VNB.n299 VNB.n298 85.559
R574 VNB.n244 VNB.n243 84.842
R575 VNB.n269 VNB.n69 76
R576 VNB.n378 VNB.n377 76
R577 VNB.n366 VNB.n365 76
R578 VNB.n361 VNB.n360 76
R579 VNB.n357 VNB.n356 76
R580 VNB.n353 VNB.n352 76
R581 VNB.n349 VNB.n348 76
R582 VNB.n345 VNB.n344 76
R583 VNB.n341 VNB.n340 76
R584 VNB.n337 VNB.n336 76
R585 VNB.n333 VNB.n332 76
R586 VNB.n311 VNB.n310 76
R587 VNB.n307 VNB.n306 76
R588 VNB.n303 VNB.n302 76
R589 VNB.n297 VNB.n296 76
R590 VNB.n293 VNB.n292 76
R591 VNB.n289 VNB.n288 76
R592 VNB.n285 VNB.n284 76
R593 VNB.n281 VNB.n280 76
R594 VNB.n277 VNB.n276 76
R595 VNB.n273 VNB.n272 76
R596 VNB.n266 VNB.n262 76
R597 VNB.n252 VNB.n251 76
R598 VNB.n248 VNB.n247 76
R599 VNB.n242 VNB.n241 76
R600 VNB.n238 VNB.n237 76
R601 VNB.n234 VNB.n233 76
R602 VNB.n230 VNB.n229 76
R603 VNB.n226 VNB.n225 76
R604 VNB.n204 VNB.n203 76
R605 VNB.n200 VNB.n199 76
R606 VNB.n196 VNB.n195 76
R607 VNB.n190 VNB.n189 76
R608 VNB.n186 VNB.n185 76
R609 VNB.n182 VNB.n181 76
R610 VNB.n178 VNB.n177 76
R611 VNB.n174 VNB.n173 76
R612 VNB.n35 VNB.n34 73.875
R613 VNB.n33 VNB.n27 64.552
R614 VNB.n128 VNB.n89 63.835
R615 VNB.n60 VNB.n7 63.835
R616 VNB.n194 VNB.n193 41.971
R617 VNB.n301 VNB.n300 41.971
R618 VNB.n125 VNB.n124 36.937
R619 VNB.n30 VNB.n29 36.937
R620 VNB.n57 VNB.n56 36.937
R621 VNB.n246 VNB.n245 36.678
R622 VNB.n169 VNB.n168 35.118
R623 VNB.n89 VNB.n88 28.421
R624 VNB.n27 VNB.n26 28.421
R625 VNB.n7 VNB.n6 28.421
R626 VNB.n131 VNB.n130 27.855
R627 VNB.n63 VNB.n62 27.855
R628 VNB.n89 VNB.n87 25.263
R629 VNB.n27 VNB.n25 25.263
R630 VNB.n7 VNB.n5 25.263
R631 VNB.n87 VNB.n86 24.383
R632 VNB.n25 VNB.n24 24.383
R633 VNB.n5 VNB.n4 24.383
R634 VNB.n158 VNB.n155 20.452
R635 VNB.n379 VNB.n378 20.452
R636 VNB.n132 VNB.n131 16.721
R637 VNB.n64 VNB.n63 16.721
R638 VNB.n167 VNB.n166 13.653
R639 VNB.n166 VNB.n165 13.653
R640 VNB.n164 VNB.n163 13.653
R641 VNB.n163 VNB.n162 13.653
R642 VNB.n161 VNB.n160 13.653
R643 VNB.n160 VNB.n159 13.653
R644 VNB.n173 VNB.n172 13.653
R645 VNB.n172 VNB.n171 13.653
R646 VNB.n177 VNB.n176 13.653
R647 VNB.n176 VNB.n175 13.653
R648 VNB.n181 VNB.n180 13.653
R649 VNB.n180 VNB.n179 13.653
R650 VNB.n185 VNB.n184 13.653
R651 VNB.n184 VNB.n183 13.653
R652 VNB.n189 VNB.n188 13.653
R653 VNB.n188 VNB.n187 13.653
R654 VNB.n195 VNB.n194 13.653
R655 VNB.n199 VNB.n198 13.653
R656 VNB.n198 VNB.n197 13.653
R657 VNB.n203 VNB.n202 13.653
R658 VNB.n202 VNB.n201 13.653
R659 VNB.n225 VNB.n224 13.653
R660 VNB.n224 VNB.n223 13.653
R661 VNB.n229 VNB.n228 13.653
R662 VNB.n228 VNB.n227 13.653
R663 VNB.n233 VNB.n232 13.653
R664 VNB.n232 VNB.n231 13.653
R665 VNB.n237 VNB.n236 13.653
R666 VNB.n236 VNB.n235 13.653
R667 VNB.n241 VNB.n240 13.653
R668 VNB.n240 VNB.n239 13.653
R669 VNB.n247 VNB.n246 13.653
R670 VNB.n251 VNB.n250 13.653
R671 VNB.n250 VNB.n249 13.653
R672 VNB.n108 VNB.n107 13.653
R673 VNB.n107 VNB.n106 13.653
R674 VNB.n113 VNB.n112 13.653
R675 VNB.n112 VNB.n111 13.653
R676 VNB.n116 VNB.n115 13.653
R677 VNB.n115 VNB.n114 13.653
R678 VNB.n119 VNB.n118 13.653
R679 VNB.n118 VNB.n117 13.653
R680 VNB.n122 VNB.n121 13.653
R681 VNB.n121 VNB.n120 13.653
R682 VNB.n127 VNB.n126 13.653
R683 VNB.n126 VNB.n125 13.653
R684 VNB.n133 VNB.n132 13.653
R685 VNB.n136 VNB.n135 13.653
R686 VNB.n135 VNB.n134 13.653
R687 VNB.n139 VNB.n138 13.653
R688 VNB.n138 VNB.n137 13.653
R689 VNB.n266 VNB.n265 13.653
R690 VNB.n265 VNB.n264 13.653
R691 VNB.n269 VNB.n268 13.653
R692 VNB.n268 VNB.n267 13.653
R693 VNB.n272 VNB.n271 13.653
R694 VNB.n271 VNB.n270 13.653
R695 VNB.n276 VNB.n275 13.653
R696 VNB.n275 VNB.n274 13.653
R697 VNB.n280 VNB.n279 13.653
R698 VNB.n279 VNB.n278 13.653
R699 VNB.n284 VNB.n283 13.653
R700 VNB.n283 VNB.n282 13.653
R701 VNB.n288 VNB.n287 13.653
R702 VNB.n287 VNB.n286 13.653
R703 VNB.n292 VNB.n291 13.653
R704 VNB.n291 VNB.n290 13.653
R705 VNB.n296 VNB.n295 13.653
R706 VNB.n295 VNB.n294 13.653
R707 VNB.n302 VNB.n301 13.653
R708 VNB.n306 VNB.n305 13.653
R709 VNB.n305 VNB.n304 13.653
R710 VNB.n310 VNB.n309 13.653
R711 VNB.n309 VNB.n308 13.653
R712 VNB.n332 VNB.n331 13.653
R713 VNB.n331 VNB.n330 13.653
R714 VNB.n336 VNB.n335 13.653
R715 VNB.n335 VNB.n334 13.653
R716 VNB.n340 VNB.n339 13.653
R717 VNB.n339 VNB.n338 13.653
R718 VNB.n344 VNB.n343 13.653
R719 VNB.n343 VNB.n342 13.653
R720 VNB.n348 VNB.n347 13.653
R721 VNB.n347 VNB.n346 13.653
R722 VNB.n352 VNB.n351 13.653
R723 VNB.n351 VNB.n350 13.653
R724 VNB.n356 VNB.n355 13.653
R725 VNB.n355 VNB.n354 13.653
R726 VNB.n360 VNB.n359 13.653
R727 VNB.n359 VNB.n358 13.653
R728 VNB.n365 VNB.n364 13.653
R729 VNB.n364 VNB.n363 13.653
R730 VNB.n32 VNB.n31 13.653
R731 VNB.n31 VNB.n30 13.653
R732 VNB.n37 VNB.n36 13.653
R733 VNB.n36 VNB.n35 13.653
R734 VNB.n40 VNB.n39 13.653
R735 VNB.n39 VNB.n38 13.653
R736 VNB.n45 VNB.n44 13.653
R737 VNB.n44 VNB.n43 13.653
R738 VNB.n48 VNB.n47 13.653
R739 VNB.n47 VNB.n46 13.653
R740 VNB.n51 VNB.n50 13.653
R741 VNB.n50 VNB.n49 13.653
R742 VNB.n54 VNB.n53 13.653
R743 VNB.n53 VNB.n52 13.653
R744 VNB.n59 VNB.n58 13.653
R745 VNB.n58 VNB.n57 13.653
R746 VNB.n65 VNB.n64 13.653
R747 VNB.n68 VNB.n67 13.653
R748 VNB.n67 VNB.n66 13.653
R749 VNB.n378 VNB.n0 13.653
R750 VNB VNB.n0 13.653
R751 VNB.n158 VNB.n157 13.653
R752 VNB.n157 VNB.n156 13.653
R753 VNB.n386 VNB.n383 13.577
R754 VNB.n143 VNB.n141 13.276
R755 VNB.n155 VNB.n143 13.276
R756 VNB.n207 VNB.n205 13.276
R757 VNB.n220 VNB.n207 13.276
R758 VNB.n92 VNB.n90 13.276
R759 VNB.n105 VNB.n92 13.276
R760 VNB.n72 VNB.n70 13.276
R761 VNB.n85 VNB.n72 13.276
R762 VNB.n314 VNB.n312 13.276
R763 VNB.n327 VNB.n314 13.276
R764 VNB.n10 VNB.n8 13.276
R765 VNB.n23 VNB.n10 13.276
R766 VNB.n167 VNB.n164 13.276
R767 VNB.n164 VNB.n161 13.276
R768 VNB.n225 VNB.n221 13.276
R769 VNB.n109 VNB.n108 13.276
R770 VNB.n113 VNB.n109 13.276
R771 VNB.n116 VNB.n113 13.276
R772 VNB.n119 VNB.n116 13.276
R773 VNB.n122 VNB.n119 13.276
R774 VNB.n127 VNB.n122 13.276
R775 VNB.n136 VNB.n133 13.276
R776 VNB.n139 VNB.n136 13.276
R777 VNB.n140 VNB.n139 13.276
R778 VNB.n266 VNB.n140 13.276
R779 VNB.n269 VNB.n266 13.276
R780 VNB.n272 VNB.n269 13.276
R781 VNB.n332 VNB.n328 13.276
R782 VNB.n40 VNB.n37 13.276
R783 VNB.n41 VNB.n40 13.276
R784 VNB.n45 VNB.n41 13.276
R785 VNB.n48 VNB.n45 13.276
R786 VNB.n51 VNB.n48 13.276
R787 VNB.n54 VNB.n51 13.276
R788 VNB.n59 VNB.n54 13.276
R789 VNB.n68 VNB.n65 13.276
R790 VNB.n378 VNB.n68 13.276
R791 VNB.n3 VNB.n1 13.276
R792 VNB.n379 VNB.n3 13.276
R793 VNB.n37 VNB.n33 12.02
R794 VNB.n128 VNB.n127 10.764
R795 VNB.n60 VNB.n59 10.764
R796 VNB.n388 VNB.n387 7.5
R797 VNB.n213 VNB.n212 7.5
R798 VNB.n209 VNB.n208 7.5
R799 VNB.n207 VNB.n206 7.5
R800 VNB.n220 VNB.n219 7.5
R801 VNB.n98 VNB.n97 7.5
R802 VNB.n94 VNB.n93 7.5
R803 VNB.n92 VNB.n91 7.5
R804 VNB.n105 VNB.n104 7.5
R805 VNB.n78 VNB.n77 7.5
R806 VNB.n74 VNB.n73 7.5
R807 VNB.n72 VNB.n71 7.5
R808 VNB.n85 VNB.n84 7.5
R809 VNB.n320 VNB.n319 7.5
R810 VNB.n316 VNB.n315 7.5
R811 VNB.n314 VNB.n313 7.5
R812 VNB.n327 VNB.n326 7.5
R813 VNB.n16 VNB.n15 7.5
R814 VNB.n12 VNB.n11 7.5
R815 VNB.n10 VNB.n9 7.5
R816 VNB.n23 VNB.n22 7.5
R817 VNB.n380 VNB.n379 7.5
R818 VNB.n3 VNB.n2 7.5
R819 VNB.n385 VNB.n384 7.5
R820 VNB.n149 VNB.n148 7.5
R821 VNB.n145 VNB.n144 7.5
R822 VNB.n143 VNB.n142 7.5
R823 VNB.n155 VNB.n154 7.5
R824 VNB.n221 VNB.n220 7.176
R825 VNB.n109 VNB.n105 7.176
R826 VNB.n140 VNB.n85 7.176
R827 VNB.n328 VNB.n327 7.176
R828 VNB.n41 VNB.n23 7.176
R829 VNB.n390 VNB.n388 7.011
R830 VNB.n216 VNB.n213 7.011
R831 VNB.n211 VNB.n209 7.011
R832 VNB.n101 VNB.n98 7.011
R833 VNB.n96 VNB.n94 7.011
R834 VNB.n81 VNB.n78 7.011
R835 VNB.n76 VNB.n74 7.011
R836 VNB.n323 VNB.n320 7.011
R837 VNB.n318 VNB.n316 7.011
R838 VNB.n19 VNB.n16 7.011
R839 VNB.n14 VNB.n12 7.011
R840 VNB.n151 VNB.n149 7.011
R841 VNB.n147 VNB.n145 7.011
R842 VNB.n219 VNB.n218 7.01
R843 VNB.n211 VNB.n210 7.01
R844 VNB.n216 VNB.n215 7.01
R845 VNB.n104 VNB.n103 7.01
R846 VNB.n96 VNB.n95 7.01
R847 VNB.n101 VNB.n100 7.01
R848 VNB.n84 VNB.n83 7.01
R849 VNB.n76 VNB.n75 7.01
R850 VNB.n81 VNB.n80 7.01
R851 VNB.n326 VNB.n325 7.01
R852 VNB.n318 VNB.n317 7.01
R853 VNB.n323 VNB.n322 7.01
R854 VNB.n22 VNB.n21 7.01
R855 VNB.n14 VNB.n13 7.01
R856 VNB.n19 VNB.n18 7.01
R857 VNB.n154 VNB.n153 7.01
R858 VNB.n147 VNB.n146 7.01
R859 VNB.n151 VNB.n150 7.01
R860 VNB.n390 VNB.n389 7.01
R861 VNB.n386 VNB.n385 6.788
R862 VNB.n381 VNB.n380 6.788
R863 VNB.n168 VNB.n158 6.111
R864 VNB.n168 VNB.n167 6.1
R865 VNB.n247 VNB.n244 2.511
R866 VNB.n133 VNB.n128 2.511
R867 VNB.n65 VNB.n60 2.511
R868 VNB.n131 VNB.n129 1.99
R869 VNB.n63 VNB.n61 1.99
R870 VNB.n195 VNB.n192 1.255
R871 VNB.n302 VNB.n299 1.255
R872 VNB.n33 VNB.n32 1.255
R873 VNB.n391 VNB.n382 0.921
R874 VNB.n391 VNB.n386 0.476
R875 VNB.n391 VNB.n381 0.475
R876 VNB.n226 VNB.n204 0.272
R877 VNB.n254 VNB.n253 0.272
R878 VNB.n262 VNB.n261 0.272
R879 VNB.n333 VNB.n311 0.272
R880 VNB.n370 VNB.n369 0.272
R881 VNB.n217 VNB.n211 0.246
R882 VNB.n218 VNB.n217 0.246
R883 VNB.n217 VNB.n216 0.246
R884 VNB.n102 VNB.n96 0.246
R885 VNB.n103 VNB.n102 0.246
R886 VNB.n102 VNB.n101 0.246
R887 VNB.n82 VNB.n76 0.246
R888 VNB.n83 VNB.n82 0.246
R889 VNB.n82 VNB.n81 0.246
R890 VNB.n324 VNB.n318 0.246
R891 VNB.n325 VNB.n324 0.246
R892 VNB.n324 VNB.n323 0.246
R893 VNB.n20 VNB.n14 0.246
R894 VNB.n21 VNB.n20 0.246
R895 VNB.n20 VNB.n19 0.246
R896 VNB.n152 VNB.n147 0.246
R897 VNB.n153 VNB.n152 0.246
R898 VNB.n152 VNB.n151 0.246
R899 VNB.n391 VNB.n390 0.246
R900 VNB.n377 VNB 0.198
R901 VNB.n170 VNB.n169 0.136
R902 VNB.n174 VNB.n170 0.136
R903 VNB.n178 VNB.n174 0.136
R904 VNB.n182 VNB.n178 0.136
R905 VNB.n186 VNB.n182 0.136
R906 VNB.n190 VNB.n186 0.136
R907 VNB.n196 VNB.n190 0.136
R908 VNB.n200 VNB.n196 0.136
R909 VNB.n204 VNB.n200 0.136
R910 VNB.n230 VNB.n226 0.136
R911 VNB.n234 VNB.n230 0.136
R912 VNB.n238 VNB.n234 0.136
R913 VNB.n242 VNB.n238 0.136
R914 VNB.n248 VNB.n242 0.136
R915 VNB.n252 VNB.n248 0.136
R916 VNB.n253 VNB.n252 0.136
R917 VNB.n255 VNB.n254 0.136
R918 VNB.n256 VNB.n255 0.136
R919 VNB.n257 VNB.n256 0.136
R920 VNB.n258 VNB.n257 0.136
R921 VNB.n259 VNB.n258 0.136
R922 VNB.n260 VNB.n259 0.136
R923 VNB.n261 VNB.n260 0.136
R924 VNB.n262 VNB.n69 0.136
R925 VNB.n273 VNB.n69 0.136
R926 VNB.n277 VNB.n273 0.136
R927 VNB.n281 VNB.n277 0.136
R928 VNB.n285 VNB.n281 0.136
R929 VNB.n289 VNB.n285 0.136
R930 VNB.n293 VNB.n289 0.136
R931 VNB.n297 VNB.n293 0.136
R932 VNB.n303 VNB.n297 0.136
R933 VNB.n307 VNB.n303 0.136
R934 VNB.n311 VNB.n307 0.136
R935 VNB.n337 VNB.n333 0.136
R936 VNB.n341 VNB.n337 0.136
R937 VNB.n345 VNB.n341 0.136
R938 VNB.n349 VNB.n345 0.136
R939 VNB.n353 VNB.n349 0.136
R940 VNB.n357 VNB.n353 0.136
R941 VNB.n361 VNB.n357 0.136
R942 VNB.n366 VNB.n361 0.136
R943 VNB.n367 VNB.n366 0.136
R944 VNB.n368 VNB.n367 0.136
R945 VNB.n369 VNB.n368 0.136
R946 VNB.n371 VNB.n370 0.136
R947 VNB.n372 VNB.n371 0.136
R948 VNB.n373 VNB.n372 0.136
R949 VNB.n374 VNB.n373 0.136
R950 VNB.n375 VNB.n374 0.136
R951 VNB.n376 VNB.n375 0.136
R952 VNB.n377 VNB.n376 0.136
R953 a_757_75.n4 a_757_75.n3 19.724
R954 a_757_75.t0 a_757_75.n5 11.595
R955 a_757_75.t0 a_757_75.n4 9.207
R956 a_757_75.n2 a_757_75.n0 8.543
R957 a_757_75.t0 a_757_75.n2 3.034
R958 a_757_75.n2 a_757_75.n1 0.443
R959 a_1038_182.n12 a_1038_182.n5 96.467
R960 a_1038_182.t0 a_1038_182.n1 46.91
R961 a_1038_182.n9 a_1038_182.n7 34.805
R962 a_1038_182.n9 a_1038_182.n8 32.622
R963 a_1038_182.t0 a_1038_182.n12 32.417
R964 a_1038_182.n5 a_1038_182.n4 22.349
R965 a_1038_182.n11 a_1038_182.n9 19.017
R966 a_1038_182.n1 a_1038_182.n0 17.006
R967 a_1038_182.n5 a_1038_182.n3 8.443
R968 a_1038_182.t0 a_1038_182.n2 8.137
R969 a_1038_182.n7 a_1038_182.n6 7.5
R970 a_1038_182.n11 a_1038_182.n10 7.5
R971 a_1038_182.n12 a_1038_182.n11 1.435
R972 a_343_383.n6 a_343_383.t11 480.392
R973 a_343_383.n8 a_343_383.t7 472.359
R974 a_343_383.n6 a_343_383.t9 403.272
R975 a_343_383.n8 a_343_383.t10 384.527
R976 a_343_383.n7 a_343_383.t12 320.08
R977 a_343_383.n9 a_343_383.t8 277.772
R978 a_343_383.n13 a_343_383.n11 249.364
R979 a_343_383.n11 a_343_383.n5 127.401
R980 a_343_383.n10 a_343_383.n7 83.304
R981 a_343_383.n10 a_343_383.n9 80.032
R982 a_343_383.n4 a_343_383.n3 79.232
R983 a_343_383.n11 a_343_383.n10 76
R984 a_343_383.n9 a_343_383.n8 67.001
R985 a_343_383.n5 a_343_383.n4 63.152
R986 a_343_383.n7 a_343_383.n6 55.388
R987 a_343_383.n14 a_343_383.n0 55.263
R988 a_343_383.n13 a_343_383.n12 30
R989 a_343_383.n14 a_343_383.n13 23.684
R990 a_343_383.n5 a_343_383.n1 16.08
R991 a_343_383.n4 a_343_383.n2 16.08
R992 a_343_383.n1 a_343_383.t3 14.282
R993 a_343_383.n1 a_343_383.t2 14.282
R994 a_343_383.n2 a_343_383.t6 14.282
R995 a_343_383.n2 a_343_383.t5 14.282
R996 a_343_383.n3 a_343_383.t1 14.282
R997 a_343_383.n3 a_343_383.t0 14.282
R998 a_2702_73.n12 a_2702_73.n11 26.811
R999 a_2702_73.n6 a_2702_73.n5 24.977
R1000 a_2702_73.n2 a_2702_73.n1 24.877
R1001 a_2702_73.t0 a_2702_73.n2 12.677
R1002 a_2702_73.t0 a_2702_73.n3 11.595
R1003 a_2702_73.t1 a_2702_73.n8 8.137
R1004 a_2702_73.t0 a_2702_73.n4 7.273
R1005 a_2702_73.t0 a_2702_73.n0 6.109
R1006 a_2702_73.t1 a_2702_73.n7 4.864
R1007 a_2702_73.t0 a_2702_73.n12 2.074
R1008 a_2702_73.n7 a_2702_73.n6 1.13
R1009 a_2702_73.n12 a_2702_73.t1 0.937
R1010 a_2702_73.t1 a_2702_73.n10 0.804
R1011 a_2702_73.n10 a_2702_73.n9 0.136
R1012 a_3473_1004.n4 a_3473_1004.t6 512.525
R1013 a_3473_1004.n4 a_3473_1004.t7 371.139
R1014 a_3473_1004.n5 a_3473_1004.t5 244.609
R1015 a_3473_1004.n5 a_3473_1004.n4 199.313
R1016 a_3473_1004.n6 a_3473_1004.n3 189.099
R1017 a_3473_1004.n8 a_3473_1004.n6 167.533
R1018 a_3473_1004.n6 a_3473_1004.n5 153.315
R1019 a_3473_1004.n3 a_3473_1004.n2 76.002
R1020 a_3473_1004.n8 a_3473_1004.n7 30
R1021 a_3473_1004.n9 a_3473_1004.n0 24.383
R1022 a_3473_1004.n9 a_3473_1004.n8 23.684
R1023 a_3473_1004.n1 a_3473_1004.t2 14.282
R1024 a_3473_1004.n1 a_3473_1004.t3 14.282
R1025 a_3473_1004.n2 a_3473_1004.t0 14.282
R1026 a_3473_1004.n2 a_3473_1004.t1 14.282
R1027 a_3473_1004.n3 a_3473_1004.n1 12.85
R1028 a_112_73.t0 a_112_73.n1 34.62
R1029 a_112_73.t0 a_112_73.n0 8.137
R1030 a_112_73.t0 a_112_73.n2 4.69
R1031 a_4294_182.n10 a_4294_182.n8 82.852
R1032 a_4294_182.n7 a_4294_182.n6 32.833
R1033 a_4294_182.n8 a_4294_182.t1 32.416
R1034 a_4294_182.n10 a_4294_182.n9 27.2
R1035 a_4294_182.n11 a_4294_182.n0 23.498
R1036 a_4294_182.n3 a_4294_182.n2 23.284
R1037 a_4294_182.n11 a_4294_182.n10 22.4
R1038 a_4294_182.n7 a_4294_182.n4 19.017
R1039 a_4294_182.n6 a_4294_182.n5 13.494
R1040 a_4294_182.t1 a_4294_182.n1 7.04
R1041 a_4294_182.t1 a_4294_182.n3 5.727
R1042 a_4294_182.n8 a_4294_182.n7 1.435
R1043 a_2000_182.n10 a_2000_182.n8 82.852
R1044 a_2000_182.n11 a_2000_182.n0 49.6
R1045 a_2000_182.n7 a_2000_182.n6 32.833
R1046 a_2000_182.n8 a_2000_182.t1 32.416
R1047 a_2000_182.n10 a_2000_182.n9 27.2
R1048 a_2000_182.n3 a_2000_182.n2 23.284
R1049 a_2000_182.n11 a_2000_182.n10 22.4
R1050 a_2000_182.n7 a_2000_182.n4 19.017
R1051 a_2000_182.n6 a_2000_182.n5 13.494
R1052 a_2000_182.t1 a_2000_182.n1 7.04
R1053 a_2000_182.t1 a_2000_182.n3 5.727
R1054 a_2000_182.n8 a_2000_182.n7 1.435
R1055 a_3368_73.n12 a_3368_73.n11 26.811
R1056 a_3368_73.n6 a_3368_73.n5 24.977
R1057 a_3368_73.n2 a_3368_73.n1 24.877
R1058 a_3368_73.t0 a_3368_73.n2 12.677
R1059 a_3368_73.t0 a_3368_73.n3 11.595
R1060 a_3368_73.t1 a_3368_73.n8 8.137
R1061 a_3368_73.t0 a_3368_73.n4 7.273
R1062 a_3368_73.t0 a_3368_73.n0 6.109
R1063 a_3368_73.t1 a_3368_73.n7 4.864
R1064 a_3368_73.t0 a_3368_73.n12 2.074
R1065 a_3368_73.n7 a_3368_73.n6 1.13
R1066 a_3368_73.n12 a_3368_73.t1 0.937
R1067 a_3368_73.t1 a_3368_73.n10 0.804
R1068 a_3368_73.n10 a_3368_73.n9 0.136
R1069 a_4013_75.n5 a_4013_75.n4 19.724
R1070 a_4013_75.t0 a_4013_75.n3 11.595
R1071 a_4013_75.t0 a_4013_75.n5 9.207
R1072 a_4013_75.n2 a_4013_75.n1 2.455
R1073 a_4013_75.n2 a_4013_75.n0 1.32
R1074 a_4013_75.t0 a_4013_75.n2 0.246
C6 VPB VNB 18.74fF
C7 a_4013_75.n0 VNB 0.10fF
C8 a_4013_75.n1 VNB 0.04fF
C9 a_4013_75.n2 VNB 0.03fF
C10 a_4013_75.n3 VNB 0.07fF
C11 a_4013_75.n4 VNB 0.08fF
C12 a_4013_75.n5 VNB 0.06fF
C13 a_3368_73.n0 VNB 0.02fF
C14 a_3368_73.n1 VNB 0.10fF
C15 a_3368_73.n2 VNB 0.06fF
C16 a_3368_73.n3 VNB 0.06fF
C17 a_3368_73.n4 VNB 0.00fF
C18 a_3368_73.n5 VNB 0.04fF
C19 a_3368_73.n6 VNB 0.05fF
C20 a_3368_73.n7 VNB 0.02fF
C21 a_3368_73.n8 VNB 0.05fF
C22 a_3368_73.n9 VNB 0.08fF
C23 a_3368_73.n10 VNB 0.17fF
C24 a_3368_73.t1 VNB 0.23fF
C25 a_3368_73.n11 VNB 0.09fF
C26 a_3368_73.n12 VNB 0.00fF
C27 a_2000_182.n0 VNB 0.02fF
C28 a_2000_182.n1 VNB 0.09fF
C29 a_2000_182.n2 VNB 0.13fF
C30 a_2000_182.n3 VNB 0.11fF
C31 a_2000_182.t1 VNB 0.30fF
C32 a_2000_182.n4 VNB 0.09fF
C33 a_2000_182.n5 VNB 0.06fF
C34 a_2000_182.n6 VNB 0.01fF
C35 a_2000_182.n7 VNB 0.03fF
C36 a_2000_182.n8 VNB 0.11fF
C37 a_2000_182.n9 VNB 0.02fF
C38 a_2000_182.n10 VNB 0.05fF
C39 a_2000_182.n11 VNB 0.02fF
C40 a_4294_182.n0 VNB 0.02fF
C41 a_4294_182.n1 VNB 0.09fF
C42 a_4294_182.n2 VNB 0.13fF
C43 a_4294_182.n3 VNB 0.11fF
C44 a_4294_182.n4 VNB 0.09fF
C45 a_4294_182.n5 VNB 0.05fF
C46 a_4294_182.n6 VNB 0.01fF
C47 a_4294_182.n7 VNB 0.03fF
C48 a_4294_182.n8 VNB 0.11fF
C49 a_4294_182.n9 VNB 0.02fF
C50 a_4294_182.n10 VNB 0.05fF
C51 a_4294_182.n11 VNB 0.03fF
C52 a_112_73.n0 VNB 0.05fF
C53 a_112_73.n1 VNB 0.12fF
C54 a_112_73.n2 VNB 0.04fF
C55 a_3473_1004.n0 VNB 0.04fF
C56 a_3473_1004.n1 VNB 0.51fF
C57 a_3473_1004.n2 VNB 0.61fF
C58 a_3473_1004.n3 VNB 0.34fF
C59 a_3473_1004.n4 VNB 0.37fF
C60 a_3473_1004.n5 VNB 0.62fF
C61 a_3473_1004.n6 VNB 0.58fF
C62 a_3473_1004.n7 VNB 0.03fF
C63 a_3473_1004.n8 VNB 0.24fF
C64 a_3473_1004.n9 VNB 0.05fF
C65 a_2702_73.n0 VNB 0.02fF
C66 a_2702_73.n1 VNB 0.10fF
C67 a_2702_73.n2 VNB 0.06fF
C68 a_2702_73.n3 VNB 0.06fF
C69 a_2702_73.n4 VNB 0.00fF
C70 a_2702_73.n5 VNB 0.04fF
C71 a_2702_73.n6 VNB 0.05fF
C72 a_2702_73.n7 VNB 0.02fF
C73 a_2702_73.n8 VNB 0.05fF
C74 a_2702_73.n9 VNB 0.08fF
C75 a_2702_73.n10 VNB 0.17fF
C76 a_2702_73.t1 VNB 0.23fF
C77 a_2702_73.n11 VNB 0.09fF
C78 a_2702_73.n12 VNB 0.00fF
C79 a_343_383.n0 VNB 0.05fF
C80 a_343_383.n1 VNB 0.68fF
C81 a_343_383.n2 VNB 0.68fF
C82 a_343_383.n3 VNB 0.80fF
C83 a_343_383.n4 VNB 0.25fF
C84 a_343_383.n5 VNB 0.32fF
C85 a_343_383.n6 VNB 0.41fF
C86 a_343_383.n7 VNB 0.59fF
C87 a_343_383.n8 VNB 0.36fF
C88 a_343_383.t8 VNB 0.72fF
C89 a_343_383.n9 VNB 0.50fF
C90 a_343_383.n10 VNB 3.16fF
C91 a_343_383.n11 VNB 0.56fF
C92 a_343_383.n12 VNB 0.05fF
C93 a_343_383.n13 VNB 0.43fF
C94 a_343_383.n14 VNB 0.06fF
C95 a_1038_182.n0 VNB 0.07fF
C96 a_1038_182.n1 VNB 0.13fF
C97 a_1038_182.n2 VNB 0.07fF
C98 a_1038_182.n3 VNB 0.02fF
C99 a_1038_182.n4 VNB 0.03fF
C100 a_1038_182.n5 VNB 0.06fF
C101 a_1038_182.n6 VNB 0.05fF
C102 a_1038_182.n7 VNB 0.06fF
C103 a_1038_182.n8 VNB 0.07fF
C104 a_1038_182.n9 VNB 0.07fF
C105 a_1038_182.n10 VNB 0.03fF
C106 a_1038_182.n11 VNB 0.01fF
C107 a_1038_182.n12 VNB 0.12fF
C108 a_1038_182.t0 VNB 0.28fF
C109 a_757_75.n0 VNB 0.20fF
C110 a_757_75.n1 VNB 0.04fF
C111 a_757_75.n2 VNB 0.01fF
C112 a_757_75.n3 VNB 0.08fF
C113 a_757_75.n4 VNB 0.06fF
C114 a_757_75.n5 VNB 0.07fF
C115 a_1719_75.n0 VNB 0.20fF
C116 a_1719_75.n1 VNB 0.04fF
C117 a_1719_75.n2 VNB 0.01fF
C118 a_1719_75.n3 VNB 0.03fF
C119 a_1719_75.n4 VNB 0.05fF
C120 a_1719_75.n5 VNB 0.09fF
C121 a_1719_75.n6 VNB 0.07fF
C122 a_1905_1004.n0 VNB 0.04fF
C123 a_1905_1004.n1 VNB 0.48fF
C124 a_1905_1004.n2 VNB 0.48fF
C125 a_1905_1004.n3 VNB 0.57fF
C126 a_1905_1004.n4 VNB 0.18fF
C127 a_1905_1004.n5 VNB 0.34fF
C128 a_1905_1004.n6 VNB 0.40fF
C129 a_1905_1004.n7 VNB 0.49fF
C130 a_1905_1004.n8 VNB 0.56fF
C131 a_1905_1004.n9 VNB 0.03fF
C132 a_1905_1004.n10 VNB 0.20fF
C133 a_1905_1004.n11 VNB 0.05fF
C134 a_1265_943.n0 VNB 0.05fF
C135 a_1265_943.n1 VNB 0.65fF
C136 a_1265_943.n2 VNB 0.76fF
C137 a_1265_943.n3 VNB 0.35fF
C138 a_1265_943.n4 VNB 0.43fF
C139 a_1265_943.n5 VNB 0.49fF
C140 a_1265_943.n6 VNB 0.43fF
C141 a_1265_943.t11 VNB 0.66fF
C142 a_1265_943.n7 VNB 0.44fF
C143 a_1265_943.n8 VNB 0.43fF
C144 a_1265_943.t12 VNB 0.66fF
C145 a_1265_943.n9 VNB 0.46fF
C146 a_1265_943.n10 VNB 1.39fF
C147 a_1265_943.n11 VNB 1.87fF
C148 a_1265_943.n12 VNB 0.51fF
C149 a_1265_943.n13 VNB 0.04fF
C150 a_1265_943.n14 VNB 0.38fF
C151 a_1265_943.n15 VNB 0.07fF
C152 a_217_1004.n0 VNB 0.42fF
C153 a_217_1004.n1 VNB 0.50fF
C154 a_217_1004.n2 VNB 0.30fF
C155 a_217_1004.n3 VNB 0.33fF
C156 a_217_1004.n4 VNB 0.38fF
C157 a_217_1004.n5 VNB 0.33fF
C158 a_217_1004.n6 VNB 0.36fF
C159 a_217_1004.n7 VNB 0.90fF
C160 a_217_1004.n8 VNB 0.34fF
C161 a_217_1004.n9 VNB 0.07fF
C162 a_217_1004.n10 VNB 0.16fF
C163 a_217_1004.n11 VNB 0.04fF
C164 VPB.n0 VNB 0.18fF
C165 VPB.n1 VNB 0.03fF
C166 VPB.n2 VNB 0.02fF
C167 VPB.n3 VNB 0.05fF
C168 VPB.n4 VNB 0.01fF
C169 VPB.n6 VNB 0.02fF
C170 VPB.n7 VNB 0.02fF
C171 VPB.n8 VNB 0.02fF
C172 VPB.n9 VNB 0.02fF
C173 VPB.n11 VNB 0.02fF
C174 VPB.n14 VNB 0.45fF
C175 VPB.n16 VNB 0.04fF
C176 VPB.n17 VNB 0.02fF
C177 VPB.n18 VNB 0.02fF
C178 VPB.n19 VNB 0.02fF
C179 VPB.n20 VNB 0.04fF
C180 VPB.n21 VNB 0.27fF
C181 VPB.n22 VNB 0.03fF
C182 VPB.n23 VNB 0.03fF
C183 VPB.n24 VNB 0.13fF
C184 VPB.n25 VNB 0.20fF
C185 VPB.n26 VNB 0.02fF
C186 VPB.n27 VNB 0.16fF
C187 VPB.n28 VNB 0.02fF
C188 VPB.n29 VNB 0.02fF
C189 VPB.n30 VNB 0.01fF
C190 VPB.n31 VNB 0.05fF
C191 VPB.n32 VNB 0.27fF
C192 VPB.n33 VNB 0.02fF
C193 VPB.n34 VNB 0.02fF
C194 VPB.n35 VNB 0.00fF
C195 VPB.n36 VNB 0.09fF
C196 VPB.n37 VNB 0.02fF
C197 VPB.n38 VNB 0.13fF
C198 VPB.n39 VNB 0.16fF
C199 VPB.n40 VNB 0.02fF
C200 VPB.n41 VNB 0.10fF
C201 VPB.n42 VNB 0.02fF
C202 VPB.n43 VNB 0.02fF
C203 VPB.n44 VNB 0.02fF
C204 VPB.n45 VNB 0.13fF
C205 VPB.n46 VNB 0.15fF
C206 VPB.n47 VNB 0.02fF
C207 VPB.n48 VNB 0.02fF
C208 VPB.n49 VNB 0.02fF
C209 VPB.n50 VNB 0.13fF
C210 VPB.n51 VNB 0.14fF
C211 VPB.n52 VNB 0.02fF
C212 VPB.n53 VNB 0.02fF
C213 VPB.n54 VNB 0.02fF
C214 VPB.n55 VNB 0.10fF
C215 VPB.n56 VNB 0.02fF
C216 VPB.n57 VNB 0.13fF
C217 VPB.n58 VNB 0.16fF
C218 VPB.n59 VNB 0.02fF
C219 VPB.n60 VNB 0.02fF
C220 VPB.n61 VNB 0.02fF
C221 VPB.n62 VNB 0.13fF
C222 VPB.n63 VNB 0.16fF
C223 VPB.n64 VNB 0.02fF
C224 VPB.n65 VNB 0.02fF
C225 VPB.n66 VNB 0.02fF
C226 VPB.n67 VNB 0.06fF
C227 VPB.n68 VNB 0.21fF
C228 VPB.n69 VNB 0.02fF
C229 VPB.n70 VNB 0.01fF
C230 VPB.n71 VNB 0.02fF
C231 VPB.n72 VNB 0.27fF
C232 VPB.n73 VNB 0.02fF
C233 VPB.n74 VNB 0.02fF
C234 VPB.n75 VNB 0.02fF
C235 VPB.n76 VNB 0.27fF
C236 VPB.n77 VNB 0.01fF
C237 VPB.n78 VNB 0.02fF
C238 VPB.n79 VNB 0.04fF
C239 VPB.n80 VNB 0.02fF
C240 VPB.n81 VNB 0.02fF
C241 VPB.n82 VNB 0.02fF
C242 VPB.n83 VNB 0.24fF
C243 VPB.n84 VNB 0.04fF
C244 VPB.n85 VNB 0.03fF
C245 VPB.n86 VNB 0.02fF
C246 VPB.n87 VNB 0.02fF
C247 VPB.n88 VNB 0.02fF
C248 VPB.n89 VNB 0.03fF
C249 VPB.n90 VNB 0.02fF
C250 VPB.n92 VNB 0.02fF
C251 VPB.n93 VNB 0.02fF
C252 VPB.n94 VNB 0.02fF
C253 VPB.n96 VNB 0.27fF
C254 VPB.n98 VNB 0.03fF
C255 VPB.n99 VNB 0.02fF
C256 VPB.n100 VNB 0.03fF
C257 VPB.n101 VNB 0.03fF
C258 VPB.n102 VNB 0.27fF
C259 VPB.n103 VNB 0.01fF
C260 VPB.n104 VNB 0.02fF
C261 VPB.n105 VNB 0.04fF
C262 VPB.n106 VNB 0.05fF
C263 VPB.n107 VNB 0.23fF
C264 VPB.n108 VNB 0.02fF
C265 VPB.n109 VNB 0.01fF
C266 VPB.n110 VNB 0.02fF
C267 VPB.n111 VNB 0.13fF
C268 VPB.n112 VNB 0.16fF
C269 VPB.n113 VNB 0.02fF
C270 VPB.n114 VNB 0.02fF
C271 VPB.n115 VNB 0.02fF
C272 VPB.n116 VNB 0.10fF
C273 VPB.n117 VNB 0.02fF
C274 VPB.n118 VNB 0.13fF
C275 VPB.n119 VNB 0.15fF
C276 VPB.n120 VNB 0.02fF
C277 VPB.n121 VNB 0.02fF
C278 VPB.n122 VNB 0.02fF
C279 VPB.n123 VNB 0.13fF
C280 VPB.n124 VNB 0.14fF
C281 VPB.n125 VNB 0.02fF
C282 VPB.n126 VNB 0.02fF
C283 VPB.n127 VNB 0.02fF
C284 VPB.n128 VNB 0.13fF
C285 VPB.n129 VNB 0.16fF
C286 VPB.n130 VNB 0.02fF
C287 VPB.n131 VNB 0.02fF
C288 VPB.n132 VNB 0.02fF
C289 VPB.n133 VNB 0.06fF
C290 VPB.n134 VNB 0.23fF
C291 VPB.n135 VNB 0.02fF
C292 VPB.n136 VNB 0.01fF
C293 VPB.n137 VNB 0.02fF
C294 VPB.n138 VNB 0.27fF
C295 VPB.n139 VNB 0.01fF
C296 VPB.n140 VNB 0.02fF
C297 VPB.n141 VNB 0.04fF
C298 VPB.n142 VNB 0.02fF
C299 VPB.n143 VNB 0.02fF
C300 VPB.n144 VNB 0.02fF
C301 VPB.n145 VNB 0.19fF
C302 VPB.n146 VNB 0.04fF
C303 VPB.n147 VNB 0.03fF
C304 VPB.n148 VNB 0.02fF
C305 VPB.n149 VNB 0.02fF
C306 VPB.n150 VNB 0.02fF
C307 VPB.n151 VNB 0.03fF
C308 VPB.n152 VNB 0.02fF
C309 VPB.n154 VNB 0.02fF
C310 VPB.n155 VNB 0.02fF
C311 VPB.n156 VNB 0.02fF
C312 VPB.n158 VNB 0.27fF
C313 VPB.n160 VNB 0.03fF
C314 VPB.n161 VNB 0.02fF
C315 VPB.n162 VNB 0.03fF
C316 VPB.n163 VNB 0.03fF
C317 VPB.n164 VNB 0.27fF
C318 VPB.n165 VNB 0.01fF
C319 VPB.n166 VNB 0.02fF
C320 VPB.n167 VNB 0.04fF
C321 VPB.n168 VNB 0.05fF
C322 VPB.n169 VNB 0.23fF
C323 VPB.n170 VNB 0.02fF
C324 VPB.n171 VNB 0.01fF
C325 VPB.n172 VNB 0.02fF
C326 VPB.n173 VNB 0.13fF
C327 VPB.n174 VNB 0.16fF
C328 VPB.n175 VNB 0.02fF
C329 VPB.n176 VNB 0.02fF
C330 VPB.n177 VNB 0.02fF
C331 VPB.n178 VNB 0.10fF
C332 VPB.n179 VNB 0.02fF
C333 VPB.n180 VNB 0.13fF
C334 VPB.n181 VNB 0.15fF
C335 VPB.n182 VNB 0.02fF
C336 VPB.n183 VNB 0.02fF
C337 VPB.n184 VNB 0.02fF
C338 VPB.n185 VNB 0.13fF
C339 VPB.n186 VNB 0.14fF
C340 VPB.n187 VNB 0.02fF
C341 VPB.n188 VNB 0.02fF
C342 VPB.n189 VNB 0.02fF
C343 VPB.n190 VNB 0.13fF
C344 VPB.n191 VNB 0.16fF
C345 VPB.n192 VNB 0.02fF
C346 VPB.n193 VNB 0.02fF
C347 VPB.n194 VNB 0.02fF
C348 VPB.n195 VNB 0.06fF
C349 VPB.n196 VNB 0.23fF
C350 VPB.n197 VNB 0.02fF
C351 VPB.n198 VNB 0.01fF
C352 VPB.n199 VNB 0.02fF
C353 VPB.n200 VNB 0.27fF
C354 VPB.n201 VNB 0.01fF
C355 VPB.n202 VNB 0.02fF
C356 VPB.n203 VNB 0.04fF
C357 VPB.n204 VNB 0.02fF
C358 VPB.n205 VNB 0.02fF
C359 VPB.n206 VNB 0.02fF
C360 VPB.n207 VNB 0.23fF
C361 VPB.n208 VNB 0.04fF
C362 VPB.n209 VNB 0.03fF
C363 VPB.n210 VNB 0.02fF
C364 VPB.n211 VNB 0.02fF
C365 VPB.n212 VNB 0.02fF
C366 VPB.n213 VNB 0.03fF
C367 VPB.n214 VNB 0.02fF
C368 VPB.n216 VNB 0.02fF
C369 VPB.n217 VNB 0.02fF
C370 VPB.n218 VNB 0.02fF
C371 VPB.n220 VNB 0.27fF
C372 VPB.n222 VNB 0.03fF
C373 VPB.n223 VNB 0.02fF
C374 VPB.n224 VNB 0.03fF
C375 VPB.n225 VNB 0.03fF
C376 VPB.n226 VNB 0.27fF
C377 VPB.n227 VNB 0.01fF
C378 VPB.n228 VNB 0.02fF
C379 VPB.n229 VNB 0.04fF
C380 VPB.n230 VNB 0.01fF
C381 VPB.n231 VNB 0.06fF
C382 VPB.n232 VNB 0.23fF
C383 VPB.n233 VNB 0.02fF
C384 VPB.n234 VNB 0.02fF
C385 VPB.n235 VNB 0.02fF
C386 VPB.n236 VNB 0.02fF
C387 VPB.n237 VNB 0.02fF
C388 VPB.n238 VNB 0.02fF
C389 VPB.n239 VNB 0.02fF
C390 VPB.n241 VNB 0.02fF
C391 VPB.n242 VNB 0.02fF
C392 VPB.n243 VNB 0.02fF
C393 VPB.n244 VNB 0.02fF
C394 VPB.n246 VNB 0.04fF
C395 VPB.n247 VNB 0.02fF
C396 VPB.n248 VNB 0.14fF
C397 VPB.n250 VNB 0.45fF
C398 VPB.n252 VNB 0.04fF
C399 VPB.n253 VNB 0.04fF
C400 VPB.n254 VNB 0.27fF
C401 VPB.n255 VNB 0.03fF
C402 VPB.n256 VNB 0.03fF
C403 VPB.n257 VNB 0.01fF
C404 VPB.n258 VNB 0.02fF
C405 VPB.n259 VNB 0.13fF
C406 VPB.n260 VNB 0.16fF
C407 VPB.n261 VNB 0.02fF
C408 VPB.n262 VNB 0.02fF
C409 VPB.n263 VNB 0.02fF
C410 VPB.n264 VNB 0.13fF
C411 VPB.n265 VNB 0.14fF
C412 VPB.n266 VNB 0.02fF
C413 VPB.n267 VNB 0.02fF
C414 VPB.n268 VNB 0.02fF
C415 VPB.n269 VNB 0.10fF
C416 VPB.n270 VNB 0.02fF
C417 VPB.n271 VNB 0.13fF
C418 VPB.n272 VNB 0.15fF
C419 VPB.n273 VNB 0.02fF
C420 VPB.n274 VNB 0.02fF
C421 VPB.n275 VNB 0.02fF
C422 VPB.n276 VNB 0.13fF
C423 VPB.n277 VNB 0.16fF
C424 VPB.n278 VNB 0.02fF
C425 VPB.n279 VNB 0.02fF
C426 VPB.n280 VNB 0.02fF
C427 VPB.n281 VNB 0.05fF
C428 VPB.n282 VNB 0.23fF
C429 VPB.n283 VNB 0.02fF
C430 VPB.n284 VNB 0.01fF
C431 VPB.n285 VNB 0.02fF
C432 VPB.n286 VNB 0.27fF
C433 VPB.n287 VNB 0.01fF
C434 VPB.n288 VNB 0.02fF
C435 VPB.n289 VNB 0.04fF
C436 VPB.n290 VNB 0.02fF
C437 VPB.n291 VNB 0.02fF
C438 VPB.n292 VNB 0.02fF
C439 VPB.n293 VNB 0.24fF
C440 VPB.n294 VNB 0.04fF
C441 VPB.n295 VNB 0.03fF
C442 VPB.n296 VNB 0.02fF
C443 VPB.n297 VNB 0.02fF
C444 VPB.n298 VNB 0.02fF
C445 VPB.n299 VNB 0.03fF
C446 VPB.n300 VNB 0.02fF
C447 VPB.n302 VNB 0.02fF
C448 VPB.n303 VNB 0.02fF
C449 VPB.n304 VNB 0.02fF
C450 VPB.n306 VNB 0.27fF
C451 VPB.n308 VNB 0.03fF
C452 VPB.n309 VNB 0.02fF
C453 VPB.n310 VNB 0.03fF
C454 VPB.n311 VNB 0.03fF
C455 VPB.n312 VNB 0.27fF
C456 VPB.n313 VNB 0.01fF
C457 VPB.n314 VNB 0.02fF
C458 VPB.n315 VNB 0.04fF
C459 VPB.n316 VNB 0.27fF
C460 VPB.n317 VNB 0.02fF
C461 VPB.n318 VNB 0.02fF
C462 VPB.n319 VNB 0.02fF
C463 VPB.n320 VNB 0.06fF
C464 VPB.n321 VNB 0.21fF
C465 VPB.n322 VNB 0.02fF
C466 VPB.n323 VNB 0.01fF
C467 VPB.n324 VNB 0.02fF
C468 VPB.n325 VNB 0.13fF
C469 VPB.n326 VNB 0.16fF
C470 VPB.n327 VNB 0.02fF
C471 VPB.n328 VNB 0.02fF
C472 VPB.n329 VNB 0.02fF
C473 VPB.n330 VNB 0.10fF
C474 VPB.n331 VNB 0.02fF
C475 VPB.n332 VNB 0.13fF
C476 VPB.n333 VNB 0.16fF
C477 VPB.n334 VNB 0.02fF
C478 VPB.n335 VNB 0.02fF
C479 VPB.n336 VNB 0.02fF
C480 VPB.n337 VNB 0.13fF
C481 VPB.n338 VNB 0.14fF
C482 VPB.n339 VNB 0.02fF
C483 VPB.n340 VNB 0.02fF
C484 VPB.n341 VNB 0.02fF
C485 VPB.n342 VNB 0.13fF
C486 VPB.n343 VNB 0.15fF
C487 VPB.n344 VNB 0.02fF
C488 VPB.n345 VNB 0.02fF
C489 VPB.n346 VNB 0.02fF
C490 VPB.n347 VNB 0.13fF
C491 VPB.n348 VNB 0.16fF
C492 VPB.n349 VNB 0.02fF
C493 VPB.n350 VNB 0.10fF
C494 VPB.n351 VNB 0.02fF
C495 VPB.n352 VNB 0.02fF
C496 VPB.n353 VNB 0.02fF
C497 VPB.n354 VNB 0.13fF
C498 VPB.n355 VNB 0.16fF
C499 VPB.n356 VNB 0.02fF
C500 VPB.n357 VNB 0.02fF
C501 VPB.n358 VNB 0.02fF
C502 VPB.n359 VNB 0.05fF
C503 VPB.n360 VNB 0.20fF
C504 VPB.n361 VNB 0.02fF
C505 VPB.n362 VNB 0.01fF
C506 VPB.n363 VNB 0.02fF
C507 VPB.n364 VNB 0.27fF
C508 VPB.n365 VNB 0.02fF
C509 VPB.n366 VNB 0.02fF
C510 VPB.n367 VNB 0.02fF
C511 VPB.n368 VNB 0.27fF
C512 VPB.n369 VNB 0.01fF
C513 VPB.n370 VNB 0.02fF
C514 VPB.n371 VNB 0.04fF
C515 VPB.n372 VNB 0.02fF
C516 VPB.n373 VNB 0.02fF
C517 VPB.n374 VNB 0.02fF
C518 VPB.n375 VNB 0.28fF
C519 VPB.n376 VNB 0.04fF
C520 VPB.n377 VNB 0.03fF
C521 VPB.n378 VNB 0.02fF
C522 VPB.n379 VNB 0.02fF
C523 VPB.n380 VNB 0.02fF
C524 VPB.n381 VNB 0.03fF
C525 VPB.n382 VNB 0.02fF
C526 VPB.n384 VNB 0.02fF
C527 VPB.n385 VNB 0.02fF
C528 VPB.n386 VNB 0.02fF
C529 VPB.n388 VNB 0.27fF
C530 VPB.n390 VNB 0.03fF
C531 VPB.n391 VNB 0.02fF
C532 VPB.n392 VNB 0.03fF
C533 VPB.n393 VNB 0.03fF
C534 VPB.n394 VNB 0.27fF
C535 VPB.n395 VNB 0.01fF
C536 VPB.n396 VNB 0.02fF
C537 VPB.n397 VNB 0.04fF
C538 VPB.n398 VNB 0.27fF
C539 VPB.n399 VNB 0.02fF
C540 VPB.n400 VNB 0.02fF
C541 VPB.n401 VNB 0.02fF
C542 VPB.n402 VNB 0.06fF
C543 VPB.n403 VNB 0.21fF
C544 VPB.n404 VNB 0.02fF
C545 VPB.n405 VNB 0.01fF
C546 VPB.n406 VNB 0.02fF
C547 VPB.n407 VNB 0.13fF
C548 VPB.n408 VNB 0.16fF
C549 VPB.n409 VNB 0.02fF
C550 VPB.n410 VNB 0.02fF
C551 VPB.n411 VNB 0.02fF
C552 VPB.n412 VNB 0.10fF
C553 VPB.n413 VNB 0.02fF
C554 VPB.n414 VNB 0.13fF
C555 VPB.n415 VNB 0.16fF
C556 VPB.n416 VNB 0.02fF
C557 VPB.n417 VNB 0.02fF
C558 VPB.n418 VNB 0.02fF
C559 VPB.n419 VNB 0.13fF
C560 VPB.n420 VNB 0.14fF
C561 VPB.n421 VNB 0.02fF
C562 VPB.n422 VNB 0.02fF
C563 VPB.n423 VNB 0.02fF
C564 VPB.n424 VNB 0.13fF
C565 VPB.n425 VNB 0.15fF
C566 VPB.n426 VNB 0.02fF
C567 VPB.n427 VNB 0.02fF
C568 VPB.n428 VNB 0.02fF
C569 VPB.n429 VNB 0.13fF
C570 VPB.n430 VNB 0.16fF
C571 VPB.n431 VNB 0.02fF
C572 VPB.n432 VNB 0.10fF
C573 VPB.n433 VNB 0.02fF
C574 VPB.n434 VNB 0.02fF
C575 VPB.n435 VNB 0.02fF
C576 VPB.n436 VNB 0.13fF
C577 VPB.n437 VNB 0.16fF
C578 VPB.n438 VNB 0.02fF
C579 VPB.n439 VNB 0.02fF
C580 VPB.n440 VNB 0.02fF
C581 VPB.n441 VNB 0.05fF
C582 VPB.n442 VNB 0.20fF
C583 VPB.n443 VNB 0.02fF
C584 VPB.n444 VNB 0.01fF
C585 VPB.n445 VNB 0.02fF
C586 VPB.n446 VNB 0.27fF
C587 VPB.n447 VNB 0.02fF
C588 VPB.n448 VNB 0.02fF
C589 VPB.n449 VNB 0.02fF
.ends
