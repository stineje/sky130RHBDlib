magic
tech sky130A
magscale 1 2
timestamp 1645210163
use sky130_fd_pr__hvdfm1sd__example_55959141808200  sky130_fd_pr__hvdfm1sd__example_55959141808200_0
timestamp 1645210163
transform 1 0 296 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808449  sky130_fd_pr__hvdfm1sd2__example_55959141808449_0
timestamp 1645210163
transform 1 0 120 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 324 85 324 85 0 FreeSans 300 0 0 0 S
flabel comment s 148 85 148 85 0 FreeSans 300 0 0 0 D
flabel comment s -25 100 -25 100 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 48852408
string GDS_START 48850988
<< end >>
