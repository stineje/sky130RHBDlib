magic
tech sky130A
magscale 1 2
timestamp 1652474524
<< nwell >>
rect 57 1463 91 1497
<< pwell >>
rect 57 -17 91 17
<< locali >>
rect 4349 945 4383 979
rect 5015 945 5049 979
rect 427 871 461 905
rect 3017 871 3051 905
rect 4201 871 4235 905
rect 4349 871 4383 905
rect 4719 871 4753 905
rect 5015 871 5049 905
rect 5015 797 5049 831
rect 427 723 461 757
rect 3979 723 4013 757
rect 4201 723 4235 757
rect 5015 723 5049 757
rect 427 649 461 683
rect 3017 649 3051 683
rect 3979 649 4013 683
rect 4201 649 4235 683
rect 4349 649 4383 683
rect 4719 649 4753 683
rect 5015 649 5049 683
rect 427 575 461 609
rect 1389 575 1423 609
rect 1611 575 1645 609
rect 3017 575 3051 609
rect 3979 575 4013 609
rect 4201 575 4235 609
rect 4349 575 4383 609
rect 4719 575 4753 609
rect 5015 575 5049 609
rect 427 501 461 535
rect 1389 501 1423 535
rect 1611 501 1645 535
rect 3017 501 3051 535
rect 3979 501 4013 535
rect 4201 501 4235 535
rect 4349 501 4383 535
rect 4719 501 4753 535
rect 5015 501 5049 535
rect 427 427 461 461
rect 1389 427 1423 461
rect 1611 427 1645 461
rect 3017 427 3051 461
rect 3979 427 4013 461
rect 4201 427 4235 461
rect 4349 427 4383 461
rect 5015 427 5049 461
<< metal1 >>
rect -34 1446 5214 1514
rect 4271 723 4979 757
rect 4419 649 4683 683
rect -34 -34 5214 34
use li1_M1_contact  li1_M1_contact_2 pcells
timestamp 1648061256
transform -1 0 4366 0 -1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_1
timestamp 1648061256
transform 1 0 4736 0 1 666
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_13
timestamp 1648061256
transform 1 0 5032 0 1 740
box -53 -33 29 33
use li1_M1_contact  li1_M1_contact_0
timestamp 1648061256
transform -1 0 4218 0 -1 740
box -53 -33 29 33
use dffrnx1_pcell  dffrnx1_pcell_0 pcells
timestamp 1652425808
transform 1 0 0 0 1 0
box -87 -34 5267 1550
<< labels >>
rlabel locali 5015 723 5049 757 1 Q
port 1 nsew signal output
rlabel locali 4349 649 4383 683 1 QN
port 2 nsew signal output
rlabel locali 1389 575 1423 609 1 D
port 3 nsew signal input
rlabel locali 427 871 461 905 1 CLK
port 4 nsew signal input
rlabel locali 1611 427 1645 461 1 RN
port 5 nsew signal input
rlabel locali 427 723 461 757 1 CLK
port 4 nsew signal input
rlabel locali 427 649 461 683 1 CLK
port 4 nsew signal input
rlabel locali 427 575 461 609 1 CLK
port 4 nsew signal input
rlabel locali 427 501 461 535 1 CLK
port 4 nsew signal input
rlabel locali 427 427 461 461 1 CLK
port 4 nsew signal input
rlabel locali 3017 649 3051 683 1 CLK
port 4 nsew signal input
rlabel locali 3017 575 3051 609 1 CLK
port 4 nsew signal input
rlabel locali 3017 501 3051 535 1 CLK
port 4 nsew signal input
rlabel locali 3017 427 3051 461 1 CLK
port 4 nsew signal input
rlabel locali 3017 871 3051 905 1 CLK
port 4 nsew signal input
rlabel locali 1389 501 1423 535 1 D
port 3 nsew signal input
rlabel locali 1389 427 1423 461 1 D
port 3 nsew signal input
rlabel locali 5015 797 5049 831 1 Q
port 1 nsew signal output
rlabel locali 5015 871 5049 905 1 Q
port 1 nsew signal output
rlabel locali 5015 945 5049 979 1 Q
port 1 nsew signal output
rlabel locali 5015 649 5049 683 1 Q
port 1 nsew signal output
rlabel locali 5015 575 5049 609 1 Q
port 1 nsew signal output
rlabel locali 5015 501 5049 535 1 Q
port 1 nsew signal output
rlabel locali 5015 427 5049 461 1 Q
port 1 nsew signal output
rlabel locali 4201 871 4235 905 1 Q
port 1 nsew signal output
rlabel locali 4201 723 4235 757 1 Q
port 1 nsew signal output
rlabel locali 4201 649 4235 683 1 Q
port 1 nsew signal output
rlabel locali 4201 575 4235 609 1 Q
port 1 nsew signal output
rlabel locali 4201 501 4235 535 1 Q
port 1 nsew signal output
rlabel locali 4201 427 4235 461 1 Q
port 1 nsew signal output
rlabel locali 4349 575 4383 609 1 QN
port 2 nsew signal output
rlabel locali 4349 501 4383 535 1 QN
port 2 nsew signal output
rlabel locali 4349 427 4383 461 1 QN
port 2 nsew signal output
rlabel locali 4349 945 4383 979 1 QN
port 2 nsew signal output
rlabel locali 4349 871 4383 905 1 QN
port 2 nsew signal output
rlabel locali 4719 649 4753 683 1 QN
port 2 nsew signal output
rlabel locali 4719 575 4753 609 1 QN
port 2 nsew signal output
rlabel locali 4719 501 4753 535 1 QN
port 2 nsew signal output
rlabel locali 4719 871 4753 905 1 QN
port 2 nsew signal output
rlabel locali 1611 501 1645 535 1 RN
port 5 nsew signal input
rlabel locali 1611 575 1645 609 1 RN
port 5 nsew signal input
rlabel locali 3979 427 4013 461 1 RN
port 5 nsew signal input
rlabel locali 3979 501 4013 535 1 RN
port 5 nsew signal input
rlabel locali 3979 575 4013 609 1 RN
port 5 nsew signal input
rlabel locali 3979 649 4013 683 1 RN
port 5 nsew signal input
rlabel locali 3979 723 4013 757 1 RN
port 5 nsew signal input
rlabel metal1 -34 1446 5214 1514 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 -34 -34 5214 34 1 GND
port 6 nsew ground bidirectional abutment
<< properties >>
string LEFclass CORE
string LEFsite unitrh
string FIXED_BBOX 0 0 5180 1480
string LEFsymmetry X Y R90
<< end >>
