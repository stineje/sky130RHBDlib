* SPICE3 file created from TMRDFFSNRNQNX1.ext - technology: sky130A

.subckt TMRDFFSNRNQNX1 QN D CLK SN RN VDD GND
M1000 VDD.t48 a_10219_989.t7 a_17533_1051.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1001 a_15669_1050.t5 a_15991_989.t7 VDD.t43 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1002 GND a_6049_1050.t8 a_7787_103.t0 nshort w=-1.605u l=1.765u
+  ad=3.7611p pd=32.97u as=0p ps=0u
M1003 VDD.t102 a_11821_1050.t7 a_12143_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_13105_989.t2 CLK.t1 VDD.t34 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1005 GND a_6371_989.t8 a_9711_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1006 QN a_10219_989.t10 a_18760_101.t0 nshort w=-1.83u l=2.06u
+  ad=0.5373p pd=4.72u as=0p ps=0u
M1007 VDD.t111 SN.t0 a_15991_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1008 GND D.t4 a_5863_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1009 VDD.t68 SN.t1 a_10219_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1010 VDD.t36 a_12143_989.t7 a_15669_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_13745_1050.t6 a_11821_1050.t8 VDD.t103 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_6049_1050.t2 a_6371_989.t7 VDD.t20 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1013 VDD.t1 a_2201_1050.t7 a_1561_989.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1014 VDD.t71 a_7333_989.t7 a_7973_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1015 VDD.t50 a_10219_989.t8 a_9897_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_4447_989.t3 SN.t2 VDD.t8 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1017 QN.t6 a_4447_989.t8 a_18197_1051.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_17533_1051.t7 a_4447_989.t9 a_18197_1051.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1019 VDD.t23 CLK.t2 a_6371_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_7333_989.t6 RN.t0 VDD.t108 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1021 GND a_11821_1050.t9 a_12597_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1022 VDD.t16 D.t1 a_6049_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1023 GND a_13745_1050.t7 a_14521_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_7973_1050.t4 SN.t4 VDD.t90 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_18197_1051.t0 a_10219_989.t9 QN.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1026 VDD.t39 a_15991_989.t9 a_17533_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1027 GND a_9897_1050.t7 a_10673_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1028 GND a_7973_1050.t7 a_8749_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1029 VDD.t55 D.t2 a_277_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1030 VDD.t52 D.t3 a_11821_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1031 GND D.t5 a_91_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1032 VDD.t80 RN.t2 a_15669_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_599_989.t4 CLK.t3 VDD.t27 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1034 VDD.t107 RN.t3 a_9897_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_11821_1050.t1 a_12143_989.t8 VDD.t37 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1036 VDD.t30 CLK.t4 a_1561_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1037 VDD.t97 a_13105_989.t9 a_13745_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1038 GND a_15991_989.t11 a_17428_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1039 VDD.t15 a_277_1050.t7 a_2201_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_7333_989.t1 CLK.t6 VDD.t29 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_10219_989.t1 SN.t5 VDD.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1042 VDD.t4 a_7333_989.t8 a_6371_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1043 VDD.t25 CLK.t7 a_12143_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_13105_989.t1 RN.t4 VDD.t12 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1045 GND a_11821_1050.t10 a_13559_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1046 GND a_12143_989.t9 a_15483_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1047 QN a_4447_989.t11 a_18094_101.t0 nshort w=-1.235u l=1.535u
+  ad=0p pd=0u as=0p ps=0u
M1048 VDD.t75 RN.t5 a_277_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_6371_989.t4 a_6049_1050.t9 VDD.t58 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_17533_1051.t3 a_15991_989.t10 VDD.t40 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1051 VDD.t93 a_7973_1050.t8 a_7333_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1052 VDD.t91 a_9897_1050.t8 a_10219_989.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1053 a_12143_989.t0 CLK.t8 VDD.t24 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_599_989.t1 a_1561_989.t7 VDD.t67 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1055 a_15991_989.t2 a_15669_1050.t7 VDD.t45 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1056 VDD.t106 RN.t7 a_1561_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_9897_1050.t1 a_6371_989.t9 VDD.t73 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1058 GND a_15669_1050.t8 a_16445_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1059 a_4125_1050.t6 a_599_989.t8 VDD.t109 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1060 VDD.t83 SN.t6 a_2201_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1061 a_4125_1050.t5 a_4447_989.t10 VDD.t87 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1062 VDD.t53 a_6371_989.t10 a_6049_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1063 a_18197_1051.t3 a_15991_989.t12 a_17533_1051.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1064 a_1561_989.t1 CLK.t9 VDD.t32 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1065 VDD.t46 a_599_989.t9 a_277_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1066 a_13745_1050.t1 SN.t7 VDD.t70 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1067 a_17533_1051.t5 a_10219_989.t11 VDD.t47 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1068 a_12143_989.t2 a_11821_1050.t11 VDD.t13 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1069 VDD.t22 a_13745_1050.t8 a_13105_989.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1070 a_15991_989.t0 SN.t10 VDD.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1071 a_15669_1050.t1 a_12143_989.t10 VDD.t35 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1072 a_4125_1050.t2 RN.t9 VDD.t74 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1073 GND a_277_1050.t8 a_2015_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1074 VDD.t92 a_1561_989.t8 a_2201_1050.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1075 VDD.t79 RN.t10 a_6049_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1076 a_7333_989.t4 a_7973_1050.t9 VDD.t95 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1077 a_7973_1050.t1 a_7333_989.t9 VDD.t89 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1078 a_9897_1050.t2 a_10219_989.t12 VDD.t49 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1079 VDD.t101 a_13105_989.t10 a_15991_989.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1080 a_1561_989.t3 a_2201_1050.t8 VDD.t9 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1081 a_18197_1051.t4 a_4447_989.t13 a_17533_1051.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1082 VDD.t42 a_4125_1050.t8 a_4447_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1083 a_6371_989.t1 CLK.t12 VDD.t31 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1084 VDD.t28 CLK.t13 a_7333_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1085 a_6049_1050.t5 D.t6 VDD.t77 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1086 QN.t2 a_10219_989.t13 a_18197_1051.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1087 a_277_1050.t2 D.t7 VDD.t78 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1088 VDD.t33 CLK.t14 a_13105_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1089 a_15991_989.t4 a_13105_989.t11 VDD.t98 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1090 a_10219_989.t0 a_7333_989.t10 VDD.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1091 VDD.t14 a_11821_1050.t12 a_13745_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1092 QN a_10219_989.t14 a_17428_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1093 VDD.t100 a_13105_989.t12 a_12143_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1094 a_15669_1050.t0 RN.t13 VDD.t11 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1095 GND a_2201_1050.t9 a_2977_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1096 VDD.t63 a_277_1050.t9 a_599_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1097 a_9897_1050.t5 RN.t14 VDD.t51 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1098 VDD.t6 RN.t15 a_11821_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1099 VDD.t110 a_1561_989.t11 a_599_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1100 a_13745_1050.t5 a_13105_989.t13 VDD.t96 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1101 GND a_277_1050.t10 a_1053_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1102 VDD.t94 SN.t12 a_4447_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1103 a_18197_1051.t7 a_4447_989.t14 QN.t5 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1104 VDD.t17 a_15991_989.t13 a_15669_1050.t4 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1105 a_6371_989.t5 a_7333_989.t12 VDD.t66 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1106 VDD.t65 RN.t17 a_7333_989.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1107 VDD.t88 SN.t13 a_7973_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1108 a_277_1050.t0 RN.t18 VDD.t44 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1109 a_11821_1050.t3 RN.t19 VDD.t64 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1110 VDD.t85 SN.t14 a_13745_1050.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1111 a_10219_989.t4 a_9897_1050.t9 VDD.t84 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1112 GND a_599_989.t11 a_3939_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1113 VDD.t26 CLK.t15 a_599_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1114 a_1561_989.t5 RN.t20 VDD.t105 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1115 VDD.t82 a_12143_989.t12 a_11821_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1116 VDD.t86 a_1561_989.t13 a_4447_989.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1117 a_2201_1050.t2 SN.t15 VDD.t19 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1118 a_12143_989.t5 a_13105_989.t14 VDD.t99 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1119 VDD.t5 RN.t21 a_4125_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1120 VDD.t10 RN.t22 a_13105_989.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1121 a_599_989.t5 a_277_1050.t11 VDD.t57 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1122 VDD.t60 a_6049_1050.t10 a_7973_1050.t6 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1123 a_277_1050.t4 a_599_989.t10 VDD.t18 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1124 a_11821_1050.t4 D.t8 VDD.t76 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1125 GND a_6049_1050.t7 a_6825_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1126 a_13105_989.t6 a_13745_1050.t9 VDD.t21 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1127 GND a_4125_1050.t7 a_4901_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1128 VDD.t41 a_15669_1050.t9 a_15991_989.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1129 a_7973_1050.t5 a_6049_1050.t11 VDD.t61 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1130 VDD.t69 a_6371_989.t12 a_9897_1050.t0 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1131 a_2201_1050.t6 a_277_1050.t12 VDD.t104 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1132 VDD.t72 a_7333_989.t15 a_10219_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1133 a_2201_1050.t4 a_1561_989.t14 VDD.t54 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1134 VDD.t81 a_599_989.t12 a_4125_1050.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1135 a_6049_1050.t4 RN.t26 VDD.t62 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1136 GND a_4447_989.t7 a_18760_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1137 GND a_15991_989.t8 a_18094_101.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
M1138 VDD.t7 a_4447_989.t15 a_4125_1050.t1 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1139 a_17533_1051.t1 a_15991_989.t14 a_18197_1051.t2 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1140 a_4447_989.t0 a_4125_1050.t9 VDD.t38 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1141 VDD.t59 a_6049_1050.t12 a_6371_989.t3 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1142 a_4447_989.t4 a_1561_989.t15 VDD.t56 pshort w=2u l=0.15u
+  ad=0p pd=0u as=0p ps=0u
M1143 GND D.t0 a_11635_103.t0 nshort w=-1.605u l=1.765u
+  ad=0p pd=0u as=0p ps=0u
C0 VDD RN 0.48fF
C1 VDD CLK 1.65fF
C2 D RN 2.36fF
C3 VDD SN 0.30fF
C4 D CLK 12.06fF
C5 VDD QN 0.29fF
C6 RN CLK 1.11fF
C7 D SN 0.31fF
C8 RN SN 16.07fF
C9 CLK SN 0.63fF
C10 VDD D 5.87fF
R0 CLK.n18 CLK.t15 459.505
R1 CLK.n15 CLK.t4 459.505
R2 CLK.n12 CLK.t2 459.505
R3 CLK.n7 CLK.t13 459.505
R4 CLK.n4 CLK.t7 459.505
R5 CLK.n0 CLK.t14 459.505
R6 CLK.n18 CLK.t3 384.527
R7 CLK.n15 CLK.t9 384.527
R8 CLK.n12 CLK.t12 384.527
R9 CLK.n7 CLK.t6 384.527
R10 CLK.n4 CLK.t8 384.527
R11 CLK.n0 CLK.t1 384.527
R12 CLK.n16 CLK.t0 322.151
R13 CLK.n8 CLK.t5 322.151
R14 CLK.n1 CLK.t10 322.151
R15 CLK.n20 CLK.t17 321.792
R16 CLK.n10 CLK.t16 320.152
R17 CLK.n2 CLK.t11 320.152
R18 CLK.n19 CLK 152
R19 CLK.n6 CLK.n5 75.989
R20 CLK.n14 CLK.n13 75.989
R21 CLK.n3 CLK.n2 75.568
R22 CLK.n11 CLK.n10 75.568
R23 CLK.n3 CLK.n1 56.374
R24 CLK.n21 CLK.n20 49.379
R25 CLK.n9 CLK.n8 49.342
R26 CLK.n17 CLK.n16 49.342
R27 CLK.n1 CLK.n0 27.599
R28 CLK.n8 CLK.n7 27.599
R29 CLK.n16 CLK.n15 27.599
R30 CLK.n19 CLK.n18 21.475
R31 CLK.n13 CLK.n12 21.475
R32 CLK.n5 CLK.n4 21.475
R33 CLK.n9 CLK.n6 14.076
R34 CLK.n17 CLK.n14 14.076
R35 CLK.n11 CLK.n9 7.032
R36 CLK.n21 CLK.n17 7.032
R37 CLK.n20 CLK.n19 3.3
R38 CLK.n21 CLK 0.046
R39 CLK.n6 CLK.n3 0.023
R40 CLK.n14 CLK.n11 0.023
R41 a_2977_103.t0 a_2977_103.n0 117.777
R42 a_2977_103.n2 a_2977_103.n1 55.228
R43 a_2977_103.n4 a_2977_103.n3 9.111
R44 a_2977_103.n8 a_2977_103.n6 7.859
R45 a_2977_103.t0 a_2977_103.n2 4.04
R46 a_2977_103.t0 a_2977_103.n8 3.034
R47 a_2977_103.n6 a_2977_103.n4 1.964
R48 a_2977_103.n6 a_2977_103.n5 1.964
R49 a_2977_103.n8 a_2977_103.n7 0.443
R50 a_3258_210.n12 a_3258_210.n5 96.467
R51 a_3258_210.t0 a_3258_210.n1 46.91
R52 a_3258_210.n9 a_3258_210.n7 34.805
R53 a_3258_210.n9 a_3258_210.n8 32.622
R54 a_3258_210.t0 a_3258_210.n12 32.417
R55 a_3258_210.n5 a_3258_210.n4 22.349
R56 a_3258_210.n11 a_3258_210.n9 19.017
R57 a_3258_210.n1 a_3258_210.n0 17.006
R58 a_3258_210.n5 a_3258_210.n3 8.443
R59 a_3258_210.t0 a_3258_210.n2 8.137
R60 a_3258_210.n7 a_3258_210.n6 7.5
R61 a_3258_210.n11 a_3258_210.n10 7.5
R62 a_3258_210.n12 a_3258_210.n11 1.435
R63 a_13105_989.n7 a_13105_989.t13 454.685
R64 a_13105_989.n9 a_13105_989.t14 454.685
R65 a_13105_989.n5 a_13105_989.t11 454.685
R66 a_13105_989.n7 a_13105_989.t9 428.979
R67 a_13105_989.n9 a_13105_989.t12 428.979
R68 a_13105_989.n5 a_13105_989.t10 428.979
R69 a_13105_989.n8 a_13105_989.t7 264.512
R70 a_13105_989.n6 a_13105_989.t8 264.512
R71 a_13105_989.n10 a_13105_989.t15 264.173
R72 a_13105_989.n15 a_13105_989.n13 246.179
R73 a_13105_989.n13 a_13105_989.n4 144.246
R74 a_13105_989.n12 a_13105_989.n6 82.484
R75 a_13105_989.n11 a_13105_989.n10 79.495
R76 a_13105_989.n3 a_13105_989.n2 79.232
R77 a_13105_989.n11 a_13105_989.n8 76
R78 a_13105_989.n13 a_13105_989.n12 76
R79 a_13105_989.n8 a_13105_989.n7 71.894
R80 a_13105_989.n6 a_13105_989.n5 71.894
R81 a_13105_989.n10 a_13105_989.n9 71.555
R82 a_13105_989.n4 a_13105_989.n3 63.152
R83 a_13105_989.n4 a_13105_989.n0 16.08
R84 a_13105_989.n3 a_13105_989.n1 16.08
R85 a_13105_989.n15 a_13105_989.n14 15.218
R86 a_13105_989.n0 a_13105_989.t0 14.282
R87 a_13105_989.n0 a_13105_989.t1 14.282
R88 a_13105_989.n1 a_13105_989.t3 14.282
R89 a_13105_989.n1 a_13105_989.t2 14.282
R90 a_13105_989.n2 a_13105_989.t5 14.282
R91 a_13105_989.n2 a_13105_989.t6 14.282
R92 a_13105_989.n16 a_13105_989.n15 12.014
R93 a_13105_989.n12 a_13105_989.n11 4.035
R94 a_13840_210.n12 a_13840_210.n5 96.467
R95 a_13840_210.t0 a_13840_210.n1 46.91
R96 a_13840_210.n9 a_13840_210.n7 34.805
R97 a_13840_210.n9 a_13840_210.n8 32.622
R98 a_13840_210.t0 a_13840_210.n12 32.417
R99 a_13840_210.n5 a_13840_210.n4 22.349
R100 a_13840_210.n11 a_13840_210.n9 19.017
R101 a_13840_210.n1 a_13840_210.n0 17.006
R102 a_13840_210.n5 a_13840_210.n3 8.443
R103 a_13840_210.t0 a_13840_210.n2 8.137
R104 a_13840_210.n7 a_13840_210.n6 7.5
R105 a_13840_210.n11 a_13840_210.n10 7.5
R106 a_13840_210.n12 a_13840_210.n11 1.435
R107 a_13745_1050.n5 a_13745_1050.t8 512.525
R108 a_13745_1050.n5 a_13745_1050.t9 371.139
R109 a_13745_1050.n6 a_13745_1050.t7 234.562
R110 a_13745_1050.n7 a_13745_1050.n4 223.905
R111 a_13745_1050.n6 a_13745_1050.n5 215.819
R112 a_13745_1050.n9 a_13745_1050.n7 166.52
R113 a_13745_1050.n7 a_13745_1050.n6 153.315
R114 a_13745_1050.n3 a_13745_1050.n2 79.232
R115 a_13745_1050.n4 a_13745_1050.n3 63.152
R116 a_13745_1050.n4 a_13745_1050.n0 16.08
R117 a_13745_1050.n3 a_13745_1050.n1 16.08
R118 a_13745_1050.n9 a_13745_1050.n8 15.218
R119 a_13745_1050.n0 a_13745_1050.t4 14.282
R120 a_13745_1050.n0 a_13745_1050.t5 14.282
R121 a_13745_1050.n1 a_13745_1050.t2 14.282
R122 a_13745_1050.n1 a_13745_1050.t1 14.282
R123 a_13745_1050.n2 a_13745_1050.t0 14.282
R124 a_13745_1050.n2 a_13745_1050.t6 14.282
R125 a_13745_1050.n10 a_13745_1050.n9 12.014
R126 a_6049_1050.n7 a_6049_1050.t12 512.525
R127 a_6049_1050.n5 a_6049_1050.t10 512.525
R128 a_6049_1050.n7 a_6049_1050.t9 371.139
R129 a_6049_1050.n5 a_6049_1050.t11 371.139
R130 a_6049_1050.n8 a_6049_1050.t7 234.921
R131 a_6049_1050.n6 a_6049_1050.t8 234.921
R132 a_6049_1050.n10 a_6049_1050.n4 223.546
R133 a_6049_1050.n8 a_6049_1050.n7 215.46
R134 a_6049_1050.n6 a_6049_1050.n5 215.46
R135 a_6049_1050.n12 a_6049_1050.n10 166.879
R136 a_6049_1050.n9 a_6049_1050.n6 79.491
R137 a_6049_1050.n3 a_6049_1050.n2 79.232
R138 a_6049_1050.n10 a_6049_1050.n9 77.315
R139 a_6049_1050.n9 a_6049_1050.n8 76
R140 a_6049_1050.n4 a_6049_1050.n3 63.152
R141 a_6049_1050.n4 a_6049_1050.n0 16.08
R142 a_6049_1050.n3 a_6049_1050.n1 16.08
R143 a_6049_1050.n12 a_6049_1050.n11 15.218
R144 a_6049_1050.n0 a_6049_1050.t3 14.282
R145 a_6049_1050.n0 a_6049_1050.t2 14.282
R146 a_6049_1050.n1 a_6049_1050.t6 14.282
R147 a_6049_1050.n1 a_6049_1050.t4 14.282
R148 a_6049_1050.n2 a_6049_1050.t1 14.282
R149 a_6049_1050.n2 a_6049_1050.t5 14.282
R150 a_6049_1050.n13 a_6049_1050.n12 12.014
R151 a_6825_103.t0 a_6825_103.n0 117.777
R152 a_6825_103.n2 a_6825_103.n1 55.228
R153 a_6825_103.n4 a_6825_103.n3 9.111
R154 a_6825_103.n8 a_6825_103.n6 7.859
R155 a_6825_103.t0 a_6825_103.n2 4.04
R156 a_6825_103.t0 a_6825_103.n8 3.034
R157 a_6825_103.n6 a_6825_103.n4 1.964
R158 a_6825_103.n6 a_6825_103.n5 1.964
R159 a_6825_103.n8 a_6825_103.n7 0.443
R160 GND.n26 GND.n24 219.745
R161 GND.n56 GND.n54 219.745
R162 GND.n468 GND.n467 219.745
R163 GND.n510 GND.n508 219.745
R164 GND.n552 GND.n550 219.745
R165 GND.n594 GND.n592 219.745
R166 GND.n636 GND.n634 219.745
R167 GND.n678 GND.n676 219.745
R168 GND.n723 GND.n721 219.745
R169 GND.n765 GND.n763 219.745
R170 GND.n810 GND.n808 219.745
R171 GND.n423 GND.n421 219.745
R172 GND.n383 GND.n381 219.745
R173 GND.n341 GND.n339 219.745
R174 GND.n299 GND.n297 219.745
R175 GND.n257 GND.n255 219.745
R176 GND.n215 GND.n213 219.745
R177 GND.n170 GND.n168 219.745
R178 GND.n128 GND.n126 219.745
R179 GND.n86 GND.n85 219.745
R180 GND.n117 GND.n116 85.559
R181 GND.n159 GND.n158 85.559
R182 GND.n246 GND.n245 85.559
R183 GND.n288 GND.n287 85.559
R184 GND.n330 GND.n329 85.559
R185 GND.n372 GND.n371 85.559
R186 GND.n414 GND.n413 85.559
R187 GND.n819 GND.n818 85.559
R188 GND.n732 GND.n731 85.559
R189 GND.n645 GND.n644 85.559
R190 GND.n603 GND.n602 85.559
R191 GND.n561 GND.n560 85.559
R192 GND.n519 GND.n518 85.559
R193 GND.n477 GND.n476 85.559
R194 GND.n435 GND.n434 85.559
R195 GND.n26 GND.n25 85.529
R196 GND.n56 GND.n55 85.529
R197 GND.n468 GND.n466 85.529
R198 GND.n510 GND.n509 85.529
R199 GND.n552 GND.n551 85.529
R200 GND.n594 GND.n593 85.529
R201 GND.n636 GND.n635 85.529
R202 GND.n678 GND.n677 85.529
R203 GND.n723 GND.n722 85.529
R204 GND.n765 GND.n764 85.529
R205 GND.n810 GND.n809 85.529
R206 GND.n423 GND.n422 85.529
R207 GND.n383 GND.n382 85.529
R208 GND.n341 GND.n340 85.529
R209 GND.n299 GND.n298 85.529
R210 GND.n257 GND.n256 85.529
R211 GND.n215 GND.n214 85.529
R212 GND.n170 GND.n169 85.529
R213 GND.n128 GND.n127 85.529
R214 GND.n86 GND.n84 85.529
R215 GND.n44 GND.n43 84.842
R216 GND.n74 GND.n73 84.842
R217 GND.n14 GND.n13 84.842
R218 GND.n429 GND.n428 76
R219 GND.n39 GND.n38 76
R220 GND.n42 GND.n41 76
R221 GND.n47 GND.n46 76
R222 GND.n50 GND.n49 76
R223 GND.n53 GND.n52 76
R224 GND.n60 GND.n59 76
R225 GND.n63 GND.n62 76
R226 GND.n66 GND.n65 76
R227 GND.n69 GND.n68 76
R228 GND.n72 GND.n71 76
R229 GND.n77 GND.n76 76
R230 GND.n80 GND.n79 76
R231 GND.n83 GND.n82 76
R232 GND.n90 GND.n89 76
R233 GND.n93 GND.n92 76
R234 GND.n96 GND.n95 76
R235 GND.n99 GND.n98 76
R236 GND.n102 GND.n101 76
R237 GND.n105 GND.n104 76
R238 GND.n108 GND.n107 76
R239 GND.n111 GND.n110 76
R240 GND.n114 GND.n113 76
R241 GND.n119 GND.n118 76
R242 GND.n122 GND.n121 76
R243 GND.n125 GND.n124 76
R244 GND.n132 GND.n131 76
R245 GND.n135 GND.n134 76
R246 GND.n138 GND.n137 76
R247 GND.n141 GND.n140 76
R248 GND.n144 GND.n143 76
R249 GND.n147 GND.n146 76
R250 GND.n150 GND.n149 76
R251 GND.n153 GND.n152 76
R252 GND.n156 GND.n155 76
R253 GND.n161 GND.n160 76
R254 GND.n164 GND.n163 76
R255 GND.n167 GND.n166 76
R256 GND.n174 GND.n173 76
R257 GND.n177 GND.n176 76
R258 GND.n180 GND.n179 76
R259 GND.n183 GND.n182 76
R260 GND.n186 GND.n185 76
R261 GND.n189 GND.n188 76
R262 GND.n192 GND.n191 76
R263 GND.n195 GND.n194 76
R264 GND.n198 GND.n197 76
R265 GND.n206 GND.n205 76
R266 GND.n209 GND.n208 76
R267 GND.n212 GND.n211 76
R268 GND.n219 GND.n218 76
R269 GND.n222 GND.n221 76
R270 GND.n225 GND.n224 76
R271 GND.n228 GND.n227 76
R272 GND.n231 GND.n230 76
R273 GND.n234 GND.n233 76
R274 GND.n237 GND.n236 76
R275 GND.n240 GND.n239 76
R276 GND.n243 GND.n242 76
R277 GND.n248 GND.n247 76
R278 GND.n251 GND.n250 76
R279 GND.n254 GND.n253 76
R280 GND.n261 GND.n260 76
R281 GND.n264 GND.n263 76
R282 GND.n267 GND.n266 76
R283 GND.n270 GND.n269 76
R284 GND.n273 GND.n272 76
R285 GND.n276 GND.n275 76
R286 GND.n279 GND.n278 76
R287 GND.n282 GND.n281 76
R288 GND.n285 GND.n284 76
R289 GND.n290 GND.n289 76
R290 GND.n293 GND.n292 76
R291 GND.n296 GND.n295 76
R292 GND.n303 GND.n302 76
R293 GND.n306 GND.n305 76
R294 GND.n309 GND.n308 76
R295 GND.n312 GND.n311 76
R296 GND.n315 GND.n314 76
R297 GND.n318 GND.n317 76
R298 GND.n321 GND.n320 76
R299 GND.n324 GND.n323 76
R300 GND.n327 GND.n326 76
R301 GND.n332 GND.n331 76
R302 GND.n335 GND.n334 76
R303 GND.n338 GND.n337 76
R304 GND.n345 GND.n344 76
R305 GND.n348 GND.n347 76
R306 GND.n351 GND.n350 76
R307 GND.n354 GND.n353 76
R308 GND.n357 GND.n356 76
R309 GND.n360 GND.n359 76
R310 GND.n363 GND.n362 76
R311 GND.n366 GND.n365 76
R312 GND.n369 GND.n368 76
R313 GND.n374 GND.n373 76
R314 GND.n377 GND.n376 76
R315 GND.n380 GND.n379 76
R316 GND.n387 GND.n386 76
R317 GND.n390 GND.n389 76
R318 GND.n393 GND.n392 76
R319 GND.n396 GND.n395 76
R320 GND.n399 GND.n398 76
R321 GND.n402 GND.n401 76
R322 GND.n405 GND.n404 76
R323 GND.n408 GND.n407 76
R324 GND.n411 GND.n410 76
R325 GND.n416 GND.n415 76
R326 GND.n419 GND.n418 76
R327 GND.n426 GND.n425 76
R328 GND.n848 GND.n847 76
R329 GND.n845 GND.n844 76
R330 GND.n842 GND.n841 76
R331 GND.n839 GND.n838 76
R332 GND.n836 GND.n835 76
R333 GND.n833 GND.n832 76
R334 GND.n830 GND.n829 76
R335 GND.n827 GND.n826 76
R336 GND.n824 GND.n823 76
R337 GND.n821 GND.n820 76
R338 GND.n816 GND.n815 76
R339 GND.n813 GND.n812 76
R340 GND.n806 GND.n805 76
R341 GND.n803 GND.n802 76
R342 GND.n800 GND.n799 76
R343 GND.n797 GND.n796 76
R344 GND.n794 GND.n793 76
R345 GND.n791 GND.n790 76
R346 GND.n788 GND.n787 76
R347 GND.n785 GND.n784 76
R348 GND.n782 GND.n781 76
R349 GND.n779 GND.n778 76
R350 GND.n771 GND.n770 76
R351 GND.n768 GND.n767 76
R352 GND.n761 GND.n760 76
R353 GND.n758 GND.n757 76
R354 GND.n755 GND.n754 76
R355 GND.n752 GND.n751 76
R356 GND.n749 GND.n748 76
R357 GND.n746 GND.n745 76
R358 GND.n743 GND.n742 76
R359 GND.n740 GND.n739 76
R360 GND.n737 GND.n736 76
R361 GND.n734 GND.n733 76
R362 GND.n729 GND.n728 76
R363 GND.n726 GND.n725 76
R364 GND.n719 GND.n718 76
R365 GND.n716 GND.n715 76
R366 GND.n713 GND.n712 76
R367 GND.n710 GND.n709 76
R368 GND.n707 GND.n706 76
R369 GND.n704 GND.n703 76
R370 GND.n701 GND.n700 76
R371 GND.n698 GND.n697 76
R372 GND.n695 GND.n694 76
R373 GND.n692 GND.n691 76
R374 GND.n684 GND.n683 76
R375 GND.n681 GND.n680 76
R376 GND.n674 GND.n673 76
R377 GND.n671 GND.n670 76
R378 GND.n668 GND.n667 76
R379 GND.n665 GND.n664 76
R380 GND.n662 GND.n661 76
R381 GND.n659 GND.n658 76
R382 GND.n656 GND.n655 76
R383 GND.n653 GND.n652 76
R384 GND.n650 GND.n649 76
R385 GND.n647 GND.n646 76
R386 GND.n642 GND.n641 76
R387 GND.n639 GND.n638 76
R388 GND.n632 GND.n631 76
R389 GND.n629 GND.n628 76
R390 GND.n626 GND.n625 76
R391 GND.n623 GND.n622 76
R392 GND.n620 GND.n619 76
R393 GND.n617 GND.n616 76
R394 GND.n614 GND.n613 76
R395 GND.n611 GND.n610 76
R396 GND.n608 GND.n607 76
R397 GND.n605 GND.n604 76
R398 GND.n600 GND.n599 76
R399 GND.n597 GND.n596 76
R400 GND.n590 GND.n589 76
R401 GND.n587 GND.n586 76
R402 GND.n584 GND.n583 76
R403 GND.n581 GND.n580 76
R404 GND.n578 GND.n577 76
R405 GND.n575 GND.n574 76
R406 GND.n572 GND.n571 76
R407 GND.n569 GND.n568 76
R408 GND.n566 GND.n565 76
R409 GND.n563 GND.n562 76
R410 GND.n558 GND.n557 76
R411 GND.n555 GND.n554 76
R412 GND.n548 GND.n547 76
R413 GND.n545 GND.n544 76
R414 GND.n542 GND.n541 76
R415 GND.n539 GND.n538 76
R416 GND.n536 GND.n535 76
R417 GND.n533 GND.n532 76
R418 GND.n530 GND.n529 76
R419 GND.n527 GND.n526 76
R420 GND.n524 GND.n523 76
R421 GND.n521 GND.n520 76
R422 GND.n516 GND.n515 76
R423 GND.n513 GND.n512 76
R424 GND.n506 GND.n505 76
R425 GND.n503 GND.n502 76
R426 GND.n500 GND.n499 76
R427 GND.n497 GND.n496 76
R428 GND.n494 GND.n493 76
R429 GND.n491 GND.n490 76
R430 GND.n488 GND.n487 76
R431 GND.n485 GND.n484 76
R432 GND.n482 GND.n481 76
R433 GND.n479 GND.n478 76
R434 GND.n474 GND.n473 76
R435 GND.n471 GND.n470 76
R436 GND.n464 GND.n463 76
R437 GND.n461 GND.n460 76
R438 GND.n458 GND.n457 76
R439 GND.n455 GND.n454 76
R440 GND.n452 GND.n451 76
R441 GND.n449 GND.n448 76
R442 GND.n446 GND.n445 76
R443 GND.n443 GND.n442 76
R444 GND.n440 GND.n439 76
R445 GND.n437 GND.n436 76
R446 GND.n432 GND.n431 76
R447 GND.n12 GND.n11 76
R448 GND.n17 GND.n16 76
R449 GND.n20 GND.n19 76
R450 GND.n23 GND.n22 76
R451 GND.n30 GND.n29 76
R452 GND.n33 GND.n32 76
R453 GND.n36 GND.n35 76
R454 GND.n204 GND.n203 64.552
R455 GND.n777 GND.n776 64.552
R456 GND.n690 GND.n689 64.552
R457 GND.n8 GND.n7 34.942
R458 GND.n203 GND.n202 28.421
R459 GND.n776 GND.n775 28.421
R460 GND.n689 GND.n688 28.421
R461 GND.n203 GND.n201 25.263
R462 GND.n776 GND.n774 25.263
R463 GND.n689 GND.n687 25.263
R464 GND.n201 GND.n200 24.383
R465 GND.n774 GND.n773 24.383
R466 GND.n687 GND.n686 24.383
R467 GND.n5 GND.n4 14.167
R468 GND.n4 GND.n2 14.167
R469 GND.n29 GND.n27 14.167
R470 GND.n59 GND.n57 14.167
R471 GND.n89 GND.n87 14.167
R472 GND.n131 GND.n129 14.167
R473 GND.n173 GND.n171 14.167
R474 GND.n218 GND.n216 14.167
R475 GND.n260 GND.n258 14.167
R476 GND.n302 GND.n300 14.167
R477 GND.n344 GND.n342 14.167
R478 GND.n386 GND.n384 14.167
R479 GND.n425 GND.n424 14.167
R480 GND.n812 GND.n811 14.167
R481 GND.n767 GND.n766 14.167
R482 GND.n725 GND.n724 14.167
R483 GND.n680 GND.n679 14.167
R484 GND.n638 GND.n637 14.167
R485 GND.n596 GND.n595 14.167
R486 GND.n554 GND.n553 14.167
R487 GND.n512 GND.n511 14.167
R488 GND.n470 GND.n469 14.167
R489 GND.n431 GND.n430 13.653
R490 GND.n436 GND.n433 13.653
R491 GND.n439 GND.n438 13.653
R492 GND.n442 GND.n441 13.653
R493 GND.n445 GND.n444 13.653
R494 GND.n448 GND.n447 13.653
R495 GND.n451 GND.n450 13.653
R496 GND.n454 GND.n453 13.653
R497 GND.n457 GND.n456 13.653
R498 GND.n460 GND.n459 13.653
R499 GND.n463 GND.n462 13.653
R500 GND.n470 GND.n465 13.653
R501 GND.n473 GND.n472 13.653
R502 GND.n478 GND.n475 13.653
R503 GND.n481 GND.n480 13.653
R504 GND.n484 GND.n483 13.653
R505 GND.n487 GND.n486 13.653
R506 GND.n490 GND.n489 13.653
R507 GND.n493 GND.n492 13.653
R508 GND.n496 GND.n495 13.653
R509 GND.n499 GND.n498 13.653
R510 GND.n502 GND.n501 13.653
R511 GND.n505 GND.n504 13.653
R512 GND.n512 GND.n507 13.653
R513 GND.n515 GND.n514 13.653
R514 GND.n520 GND.n517 13.653
R515 GND.n523 GND.n522 13.653
R516 GND.n526 GND.n525 13.653
R517 GND.n529 GND.n528 13.653
R518 GND.n532 GND.n531 13.653
R519 GND.n535 GND.n534 13.653
R520 GND.n538 GND.n537 13.653
R521 GND.n541 GND.n540 13.653
R522 GND.n544 GND.n543 13.653
R523 GND.n547 GND.n546 13.653
R524 GND.n554 GND.n549 13.653
R525 GND.n557 GND.n556 13.653
R526 GND.n562 GND.n559 13.653
R527 GND.n565 GND.n564 13.653
R528 GND.n568 GND.n567 13.653
R529 GND.n571 GND.n570 13.653
R530 GND.n574 GND.n573 13.653
R531 GND.n577 GND.n576 13.653
R532 GND.n580 GND.n579 13.653
R533 GND.n583 GND.n582 13.653
R534 GND.n586 GND.n585 13.653
R535 GND.n589 GND.n588 13.653
R536 GND.n596 GND.n591 13.653
R537 GND.n599 GND.n598 13.653
R538 GND.n604 GND.n601 13.653
R539 GND.n607 GND.n606 13.653
R540 GND.n610 GND.n609 13.653
R541 GND.n613 GND.n612 13.653
R542 GND.n616 GND.n615 13.653
R543 GND.n619 GND.n618 13.653
R544 GND.n622 GND.n621 13.653
R545 GND.n625 GND.n624 13.653
R546 GND.n628 GND.n627 13.653
R547 GND.n631 GND.n630 13.653
R548 GND.n638 GND.n633 13.653
R549 GND.n641 GND.n640 13.653
R550 GND.n646 GND.n643 13.653
R551 GND.n649 GND.n648 13.653
R552 GND.n652 GND.n651 13.653
R553 GND.n655 GND.n654 13.653
R554 GND.n658 GND.n657 13.653
R555 GND.n661 GND.n660 13.653
R556 GND.n664 GND.n663 13.653
R557 GND.n667 GND.n666 13.653
R558 GND.n670 GND.n669 13.653
R559 GND.n673 GND.n672 13.653
R560 GND.n680 GND.n675 13.653
R561 GND.n683 GND.n682 13.653
R562 GND.n691 GND.n685 13.653
R563 GND.n694 GND.n693 13.653
R564 GND.n697 GND.n696 13.653
R565 GND.n700 GND.n699 13.653
R566 GND.n703 GND.n702 13.653
R567 GND.n706 GND.n705 13.653
R568 GND.n709 GND.n708 13.653
R569 GND.n712 GND.n711 13.653
R570 GND.n715 GND.n714 13.653
R571 GND.n718 GND.n717 13.653
R572 GND.n725 GND.n720 13.653
R573 GND.n728 GND.n727 13.653
R574 GND.n733 GND.n730 13.653
R575 GND.n736 GND.n735 13.653
R576 GND.n739 GND.n738 13.653
R577 GND.n742 GND.n741 13.653
R578 GND.n745 GND.n744 13.653
R579 GND.n748 GND.n747 13.653
R580 GND.n751 GND.n750 13.653
R581 GND.n754 GND.n753 13.653
R582 GND.n757 GND.n756 13.653
R583 GND.n760 GND.n759 13.653
R584 GND.n767 GND.n762 13.653
R585 GND.n770 GND.n769 13.653
R586 GND.n778 GND.n772 13.653
R587 GND.n781 GND.n780 13.653
R588 GND.n784 GND.n783 13.653
R589 GND.n787 GND.n786 13.653
R590 GND.n790 GND.n789 13.653
R591 GND.n793 GND.n792 13.653
R592 GND.n796 GND.n795 13.653
R593 GND.n799 GND.n798 13.653
R594 GND.n802 GND.n801 13.653
R595 GND.n805 GND.n804 13.653
R596 GND.n812 GND.n807 13.653
R597 GND.n815 GND.n814 13.653
R598 GND.n820 GND.n817 13.653
R599 GND.n823 GND.n822 13.653
R600 GND.n826 GND.n825 13.653
R601 GND.n829 GND.n828 13.653
R602 GND.n832 GND.n831 13.653
R603 GND.n835 GND.n834 13.653
R604 GND.n838 GND.n837 13.653
R605 GND.n841 GND.n840 13.653
R606 GND.n844 GND.n843 13.653
R607 GND.n847 GND.n846 13.653
R608 GND.n425 GND.n420 13.653
R609 GND.n418 GND.n417 13.653
R610 GND.n415 GND.n412 13.653
R611 GND.n410 GND.n409 13.653
R612 GND.n407 GND.n406 13.653
R613 GND.n404 GND.n403 13.653
R614 GND.n401 GND.n400 13.653
R615 GND.n398 GND.n397 13.653
R616 GND.n395 GND.n394 13.653
R617 GND.n392 GND.n391 13.653
R618 GND.n389 GND.n388 13.653
R619 GND.n386 GND.n385 13.653
R620 GND.n379 GND.n378 13.653
R621 GND.n376 GND.n375 13.653
R622 GND.n373 GND.n370 13.653
R623 GND.n368 GND.n367 13.653
R624 GND.n365 GND.n364 13.653
R625 GND.n362 GND.n361 13.653
R626 GND.n359 GND.n358 13.653
R627 GND.n356 GND.n355 13.653
R628 GND.n353 GND.n352 13.653
R629 GND.n350 GND.n349 13.653
R630 GND.n347 GND.n346 13.653
R631 GND.n344 GND.n343 13.653
R632 GND.n337 GND.n336 13.653
R633 GND.n334 GND.n333 13.653
R634 GND.n331 GND.n328 13.653
R635 GND.n326 GND.n325 13.653
R636 GND.n323 GND.n322 13.653
R637 GND.n320 GND.n319 13.653
R638 GND.n317 GND.n316 13.653
R639 GND.n314 GND.n313 13.653
R640 GND.n311 GND.n310 13.653
R641 GND.n308 GND.n307 13.653
R642 GND.n305 GND.n304 13.653
R643 GND.n302 GND.n301 13.653
R644 GND.n295 GND.n294 13.653
R645 GND.n292 GND.n291 13.653
R646 GND.n289 GND.n286 13.653
R647 GND.n284 GND.n283 13.653
R648 GND.n281 GND.n280 13.653
R649 GND.n278 GND.n277 13.653
R650 GND.n275 GND.n274 13.653
R651 GND.n272 GND.n271 13.653
R652 GND.n269 GND.n268 13.653
R653 GND.n266 GND.n265 13.653
R654 GND.n263 GND.n262 13.653
R655 GND.n260 GND.n259 13.653
R656 GND.n253 GND.n252 13.653
R657 GND.n250 GND.n249 13.653
R658 GND.n247 GND.n244 13.653
R659 GND.n242 GND.n241 13.653
R660 GND.n239 GND.n238 13.653
R661 GND.n236 GND.n235 13.653
R662 GND.n233 GND.n232 13.653
R663 GND.n230 GND.n229 13.653
R664 GND.n227 GND.n226 13.653
R665 GND.n224 GND.n223 13.653
R666 GND.n221 GND.n220 13.653
R667 GND.n218 GND.n217 13.653
R668 GND.n211 GND.n210 13.653
R669 GND.n208 GND.n207 13.653
R670 GND.n205 GND.n199 13.653
R671 GND.n197 GND.n196 13.653
R672 GND.n194 GND.n193 13.653
R673 GND.n191 GND.n190 13.653
R674 GND.n188 GND.n187 13.653
R675 GND.n185 GND.n184 13.653
R676 GND.n182 GND.n181 13.653
R677 GND.n179 GND.n178 13.653
R678 GND.n176 GND.n175 13.653
R679 GND.n173 GND.n172 13.653
R680 GND.n166 GND.n165 13.653
R681 GND.n163 GND.n162 13.653
R682 GND.n160 GND.n157 13.653
R683 GND.n155 GND.n154 13.653
R684 GND.n152 GND.n151 13.653
R685 GND.n149 GND.n148 13.653
R686 GND.n146 GND.n145 13.653
R687 GND.n143 GND.n142 13.653
R688 GND.n140 GND.n139 13.653
R689 GND.n137 GND.n136 13.653
R690 GND.n134 GND.n133 13.653
R691 GND.n131 GND.n130 13.653
R692 GND.n124 GND.n123 13.653
R693 GND.n121 GND.n120 13.653
R694 GND.n118 GND.n115 13.653
R695 GND.n113 GND.n112 13.653
R696 GND.n110 GND.n109 13.653
R697 GND.n107 GND.n106 13.653
R698 GND.n104 GND.n103 13.653
R699 GND.n101 GND.n100 13.653
R700 GND.n98 GND.n97 13.653
R701 GND.n95 GND.n94 13.653
R702 GND.n92 GND.n91 13.653
R703 GND.n89 GND.n88 13.653
R704 GND.n82 GND.n81 13.653
R705 GND.n79 GND.n78 13.653
R706 GND.n76 GND.n75 13.653
R707 GND.n71 GND.n70 13.653
R708 GND.n68 GND.n67 13.653
R709 GND.n65 GND.n64 13.653
R710 GND.n62 GND.n61 13.653
R711 GND.n59 GND.n58 13.653
R712 GND.n52 GND.n51 13.653
R713 GND.n49 GND.n48 13.653
R714 GND.n46 GND.n45 13.653
R715 GND.n41 GND.n40 13.653
R716 GND.n38 GND.n37 13.653
R717 GND.n5 GND.n0 13.653
R718 GND.n4 GND.n3 13.653
R719 GND.n2 GND.n1 13.653
R720 GND.n11 GND.n10 13.653
R721 GND.n16 GND.n15 13.653
R722 GND.n19 GND.n18 13.653
R723 GND.n22 GND.n21 13.653
R724 GND.n29 GND.n28 13.653
R725 GND.n32 GND.n31 13.653
R726 GND.n35 GND.n34 13.653
R727 GND.n27 GND.n26 7.312
R728 GND.n57 GND.n56 7.312
R729 GND.n469 GND.n468 7.312
R730 GND.n511 GND.n510 7.312
R731 GND.n553 GND.n552 7.312
R732 GND.n595 GND.n594 7.312
R733 GND.n637 GND.n636 7.312
R734 GND.n679 GND.n678 7.312
R735 GND.n724 GND.n723 7.312
R736 GND.n766 GND.n765 7.312
R737 GND.n811 GND.n810 7.312
R738 GND.n424 GND.n423 7.312
R739 GND.n384 GND.n383 7.312
R740 GND.n342 GND.n341 7.312
R741 GND.n300 GND.n299 7.312
R742 GND.n258 GND.n257 7.312
R743 GND.n216 GND.n215 7.312
R744 GND.n171 GND.n170 7.312
R745 GND.n129 GND.n128 7.312
R746 GND.n87 GND.n86 7.312
R747 GND.n7 GND.n6 7.084
R748 GND.n7 GND.n5 6.475
R749 GND.n16 GND.n14 3.935
R750 GND.n46 GND.n44 3.935
R751 GND.n76 GND.n74 3.935
R752 GND.n428 GND.n427 0.596
R753 GND.n30 GND.n23 0.29
R754 GND.n60 GND.n53 0.29
R755 GND.n90 GND.n83 0.29
R756 GND.n132 GND.n125 0.29
R757 GND.n174 GND.n167 0.29
R758 GND.n219 GND.n212 0.29
R759 GND.n261 GND.n254 0.29
R760 GND.n303 GND.n296 0.29
R761 GND.n345 GND.n338 0.29
R762 GND.n387 GND.n380 0.29
R763 GND.n813 GND.n806 0.29
R764 GND.n768 GND.n761 0.29
R765 GND.n726 GND.n719 0.29
R766 GND.n681 GND.n674 0.29
R767 GND.n639 GND.n632 0.29
R768 GND.n597 GND.n590 0.29
R769 GND.n555 GND.n548 0.29
R770 GND.n513 GND.n506 0.29
R771 GND.n471 GND.n464 0.29
R772 GND GND.n848 0.219
R773 GND.n429 GND 0.207
R774 GND.n108 GND.n105 0.197
R775 GND.n150 GND.n147 0.197
R776 GND.n192 GND.n189 0.197
R777 GND.n237 GND.n234 0.197
R778 GND.n279 GND.n276 0.197
R779 GND.n321 GND.n318 0.197
R780 GND.n363 GND.n360 0.197
R781 GND.n405 GND.n402 0.197
R782 GND.n833 GND.n830 0.197
R783 GND.n791 GND.n788 0.197
R784 GND.n746 GND.n743 0.197
R785 GND.n704 GND.n701 0.197
R786 GND.n659 GND.n656 0.197
R787 GND.n617 GND.n614 0.197
R788 GND.n575 GND.n572 0.197
R789 GND.n533 GND.n530 0.197
R790 GND.n491 GND.n488 0.197
R791 GND.n449 GND.n446 0.197
R792 GND.n118 GND.n117 0.196
R793 GND.n160 GND.n159 0.196
R794 GND.n205 GND.n204 0.196
R795 GND.n247 GND.n246 0.196
R796 GND.n289 GND.n288 0.196
R797 GND.n331 GND.n330 0.196
R798 GND.n373 GND.n372 0.196
R799 GND.n415 GND.n414 0.196
R800 GND.n820 GND.n819 0.196
R801 GND.n778 GND.n777 0.196
R802 GND.n733 GND.n732 0.196
R803 GND.n691 GND.n690 0.196
R804 GND.n646 GND.n645 0.196
R805 GND.n604 GND.n603 0.196
R806 GND.n562 GND.n561 0.196
R807 GND.n520 GND.n519 0.196
R808 GND.n478 GND.n477 0.196
R809 GND.n436 GND.n435 0.196
R810 GND.n12 GND.n9 0.181
R811 GND.n42 GND.n39 0.181
R812 GND.n72 GND.n69 0.181
R813 GND.n9 GND.n8 0.145
R814 GND.n17 GND.n12 0.145
R815 GND.n20 GND.n17 0.145
R816 GND.n23 GND.n20 0.145
R817 GND.n33 GND.n30 0.145
R818 GND.n36 GND.n33 0.145
R819 GND.n39 GND.n36 0.145
R820 GND.n47 GND.n42 0.145
R821 GND.n50 GND.n47 0.145
R822 GND.n53 GND.n50 0.145
R823 GND.n63 GND.n60 0.145
R824 GND.n66 GND.n63 0.145
R825 GND.n69 GND.n66 0.145
R826 GND.n77 GND.n72 0.145
R827 GND.n80 GND.n77 0.145
R828 GND.n83 GND.n80 0.145
R829 GND.n93 GND.n90 0.145
R830 GND.n96 GND.n93 0.145
R831 GND.n99 GND.n96 0.145
R832 GND.n102 GND.n99 0.145
R833 GND.n105 GND.n102 0.145
R834 GND.n111 GND.n108 0.145
R835 GND.n114 GND.n111 0.145
R836 GND.n119 GND.n114 0.145
R837 GND.n122 GND.n119 0.145
R838 GND.n125 GND.n122 0.145
R839 GND.n135 GND.n132 0.145
R840 GND.n138 GND.n135 0.145
R841 GND.n141 GND.n138 0.145
R842 GND.n144 GND.n141 0.145
R843 GND.n147 GND.n144 0.145
R844 GND.n153 GND.n150 0.145
R845 GND.n156 GND.n153 0.145
R846 GND.n161 GND.n156 0.145
R847 GND.n164 GND.n161 0.145
R848 GND.n167 GND.n164 0.145
R849 GND.n177 GND.n174 0.145
R850 GND.n180 GND.n177 0.145
R851 GND.n183 GND.n180 0.145
R852 GND.n186 GND.n183 0.145
R853 GND.n189 GND.n186 0.145
R854 GND.n195 GND.n192 0.145
R855 GND.n198 GND.n195 0.145
R856 GND.n206 GND.n198 0.145
R857 GND.n209 GND.n206 0.145
R858 GND.n212 GND.n209 0.145
R859 GND.n222 GND.n219 0.145
R860 GND.n225 GND.n222 0.145
R861 GND.n228 GND.n225 0.145
R862 GND.n231 GND.n228 0.145
R863 GND.n234 GND.n231 0.145
R864 GND.n240 GND.n237 0.145
R865 GND.n243 GND.n240 0.145
R866 GND.n248 GND.n243 0.145
R867 GND.n251 GND.n248 0.145
R868 GND.n254 GND.n251 0.145
R869 GND.n264 GND.n261 0.145
R870 GND.n267 GND.n264 0.145
R871 GND.n270 GND.n267 0.145
R872 GND.n273 GND.n270 0.145
R873 GND.n276 GND.n273 0.145
R874 GND.n282 GND.n279 0.145
R875 GND.n285 GND.n282 0.145
R876 GND.n290 GND.n285 0.145
R877 GND.n293 GND.n290 0.145
R878 GND.n296 GND.n293 0.145
R879 GND.n306 GND.n303 0.145
R880 GND.n309 GND.n306 0.145
R881 GND.n312 GND.n309 0.145
R882 GND.n315 GND.n312 0.145
R883 GND.n318 GND.n315 0.145
R884 GND.n324 GND.n321 0.145
R885 GND.n327 GND.n324 0.145
R886 GND.n332 GND.n327 0.145
R887 GND.n335 GND.n332 0.145
R888 GND.n338 GND.n335 0.145
R889 GND.n348 GND.n345 0.145
R890 GND.n351 GND.n348 0.145
R891 GND.n354 GND.n351 0.145
R892 GND.n357 GND.n354 0.145
R893 GND.n360 GND.n357 0.145
R894 GND.n366 GND.n363 0.145
R895 GND.n369 GND.n366 0.145
R896 GND.n374 GND.n369 0.145
R897 GND.n377 GND.n374 0.145
R898 GND.n380 GND.n377 0.145
R899 GND.n390 GND.n387 0.145
R900 GND.n393 GND.n390 0.145
R901 GND.n396 GND.n393 0.145
R902 GND.n399 GND.n396 0.145
R903 GND.n402 GND.n399 0.145
R904 GND.n408 GND.n405 0.145
R905 GND.n411 GND.n408 0.145
R906 GND.n416 GND.n411 0.145
R907 GND.n419 GND.n416 0.145
R908 GND.n426 GND.n419 0.145
R909 GND.n848 GND.n845 0.145
R910 GND.n845 GND.n842 0.145
R911 GND.n842 GND.n839 0.145
R912 GND.n839 GND.n836 0.145
R913 GND.n836 GND.n833 0.145
R914 GND.n830 GND.n827 0.145
R915 GND.n827 GND.n824 0.145
R916 GND.n824 GND.n821 0.145
R917 GND.n821 GND.n816 0.145
R918 GND.n816 GND.n813 0.145
R919 GND.n806 GND.n803 0.145
R920 GND.n803 GND.n800 0.145
R921 GND.n800 GND.n797 0.145
R922 GND.n797 GND.n794 0.145
R923 GND.n794 GND.n791 0.145
R924 GND.n788 GND.n785 0.145
R925 GND.n785 GND.n782 0.145
R926 GND.n782 GND.n779 0.145
R927 GND.n779 GND.n771 0.145
R928 GND.n771 GND.n768 0.145
R929 GND.n761 GND.n758 0.145
R930 GND.n758 GND.n755 0.145
R931 GND.n755 GND.n752 0.145
R932 GND.n752 GND.n749 0.145
R933 GND.n749 GND.n746 0.145
R934 GND.n743 GND.n740 0.145
R935 GND.n740 GND.n737 0.145
R936 GND.n737 GND.n734 0.145
R937 GND.n734 GND.n729 0.145
R938 GND.n729 GND.n726 0.145
R939 GND.n719 GND.n716 0.145
R940 GND.n716 GND.n713 0.145
R941 GND.n713 GND.n710 0.145
R942 GND.n710 GND.n707 0.145
R943 GND.n707 GND.n704 0.145
R944 GND.n701 GND.n698 0.145
R945 GND.n698 GND.n695 0.145
R946 GND.n695 GND.n692 0.145
R947 GND.n692 GND.n684 0.145
R948 GND.n684 GND.n681 0.145
R949 GND.n674 GND.n671 0.145
R950 GND.n671 GND.n668 0.145
R951 GND.n668 GND.n665 0.145
R952 GND.n665 GND.n662 0.145
R953 GND.n662 GND.n659 0.145
R954 GND.n656 GND.n653 0.145
R955 GND.n653 GND.n650 0.145
R956 GND.n650 GND.n647 0.145
R957 GND.n647 GND.n642 0.145
R958 GND.n642 GND.n639 0.145
R959 GND.n632 GND.n629 0.145
R960 GND.n629 GND.n626 0.145
R961 GND.n626 GND.n623 0.145
R962 GND.n623 GND.n620 0.145
R963 GND.n620 GND.n617 0.145
R964 GND.n614 GND.n611 0.145
R965 GND.n611 GND.n608 0.145
R966 GND.n608 GND.n605 0.145
R967 GND.n605 GND.n600 0.145
R968 GND.n600 GND.n597 0.145
R969 GND.n590 GND.n587 0.145
R970 GND.n587 GND.n584 0.145
R971 GND.n584 GND.n581 0.145
R972 GND.n581 GND.n578 0.145
R973 GND.n578 GND.n575 0.145
R974 GND.n572 GND.n569 0.145
R975 GND.n569 GND.n566 0.145
R976 GND.n566 GND.n563 0.145
R977 GND.n563 GND.n558 0.145
R978 GND.n558 GND.n555 0.145
R979 GND.n548 GND.n545 0.145
R980 GND.n545 GND.n542 0.145
R981 GND.n542 GND.n539 0.145
R982 GND.n539 GND.n536 0.145
R983 GND.n536 GND.n533 0.145
R984 GND.n530 GND.n527 0.145
R985 GND.n527 GND.n524 0.145
R986 GND.n524 GND.n521 0.145
R987 GND.n521 GND.n516 0.145
R988 GND.n516 GND.n513 0.145
R989 GND.n506 GND.n503 0.145
R990 GND.n503 GND.n500 0.145
R991 GND.n500 GND.n497 0.145
R992 GND.n497 GND.n494 0.145
R993 GND.n494 GND.n491 0.145
R994 GND.n488 GND.n485 0.145
R995 GND.n485 GND.n482 0.145
R996 GND.n482 GND.n479 0.145
R997 GND.n479 GND.n474 0.145
R998 GND.n474 GND.n471 0.145
R999 GND.n464 GND.n461 0.145
R1000 GND.n461 GND.n458 0.145
R1001 GND.n458 GND.n455 0.145
R1002 GND.n455 GND.n452 0.145
R1003 GND.n452 GND.n449 0.145
R1004 GND.n446 GND.n443 0.145
R1005 GND.n443 GND.n440 0.145
R1006 GND.n440 GND.n437 0.145
R1007 GND.n437 GND.n432 0.145
R1008 GND.n432 GND.n429 0.145
R1009 GND GND.n426 0.07
R1010 a_10219_989.n5 a_10219_989.t9 475.572
R1011 a_10219_989.n7 a_10219_989.t7 469.145
R1012 a_10219_989.n11 a_10219_989.t12 454.685
R1013 a_10219_989.n11 a_10219_989.t8 428.979
R1014 a_10219_989.n7 a_10219_989.t11 384.527
R1015 a_10219_989.n5 a_10219_989.t13 384.527
R1016 a_10219_989.n8 a_10219_989.t14 294.278
R1017 a_10219_989.n6 a_10219_989.t10 294.278
R1018 a_10219_989.n12 a_10219_989.t15 184.853
R1019 a_10219_989.n15 a_10219_989.n13 166.52
R1020 a_10219_989.n13 a_10219_989.n12 156.035
R1021 a_10219_989.n12 a_10219_989.n11 151.553
R1022 a_10219_989.n10 a_10219_989.n4 144.246
R1023 a_10219_989.n10 a_10219_989.n9 99.225
R1024 a_10219_989.n9 a_10219_989.n6 80.851
R1025 a_10219_989.n13 a_10219_989.n10 79.658
R1026 a_10219_989.n3 a_10219_989.n2 79.232
R1027 a_10219_989.n9 a_10219_989.n8 76
R1028 a_10219_989.n4 a_10219_989.n3 63.152
R1029 a_10219_989.n6 a_10219_989.n5 57.842
R1030 a_10219_989.n8 a_10219_989.n7 56.833
R1031 a_10219_989.n4 a_10219_989.n0 16.08
R1032 a_10219_989.n3 a_10219_989.n1 16.08
R1033 a_10219_989.n15 a_10219_989.n14 15.218
R1034 a_10219_989.n0 a_10219_989.t3 14.282
R1035 a_10219_989.n0 a_10219_989.t0 14.282
R1036 a_10219_989.n1 a_10219_989.t2 14.282
R1037 a_10219_989.n1 a_10219_989.t1 14.282
R1038 a_10219_989.n2 a_10219_989.t5 14.282
R1039 a_10219_989.n2 a_10219_989.t4 14.282
R1040 a_10219_989.n16 a_10219_989.n15 12.014
R1041 a_17533_1051.n3 a_17533_1051.n2 195.987
R1042 a_17533_1051.n4 a_17533_1051.t7 89.553
R1043 a_17533_1051.n2 a_17533_1051.n1 75.271
R1044 a_17533_1051.n4 a_17533_1051.n3 75.214
R1045 a_17533_1051.n2 a_17533_1051.n0 36.519
R1046 a_17533_1051.n3 a_17533_1051.t6 14.338
R1047 a_17533_1051.n0 a_17533_1051.t4 14.282
R1048 a_17533_1051.n0 a_17533_1051.t5 14.282
R1049 a_17533_1051.n1 a_17533_1051.t2 14.282
R1050 a_17533_1051.n1 a_17533_1051.t3 14.282
R1051 a_17533_1051.t0 a_17533_1051.n5 14.282
R1052 a_17533_1051.n5 a_17533_1051.t1 14.282
R1053 a_17533_1051.n5 a_17533_1051.n4 12.122
R1054 VDD.n940 VDD.n938 144.705
R1055 VDD.n1021 VDD.n1019 144.705
R1056 VDD.n1102 VDD.n1100 144.705
R1057 VDD.n1183 VDD.n1181 144.705
R1058 VDD.n1264 VDD.n1262 144.705
R1059 VDD.n1345 VDD.n1343 144.705
R1060 VDD.n1426 VDD.n1424 144.705
R1061 VDD.n1507 VDD.n1505 144.705
R1062 VDD.n1588 VDD.n1586 144.705
R1063 VDD.n758 VDD.n756 144.705
R1064 VDD.n835 VDD.n833 144.705
R1065 VDD.n677 VDD.n675 144.705
R1066 VDD.n596 VDD.n594 144.705
R1067 VDD.n515 VDD.n513 144.705
R1068 VDD.n434 VDD.n432 144.705
R1069 VDD.n353 VDD.n351 144.705
R1070 VDD.n272 VDD.n270 144.705
R1071 VDD.n191 VDD.n189 144.705
R1072 VDD.n130 VDD.n128 144.705
R1073 VDD.n76 VDD.n74 144.705
R1074 VDD.n39 VDD.n38 76
R1075 VDD.n43 VDD.n42 76
R1076 VDD.n47 VDD.n46 76
R1077 VDD.n51 VDD.n50 76
R1078 VDD.n78 VDD.n77 76
R1079 VDD.n82 VDD.n81 76
R1080 VDD.n86 VDD.n85 76
R1081 VDD.n90 VDD.n89 76
R1082 VDD.n94 VDD.n93 76
R1083 VDD.n98 VDD.n97 76
R1084 VDD.n102 VDD.n101 76
R1085 VDD.n106 VDD.n105 76
R1086 VDD.n132 VDD.n131 76
R1087 VDD.n137 VDD.n136 76
R1088 VDD.n142 VDD.n141 76
R1089 VDD.n148 VDD.n147 76
R1090 VDD.n153 VDD.n152 76
R1091 VDD.n158 VDD.n157 76
R1092 VDD.n163 VDD.n162 76
R1093 VDD.n167 VDD.n166 76
R1094 VDD.n193 VDD.n192 76
R1095 VDD.n197 VDD.n196 76
R1096 VDD.n201 VDD.n200 76
R1097 VDD.n206 VDD.n205 76
R1098 VDD.n213 VDD.n212 76
R1099 VDD.n218 VDD.n217 76
R1100 VDD.n223 VDD.n222 76
R1101 VDD.n230 VDD.n229 76
R1102 VDD.n235 VDD.n234 76
R1103 VDD.n240 VDD.n239 76
R1104 VDD.n244 VDD.n243 76
R1105 VDD.n248 VDD.n247 76
R1106 VDD.n274 VDD.n273 76
R1107 VDD.n278 VDD.n277 76
R1108 VDD.n282 VDD.n281 76
R1109 VDD.n287 VDD.n286 76
R1110 VDD.n294 VDD.n293 76
R1111 VDD.n299 VDD.n298 76
R1112 VDD.n304 VDD.n303 76
R1113 VDD.n311 VDD.n310 76
R1114 VDD.n316 VDD.n315 76
R1115 VDD.n321 VDD.n320 76
R1116 VDD.n325 VDD.n324 76
R1117 VDD.n329 VDD.n328 76
R1118 VDD.n355 VDD.n354 76
R1119 VDD.n359 VDD.n358 76
R1120 VDD.n363 VDD.n362 76
R1121 VDD.n368 VDD.n367 76
R1122 VDD.n375 VDD.n374 76
R1123 VDD.n380 VDD.n379 76
R1124 VDD.n385 VDD.n384 76
R1125 VDD.n392 VDD.n391 76
R1126 VDD.n397 VDD.n396 76
R1127 VDD.n402 VDD.n401 76
R1128 VDD.n406 VDD.n405 76
R1129 VDD.n410 VDD.n409 76
R1130 VDD.n436 VDD.n435 76
R1131 VDD.n440 VDD.n439 76
R1132 VDD.n444 VDD.n443 76
R1133 VDD.n449 VDD.n448 76
R1134 VDD.n456 VDD.n455 76
R1135 VDD.n461 VDD.n460 76
R1136 VDD.n466 VDD.n465 76
R1137 VDD.n473 VDD.n472 76
R1138 VDD.n478 VDD.n477 76
R1139 VDD.n483 VDD.n482 76
R1140 VDD.n487 VDD.n486 76
R1141 VDD.n491 VDD.n490 76
R1142 VDD.n517 VDD.n516 76
R1143 VDD.n521 VDD.n520 76
R1144 VDD.n525 VDD.n524 76
R1145 VDD.n530 VDD.n529 76
R1146 VDD.n537 VDD.n536 76
R1147 VDD.n542 VDD.n541 76
R1148 VDD.n547 VDD.n546 76
R1149 VDD.n554 VDD.n553 76
R1150 VDD.n559 VDD.n558 76
R1151 VDD.n564 VDD.n563 76
R1152 VDD.n568 VDD.n567 76
R1153 VDD.n572 VDD.n571 76
R1154 VDD.n598 VDD.n597 76
R1155 VDD.n602 VDD.n601 76
R1156 VDD.n606 VDD.n605 76
R1157 VDD.n611 VDD.n610 76
R1158 VDD.n618 VDD.n617 76
R1159 VDD.n623 VDD.n622 76
R1160 VDD.n628 VDD.n627 76
R1161 VDD.n635 VDD.n634 76
R1162 VDD.n640 VDD.n639 76
R1163 VDD.n645 VDD.n644 76
R1164 VDD.n649 VDD.n648 76
R1165 VDD.n653 VDD.n652 76
R1166 VDD.n679 VDD.n678 76
R1167 VDD.n683 VDD.n682 76
R1168 VDD.n687 VDD.n686 76
R1169 VDD.n692 VDD.n691 76
R1170 VDD.n699 VDD.n698 76
R1171 VDD.n704 VDD.n703 76
R1172 VDD.n709 VDD.n708 76
R1173 VDD.n716 VDD.n715 76
R1174 VDD.n721 VDD.n720 76
R1175 VDD.n726 VDD.n725 76
R1176 VDD.n730 VDD.n729 76
R1177 VDD.n734 VDD.n733 76
R1178 VDD.n760 VDD.n759 76
R1179 VDD.n764 VDD.n763 76
R1180 VDD.n768 VDD.n767 76
R1181 VDD.n773 VDD.n772 76
R1182 VDD.n780 VDD.n779 76
R1183 VDD.n785 VDD.n784 76
R1184 VDD.n790 VDD.n789 76
R1185 VDD.n797 VDD.n796 76
R1186 VDD.n802 VDD.n801 76
R1187 VDD.n807 VDD.n806 76
R1188 VDD.n811 VDD.n810 76
R1189 VDD.n837 VDD.n836 76
R1190 VDD.n1645 VDD.n1644 76
R1191 VDD.n1641 VDD.n1640 76
R1192 VDD.n1637 VDD.n1636 76
R1193 VDD.n1633 VDD.n1632 76
R1194 VDD.n1628 VDD.n1627 76
R1195 VDD.n1621 VDD.n1620 76
R1196 VDD.n1616 VDD.n1615 76
R1197 VDD.n1611 VDD.n1610 76
R1198 VDD.n1604 VDD.n1603 76
R1199 VDD.n1599 VDD.n1598 76
R1200 VDD.n1594 VDD.n1593 76
R1201 VDD.n1590 VDD.n1589 76
R1202 VDD.n1564 VDD.n1563 76
R1203 VDD.n1560 VDD.n1559 76
R1204 VDD.n1556 VDD.n1555 76
R1205 VDD.n1552 VDD.n1551 76
R1206 VDD.n1547 VDD.n1546 76
R1207 VDD.n1540 VDD.n1539 76
R1208 VDD.n1535 VDD.n1534 76
R1209 VDD.n1530 VDD.n1529 76
R1210 VDD.n1523 VDD.n1522 76
R1211 VDD.n1518 VDD.n1517 76
R1212 VDD.n1513 VDD.n1512 76
R1213 VDD.n1509 VDD.n1508 76
R1214 VDD.n1483 VDD.n1482 76
R1215 VDD.n1479 VDD.n1478 76
R1216 VDD.n1475 VDD.n1474 76
R1217 VDD.n1471 VDD.n1470 76
R1218 VDD.n1466 VDD.n1465 76
R1219 VDD.n1459 VDD.n1458 76
R1220 VDD.n1454 VDD.n1453 76
R1221 VDD.n1449 VDD.n1448 76
R1222 VDD.n1442 VDD.n1441 76
R1223 VDD.n1437 VDD.n1436 76
R1224 VDD.n1432 VDD.n1431 76
R1225 VDD.n1428 VDD.n1427 76
R1226 VDD.n1402 VDD.n1401 76
R1227 VDD.n1398 VDD.n1397 76
R1228 VDD.n1394 VDD.n1393 76
R1229 VDD.n1390 VDD.n1389 76
R1230 VDD.n1385 VDD.n1384 76
R1231 VDD.n1378 VDD.n1377 76
R1232 VDD.n1373 VDD.n1372 76
R1233 VDD.n1368 VDD.n1367 76
R1234 VDD.n1361 VDD.n1360 76
R1235 VDD.n1356 VDD.n1355 76
R1236 VDD.n1351 VDD.n1350 76
R1237 VDD.n1347 VDD.n1346 76
R1238 VDD.n1321 VDD.n1320 76
R1239 VDD.n1317 VDD.n1316 76
R1240 VDD.n1313 VDD.n1312 76
R1241 VDD.n1309 VDD.n1308 76
R1242 VDD.n1304 VDD.n1303 76
R1243 VDD.n1297 VDD.n1296 76
R1244 VDD.n1292 VDD.n1291 76
R1245 VDD.n1287 VDD.n1286 76
R1246 VDD.n1280 VDD.n1279 76
R1247 VDD.n1275 VDD.n1274 76
R1248 VDD.n1270 VDD.n1269 76
R1249 VDD.n1266 VDD.n1265 76
R1250 VDD.n1240 VDD.n1239 76
R1251 VDD.n1236 VDD.n1235 76
R1252 VDD.n1232 VDD.n1231 76
R1253 VDD.n1228 VDD.n1227 76
R1254 VDD.n1223 VDD.n1222 76
R1255 VDD.n1216 VDD.n1215 76
R1256 VDD.n1211 VDD.n1210 76
R1257 VDD.n1206 VDD.n1205 76
R1258 VDD.n1199 VDD.n1198 76
R1259 VDD.n1194 VDD.n1193 76
R1260 VDD.n1189 VDD.n1188 76
R1261 VDD.n1185 VDD.n1184 76
R1262 VDD.n1159 VDD.n1158 76
R1263 VDD.n1155 VDD.n1154 76
R1264 VDD.n1151 VDD.n1150 76
R1265 VDD.n1147 VDD.n1146 76
R1266 VDD.n1142 VDD.n1141 76
R1267 VDD.n1135 VDD.n1134 76
R1268 VDD.n1130 VDD.n1129 76
R1269 VDD.n1125 VDD.n1124 76
R1270 VDD.n1118 VDD.n1117 76
R1271 VDD.n1113 VDD.n1112 76
R1272 VDD.n1108 VDD.n1107 76
R1273 VDD.n1104 VDD.n1103 76
R1274 VDD.n1078 VDD.n1077 76
R1275 VDD.n1074 VDD.n1073 76
R1276 VDD.n1070 VDD.n1069 76
R1277 VDD.n1066 VDD.n1065 76
R1278 VDD.n1061 VDD.n1060 76
R1279 VDD.n1054 VDD.n1053 76
R1280 VDD.n1049 VDD.n1048 76
R1281 VDD.n1044 VDD.n1043 76
R1282 VDD.n1037 VDD.n1036 76
R1283 VDD.n1032 VDD.n1031 76
R1284 VDD.n1027 VDD.n1026 76
R1285 VDD.n1023 VDD.n1022 76
R1286 VDD.n997 VDD.n996 76
R1287 VDD.n993 VDD.n992 76
R1288 VDD.n989 VDD.n988 76
R1289 VDD.n985 VDD.n984 76
R1290 VDD.n980 VDD.n979 76
R1291 VDD.n973 VDD.n972 76
R1292 VDD.n968 VDD.n967 76
R1293 VDD.n963 VDD.n962 76
R1294 VDD.n956 VDD.n955 76
R1295 VDD.n951 VDD.n950 76
R1296 VDD.n946 VDD.n945 76
R1297 VDD.n942 VDD.n941 76
R1298 VDD.n915 VDD.n914 76
R1299 VDD.n911 VDD.n910 76
R1300 VDD.n907 VDD.n906 76
R1301 VDD.n903 VDD.n902 76
R1302 VDD.n898 VDD.n897 76
R1303 VDD.n891 VDD.n890 76
R1304 VDD.n886 VDD.n885 76
R1305 VDD.n881 VDD.n880 76
R1306 VDD.n874 VDD.n873 76
R1307 VDD.n869 VDD.n868 76
R1308 VDD.n864 VDD.n863 76
R1309 VDD.n860 VDD.n859 76
R1310 VDD.n203 VDD.n202 64.064
R1311 VDD.n284 VDD.n283 64.064
R1312 VDD.n365 VDD.n364 64.064
R1313 VDD.n446 VDD.n445 64.064
R1314 VDD.n527 VDD.n526 64.064
R1315 VDD.n608 VDD.n607 64.064
R1316 VDD.n689 VDD.n688 64.064
R1317 VDD.n770 VDD.n769 64.064
R1318 VDD.n1630 VDD.n1629 64.064
R1319 VDD.n1549 VDD.n1548 64.064
R1320 VDD.n1468 VDD.n1467 64.064
R1321 VDD.n1387 VDD.n1386 64.064
R1322 VDD.n1306 VDD.n1305 64.064
R1323 VDD.n1225 VDD.n1224 64.064
R1324 VDD.n1144 VDD.n1143 64.064
R1325 VDD.n1063 VDD.n1062 64.064
R1326 VDD.n982 VDD.n981 64.064
R1327 VDD.n900 VDD.n899 64.064
R1328 VDD.n232 VDD.n231 59.488
R1329 VDD.n313 VDD.n312 59.488
R1330 VDD.n394 VDD.n393 59.488
R1331 VDD.n475 VDD.n474 59.488
R1332 VDD.n556 VDD.n555 59.488
R1333 VDD.n637 VDD.n636 59.488
R1334 VDD.n718 VDD.n717 59.488
R1335 VDD.n799 VDD.n798 59.488
R1336 VDD.n1601 VDD.n1600 59.488
R1337 VDD.n1520 VDD.n1519 59.488
R1338 VDD.n1439 VDD.n1438 59.488
R1339 VDD.n1358 VDD.n1357 59.488
R1340 VDD.n1277 VDD.n1276 59.488
R1341 VDD.n1196 VDD.n1195 59.488
R1342 VDD.n1115 VDD.n1114 59.488
R1343 VDD.n1034 VDD.n1033 59.488
R1344 VDD.n953 VDD.n952 59.488
R1345 VDD.n871 VDD.n870 59.488
R1346 VDD.n159 VDD.t40 55.465
R1347 VDD.n133 VDD.t48 55.465
R1348 VDD.n865 VDD.t78 55.106
R1349 VDD.n947 VDD.t57 55.106
R1350 VDD.n1028 VDD.t104 55.106
R1351 VDD.n1109 VDD.t9 55.106
R1352 VDD.n1190 VDD.t109 55.106
R1353 VDD.n1271 VDD.t38 55.106
R1354 VDD.n1352 VDD.t77 55.106
R1355 VDD.n1433 VDD.t58 55.106
R1356 VDD.n1514 VDD.t61 55.106
R1357 VDD.n1595 VDD.t95 55.106
R1358 VDD.n803 VDD.t73 55.106
R1359 VDD.n722 VDD.t84 55.106
R1360 VDD.n641 VDD.t76 55.106
R1361 VDD.n560 VDD.t13 55.106
R1362 VDD.n479 VDD.t103 55.106
R1363 VDD.n398 VDD.t21 55.106
R1364 VDD.n317 VDD.t35 55.106
R1365 VDD.n236 VDD.t45 55.106
R1366 VDD.n906 VDD.t46 55.106
R1367 VDD.n988 VDD.t110 55.106
R1368 VDD.n1069 VDD.t92 55.106
R1369 VDD.n1150 VDD.t106 55.106
R1370 VDD.n1231 VDD.t7 55.106
R1371 VDD.n1312 VDD.t86 55.106
R1372 VDD.n1393 VDD.t53 55.106
R1373 VDD.n1474 VDD.t4 55.106
R1374 VDD.n1555 VDD.t71 55.106
R1375 VDD.n1636 VDD.t65 55.106
R1376 VDD.n767 VDD.t50 55.106
R1377 VDD.n686 VDD.t72 55.106
R1378 VDD.n605 VDD.t82 55.106
R1379 VDD.n524 VDD.t100 55.106
R1380 VDD.n443 VDD.t97 55.106
R1381 VDD.n362 VDD.t10 55.106
R1382 VDD.n281 VDD.t17 55.106
R1383 VDD.n200 VDD.t101 55.106
R1384 VDD.n144 VDD.n143 41.183
R1385 VDD.n876 VDD.n875 40.824
R1386 VDD.n896 VDD.n895 40.824
R1387 VDD.n958 VDD.n957 40.824
R1388 VDD.n978 VDD.n977 40.824
R1389 VDD.n1039 VDD.n1038 40.824
R1390 VDD.n1059 VDD.n1058 40.824
R1391 VDD.n1120 VDD.n1119 40.824
R1392 VDD.n1140 VDD.n1139 40.824
R1393 VDD.n1201 VDD.n1200 40.824
R1394 VDD.n1221 VDD.n1220 40.824
R1395 VDD.n1282 VDD.n1281 40.824
R1396 VDD.n1302 VDD.n1301 40.824
R1397 VDD.n1363 VDD.n1362 40.824
R1398 VDD.n1383 VDD.n1382 40.824
R1399 VDD.n1444 VDD.n1443 40.824
R1400 VDD.n1464 VDD.n1463 40.824
R1401 VDD.n1525 VDD.n1524 40.824
R1402 VDD.n1545 VDD.n1544 40.824
R1403 VDD.n1606 VDD.n1605 40.824
R1404 VDD.n1626 VDD.n1625 40.824
R1405 VDD.n792 VDD.n791 40.824
R1406 VDD.n778 VDD.n777 40.824
R1407 VDD.n711 VDD.n710 40.824
R1408 VDD.n697 VDD.n696 40.824
R1409 VDD.n630 VDD.n629 40.824
R1410 VDD.n616 VDD.n615 40.824
R1411 VDD.n549 VDD.n548 40.824
R1412 VDD.n535 VDD.n534 40.824
R1413 VDD.n468 VDD.n467 40.824
R1414 VDD.n454 VDD.n453 40.824
R1415 VDD.n387 VDD.n386 40.824
R1416 VDD.n373 VDD.n372 40.824
R1417 VDD.n306 VDD.n305 40.824
R1418 VDD.n292 VDD.n291 40.824
R1419 VDD.n225 VDD.n224 40.824
R1420 VDD.n211 VDD.n210 40.824
R1421 VDD.n1002 VDD.n1001 36.774
R1422 VDD.n1083 VDD.n1082 36.774
R1423 VDD.n1164 VDD.n1163 36.774
R1424 VDD.n1245 VDD.n1244 36.774
R1425 VDD.n1326 VDD.n1325 36.774
R1426 VDD.n1407 VDD.n1406 36.774
R1427 VDD.n1488 VDD.n1487 36.774
R1428 VDD.n1569 VDD.n1568 36.774
R1429 VDD.n816 VDD.n815 36.774
R1430 VDD.n739 VDD.n738 36.774
R1431 VDD.n658 VDD.n657 36.774
R1432 VDD.n577 VDD.n576 36.774
R1433 VDD.n496 VDD.n495 36.774
R1434 VDD.n415 VDD.n414 36.774
R1435 VDD.n334 VDD.n333 36.774
R1436 VDD.n253 VDD.n252 36.774
R1437 VDD.n172 VDD.n171 36.774
R1438 VDD.n111 VDD.n110 36.774
R1439 VDD.n56 VDD.n55 36.774
R1440 VDD.n931 VDD.n930 36.774
R1441 VDD.n139 VDD.n138 36.608
R1442 VDD.n34 VDD.n33 34.942
R1443 VDD.n155 VDD.n154 32.032
R1444 VDD.n208 VDD.n207 27.456
R1445 VDD.n289 VDD.n288 27.456
R1446 VDD.n370 VDD.n369 27.456
R1447 VDD.n451 VDD.n450 27.456
R1448 VDD.n532 VDD.n531 27.456
R1449 VDD.n613 VDD.n612 27.456
R1450 VDD.n694 VDD.n693 27.456
R1451 VDD.n775 VDD.n774 27.456
R1452 VDD.n1623 VDD.n1622 27.456
R1453 VDD.n1542 VDD.n1541 27.456
R1454 VDD.n1461 VDD.n1460 27.456
R1455 VDD.n1380 VDD.n1379 27.456
R1456 VDD.n1299 VDD.n1298 27.456
R1457 VDD.n1218 VDD.n1217 27.456
R1458 VDD.n1137 VDD.n1136 27.456
R1459 VDD.n1056 VDD.n1055 27.456
R1460 VDD.n975 VDD.n974 27.456
R1461 VDD.n893 VDD.n892 27.456
R1462 VDD.n227 VDD.n226 22.88
R1463 VDD.n308 VDD.n307 22.88
R1464 VDD.n389 VDD.n388 22.88
R1465 VDD.n470 VDD.n469 22.88
R1466 VDD.n551 VDD.n550 22.88
R1467 VDD.n632 VDD.n631 22.88
R1468 VDD.n713 VDD.n712 22.88
R1469 VDD.n794 VDD.n793 22.88
R1470 VDD.n1608 VDD.n1607 22.88
R1471 VDD.n1527 VDD.n1526 22.88
R1472 VDD.n1446 VDD.n1445 22.88
R1473 VDD.n1365 VDD.n1364 22.88
R1474 VDD.n1284 VDD.n1283 22.88
R1475 VDD.n1203 VDD.n1202 22.88
R1476 VDD.n1122 VDD.n1121 22.88
R1477 VDD.n1041 VDD.n1040 22.88
R1478 VDD.n960 VDD.n959 22.88
R1479 VDD.n878 VDD.n877 22.88
R1480 VDD.n859 VDD.n856 21.841
R1481 VDD.n23 VDD.n20 21.841
R1482 VDD.n875 VDD.t44 14.282
R1483 VDD.n875 VDD.t55 14.282
R1484 VDD.n895 VDD.t18 14.282
R1485 VDD.n895 VDD.t75 14.282
R1486 VDD.n957 VDD.t27 14.282
R1487 VDD.n957 VDD.t63 14.282
R1488 VDD.n977 VDD.t67 14.282
R1489 VDD.n977 VDD.t26 14.282
R1490 VDD.n1038 VDD.t19 14.282
R1491 VDD.n1038 VDD.t15 14.282
R1492 VDD.n1058 VDD.t54 14.282
R1493 VDD.n1058 VDD.t83 14.282
R1494 VDD.n1119 VDD.t32 14.282
R1495 VDD.n1119 VDD.t1 14.282
R1496 VDD.n1139 VDD.t105 14.282
R1497 VDD.n1139 VDD.t30 14.282
R1498 VDD.n1200 VDD.t74 14.282
R1499 VDD.n1200 VDD.t81 14.282
R1500 VDD.n1220 VDD.t87 14.282
R1501 VDD.n1220 VDD.t5 14.282
R1502 VDD.n1281 VDD.t8 14.282
R1503 VDD.n1281 VDD.t42 14.282
R1504 VDD.n1301 VDD.t56 14.282
R1505 VDD.n1301 VDD.t94 14.282
R1506 VDD.n1362 VDD.t62 14.282
R1507 VDD.n1362 VDD.t16 14.282
R1508 VDD.n1382 VDD.t20 14.282
R1509 VDD.n1382 VDD.t79 14.282
R1510 VDD.n1443 VDD.t31 14.282
R1511 VDD.n1443 VDD.t59 14.282
R1512 VDD.n1463 VDD.t66 14.282
R1513 VDD.n1463 VDD.t23 14.282
R1514 VDD.n1524 VDD.t90 14.282
R1515 VDD.n1524 VDD.t60 14.282
R1516 VDD.n1544 VDD.t89 14.282
R1517 VDD.n1544 VDD.t88 14.282
R1518 VDD.n1605 VDD.t29 14.282
R1519 VDD.n1605 VDD.t93 14.282
R1520 VDD.n1625 VDD.t108 14.282
R1521 VDD.n1625 VDD.t28 14.282
R1522 VDD.n791 VDD.t51 14.282
R1523 VDD.n791 VDD.t69 14.282
R1524 VDD.n777 VDD.t49 14.282
R1525 VDD.n777 VDD.t107 14.282
R1526 VDD.n710 VDD.t2 14.282
R1527 VDD.n710 VDD.t91 14.282
R1528 VDD.n696 VDD.t0 14.282
R1529 VDD.n696 VDD.t68 14.282
R1530 VDD.n629 VDD.t64 14.282
R1531 VDD.n629 VDD.t52 14.282
R1532 VDD.n615 VDD.t37 14.282
R1533 VDD.n615 VDD.t6 14.282
R1534 VDD.n548 VDD.t24 14.282
R1535 VDD.n548 VDD.t102 14.282
R1536 VDD.n534 VDD.t99 14.282
R1537 VDD.n534 VDD.t25 14.282
R1538 VDD.n467 VDD.t70 14.282
R1539 VDD.n467 VDD.t14 14.282
R1540 VDD.n453 VDD.t96 14.282
R1541 VDD.n453 VDD.t85 14.282
R1542 VDD.n386 VDD.t34 14.282
R1543 VDD.n386 VDD.t22 14.282
R1544 VDD.n372 VDD.t12 14.282
R1545 VDD.n372 VDD.t33 14.282
R1546 VDD.n305 VDD.t11 14.282
R1547 VDD.n305 VDD.t36 14.282
R1548 VDD.n291 VDD.t43 14.282
R1549 VDD.n291 VDD.t80 14.282
R1550 VDD.n224 VDD.t3 14.282
R1551 VDD.n224 VDD.t41 14.282
R1552 VDD.n210 VDD.t98 14.282
R1553 VDD.n210 VDD.t111 14.282
R1554 VDD.n143 VDD.t47 14.282
R1555 VDD.n143 VDD.t39 14.282
R1556 VDD.n856 VDD.n839 14.167
R1557 VDD.n839 VDD.n838 14.167
R1558 VDD.n1017 VDD.n999 14.167
R1559 VDD.n999 VDD.n998 14.167
R1560 VDD.n1098 VDD.n1080 14.167
R1561 VDD.n1080 VDD.n1079 14.167
R1562 VDD.n1179 VDD.n1161 14.167
R1563 VDD.n1161 VDD.n1160 14.167
R1564 VDD.n1260 VDD.n1242 14.167
R1565 VDD.n1242 VDD.n1241 14.167
R1566 VDD.n1341 VDD.n1323 14.167
R1567 VDD.n1323 VDD.n1322 14.167
R1568 VDD.n1422 VDD.n1404 14.167
R1569 VDD.n1404 VDD.n1403 14.167
R1570 VDD.n1503 VDD.n1485 14.167
R1571 VDD.n1485 VDD.n1484 14.167
R1572 VDD.n1584 VDD.n1566 14.167
R1573 VDD.n1566 VDD.n1565 14.167
R1574 VDD.n831 VDD.n813 14.167
R1575 VDD.n813 VDD.n812 14.167
R1576 VDD.n754 VDD.n736 14.167
R1577 VDD.n736 VDD.n735 14.167
R1578 VDD.n673 VDD.n655 14.167
R1579 VDD.n655 VDD.n654 14.167
R1580 VDD.n592 VDD.n574 14.167
R1581 VDD.n574 VDD.n573 14.167
R1582 VDD.n511 VDD.n493 14.167
R1583 VDD.n493 VDD.n492 14.167
R1584 VDD.n430 VDD.n412 14.167
R1585 VDD.n412 VDD.n411 14.167
R1586 VDD.n349 VDD.n331 14.167
R1587 VDD.n331 VDD.n330 14.167
R1588 VDD.n268 VDD.n250 14.167
R1589 VDD.n250 VDD.n249 14.167
R1590 VDD.n187 VDD.n169 14.167
R1591 VDD.n169 VDD.n168 14.167
R1592 VDD.n126 VDD.n108 14.167
R1593 VDD.n108 VDD.n107 14.167
R1594 VDD.n72 VDD.n53 14.167
R1595 VDD.n53 VDD.n52 14.167
R1596 VDD.n936 VDD.n917 14.167
R1597 VDD.n917 VDD.n916 14.167
R1598 VDD.n20 VDD.n19 14.167
R1599 VDD.n19 VDD.n17 14.167
R1600 VDD.n32 VDD.n29 14.167
R1601 VDD.n29 VDD.n28 14.167
R1602 VDD.n77 VDD.n73 14.167
R1603 VDD.n131 VDD.n127 14.167
R1604 VDD.n192 VDD.n188 14.167
R1605 VDD.n273 VDD.n269 14.167
R1606 VDD.n354 VDD.n350 14.167
R1607 VDD.n435 VDD.n431 14.167
R1608 VDD.n516 VDD.n512 14.167
R1609 VDD.n597 VDD.n593 14.167
R1610 VDD.n678 VDD.n674 14.167
R1611 VDD.n759 VDD.n755 14.167
R1612 VDD.n836 VDD.n832 14.167
R1613 VDD.n1589 VDD.n1585 14.167
R1614 VDD.n1508 VDD.n1504 14.167
R1615 VDD.n1427 VDD.n1423 14.167
R1616 VDD.n1346 VDD.n1342 14.167
R1617 VDD.n1265 VDD.n1261 14.167
R1618 VDD.n1184 VDD.n1180 14.167
R1619 VDD.n1103 VDD.n1099 14.167
R1620 VDD.n1022 VDD.n1018 14.167
R1621 VDD.n941 VDD.n937 14.167
R1622 VDD.n220 VDD.n219 13.728
R1623 VDD.n301 VDD.n300 13.728
R1624 VDD.n382 VDD.n381 13.728
R1625 VDD.n463 VDD.n462 13.728
R1626 VDD.n544 VDD.n543 13.728
R1627 VDD.n625 VDD.n624 13.728
R1628 VDD.n706 VDD.n705 13.728
R1629 VDD.n787 VDD.n786 13.728
R1630 VDD.n1613 VDD.n1612 13.728
R1631 VDD.n1532 VDD.n1531 13.728
R1632 VDD.n1451 VDD.n1450 13.728
R1633 VDD.n1370 VDD.n1369 13.728
R1634 VDD.n1289 VDD.n1288 13.728
R1635 VDD.n1208 VDD.n1207 13.728
R1636 VDD.n1127 VDD.n1126 13.728
R1637 VDD.n1046 VDD.n1045 13.728
R1638 VDD.n965 VDD.n964 13.728
R1639 VDD.n883 VDD.n882 13.728
R1640 VDD.n23 VDD.n22 13.653
R1641 VDD.n22 VDD.n21 13.653
R1642 VDD.n32 VDD.n31 13.653
R1643 VDD.n31 VDD.n30 13.653
R1644 VDD.n29 VDD.n25 13.653
R1645 VDD.n25 VDD.n24 13.653
R1646 VDD.n28 VDD.n27 13.653
R1647 VDD.n27 VDD.n26 13.653
R1648 VDD.n38 VDD.n37 13.653
R1649 VDD.n37 VDD.n36 13.653
R1650 VDD.n42 VDD.n41 13.653
R1651 VDD.n41 VDD.n40 13.653
R1652 VDD.n46 VDD.n45 13.653
R1653 VDD.n45 VDD.n44 13.653
R1654 VDD.n50 VDD.n49 13.653
R1655 VDD.n49 VDD.n48 13.653
R1656 VDD.n77 VDD.n76 13.653
R1657 VDD.n76 VDD.n75 13.653
R1658 VDD.n81 VDD.n80 13.653
R1659 VDD.n80 VDD.n79 13.653
R1660 VDD.n85 VDD.n84 13.653
R1661 VDD.n84 VDD.n83 13.653
R1662 VDD.n89 VDD.n88 13.653
R1663 VDD.n88 VDD.n87 13.653
R1664 VDD.n93 VDD.n92 13.653
R1665 VDD.n92 VDD.n91 13.653
R1666 VDD.n97 VDD.n96 13.653
R1667 VDD.n96 VDD.n95 13.653
R1668 VDD.n101 VDD.n100 13.653
R1669 VDD.n100 VDD.n99 13.653
R1670 VDD.n105 VDD.n104 13.653
R1671 VDD.n104 VDD.n103 13.653
R1672 VDD.n131 VDD.n130 13.653
R1673 VDD.n130 VDD.n129 13.653
R1674 VDD.n136 VDD.n135 13.653
R1675 VDD.n135 VDD.n134 13.653
R1676 VDD.n141 VDD.n140 13.653
R1677 VDD.n140 VDD.n139 13.653
R1678 VDD.n147 VDD.n146 13.653
R1679 VDD.n146 VDD.n145 13.653
R1680 VDD.n152 VDD.n151 13.653
R1681 VDD.n151 VDD.n150 13.653
R1682 VDD.n157 VDD.n156 13.653
R1683 VDD.n156 VDD.n155 13.653
R1684 VDD.n162 VDD.n161 13.653
R1685 VDD.n161 VDD.n160 13.653
R1686 VDD.n166 VDD.n165 13.653
R1687 VDD.n165 VDD.n164 13.653
R1688 VDD.n192 VDD.n191 13.653
R1689 VDD.n191 VDD.n190 13.653
R1690 VDD.n196 VDD.n195 13.653
R1691 VDD.n195 VDD.n194 13.653
R1692 VDD.n200 VDD.n199 13.653
R1693 VDD.n199 VDD.n198 13.653
R1694 VDD.n205 VDD.n204 13.653
R1695 VDD.n204 VDD.n203 13.653
R1696 VDD.n212 VDD.n209 13.653
R1697 VDD.n209 VDD.n208 13.653
R1698 VDD.n217 VDD.n216 13.653
R1699 VDD.n216 VDD.n215 13.653
R1700 VDD.n222 VDD.n221 13.653
R1701 VDD.n221 VDD.n220 13.653
R1702 VDD.n229 VDD.n228 13.653
R1703 VDD.n228 VDD.n227 13.653
R1704 VDD.n234 VDD.n233 13.653
R1705 VDD.n233 VDD.n232 13.653
R1706 VDD.n239 VDD.n238 13.653
R1707 VDD.n238 VDD.n237 13.653
R1708 VDD.n243 VDD.n242 13.653
R1709 VDD.n242 VDD.n241 13.653
R1710 VDD.n247 VDD.n246 13.653
R1711 VDD.n246 VDD.n245 13.653
R1712 VDD.n273 VDD.n272 13.653
R1713 VDD.n272 VDD.n271 13.653
R1714 VDD.n277 VDD.n276 13.653
R1715 VDD.n276 VDD.n275 13.653
R1716 VDD.n281 VDD.n280 13.653
R1717 VDD.n280 VDD.n279 13.653
R1718 VDD.n286 VDD.n285 13.653
R1719 VDD.n285 VDD.n284 13.653
R1720 VDD.n293 VDD.n290 13.653
R1721 VDD.n290 VDD.n289 13.653
R1722 VDD.n298 VDD.n297 13.653
R1723 VDD.n297 VDD.n296 13.653
R1724 VDD.n303 VDD.n302 13.653
R1725 VDD.n302 VDD.n301 13.653
R1726 VDD.n310 VDD.n309 13.653
R1727 VDD.n309 VDD.n308 13.653
R1728 VDD.n315 VDD.n314 13.653
R1729 VDD.n314 VDD.n313 13.653
R1730 VDD.n320 VDD.n319 13.653
R1731 VDD.n319 VDD.n318 13.653
R1732 VDD.n324 VDD.n323 13.653
R1733 VDD.n323 VDD.n322 13.653
R1734 VDD.n328 VDD.n327 13.653
R1735 VDD.n327 VDD.n326 13.653
R1736 VDD.n354 VDD.n353 13.653
R1737 VDD.n353 VDD.n352 13.653
R1738 VDD.n358 VDD.n357 13.653
R1739 VDD.n357 VDD.n356 13.653
R1740 VDD.n362 VDD.n361 13.653
R1741 VDD.n361 VDD.n360 13.653
R1742 VDD.n367 VDD.n366 13.653
R1743 VDD.n366 VDD.n365 13.653
R1744 VDD.n374 VDD.n371 13.653
R1745 VDD.n371 VDD.n370 13.653
R1746 VDD.n379 VDD.n378 13.653
R1747 VDD.n378 VDD.n377 13.653
R1748 VDD.n384 VDD.n383 13.653
R1749 VDD.n383 VDD.n382 13.653
R1750 VDD.n391 VDD.n390 13.653
R1751 VDD.n390 VDD.n389 13.653
R1752 VDD.n396 VDD.n395 13.653
R1753 VDD.n395 VDD.n394 13.653
R1754 VDD.n401 VDD.n400 13.653
R1755 VDD.n400 VDD.n399 13.653
R1756 VDD.n405 VDD.n404 13.653
R1757 VDD.n404 VDD.n403 13.653
R1758 VDD.n409 VDD.n408 13.653
R1759 VDD.n408 VDD.n407 13.653
R1760 VDD.n435 VDD.n434 13.653
R1761 VDD.n434 VDD.n433 13.653
R1762 VDD.n439 VDD.n438 13.653
R1763 VDD.n438 VDD.n437 13.653
R1764 VDD.n443 VDD.n442 13.653
R1765 VDD.n442 VDD.n441 13.653
R1766 VDD.n448 VDD.n447 13.653
R1767 VDD.n447 VDD.n446 13.653
R1768 VDD.n455 VDD.n452 13.653
R1769 VDD.n452 VDD.n451 13.653
R1770 VDD.n460 VDD.n459 13.653
R1771 VDD.n459 VDD.n458 13.653
R1772 VDD.n465 VDD.n464 13.653
R1773 VDD.n464 VDD.n463 13.653
R1774 VDD.n472 VDD.n471 13.653
R1775 VDD.n471 VDD.n470 13.653
R1776 VDD.n477 VDD.n476 13.653
R1777 VDD.n476 VDD.n475 13.653
R1778 VDD.n482 VDD.n481 13.653
R1779 VDD.n481 VDD.n480 13.653
R1780 VDD.n486 VDD.n485 13.653
R1781 VDD.n485 VDD.n484 13.653
R1782 VDD.n490 VDD.n489 13.653
R1783 VDD.n489 VDD.n488 13.653
R1784 VDD.n516 VDD.n515 13.653
R1785 VDD.n515 VDD.n514 13.653
R1786 VDD.n520 VDD.n519 13.653
R1787 VDD.n519 VDD.n518 13.653
R1788 VDD.n524 VDD.n523 13.653
R1789 VDD.n523 VDD.n522 13.653
R1790 VDD.n529 VDD.n528 13.653
R1791 VDD.n528 VDD.n527 13.653
R1792 VDD.n536 VDD.n533 13.653
R1793 VDD.n533 VDD.n532 13.653
R1794 VDD.n541 VDD.n540 13.653
R1795 VDD.n540 VDD.n539 13.653
R1796 VDD.n546 VDD.n545 13.653
R1797 VDD.n545 VDD.n544 13.653
R1798 VDD.n553 VDD.n552 13.653
R1799 VDD.n552 VDD.n551 13.653
R1800 VDD.n558 VDD.n557 13.653
R1801 VDD.n557 VDD.n556 13.653
R1802 VDD.n563 VDD.n562 13.653
R1803 VDD.n562 VDD.n561 13.653
R1804 VDD.n567 VDD.n566 13.653
R1805 VDD.n566 VDD.n565 13.653
R1806 VDD.n571 VDD.n570 13.653
R1807 VDD.n570 VDD.n569 13.653
R1808 VDD.n597 VDD.n596 13.653
R1809 VDD.n596 VDD.n595 13.653
R1810 VDD.n601 VDD.n600 13.653
R1811 VDD.n600 VDD.n599 13.653
R1812 VDD.n605 VDD.n604 13.653
R1813 VDD.n604 VDD.n603 13.653
R1814 VDD.n610 VDD.n609 13.653
R1815 VDD.n609 VDD.n608 13.653
R1816 VDD.n617 VDD.n614 13.653
R1817 VDD.n614 VDD.n613 13.653
R1818 VDD.n622 VDD.n621 13.653
R1819 VDD.n621 VDD.n620 13.653
R1820 VDD.n627 VDD.n626 13.653
R1821 VDD.n626 VDD.n625 13.653
R1822 VDD.n634 VDD.n633 13.653
R1823 VDD.n633 VDD.n632 13.653
R1824 VDD.n639 VDD.n638 13.653
R1825 VDD.n638 VDD.n637 13.653
R1826 VDD.n644 VDD.n643 13.653
R1827 VDD.n643 VDD.n642 13.653
R1828 VDD.n648 VDD.n647 13.653
R1829 VDD.n647 VDD.n646 13.653
R1830 VDD.n652 VDD.n651 13.653
R1831 VDD.n651 VDD.n650 13.653
R1832 VDD.n678 VDD.n677 13.653
R1833 VDD.n677 VDD.n676 13.653
R1834 VDD.n682 VDD.n681 13.653
R1835 VDD.n681 VDD.n680 13.653
R1836 VDD.n686 VDD.n685 13.653
R1837 VDD.n685 VDD.n684 13.653
R1838 VDD.n691 VDD.n690 13.653
R1839 VDD.n690 VDD.n689 13.653
R1840 VDD.n698 VDD.n695 13.653
R1841 VDD.n695 VDD.n694 13.653
R1842 VDD.n703 VDD.n702 13.653
R1843 VDD.n702 VDD.n701 13.653
R1844 VDD.n708 VDD.n707 13.653
R1845 VDD.n707 VDD.n706 13.653
R1846 VDD.n715 VDD.n714 13.653
R1847 VDD.n714 VDD.n713 13.653
R1848 VDD.n720 VDD.n719 13.653
R1849 VDD.n719 VDD.n718 13.653
R1850 VDD.n725 VDD.n724 13.653
R1851 VDD.n724 VDD.n723 13.653
R1852 VDD.n729 VDD.n728 13.653
R1853 VDD.n728 VDD.n727 13.653
R1854 VDD.n733 VDD.n732 13.653
R1855 VDD.n732 VDD.n731 13.653
R1856 VDD.n759 VDD.n758 13.653
R1857 VDD.n758 VDD.n757 13.653
R1858 VDD.n763 VDD.n762 13.653
R1859 VDD.n762 VDD.n761 13.653
R1860 VDD.n767 VDD.n766 13.653
R1861 VDD.n766 VDD.n765 13.653
R1862 VDD.n772 VDD.n771 13.653
R1863 VDD.n771 VDD.n770 13.653
R1864 VDD.n779 VDD.n776 13.653
R1865 VDD.n776 VDD.n775 13.653
R1866 VDD.n784 VDD.n783 13.653
R1867 VDD.n783 VDD.n782 13.653
R1868 VDD.n789 VDD.n788 13.653
R1869 VDD.n788 VDD.n787 13.653
R1870 VDD.n796 VDD.n795 13.653
R1871 VDD.n795 VDD.n794 13.653
R1872 VDD.n801 VDD.n800 13.653
R1873 VDD.n800 VDD.n799 13.653
R1874 VDD.n806 VDD.n805 13.653
R1875 VDD.n805 VDD.n804 13.653
R1876 VDD.n810 VDD.n809 13.653
R1877 VDD.n809 VDD.n808 13.653
R1878 VDD.n836 VDD.n835 13.653
R1879 VDD.n835 VDD.n834 13.653
R1880 VDD.n1644 VDD.n1643 13.653
R1881 VDD.n1643 VDD.n1642 13.653
R1882 VDD.n1640 VDD.n1639 13.653
R1883 VDD.n1639 VDD.n1638 13.653
R1884 VDD.n1636 VDD.n1635 13.653
R1885 VDD.n1635 VDD.n1634 13.653
R1886 VDD.n1632 VDD.n1631 13.653
R1887 VDD.n1631 VDD.n1630 13.653
R1888 VDD.n1627 VDD.n1624 13.653
R1889 VDD.n1624 VDD.n1623 13.653
R1890 VDD.n1620 VDD.n1619 13.653
R1891 VDD.n1619 VDD.n1618 13.653
R1892 VDD.n1615 VDD.n1614 13.653
R1893 VDD.n1614 VDD.n1613 13.653
R1894 VDD.n1610 VDD.n1609 13.653
R1895 VDD.n1609 VDD.n1608 13.653
R1896 VDD.n1603 VDD.n1602 13.653
R1897 VDD.n1602 VDD.n1601 13.653
R1898 VDD.n1598 VDD.n1597 13.653
R1899 VDD.n1597 VDD.n1596 13.653
R1900 VDD.n1593 VDD.n1592 13.653
R1901 VDD.n1592 VDD.n1591 13.653
R1902 VDD.n1589 VDD.n1588 13.653
R1903 VDD.n1588 VDD.n1587 13.653
R1904 VDD.n1563 VDD.n1562 13.653
R1905 VDD.n1562 VDD.n1561 13.653
R1906 VDD.n1559 VDD.n1558 13.653
R1907 VDD.n1558 VDD.n1557 13.653
R1908 VDD.n1555 VDD.n1554 13.653
R1909 VDD.n1554 VDD.n1553 13.653
R1910 VDD.n1551 VDD.n1550 13.653
R1911 VDD.n1550 VDD.n1549 13.653
R1912 VDD.n1546 VDD.n1543 13.653
R1913 VDD.n1543 VDD.n1542 13.653
R1914 VDD.n1539 VDD.n1538 13.653
R1915 VDD.n1538 VDD.n1537 13.653
R1916 VDD.n1534 VDD.n1533 13.653
R1917 VDD.n1533 VDD.n1532 13.653
R1918 VDD.n1529 VDD.n1528 13.653
R1919 VDD.n1528 VDD.n1527 13.653
R1920 VDD.n1522 VDD.n1521 13.653
R1921 VDD.n1521 VDD.n1520 13.653
R1922 VDD.n1517 VDD.n1516 13.653
R1923 VDD.n1516 VDD.n1515 13.653
R1924 VDD.n1512 VDD.n1511 13.653
R1925 VDD.n1511 VDD.n1510 13.653
R1926 VDD.n1508 VDD.n1507 13.653
R1927 VDD.n1507 VDD.n1506 13.653
R1928 VDD.n1482 VDD.n1481 13.653
R1929 VDD.n1481 VDD.n1480 13.653
R1930 VDD.n1478 VDD.n1477 13.653
R1931 VDD.n1477 VDD.n1476 13.653
R1932 VDD.n1474 VDD.n1473 13.653
R1933 VDD.n1473 VDD.n1472 13.653
R1934 VDD.n1470 VDD.n1469 13.653
R1935 VDD.n1469 VDD.n1468 13.653
R1936 VDD.n1465 VDD.n1462 13.653
R1937 VDD.n1462 VDD.n1461 13.653
R1938 VDD.n1458 VDD.n1457 13.653
R1939 VDD.n1457 VDD.n1456 13.653
R1940 VDD.n1453 VDD.n1452 13.653
R1941 VDD.n1452 VDD.n1451 13.653
R1942 VDD.n1448 VDD.n1447 13.653
R1943 VDD.n1447 VDD.n1446 13.653
R1944 VDD.n1441 VDD.n1440 13.653
R1945 VDD.n1440 VDD.n1439 13.653
R1946 VDD.n1436 VDD.n1435 13.653
R1947 VDD.n1435 VDD.n1434 13.653
R1948 VDD.n1431 VDD.n1430 13.653
R1949 VDD.n1430 VDD.n1429 13.653
R1950 VDD.n1427 VDD.n1426 13.653
R1951 VDD.n1426 VDD.n1425 13.653
R1952 VDD.n1401 VDD.n1400 13.653
R1953 VDD.n1400 VDD.n1399 13.653
R1954 VDD.n1397 VDD.n1396 13.653
R1955 VDD.n1396 VDD.n1395 13.653
R1956 VDD.n1393 VDD.n1392 13.653
R1957 VDD.n1392 VDD.n1391 13.653
R1958 VDD.n1389 VDD.n1388 13.653
R1959 VDD.n1388 VDD.n1387 13.653
R1960 VDD.n1384 VDD.n1381 13.653
R1961 VDD.n1381 VDD.n1380 13.653
R1962 VDD.n1377 VDD.n1376 13.653
R1963 VDD.n1376 VDD.n1375 13.653
R1964 VDD.n1372 VDD.n1371 13.653
R1965 VDD.n1371 VDD.n1370 13.653
R1966 VDD.n1367 VDD.n1366 13.653
R1967 VDD.n1366 VDD.n1365 13.653
R1968 VDD.n1360 VDD.n1359 13.653
R1969 VDD.n1359 VDD.n1358 13.653
R1970 VDD.n1355 VDD.n1354 13.653
R1971 VDD.n1354 VDD.n1353 13.653
R1972 VDD.n1350 VDD.n1349 13.653
R1973 VDD.n1349 VDD.n1348 13.653
R1974 VDD.n1346 VDD.n1345 13.653
R1975 VDD.n1345 VDD.n1344 13.653
R1976 VDD.n1320 VDD.n1319 13.653
R1977 VDD.n1319 VDD.n1318 13.653
R1978 VDD.n1316 VDD.n1315 13.653
R1979 VDD.n1315 VDD.n1314 13.653
R1980 VDD.n1312 VDD.n1311 13.653
R1981 VDD.n1311 VDD.n1310 13.653
R1982 VDD.n1308 VDD.n1307 13.653
R1983 VDD.n1307 VDD.n1306 13.653
R1984 VDD.n1303 VDD.n1300 13.653
R1985 VDD.n1300 VDD.n1299 13.653
R1986 VDD.n1296 VDD.n1295 13.653
R1987 VDD.n1295 VDD.n1294 13.653
R1988 VDD.n1291 VDD.n1290 13.653
R1989 VDD.n1290 VDD.n1289 13.653
R1990 VDD.n1286 VDD.n1285 13.653
R1991 VDD.n1285 VDD.n1284 13.653
R1992 VDD.n1279 VDD.n1278 13.653
R1993 VDD.n1278 VDD.n1277 13.653
R1994 VDD.n1274 VDD.n1273 13.653
R1995 VDD.n1273 VDD.n1272 13.653
R1996 VDD.n1269 VDD.n1268 13.653
R1997 VDD.n1268 VDD.n1267 13.653
R1998 VDD.n1265 VDD.n1264 13.653
R1999 VDD.n1264 VDD.n1263 13.653
R2000 VDD.n1239 VDD.n1238 13.653
R2001 VDD.n1238 VDD.n1237 13.653
R2002 VDD.n1235 VDD.n1234 13.653
R2003 VDD.n1234 VDD.n1233 13.653
R2004 VDD.n1231 VDD.n1230 13.653
R2005 VDD.n1230 VDD.n1229 13.653
R2006 VDD.n1227 VDD.n1226 13.653
R2007 VDD.n1226 VDD.n1225 13.653
R2008 VDD.n1222 VDD.n1219 13.653
R2009 VDD.n1219 VDD.n1218 13.653
R2010 VDD.n1215 VDD.n1214 13.653
R2011 VDD.n1214 VDD.n1213 13.653
R2012 VDD.n1210 VDD.n1209 13.653
R2013 VDD.n1209 VDD.n1208 13.653
R2014 VDD.n1205 VDD.n1204 13.653
R2015 VDD.n1204 VDD.n1203 13.653
R2016 VDD.n1198 VDD.n1197 13.653
R2017 VDD.n1197 VDD.n1196 13.653
R2018 VDD.n1193 VDD.n1192 13.653
R2019 VDD.n1192 VDD.n1191 13.653
R2020 VDD.n1188 VDD.n1187 13.653
R2021 VDD.n1187 VDD.n1186 13.653
R2022 VDD.n1184 VDD.n1183 13.653
R2023 VDD.n1183 VDD.n1182 13.653
R2024 VDD.n1158 VDD.n1157 13.653
R2025 VDD.n1157 VDD.n1156 13.653
R2026 VDD.n1154 VDD.n1153 13.653
R2027 VDD.n1153 VDD.n1152 13.653
R2028 VDD.n1150 VDD.n1149 13.653
R2029 VDD.n1149 VDD.n1148 13.653
R2030 VDD.n1146 VDD.n1145 13.653
R2031 VDD.n1145 VDD.n1144 13.653
R2032 VDD.n1141 VDD.n1138 13.653
R2033 VDD.n1138 VDD.n1137 13.653
R2034 VDD.n1134 VDD.n1133 13.653
R2035 VDD.n1133 VDD.n1132 13.653
R2036 VDD.n1129 VDD.n1128 13.653
R2037 VDD.n1128 VDD.n1127 13.653
R2038 VDD.n1124 VDD.n1123 13.653
R2039 VDD.n1123 VDD.n1122 13.653
R2040 VDD.n1117 VDD.n1116 13.653
R2041 VDD.n1116 VDD.n1115 13.653
R2042 VDD.n1112 VDD.n1111 13.653
R2043 VDD.n1111 VDD.n1110 13.653
R2044 VDD.n1107 VDD.n1106 13.653
R2045 VDD.n1106 VDD.n1105 13.653
R2046 VDD.n1103 VDD.n1102 13.653
R2047 VDD.n1102 VDD.n1101 13.653
R2048 VDD.n1077 VDD.n1076 13.653
R2049 VDD.n1076 VDD.n1075 13.653
R2050 VDD.n1073 VDD.n1072 13.653
R2051 VDD.n1072 VDD.n1071 13.653
R2052 VDD.n1069 VDD.n1068 13.653
R2053 VDD.n1068 VDD.n1067 13.653
R2054 VDD.n1065 VDD.n1064 13.653
R2055 VDD.n1064 VDD.n1063 13.653
R2056 VDD.n1060 VDD.n1057 13.653
R2057 VDD.n1057 VDD.n1056 13.653
R2058 VDD.n1053 VDD.n1052 13.653
R2059 VDD.n1052 VDD.n1051 13.653
R2060 VDD.n1048 VDD.n1047 13.653
R2061 VDD.n1047 VDD.n1046 13.653
R2062 VDD.n1043 VDD.n1042 13.653
R2063 VDD.n1042 VDD.n1041 13.653
R2064 VDD.n1036 VDD.n1035 13.653
R2065 VDD.n1035 VDD.n1034 13.653
R2066 VDD.n1031 VDD.n1030 13.653
R2067 VDD.n1030 VDD.n1029 13.653
R2068 VDD.n1026 VDD.n1025 13.653
R2069 VDD.n1025 VDD.n1024 13.653
R2070 VDD.n1022 VDD.n1021 13.653
R2071 VDD.n1021 VDD.n1020 13.653
R2072 VDD.n996 VDD.n995 13.653
R2073 VDD.n995 VDD.n994 13.653
R2074 VDD.n992 VDD.n991 13.653
R2075 VDD.n991 VDD.n990 13.653
R2076 VDD.n988 VDD.n987 13.653
R2077 VDD.n987 VDD.n986 13.653
R2078 VDD.n984 VDD.n983 13.653
R2079 VDD.n983 VDD.n982 13.653
R2080 VDD.n979 VDD.n976 13.653
R2081 VDD.n976 VDD.n975 13.653
R2082 VDD.n972 VDD.n971 13.653
R2083 VDD.n971 VDD.n970 13.653
R2084 VDD.n967 VDD.n966 13.653
R2085 VDD.n966 VDD.n965 13.653
R2086 VDD.n962 VDD.n961 13.653
R2087 VDD.n961 VDD.n960 13.653
R2088 VDD.n955 VDD.n954 13.653
R2089 VDD.n954 VDD.n953 13.653
R2090 VDD.n950 VDD.n949 13.653
R2091 VDD.n949 VDD.n948 13.653
R2092 VDD.n945 VDD.n944 13.653
R2093 VDD.n944 VDD.n943 13.653
R2094 VDD.n941 VDD.n940 13.653
R2095 VDD.n940 VDD.n939 13.653
R2096 VDD.n914 VDD.n913 13.653
R2097 VDD.n913 VDD.n912 13.653
R2098 VDD.n910 VDD.n909 13.653
R2099 VDD.n909 VDD.n908 13.653
R2100 VDD.n906 VDD.n905 13.653
R2101 VDD.n905 VDD.n904 13.653
R2102 VDD.n902 VDD.n901 13.653
R2103 VDD.n901 VDD.n900 13.653
R2104 VDD.n897 VDD.n894 13.653
R2105 VDD.n894 VDD.n893 13.653
R2106 VDD.n890 VDD.n889 13.653
R2107 VDD.n889 VDD.n888 13.653
R2108 VDD.n885 VDD.n884 13.653
R2109 VDD.n884 VDD.n883 13.653
R2110 VDD.n880 VDD.n879 13.653
R2111 VDD.n879 VDD.n878 13.653
R2112 VDD.n873 VDD.n872 13.653
R2113 VDD.n872 VDD.n871 13.653
R2114 VDD.n868 VDD.n867 13.653
R2115 VDD.n867 VDD.n866 13.653
R2116 VDD.n863 VDD.n862 13.653
R2117 VDD.n862 VDD.n861 13.653
R2118 VDD.n859 VDD.n858 13.653
R2119 VDD.n858 VDD.n857 13.653
R2120 VDD.n4 VDD.n2 12.915
R2121 VDD.n4 VDD.n3 12.66
R2122 VDD.n13 VDD.n12 12.343
R2123 VDD.n11 VDD.n10 12.343
R2124 VDD.n7 VDD.n6 12.343
R2125 VDD.n215 VDD.n214 9.152
R2126 VDD.n296 VDD.n295 9.152
R2127 VDD.n377 VDD.n376 9.152
R2128 VDD.n458 VDD.n457 9.152
R2129 VDD.n539 VDD.n538 9.152
R2130 VDD.n620 VDD.n619 9.152
R2131 VDD.n701 VDD.n700 9.152
R2132 VDD.n782 VDD.n781 9.152
R2133 VDD.n1618 VDD.n1617 9.152
R2134 VDD.n1537 VDD.n1536 9.152
R2135 VDD.n1456 VDD.n1455 9.152
R2136 VDD.n1375 VDD.n1374 9.152
R2137 VDD.n1294 VDD.n1293 9.152
R2138 VDD.n1213 VDD.n1212 9.152
R2139 VDD.n1132 VDD.n1131 9.152
R2140 VDD.n1051 VDD.n1050 9.152
R2141 VDD.n970 VDD.n969 9.152
R2142 VDD.n888 VDD.n887 9.152
R2143 VDD.n147 VDD.n144 8.658
R2144 VDD.n1018 VDD.n1017 7.674
R2145 VDD.n1099 VDD.n1098 7.674
R2146 VDD.n1180 VDD.n1179 7.674
R2147 VDD.n1261 VDD.n1260 7.674
R2148 VDD.n1342 VDD.n1341 7.674
R2149 VDD.n1423 VDD.n1422 7.674
R2150 VDD.n1504 VDD.n1503 7.674
R2151 VDD.n1585 VDD.n1584 7.674
R2152 VDD.n832 VDD.n831 7.674
R2153 VDD.n755 VDD.n754 7.674
R2154 VDD.n674 VDD.n673 7.674
R2155 VDD.n593 VDD.n592 7.674
R2156 VDD.n512 VDD.n511 7.674
R2157 VDD.n431 VDD.n430 7.674
R2158 VDD.n350 VDD.n349 7.674
R2159 VDD.n269 VDD.n268 7.674
R2160 VDD.n188 VDD.n187 7.674
R2161 VDD.n127 VDD.n126 7.674
R2162 VDD.n73 VDD.n72 7.674
R2163 VDD.n937 VDD.n936 7.674
R2164 VDD.n67 VDD.n66 7.5
R2165 VDD.n61 VDD.n60 7.5
R2166 VDD.n63 VDD.n62 7.5
R2167 VDD.n58 VDD.n57 7.5
R2168 VDD.n72 VDD.n71 7.5
R2169 VDD.n121 VDD.n120 7.5
R2170 VDD.n115 VDD.n114 7.5
R2171 VDD.n117 VDD.n116 7.5
R2172 VDD.n123 VDD.n113 7.5
R2173 VDD.n123 VDD.n111 7.5
R2174 VDD.n126 VDD.n125 7.5
R2175 VDD.n182 VDD.n181 7.5
R2176 VDD.n176 VDD.n175 7.5
R2177 VDD.n178 VDD.n177 7.5
R2178 VDD.n184 VDD.n174 7.5
R2179 VDD.n184 VDD.n172 7.5
R2180 VDD.n187 VDD.n186 7.5
R2181 VDD.n263 VDD.n262 7.5
R2182 VDD.n257 VDD.n256 7.5
R2183 VDD.n259 VDD.n258 7.5
R2184 VDD.n265 VDD.n255 7.5
R2185 VDD.n265 VDD.n253 7.5
R2186 VDD.n268 VDD.n267 7.5
R2187 VDD.n344 VDD.n343 7.5
R2188 VDD.n338 VDD.n337 7.5
R2189 VDD.n340 VDD.n339 7.5
R2190 VDD.n346 VDD.n336 7.5
R2191 VDD.n346 VDD.n334 7.5
R2192 VDD.n349 VDD.n348 7.5
R2193 VDD.n425 VDD.n424 7.5
R2194 VDD.n419 VDD.n418 7.5
R2195 VDD.n421 VDD.n420 7.5
R2196 VDD.n427 VDD.n417 7.5
R2197 VDD.n427 VDD.n415 7.5
R2198 VDD.n430 VDD.n429 7.5
R2199 VDD.n506 VDD.n505 7.5
R2200 VDD.n500 VDD.n499 7.5
R2201 VDD.n502 VDD.n501 7.5
R2202 VDD.n508 VDD.n498 7.5
R2203 VDD.n508 VDD.n496 7.5
R2204 VDD.n511 VDD.n510 7.5
R2205 VDD.n587 VDD.n586 7.5
R2206 VDD.n581 VDD.n580 7.5
R2207 VDD.n583 VDD.n582 7.5
R2208 VDD.n589 VDD.n579 7.5
R2209 VDD.n589 VDD.n577 7.5
R2210 VDD.n592 VDD.n591 7.5
R2211 VDD.n668 VDD.n667 7.5
R2212 VDD.n662 VDD.n661 7.5
R2213 VDD.n664 VDD.n663 7.5
R2214 VDD.n670 VDD.n660 7.5
R2215 VDD.n670 VDD.n658 7.5
R2216 VDD.n673 VDD.n672 7.5
R2217 VDD.n749 VDD.n748 7.5
R2218 VDD.n743 VDD.n742 7.5
R2219 VDD.n745 VDD.n744 7.5
R2220 VDD.n751 VDD.n741 7.5
R2221 VDD.n751 VDD.n739 7.5
R2222 VDD.n754 VDD.n753 7.5
R2223 VDD.n826 VDD.n825 7.5
R2224 VDD.n820 VDD.n819 7.5
R2225 VDD.n822 VDD.n821 7.5
R2226 VDD.n828 VDD.n818 7.5
R2227 VDD.n828 VDD.n816 7.5
R2228 VDD.n831 VDD.n830 7.5
R2229 VDD.n1579 VDD.n1578 7.5
R2230 VDD.n1573 VDD.n1572 7.5
R2231 VDD.n1575 VDD.n1574 7.5
R2232 VDD.n1581 VDD.n1571 7.5
R2233 VDD.n1581 VDD.n1569 7.5
R2234 VDD.n1584 VDD.n1583 7.5
R2235 VDD.n1498 VDD.n1497 7.5
R2236 VDD.n1492 VDD.n1491 7.5
R2237 VDD.n1494 VDD.n1493 7.5
R2238 VDD.n1500 VDD.n1490 7.5
R2239 VDD.n1500 VDD.n1488 7.5
R2240 VDD.n1503 VDD.n1502 7.5
R2241 VDD.n1417 VDD.n1416 7.5
R2242 VDD.n1411 VDD.n1410 7.5
R2243 VDD.n1413 VDD.n1412 7.5
R2244 VDD.n1419 VDD.n1409 7.5
R2245 VDD.n1419 VDD.n1407 7.5
R2246 VDD.n1422 VDD.n1421 7.5
R2247 VDD.n1336 VDD.n1335 7.5
R2248 VDD.n1330 VDD.n1329 7.5
R2249 VDD.n1332 VDD.n1331 7.5
R2250 VDD.n1338 VDD.n1328 7.5
R2251 VDD.n1338 VDD.n1326 7.5
R2252 VDD.n1341 VDD.n1340 7.5
R2253 VDD.n1255 VDD.n1254 7.5
R2254 VDD.n1249 VDD.n1248 7.5
R2255 VDD.n1251 VDD.n1250 7.5
R2256 VDD.n1257 VDD.n1247 7.5
R2257 VDD.n1257 VDD.n1245 7.5
R2258 VDD.n1260 VDD.n1259 7.5
R2259 VDD.n1174 VDD.n1173 7.5
R2260 VDD.n1168 VDD.n1167 7.5
R2261 VDD.n1170 VDD.n1169 7.5
R2262 VDD.n1176 VDD.n1166 7.5
R2263 VDD.n1176 VDD.n1164 7.5
R2264 VDD.n1179 VDD.n1178 7.5
R2265 VDD.n1093 VDD.n1092 7.5
R2266 VDD.n1087 VDD.n1086 7.5
R2267 VDD.n1089 VDD.n1088 7.5
R2268 VDD.n1095 VDD.n1085 7.5
R2269 VDD.n1095 VDD.n1083 7.5
R2270 VDD.n1098 VDD.n1097 7.5
R2271 VDD.n1012 VDD.n1011 7.5
R2272 VDD.n1006 VDD.n1005 7.5
R2273 VDD.n1008 VDD.n1007 7.5
R2274 VDD.n1014 VDD.n1004 7.5
R2275 VDD.n1014 VDD.n1002 7.5
R2276 VDD.n1017 VDD.n1016 7.5
R2277 VDD.n921 VDD.n920 7.5
R2278 VDD.n924 VDD.n923 7.5
R2279 VDD.n926 VDD.n925 7.5
R2280 VDD.n929 VDD.n928 7.5
R2281 VDD.n936 VDD.n935 7.5
R2282 VDD.n851 VDD.n850 7.5
R2283 VDD.n845 VDD.n844 7.5
R2284 VDD.n847 VDD.n846 7.5
R2285 VDD.n853 VDD.n843 7.5
R2286 VDD.n853 VDD.n841 7.5
R2287 VDD.n856 VDD.n855 7.5
R2288 VDD.n20 VDD.n16 7.5
R2289 VDD.n2 VDD.n1 7.5
R2290 VDD.n6 VDD.n5 7.5
R2291 VDD.n10 VDD.n9 7.5
R2292 VDD.n19 VDD.n18 7.5
R2293 VDD.n14 VDD.n0 7.5
R2294 VDD.n59 VDD.n56 6.772
R2295 VDD.n70 VDD.n54 6.772
R2296 VDD.n68 VDD.n65 6.772
R2297 VDD.n64 VDD.n61 6.772
R2298 VDD.n124 VDD.n109 6.772
R2299 VDD.n122 VDD.n119 6.772
R2300 VDD.n118 VDD.n115 6.772
R2301 VDD.n185 VDD.n170 6.772
R2302 VDD.n183 VDD.n180 6.772
R2303 VDD.n179 VDD.n176 6.772
R2304 VDD.n266 VDD.n251 6.772
R2305 VDD.n264 VDD.n261 6.772
R2306 VDD.n260 VDD.n257 6.772
R2307 VDD.n347 VDD.n332 6.772
R2308 VDD.n345 VDD.n342 6.772
R2309 VDD.n341 VDD.n338 6.772
R2310 VDD.n428 VDD.n413 6.772
R2311 VDD.n426 VDD.n423 6.772
R2312 VDD.n422 VDD.n419 6.772
R2313 VDD.n509 VDD.n494 6.772
R2314 VDD.n507 VDD.n504 6.772
R2315 VDD.n503 VDD.n500 6.772
R2316 VDD.n590 VDD.n575 6.772
R2317 VDD.n588 VDD.n585 6.772
R2318 VDD.n584 VDD.n581 6.772
R2319 VDD.n671 VDD.n656 6.772
R2320 VDD.n669 VDD.n666 6.772
R2321 VDD.n665 VDD.n662 6.772
R2322 VDD.n752 VDD.n737 6.772
R2323 VDD.n750 VDD.n747 6.772
R2324 VDD.n746 VDD.n743 6.772
R2325 VDD.n829 VDD.n814 6.772
R2326 VDD.n827 VDD.n824 6.772
R2327 VDD.n823 VDD.n820 6.772
R2328 VDD.n1582 VDD.n1567 6.772
R2329 VDD.n1580 VDD.n1577 6.772
R2330 VDD.n1576 VDD.n1573 6.772
R2331 VDD.n1501 VDD.n1486 6.772
R2332 VDD.n1499 VDD.n1496 6.772
R2333 VDD.n1495 VDD.n1492 6.772
R2334 VDD.n1420 VDD.n1405 6.772
R2335 VDD.n1418 VDD.n1415 6.772
R2336 VDD.n1414 VDD.n1411 6.772
R2337 VDD.n1339 VDD.n1324 6.772
R2338 VDD.n1337 VDD.n1334 6.772
R2339 VDD.n1333 VDD.n1330 6.772
R2340 VDD.n1258 VDD.n1243 6.772
R2341 VDD.n1256 VDD.n1253 6.772
R2342 VDD.n1252 VDD.n1249 6.772
R2343 VDD.n1177 VDD.n1162 6.772
R2344 VDD.n1175 VDD.n1172 6.772
R2345 VDD.n1171 VDD.n1168 6.772
R2346 VDD.n1096 VDD.n1081 6.772
R2347 VDD.n1094 VDD.n1091 6.772
R2348 VDD.n1090 VDD.n1087 6.772
R2349 VDD.n1015 VDD.n1000 6.772
R2350 VDD.n1013 VDD.n1010 6.772
R2351 VDD.n1009 VDD.n1006 6.772
R2352 VDD.n854 VDD.n840 6.772
R2353 VDD.n852 VDD.n849 6.772
R2354 VDD.n848 VDD.n845 6.772
R2355 VDD.n59 VDD.n58 6.772
R2356 VDD.n64 VDD.n63 6.772
R2357 VDD.n68 VDD.n67 6.772
R2358 VDD.n71 VDD.n70 6.772
R2359 VDD.n118 VDD.n117 6.772
R2360 VDD.n122 VDD.n121 6.772
R2361 VDD.n125 VDD.n124 6.772
R2362 VDD.n179 VDD.n178 6.772
R2363 VDD.n183 VDD.n182 6.772
R2364 VDD.n186 VDD.n185 6.772
R2365 VDD.n260 VDD.n259 6.772
R2366 VDD.n264 VDD.n263 6.772
R2367 VDD.n267 VDD.n266 6.772
R2368 VDD.n341 VDD.n340 6.772
R2369 VDD.n345 VDD.n344 6.772
R2370 VDD.n348 VDD.n347 6.772
R2371 VDD.n422 VDD.n421 6.772
R2372 VDD.n426 VDD.n425 6.772
R2373 VDD.n429 VDD.n428 6.772
R2374 VDD.n503 VDD.n502 6.772
R2375 VDD.n507 VDD.n506 6.772
R2376 VDD.n510 VDD.n509 6.772
R2377 VDD.n584 VDD.n583 6.772
R2378 VDD.n588 VDD.n587 6.772
R2379 VDD.n591 VDD.n590 6.772
R2380 VDD.n665 VDD.n664 6.772
R2381 VDD.n669 VDD.n668 6.772
R2382 VDD.n672 VDD.n671 6.772
R2383 VDD.n746 VDD.n745 6.772
R2384 VDD.n750 VDD.n749 6.772
R2385 VDD.n753 VDD.n752 6.772
R2386 VDD.n823 VDD.n822 6.772
R2387 VDD.n827 VDD.n826 6.772
R2388 VDD.n830 VDD.n829 6.772
R2389 VDD.n1576 VDD.n1575 6.772
R2390 VDD.n1580 VDD.n1579 6.772
R2391 VDD.n1583 VDD.n1582 6.772
R2392 VDD.n1495 VDD.n1494 6.772
R2393 VDD.n1499 VDD.n1498 6.772
R2394 VDD.n1502 VDD.n1501 6.772
R2395 VDD.n1414 VDD.n1413 6.772
R2396 VDD.n1418 VDD.n1417 6.772
R2397 VDD.n1421 VDD.n1420 6.772
R2398 VDD.n1333 VDD.n1332 6.772
R2399 VDD.n1337 VDD.n1336 6.772
R2400 VDD.n1340 VDD.n1339 6.772
R2401 VDD.n1252 VDD.n1251 6.772
R2402 VDD.n1256 VDD.n1255 6.772
R2403 VDD.n1259 VDD.n1258 6.772
R2404 VDD.n1171 VDD.n1170 6.772
R2405 VDD.n1175 VDD.n1174 6.772
R2406 VDD.n1178 VDD.n1177 6.772
R2407 VDD.n1090 VDD.n1089 6.772
R2408 VDD.n1094 VDD.n1093 6.772
R2409 VDD.n1097 VDD.n1096 6.772
R2410 VDD.n1009 VDD.n1008 6.772
R2411 VDD.n1013 VDD.n1012 6.772
R2412 VDD.n1016 VDD.n1015 6.772
R2413 VDD.n848 VDD.n847 6.772
R2414 VDD.n852 VDD.n851 6.772
R2415 VDD.n855 VDD.n854 6.772
R2416 VDD.n935 VDD.n934 6.772
R2417 VDD.n922 VDD.n919 6.772
R2418 VDD.n927 VDD.n924 6.772
R2419 VDD.n932 VDD.n929 6.772
R2420 VDD.n932 VDD.n931 6.772
R2421 VDD.n927 VDD.n926 6.772
R2422 VDD.n922 VDD.n921 6.772
R2423 VDD.n934 VDD.n918 6.772
R2424 VDD.n229 VDD.n225 6.69
R2425 VDD.n310 VDD.n306 6.69
R2426 VDD.n391 VDD.n387 6.69
R2427 VDD.n472 VDD.n468 6.69
R2428 VDD.n553 VDD.n549 6.69
R2429 VDD.n634 VDD.n630 6.69
R2430 VDD.n715 VDD.n711 6.69
R2431 VDD.n796 VDD.n792 6.69
R2432 VDD.n1610 VDD.n1606 6.69
R2433 VDD.n1529 VDD.n1525 6.69
R2434 VDD.n1448 VDD.n1444 6.69
R2435 VDD.n1367 VDD.n1363 6.69
R2436 VDD.n1286 VDD.n1282 6.69
R2437 VDD.n1205 VDD.n1201 6.69
R2438 VDD.n1124 VDD.n1120 6.69
R2439 VDD.n1043 VDD.n1039 6.69
R2440 VDD.n962 VDD.n958 6.69
R2441 VDD.n880 VDD.n876 6.69
R2442 VDD.n33 VDD.n23 6.487
R2443 VDD.n33 VDD.n32 6.475
R2444 VDD.n16 VDD.n15 6.458
R2445 VDD.n212 VDD.n211 6.296
R2446 VDD.n293 VDD.n292 6.296
R2447 VDD.n374 VDD.n373 6.296
R2448 VDD.n455 VDD.n454 6.296
R2449 VDD.n536 VDD.n535 6.296
R2450 VDD.n617 VDD.n616 6.296
R2451 VDD.n698 VDD.n697 6.296
R2452 VDD.n779 VDD.n778 6.296
R2453 VDD.n1627 VDD.n1626 6.296
R2454 VDD.n1546 VDD.n1545 6.296
R2455 VDD.n1465 VDD.n1464 6.296
R2456 VDD.n1384 VDD.n1383 6.296
R2457 VDD.n1303 VDD.n1302 6.296
R2458 VDD.n1222 VDD.n1221 6.296
R2459 VDD.n1141 VDD.n1140 6.296
R2460 VDD.n1060 VDD.n1059 6.296
R2461 VDD.n979 VDD.n978 6.296
R2462 VDD.n897 VDD.n896 6.296
R2463 VDD.n113 VDD.n112 6.202
R2464 VDD.n174 VDD.n173 6.202
R2465 VDD.n255 VDD.n254 6.202
R2466 VDD.n336 VDD.n335 6.202
R2467 VDD.n417 VDD.n416 6.202
R2468 VDD.n498 VDD.n497 6.202
R2469 VDD.n579 VDD.n578 6.202
R2470 VDD.n660 VDD.n659 6.202
R2471 VDD.n741 VDD.n740 6.202
R2472 VDD.n818 VDD.n817 6.202
R2473 VDD.n1571 VDD.n1570 6.202
R2474 VDD.n1490 VDD.n1489 6.202
R2475 VDD.n1409 VDD.n1408 6.202
R2476 VDD.n1328 VDD.n1327 6.202
R2477 VDD.n1247 VDD.n1246 6.202
R2478 VDD.n1166 VDD.n1165 6.202
R2479 VDD.n1085 VDD.n1084 6.202
R2480 VDD.n1004 VDD.n1003 6.202
R2481 VDD.n843 VDD.n842 6.202
R2482 VDD.n150 VDD.n149 4.576
R2483 VDD.n162 VDD.n159 2.754
R2484 VDD.n136 VDD.n133 2.361
R2485 VDD.n14 VDD.n7 1.329
R2486 VDD.n14 VDD.n8 1.329
R2487 VDD.n14 VDD.n11 1.329
R2488 VDD.n14 VDD.n13 1.329
R2489 VDD.n15 VDD.n14 0.696
R2490 VDD.n14 VDD.n4 0.696
R2491 VDD.n239 VDD.n236 0.393
R2492 VDD.n320 VDD.n317 0.393
R2493 VDD.n401 VDD.n398 0.393
R2494 VDD.n482 VDD.n479 0.393
R2495 VDD.n563 VDD.n560 0.393
R2496 VDD.n644 VDD.n641 0.393
R2497 VDD.n725 VDD.n722 0.393
R2498 VDD.n806 VDD.n803 0.393
R2499 VDD.n1598 VDD.n1595 0.393
R2500 VDD.n1517 VDD.n1514 0.393
R2501 VDD.n1436 VDD.n1433 0.393
R2502 VDD.n1355 VDD.n1352 0.393
R2503 VDD.n1274 VDD.n1271 0.393
R2504 VDD.n1193 VDD.n1190 0.393
R2505 VDD.n1112 VDD.n1109 0.393
R2506 VDD.n1031 VDD.n1028 0.393
R2507 VDD.n950 VDD.n947 0.393
R2508 VDD.n868 VDD.n865 0.393
R2509 VDD.n69 VDD.n68 0.365
R2510 VDD.n69 VDD.n64 0.365
R2511 VDD.n69 VDD.n59 0.365
R2512 VDD.n70 VDD.n69 0.365
R2513 VDD.n123 VDD.n122 0.365
R2514 VDD.n123 VDD.n118 0.365
R2515 VDD.n124 VDD.n123 0.365
R2516 VDD.n184 VDD.n183 0.365
R2517 VDD.n184 VDD.n179 0.365
R2518 VDD.n185 VDD.n184 0.365
R2519 VDD.n265 VDD.n264 0.365
R2520 VDD.n265 VDD.n260 0.365
R2521 VDD.n266 VDD.n265 0.365
R2522 VDD.n346 VDD.n345 0.365
R2523 VDD.n346 VDD.n341 0.365
R2524 VDD.n347 VDD.n346 0.365
R2525 VDD.n427 VDD.n426 0.365
R2526 VDD.n427 VDD.n422 0.365
R2527 VDD.n428 VDD.n427 0.365
R2528 VDD.n508 VDD.n507 0.365
R2529 VDD.n508 VDD.n503 0.365
R2530 VDD.n509 VDD.n508 0.365
R2531 VDD.n589 VDD.n588 0.365
R2532 VDD.n589 VDD.n584 0.365
R2533 VDD.n590 VDD.n589 0.365
R2534 VDD.n670 VDD.n669 0.365
R2535 VDD.n670 VDD.n665 0.365
R2536 VDD.n671 VDD.n670 0.365
R2537 VDD.n751 VDD.n750 0.365
R2538 VDD.n751 VDD.n746 0.365
R2539 VDD.n752 VDD.n751 0.365
R2540 VDD.n828 VDD.n827 0.365
R2541 VDD.n828 VDD.n823 0.365
R2542 VDD.n829 VDD.n828 0.365
R2543 VDD.n1581 VDD.n1580 0.365
R2544 VDD.n1581 VDD.n1576 0.365
R2545 VDD.n1582 VDD.n1581 0.365
R2546 VDD.n1500 VDD.n1499 0.365
R2547 VDD.n1500 VDD.n1495 0.365
R2548 VDD.n1501 VDD.n1500 0.365
R2549 VDD.n1419 VDD.n1418 0.365
R2550 VDD.n1419 VDD.n1414 0.365
R2551 VDD.n1420 VDD.n1419 0.365
R2552 VDD.n1338 VDD.n1337 0.365
R2553 VDD.n1338 VDD.n1333 0.365
R2554 VDD.n1339 VDD.n1338 0.365
R2555 VDD.n1257 VDD.n1256 0.365
R2556 VDD.n1257 VDD.n1252 0.365
R2557 VDD.n1258 VDD.n1257 0.365
R2558 VDD.n1176 VDD.n1175 0.365
R2559 VDD.n1176 VDD.n1171 0.365
R2560 VDD.n1177 VDD.n1176 0.365
R2561 VDD.n1095 VDD.n1094 0.365
R2562 VDD.n1095 VDD.n1090 0.365
R2563 VDD.n1096 VDD.n1095 0.365
R2564 VDD.n1014 VDD.n1013 0.365
R2565 VDD.n1014 VDD.n1009 0.365
R2566 VDD.n1015 VDD.n1014 0.365
R2567 VDD.n853 VDD.n852 0.365
R2568 VDD.n853 VDD.n848 0.365
R2569 VDD.n854 VDD.n853 0.365
R2570 VDD.n933 VDD.n932 0.365
R2571 VDD.n933 VDD.n927 0.365
R2572 VDD.n933 VDD.n922 0.365
R2573 VDD.n934 VDD.n933 0.365
R2574 VDD.n78 VDD.n51 0.29
R2575 VDD.n132 VDD.n106 0.29
R2576 VDD.n193 VDD.n167 0.29
R2577 VDD.n274 VDD.n248 0.29
R2578 VDD.n355 VDD.n329 0.29
R2579 VDD.n436 VDD.n410 0.29
R2580 VDD.n517 VDD.n491 0.29
R2581 VDD.n598 VDD.n572 0.29
R2582 VDD.n679 VDD.n653 0.29
R2583 VDD.n760 VDD.n734 0.29
R2584 VDD.n1590 VDD.n1564 0.29
R2585 VDD.n1509 VDD.n1483 0.29
R2586 VDD.n1428 VDD.n1402 0.29
R2587 VDD.n1347 VDD.n1321 0.29
R2588 VDD.n1266 VDD.n1240 0.29
R2589 VDD.n1185 VDD.n1159 0.29
R2590 VDD.n1104 VDD.n1078 0.29
R2591 VDD.n1023 VDD.n997 0.29
R2592 VDD.n942 VDD.n915 0.29
R2593 VDD VDD.n1645 0.219
R2594 VDD.n860 VDD 0.207
R2595 VDD.n223 VDD.n218 0.197
R2596 VDD.n304 VDD.n299 0.197
R2597 VDD.n385 VDD.n380 0.197
R2598 VDD.n466 VDD.n461 0.197
R2599 VDD.n547 VDD.n542 0.197
R2600 VDD.n628 VDD.n623 0.197
R2601 VDD.n709 VDD.n704 0.197
R2602 VDD.n790 VDD.n785 0.197
R2603 VDD.n1621 VDD.n1616 0.197
R2604 VDD.n1540 VDD.n1535 0.197
R2605 VDD.n1459 VDD.n1454 0.197
R2606 VDD.n1378 VDD.n1373 0.197
R2607 VDD.n1297 VDD.n1292 0.197
R2608 VDD.n1216 VDD.n1211 0.197
R2609 VDD.n1135 VDD.n1130 0.197
R2610 VDD.n1054 VDD.n1049 0.197
R2611 VDD.n973 VDD.n968 0.197
R2612 VDD.n891 VDD.n886 0.197
R2613 VDD.n39 VDD.n35 0.181
R2614 VDD.n94 VDD.n90 0.181
R2615 VDD.n153 VDD.n148 0.181
R2616 VDD.n35 VDD.n34 0.145
R2617 VDD.n43 VDD.n39 0.145
R2618 VDD.n47 VDD.n43 0.145
R2619 VDD.n51 VDD.n47 0.145
R2620 VDD.n82 VDD.n78 0.145
R2621 VDD.n86 VDD.n82 0.145
R2622 VDD.n90 VDD.n86 0.145
R2623 VDD.n98 VDD.n94 0.145
R2624 VDD.n102 VDD.n98 0.145
R2625 VDD.n106 VDD.n102 0.145
R2626 VDD.n137 VDD.n132 0.145
R2627 VDD.n142 VDD.n137 0.145
R2628 VDD.n148 VDD.n142 0.145
R2629 VDD.n158 VDD.n153 0.145
R2630 VDD.n163 VDD.n158 0.145
R2631 VDD.n167 VDD.n163 0.145
R2632 VDD.n197 VDD.n193 0.145
R2633 VDD.n201 VDD.n197 0.145
R2634 VDD.n206 VDD.n201 0.145
R2635 VDD.n213 VDD.n206 0.145
R2636 VDD.n218 VDD.n213 0.145
R2637 VDD.n230 VDD.n223 0.145
R2638 VDD.n235 VDD.n230 0.145
R2639 VDD.n240 VDD.n235 0.145
R2640 VDD.n244 VDD.n240 0.145
R2641 VDD.n248 VDD.n244 0.145
R2642 VDD.n278 VDD.n274 0.145
R2643 VDD.n282 VDD.n278 0.145
R2644 VDD.n287 VDD.n282 0.145
R2645 VDD.n294 VDD.n287 0.145
R2646 VDD.n299 VDD.n294 0.145
R2647 VDD.n311 VDD.n304 0.145
R2648 VDD.n316 VDD.n311 0.145
R2649 VDD.n321 VDD.n316 0.145
R2650 VDD.n325 VDD.n321 0.145
R2651 VDD.n329 VDD.n325 0.145
R2652 VDD.n359 VDD.n355 0.145
R2653 VDD.n363 VDD.n359 0.145
R2654 VDD.n368 VDD.n363 0.145
R2655 VDD.n375 VDD.n368 0.145
R2656 VDD.n380 VDD.n375 0.145
R2657 VDD.n392 VDD.n385 0.145
R2658 VDD.n397 VDD.n392 0.145
R2659 VDD.n402 VDD.n397 0.145
R2660 VDD.n406 VDD.n402 0.145
R2661 VDD.n410 VDD.n406 0.145
R2662 VDD.n440 VDD.n436 0.145
R2663 VDD.n444 VDD.n440 0.145
R2664 VDD.n449 VDD.n444 0.145
R2665 VDD.n456 VDD.n449 0.145
R2666 VDD.n461 VDD.n456 0.145
R2667 VDD.n473 VDD.n466 0.145
R2668 VDD.n478 VDD.n473 0.145
R2669 VDD.n483 VDD.n478 0.145
R2670 VDD.n487 VDD.n483 0.145
R2671 VDD.n491 VDD.n487 0.145
R2672 VDD.n521 VDD.n517 0.145
R2673 VDD.n525 VDD.n521 0.145
R2674 VDD.n530 VDD.n525 0.145
R2675 VDD.n537 VDD.n530 0.145
R2676 VDD.n542 VDD.n537 0.145
R2677 VDD.n554 VDD.n547 0.145
R2678 VDD.n559 VDD.n554 0.145
R2679 VDD.n564 VDD.n559 0.145
R2680 VDD.n568 VDD.n564 0.145
R2681 VDD.n572 VDD.n568 0.145
R2682 VDD.n602 VDD.n598 0.145
R2683 VDD.n606 VDD.n602 0.145
R2684 VDD.n611 VDD.n606 0.145
R2685 VDD.n618 VDD.n611 0.145
R2686 VDD.n623 VDD.n618 0.145
R2687 VDD.n635 VDD.n628 0.145
R2688 VDD.n640 VDD.n635 0.145
R2689 VDD.n645 VDD.n640 0.145
R2690 VDD.n649 VDD.n645 0.145
R2691 VDD.n653 VDD.n649 0.145
R2692 VDD.n683 VDD.n679 0.145
R2693 VDD.n687 VDD.n683 0.145
R2694 VDD.n692 VDD.n687 0.145
R2695 VDD.n699 VDD.n692 0.145
R2696 VDD.n704 VDD.n699 0.145
R2697 VDD.n716 VDD.n709 0.145
R2698 VDD.n721 VDD.n716 0.145
R2699 VDD.n726 VDD.n721 0.145
R2700 VDD.n730 VDD.n726 0.145
R2701 VDD.n734 VDD.n730 0.145
R2702 VDD.n764 VDD.n760 0.145
R2703 VDD.n768 VDD.n764 0.145
R2704 VDD.n773 VDD.n768 0.145
R2705 VDD.n780 VDD.n773 0.145
R2706 VDD.n785 VDD.n780 0.145
R2707 VDD.n797 VDD.n790 0.145
R2708 VDD.n802 VDD.n797 0.145
R2709 VDD.n807 VDD.n802 0.145
R2710 VDD.n811 VDD.n807 0.145
R2711 VDD.n837 VDD.n811 0.145
R2712 VDD.n1645 VDD.n1641 0.145
R2713 VDD.n1641 VDD.n1637 0.145
R2714 VDD.n1637 VDD.n1633 0.145
R2715 VDD.n1633 VDD.n1628 0.145
R2716 VDD.n1628 VDD.n1621 0.145
R2717 VDD.n1616 VDD.n1611 0.145
R2718 VDD.n1611 VDD.n1604 0.145
R2719 VDD.n1604 VDD.n1599 0.145
R2720 VDD.n1599 VDD.n1594 0.145
R2721 VDD.n1594 VDD.n1590 0.145
R2722 VDD.n1564 VDD.n1560 0.145
R2723 VDD.n1560 VDD.n1556 0.145
R2724 VDD.n1556 VDD.n1552 0.145
R2725 VDD.n1552 VDD.n1547 0.145
R2726 VDD.n1547 VDD.n1540 0.145
R2727 VDD.n1535 VDD.n1530 0.145
R2728 VDD.n1530 VDD.n1523 0.145
R2729 VDD.n1523 VDD.n1518 0.145
R2730 VDD.n1518 VDD.n1513 0.145
R2731 VDD.n1513 VDD.n1509 0.145
R2732 VDD.n1483 VDD.n1479 0.145
R2733 VDD.n1479 VDD.n1475 0.145
R2734 VDD.n1475 VDD.n1471 0.145
R2735 VDD.n1471 VDD.n1466 0.145
R2736 VDD.n1466 VDD.n1459 0.145
R2737 VDD.n1454 VDD.n1449 0.145
R2738 VDD.n1449 VDD.n1442 0.145
R2739 VDD.n1442 VDD.n1437 0.145
R2740 VDD.n1437 VDD.n1432 0.145
R2741 VDD.n1432 VDD.n1428 0.145
R2742 VDD.n1402 VDD.n1398 0.145
R2743 VDD.n1398 VDD.n1394 0.145
R2744 VDD.n1394 VDD.n1390 0.145
R2745 VDD.n1390 VDD.n1385 0.145
R2746 VDD.n1385 VDD.n1378 0.145
R2747 VDD.n1373 VDD.n1368 0.145
R2748 VDD.n1368 VDD.n1361 0.145
R2749 VDD.n1361 VDD.n1356 0.145
R2750 VDD.n1356 VDD.n1351 0.145
R2751 VDD.n1351 VDD.n1347 0.145
R2752 VDD.n1321 VDD.n1317 0.145
R2753 VDD.n1317 VDD.n1313 0.145
R2754 VDD.n1313 VDD.n1309 0.145
R2755 VDD.n1309 VDD.n1304 0.145
R2756 VDD.n1304 VDD.n1297 0.145
R2757 VDD.n1292 VDD.n1287 0.145
R2758 VDD.n1287 VDD.n1280 0.145
R2759 VDD.n1280 VDD.n1275 0.145
R2760 VDD.n1275 VDD.n1270 0.145
R2761 VDD.n1270 VDD.n1266 0.145
R2762 VDD.n1240 VDD.n1236 0.145
R2763 VDD.n1236 VDD.n1232 0.145
R2764 VDD.n1232 VDD.n1228 0.145
R2765 VDD.n1228 VDD.n1223 0.145
R2766 VDD.n1223 VDD.n1216 0.145
R2767 VDD.n1211 VDD.n1206 0.145
R2768 VDD.n1206 VDD.n1199 0.145
R2769 VDD.n1199 VDD.n1194 0.145
R2770 VDD.n1194 VDD.n1189 0.145
R2771 VDD.n1189 VDD.n1185 0.145
R2772 VDD.n1159 VDD.n1155 0.145
R2773 VDD.n1155 VDD.n1151 0.145
R2774 VDD.n1151 VDD.n1147 0.145
R2775 VDD.n1147 VDD.n1142 0.145
R2776 VDD.n1142 VDD.n1135 0.145
R2777 VDD.n1130 VDD.n1125 0.145
R2778 VDD.n1125 VDD.n1118 0.145
R2779 VDD.n1118 VDD.n1113 0.145
R2780 VDD.n1113 VDD.n1108 0.145
R2781 VDD.n1108 VDD.n1104 0.145
R2782 VDD.n1078 VDD.n1074 0.145
R2783 VDD.n1074 VDD.n1070 0.145
R2784 VDD.n1070 VDD.n1066 0.145
R2785 VDD.n1066 VDD.n1061 0.145
R2786 VDD.n1061 VDD.n1054 0.145
R2787 VDD.n1049 VDD.n1044 0.145
R2788 VDD.n1044 VDD.n1037 0.145
R2789 VDD.n1037 VDD.n1032 0.145
R2790 VDD.n1032 VDD.n1027 0.145
R2791 VDD.n1027 VDD.n1023 0.145
R2792 VDD.n997 VDD.n993 0.145
R2793 VDD.n993 VDD.n989 0.145
R2794 VDD.n989 VDD.n985 0.145
R2795 VDD.n985 VDD.n980 0.145
R2796 VDD.n980 VDD.n973 0.145
R2797 VDD.n968 VDD.n963 0.145
R2798 VDD.n963 VDD.n956 0.145
R2799 VDD.n956 VDD.n951 0.145
R2800 VDD.n951 VDD.n946 0.145
R2801 VDD.n946 VDD.n942 0.145
R2802 VDD.n915 VDD.n911 0.145
R2803 VDD.n911 VDD.n907 0.145
R2804 VDD.n907 VDD.n903 0.145
R2805 VDD.n903 VDD.n898 0.145
R2806 VDD.n898 VDD.n891 0.145
R2807 VDD.n886 VDD.n881 0.145
R2808 VDD.n881 VDD.n874 0.145
R2809 VDD.n874 VDD.n869 0.145
R2810 VDD.n869 VDD.n864 0.145
R2811 VDD.n864 VDD.n860 0.145
R2812 VDD VDD.n837 0.07
R2813 a_15991_989.n2 a_15991_989.t9 512.525
R2814 a_15991_989.n0 a_15991_989.t14 477.179
R2815 a_15991_989.n5 a_15991_989.t7 454.685
R2816 a_15991_989.n5 a_15991_989.t13 428.979
R2817 a_15991_989.n0 a_15991_989.t12 406.485
R2818 a_15991_989.n2 a_15991_989.t10 371.139
R2819 a_15991_989.n1 a_15991_989.t8 363.924
R2820 a_15991_989.n4 a_15991_989.t11 303.606
R2821 a_15991_989.n6 a_15991_989.t15 184.853
R2822 a_15991_989.n11 a_15991_989.n10 159.998
R2823 a_15991_989.n11 a_15991_989.n6 156.035
R2824 a_15991_989.n12 a_15991_989.n4 153.043
R2825 a_15991_989.n6 a_15991_989.n5 151.553
R2826 a_15991_989.n16 a_15991_989.n12 144.246
R2827 a_15991_989.n3 a_15991_989.n1 101.359
R2828 a_15991_989.n12 a_15991_989.n11 79.658
R2829 a_15991_989.n15 a_15991_989.n14 79.232
R2830 a_15991_989.n3 a_15991_989.n2 71.88
R2831 a_15991_989.n16 a_15991_989.n15 63.152
R2832 a_15991_989.n4 a_15991_989.n3 53.891
R2833 a_15991_989.n10 a_15991_989.n9 30
R2834 a_15991_989.n8 a_15991_989.n7 24.383
R2835 a_15991_989.n10 a_15991_989.n8 23.684
R2836 a_15991_989.n15 a_15991_989.n13 16.08
R2837 a_15991_989.n17 a_15991_989.n16 16.078
R2838 a_15991_989.n1 a_15991_989.n0 15.776
R2839 a_15991_989.n13 a_15991_989.t6 14.282
R2840 a_15991_989.n13 a_15991_989.t0 14.282
R2841 a_15991_989.n14 a_15991_989.t1 14.282
R2842 a_15991_989.n14 a_15991_989.t2 14.282
R2843 a_15991_989.t5 a_15991_989.n17 14.282
R2844 a_15991_989.n17 a_15991_989.t4 14.282
R2845 a_15669_1050.n0 a_15669_1050.t9 512.525
R2846 a_15669_1050.n0 a_15669_1050.t7 371.139
R2847 a_15669_1050.n1 a_15669_1050.t8 287.668
R2848 a_15669_1050.n6 a_15669_1050.n5 213.104
R2849 a_15669_1050.n10 a_15669_1050.n6 170.799
R2850 a_15669_1050.n1 a_15669_1050.n0 162.713
R2851 a_15669_1050.n6 a_15669_1050.n1 153.315
R2852 a_15669_1050.n9 a_15669_1050.n8 79.232
R2853 a_15669_1050.n10 a_15669_1050.n9 63.152
R2854 a_15669_1050.n5 a_15669_1050.n4 30
R2855 a_15669_1050.n3 a_15669_1050.n2 24.383
R2856 a_15669_1050.n5 a_15669_1050.n3 23.684
R2857 a_15669_1050.n9 a_15669_1050.n7 16.08
R2858 a_15669_1050.n11 a_15669_1050.n10 16.078
R2859 a_15669_1050.n7 a_15669_1050.t6 14.282
R2860 a_15669_1050.n7 a_15669_1050.t0 14.282
R2861 a_15669_1050.n8 a_15669_1050.t2 14.282
R2862 a_15669_1050.n8 a_15669_1050.t1 14.282
R2863 a_15669_1050.n11 a_15669_1050.t4 14.282
R2864 a_15669_1050.t5 a_15669_1050.n11 14.282
R2865 a_11821_1050.n7 a_11821_1050.t7 512.525
R2866 a_11821_1050.n5 a_11821_1050.t12 512.525
R2867 a_11821_1050.n7 a_11821_1050.t11 371.139
R2868 a_11821_1050.n5 a_11821_1050.t8 371.139
R2869 a_11821_1050.n8 a_11821_1050.t9 234.921
R2870 a_11821_1050.n6 a_11821_1050.t10 234.921
R2871 a_11821_1050.n10 a_11821_1050.n4 223.546
R2872 a_11821_1050.n8 a_11821_1050.n7 215.46
R2873 a_11821_1050.n6 a_11821_1050.n5 215.46
R2874 a_11821_1050.n12 a_11821_1050.n10 166.879
R2875 a_11821_1050.n9 a_11821_1050.n6 79.491
R2876 a_11821_1050.n3 a_11821_1050.n2 79.232
R2877 a_11821_1050.n10 a_11821_1050.n9 77.315
R2878 a_11821_1050.n9 a_11821_1050.n8 76
R2879 a_11821_1050.n4 a_11821_1050.n3 63.152
R2880 a_11821_1050.n4 a_11821_1050.n0 16.08
R2881 a_11821_1050.n3 a_11821_1050.n1 16.08
R2882 a_11821_1050.n12 a_11821_1050.n11 15.218
R2883 a_11821_1050.n0 a_11821_1050.t6 14.282
R2884 a_11821_1050.n0 a_11821_1050.t1 14.282
R2885 a_11821_1050.n1 a_11821_1050.t0 14.282
R2886 a_11821_1050.n1 a_11821_1050.t3 14.282
R2887 a_11821_1050.n2 a_11821_1050.t2 14.282
R2888 a_11821_1050.n2 a_11821_1050.t4 14.282
R2889 a_11821_1050.n13 a_11821_1050.n12 12.014
R2890 a_12143_989.n1 a_12143_989.t7 512.525
R2891 a_12143_989.n3 a_12143_989.t8 454.685
R2892 a_12143_989.n3 a_12143_989.t12 428.979
R2893 a_12143_989.n1 a_12143_989.t10 371.139
R2894 a_12143_989.n2 a_12143_989.t9 287.668
R2895 a_12143_989.n4 a_12143_989.t11 237.959
R2896 a_12143_989.n10 a_12143_989.n9 213.104
R2897 a_12143_989.n11 a_12143_989.n10 170.799
R2898 a_12143_989.n2 a_12143_989.n1 162.713
R2899 a_12143_989.n4 a_12143_989.n3 98.447
R2900 a_12143_989.n5 a_12143_989.n2 84.388
R2901 a_12143_989.n5 a_12143_989.n4 80.035
R2902 a_12143_989.n13 a_12143_989.n12 79.232
R2903 a_12143_989.n10 a_12143_989.n5 76
R2904 a_12143_989.n13 a_12143_989.n11 63.152
R2905 a_12143_989.n9 a_12143_989.n8 30
R2906 a_12143_989.n7 a_12143_989.n6 24.383
R2907 a_12143_989.n9 a_12143_989.n7 23.684
R2908 a_12143_989.n11 a_12143_989.n0 16.08
R2909 a_12143_989.n14 a_12143_989.n13 16.078
R2910 a_12143_989.n0 a_12143_989.t6 14.282
R2911 a_12143_989.n0 a_12143_989.t5 14.282
R2912 a_12143_989.n12 a_12143_989.t3 14.282
R2913 a_12143_989.n12 a_12143_989.t2 14.282
R2914 a_12143_989.t1 a_12143_989.n14 14.282
R2915 a_12143_989.n14 a_12143_989.t0 14.282
R2916 a_4125_1050.n5 a_4125_1050.t8 512.525
R2917 a_4125_1050.n5 a_4125_1050.t9 371.139
R2918 a_4125_1050.n6 a_4125_1050.t7 287.668
R2919 a_4125_1050.n9 a_4125_1050.n7 219.626
R2920 a_4125_1050.n7 a_4125_1050.n4 170.799
R2921 a_4125_1050.n6 a_4125_1050.n5 162.713
R2922 a_4125_1050.n7 a_4125_1050.n6 153.315
R2923 a_4125_1050.n3 a_4125_1050.n2 79.232
R2924 a_4125_1050.n4 a_4125_1050.n3 63.152
R2925 a_4125_1050.n4 a_4125_1050.n0 16.08
R2926 a_4125_1050.n3 a_4125_1050.n1 16.08
R2927 a_4125_1050.n9 a_4125_1050.n8 15.218
R2928 a_4125_1050.n0 a_4125_1050.t1 14.282
R2929 a_4125_1050.n0 a_4125_1050.t5 14.282
R2930 a_4125_1050.n1 a_4125_1050.t0 14.282
R2931 a_4125_1050.n1 a_4125_1050.t2 14.282
R2932 a_4125_1050.n2 a_4125_1050.t3 14.282
R2933 a_4125_1050.n2 a_4125_1050.t6 14.282
R2934 a_4125_1050.n10 a_4125_1050.n9 12.014
R2935 a_4901_103.n5 a_4901_103.n4 19.724
R2936 a_4901_103.t0 a_4901_103.n3 11.595
R2937 a_4901_103.t0 a_4901_103.n5 9.207
R2938 a_4901_103.n2 a_4901_103.n1 2.455
R2939 a_4901_103.n2 a_4901_103.n0 1.32
R2940 a_4901_103.t0 a_4901_103.n2 0.246
R2941 SN.n14 SN.t6 479.223
R2942 SN.n11 SN.t12 479.223
R2943 SN.n8 SN.t13 479.223
R2944 SN.n5 SN.t1 479.223
R2945 SN.n2 SN.t14 479.223
R2946 SN.n0 SN.t0 479.223
R2947 SN.n14 SN.t15 375.52
R2948 SN.n11 SN.t2 375.52
R2949 SN.n8 SN.t4 375.52
R2950 SN.n5 SN.t5 375.52
R2951 SN.n2 SN.t7 375.52
R2952 SN.n0 SN.t10 375.52
R2953 SN.n12 SN.n11 201.982
R2954 SN.n6 SN.n5 201.982
R2955 SN.n1 SN.n0 201.982
R2956 SN.n3 SN.n2 199.731
R2957 SN.n9 SN.n8 199.731
R2958 SN.n15 SN.n14 199.731
R2959 SN.n12 SN.t17 141.649
R2960 SN.n6 SN.t8 141.649
R2961 SN.n1 SN.t9 141.649
R2962 SN.n15 SN.t16 128.128
R2963 SN.n9 SN.t3 128.128
R2964 SN.n3 SN.t11 128.128
R2965 SN.n4 SN.n1 86.561
R2966 SN.n7 SN.n6 76
R2967 SN.n13 SN.n12 76
R2968 SN.n4 SN.n3 49.346
R2969 SN.n10 SN.n9 49.346
R2970 SN.n16 SN.n15 49.346
R2971 SN.n7 SN.n4 10.564
R2972 SN.n13 SN.n10 10.564
R2973 SN.n10 SN.n7 10.561
R2974 SN.n16 SN.n13 10.561
R2975 SN.n16 SN 0.046
R2976 a_6371_989.n1 a_6371_989.t12 512.525
R2977 a_6371_989.n3 a_6371_989.t7 454.685
R2978 a_6371_989.n3 a_6371_989.t10 428.979
R2979 a_6371_989.n1 a_6371_989.t9 371.139
R2980 a_6371_989.n2 a_6371_989.t8 287.668
R2981 a_6371_989.n4 a_6371_989.t11 237.959
R2982 a_6371_989.n7 a_6371_989.n6 234.843
R2983 a_6371_989.n8 a_6371_989.n7 170.799
R2984 a_6371_989.n2 a_6371_989.n1 162.713
R2985 a_6371_989.n4 a_6371_989.n3 98.447
R2986 a_6371_989.n5 a_6371_989.n2 84.388
R2987 a_6371_989.n5 a_6371_989.n4 80.035
R2988 a_6371_989.n10 a_6371_989.n9 79.232
R2989 a_6371_989.n7 a_6371_989.n5 76
R2990 a_6371_989.n10 a_6371_989.n8 63.152
R2991 a_6371_989.n8 a_6371_989.n0 16.08
R2992 a_6371_989.n11 a_6371_989.n10 16.078
R2993 a_6371_989.n0 a_6371_989.t0 14.282
R2994 a_6371_989.n0 a_6371_989.t5 14.282
R2995 a_6371_989.n9 a_6371_989.t3 14.282
R2996 a_6371_989.n9 a_6371_989.t4 14.282
R2997 a_6371_989.t2 a_6371_989.n11 14.282
R2998 a_6371_989.n11 a_6371_989.t1 14.282
R2999 a_4447_989.n3 a_4447_989.t14 512.525
R3000 a_4447_989.n2 a_4447_989.t13 512.525
R3001 a_4447_989.n7 a_4447_989.t10 454.685
R3002 a_4447_989.n7 a_4447_989.t15 428.979
R3003 a_4447_989.n3 a_4447_989.t8 371.139
R3004 a_4447_989.n2 a_4447_989.t9 371.139
R3005 a_4447_989.n4 a_4447_989.n3 265.439
R3006 a_4447_989.n13 a_4447_989.n12 202.074
R3007 a_4447_989.n8 a_4447_989.t12 200.159
R3008 a_4447_989.n14 a_4447_989.n13 197.352
R3009 a_4447_989.n6 a_4447_989.n2 185.78
R3010 a_4447_989.n4 a_4447_989.t7 176.995
R3011 a_4447_989.n5 a_4447_989.t11 170.569
R3012 a_4447_989.n5 a_4447_989.n4 153.043
R3013 a_4447_989.n8 a_4447_989.n7 125
R3014 a_4447_989.n9 a_4447_989.n6 123.293
R3015 a_4447_989.n9 a_4447_989.n8 80.035
R3016 a_4447_989.n6 a_4447_989.n5 79.658
R3017 a_4447_989.n16 a_4447_989.n15 79.231
R3018 a_4447_989.n13 a_4447_989.n9 76
R3019 a_4447_989.n15 a_4447_989.n14 63.152
R3020 a_4447_989.n12 a_4447_989.n11 22.578
R3021 a_4447_989.n14 a_4447_989.n1 16.08
R3022 a_4447_989.n15 a_4447_989.n0 16.08
R3023 a_4447_989.n1 a_4447_989.t6 14.282
R3024 a_4447_989.n1 a_4447_989.t4 14.282
R3025 a_4447_989.n0 a_4447_989.t2 14.282
R3026 a_4447_989.n0 a_4447_989.t3 14.282
R3027 a_4447_989.t1 a_4447_989.n16 14.282
R3028 a_4447_989.n16 a_4447_989.t0 14.282
R3029 a_4447_989.n12 a_4447_989.n10 8.58
R3030 a_18760_101.t0 a_18760_101.n1 34.62
R3031 a_18760_101.t0 a_18760_101.n0 8.137
R3032 a_18760_101.t0 a_18760_101.n2 4.69
R3033 a_18094_101.t0 a_18094_101.n0 34.606
R3034 a_18094_101.t0 a_18094_101.n1 2.115
R3035 a_2201_1050.n1 a_2201_1050.t7 512.525
R3036 a_2201_1050.n1 a_2201_1050.t8 371.139
R3037 a_2201_1050.n2 a_2201_1050.t9 234.562
R3038 a_2201_1050.n5 a_2201_1050.n4 223.905
R3039 a_2201_1050.n2 a_2201_1050.n1 215.819
R3040 a_2201_1050.n4 a_2201_1050.n3 181.737
R3041 a_2201_1050.n4 a_2201_1050.n2 153.315
R3042 a_2201_1050.n7 a_2201_1050.n6 79.232
R3043 a_2201_1050.n7 a_2201_1050.n5 63.152
R3044 a_2201_1050.n5 a_2201_1050.n0 16.08
R3045 a_2201_1050.n8 a_2201_1050.n7 16.078
R3046 a_2201_1050.n0 a_2201_1050.t5 14.282
R3047 a_2201_1050.n0 a_2201_1050.t4 14.282
R3048 a_2201_1050.n6 a_2201_1050.t1 14.282
R3049 a_2201_1050.n6 a_2201_1050.t6 14.282
R3050 a_2201_1050.t3 a_2201_1050.n8 14.282
R3051 a_2201_1050.n8 a_2201_1050.t2 14.282
R3052 a_1561_989.n3 a_1561_989.t14 454.685
R3053 a_1561_989.n5 a_1561_989.t7 454.685
R3054 a_1561_989.n1 a_1561_989.t15 454.685
R3055 a_1561_989.n3 a_1561_989.t8 428.979
R3056 a_1561_989.n5 a_1561_989.t11 428.979
R3057 a_1561_989.n1 a_1561_989.t13 428.979
R3058 a_1561_989.n4 a_1561_989.t9 264.512
R3059 a_1561_989.n2 a_1561_989.t12 264.512
R3060 a_1561_989.n6 a_1561_989.t10 264.173
R3061 a_1561_989.n10 a_1561_989.n9 261.396
R3062 a_1561_989.n11 a_1561_989.n10 144.246
R3063 a_1561_989.n8 a_1561_989.n2 82.484
R3064 a_1561_989.n7 a_1561_989.n6 79.495
R3065 a_1561_989.n13 a_1561_989.n12 79.232
R3066 a_1561_989.n7 a_1561_989.n4 76
R3067 a_1561_989.n10 a_1561_989.n8 76
R3068 a_1561_989.n4 a_1561_989.n3 71.894
R3069 a_1561_989.n2 a_1561_989.n1 71.894
R3070 a_1561_989.n6 a_1561_989.n5 71.555
R3071 a_1561_989.n13 a_1561_989.n11 63.152
R3072 a_1561_989.n11 a_1561_989.n0 16.08
R3073 a_1561_989.n14 a_1561_989.n13 16.078
R3074 a_1561_989.n0 a_1561_989.t6 14.282
R3075 a_1561_989.n0 a_1561_989.t5 14.282
R3076 a_1561_989.n12 a_1561_989.t4 14.282
R3077 a_1561_989.n12 a_1561_989.t3 14.282
R3078 a_1561_989.t2 a_1561_989.n14 14.282
R3079 a_1561_989.n14 a_1561_989.t1 14.282
R3080 a_1561_989.n8 a_1561_989.n7 4.035
R3081 a_7333_989.n3 a_7333_989.t9 454.685
R3082 a_7333_989.n5 a_7333_989.t12 454.685
R3083 a_7333_989.n1 a_7333_989.t10 454.685
R3084 a_7333_989.n3 a_7333_989.t7 428.979
R3085 a_7333_989.n5 a_7333_989.t8 428.979
R3086 a_7333_989.n1 a_7333_989.t15 428.979
R3087 a_7333_989.n4 a_7333_989.t13 264.512
R3088 a_7333_989.n2 a_7333_989.t14 264.512
R3089 a_7333_989.n6 a_7333_989.t11 264.173
R3090 a_7333_989.n10 a_7333_989.n9 261.396
R3091 a_7333_989.n11 a_7333_989.n10 144.246
R3092 a_7333_989.n8 a_7333_989.n2 82.484
R3093 a_7333_989.n7 a_7333_989.n6 79.495
R3094 a_7333_989.n13 a_7333_989.n12 79.232
R3095 a_7333_989.n7 a_7333_989.n4 76
R3096 a_7333_989.n10 a_7333_989.n8 76
R3097 a_7333_989.n4 a_7333_989.n3 71.894
R3098 a_7333_989.n2 a_7333_989.n1 71.894
R3099 a_7333_989.n6 a_7333_989.n5 71.555
R3100 a_7333_989.n13 a_7333_989.n11 63.152
R3101 a_7333_989.n11 a_7333_989.n0 16.08
R3102 a_7333_989.n14 a_7333_989.n13 16.078
R3103 a_7333_989.n0 a_7333_989.t2 14.282
R3104 a_7333_989.n0 a_7333_989.t6 14.282
R3105 a_7333_989.n12 a_7333_989.t3 14.282
R3106 a_7333_989.n12 a_7333_989.t4 14.282
R3107 a_7333_989.n14 a_7333_989.t0 14.282
R3108 a_7333_989.t1 a_7333_989.n14 14.282
R3109 a_7333_989.n8 a_7333_989.n7 4.035
R3110 a_7973_1050.n0 a_7973_1050.t8 512.525
R3111 a_7973_1050.n0 a_7973_1050.t9 371.139
R3112 a_7973_1050.n1 a_7973_1050.t7 234.562
R3113 a_7973_1050.n10 a_7973_1050.n6 223.905
R3114 a_7973_1050.n1 a_7973_1050.n0 215.819
R3115 a_7973_1050.n6 a_7973_1050.n5 159.998
R3116 a_7973_1050.n6 a_7973_1050.n1 153.315
R3117 a_7973_1050.n9 a_7973_1050.n8 79.232
R3118 a_7973_1050.n10 a_7973_1050.n9 63.152
R3119 a_7973_1050.n5 a_7973_1050.n4 30
R3120 a_7973_1050.n3 a_7973_1050.n2 24.383
R3121 a_7973_1050.n5 a_7973_1050.n3 23.684
R3122 a_7973_1050.n9 a_7973_1050.n7 16.08
R3123 a_7973_1050.n11 a_7973_1050.n10 16.078
R3124 a_7973_1050.n7 a_7973_1050.t3 14.282
R3125 a_7973_1050.n7 a_7973_1050.t4 14.282
R3126 a_7973_1050.n8 a_7973_1050.t6 14.282
R3127 a_7973_1050.n8 a_7973_1050.t5 14.282
R3128 a_7973_1050.t2 a_7973_1050.n11 14.282
R3129 a_7973_1050.n11 a_7973_1050.t1 14.282
R3130 a_9897_1050.n2 a_9897_1050.t8 512.525
R3131 a_9897_1050.n2 a_9897_1050.t9 371.139
R3132 a_9897_1050.n3 a_9897_1050.t7 287.668
R3133 a_9897_1050.n8 a_9897_1050.n7 213.104
R3134 a_9897_1050.n9 a_9897_1050.n8 170.799
R3135 a_9897_1050.n3 a_9897_1050.n2 162.713
R3136 a_9897_1050.n8 a_9897_1050.n3 153.315
R3137 a_9897_1050.n11 a_9897_1050.n10 79.231
R3138 a_9897_1050.n10 a_9897_1050.n9 63.152
R3139 a_9897_1050.n7 a_9897_1050.n6 30
R3140 a_9897_1050.n5 a_9897_1050.n4 24.383
R3141 a_9897_1050.n7 a_9897_1050.n5 23.684
R3142 a_9897_1050.n9 a_9897_1050.n1 16.08
R3143 a_9897_1050.n10 a_9897_1050.n0 16.08
R3144 a_9897_1050.n1 a_9897_1050.t3 14.282
R3145 a_9897_1050.n1 a_9897_1050.t2 14.282
R3146 a_9897_1050.n0 a_9897_1050.t6 14.282
R3147 a_9897_1050.n0 a_9897_1050.t5 14.282
R3148 a_9897_1050.n11 a_9897_1050.t0 14.282
R3149 a_9897_1050.t1 a_9897_1050.n11 14.282
R3150 a_18197_1051.n4 a_18197_1051.n3 196.002
R3151 a_18197_1051.n2 a_18197_1051.t0 89.553
R3152 a_18197_1051.n5 a_18197_1051.n4 75.27
R3153 a_18197_1051.n3 a_18197_1051.n2 75.214
R3154 a_18197_1051.n4 a_18197_1051.n0 36.52
R3155 a_18197_1051.n3 a_18197_1051.t6 14.338
R3156 a_18197_1051.n0 a_18197_1051.t5 14.282
R3157 a_18197_1051.n0 a_18197_1051.t4 14.282
R3158 a_18197_1051.n1 a_18197_1051.t1 14.282
R3159 a_18197_1051.n1 a_18197_1051.t7 14.282
R3160 a_18197_1051.n5 a_18197_1051.t2 14.282
R3161 a_18197_1051.t3 a_18197_1051.n5 14.282
R3162 a_18197_1051.n2 a_18197_1051.n1 12.119
R3163 QN.n13 QN.n12 216.728
R3164 QN.n13 QN.n2 126.664
R3165 QN.n10 QN.n5 111.94
R3166 QN.n10 QN.n9 98.501
R3167 QN.n12 QN.n10 78.403
R3168 QN.n14 QN.n13 76
R3169 QN.n2 QN.n1 75.271
R3170 QN.n12 QN.n11 42.274
R3171 QN.n9 QN.n8 30
R3172 QN.n7 QN.n6 24.383
R3173 QN.n9 QN.n7 23.684
R3174 QN.n5 QN.n4 22.578
R3175 QN.n0 QN.t3 14.282
R3176 QN.n0 QN.t2 14.282
R3177 QN.n1 QN.t5 14.282
R3178 QN.n1 QN.t6 14.282
R3179 QN.n2 QN.n0 12.119
R3180 QN.n5 QN.n3 8.58
R3181 QN.n14 QN 0.046
R3182 RN.n23 RN.t5 479.223
R3183 RN.n17 RN.t21 479.223
R3184 RN.n14 RN.t10 479.223
R3185 RN.n8 RN.t3 479.223
R3186 RN.n5 RN.t15 479.223
R3187 RN.n0 RN.t2 479.223
R3188 RN.n20 RN.t20 454.685
R3189 RN.n11 RN.t0 454.685
R3190 RN.n2 RN.t4 454.685
R3191 RN.n20 RN.t7 428.979
R3192 RN.n11 RN.t17 428.979
R3193 RN.n2 RN.t22 428.979
R3194 RN.n23 RN.t18 375.52
R3195 RN.n17 RN.t9 375.52
R3196 RN.n14 RN.t26 375.52
R3197 RN.n8 RN.t14 375.52
R3198 RN.n5 RN.t19 375.52
R3199 RN.n0 RN.t13 375.52
R3200 RN.n21 RN.n20 178.106
R3201 RN.n12 RN.n11 178.106
R3202 RN.n3 RN.n2 178.106
R3203 RN.n24 RN.n23 175.429
R3204 RN.n18 RN.n17 175.429
R3205 RN.n15 RN.n14 175.429
R3206 RN.n9 RN.n8 175.429
R3207 RN.n6 RN.n5 175.429
R3208 RN.n1 RN.n0 175.429
R3209 RN.n24 RN.t11 162.048
R3210 RN.n18 RN.t23 162.048
R3211 RN.n15 RN.t1 162.048
R3212 RN.n9 RN.t8 162.048
R3213 RN.n6 RN.t6 162.048
R3214 RN.n1 RN.t12 162.048
R3215 RN.n21 RN.t16 158.3
R3216 RN.n12 RN.t25 158.3
R3217 RN.n3 RN.t24 158.3
R3218 RN.n4 RN.n1 78.675
R3219 RN.n4 RN.n3 76
R3220 RN.n7 RN.n6 76
R3221 RN.n10 RN.n9 76
R3222 RN.n13 RN.n12 76
R3223 RN.n16 RN.n15 76
R3224 RN.n19 RN.n18 76
R3225 RN.n22 RN.n21 76
R3226 RN.n25 RN.n24 76
R3227 RN.n7 RN.n4 11.381
R3228 RN.n16 RN.n13 11.381
R3229 RN.n25 RN.n22 11.381
R3230 RN.n10 RN.n7 7.028
R3231 RN.n19 RN.n16 7.028
R3232 RN.n13 RN.n10 2.675
R3233 RN.n22 RN.n19 2.675
R3234 RN.n25 RN 0.046
R3235 a_5863_103.n1 a_5863_103.n0 25.576
R3236 a_5863_103.n3 a_5863_103.n2 9.111
R3237 a_5863_103.n7 a_5863_103.n5 7.859
R3238 a_5863_103.t0 a_5863_103.n7 3.034
R3239 a_5863_103.n5 a_5863_103.n3 1.964
R3240 a_5863_103.n5 a_5863_103.n4 1.964
R3241 a_5863_103.t0 a_5863_103.n1 1.871
R3242 a_5863_103.n7 a_5863_103.n6 0.443
R3243 a_6144_210.n10 a_6144_210.n8 82.852
R3244 a_6144_210.n11 a_6144_210.n0 49.6
R3245 a_6144_210.n7 a_6144_210.n6 32.833
R3246 a_6144_210.n8 a_6144_210.t1 32.416
R3247 a_6144_210.n10 a_6144_210.n9 27.2
R3248 a_6144_210.n3 a_6144_210.n2 23.284
R3249 a_6144_210.n11 a_6144_210.n10 22.4
R3250 a_6144_210.n7 a_6144_210.n4 19.017
R3251 a_6144_210.n6 a_6144_210.n5 13.494
R3252 a_6144_210.t1 a_6144_210.n1 7.04
R3253 a_6144_210.t1 a_6144_210.n3 5.727
R3254 a_6144_210.n8 a_6144_210.n7 1.435
R3255 D.n5 D.t2 512.525
R3256 D.n2 D.t1 512.525
R3257 D.n0 D.t3 512.525
R3258 D.n5 D.t7 371.139
R3259 D.n2 D.t6 371.139
R3260 D.n0 D.t8 371.139
R3261 D.n6 D.t5 340.774
R3262 D.n3 D.t4 340.774
R3263 D.n1 D.t0 340.774
R3264 D.n6 D.n5 109.607
R3265 D.n3 D.n2 109.607
R3266 D.n1 D.n0 109.607
R3267 D.n4 D.n1 97.175
R3268 D.n4 D.n3 76
R3269 D.n7 D.n6 76
R3270 D.n7 D.n4 21.175
R3271 D.n7 D 0.046
R3272 a_11635_103.n1 a_11635_103.n0 25.576
R3273 a_11635_103.n3 a_11635_103.n2 9.111
R3274 a_11635_103.n7 a_11635_103.n5 7.859
R3275 a_11635_103.t0 a_11635_103.n7 3.034
R3276 a_11635_103.n5 a_11635_103.n3 1.964
R3277 a_11635_103.n5 a_11635_103.n4 1.964
R3278 a_11635_103.t0 a_11635_103.n1 1.871
R3279 a_11635_103.n7 a_11635_103.n6 0.443
R3280 a_16726_210.n10 a_16726_210.n8 82.852
R3281 a_16726_210.n7 a_16726_210.n6 32.833
R3282 a_16726_210.n8 a_16726_210.t1 32.416
R3283 a_16726_210.n10 a_16726_210.n9 27.2
R3284 a_16726_210.n11 a_16726_210.n0 23.498
R3285 a_16726_210.n3 a_16726_210.n2 23.284
R3286 a_16726_210.n11 a_16726_210.n10 22.4
R3287 a_16726_210.n7 a_16726_210.n4 19.017
R3288 a_16726_210.n6 a_16726_210.n5 13.494
R3289 a_16726_210.t1 a_16726_210.n1 7.04
R3290 a_16726_210.t1 a_16726_210.n3 5.727
R3291 a_16726_210.n8 a_16726_210.n7 1.435
R3292 a_7787_103.n1 a_7787_103.n0 25.576
R3293 a_7787_103.n3 a_7787_103.n2 9.111
R3294 a_7787_103.n7 a_7787_103.n5 7.859
R3295 a_7787_103.t0 a_7787_103.n7 3.034
R3296 a_7787_103.n5 a_7787_103.n3 1.964
R3297 a_7787_103.n5 a_7787_103.n4 1.964
R3298 a_7787_103.t0 a_7787_103.n1 1.871
R3299 a_7787_103.n7 a_7787_103.n6 0.443
R3300 a_8068_210.n8 a_8068_210.n6 96.467
R3301 a_8068_210.n3 a_8068_210.n1 44.628
R3302 a_8068_210.t0 a_8068_210.n8 32.417
R3303 a_8068_210.n3 a_8068_210.n2 23.284
R3304 a_8068_210.n6 a_8068_210.n5 22.349
R3305 a_8068_210.t0 a_8068_210.n10 20.241
R3306 a_8068_210.n10 a_8068_210.n9 13.494
R3307 a_8068_210.n6 a_8068_210.n4 8.443
R3308 a_8068_210.t0 a_8068_210.n0 8.137
R3309 a_8068_210.t0 a_8068_210.n3 5.727
R3310 a_8068_210.n8 a_8068_210.n7 1.435
R3311 a_277_1050.n3 a_277_1050.t9 512.525
R3312 a_277_1050.n1 a_277_1050.t7 512.525
R3313 a_277_1050.n3 a_277_1050.t11 371.139
R3314 a_277_1050.n1 a_277_1050.t12 371.139
R3315 a_277_1050.n4 a_277_1050.t10 234.921
R3316 a_277_1050.n2 a_277_1050.t8 234.921
R3317 a_277_1050.n8 a_277_1050.n7 223.546
R3318 a_277_1050.n4 a_277_1050.n3 215.46
R3319 a_277_1050.n2 a_277_1050.n1 215.46
R3320 a_277_1050.n7 a_277_1050.n6 182.096
R3321 a_277_1050.n5 a_277_1050.n2 79.491
R3322 a_277_1050.n10 a_277_1050.n9 79.232
R3323 a_277_1050.n7 a_277_1050.n5 77.315
R3324 a_277_1050.n5 a_277_1050.n4 76
R3325 a_277_1050.n10 a_277_1050.n8 63.152
R3326 a_277_1050.n8 a_277_1050.n0 16.08
R3327 a_277_1050.n11 a_277_1050.n10 16.078
R3328 a_277_1050.n0 a_277_1050.t5 14.282
R3329 a_277_1050.n0 a_277_1050.t4 14.282
R3330 a_277_1050.n9 a_277_1050.t3 14.282
R3331 a_277_1050.n9 a_277_1050.t2 14.282
R3332 a_277_1050.t1 a_277_1050.n11 14.282
R3333 a_277_1050.n11 a_277_1050.t0 14.282
R3334 a_9711_103.n1 a_9711_103.n0 25.576
R3335 a_9711_103.n3 a_9711_103.n2 9.111
R3336 a_9711_103.n7 a_9711_103.n5 7.859
R3337 a_9711_103.t0 a_9711_103.n7 3.034
R3338 a_9711_103.n5 a_9711_103.n3 1.964
R3339 a_9711_103.n5 a_9711_103.n4 1.964
R3340 a_9711_103.t0 a_9711_103.n1 1.871
R3341 a_9711_103.n7 a_9711_103.n6 0.443
R3342 a_599_989.n0 a_599_989.t12 512.525
R3343 a_599_989.n2 a_599_989.t10 454.685
R3344 a_599_989.n2 a_599_989.t9 428.979
R3345 a_599_989.n0 a_599_989.t8 371.139
R3346 a_599_989.n1 a_599_989.t11 287.668
R3347 a_599_989.n3 a_599_989.t7 237.959
R3348 a_599_989.n9 a_599_989.n8 213.104
R3349 a_599_989.n13 a_599_989.n9 170.799
R3350 a_599_989.n1 a_599_989.n0 162.713
R3351 a_599_989.n3 a_599_989.n2 98.447
R3352 a_599_989.n4 a_599_989.n1 84.388
R3353 a_599_989.n4 a_599_989.n3 80.035
R3354 a_599_989.n12 a_599_989.n11 79.232
R3355 a_599_989.n9 a_599_989.n4 76
R3356 a_599_989.n13 a_599_989.n12 63.152
R3357 a_599_989.n8 a_599_989.n7 30
R3358 a_599_989.n6 a_599_989.n5 24.383
R3359 a_599_989.n8 a_599_989.n6 23.684
R3360 a_599_989.n12 a_599_989.n10 16.08
R3361 a_599_989.n14 a_599_989.n13 16.078
R3362 a_599_989.n10 a_599_989.t3 14.282
R3363 a_599_989.n10 a_599_989.t4 14.282
R3364 a_599_989.n11 a_599_989.t6 14.282
R3365 a_599_989.n11 a_599_989.t5 14.282
R3366 a_599_989.n14 a_599_989.t0 14.282
R3367 a_599_989.t1 a_599_989.n14 14.282
R3368 a_372_210.n10 a_372_210.n8 82.852
R3369 a_372_210.n7 a_372_210.n6 32.833
R3370 a_372_210.n8 a_372_210.t1 32.416
R3371 a_372_210.n10 a_372_210.n9 27.2
R3372 a_372_210.n11 a_372_210.n0 23.498
R3373 a_372_210.n3 a_372_210.n2 23.284
R3374 a_372_210.n11 a_372_210.n10 22.4
R3375 a_372_210.n7 a_372_210.n4 19.017
R3376 a_372_210.n6 a_372_210.n5 13.494
R3377 a_372_210.t1 a_372_210.n1 7.04
R3378 a_372_210.t1 a_372_210.n3 5.727
R3379 a_372_210.n8 a_372_210.n7 1.435
R3380 a_8749_103.n1 a_8749_103.n0 25.576
R3381 a_8749_103.n3 a_8749_103.n2 9.111
R3382 a_8749_103.n7 a_8749_103.n5 7.859
R3383 a_8749_103.t0 a_8749_103.n7 3.034
R3384 a_8749_103.n5 a_8749_103.n3 1.964
R3385 a_8749_103.n5 a_8749_103.n4 1.964
R3386 a_8749_103.t0 a_8749_103.n1 1.871
R3387 a_8749_103.n7 a_8749_103.n6 0.443
R3388 a_9030_210.n8 a_9030_210.n6 96.467
R3389 a_9030_210.n3 a_9030_210.n1 44.628
R3390 a_9030_210.t0 a_9030_210.n8 32.417
R3391 a_9030_210.n3 a_9030_210.n2 23.284
R3392 a_9030_210.n6 a_9030_210.n5 22.349
R3393 a_9030_210.t0 a_9030_210.n10 20.241
R3394 a_9030_210.n10 a_9030_210.n9 13.494
R3395 a_9030_210.n6 a_9030_210.n4 8.443
R3396 a_9030_210.t0 a_9030_210.n0 8.137
R3397 a_9030_210.t0 a_9030_210.n3 5.727
R3398 a_9030_210.n8 a_9030_210.n7 1.435
R3399 a_12597_103.n1 a_12597_103.n0 25.576
R3400 a_12597_103.n3 a_12597_103.n2 9.111
R3401 a_12597_103.n7 a_12597_103.n5 7.859
R3402 a_12597_103.t0 a_12597_103.n7 3.034
R3403 a_12597_103.n5 a_12597_103.n3 1.964
R3404 a_12597_103.n5 a_12597_103.n4 1.964
R3405 a_12597_103.t0 a_12597_103.n1 1.871
R3406 a_12597_103.n7 a_12597_103.n6 0.443
R3407 a_14521_103.n4 a_14521_103.n3 19.724
R3408 a_14521_103.t0 a_14521_103.n5 11.595
R3409 a_14521_103.t0 a_14521_103.n4 9.207
R3410 a_14521_103.n2 a_14521_103.n0 8.543
R3411 a_14521_103.t0 a_14521_103.n2 3.034
R3412 a_14521_103.n2 a_14521_103.n1 0.443
R3413 a_10673_103.n1 a_10673_103.n0 25.576
R3414 a_10673_103.n3 a_10673_103.n2 9.111
R3415 a_10673_103.n7 a_10673_103.n5 7.859
R3416 a_10673_103.t0 a_10673_103.n7 3.034
R3417 a_10673_103.n5 a_10673_103.n3 1.964
R3418 a_10673_103.n5 a_10673_103.n4 1.964
R3419 a_10673_103.t0 a_10673_103.n1 1.871
R3420 a_10673_103.n7 a_10673_103.n6 0.443
R3421 a_91_103.n1 a_91_103.n0 25.576
R3422 a_91_103.n3 a_91_103.n2 9.111
R3423 a_91_103.n7 a_91_103.n6 2.455
R3424 a_91_103.n5 a_91_103.n3 1.964
R3425 a_91_103.n5 a_91_103.n4 1.964
R3426 a_91_103.t0 a_91_103.n1 1.871
R3427 a_91_103.n7 a_91_103.n5 0.636
R3428 a_91_103.t0 a_91_103.n7 0.246
R3429 a_11916_210.n10 a_11916_210.n8 82.852
R3430 a_11916_210.n11 a_11916_210.n0 49.6
R3431 a_11916_210.n7 a_11916_210.n6 32.833
R3432 a_11916_210.n8 a_11916_210.t1 32.416
R3433 a_11916_210.n10 a_11916_210.n9 27.2
R3434 a_11916_210.n3 a_11916_210.n2 23.284
R3435 a_11916_210.n11 a_11916_210.n10 22.4
R3436 a_11916_210.n7 a_11916_210.n4 19.017
R3437 a_11916_210.n6 a_11916_210.n5 13.494
R3438 a_11916_210.t1 a_11916_210.n1 7.04
R3439 a_11916_210.t1 a_11916_210.n3 5.727
R3440 a_11916_210.n8 a_11916_210.n7 1.435
R3441 a_9992_210.n10 a_9992_210.n8 82.852
R3442 a_9992_210.n11 a_9992_210.n0 49.6
R3443 a_9992_210.n7 a_9992_210.n6 32.833
R3444 a_9992_210.n8 a_9992_210.t1 32.416
R3445 a_9992_210.n10 a_9992_210.n9 27.2
R3446 a_9992_210.n3 a_9992_210.n2 23.284
R3447 a_9992_210.n11 a_9992_210.n10 22.4
R3448 a_9992_210.n7 a_9992_210.n4 19.017
R3449 a_9992_210.n6 a_9992_210.n5 13.494
R3450 a_9992_210.t1 a_9992_210.n1 7.04
R3451 a_9992_210.t1 a_9992_210.n3 5.727
R3452 a_9992_210.n8 a_9992_210.n7 1.435
R3453 a_17428_101.n1 a_17428_101.n0 32.249
R3454 a_17428_101.t0 a_17428_101.n5 7.911
R3455 a_17428_101.n4 a_17428_101.n2 4.032
R3456 a_17428_101.n4 a_17428_101.n3 3.644
R3457 a_17428_101.t0 a_17428_101.n1 2.534
R3458 a_17428_101.t0 a_17428_101.n4 1.099
R3459 a_13559_103.n1 a_13559_103.n0 25.576
R3460 a_13559_103.n3 a_13559_103.n2 9.111
R3461 a_13559_103.n7 a_13559_103.n6 2.455
R3462 a_13559_103.n5 a_13559_103.n3 1.964
R3463 a_13559_103.n5 a_13559_103.n4 1.964
R3464 a_13559_103.t0 a_13559_103.n1 1.871
R3465 a_13559_103.n7 a_13559_103.n5 0.636
R3466 a_13559_103.t0 a_13559_103.n7 0.246
R3467 a_15483_103.n1 a_15483_103.n0 25.576
R3468 a_15483_103.n3 a_15483_103.n2 9.111
R3469 a_15483_103.n7 a_15483_103.n5 7.859
R3470 a_15483_103.t0 a_15483_103.n7 3.034
R3471 a_15483_103.n5 a_15483_103.n3 1.964
R3472 a_15483_103.n5 a_15483_103.n4 1.964
R3473 a_15483_103.t0 a_15483_103.n1 1.871
R3474 a_15483_103.n7 a_15483_103.n6 0.443
R3475 a_14802_210.n8 a_14802_210.n6 96.467
R3476 a_14802_210.n3 a_14802_210.n1 44.628
R3477 a_14802_210.t0 a_14802_210.n8 32.417
R3478 a_14802_210.n3 a_14802_210.n2 23.284
R3479 a_14802_210.n6 a_14802_210.n5 22.349
R3480 a_14802_210.t0 a_14802_210.n10 20.241
R3481 a_14802_210.n10 a_14802_210.n9 13.494
R3482 a_14802_210.n6 a_14802_210.n4 8.443
R3483 a_14802_210.t0 a_14802_210.n0 8.137
R3484 a_14802_210.t0 a_14802_210.n3 5.727
R3485 a_14802_210.n8 a_14802_210.n7 1.435
R3486 a_10954_210.n8 a_10954_210.n6 96.467
R3487 a_10954_210.n3 a_10954_210.n1 44.628
R3488 a_10954_210.t0 a_10954_210.n8 32.417
R3489 a_10954_210.n3 a_10954_210.n2 23.284
R3490 a_10954_210.n6 a_10954_210.n5 22.349
R3491 a_10954_210.t0 a_10954_210.n10 20.241
R3492 a_10954_210.n10 a_10954_210.n9 13.494
R3493 a_10954_210.n6 a_10954_210.n4 8.443
R3494 a_10954_210.t0 a_10954_210.n0 8.137
R3495 a_10954_210.t0 a_10954_210.n3 5.727
R3496 a_10954_210.n8 a_10954_210.n7 1.435
R3497 a_16445_103.n1 a_16445_103.n0 25.576
R3498 a_16445_103.n3 a_16445_103.n2 9.111
R3499 a_16445_103.n7 a_16445_103.n6 2.455
R3500 a_16445_103.n5 a_16445_103.n3 1.964
R3501 a_16445_103.n5 a_16445_103.n4 1.964
R3502 a_16445_103.t0 a_16445_103.n1 1.871
R3503 a_16445_103.n7 a_16445_103.n5 0.636
R3504 a_16445_103.t0 a_16445_103.n7 0.246
R3505 a_12878_210.n10 a_12878_210.n8 82.852
R3506 a_12878_210.n11 a_12878_210.n0 49.6
R3507 a_12878_210.n7 a_12878_210.n6 32.833
R3508 a_12878_210.n8 a_12878_210.t1 32.416
R3509 a_12878_210.n10 a_12878_210.n9 27.2
R3510 a_12878_210.n3 a_12878_210.n2 23.284
R3511 a_12878_210.n11 a_12878_210.n10 22.4
R3512 a_12878_210.n7 a_12878_210.n4 19.017
R3513 a_12878_210.n6 a_12878_210.n5 13.494
R3514 a_12878_210.t1 a_12878_210.n1 7.04
R3515 a_12878_210.t1 a_12878_210.n3 5.727
R3516 a_12878_210.n8 a_12878_210.n7 1.435
R3517 a_2296_210.n9 a_2296_210.n7 82.852
R3518 a_2296_210.n3 a_2296_210.n1 44.628
R3519 a_2296_210.t0 a_2296_210.n9 32.417
R3520 a_2296_210.n7 a_2296_210.n6 27.2
R3521 a_2296_210.n5 a_2296_210.n4 23.498
R3522 a_2296_210.n3 a_2296_210.n2 23.284
R3523 a_2296_210.n7 a_2296_210.n5 22.4
R3524 a_2296_210.t0 a_2296_210.n11 20.241
R3525 a_2296_210.n11 a_2296_210.n10 13.494
R3526 a_2296_210.t0 a_2296_210.n0 8.137
R3527 a_2296_210.t0 a_2296_210.n3 5.727
R3528 a_2296_210.n9 a_2296_210.n8 1.435
R3529 a_4220_210.n10 a_4220_210.n8 82.852
R3530 a_4220_210.n7 a_4220_210.n6 32.833
R3531 a_4220_210.n8 a_4220_210.t1 32.416
R3532 a_4220_210.n10 a_4220_210.n9 27.2
R3533 a_4220_210.n11 a_4220_210.n0 23.498
R3534 a_4220_210.n3 a_4220_210.n2 23.284
R3535 a_4220_210.n11 a_4220_210.n10 22.4
R3536 a_4220_210.n7 a_4220_210.n4 19.017
R3537 a_4220_210.n6 a_4220_210.n5 13.494
R3538 a_4220_210.t1 a_4220_210.n1 7.04
R3539 a_4220_210.t1 a_4220_210.n3 5.727
R3540 a_4220_210.n8 a_4220_210.n7 1.435
R3541 a_15764_210.n10 a_15764_210.n8 82.852
R3542 a_15764_210.n11 a_15764_210.n0 49.6
R3543 a_15764_210.n7 a_15764_210.n6 32.833
R3544 a_15764_210.n8 a_15764_210.t1 32.416
R3545 a_15764_210.n10 a_15764_210.n9 27.2
R3546 a_15764_210.n3 a_15764_210.n2 23.284
R3547 a_15764_210.n11 a_15764_210.n10 22.4
R3548 a_15764_210.n7 a_15764_210.n4 19.017
R3549 a_15764_210.n6 a_15764_210.n5 13.494
R3550 a_15764_210.t1 a_15764_210.n1 7.04
R3551 a_15764_210.t1 a_15764_210.n3 5.727
R3552 a_15764_210.n8 a_15764_210.n7 1.435
R3553 a_2015_103.n1 a_2015_103.n0 25.576
R3554 a_2015_103.n3 a_2015_103.n2 9.111
R3555 a_2015_103.n7 a_2015_103.n6 2.455
R3556 a_2015_103.n5 a_2015_103.n3 1.964
R3557 a_2015_103.n5 a_2015_103.n4 1.964
R3558 a_2015_103.t0 a_2015_103.n1 1.871
R3559 a_2015_103.n7 a_2015_103.n5 0.636
R3560 a_2015_103.t0 a_2015_103.n7 0.246
R3561 a_1334_210.n9 a_1334_210.n7 82.852
R3562 a_1334_210.n3 a_1334_210.n1 44.628
R3563 a_1334_210.t0 a_1334_210.n9 32.417
R3564 a_1334_210.n7 a_1334_210.n6 27.2
R3565 a_1334_210.n5 a_1334_210.n4 23.498
R3566 a_1334_210.n3 a_1334_210.n2 23.284
R3567 a_1334_210.n7 a_1334_210.n5 22.4
R3568 a_1334_210.t0 a_1334_210.n11 20.241
R3569 a_1334_210.n11 a_1334_210.n10 13.494
R3570 a_1334_210.t0 a_1334_210.n0 8.137
R3571 a_1334_210.t0 a_1334_210.n3 5.727
R3572 a_1334_210.n9 a_1334_210.n8 1.435
R3573 a_7106_210.n8 a_7106_210.n6 96.467
R3574 a_7106_210.n3 a_7106_210.n1 44.628
R3575 a_7106_210.t0 a_7106_210.n8 32.417
R3576 a_7106_210.n3 a_7106_210.n2 23.284
R3577 a_7106_210.n6 a_7106_210.n5 22.349
R3578 a_7106_210.t0 a_7106_210.n10 20.241
R3579 a_7106_210.n10 a_7106_210.n9 13.494
R3580 a_7106_210.n6 a_7106_210.n4 8.443
R3581 a_7106_210.t0 a_7106_210.n0 8.137
R3582 a_7106_210.t0 a_7106_210.n3 5.727
R3583 a_7106_210.n8 a_7106_210.n7 1.435
R3584 a_5182_210.n8 a_5182_210.n6 96.467
R3585 a_5182_210.n3 a_5182_210.n1 44.628
R3586 a_5182_210.t0 a_5182_210.n8 32.417
R3587 a_5182_210.n3 a_5182_210.n2 23.284
R3588 a_5182_210.n6 a_5182_210.n5 22.349
R3589 a_5182_210.t0 a_5182_210.n10 20.241
R3590 a_5182_210.n10 a_5182_210.n9 13.494
R3591 a_5182_210.n6 a_5182_210.n4 8.443
R3592 a_5182_210.t0 a_5182_210.n0 8.137
R3593 a_5182_210.t0 a_5182_210.n3 5.727
R3594 a_5182_210.n8 a_5182_210.n7 1.435
R3595 a_1053_103.n1 a_1053_103.n0 25.576
R3596 a_1053_103.n3 a_1053_103.n2 9.111
R3597 a_1053_103.n7 a_1053_103.n6 2.455
R3598 a_1053_103.n5 a_1053_103.n3 1.964
R3599 a_1053_103.n5 a_1053_103.n4 1.964
R3600 a_1053_103.t0 a_1053_103.n1 1.871
R3601 a_1053_103.n7 a_1053_103.n5 0.636
R3602 a_1053_103.t0 a_1053_103.n7 0.246
R3603 a_3939_103.n1 a_3939_103.n0 25.576
R3604 a_3939_103.n3 a_3939_103.n2 9.111
R3605 a_3939_103.n7 a_3939_103.n6 2.455
R3606 a_3939_103.n5 a_3939_103.n3 1.964
R3607 a_3939_103.n5 a_3939_103.n4 1.964
R3608 a_3939_103.t0 a_3939_103.n1 1.871
R3609 a_3939_103.n7 a_3939_103.n5 0.636
R3610 a_3939_103.t0 a_3939_103.n7 0.246
C11 SN GND 9.66fF
C12 RN GND 11.16fF
C13 VDD GND 69.06fF
C14 a_3939_103.n0 GND 0.09fF
C15 a_3939_103.n1 GND 0.10fF
C16 a_3939_103.n2 GND 0.05fF
C17 a_3939_103.n3 GND 0.03fF
C18 a_3939_103.n4 GND 0.04fF
C19 a_3939_103.n5 GND 0.03fF
C20 a_3939_103.n6 GND 0.04fF
C21 a_1053_103.n0 GND 0.09fF
C22 a_1053_103.n1 GND 0.10fF
C23 a_1053_103.n2 GND 0.05fF
C24 a_1053_103.n3 GND 0.03fF
C25 a_1053_103.n4 GND 0.04fF
C26 a_1053_103.n5 GND 0.03fF
C27 a_1053_103.n6 GND 0.04fF
C28 a_5182_210.n0 GND 0.07fF
C29 a_5182_210.n1 GND 0.09fF
C30 a_5182_210.n2 GND 0.13fF
C31 a_5182_210.n3 GND 0.11fF
C32 a_5182_210.n4 GND 0.02fF
C33 a_5182_210.n5 GND 0.03fF
C34 a_5182_210.n6 GND 0.06fF
C35 a_5182_210.n7 GND 0.03fF
C36 a_5182_210.n8 GND 0.12fF
C37 a_5182_210.n9 GND 0.06fF
C38 a_5182_210.n10 GND 0.01fF
C39 a_5182_210.t0 GND 0.33fF
C40 a_7106_210.n0 GND 0.07fF
C41 a_7106_210.n1 GND 0.09fF
C42 a_7106_210.n2 GND 0.13fF
C43 a_7106_210.n3 GND 0.11fF
C44 a_7106_210.n4 GND 0.02fF
C45 a_7106_210.n5 GND 0.03fF
C46 a_7106_210.n6 GND 0.06fF
C47 a_7106_210.n7 GND 0.03fF
C48 a_7106_210.n8 GND 0.12fF
C49 a_7106_210.n9 GND 0.06fF
C50 a_7106_210.n10 GND 0.01fF
C51 a_7106_210.t0 GND 0.33fF
C52 a_1334_210.n0 GND 0.07fF
C53 a_1334_210.n1 GND 0.09fF
C54 a_1334_210.n2 GND 0.13fF
C55 a_1334_210.n3 GND 0.11fF
C56 a_1334_210.n4 GND 0.02fF
C57 a_1334_210.n5 GND 0.03fF
C58 a_1334_210.n6 GND 0.02fF
C59 a_1334_210.n7 GND 0.05fF
C60 a_1334_210.n8 GND 0.03fF
C61 a_1334_210.n9 GND 0.11fF
C62 a_1334_210.n10 GND 0.06fF
C63 a_1334_210.n11 GND 0.01fF
C64 a_1334_210.t0 GND 0.33fF
C65 a_2015_103.n0 GND 0.09fF
C66 a_2015_103.n1 GND 0.10fF
C67 a_2015_103.n2 GND 0.05fF
C68 a_2015_103.n3 GND 0.03fF
C69 a_2015_103.n4 GND 0.04fF
C70 a_2015_103.n5 GND 0.03fF
C71 a_2015_103.n6 GND 0.04fF
C72 a_15764_210.n0 GND 0.02fF
C73 a_15764_210.n1 GND 0.09fF
C74 a_15764_210.n2 GND 0.13fF
C75 a_15764_210.n3 GND 0.11fF
C76 a_15764_210.t1 GND 0.30fF
C77 a_15764_210.n4 GND 0.09fF
C78 a_15764_210.n5 GND 0.06fF
C79 a_15764_210.n6 GND 0.01fF
C80 a_15764_210.n7 GND 0.03fF
C81 a_15764_210.n8 GND 0.11fF
C82 a_15764_210.n9 GND 0.02fF
C83 a_15764_210.n10 GND 0.05fF
C84 a_15764_210.n11 GND 0.02fF
C85 a_4220_210.n0 GND 0.02fF
C86 a_4220_210.n1 GND 0.09fF
C87 a_4220_210.n2 GND 0.13fF
C88 a_4220_210.n3 GND 0.11fF
C89 a_4220_210.t1 GND 0.30fF
C90 a_4220_210.n4 GND 0.09fF
C91 a_4220_210.n5 GND 0.06fF
C92 a_4220_210.n6 GND 0.01fF
C93 a_4220_210.n7 GND 0.03fF
C94 a_4220_210.n8 GND 0.11fF
C95 a_4220_210.n9 GND 0.02fF
C96 a_4220_210.n10 GND 0.05fF
C97 a_4220_210.n11 GND 0.03fF
C98 a_2296_210.n0 GND 0.07fF
C99 a_2296_210.n1 GND 0.09fF
C100 a_2296_210.n2 GND 0.13fF
C101 a_2296_210.n3 GND 0.11fF
C102 a_2296_210.n4 GND 0.02fF
C103 a_2296_210.n5 GND 0.03fF
C104 a_2296_210.n6 GND 0.02fF
C105 a_2296_210.n7 GND 0.05fF
C106 a_2296_210.n8 GND 0.03fF
C107 a_2296_210.n9 GND 0.11fF
C108 a_2296_210.n10 GND 0.06fF
C109 a_2296_210.n11 GND 0.01fF
C110 a_2296_210.t0 GND 0.33fF
C111 a_12878_210.n0 GND 0.02fF
C112 a_12878_210.n1 GND 0.09fF
C113 a_12878_210.n2 GND 0.13fF
C114 a_12878_210.n3 GND 0.11fF
C115 a_12878_210.t1 GND 0.30fF
C116 a_12878_210.n4 GND 0.09fF
C117 a_12878_210.n5 GND 0.06fF
C118 a_12878_210.n6 GND 0.01fF
C119 a_12878_210.n7 GND 0.03fF
C120 a_12878_210.n8 GND 0.11fF
C121 a_12878_210.n9 GND 0.02fF
C122 a_12878_210.n10 GND 0.05fF
C123 a_12878_210.n11 GND 0.02fF
C124 a_16445_103.n0 GND 0.09fF
C125 a_16445_103.n1 GND 0.10fF
C126 a_16445_103.n2 GND 0.05fF
C127 a_16445_103.n3 GND 0.03fF
C128 a_16445_103.n4 GND 0.04fF
C129 a_16445_103.n5 GND 0.03fF
C130 a_16445_103.n6 GND 0.04fF
C131 a_10954_210.n0 GND 0.07fF
C132 a_10954_210.n1 GND 0.09fF
C133 a_10954_210.n2 GND 0.13fF
C134 a_10954_210.n3 GND 0.11fF
C135 a_10954_210.n4 GND 0.02fF
C136 a_10954_210.n5 GND 0.03fF
C137 a_10954_210.n6 GND 0.06fF
C138 a_10954_210.n7 GND 0.03fF
C139 a_10954_210.n8 GND 0.12fF
C140 a_10954_210.n9 GND 0.06fF
C141 a_10954_210.n10 GND 0.01fF
C142 a_10954_210.t0 GND 0.33fF
C143 a_14802_210.n0 GND 0.07fF
C144 a_14802_210.n1 GND 0.09fF
C145 a_14802_210.n2 GND 0.13fF
C146 a_14802_210.n3 GND 0.11fF
C147 a_14802_210.n4 GND 0.02fF
C148 a_14802_210.n5 GND 0.03fF
C149 a_14802_210.n6 GND 0.06fF
C150 a_14802_210.n7 GND 0.03fF
C151 a_14802_210.n8 GND 0.12fF
C152 a_14802_210.n9 GND 0.06fF
C153 a_14802_210.n10 GND 0.01fF
C154 a_14802_210.t0 GND 0.33fF
C155 a_15483_103.n0 GND 0.09fF
C156 a_15483_103.n1 GND 0.10fF
C157 a_15483_103.n2 GND 0.05fF
C158 a_15483_103.n3 GND 0.03fF
C159 a_15483_103.n4 GND 0.04fF
C160 a_15483_103.n5 GND 0.11fF
C161 a_15483_103.n6 GND 0.04fF
C162 a_13559_103.n0 GND 0.09fF
C163 a_13559_103.n1 GND 0.10fF
C164 a_13559_103.n2 GND 0.05fF
C165 a_13559_103.n3 GND 0.03fF
C166 a_13559_103.n4 GND 0.04fF
C167 a_13559_103.n5 GND 0.03fF
C168 a_13559_103.n6 GND 0.04fF
C169 a_17428_101.n0 GND 0.11fF
C170 a_17428_101.n1 GND 0.09fF
C171 a_17428_101.n2 GND 0.08fF
C172 a_17428_101.n3 GND 0.02fF
C173 a_17428_101.n4 GND 0.01fF
C174 a_17428_101.n5 GND 0.06fF
C175 a_9992_210.n0 GND 0.02fF
C176 a_9992_210.n1 GND 0.09fF
C177 a_9992_210.n2 GND 0.13fF
C178 a_9992_210.n3 GND 0.11fF
C179 a_9992_210.t1 GND 0.30fF
C180 a_9992_210.n4 GND 0.09fF
C181 a_9992_210.n5 GND 0.06fF
C182 a_9992_210.n6 GND 0.01fF
C183 a_9992_210.n7 GND 0.03fF
C184 a_9992_210.n8 GND 0.11fF
C185 a_9992_210.n9 GND 0.02fF
C186 a_9992_210.n10 GND 0.05fF
C187 a_9992_210.n11 GND 0.02fF
C188 a_11916_210.n0 GND 0.02fF
C189 a_11916_210.n1 GND 0.09fF
C190 a_11916_210.n2 GND 0.13fF
C191 a_11916_210.n3 GND 0.11fF
C192 a_11916_210.t1 GND 0.30fF
C193 a_11916_210.n4 GND 0.09fF
C194 a_11916_210.n5 GND 0.06fF
C195 a_11916_210.n6 GND 0.01fF
C196 a_11916_210.n7 GND 0.03fF
C197 a_11916_210.n8 GND 0.11fF
C198 a_11916_210.n9 GND 0.02fF
C199 a_11916_210.n10 GND 0.05fF
C200 a_11916_210.n11 GND 0.02fF
C201 a_91_103.n0 GND 0.09fF
C202 a_91_103.n1 GND 0.09fF
C203 a_91_103.n2 GND 0.04fF
C204 a_91_103.n3 GND 0.03fF
C205 a_91_103.n4 GND 0.04fF
C206 a_91_103.n5 GND 0.03fF
C207 a_91_103.n6 GND 0.04fF
C208 a_10673_103.n0 GND 0.09fF
C209 a_10673_103.n1 GND 0.10fF
C210 a_10673_103.n2 GND 0.05fF
C211 a_10673_103.n3 GND 0.03fF
C212 a_10673_103.n4 GND 0.04fF
C213 a_10673_103.n5 GND 0.11fF
C214 a_10673_103.n6 GND 0.04fF
C215 a_14521_103.n0 GND 0.20fF
C216 a_14521_103.n1 GND 0.04fF
C217 a_14521_103.n2 GND 0.01fF
C218 a_14521_103.n3 GND 0.08fF
C219 a_14521_103.n4 GND 0.06fF
C220 a_14521_103.n5 GND 0.07fF
C221 a_12597_103.n0 GND 0.09fF
C222 a_12597_103.n1 GND 0.10fF
C223 a_12597_103.n2 GND 0.05fF
C224 a_12597_103.n3 GND 0.03fF
C225 a_12597_103.n4 GND 0.04fF
C226 a_12597_103.n5 GND 0.11fF
C227 a_12597_103.n6 GND 0.04fF
C228 a_9030_210.n0 GND 0.07fF
C229 a_9030_210.n1 GND 0.09fF
C230 a_9030_210.n2 GND 0.13fF
C231 a_9030_210.n3 GND 0.11fF
C232 a_9030_210.n4 GND 0.02fF
C233 a_9030_210.n5 GND 0.03fF
C234 a_9030_210.n6 GND 0.06fF
C235 a_9030_210.n7 GND 0.03fF
C236 a_9030_210.n8 GND 0.12fF
C237 a_9030_210.n9 GND 0.06fF
C238 a_9030_210.n10 GND 0.01fF
C239 a_9030_210.t0 GND 0.33fF
C240 a_8749_103.n0 GND 0.09fF
C241 a_8749_103.n1 GND 0.10fF
C242 a_8749_103.n2 GND 0.05fF
C243 a_8749_103.n3 GND 0.03fF
C244 a_8749_103.n4 GND 0.04fF
C245 a_8749_103.n5 GND 0.11fF
C246 a_8749_103.n6 GND 0.04fF
C247 a_372_210.n0 GND 0.02fF
C248 a_372_210.n1 GND 0.09fF
C249 a_372_210.n2 GND 0.13fF
C250 a_372_210.n3 GND 0.11fF
C251 a_372_210.t1 GND 0.30fF
C252 a_372_210.n4 GND 0.09fF
C253 a_372_210.n5 GND 0.06fF
C254 a_372_210.n6 GND 0.01fF
C255 a_372_210.n7 GND 0.03fF
C256 a_372_210.n8 GND 0.11fF
C257 a_372_210.n9 GND 0.02fF
C258 a_372_210.n10 GND 0.05fF
C259 a_372_210.n11 GND 0.03fF
C260 a_599_989.n0 GND 0.46fF
C261 a_599_989.n1 GND 0.79fF
C262 a_599_989.n2 GND 0.52fF
C263 a_599_989.t7 GND 0.74fF
C264 a_599_989.n3 GND 0.54fF
C265 a_599_989.n4 GND 3.76fF
C266 a_599_989.n5 GND 0.06fF
C267 a_599_989.n6 GND 0.07fF
C268 a_599_989.n7 GND 0.05fF
C269 a_599_989.n8 GND 0.42fF
C270 a_599_989.n9 GND 0.62fF
C271 a_599_989.n10 GND 0.74fF
C272 a_599_989.n11 GND 0.87fF
C273 a_599_989.n12 GND 0.27fF
C274 a_599_989.n13 GND 0.42fF
C275 a_599_989.n14 GND 0.74fF
C276 a_9711_103.n0 GND 0.09fF
C277 a_9711_103.n1 GND 0.10fF
C278 a_9711_103.n2 GND 0.05fF
C279 a_9711_103.n3 GND 0.03fF
C280 a_9711_103.n4 GND 0.04fF
C281 a_9711_103.n5 GND 0.11fF
C282 a_9711_103.n6 GND 0.04fF
C283 a_277_1050.n0 GND 0.54fF
C284 a_277_1050.n1 GND 0.40fF
C285 a_277_1050.n2 GND 0.49fF
C286 a_277_1050.n3 GND 0.40fF
C287 a_277_1050.n4 GND 0.47fF
C288 a_277_1050.n5 GND 1.14fF
C289 a_277_1050.n6 GND 0.34fF
C290 a_277_1050.n7 GND 0.49fF
C291 a_277_1050.n8 GND 0.37fF
C292 a_277_1050.n9 GND 0.64fF
C293 a_277_1050.n10 GND 0.20fF
C294 a_277_1050.n11 GND 0.54fF
C295 a_8068_210.n0 GND 0.07fF
C296 a_8068_210.n1 GND 0.09fF
C297 a_8068_210.n2 GND 0.13fF
C298 a_8068_210.n3 GND 0.11fF
C299 a_8068_210.n4 GND 0.02fF
C300 a_8068_210.n5 GND 0.03fF
C301 a_8068_210.n6 GND 0.06fF
C302 a_8068_210.n7 GND 0.03fF
C303 a_8068_210.n8 GND 0.12fF
C304 a_8068_210.n9 GND 0.06fF
C305 a_8068_210.n10 GND 0.01fF
C306 a_8068_210.t0 GND 0.33fF
C307 a_7787_103.n0 GND 0.09fF
C308 a_7787_103.n1 GND 0.10fF
C309 a_7787_103.n2 GND 0.05fF
C310 a_7787_103.n3 GND 0.03fF
C311 a_7787_103.n4 GND 0.04fF
C312 a_7787_103.n5 GND 0.11fF
C313 a_7787_103.n6 GND 0.04fF
C314 a_16726_210.n0 GND 0.02fF
C315 a_16726_210.n1 GND 0.09fF
C316 a_16726_210.n2 GND 0.13fF
C317 a_16726_210.n3 GND 0.11fF
C318 a_16726_210.t1 GND 0.30fF
C319 a_16726_210.n4 GND 0.09fF
C320 a_16726_210.n5 GND 0.06fF
C321 a_16726_210.n6 GND 0.01fF
C322 a_16726_210.n7 GND 0.03fF
C323 a_16726_210.n8 GND 0.11fF
C324 a_16726_210.n9 GND 0.02fF
C325 a_16726_210.n10 GND 0.05fF
C326 a_16726_210.n11 GND 0.03fF
C327 a_11635_103.n0 GND 0.09fF
C328 a_11635_103.n1 GND 0.10fF
C329 a_11635_103.n2 GND 0.05fF
C330 a_11635_103.n3 GND 0.03fF
C331 a_11635_103.n4 GND 0.04fF
C332 a_11635_103.n5 GND 0.11fF
C333 a_11635_103.n6 GND 0.04fF
C334 a_6144_210.n0 GND 0.02fF
C335 a_6144_210.n1 GND 0.09fF
C336 a_6144_210.n2 GND 0.13fF
C337 a_6144_210.n3 GND 0.11fF
C338 a_6144_210.t1 GND 0.30fF
C339 a_6144_210.n4 GND 0.09fF
C340 a_6144_210.n5 GND 0.06fF
C341 a_6144_210.n6 GND 0.01fF
C342 a_6144_210.n7 GND 0.03fF
C343 a_6144_210.n8 GND 0.11fF
C344 a_6144_210.n9 GND 0.02fF
C345 a_6144_210.n10 GND 0.05fF
C346 a_6144_210.n11 GND 0.02fF
C347 a_5863_103.n0 GND 0.09fF
C348 a_5863_103.n1 GND 0.10fF
C349 a_5863_103.n2 GND 0.05fF
C350 a_5863_103.n3 GND 0.03fF
C351 a_5863_103.n4 GND 0.04fF
C352 a_5863_103.n5 GND 0.11fF
C353 a_5863_103.n6 GND 0.04fF
C354 RN.n0 GND 0.92fF
C355 RN.t12 GND 0.84fF
C356 RN.n1 GND 0.71fF
C357 RN.n2 GND 0.90fF
C358 RN.t24 GND 0.86fF
C359 RN.n3 GND 0.69fF
C360 RN.n4 GND 3.65fF
C361 RN.n5 GND 0.92fF
C362 RN.t6 GND 0.84fF
C363 RN.n6 GND 0.69fF
C364 RN.n7 GND 3.96fF
C365 RN.n8 GND 0.92fF
C366 RN.t8 GND 0.84fF
C367 RN.n9 GND 0.69fF
C368 RN.n10 GND 2.11fF
C369 RN.n11 GND 0.90fF
C370 RN.t25 GND 0.86fF
C371 RN.n12 GND 0.69fF
C372 RN.n13 GND 3.04fF
C373 RN.n14 GND 0.92fF
C374 RN.t1 GND 0.84fF
C375 RN.n15 GND 0.69fF
C376 RN.n16 GND 3.96fF
C377 RN.n17 GND 0.92fF
C378 RN.t23 GND 0.84fF
C379 RN.n18 GND 0.69fF
C380 RN.n19 GND 2.11fF
C381 RN.n20 GND 0.90fF
C382 RN.t16 GND 0.86fF
C383 RN.n21 GND 0.69fF
C384 RN.n22 GND 3.04fF
C385 RN.n23 GND 0.92fF
C386 RN.t11 GND 0.84fF
C387 RN.n24 GND 0.69fF
C388 RN.n25 GND 2.46fF
C389 QN.n0 GND 0.42fF
C390 QN.n1 GND 0.51fF
C391 QN.n2 GND 0.25fF
C392 QN.n3 GND 0.04fF
C393 QN.n4 GND 0.05fF
C394 QN.n5 GND 0.11fF
C395 QN.n6 GND 0.04fF
C396 QN.n7 GND 0.05fF
C397 QN.n8 GND 0.03fF
C398 QN.n9 GND 0.10fF
C399 QN.n10 GND 1.08fF
C400 QN.n11 GND 0.13fF
C401 QN.n12 GND 0.32fF
C402 QN.n13 GND 0.37fF
C403 QN.n14 GND 0.01fF
C404 a_18197_1051.n0 GND 0.28fF
C405 a_18197_1051.n1 GND 0.29fF
C406 a_18197_1051.n2 GND 0.20fF
C407 a_18197_1051.n3 GND 0.56fF
C408 a_18197_1051.n4 GND 0.25fF
C409 a_18197_1051.n5 GND 0.35fF
C410 a_9897_1050.n0 GND 0.57fF
C411 a_9897_1050.n1 GND 0.57fF
C412 a_9897_1050.n2 GND 0.36fF
C413 a_9897_1050.n3 GND 0.69fF
C414 a_9897_1050.n4 GND 0.04fF
C415 a_9897_1050.n5 GND 0.06fF
C416 a_9897_1050.n6 GND 0.04fF
C417 a_9897_1050.n7 GND 0.32fF
C418 a_9897_1050.n8 GND 0.66fF
C419 a_9897_1050.n9 GND 0.32fF
C420 a_9897_1050.n10 GND 0.21fF
C421 a_9897_1050.n11 GND 0.67fF
C422 a_7973_1050.n0 GND 0.42fF
C423 a_7973_1050.n1 GND 0.67fF
C424 a_7973_1050.n2 GND 0.04fF
C425 a_7973_1050.n3 GND 0.06fF
C426 a_7973_1050.n4 GND 0.04fF
C427 a_7973_1050.n5 GND 0.25fF
C428 a_7973_1050.n6 GND 0.66fF
C429 a_7973_1050.n7 GND 0.56fF
C430 a_7973_1050.n8 GND 0.66fF
C431 a_7973_1050.n9 GND 0.21fF
C432 a_7973_1050.n10 GND 0.39fF
C433 a_7973_1050.n11 GND 0.56fF
C434 a_7333_989.n0 GND 0.95fF
C435 a_7333_989.n1 GND 0.61fF
C436 a_7333_989.t14 GND 1.00fF
C437 a_7333_989.n2 GND 0.76fF
C438 a_7333_989.n3 GND 0.61fF
C439 a_7333_989.t13 GND 1.00fF
C440 a_7333_989.n4 GND 0.66fF
C441 a_7333_989.n5 GND 0.61fF
C442 a_7333_989.t11 GND 1.00fF
C443 a_7333_989.n6 GND 0.69fF
C444 a_7333_989.n7 GND 2.24fF
C445 a_7333_989.n8 GND 3.34fF
C446 a_7333_989.n9 GND 0.77fF
C447 a_7333_989.n10 GND 0.85fF
C448 a_7333_989.n11 GND 0.49fF
C449 a_7333_989.n12 GND 1.12fF
C450 a_7333_989.n13 GND 0.35fF
C451 a_7333_989.n14 GND 0.95fF
C452 a_1561_989.n0 GND 0.88fF
C453 a_1561_989.n1 GND 0.56fF
C454 a_1561_989.t12 GND 0.92fF
C455 a_1561_989.n2 GND 0.70fF
C456 a_1561_989.n3 GND 0.56fF
C457 a_1561_989.t9 GND 0.92fF
C458 a_1561_989.n4 GND 0.61fF
C459 a_1561_989.n5 GND 0.56fF
C460 a_1561_989.t10 GND 0.92fF
C461 a_1561_989.n6 GND 0.64fF
C462 a_1561_989.n7 GND 2.06fF
C463 a_1561_989.n8 GND 3.08fF
C464 a_1561_989.n9 GND 0.70fF
C465 a_1561_989.n10 GND 0.79fF
C466 a_1561_989.n11 GND 0.45fF
C467 a_1561_989.n12 GND 1.03fF
C468 a_1561_989.n13 GND 0.32fF
C469 a_1561_989.n14 GND 0.88fF
C470 a_2201_1050.n0 GND 0.51fF
C471 a_2201_1050.n1 GND 0.38fF
C472 a_2201_1050.n2 GND 0.61fF
C473 a_2201_1050.n3 GND 0.32fF
C474 a_2201_1050.n4 GND 0.63fF
C475 a_2201_1050.n5 GND 0.35fF
C476 a_2201_1050.n6 GND 0.60fF
C477 a_2201_1050.n7 GND 0.19fF
C478 a_2201_1050.n8 GND 0.51fF
C479 a_18094_101.n0 GND 0.13fF
C480 a_18094_101.n1 GND 0.15fF
C481 a_18760_101.n0 GND 0.06fF
C482 a_18760_101.n1 GND 0.13fF
C483 a_18760_101.n2 GND 0.04fF
C484 a_4447_989.n0 GND 1.21fF
C485 a_4447_989.n1 GND 1.21fF
C486 a_4447_989.n2 GND 0.86fF
C487 a_4447_989.n3 GND 1.06fF
C488 a_4447_989.n4 GND 1.31fF
C489 a_4447_989.n5 GND 0.82fF
C490 a_4447_989.n6 GND 5.26fF
C491 a_4447_989.n7 GND 0.92fF
C492 a_4447_989.t12 GND 1.15fF
C493 a_4447_989.n8 GND 0.86fF
C494 a_4447_989.n9 GND 21.24fF
C495 a_4447_989.n10 GND 0.10fF
C496 a_4447_989.n11 GND 0.12fF
C497 a_4447_989.n12 GND 0.63fF
C498 a_4447_989.n13 GND 1.07fF
C499 a_4447_989.n14 GND 0.76fF
C500 a_4447_989.n15 GND 0.45fF
C501 a_4447_989.n16 GND 1.42fF
C502 a_6371_989.n0 GND 0.98fF
C503 a_6371_989.n1 GND 0.62fF
C504 a_6371_989.n2 GND 1.05fF
C505 a_6371_989.n3 GND 0.69fF
C506 a_6371_989.t11 GND 0.98fF
C507 a_6371_989.n4 GND 0.72fF
C508 a_6371_989.n5 GND 4.99fF
C509 a_6371_989.n6 GND 0.73fF
C510 a_6371_989.n7 GND 0.88fF
C511 a_6371_989.n8 GND 0.56fF
C512 a_6371_989.n9 GND 1.15fF
C513 a_6371_989.n10 GND 0.36fF
C514 a_6371_989.n11 GND 0.98fF
C515 SN.n0 GND 0.97fF
C516 SN.t9 GND 0.79fF
C517 SN.n1 GND 0.94fF
C518 SN.n2 GND 0.96fF
C519 SN.t11 GND 0.78fF
C520 SN.n3 GND 0.68fF
C521 SN.n4 GND 6.47fF
C522 SN.n5 GND 0.97fF
C523 SN.t8 GND 0.79fF
C524 SN.n6 GND 0.66fF
C525 SN.n7 GND 4.47fF
C526 SN.n8 GND 0.96fF
C527 SN.t3 GND 0.78fF
C528 SN.n9 GND 0.68fF
C529 SN.n10 GND 4.47fF
C530 SN.n11 GND 0.97fF
C531 SN.t17 GND 0.79fF
C532 SN.n12 GND 0.66fF
C533 SN.n13 GND 4.47fF
C534 SN.t16 GND 0.78fF
C535 SN.n14 GND 0.96fF
C536 SN.n15 GND 0.68fF
C537 SN.n16 GND 2.26fF
C538 a_4901_103.n0 GND 0.10fF
C539 a_4901_103.n1 GND 0.04fF
C540 a_4901_103.n2 GND 0.03fF
C541 a_4901_103.n3 GND 0.07fF
C542 a_4901_103.n4 GND 0.08fF
C543 a_4901_103.n5 GND 0.06fF
C544 a_4125_1050.n0 GND 0.55fF
C545 a_4125_1050.n1 GND 0.55fF
C546 a_4125_1050.n2 GND 0.64fF
C547 a_4125_1050.n3 GND 0.20fF
C548 a_4125_1050.n4 GND 0.31fF
C549 a_4125_1050.n5 GND 0.34fF
C550 a_4125_1050.n6 GND 0.67fF
C551 a_4125_1050.n7 GND 0.65fF
C552 a_4125_1050.n8 GND 0.08fF
C553 a_4125_1050.n9 GND 0.30fF
C554 a_4125_1050.n10 GND 0.05fF
C555 a_12143_989.n0 GND 0.97fF
C556 a_12143_989.n1 GND 0.61fF
C557 a_12143_989.n2 GND 1.04fF
C558 a_12143_989.n3 GND 0.68fF
C559 a_12143_989.t11 GND 0.97fF
C560 a_12143_989.n4 GND 0.71fF
C561 a_12143_989.n5 GND 4.93fF
C562 a_12143_989.n6 GND 0.07fF
C563 a_12143_989.n7 GND 0.10fF
C564 a_12143_989.n8 GND 0.06fF
C565 a_12143_989.n9 GND 0.55fF
C566 a_12143_989.n10 GND 0.81fF
C567 a_12143_989.n11 GND 0.55fF
C568 a_12143_989.n12 GND 1.14fF
C569 a_12143_989.n13 GND 0.36fF
C570 a_12143_989.n14 GND 0.97fF
C571 a_11821_1050.n0 GND 0.71fF
C572 a_11821_1050.n1 GND 0.71fF
C573 a_11821_1050.n2 GND 0.83fF
C574 a_11821_1050.n3 GND 0.26fF
C575 a_11821_1050.n4 GND 0.48fF
C576 a_11821_1050.n5 GND 0.52fF
C577 a_11821_1050.n6 GND 0.64fF
C578 a_11821_1050.n7 GND 0.52fF
C579 a_11821_1050.n8 GND 0.61fF
C580 a_11821_1050.n9 GND 1.49fF
C581 a_11821_1050.n10 GND 0.61fF
C582 a_11821_1050.n11 GND 0.11fF
C583 a_11821_1050.n12 GND 0.30fF
C584 a_11821_1050.n13 GND 0.06fF
C585 a_15669_1050.n0 GND 0.34fF
C586 a_15669_1050.n1 GND 0.65fF
C587 a_15669_1050.n2 GND 0.04fF
C588 a_15669_1050.n3 GND 0.05fF
C589 a_15669_1050.n4 GND 0.03fF
C590 a_15669_1050.n5 GND 0.30fF
C591 a_15669_1050.n6 GND 0.63fF
C592 a_15669_1050.n7 GND 0.53fF
C593 a_15669_1050.n8 GND 0.63fF
C594 a_15669_1050.n9 GND 0.20fF
C595 a_15669_1050.n10 GND 0.31fF
C596 a_15669_1050.n11 GND 0.53fF
C597 a_15991_989.n0 GND 0.29fF
C598 a_15991_989.n1 GND 0.78fF
C599 a_15991_989.n2 GND 0.26fF
C600 a_15991_989.n3 GND 0.53fF
C601 a_15991_989.n4 GND 0.55fF
C602 a_15991_989.n5 GND 0.46fF
C603 a_15991_989.t15 GND 0.51fF
C604 a_15991_989.n6 GND 0.89fF
C605 a_15991_989.n7 GND 0.04fF
C606 a_15991_989.n8 GND 0.06fF
C607 a_15991_989.n9 GND 0.04fF
C608 a_15991_989.n10 GND 0.25fF
C609 a_15991_989.n11 GND 0.81fF
C610 a_15991_989.n12 GND 0.43fF
C611 a_15991_989.n13 GND 0.57fF
C612 a_15991_989.n14 GND 0.67fF
C613 a_15991_989.n15 GND 0.21fF
C614 a_15991_989.n16 GND 0.29fF
C615 a_15991_989.n17 GND 0.57fF
C616 VDD.n0 GND 0.16fF
C617 VDD.n1 GND 0.03fF
C618 VDD.n2 GND 0.02fF
C619 VDD.n3 GND 0.05fF
C620 VDD.n4 GND 0.01fF
C621 VDD.n5 GND 0.02fF
C622 VDD.n6 GND 0.02fF
C623 VDD.n9 GND 0.02fF
C624 VDD.n10 GND 0.02fF
C625 VDD.n12 GND 0.02fF
C626 VDD.n14 GND 0.46fF
C627 VDD.n16 GND 0.03fF
C628 VDD.n17 GND 0.02fF
C629 VDD.n18 GND 0.02fF
C630 VDD.n19 GND 0.02fF
C631 VDD.n20 GND 0.04fF
C632 VDD.n21 GND 0.28fF
C633 VDD.n22 GND 0.02fF
C634 VDD.n23 GND 0.03fF
C635 VDD.n24 GND 0.28fF
C636 VDD.n25 GND 0.01fF
C637 VDD.n26 GND 0.31fF
C638 VDD.n27 GND 0.01fF
C639 VDD.n28 GND 0.03fF
C640 VDD.n29 GND 0.02fF
C641 VDD.n30 GND 0.28fF
C642 VDD.n31 GND 0.01fF
C643 VDD.n32 GND 0.02fF
C644 VDD.n33 GND 0.00fF
C645 VDD.n34 GND 0.09fF
C646 VDD.n35 GND 0.03fF
C647 VDD.n36 GND 0.31fF
C648 VDD.n37 GND 0.01fF
C649 VDD.n38 GND 0.03fF
C650 VDD.n39 GND 0.03fF
C651 VDD.n40 GND 0.28fF
C652 VDD.n41 GND 0.01fF
C653 VDD.n42 GND 0.02fF
C654 VDD.n43 GND 0.02fF
C655 VDD.n44 GND 0.28fF
C656 VDD.n45 GND 0.01fF
C657 VDD.n46 GND 0.02fF
C658 VDD.n47 GND 0.02fF
C659 VDD.n48 GND 0.28fF
C660 VDD.n49 GND 0.01fF
C661 VDD.n50 GND 0.02fF
C662 VDD.n51 GND 0.03fF
C663 VDD.n52 GND 0.02fF
C664 VDD.n53 GND 0.02fF
C665 VDD.n54 GND 0.02fF
C666 VDD.n55 GND 0.22fF
C667 VDD.n56 GND 0.04fF
C668 VDD.n57 GND 0.04fF
C669 VDD.n58 GND 0.02fF
C670 VDD.n60 GND 0.02fF
C671 VDD.n61 GND 0.02fF
C672 VDD.n62 GND 0.02fF
C673 VDD.n63 GND 0.02fF
C674 VDD.n65 GND 0.02fF
C675 VDD.n66 GND 0.02fF
C676 VDD.n67 GND 0.02fF
C677 VDD.n69 GND 0.28fF
C678 VDD.n71 GND 0.02fF
C679 VDD.n72 GND 0.02fF
C680 VDD.n73 GND 0.03fF
C681 VDD.n74 GND 0.02fF
C682 VDD.n75 GND 0.28fF
C683 VDD.n76 GND 0.01fF
C684 VDD.n77 GND 0.02fF
C685 VDD.n78 GND 0.03fF
C686 VDD.n79 GND 0.28fF
C687 VDD.n80 GND 0.01fF
C688 VDD.n81 GND 0.02fF
C689 VDD.n82 GND 0.02fF
C690 VDD.n83 GND 0.28fF
C691 VDD.n84 GND 0.01fF
C692 VDD.n85 GND 0.02fF
C693 VDD.n86 GND 0.02fF
C694 VDD.n87 GND 0.31fF
C695 VDD.n88 GND 0.01fF
C696 VDD.n89 GND 0.03fF
C697 VDD.n90 GND 0.03fF
C698 VDD.n91 GND 0.31fF
C699 VDD.n92 GND 0.01fF
C700 VDD.n93 GND 0.03fF
C701 VDD.n94 GND 0.03fF
C702 VDD.n95 GND 0.28fF
C703 VDD.n96 GND 0.01fF
C704 VDD.n97 GND 0.02fF
C705 VDD.n98 GND 0.02fF
C706 VDD.n99 GND 0.28fF
C707 VDD.n100 GND 0.01fF
C708 VDD.n101 GND 0.02fF
C709 VDD.n102 GND 0.02fF
C710 VDD.n103 GND 0.28fF
C711 VDD.n104 GND 0.01fF
C712 VDD.n105 GND 0.02fF
C713 VDD.n106 GND 0.03fF
C714 VDD.n107 GND 0.02fF
C715 VDD.n108 GND 0.02fF
C716 VDD.n109 GND 0.02fF
C717 VDD.n110 GND 0.22fF
C718 VDD.n111 GND 0.04fF
C719 VDD.n112 GND 0.03fF
C720 VDD.n113 GND 0.02fF
C721 VDD.n114 GND 0.02fF
C722 VDD.n115 GND 0.02fF
C723 VDD.n116 GND 0.03fF
C724 VDD.n117 GND 0.02fF
C725 VDD.n119 GND 0.02fF
C726 VDD.n120 GND 0.02fF
C727 VDD.n121 GND 0.02fF
C728 VDD.n123 GND 0.28fF
C729 VDD.n125 GND 0.02fF
C730 VDD.n126 GND 0.02fF
C731 VDD.n127 GND 0.03fF
C732 VDD.n128 GND 0.02fF
C733 VDD.n129 GND 0.28fF
C734 VDD.n130 GND 0.01fF
C735 VDD.n131 GND 0.02fF
C736 VDD.n132 GND 0.03fF
C737 VDD.n133 GND 0.06fF
C738 VDD.n134 GND 0.25fF
C739 VDD.n135 GND 0.01fF
C740 VDD.n136 GND 0.01fF
C741 VDD.n137 GND 0.02fF
C742 VDD.n138 GND 0.14fF
C743 VDD.n139 GND 0.17fF
C744 VDD.n140 GND 0.01fF
C745 VDD.n141 GND 0.02fF
C746 VDD.n142 GND 0.02fF
C747 VDD.n143 GND 0.11fF
C748 VDD.n144 GND 0.03fF
C749 VDD.n145 GND 0.31fF
C750 VDD.n146 GND 0.01fF
C751 VDD.n147 GND 0.02fF
C752 VDD.n148 GND 0.03fF
C753 VDD.n149 GND 0.17fF
C754 VDD.n150 GND 0.14fF
C755 VDD.n151 GND 0.01fF
C756 VDD.n152 GND 0.02fF
C757 VDD.n153 GND 0.03fF
C758 VDD.n154 GND 0.14fF
C759 VDD.n155 GND 0.16fF
C760 VDD.n156 GND 0.01fF
C761 VDD.n157 GND 0.02fF
C762 VDD.n158 GND 0.02fF
C763 VDD.n159 GND 0.06fF
C764 VDD.n160 GND 0.25fF
C765 VDD.n161 GND 0.01fF
C766 VDD.n162 GND 0.01fF
C767 VDD.n163 GND 0.02fF
C768 VDD.n164 GND 0.28fF
C769 VDD.n165 GND 0.01fF
C770 VDD.n166 GND 0.02fF
C771 VDD.n167 GND 0.03fF
C772 VDD.n168 GND 0.02fF
C773 VDD.n169 GND 0.02fF
C774 VDD.n170 GND 0.02fF
C775 VDD.n171 GND 0.26fF
C776 VDD.n172 GND 0.04fF
C777 VDD.n173 GND 0.03fF
C778 VDD.n174 GND 0.02fF
C779 VDD.n175 GND 0.02fF
C780 VDD.n176 GND 0.02fF
C781 VDD.n177 GND 0.03fF
C782 VDD.n178 GND 0.02fF
C783 VDD.n180 GND 0.02fF
C784 VDD.n181 GND 0.02fF
C785 VDD.n182 GND 0.02fF
C786 VDD.n184 GND 0.28fF
C787 VDD.n186 GND 0.02fF
C788 VDD.n187 GND 0.02fF
C789 VDD.n188 GND 0.03fF
C790 VDD.n189 GND 0.02fF
C791 VDD.n190 GND 0.28fF
C792 VDD.n191 GND 0.01fF
C793 VDD.n192 GND 0.02fF
C794 VDD.n193 GND 0.03fF
C795 VDD.n194 GND 0.28fF
C796 VDD.n195 GND 0.01fF
C797 VDD.n196 GND 0.02fF
C798 VDD.n197 GND 0.02fF
C799 VDD.n198 GND 0.22fF
C800 VDD.n199 GND 0.01fF
C801 VDD.n200 GND 0.07fF
C802 VDD.n201 GND 0.02fF
C803 VDD.n202 GND 0.14fF
C804 VDD.n203 GND 0.17fF
C805 VDD.n204 GND 0.01fF
C806 VDD.n205 GND 0.02fF
C807 VDD.n206 GND 0.02fF
C808 VDD.n207 GND 0.14fF
C809 VDD.n208 GND 0.16fF
C810 VDD.n209 GND 0.01fF
C811 VDD.n210 GND 0.11fF
C812 VDD.n211 GND 0.02fF
C813 VDD.n212 GND 0.02fF
C814 VDD.n213 GND 0.02fF
C815 VDD.n214 GND 0.18fF
C816 VDD.n215 GND 0.15fF
C817 VDD.n216 GND 0.01fF
C818 VDD.n217 GND 0.02fF
C819 VDD.n218 GND 0.03fF
C820 VDD.n219 GND 0.18fF
C821 VDD.n220 GND 0.15fF
C822 VDD.n221 GND 0.01fF
C823 VDD.n222 GND 0.02fF
C824 VDD.n223 GND 0.03fF
C825 VDD.n224 GND 0.11fF
C826 VDD.n225 GND 0.02fF
C827 VDD.n226 GND 0.14fF
C828 VDD.n227 GND 0.16fF
C829 VDD.n228 GND 0.01fF
C830 VDD.n229 GND 0.02fF
C831 VDD.n230 GND 0.02fF
C832 VDD.n231 GND 0.14fF
C833 VDD.n232 GND 0.17fF
C834 VDD.n233 GND 0.01fF
C835 VDD.n234 GND 0.02fF
C836 VDD.n235 GND 0.02fF
C837 VDD.n236 GND 0.06fF
C838 VDD.n237 GND 0.23fF
C839 VDD.n238 GND 0.01fF
C840 VDD.n239 GND 0.01fF
C841 VDD.n240 GND 0.02fF
C842 VDD.n241 GND 0.28fF
C843 VDD.n242 GND 0.01fF
C844 VDD.n243 GND 0.02fF
C845 VDD.n244 GND 0.02fF
C846 VDD.n245 GND 0.28fF
C847 VDD.n246 GND 0.01fF
C848 VDD.n247 GND 0.02fF
C849 VDD.n248 GND 0.03fF
C850 VDD.n249 GND 0.02fF
C851 VDD.n250 GND 0.02fF
C852 VDD.n251 GND 0.02fF
C853 VDD.n252 GND 0.31fF
C854 VDD.n253 GND 0.04fF
C855 VDD.n254 GND 0.03fF
C856 VDD.n255 GND 0.02fF
C857 VDD.n256 GND 0.02fF
C858 VDD.n257 GND 0.02fF
C859 VDD.n258 GND 0.03fF
C860 VDD.n259 GND 0.02fF
C861 VDD.n261 GND 0.02fF
C862 VDD.n262 GND 0.02fF
C863 VDD.n263 GND 0.02fF
C864 VDD.n265 GND 0.28fF
C865 VDD.n267 GND 0.02fF
C866 VDD.n268 GND 0.02fF
C867 VDD.n269 GND 0.03fF
C868 VDD.n270 GND 0.02fF
C869 VDD.n271 GND 0.28fF
C870 VDD.n272 GND 0.01fF
C871 VDD.n273 GND 0.02fF
C872 VDD.n274 GND 0.03fF
C873 VDD.n275 GND 0.28fF
C874 VDD.n276 GND 0.01fF
C875 VDD.n277 GND 0.02fF
C876 VDD.n278 GND 0.02fF
C877 VDD.n279 GND 0.22fF
C878 VDD.n280 GND 0.01fF
C879 VDD.n281 GND 0.07fF
C880 VDD.n282 GND 0.02fF
C881 VDD.n283 GND 0.14fF
C882 VDD.n284 GND 0.17fF
C883 VDD.n285 GND 0.01fF
C884 VDD.n286 GND 0.02fF
C885 VDD.n287 GND 0.02fF
C886 VDD.n288 GND 0.14fF
C887 VDD.n289 GND 0.16fF
C888 VDD.n290 GND 0.01fF
C889 VDD.n291 GND 0.11fF
C890 VDD.n292 GND 0.02fF
C891 VDD.n293 GND 0.02fF
C892 VDD.n294 GND 0.02fF
C893 VDD.n295 GND 0.18fF
C894 VDD.n296 GND 0.15fF
C895 VDD.n297 GND 0.01fF
C896 VDD.n298 GND 0.02fF
C897 VDD.n299 GND 0.03fF
C898 VDD.n300 GND 0.18fF
C899 VDD.n301 GND 0.15fF
C900 VDD.n302 GND 0.01fF
C901 VDD.n303 GND 0.02fF
C902 VDD.n304 GND 0.03fF
C903 VDD.n305 GND 0.11fF
C904 VDD.n306 GND 0.02fF
C905 VDD.n307 GND 0.14fF
C906 VDD.n308 GND 0.16fF
C907 VDD.n309 GND 0.01fF
C908 VDD.n310 GND 0.02fF
C909 VDD.n311 GND 0.02fF
C910 VDD.n312 GND 0.14fF
C911 VDD.n313 GND 0.17fF
C912 VDD.n314 GND 0.01fF
C913 VDD.n315 GND 0.02fF
C914 VDD.n316 GND 0.02fF
C915 VDD.n317 GND 0.06fF
C916 VDD.n318 GND 0.23fF
C917 VDD.n319 GND 0.01fF
C918 VDD.n320 GND 0.01fF
C919 VDD.n321 GND 0.02fF
C920 VDD.n322 GND 0.28fF
C921 VDD.n323 GND 0.01fF
C922 VDD.n324 GND 0.02fF
C923 VDD.n325 GND 0.02fF
C924 VDD.n326 GND 0.28fF
C925 VDD.n327 GND 0.01fF
C926 VDD.n328 GND 0.02fF
C927 VDD.n329 GND 0.03fF
C928 VDD.n330 GND 0.02fF
C929 VDD.n331 GND 0.02fF
C930 VDD.n332 GND 0.02fF
C931 VDD.n333 GND 0.31fF
C932 VDD.n334 GND 0.04fF
C933 VDD.n335 GND 0.03fF
C934 VDD.n336 GND 0.02fF
C935 VDD.n337 GND 0.02fF
C936 VDD.n338 GND 0.02fF
C937 VDD.n339 GND 0.03fF
C938 VDD.n340 GND 0.02fF
C939 VDD.n342 GND 0.02fF
C940 VDD.n343 GND 0.02fF
C941 VDD.n344 GND 0.02fF
C942 VDD.n346 GND 0.28fF
C943 VDD.n348 GND 0.02fF
C944 VDD.n349 GND 0.02fF
C945 VDD.n350 GND 0.03fF
C946 VDD.n351 GND 0.02fF
C947 VDD.n352 GND 0.28fF
C948 VDD.n353 GND 0.01fF
C949 VDD.n354 GND 0.02fF
C950 VDD.n355 GND 0.03fF
C951 VDD.n356 GND 0.28fF
C952 VDD.n357 GND 0.01fF
C953 VDD.n358 GND 0.02fF
C954 VDD.n359 GND 0.02fF
C955 VDD.n360 GND 0.22fF
C956 VDD.n361 GND 0.01fF
C957 VDD.n362 GND 0.07fF
C958 VDD.n363 GND 0.02fF
C959 VDD.n364 GND 0.14fF
C960 VDD.n365 GND 0.17fF
C961 VDD.n366 GND 0.01fF
C962 VDD.n367 GND 0.02fF
C963 VDD.n368 GND 0.02fF
C964 VDD.n369 GND 0.14fF
C965 VDD.n370 GND 0.16fF
C966 VDD.n371 GND 0.01fF
C967 VDD.n372 GND 0.11fF
C968 VDD.n373 GND 0.02fF
C969 VDD.n374 GND 0.02fF
C970 VDD.n375 GND 0.02fF
C971 VDD.n376 GND 0.18fF
C972 VDD.n377 GND 0.15fF
C973 VDD.n378 GND 0.01fF
C974 VDD.n379 GND 0.02fF
C975 VDD.n380 GND 0.03fF
C976 VDD.n381 GND 0.18fF
C977 VDD.n382 GND 0.15fF
C978 VDD.n383 GND 0.01fF
C979 VDD.n384 GND 0.02fF
C980 VDD.n385 GND 0.03fF
C981 VDD.n386 GND 0.11fF
C982 VDD.n387 GND 0.02fF
C983 VDD.n388 GND 0.14fF
C984 VDD.n389 GND 0.16fF
C985 VDD.n390 GND 0.01fF
C986 VDD.n391 GND 0.02fF
C987 VDD.n392 GND 0.02fF
C988 VDD.n393 GND 0.14fF
C989 VDD.n394 GND 0.17fF
C990 VDD.n395 GND 0.01fF
C991 VDD.n396 GND 0.02fF
C992 VDD.n397 GND 0.02fF
C993 VDD.n398 GND 0.06fF
C994 VDD.n399 GND 0.23fF
C995 VDD.n400 GND 0.01fF
C996 VDD.n401 GND 0.01fF
C997 VDD.n402 GND 0.02fF
C998 VDD.n403 GND 0.28fF
C999 VDD.n404 GND 0.01fF
C1000 VDD.n405 GND 0.02fF
C1001 VDD.n406 GND 0.02fF
C1002 VDD.n407 GND 0.28fF
C1003 VDD.n408 GND 0.01fF
C1004 VDD.n409 GND 0.02fF
C1005 VDD.n410 GND 0.03fF
C1006 VDD.n411 GND 0.02fF
C1007 VDD.n412 GND 0.02fF
C1008 VDD.n413 GND 0.02fF
C1009 VDD.n414 GND 0.31fF
C1010 VDD.n415 GND 0.04fF
C1011 VDD.n416 GND 0.03fF
C1012 VDD.n417 GND 0.02fF
C1013 VDD.n418 GND 0.02fF
C1014 VDD.n419 GND 0.02fF
C1015 VDD.n420 GND 0.03fF
C1016 VDD.n421 GND 0.02fF
C1017 VDD.n423 GND 0.02fF
C1018 VDD.n424 GND 0.02fF
C1019 VDD.n425 GND 0.02fF
C1020 VDD.n427 GND 0.28fF
C1021 VDD.n429 GND 0.02fF
C1022 VDD.n430 GND 0.02fF
C1023 VDD.n431 GND 0.03fF
C1024 VDD.n432 GND 0.02fF
C1025 VDD.n433 GND 0.28fF
C1026 VDD.n434 GND 0.01fF
C1027 VDD.n435 GND 0.02fF
C1028 VDD.n436 GND 0.03fF
C1029 VDD.n437 GND 0.28fF
C1030 VDD.n438 GND 0.01fF
C1031 VDD.n439 GND 0.02fF
C1032 VDD.n440 GND 0.02fF
C1033 VDD.n441 GND 0.22fF
C1034 VDD.n442 GND 0.01fF
C1035 VDD.n443 GND 0.07fF
C1036 VDD.n444 GND 0.02fF
C1037 VDD.n445 GND 0.14fF
C1038 VDD.n446 GND 0.17fF
C1039 VDD.n447 GND 0.01fF
C1040 VDD.n448 GND 0.02fF
C1041 VDD.n449 GND 0.02fF
C1042 VDD.n450 GND 0.14fF
C1043 VDD.n451 GND 0.16fF
C1044 VDD.n452 GND 0.01fF
C1045 VDD.n453 GND 0.11fF
C1046 VDD.n454 GND 0.02fF
C1047 VDD.n455 GND 0.02fF
C1048 VDD.n456 GND 0.02fF
C1049 VDD.n457 GND 0.18fF
C1050 VDD.n458 GND 0.15fF
C1051 VDD.n459 GND 0.01fF
C1052 VDD.n460 GND 0.02fF
C1053 VDD.n461 GND 0.03fF
C1054 VDD.n462 GND 0.18fF
C1055 VDD.n463 GND 0.15fF
C1056 VDD.n464 GND 0.01fF
C1057 VDD.n465 GND 0.02fF
C1058 VDD.n466 GND 0.03fF
C1059 VDD.n467 GND 0.11fF
C1060 VDD.n468 GND 0.02fF
C1061 VDD.n469 GND 0.14fF
C1062 VDD.n470 GND 0.16fF
C1063 VDD.n471 GND 0.01fF
C1064 VDD.n472 GND 0.02fF
C1065 VDD.n473 GND 0.02fF
C1066 VDD.n474 GND 0.14fF
C1067 VDD.n475 GND 0.17fF
C1068 VDD.n476 GND 0.01fF
C1069 VDD.n477 GND 0.02fF
C1070 VDD.n478 GND 0.02fF
C1071 VDD.n479 GND 0.06fF
C1072 VDD.n480 GND 0.23fF
C1073 VDD.n481 GND 0.01fF
C1074 VDD.n482 GND 0.01fF
C1075 VDD.n483 GND 0.02fF
C1076 VDD.n484 GND 0.28fF
C1077 VDD.n485 GND 0.01fF
C1078 VDD.n486 GND 0.02fF
C1079 VDD.n487 GND 0.02fF
C1080 VDD.n488 GND 0.28fF
C1081 VDD.n489 GND 0.01fF
C1082 VDD.n490 GND 0.02fF
C1083 VDD.n491 GND 0.03fF
C1084 VDD.n492 GND 0.02fF
C1085 VDD.n493 GND 0.02fF
C1086 VDD.n494 GND 0.02fF
C1087 VDD.n495 GND 0.31fF
C1088 VDD.n496 GND 0.04fF
C1089 VDD.n497 GND 0.03fF
C1090 VDD.n498 GND 0.02fF
C1091 VDD.n499 GND 0.02fF
C1092 VDD.n500 GND 0.02fF
C1093 VDD.n501 GND 0.03fF
C1094 VDD.n502 GND 0.02fF
C1095 VDD.n504 GND 0.02fF
C1096 VDD.n505 GND 0.02fF
C1097 VDD.n506 GND 0.02fF
C1098 VDD.n508 GND 0.28fF
C1099 VDD.n510 GND 0.02fF
C1100 VDD.n511 GND 0.02fF
C1101 VDD.n512 GND 0.03fF
C1102 VDD.n513 GND 0.02fF
C1103 VDD.n514 GND 0.28fF
C1104 VDD.n515 GND 0.01fF
C1105 VDD.n516 GND 0.02fF
C1106 VDD.n517 GND 0.03fF
C1107 VDD.n518 GND 0.28fF
C1108 VDD.n519 GND 0.01fF
C1109 VDD.n520 GND 0.02fF
C1110 VDD.n521 GND 0.02fF
C1111 VDD.n522 GND 0.22fF
C1112 VDD.n523 GND 0.01fF
C1113 VDD.n524 GND 0.07fF
C1114 VDD.n525 GND 0.02fF
C1115 VDD.n526 GND 0.14fF
C1116 VDD.n527 GND 0.17fF
C1117 VDD.n528 GND 0.01fF
C1118 VDD.n529 GND 0.02fF
C1119 VDD.n530 GND 0.02fF
C1120 VDD.n531 GND 0.14fF
C1121 VDD.n532 GND 0.16fF
C1122 VDD.n533 GND 0.01fF
C1123 VDD.n534 GND 0.11fF
C1124 VDD.n535 GND 0.02fF
C1125 VDD.n536 GND 0.02fF
C1126 VDD.n537 GND 0.02fF
C1127 VDD.n538 GND 0.18fF
C1128 VDD.n539 GND 0.15fF
C1129 VDD.n540 GND 0.01fF
C1130 VDD.n541 GND 0.02fF
C1131 VDD.n542 GND 0.03fF
C1132 VDD.n543 GND 0.18fF
C1133 VDD.n544 GND 0.15fF
C1134 VDD.n545 GND 0.01fF
C1135 VDD.n546 GND 0.02fF
C1136 VDD.n547 GND 0.03fF
C1137 VDD.n548 GND 0.11fF
C1138 VDD.n549 GND 0.02fF
C1139 VDD.n550 GND 0.14fF
C1140 VDD.n551 GND 0.16fF
C1141 VDD.n552 GND 0.01fF
C1142 VDD.n553 GND 0.02fF
C1143 VDD.n554 GND 0.02fF
C1144 VDD.n555 GND 0.14fF
C1145 VDD.n556 GND 0.17fF
C1146 VDD.n557 GND 0.01fF
C1147 VDD.n558 GND 0.02fF
C1148 VDD.n559 GND 0.02fF
C1149 VDD.n560 GND 0.06fF
C1150 VDD.n561 GND 0.23fF
C1151 VDD.n562 GND 0.01fF
C1152 VDD.n563 GND 0.01fF
C1153 VDD.n564 GND 0.02fF
C1154 VDD.n565 GND 0.28fF
C1155 VDD.n566 GND 0.01fF
C1156 VDD.n567 GND 0.02fF
C1157 VDD.n568 GND 0.02fF
C1158 VDD.n569 GND 0.28fF
C1159 VDD.n570 GND 0.01fF
C1160 VDD.n571 GND 0.02fF
C1161 VDD.n572 GND 0.03fF
C1162 VDD.n573 GND 0.02fF
C1163 VDD.n574 GND 0.02fF
C1164 VDD.n575 GND 0.02fF
C1165 VDD.n576 GND 0.31fF
C1166 VDD.n577 GND 0.04fF
C1167 VDD.n578 GND 0.03fF
C1168 VDD.n579 GND 0.02fF
C1169 VDD.n580 GND 0.02fF
C1170 VDD.n581 GND 0.02fF
C1171 VDD.n582 GND 0.03fF
C1172 VDD.n583 GND 0.02fF
C1173 VDD.n585 GND 0.02fF
C1174 VDD.n586 GND 0.02fF
C1175 VDD.n587 GND 0.02fF
C1176 VDD.n589 GND 0.28fF
C1177 VDD.n591 GND 0.02fF
C1178 VDD.n592 GND 0.02fF
C1179 VDD.n593 GND 0.03fF
C1180 VDD.n594 GND 0.02fF
C1181 VDD.n595 GND 0.28fF
C1182 VDD.n596 GND 0.01fF
C1183 VDD.n597 GND 0.02fF
C1184 VDD.n598 GND 0.03fF
C1185 VDD.n599 GND 0.28fF
C1186 VDD.n600 GND 0.01fF
C1187 VDD.n601 GND 0.02fF
C1188 VDD.n602 GND 0.02fF
C1189 VDD.n603 GND 0.22fF
C1190 VDD.n604 GND 0.01fF
C1191 VDD.n605 GND 0.07fF
C1192 VDD.n606 GND 0.02fF
C1193 VDD.n607 GND 0.14fF
C1194 VDD.n608 GND 0.17fF
C1195 VDD.n609 GND 0.01fF
C1196 VDD.n610 GND 0.02fF
C1197 VDD.n611 GND 0.02fF
C1198 VDD.n612 GND 0.14fF
C1199 VDD.n613 GND 0.16fF
C1200 VDD.n614 GND 0.01fF
C1201 VDD.n615 GND 0.11fF
C1202 VDD.n616 GND 0.02fF
C1203 VDD.n617 GND 0.02fF
C1204 VDD.n618 GND 0.02fF
C1205 VDD.n619 GND 0.18fF
C1206 VDD.n620 GND 0.15fF
C1207 VDD.n621 GND 0.01fF
C1208 VDD.n622 GND 0.02fF
C1209 VDD.n623 GND 0.03fF
C1210 VDD.n624 GND 0.18fF
C1211 VDD.n625 GND 0.15fF
C1212 VDD.n626 GND 0.01fF
C1213 VDD.n627 GND 0.02fF
C1214 VDD.n628 GND 0.03fF
C1215 VDD.n629 GND 0.11fF
C1216 VDD.n630 GND 0.02fF
C1217 VDD.n631 GND 0.14fF
C1218 VDD.n632 GND 0.16fF
C1219 VDD.n633 GND 0.01fF
C1220 VDD.n634 GND 0.02fF
C1221 VDD.n635 GND 0.02fF
C1222 VDD.n636 GND 0.14fF
C1223 VDD.n637 GND 0.17fF
C1224 VDD.n638 GND 0.01fF
C1225 VDD.n639 GND 0.02fF
C1226 VDD.n640 GND 0.02fF
C1227 VDD.n641 GND 0.06fF
C1228 VDD.n642 GND 0.23fF
C1229 VDD.n643 GND 0.01fF
C1230 VDD.n644 GND 0.01fF
C1231 VDD.n645 GND 0.02fF
C1232 VDD.n646 GND 0.28fF
C1233 VDD.n647 GND 0.01fF
C1234 VDD.n648 GND 0.02fF
C1235 VDD.n649 GND 0.02fF
C1236 VDD.n650 GND 0.28fF
C1237 VDD.n651 GND 0.01fF
C1238 VDD.n652 GND 0.02fF
C1239 VDD.n653 GND 0.03fF
C1240 VDD.n654 GND 0.02fF
C1241 VDD.n655 GND 0.02fF
C1242 VDD.n656 GND 0.02fF
C1243 VDD.n657 GND 0.31fF
C1244 VDD.n658 GND 0.04fF
C1245 VDD.n659 GND 0.03fF
C1246 VDD.n660 GND 0.02fF
C1247 VDD.n661 GND 0.02fF
C1248 VDD.n662 GND 0.02fF
C1249 VDD.n663 GND 0.03fF
C1250 VDD.n664 GND 0.02fF
C1251 VDD.n666 GND 0.02fF
C1252 VDD.n667 GND 0.02fF
C1253 VDD.n668 GND 0.02fF
C1254 VDD.n670 GND 0.28fF
C1255 VDD.n672 GND 0.02fF
C1256 VDD.n673 GND 0.02fF
C1257 VDD.n674 GND 0.03fF
C1258 VDD.n675 GND 0.02fF
C1259 VDD.n676 GND 0.28fF
C1260 VDD.n677 GND 0.01fF
C1261 VDD.n678 GND 0.02fF
C1262 VDD.n679 GND 0.03fF
C1263 VDD.n680 GND 0.28fF
C1264 VDD.n681 GND 0.01fF
C1265 VDD.n682 GND 0.02fF
C1266 VDD.n683 GND 0.02fF
C1267 VDD.n684 GND 0.22fF
C1268 VDD.n685 GND 0.01fF
C1269 VDD.n686 GND 0.07fF
C1270 VDD.n687 GND 0.02fF
C1271 VDD.n688 GND 0.14fF
C1272 VDD.n689 GND 0.17fF
C1273 VDD.n690 GND 0.01fF
C1274 VDD.n691 GND 0.02fF
C1275 VDD.n692 GND 0.02fF
C1276 VDD.n693 GND 0.14fF
C1277 VDD.n694 GND 0.16fF
C1278 VDD.n695 GND 0.01fF
C1279 VDD.n696 GND 0.11fF
C1280 VDD.n697 GND 0.02fF
C1281 VDD.n698 GND 0.02fF
C1282 VDD.n699 GND 0.02fF
C1283 VDD.n700 GND 0.18fF
C1284 VDD.n701 GND 0.15fF
C1285 VDD.n702 GND 0.01fF
C1286 VDD.n703 GND 0.02fF
C1287 VDD.n704 GND 0.03fF
C1288 VDD.n705 GND 0.18fF
C1289 VDD.n706 GND 0.15fF
C1290 VDD.n707 GND 0.01fF
C1291 VDD.n708 GND 0.02fF
C1292 VDD.n709 GND 0.03fF
C1293 VDD.n710 GND 0.11fF
C1294 VDD.n711 GND 0.02fF
C1295 VDD.n712 GND 0.14fF
C1296 VDD.n713 GND 0.16fF
C1297 VDD.n714 GND 0.01fF
C1298 VDD.n715 GND 0.02fF
C1299 VDD.n716 GND 0.02fF
C1300 VDD.n717 GND 0.14fF
C1301 VDD.n718 GND 0.17fF
C1302 VDD.n719 GND 0.01fF
C1303 VDD.n720 GND 0.02fF
C1304 VDD.n721 GND 0.02fF
C1305 VDD.n722 GND 0.06fF
C1306 VDD.n723 GND 0.23fF
C1307 VDD.n724 GND 0.01fF
C1308 VDD.n725 GND 0.01fF
C1309 VDD.n726 GND 0.02fF
C1310 VDD.n727 GND 0.28fF
C1311 VDD.n728 GND 0.01fF
C1312 VDD.n729 GND 0.02fF
C1313 VDD.n730 GND 0.02fF
C1314 VDD.n731 GND 0.28fF
C1315 VDD.n732 GND 0.01fF
C1316 VDD.n733 GND 0.02fF
C1317 VDD.n734 GND 0.03fF
C1318 VDD.n735 GND 0.02fF
C1319 VDD.n736 GND 0.02fF
C1320 VDD.n737 GND 0.02fF
C1321 VDD.n738 GND 0.31fF
C1322 VDD.n739 GND 0.04fF
C1323 VDD.n740 GND 0.03fF
C1324 VDD.n741 GND 0.02fF
C1325 VDD.n742 GND 0.02fF
C1326 VDD.n743 GND 0.02fF
C1327 VDD.n744 GND 0.03fF
C1328 VDD.n745 GND 0.02fF
C1329 VDD.n747 GND 0.02fF
C1330 VDD.n748 GND 0.02fF
C1331 VDD.n749 GND 0.02fF
C1332 VDD.n751 GND 0.28fF
C1333 VDD.n753 GND 0.02fF
C1334 VDD.n754 GND 0.02fF
C1335 VDD.n755 GND 0.03fF
C1336 VDD.n756 GND 0.02fF
C1337 VDD.n757 GND 0.28fF
C1338 VDD.n758 GND 0.01fF
C1339 VDD.n759 GND 0.02fF
C1340 VDD.n760 GND 0.03fF
C1341 VDD.n761 GND 0.28fF
C1342 VDD.n762 GND 0.01fF
C1343 VDD.n763 GND 0.02fF
C1344 VDD.n764 GND 0.02fF
C1345 VDD.n765 GND 0.22fF
C1346 VDD.n766 GND 0.01fF
C1347 VDD.n767 GND 0.07fF
C1348 VDD.n768 GND 0.02fF
C1349 VDD.n769 GND 0.14fF
C1350 VDD.n770 GND 0.17fF
C1351 VDD.n771 GND 0.01fF
C1352 VDD.n772 GND 0.02fF
C1353 VDD.n773 GND 0.02fF
C1354 VDD.n774 GND 0.14fF
C1355 VDD.n775 GND 0.16fF
C1356 VDD.n776 GND 0.01fF
C1357 VDD.n777 GND 0.11fF
C1358 VDD.n778 GND 0.02fF
C1359 VDD.n779 GND 0.02fF
C1360 VDD.n780 GND 0.02fF
C1361 VDD.n781 GND 0.18fF
C1362 VDD.n782 GND 0.15fF
C1363 VDD.n783 GND 0.01fF
C1364 VDD.n784 GND 0.02fF
C1365 VDD.n785 GND 0.03fF
C1366 VDD.n786 GND 0.18fF
C1367 VDD.n787 GND 0.15fF
C1368 VDD.n788 GND 0.01fF
C1369 VDD.n789 GND 0.02fF
C1370 VDD.n790 GND 0.03fF
C1371 VDD.n791 GND 0.11fF
C1372 VDD.n792 GND 0.02fF
C1373 VDD.n793 GND 0.14fF
C1374 VDD.n794 GND 0.16fF
C1375 VDD.n795 GND 0.01fF
C1376 VDD.n796 GND 0.02fF
C1377 VDD.n797 GND 0.02fF
C1378 VDD.n798 GND 0.14fF
C1379 VDD.n799 GND 0.17fF
C1380 VDD.n800 GND 0.01fF
C1381 VDD.n801 GND 0.02fF
C1382 VDD.n802 GND 0.02fF
C1383 VDD.n803 GND 0.06fF
C1384 VDD.n804 GND 0.23fF
C1385 VDD.n805 GND 0.01fF
C1386 VDD.n806 GND 0.01fF
C1387 VDD.n807 GND 0.02fF
C1388 VDD.n808 GND 0.28fF
C1389 VDD.n809 GND 0.01fF
C1390 VDD.n810 GND 0.02fF
C1391 VDD.n811 GND 0.02fF
C1392 VDD.n812 GND 0.02fF
C1393 VDD.n813 GND 0.02fF
C1394 VDD.n814 GND 0.02fF
C1395 VDD.n815 GND 0.31fF
C1396 VDD.n816 GND 0.04fF
C1397 VDD.n817 GND 0.03fF
C1398 VDD.n818 GND 0.02fF
C1399 VDD.n819 GND 0.02fF
C1400 VDD.n820 GND 0.02fF
C1401 VDD.n821 GND 0.03fF
C1402 VDD.n822 GND 0.02fF
C1403 VDD.n824 GND 0.02fF
C1404 VDD.n825 GND 0.02fF
C1405 VDD.n826 GND 0.02fF
C1406 VDD.n828 GND 0.28fF
C1407 VDD.n830 GND 0.02fF
C1408 VDD.n831 GND 0.02fF
C1409 VDD.n832 GND 0.03fF
C1410 VDD.n833 GND 0.02fF
C1411 VDD.n834 GND 0.28fF
C1412 VDD.n835 GND 0.01fF
C1413 VDD.n836 GND 0.02fF
C1414 VDD.n837 GND 0.02fF
C1415 VDD.n838 GND 0.02fF
C1416 VDD.n839 GND 0.02fF
C1417 VDD.n840 GND 0.02fF
C1418 VDD.n841 GND 0.20fF
C1419 VDD.n842 GND 0.03fF
C1420 VDD.n843 GND 0.02fF
C1421 VDD.n844 GND 0.02fF
C1422 VDD.n845 GND 0.02fF
C1423 VDD.n846 GND 0.03fF
C1424 VDD.n847 GND 0.02fF
C1425 VDD.n849 GND 0.02fF
C1426 VDD.n850 GND 0.02fF
C1427 VDD.n851 GND 0.02fF
C1428 VDD.n853 GND 0.46fF
C1429 VDD.n855 GND 0.03fF
C1430 VDD.n856 GND 0.04fF
C1431 VDD.n857 GND 0.28fF
C1432 VDD.n858 GND 0.02fF
C1433 VDD.n859 GND 0.03fF
C1434 VDD.n860 GND 0.03fF
C1435 VDD.n861 GND 0.28fF
C1436 VDD.n862 GND 0.01fF
C1437 VDD.n863 GND 0.02fF
C1438 VDD.n864 GND 0.02fF
C1439 VDD.n865 GND 0.06fF
C1440 VDD.n866 GND 0.23fF
C1441 VDD.n867 GND 0.01fF
C1442 VDD.n868 GND 0.01fF
C1443 VDD.n869 GND 0.02fF
C1444 VDD.n870 GND 0.14fF
C1445 VDD.n871 GND 0.17fF
C1446 VDD.n872 GND 0.01fF
C1447 VDD.n873 GND 0.02fF
C1448 VDD.n874 GND 0.02fF
C1449 VDD.n875 GND 0.11fF
C1450 VDD.n876 GND 0.02fF
C1451 VDD.n877 GND 0.14fF
C1452 VDD.n878 GND 0.16fF
C1453 VDD.n879 GND 0.01fF
C1454 VDD.n880 GND 0.02fF
C1455 VDD.n881 GND 0.02fF
C1456 VDD.n882 GND 0.18fF
C1457 VDD.n883 GND 0.15fF
C1458 VDD.n884 GND 0.01fF
C1459 VDD.n885 GND 0.02fF
C1460 VDD.n886 GND 0.03fF
C1461 VDD.n887 GND 0.18fF
C1462 VDD.n888 GND 0.15fF
C1463 VDD.n889 GND 0.01fF
C1464 VDD.n890 GND 0.02fF
C1465 VDD.n891 GND 0.03fF
C1466 VDD.n892 GND 0.14fF
C1467 VDD.n893 GND 0.16fF
C1468 VDD.n894 GND 0.01fF
C1469 VDD.n895 GND 0.11fF
C1470 VDD.n896 GND 0.02fF
C1471 VDD.n897 GND 0.02fF
C1472 VDD.n898 GND 0.02fF
C1473 VDD.n899 GND 0.14fF
C1474 VDD.n900 GND 0.17fF
C1475 VDD.n901 GND 0.01fF
C1476 VDD.n902 GND 0.02fF
C1477 VDD.n903 GND 0.02fF
C1478 VDD.n904 GND 0.22fF
C1479 VDD.n905 GND 0.01fF
C1480 VDD.n906 GND 0.07fF
C1481 VDD.n907 GND 0.02fF
C1482 VDD.n908 GND 0.28fF
C1483 VDD.n909 GND 0.01fF
C1484 VDD.n910 GND 0.02fF
C1485 VDD.n911 GND 0.02fF
C1486 VDD.n912 GND 0.28fF
C1487 VDD.n913 GND 0.01fF
C1488 VDD.n914 GND 0.02fF
C1489 VDD.n915 GND 0.03fF
C1490 VDD.n916 GND 0.02fF
C1491 VDD.n917 GND 0.02fF
C1492 VDD.n918 GND 0.02fF
C1493 VDD.n919 GND 0.02fF
C1494 VDD.n920 GND 0.02fF
C1495 VDD.n921 GND 0.02fF
C1496 VDD.n923 GND 0.02fF
C1497 VDD.n924 GND 0.02fF
C1498 VDD.n925 GND 0.02fF
C1499 VDD.n926 GND 0.02fF
C1500 VDD.n928 GND 0.04fF
C1501 VDD.n929 GND 0.02fF
C1502 VDD.n930 GND 0.31fF
C1503 VDD.n931 GND 0.04fF
C1504 VDD.n933 GND 0.28fF
C1505 VDD.n935 GND 0.02fF
C1506 VDD.n936 GND 0.02fF
C1507 VDD.n937 GND 0.03fF
C1508 VDD.n938 GND 0.02fF
C1509 VDD.n939 GND 0.28fF
C1510 VDD.n940 GND 0.01fF
C1511 VDD.n941 GND 0.02fF
C1512 VDD.n942 GND 0.03fF
C1513 VDD.n943 GND 0.28fF
C1514 VDD.n944 GND 0.01fF
C1515 VDD.n945 GND 0.02fF
C1516 VDD.n946 GND 0.02fF
C1517 VDD.n947 GND 0.06fF
C1518 VDD.n948 GND 0.23fF
C1519 VDD.n949 GND 0.01fF
C1520 VDD.n950 GND 0.01fF
C1521 VDD.n951 GND 0.02fF
C1522 VDD.n952 GND 0.14fF
C1523 VDD.n953 GND 0.17fF
C1524 VDD.n954 GND 0.01fF
C1525 VDD.n955 GND 0.02fF
C1526 VDD.n956 GND 0.02fF
C1527 VDD.n957 GND 0.11fF
C1528 VDD.n958 GND 0.02fF
C1529 VDD.n959 GND 0.14fF
C1530 VDD.n960 GND 0.16fF
C1531 VDD.n961 GND 0.01fF
C1532 VDD.n962 GND 0.02fF
C1533 VDD.n963 GND 0.02fF
C1534 VDD.n964 GND 0.18fF
C1535 VDD.n965 GND 0.15fF
C1536 VDD.n966 GND 0.01fF
C1537 VDD.n967 GND 0.02fF
C1538 VDD.n968 GND 0.03fF
C1539 VDD.n969 GND 0.18fF
C1540 VDD.n970 GND 0.15fF
C1541 VDD.n971 GND 0.01fF
C1542 VDD.n972 GND 0.02fF
C1543 VDD.n973 GND 0.03fF
C1544 VDD.n974 GND 0.14fF
C1545 VDD.n975 GND 0.16fF
C1546 VDD.n976 GND 0.01fF
C1547 VDD.n977 GND 0.11fF
C1548 VDD.n978 GND 0.02fF
C1549 VDD.n979 GND 0.02fF
C1550 VDD.n980 GND 0.02fF
C1551 VDD.n981 GND 0.14fF
C1552 VDD.n982 GND 0.17fF
C1553 VDD.n983 GND 0.01fF
C1554 VDD.n984 GND 0.02fF
C1555 VDD.n985 GND 0.02fF
C1556 VDD.n986 GND 0.22fF
C1557 VDD.n987 GND 0.01fF
C1558 VDD.n988 GND 0.07fF
C1559 VDD.n989 GND 0.02fF
C1560 VDD.n990 GND 0.28fF
C1561 VDD.n991 GND 0.01fF
C1562 VDD.n992 GND 0.02fF
C1563 VDD.n993 GND 0.02fF
C1564 VDD.n994 GND 0.28fF
C1565 VDD.n995 GND 0.01fF
C1566 VDD.n996 GND 0.02fF
C1567 VDD.n997 GND 0.03fF
C1568 VDD.n998 GND 0.02fF
C1569 VDD.n999 GND 0.02fF
C1570 VDD.n1000 GND 0.02fF
C1571 VDD.n1001 GND 0.31fF
C1572 VDD.n1002 GND 0.04fF
C1573 VDD.n1003 GND 0.03fF
C1574 VDD.n1004 GND 0.02fF
C1575 VDD.n1005 GND 0.02fF
C1576 VDD.n1006 GND 0.02fF
C1577 VDD.n1007 GND 0.03fF
C1578 VDD.n1008 GND 0.02fF
C1579 VDD.n1010 GND 0.02fF
C1580 VDD.n1011 GND 0.02fF
C1581 VDD.n1012 GND 0.02fF
C1582 VDD.n1014 GND 0.28fF
C1583 VDD.n1016 GND 0.02fF
C1584 VDD.n1017 GND 0.02fF
C1585 VDD.n1018 GND 0.03fF
C1586 VDD.n1019 GND 0.02fF
C1587 VDD.n1020 GND 0.28fF
C1588 VDD.n1021 GND 0.01fF
C1589 VDD.n1022 GND 0.02fF
C1590 VDD.n1023 GND 0.03fF
C1591 VDD.n1024 GND 0.28fF
C1592 VDD.n1025 GND 0.01fF
C1593 VDD.n1026 GND 0.02fF
C1594 VDD.n1027 GND 0.02fF
C1595 VDD.n1028 GND 0.06fF
C1596 VDD.n1029 GND 0.23fF
C1597 VDD.n1030 GND 0.01fF
C1598 VDD.n1031 GND 0.01fF
C1599 VDD.n1032 GND 0.02fF
C1600 VDD.n1033 GND 0.14fF
C1601 VDD.n1034 GND 0.17fF
C1602 VDD.n1035 GND 0.01fF
C1603 VDD.n1036 GND 0.02fF
C1604 VDD.n1037 GND 0.02fF
C1605 VDD.n1038 GND 0.11fF
C1606 VDD.n1039 GND 0.02fF
C1607 VDD.n1040 GND 0.14fF
C1608 VDD.n1041 GND 0.16fF
C1609 VDD.n1042 GND 0.01fF
C1610 VDD.n1043 GND 0.02fF
C1611 VDD.n1044 GND 0.02fF
C1612 VDD.n1045 GND 0.18fF
C1613 VDD.n1046 GND 0.15fF
C1614 VDD.n1047 GND 0.01fF
C1615 VDD.n1048 GND 0.02fF
C1616 VDD.n1049 GND 0.03fF
C1617 VDD.n1050 GND 0.18fF
C1618 VDD.n1051 GND 0.15fF
C1619 VDD.n1052 GND 0.01fF
C1620 VDD.n1053 GND 0.02fF
C1621 VDD.n1054 GND 0.03fF
C1622 VDD.n1055 GND 0.14fF
C1623 VDD.n1056 GND 0.16fF
C1624 VDD.n1057 GND 0.01fF
C1625 VDD.n1058 GND 0.11fF
C1626 VDD.n1059 GND 0.02fF
C1627 VDD.n1060 GND 0.02fF
C1628 VDD.n1061 GND 0.02fF
C1629 VDD.n1062 GND 0.14fF
C1630 VDD.n1063 GND 0.17fF
C1631 VDD.n1064 GND 0.01fF
C1632 VDD.n1065 GND 0.02fF
C1633 VDD.n1066 GND 0.02fF
C1634 VDD.n1067 GND 0.22fF
C1635 VDD.n1068 GND 0.01fF
C1636 VDD.n1069 GND 0.07fF
C1637 VDD.n1070 GND 0.02fF
C1638 VDD.n1071 GND 0.28fF
C1639 VDD.n1072 GND 0.01fF
C1640 VDD.n1073 GND 0.02fF
C1641 VDD.n1074 GND 0.02fF
C1642 VDD.n1075 GND 0.28fF
C1643 VDD.n1076 GND 0.01fF
C1644 VDD.n1077 GND 0.02fF
C1645 VDD.n1078 GND 0.03fF
C1646 VDD.n1079 GND 0.02fF
C1647 VDD.n1080 GND 0.02fF
C1648 VDD.n1081 GND 0.02fF
C1649 VDD.n1082 GND 0.31fF
C1650 VDD.n1083 GND 0.04fF
C1651 VDD.n1084 GND 0.03fF
C1652 VDD.n1085 GND 0.02fF
C1653 VDD.n1086 GND 0.02fF
C1654 VDD.n1087 GND 0.02fF
C1655 VDD.n1088 GND 0.03fF
C1656 VDD.n1089 GND 0.02fF
C1657 VDD.n1091 GND 0.02fF
C1658 VDD.n1092 GND 0.02fF
C1659 VDD.n1093 GND 0.02fF
C1660 VDD.n1095 GND 0.28fF
C1661 VDD.n1097 GND 0.02fF
C1662 VDD.n1098 GND 0.02fF
C1663 VDD.n1099 GND 0.03fF
C1664 VDD.n1100 GND 0.02fF
C1665 VDD.n1101 GND 0.28fF
C1666 VDD.n1102 GND 0.01fF
C1667 VDD.n1103 GND 0.02fF
C1668 VDD.n1104 GND 0.03fF
C1669 VDD.n1105 GND 0.28fF
C1670 VDD.n1106 GND 0.01fF
C1671 VDD.n1107 GND 0.02fF
C1672 VDD.n1108 GND 0.02fF
C1673 VDD.n1109 GND 0.06fF
C1674 VDD.n1110 GND 0.23fF
C1675 VDD.n1111 GND 0.01fF
C1676 VDD.n1112 GND 0.01fF
C1677 VDD.n1113 GND 0.02fF
C1678 VDD.n1114 GND 0.14fF
C1679 VDD.n1115 GND 0.17fF
C1680 VDD.n1116 GND 0.01fF
C1681 VDD.n1117 GND 0.02fF
C1682 VDD.n1118 GND 0.02fF
C1683 VDD.n1119 GND 0.11fF
C1684 VDD.n1120 GND 0.02fF
C1685 VDD.n1121 GND 0.14fF
C1686 VDD.n1122 GND 0.16fF
C1687 VDD.n1123 GND 0.01fF
C1688 VDD.n1124 GND 0.02fF
C1689 VDD.n1125 GND 0.02fF
C1690 VDD.n1126 GND 0.18fF
C1691 VDD.n1127 GND 0.15fF
C1692 VDD.n1128 GND 0.01fF
C1693 VDD.n1129 GND 0.02fF
C1694 VDD.n1130 GND 0.03fF
C1695 VDD.n1131 GND 0.18fF
C1696 VDD.n1132 GND 0.15fF
C1697 VDD.n1133 GND 0.01fF
C1698 VDD.n1134 GND 0.02fF
C1699 VDD.n1135 GND 0.03fF
C1700 VDD.n1136 GND 0.14fF
C1701 VDD.n1137 GND 0.16fF
C1702 VDD.n1138 GND 0.01fF
C1703 VDD.n1139 GND 0.11fF
C1704 VDD.n1140 GND 0.02fF
C1705 VDD.n1141 GND 0.02fF
C1706 VDD.n1142 GND 0.02fF
C1707 VDD.n1143 GND 0.14fF
C1708 VDD.n1144 GND 0.17fF
C1709 VDD.n1145 GND 0.01fF
C1710 VDD.n1146 GND 0.02fF
C1711 VDD.n1147 GND 0.02fF
C1712 VDD.n1148 GND 0.22fF
C1713 VDD.n1149 GND 0.01fF
C1714 VDD.n1150 GND 0.07fF
C1715 VDD.n1151 GND 0.02fF
C1716 VDD.n1152 GND 0.28fF
C1717 VDD.n1153 GND 0.01fF
C1718 VDD.n1154 GND 0.02fF
C1719 VDD.n1155 GND 0.02fF
C1720 VDD.n1156 GND 0.28fF
C1721 VDD.n1157 GND 0.01fF
C1722 VDD.n1158 GND 0.02fF
C1723 VDD.n1159 GND 0.03fF
C1724 VDD.n1160 GND 0.02fF
C1725 VDD.n1161 GND 0.02fF
C1726 VDD.n1162 GND 0.02fF
C1727 VDD.n1163 GND 0.31fF
C1728 VDD.n1164 GND 0.04fF
C1729 VDD.n1165 GND 0.03fF
C1730 VDD.n1166 GND 0.02fF
C1731 VDD.n1167 GND 0.02fF
C1732 VDD.n1168 GND 0.02fF
C1733 VDD.n1169 GND 0.03fF
C1734 VDD.n1170 GND 0.02fF
C1735 VDD.n1172 GND 0.02fF
C1736 VDD.n1173 GND 0.02fF
C1737 VDD.n1174 GND 0.02fF
C1738 VDD.n1176 GND 0.28fF
C1739 VDD.n1178 GND 0.02fF
C1740 VDD.n1179 GND 0.02fF
C1741 VDD.n1180 GND 0.03fF
C1742 VDD.n1181 GND 0.02fF
C1743 VDD.n1182 GND 0.28fF
C1744 VDD.n1183 GND 0.01fF
C1745 VDD.n1184 GND 0.02fF
C1746 VDD.n1185 GND 0.03fF
C1747 VDD.n1186 GND 0.28fF
C1748 VDD.n1187 GND 0.01fF
C1749 VDD.n1188 GND 0.02fF
C1750 VDD.n1189 GND 0.02fF
C1751 VDD.n1190 GND 0.06fF
C1752 VDD.n1191 GND 0.23fF
C1753 VDD.n1192 GND 0.01fF
C1754 VDD.n1193 GND 0.01fF
C1755 VDD.n1194 GND 0.02fF
C1756 VDD.n1195 GND 0.14fF
C1757 VDD.n1196 GND 0.17fF
C1758 VDD.n1197 GND 0.01fF
C1759 VDD.n1198 GND 0.02fF
C1760 VDD.n1199 GND 0.02fF
C1761 VDD.n1200 GND 0.11fF
C1762 VDD.n1201 GND 0.02fF
C1763 VDD.n1202 GND 0.14fF
C1764 VDD.n1203 GND 0.16fF
C1765 VDD.n1204 GND 0.01fF
C1766 VDD.n1205 GND 0.02fF
C1767 VDD.n1206 GND 0.02fF
C1768 VDD.n1207 GND 0.18fF
C1769 VDD.n1208 GND 0.15fF
C1770 VDD.n1209 GND 0.01fF
C1771 VDD.n1210 GND 0.02fF
C1772 VDD.n1211 GND 0.03fF
C1773 VDD.n1212 GND 0.18fF
C1774 VDD.n1213 GND 0.15fF
C1775 VDD.n1214 GND 0.01fF
C1776 VDD.n1215 GND 0.02fF
C1777 VDD.n1216 GND 0.03fF
C1778 VDD.n1217 GND 0.14fF
C1779 VDD.n1218 GND 0.16fF
C1780 VDD.n1219 GND 0.01fF
C1781 VDD.n1220 GND 0.11fF
C1782 VDD.n1221 GND 0.02fF
C1783 VDD.n1222 GND 0.02fF
C1784 VDD.n1223 GND 0.02fF
C1785 VDD.n1224 GND 0.14fF
C1786 VDD.n1225 GND 0.17fF
C1787 VDD.n1226 GND 0.01fF
C1788 VDD.n1227 GND 0.02fF
C1789 VDD.n1228 GND 0.02fF
C1790 VDD.n1229 GND 0.22fF
C1791 VDD.n1230 GND 0.01fF
C1792 VDD.n1231 GND 0.07fF
C1793 VDD.n1232 GND 0.02fF
C1794 VDD.n1233 GND 0.28fF
C1795 VDD.n1234 GND 0.01fF
C1796 VDD.n1235 GND 0.02fF
C1797 VDD.n1236 GND 0.02fF
C1798 VDD.n1237 GND 0.28fF
C1799 VDD.n1238 GND 0.01fF
C1800 VDD.n1239 GND 0.02fF
C1801 VDD.n1240 GND 0.03fF
C1802 VDD.n1241 GND 0.02fF
C1803 VDD.n1242 GND 0.02fF
C1804 VDD.n1243 GND 0.02fF
C1805 VDD.n1244 GND 0.31fF
C1806 VDD.n1245 GND 0.04fF
C1807 VDD.n1246 GND 0.03fF
C1808 VDD.n1247 GND 0.02fF
C1809 VDD.n1248 GND 0.02fF
C1810 VDD.n1249 GND 0.02fF
C1811 VDD.n1250 GND 0.03fF
C1812 VDD.n1251 GND 0.02fF
C1813 VDD.n1253 GND 0.02fF
C1814 VDD.n1254 GND 0.02fF
C1815 VDD.n1255 GND 0.02fF
C1816 VDD.n1257 GND 0.28fF
C1817 VDD.n1259 GND 0.02fF
C1818 VDD.n1260 GND 0.02fF
C1819 VDD.n1261 GND 0.03fF
C1820 VDD.n1262 GND 0.02fF
C1821 VDD.n1263 GND 0.28fF
C1822 VDD.n1264 GND 0.01fF
C1823 VDD.n1265 GND 0.02fF
C1824 VDD.n1266 GND 0.03fF
C1825 VDD.n1267 GND 0.28fF
C1826 VDD.n1268 GND 0.01fF
C1827 VDD.n1269 GND 0.02fF
C1828 VDD.n1270 GND 0.02fF
C1829 VDD.n1271 GND 0.06fF
C1830 VDD.n1272 GND 0.23fF
C1831 VDD.n1273 GND 0.01fF
C1832 VDD.n1274 GND 0.01fF
C1833 VDD.n1275 GND 0.02fF
C1834 VDD.n1276 GND 0.14fF
C1835 VDD.n1277 GND 0.17fF
C1836 VDD.n1278 GND 0.01fF
C1837 VDD.n1279 GND 0.02fF
C1838 VDD.n1280 GND 0.02fF
C1839 VDD.n1281 GND 0.11fF
C1840 VDD.n1282 GND 0.02fF
C1841 VDD.n1283 GND 0.14fF
C1842 VDD.n1284 GND 0.16fF
C1843 VDD.n1285 GND 0.01fF
C1844 VDD.n1286 GND 0.02fF
C1845 VDD.n1287 GND 0.02fF
C1846 VDD.n1288 GND 0.18fF
C1847 VDD.n1289 GND 0.15fF
C1848 VDD.n1290 GND 0.01fF
C1849 VDD.n1291 GND 0.02fF
C1850 VDD.n1292 GND 0.03fF
C1851 VDD.n1293 GND 0.18fF
C1852 VDD.n1294 GND 0.15fF
C1853 VDD.n1295 GND 0.01fF
C1854 VDD.n1296 GND 0.02fF
C1855 VDD.n1297 GND 0.03fF
C1856 VDD.n1298 GND 0.14fF
C1857 VDD.n1299 GND 0.16fF
C1858 VDD.n1300 GND 0.01fF
C1859 VDD.n1301 GND 0.11fF
C1860 VDD.n1302 GND 0.02fF
C1861 VDD.n1303 GND 0.02fF
C1862 VDD.n1304 GND 0.02fF
C1863 VDD.n1305 GND 0.14fF
C1864 VDD.n1306 GND 0.17fF
C1865 VDD.n1307 GND 0.01fF
C1866 VDD.n1308 GND 0.02fF
C1867 VDD.n1309 GND 0.02fF
C1868 VDD.n1310 GND 0.22fF
C1869 VDD.n1311 GND 0.01fF
C1870 VDD.n1312 GND 0.07fF
C1871 VDD.n1313 GND 0.02fF
C1872 VDD.n1314 GND 0.28fF
C1873 VDD.n1315 GND 0.01fF
C1874 VDD.n1316 GND 0.02fF
C1875 VDD.n1317 GND 0.02fF
C1876 VDD.n1318 GND 0.28fF
C1877 VDD.n1319 GND 0.01fF
C1878 VDD.n1320 GND 0.02fF
C1879 VDD.n1321 GND 0.03fF
C1880 VDD.n1322 GND 0.02fF
C1881 VDD.n1323 GND 0.02fF
C1882 VDD.n1324 GND 0.02fF
C1883 VDD.n1325 GND 0.31fF
C1884 VDD.n1326 GND 0.04fF
C1885 VDD.n1327 GND 0.03fF
C1886 VDD.n1328 GND 0.02fF
C1887 VDD.n1329 GND 0.02fF
C1888 VDD.n1330 GND 0.02fF
C1889 VDD.n1331 GND 0.03fF
C1890 VDD.n1332 GND 0.02fF
C1891 VDD.n1334 GND 0.02fF
C1892 VDD.n1335 GND 0.02fF
C1893 VDD.n1336 GND 0.02fF
C1894 VDD.n1338 GND 0.28fF
C1895 VDD.n1340 GND 0.02fF
C1896 VDD.n1341 GND 0.02fF
C1897 VDD.n1342 GND 0.03fF
C1898 VDD.n1343 GND 0.02fF
C1899 VDD.n1344 GND 0.28fF
C1900 VDD.n1345 GND 0.01fF
C1901 VDD.n1346 GND 0.02fF
C1902 VDD.n1347 GND 0.03fF
C1903 VDD.n1348 GND 0.28fF
C1904 VDD.n1349 GND 0.01fF
C1905 VDD.n1350 GND 0.02fF
C1906 VDD.n1351 GND 0.02fF
C1907 VDD.n1352 GND 0.06fF
C1908 VDD.n1353 GND 0.23fF
C1909 VDD.n1354 GND 0.01fF
C1910 VDD.n1355 GND 0.01fF
C1911 VDD.n1356 GND 0.02fF
C1912 VDD.n1357 GND 0.14fF
C1913 VDD.n1358 GND 0.17fF
C1914 VDD.n1359 GND 0.01fF
C1915 VDD.n1360 GND 0.02fF
C1916 VDD.n1361 GND 0.02fF
C1917 VDD.n1362 GND 0.11fF
C1918 VDD.n1363 GND 0.02fF
C1919 VDD.n1364 GND 0.14fF
C1920 VDD.n1365 GND 0.16fF
C1921 VDD.n1366 GND 0.01fF
C1922 VDD.n1367 GND 0.02fF
C1923 VDD.n1368 GND 0.02fF
C1924 VDD.n1369 GND 0.18fF
C1925 VDD.n1370 GND 0.15fF
C1926 VDD.n1371 GND 0.01fF
C1927 VDD.n1372 GND 0.02fF
C1928 VDD.n1373 GND 0.03fF
C1929 VDD.n1374 GND 0.18fF
C1930 VDD.n1375 GND 0.15fF
C1931 VDD.n1376 GND 0.01fF
C1932 VDD.n1377 GND 0.02fF
C1933 VDD.n1378 GND 0.03fF
C1934 VDD.n1379 GND 0.14fF
C1935 VDD.n1380 GND 0.16fF
C1936 VDD.n1381 GND 0.01fF
C1937 VDD.n1382 GND 0.11fF
C1938 VDD.n1383 GND 0.02fF
C1939 VDD.n1384 GND 0.02fF
C1940 VDD.n1385 GND 0.02fF
C1941 VDD.n1386 GND 0.14fF
C1942 VDD.n1387 GND 0.17fF
C1943 VDD.n1388 GND 0.01fF
C1944 VDD.n1389 GND 0.02fF
C1945 VDD.n1390 GND 0.02fF
C1946 VDD.n1391 GND 0.22fF
C1947 VDD.n1392 GND 0.01fF
C1948 VDD.n1393 GND 0.07fF
C1949 VDD.n1394 GND 0.02fF
C1950 VDD.n1395 GND 0.28fF
C1951 VDD.n1396 GND 0.01fF
C1952 VDD.n1397 GND 0.02fF
C1953 VDD.n1398 GND 0.02fF
C1954 VDD.n1399 GND 0.28fF
C1955 VDD.n1400 GND 0.01fF
C1956 VDD.n1401 GND 0.02fF
C1957 VDD.n1402 GND 0.03fF
C1958 VDD.n1403 GND 0.02fF
C1959 VDD.n1404 GND 0.02fF
C1960 VDD.n1405 GND 0.02fF
C1961 VDD.n1406 GND 0.31fF
C1962 VDD.n1407 GND 0.04fF
C1963 VDD.n1408 GND 0.03fF
C1964 VDD.n1409 GND 0.02fF
C1965 VDD.n1410 GND 0.02fF
C1966 VDD.n1411 GND 0.02fF
C1967 VDD.n1412 GND 0.03fF
C1968 VDD.n1413 GND 0.02fF
C1969 VDD.n1415 GND 0.02fF
C1970 VDD.n1416 GND 0.02fF
C1971 VDD.n1417 GND 0.02fF
C1972 VDD.n1419 GND 0.28fF
C1973 VDD.n1421 GND 0.02fF
C1974 VDD.n1422 GND 0.02fF
C1975 VDD.n1423 GND 0.03fF
C1976 VDD.n1424 GND 0.02fF
C1977 VDD.n1425 GND 0.28fF
C1978 VDD.n1426 GND 0.01fF
C1979 VDD.n1427 GND 0.02fF
C1980 VDD.n1428 GND 0.03fF
C1981 VDD.n1429 GND 0.28fF
C1982 VDD.n1430 GND 0.01fF
C1983 VDD.n1431 GND 0.02fF
C1984 VDD.n1432 GND 0.02fF
C1985 VDD.n1433 GND 0.06fF
C1986 VDD.n1434 GND 0.23fF
C1987 VDD.n1435 GND 0.01fF
C1988 VDD.n1436 GND 0.01fF
C1989 VDD.n1437 GND 0.02fF
C1990 VDD.n1438 GND 0.14fF
C1991 VDD.n1439 GND 0.17fF
C1992 VDD.n1440 GND 0.01fF
C1993 VDD.n1441 GND 0.02fF
C1994 VDD.n1442 GND 0.02fF
C1995 VDD.n1443 GND 0.11fF
C1996 VDD.n1444 GND 0.02fF
C1997 VDD.n1445 GND 0.14fF
C1998 VDD.n1446 GND 0.16fF
C1999 VDD.n1447 GND 0.01fF
C2000 VDD.n1448 GND 0.02fF
C2001 VDD.n1449 GND 0.02fF
C2002 VDD.n1450 GND 0.18fF
C2003 VDD.n1451 GND 0.15fF
C2004 VDD.n1452 GND 0.01fF
C2005 VDD.n1453 GND 0.02fF
C2006 VDD.n1454 GND 0.03fF
C2007 VDD.n1455 GND 0.18fF
C2008 VDD.n1456 GND 0.15fF
C2009 VDD.n1457 GND 0.01fF
C2010 VDD.n1458 GND 0.02fF
C2011 VDD.n1459 GND 0.03fF
C2012 VDD.n1460 GND 0.14fF
C2013 VDD.n1461 GND 0.16fF
C2014 VDD.n1462 GND 0.01fF
C2015 VDD.n1463 GND 0.11fF
C2016 VDD.n1464 GND 0.02fF
C2017 VDD.n1465 GND 0.02fF
C2018 VDD.n1466 GND 0.02fF
C2019 VDD.n1467 GND 0.14fF
C2020 VDD.n1468 GND 0.17fF
C2021 VDD.n1469 GND 0.01fF
C2022 VDD.n1470 GND 0.02fF
C2023 VDD.n1471 GND 0.02fF
C2024 VDD.n1472 GND 0.22fF
C2025 VDD.n1473 GND 0.01fF
C2026 VDD.n1474 GND 0.07fF
C2027 VDD.n1475 GND 0.02fF
C2028 VDD.n1476 GND 0.28fF
C2029 VDD.n1477 GND 0.01fF
C2030 VDD.n1478 GND 0.02fF
C2031 VDD.n1479 GND 0.02fF
C2032 VDD.n1480 GND 0.28fF
C2033 VDD.n1481 GND 0.01fF
C2034 VDD.n1482 GND 0.02fF
C2035 VDD.n1483 GND 0.03fF
C2036 VDD.n1484 GND 0.02fF
C2037 VDD.n1485 GND 0.02fF
C2038 VDD.n1486 GND 0.02fF
C2039 VDD.n1487 GND 0.31fF
C2040 VDD.n1488 GND 0.04fF
C2041 VDD.n1489 GND 0.03fF
C2042 VDD.n1490 GND 0.02fF
C2043 VDD.n1491 GND 0.02fF
C2044 VDD.n1492 GND 0.02fF
C2045 VDD.n1493 GND 0.03fF
C2046 VDD.n1494 GND 0.02fF
C2047 VDD.n1496 GND 0.02fF
C2048 VDD.n1497 GND 0.02fF
C2049 VDD.n1498 GND 0.02fF
C2050 VDD.n1500 GND 0.28fF
C2051 VDD.n1502 GND 0.02fF
C2052 VDD.n1503 GND 0.02fF
C2053 VDD.n1504 GND 0.03fF
C2054 VDD.n1505 GND 0.02fF
C2055 VDD.n1506 GND 0.28fF
C2056 VDD.n1507 GND 0.01fF
C2057 VDD.n1508 GND 0.02fF
C2058 VDD.n1509 GND 0.03fF
C2059 VDD.n1510 GND 0.28fF
C2060 VDD.n1511 GND 0.01fF
C2061 VDD.n1512 GND 0.02fF
C2062 VDD.n1513 GND 0.02fF
C2063 VDD.n1514 GND 0.06fF
C2064 VDD.n1515 GND 0.23fF
C2065 VDD.n1516 GND 0.01fF
C2066 VDD.n1517 GND 0.01fF
C2067 VDD.n1518 GND 0.02fF
C2068 VDD.n1519 GND 0.14fF
C2069 VDD.n1520 GND 0.17fF
C2070 VDD.n1521 GND 0.01fF
C2071 VDD.n1522 GND 0.02fF
C2072 VDD.n1523 GND 0.02fF
C2073 VDD.n1524 GND 0.11fF
C2074 VDD.n1525 GND 0.02fF
C2075 VDD.n1526 GND 0.14fF
C2076 VDD.n1527 GND 0.16fF
C2077 VDD.n1528 GND 0.01fF
C2078 VDD.n1529 GND 0.02fF
C2079 VDD.n1530 GND 0.02fF
C2080 VDD.n1531 GND 0.18fF
C2081 VDD.n1532 GND 0.15fF
C2082 VDD.n1533 GND 0.01fF
C2083 VDD.n1534 GND 0.02fF
C2084 VDD.n1535 GND 0.03fF
C2085 VDD.n1536 GND 0.18fF
C2086 VDD.n1537 GND 0.15fF
C2087 VDD.n1538 GND 0.01fF
C2088 VDD.n1539 GND 0.02fF
C2089 VDD.n1540 GND 0.03fF
C2090 VDD.n1541 GND 0.14fF
C2091 VDD.n1542 GND 0.16fF
C2092 VDD.n1543 GND 0.01fF
C2093 VDD.n1544 GND 0.11fF
C2094 VDD.n1545 GND 0.02fF
C2095 VDD.n1546 GND 0.02fF
C2096 VDD.n1547 GND 0.02fF
C2097 VDD.n1548 GND 0.14fF
C2098 VDD.n1549 GND 0.17fF
C2099 VDD.n1550 GND 0.01fF
C2100 VDD.n1551 GND 0.02fF
C2101 VDD.n1552 GND 0.02fF
C2102 VDD.n1553 GND 0.22fF
C2103 VDD.n1554 GND 0.01fF
C2104 VDD.n1555 GND 0.07fF
C2105 VDD.n1556 GND 0.02fF
C2106 VDD.n1557 GND 0.28fF
C2107 VDD.n1558 GND 0.01fF
C2108 VDD.n1559 GND 0.02fF
C2109 VDD.n1560 GND 0.02fF
C2110 VDD.n1561 GND 0.28fF
C2111 VDD.n1562 GND 0.01fF
C2112 VDD.n1563 GND 0.02fF
C2113 VDD.n1564 GND 0.03fF
C2114 VDD.n1565 GND 0.02fF
C2115 VDD.n1566 GND 0.02fF
C2116 VDD.n1567 GND 0.02fF
C2117 VDD.n1568 GND 0.31fF
C2118 VDD.n1569 GND 0.04fF
C2119 VDD.n1570 GND 0.03fF
C2120 VDD.n1571 GND 0.02fF
C2121 VDD.n1572 GND 0.02fF
C2122 VDD.n1573 GND 0.02fF
C2123 VDD.n1574 GND 0.03fF
C2124 VDD.n1575 GND 0.02fF
C2125 VDD.n1577 GND 0.02fF
C2126 VDD.n1578 GND 0.02fF
C2127 VDD.n1579 GND 0.02fF
C2128 VDD.n1581 GND 0.28fF
C2129 VDD.n1583 GND 0.02fF
C2130 VDD.n1584 GND 0.02fF
C2131 VDD.n1585 GND 0.03fF
C2132 VDD.n1586 GND 0.02fF
C2133 VDD.n1587 GND 0.28fF
C2134 VDD.n1588 GND 0.01fF
C2135 VDD.n1589 GND 0.02fF
C2136 VDD.n1590 GND 0.03fF
C2137 VDD.n1591 GND 0.28fF
C2138 VDD.n1592 GND 0.01fF
C2139 VDD.n1593 GND 0.02fF
C2140 VDD.n1594 GND 0.02fF
C2141 VDD.n1595 GND 0.06fF
C2142 VDD.n1596 GND 0.23fF
C2143 VDD.n1597 GND 0.01fF
C2144 VDD.n1598 GND 0.01fF
C2145 VDD.n1599 GND 0.02fF
C2146 VDD.n1600 GND 0.14fF
C2147 VDD.n1601 GND 0.17fF
C2148 VDD.n1602 GND 0.01fF
C2149 VDD.n1603 GND 0.02fF
C2150 VDD.n1604 GND 0.02fF
C2151 VDD.n1605 GND 0.11fF
C2152 VDD.n1606 GND 0.02fF
C2153 VDD.n1607 GND 0.14fF
C2154 VDD.n1608 GND 0.16fF
C2155 VDD.n1609 GND 0.01fF
C2156 VDD.n1610 GND 0.02fF
C2157 VDD.n1611 GND 0.02fF
C2158 VDD.n1612 GND 0.18fF
C2159 VDD.n1613 GND 0.15fF
C2160 VDD.n1614 GND 0.01fF
C2161 VDD.n1615 GND 0.02fF
C2162 VDD.n1616 GND 0.03fF
C2163 VDD.n1617 GND 0.18fF
C2164 VDD.n1618 GND 0.15fF
C2165 VDD.n1619 GND 0.01fF
C2166 VDD.n1620 GND 0.02fF
C2167 VDD.n1621 GND 0.03fF
C2168 VDD.n1622 GND 0.14fF
C2169 VDD.n1623 GND 0.16fF
C2170 VDD.n1624 GND 0.01fF
C2171 VDD.n1625 GND 0.11fF
C2172 VDD.n1626 GND 0.02fF
C2173 VDD.n1627 GND 0.02fF
C2174 VDD.n1628 GND 0.02fF
C2175 VDD.n1629 GND 0.14fF
C2176 VDD.n1630 GND 0.17fF
C2177 VDD.n1631 GND 0.01fF
C2178 VDD.n1632 GND 0.02fF
C2179 VDD.n1633 GND 0.02fF
C2180 VDD.n1634 GND 0.22fF
C2181 VDD.n1635 GND 0.01fF
C2182 VDD.n1636 GND 0.07fF
C2183 VDD.n1637 GND 0.02fF
C2184 VDD.n1638 GND 0.28fF
C2185 VDD.n1639 GND 0.01fF
C2186 VDD.n1640 GND 0.02fF
C2187 VDD.n1641 GND 0.02fF
C2188 VDD.n1642 GND 0.28fF
C2189 VDD.n1643 GND 0.01fF
C2190 VDD.n1644 GND 0.02fF
C2191 VDD.n1645 GND 0.03fF
C2192 a_17533_1051.n0 GND 0.37fF
C2193 a_17533_1051.n1 GND 0.41fF
C2194 a_17533_1051.n2 GND 0.28fF
C2195 a_17533_1051.n3 GND 0.63fF
C2196 a_17533_1051.n4 GND 0.23fF
C2197 a_17533_1051.n5 GND 0.33fF
C2198 a_10219_989.n0 GND 0.99fF
C2199 a_10219_989.n1 GND 0.99fF
C2200 a_10219_989.n2 GND 1.16fF
C2201 a_10219_989.n3 GND 0.37fF
C2202 a_10219_989.n4 GND 0.51fF
C2203 a_10219_989.n5 GND 0.57fF
C2204 a_10219_989.n6 GND 0.81fF
C2205 a_10219_989.n7 GND 0.51fF
C2206 a_10219_989.n8 GND 0.70fF
C2207 a_10219_989.n9 GND 10.47fF
C2208 a_10219_989.n10 GND 1.61fF
C2209 a_10219_989.n11 GND 0.80fF
C2210 a_10219_989.t15 GND 0.88fF
C2211 a_10219_989.n12 GND 1.55fF
C2212 a_10219_989.n13 GND 1.42fF
C2213 a_10219_989.n14 GND 0.15fF
C2214 a_10219_989.n15 GND 0.42fF
C2215 a_10219_989.n16 GND 0.08fF
C2216 a_6825_103.n0 GND 0.03fF
C2217 a_6825_103.n1 GND 0.10fF
C2218 a_6825_103.n2 GND 0.10fF
C2219 a_6825_103.n3 GND 0.05fF
C2220 a_6825_103.n4 GND 0.03fF
C2221 a_6825_103.n5 GND 0.04fF
C2222 a_6825_103.n6 GND 0.11fF
C2223 a_6825_103.n7 GND 0.04fF
C2224 a_6049_1050.n0 GND 0.71fF
C2225 a_6049_1050.n1 GND 0.71fF
C2226 a_6049_1050.n2 GND 0.83fF
C2227 a_6049_1050.n3 GND 0.26fF
C2228 a_6049_1050.n4 GND 0.48fF
C2229 a_6049_1050.n5 GND 0.52fF
C2230 a_6049_1050.n6 GND 0.64fF
C2231 a_6049_1050.n7 GND 0.52fF
C2232 a_6049_1050.n8 GND 0.61fF
C2233 a_6049_1050.n9 GND 1.49fF
C2234 a_6049_1050.n10 GND 0.61fF
C2235 a_6049_1050.n11 GND 0.11fF
C2236 a_6049_1050.n12 GND 0.30fF
C2237 a_6049_1050.n13 GND 0.06fF
C2238 a_13745_1050.n0 GND 0.56fF
C2239 a_13745_1050.n1 GND 0.56fF
C2240 a_13745_1050.n2 GND 0.66fF
C2241 a_13745_1050.n3 GND 0.21fF
C2242 a_13745_1050.n4 GND 0.39fF
C2243 a_13745_1050.n5 GND 0.42fF
C2244 a_13745_1050.n6 GND 0.67fF
C2245 a_13745_1050.n7 GND 0.67fF
C2246 a_13745_1050.n8 GND 0.09fF
C2247 a_13745_1050.n9 GND 0.24fF
C2248 a_13745_1050.n10 GND 0.05fF
C2249 a_13840_210.n0 GND 0.07fF
C2250 a_13840_210.n1 GND 0.13fF
C2251 a_13840_210.n2 GND 0.07fF
C2252 a_13840_210.n3 GND 0.02fF
C2253 a_13840_210.n4 GND 0.03fF
C2254 a_13840_210.n5 GND 0.06fF
C2255 a_13840_210.n6 GND 0.05fF
C2256 a_13840_210.n7 GND 0.06fF
C2257 a_13840_210.n8 GND 0.07fF
C2258 a_13840_210.n9 GND 0.07fF
C2259 a_13840_210.n10 GND 0.03fF
C2260 a_13840_210.n11 GND 0.01fF
C2261 a_13840_210.n12 GND 0.12fF
C2262 a_13840_210.t0 GND 0.28fF
C2263 a_13105_989.n0 GND 0.90fF
C2264 a_13105_989.n1 GND 0.90fF
C2265 a_13105_989.n2 GND 1.05fF
C2266 a_13105_989.n3 GND 0.33fF
C2267 a_13105_989.n4 GND 0.46fF
C2268 a_13105_989.n5 GND 0.58fF
C2269 a_13105_989.t8 GND 0.94fF
C2270 a_13105_989.n6 GND 0.72fF
C2271 a_13105_989.n7 GND 0.58fF
C2272 a_13105_989.t7 GND 0.94fF
C2273 a_13105_989.n8 GND 0.62fF
C2274 a_13105_989.n9 GND 0.57fF
C2275 a_13105_989.t15 GND 0.94fF
C2276 a_13105_989.n10 GND 0.65fF
C2277 a_13105_989.n11 GND 2.11fF
C2278 a_13105_989.n12 GND 3.15fF
C2279 a_13105_989.n13 GND 0.77fF
C2280 a_13105_989.n14 GND 0.14fF
C2281 a_13105_989.n15 GND 0.54fF
C2282 a_13105_989.n16 GND 0.08fF
C2283 a_3258_210.n0 GND 0.07fF
C2284 a_3258_210.n1 GND 0.13fF
C2285 a_3258_210.n2 GND 0.07fF
C2286 a_3258_210.n3 GND 0.02fF
C2287 a_3258_210.n4 GND 0.03fF
C2288 a_3258_210.n5 GND 0.06fF
C2289 a_3258_210.n6 GND 0.05fF
C2290 a_3258_210.n7 GND 0.06fF
C2291 a_3258_210.n8 GND 0.07fF
C2292 a_3258_210.n9 GND 0.07fF
C2293 a_3258_210.n10 GND 0.03fF
C2294 a_3258_210.n11 GND 0.01fF
C2295 a_3258_210.n12 GND 0.12fF
C2296 a_3258_210.t0 GND 0.28fF
C2297 a_2977_103.n0 GND 0.03fF
C2298 a_2977_103.n1 GND 0.10fF
C2299 a_2977_103.n2 GND 0.10fF
C2300 a_2977_103.n3 GND 0.05fF
C2301 a_2977_103.n4 GND 0.03fF
C2302 a_2977_103.n5 GND 0.04fF
C2303 a_2977_103.n6 GND 0.11fF
C2304 a_2977_103.n7 GND 0.04fF
.ends
