* SPICE3 file created from DFFSNRNQX1.ext - technology: sky130A

.subckt DFFSNRNQX1 Q D CLK SN RN VDD GND
X0 li1_M1_contact_8/VSUBS D nand3x1_pcell_0/nmos_bottom_0/a_0_0# li1_M1_contact_8/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15
X1 m1_831_576# m1_716_723# nand3x1_pcell_0/li_393_182# li1_M1_contact_8/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15
X2 nand3x1_pcell_0/li_393_182# RN nand3x1_pcell_0/nmos_bottom_0/a_0_0# li1_M1_contact_8/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15

X3 VDD D m1_831_576# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X4 m1_831_576# D VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X5 VDD RN m1_831_576# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X6 m1_831_576# RN VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X7 VDD m1_716_723# m1_831_576# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X8 m1_831_576# m1_716_723# VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X9 GND m1_831_576# nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 w=3 l=0.15
X10 m1_716_723# m1_1660_797# nand3x1_pcell_1/li_393_182# GND sky130_fd_pr__nfet_01v8 w=3 l=0.15
X11 nand3x1_pcell_1/li_393_182# CLK nand3x1_pcell_1/nmos_bottom_0/a_0_0# GND sky130_fd_pr__nfet_01v8 w=3 l=0.15

X12 VDD m1_831_576# m1_716_723# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X13 m1_716_723# m1_831_576# VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X14 VDD CLK m1_716_723# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X15 m1_716_723# CLK VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X16 VDD m1_1660_797# m1_716_723# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X17 m1_716_723# m1_1660_797# VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X18 li1_M1_contact_9/VSUBS m1_831_576# nand3x1_pcell_2/nmos_bottom_0/a_0_0# li1_M1_contact_9/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15
X19 m1_2757_575# m1_1660_797# nand3x1_pcell_2/li_393_182# li1_M1_contact_9/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15
X20 nand3x1_pcell_2/li_393_182# SN nand3x1_pcell_2/nmos_bottom_0/a_0_0# li1_M1_contact_9/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15

X21 VDD m1_831_576# m1_2757_575# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X22 m1_2757_575# m1_831_576# VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X23 VDD SN m1_2757_575# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X24 m1_2757_575# SN VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X25 VDD m1_1660_797# m1_2757_575# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X26 m1_2757_575# m1_1660_797# VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X27 li1_M1_contact_9/VSUBS m1_2757_575# nand3x1_pcell_3/nmos_bottom_0/a_0_0# li1_M1_contact_9/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15
X28 m1_1660_797# RN nand3x1_pcell_3/li_393_182# li1_M1_contact_9/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15
X29 nand3x1_pcell_3/li_393_182# CLK nand3x1_pcell_3/nmos_bottom_0/a_0_0# li1_M1_contact_9/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15

X30 VDD m1_2757_575# m1_1660_797# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X31 m1_1660_797# m1_2757_575# VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X32 VDD CLK m1_1660_797# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X33 m1_1660_797# CLK VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X34 VDD RN m1_1660_797# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X35 m1_1660_797# RN VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X36 li1_M1_contact_23/VSUBS m1_716_723# nand3x1_pcell_4/nmos_bottom_0/a_0_0# li1_M1_contact_23/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15
X37 m1_4645_649# Q nand3x1_pcell_4/li_393_182# li1_M1_contact_23/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15
X38 nand3x1_pcell_4/li_393_182# RN nand3x1_pcell_4/nmos_bottom_0/a_0_0# li1_M1_contact_23/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15

X39 VDD m1_716_723# m1_4645_649# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X40 m1_4645_649# m1_716_723# VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X41 VDD RN m1_4645_649# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X42 m1_4645_649# RN VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X43 VDD Q m1_4645_649# VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X44 m1_4645_649# Q VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X45 nand3x1_pcell_5/pmos2_2/VSUBS m1_4645_649# nand3x1_pcell_5/nmos_bottom_0/a_0_0# nand3x1_pcell_5/pmos2_2/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15
X46 Q m1_1660_797# nand3x1_pcell_5/li_393_182# nand3x1_pcell_5/pmos2_2/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15
X47 nand3x1_pcell_5/li_393_182# SN nand3x1_pcell_5/nmos_bottom_0/a_0_0# nand3x1_pcell_5/pmos2_2/VSUBS sky130_fd_pr__nfet_01v8 w=3 l=0.15

X48 VDD m1_4645_649# Q VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X49 Q m1_4645_649# VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X50 VDD SN Q VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X51 Q SN VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

X52 VDD m1_1660_797# Q VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15
X53 Q m1_1660_797# VDD VDD sky130_fd_pr__pfet_01v8 w=2 l=0.15

C0 m1_1660_797# VDD 2.59fF
C1 m1_1660_797# m1_716_723# 3.20fF
C2 m1_716_723# CLK 2.42fF
C3 m1_1660_797# RN 3.42fF
C4 VDD RN 2.48fF
.ends
