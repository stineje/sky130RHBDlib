* SPICE3 file created from INVX1.ext - technology: sky130A

.subckt INVX1 Y A VDD GND
X0 Y A GND GND nshort w=3 l=0.15
X1 VDD A Y VDD pshort w=2 l=0.15 M=2
.ends
