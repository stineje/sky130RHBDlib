* SPICE3 file created from BUFX1.ext - technology: sky130A

.subckt BUFX1 Y A VDD GND
X0 bufx1_0/m1_315_501# A GND GND nshort w=3 l=0.15
X1 VDD A bufx1_0/m1_315_501# VDD pshort w=2 l=0.15
X2 Y bufx1_0/m1_315_501# GND GND nshort w=3 l=0.15
X3 VDD bufx1_0/m1_315_501# Y VDD pshort w=2 l=0.15
C0 VDD GND 2.67fF
.ends
