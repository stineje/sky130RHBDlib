// File: nand3x1_pcell.spi.pex
// Created: Tue Oct 15 15:57:52 2024
// Program "Calibre xRC"
// Version "v2023.2_27.15"
// Nominal Temperature: 30C
// Circuit Temperature: 30C
// 
simulator lang=spectre
subckt PM_NAND3X1_PCELL\%noxref_2 ( 9 16 23 33 41 54 61 62 63 64 )
c47 ( 64 0 ) capacitor c=0.0455453f //x=3.585 //y=5.02
c48 ( 63 0 ) capacitor c=0.0244794f //x=2.705 //y=5.02
c49 ( 62 0 ) capacitor c=0.0244794f //x=1.825 //y=5.02
c50 ( 61 0 ) capacitor c=0.0533644f //x=0.955 //y=5.02
c51 ( 60 0 ) capacitor c=0.00591168f //x=3.73 //y=7.4
c52 ( 59 0 ) capacitor c=0.00591168f //x=2.85 //y=7.4
c53 ( 58 0 ) capacitor c=0.00591168f //x=1.97 //y=7.4
c54 ( 57 0 ) capacitor c=0.00591168f //x=1.09 //y=7.4
c55 ( 54 0 ) capacitor c=0.272255f //x=4.07 //y=7.4
c56 ( 41 0 ) capacitor c=0.028513f //x=3.645 //y=7.4
c57 ( 33 0 ) capacitor c=0.0287069f //x=2.765 //y=7.4
c58 ( 23 0 ) capacitor c=0.0292055f //x=1.885 //y=7.4
c59 ( 16 0 ) capacitor c=0.235022f //x=0.74 //y=7.4
c60 ( 13 0 ) capacitor c=0.0452081f //x=1.005 //y=7.4
c61 ( 9 0 ) capacitor c=0.214792f //x=4.07 //y=7.4
r62 (  52 60 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=3.73 //y2=7.4
r63 (  52 54 ) resistor r=9.14286 //w=0.357 //l=0.255 //layer=li \
 //thickness=0.1 //x=3.815 //y=7.4 //x2=4.07 //y2=7.4
r64 (  45 60 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=3.73 //y=7.23 //x2=3.73 //y2=7.4
r65 (  45 64 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.73 //y=7.23 //x2=3.73 //y2=6.745
r66 (  42 59 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.85 //y2=7.4
r67 (  42 44 ) resistor r=0.896359 //w=0.357 //l=0.025 //layer=li \
 //thickness=0.1 //x=2.935 //y=7.4 //x2=2.96 //y2=7.4
r68 (  41 60 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=3.73 //y2=7.4
r69 (  41 44 ) resistor r=24.5602 //w=0.357 //l=0.685 //layer=li \
 //thickness=0.1 //x=3.645 //y=7.4 //x2=2.96 //y2=7.4
r70 (  35 59 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=2.85 //y=7.23 //x2=2.85 //y2=7.4
r71 (  35 63 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.85 //y=7.23 //x2=2.85 //y2=6.745
r72 (  34 58 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.055 //y=7.4 //x2=1.97 //y2=7.4
r73 (  33 59 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.85 //y2=7.4
r74 (  33 34 ) resistor r=25.4566 //w=0.357 //l=0.71 //layer=li \
 //thickness=0.1 //x=2.765 //y=7.4 //x2=2.055 //y2=7.4
r75 (  27 58 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.97 //y=7.23 //x2=1.97 //y2=7.4
r76 (  27 62 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.97 //y=7.23 //x2=1.97 //y2=6.745
r77 (  24 57 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.09 //y2=7.4
r78 (  24 26 ) resistor r=24.2017 //w=0.357 //l=0.675 //layer=li \
 //thickness=0.1 //x=1.175 //y=7.4 //x2=1.85 //y2=7.4
r79 (  23 58 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.97 //y2=7.4
r80 (  23 26 ) resistor r=1.2549 //w=0.357 //l=0.035 //layer=li \
 //thickness=0.1 //x=1.885 //y=7.4 //x2=1.85 //y2=7.4
r81 (  17 57 ) resistor r=4.11603 //w=0.68 //l=0.17 //layer=li //thickness=0.1 \
 //x=1.09 //y=7.23 //x2=1.09 //y2=7.4
r82 (  17 61 ) resistor r=56.4706 //w=0.187 //l=0.825 //layer=li \
 //thickness=0.1 //x=1.09 //y=7.23 //x2=1.09 //y2=6.405
r83 (  13 57 ) resistor r=2.94794 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=1.09 //y2=7.4
r84 (  13 16 ) resistor r=9.5014 //w=0.357 //l=0.265 //layer=li \
 //thickness=0.1 //x=1.005 //y=7.4 //x2=0.74 //y2=7.4
r85 (  9 54 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=4.07 \
 //y=7.4 //x2=4.07 //y2=7.4
r86 (  7 44 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=2.96 \
 //y=7.4 //x2=2.96 //y2=7.4
r87 (  7 9 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=2.96 //y=7.4 //x2=4.07 //y2=7.4
r88 (  5 26 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=1.85 \
 //y=7.4 //x2=1.85 //y2=7.4
r89 (  5 7 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=1.85 //y=7.4 //x2=2.96 //y2=7.4
r90 (  2 16 ) resistor r=3.1 //w=0.17 //l=0.51 //layer=mcon //count=3 //x=0.74 \
 //y=7.4 //x2=0.74 //y2=7.4
r91 (  2 5 ) resistor r=0.460963 //w=0.301 //l=1.11 //layer=m1 \
 //thickness=0.36 //x=0.74 //y=7.4 //x2=1.85 //y2=7.4
ends PM_NAND3X1_PCELL\%noxref_2

subckt PM_NAND3X1_PCELL\%noxref_3 ( 2 7 8 9 10 11 12 13 14 16 22 23 24 25 )
c52 ( 25 0 ) capacitor c=0.0598646f //x=1.385 //y=4.79
c53 ( 24 0 ) capacitor c=0.0375015f //x=1.675 //y=4.79
c54 ( 23 0 ) capacitor c=0.0347816f //x=1.34 //y=1.22
c55 ( 22 0 ) capacitor c=0.0187487f //x=1.34 //y=0.875
c56 ( 16 0 ) capacitor c=0.0137055f //x=1.185 //y=1.375
c57 ( 14 0 ) capacitor c=0.0149861f //x=1.185 //y=0.72
c58 ( 13 0 ) capacitor c=0.102158f //x=0.81 //y=1.915
c59 ( 12 0 ) capacitor c=0.0229444f //x=0.81 //y=1.53
c60 ( 11 0 ) capacitor c=0.0234352f //x=0.81 //y=1.22
c61 ( 10 0 ) capacitor c=0.0198724f //x=0.81 //y=0.875
c62 ( 9 0 ) capacitor c=0.110114f //x=1.75 //y=6.02
c63 ( 8 0 ) capacitor c=0.158956f //x=1.31 //y=6.02
c64 ( 2 0 ) capacitor c=0.128848f //x=1.11 //y=2.08
r65 (  24 26 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.75 //y2=4.865
r66 (  24 25 ) resistor r=148.702 //w=0.094 //l=0.29 //layer=ply \
 //thickness=0.18 //x=1.675 //y=4.79 //x2=1.385 //y2=4.79
r67 (  23 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=1.22 //x2=1.3 //y2=1.375
r68 (  22 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.3 //y2=0.72
r69 (  22 23 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=1.34 //y=0.875 //x2=1.34 //y2=1.22
r70 (  19 25 ) resistor r=22.7971 //w=0.269 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.385 //y2=4.79
r71 (  19 34 ) resistor r=35.8364 //w=0.269 //l=0.270185 //layer=ply \
 //thickness=0.18 //x=1.31 //y=4.865 //x2=1.11 //y2=4.7
r72 (  17 30 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=1.375 //x2=0.85 //y2=1.375
r73 (  16 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=1.375 //x2=1.3 //y2=1.375
r74 (  15 29 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=0.965 //y=0.72 //x2=0.85 //y2=0.72
r75 (  14 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=1.3 //y2=0.72
r76 (  14 15 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=1.185 //y=0.72 //x2=0.965 //y2=0.72
r77 (  13 32 ) resistor r=58.7805 //w=0.246 //l=0.373497 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.915 //x2=1.11 //y2=2.08
r78 (  12 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.85 //y2=1.375
r79 (  12 13 ) resistor r=197.415 //w=0.094 //l=0.385 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.53 //x2=0.81 //y2=1.915
r80 (  11 30 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=1.22 //x2=0.85 //y2=1.375
r81 (  10 29 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.85 //y2=0.72
r82 (  10 11 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=0.81 //y=0.875 //x2=0.81 //y2=1.22
r83 (  9 26 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.75 //y=6.02 //x2=1.75 //y2=4.865
r84 (  8 19 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=1.31 //y=6.02 //x2=1.31 //y2=4.865
r85 (  7 16 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=1.185 //y2=1.375
r86 (  7 17 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=1.075 //y=1.375 //x2=0.965 //y2=1.375
r87 (  5 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=4.7 //x2=1.11 //y2=4.7
r88 (  2 32 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=2.08
r89 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=1.11 //y=2.08 //x2=1.11 //y2=4.7
ends PM_NAND3X1_PCELL\%noxref_3

subckt PM_NAND3X1_PCELL\%noxref_4 ( 2 7 8 9 10 11 12 14 20 21 22 23 24 32 )
c69 ( 32 0 ) capacitor c=0.0354872f //x=2.22 //y=4.7
c70 ( 24 0 ) capacitor c=0.0307682f //x=2.555 //y=4.79
c71 ( 23 0 ) capacitor c=0.0850619f //x=2.31 //y=1.915
c72 ( 22 0 ) capacitor c=0.0170266f //x=2.31 //y=1.45
c73 ( 21 0 ) capacitor c=0.018609f //x=2.31 //y=1.22
c74 ( 20 0 ) capacitor c=0.0187309f //x=2.31 //y=0.91
c75 ( 14 0 ) capacitor c=0.014725f //x=2.155 //y=1.375
c76 ( 12 0 ) capacitor c=0.0146567f //x=2.155 //y=0.755
c77 ( 11 0 ) capacitor c=0.0335408f //x=1.785 //y=1.22
c78 ( 10 0 ) capacitor c=0.0173761f //x=1.785 //y=0.91
c79 ( 9 0 ) capacitor c=0.110114f //x=2.63 //y=6.02
c80 ( 8 0 ) capacitor c=0.11012f //x=2.19 //y=6.02
c81 ( 2 0 ) capacitor c=0.106919f //x=2.22 //y=2.08
r82 (  34 35 ) resistor r=32.4568 //w=0.214 //l=0.075 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.79 //x2=2.22 //y2=4.865
r83 (  32 34 ) resistor r=20.271 //w=0.214 //l=0.09 //layer=ply \
 //thickness=0.18 //x=2.22 //y=4.7 //x2=2.22 //y2=4.79
r84 (  25 34 ) resistor r=16.5046 //w=0.27 //l=0.135 //layer=ply \
 //thickness=0.18 //x=2.355 //y=4.79 //x2=2.22 //y2=4.79
r85 (  24 26 ) resistor r=26.9307 //w=0.15 //l=0.106066 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.63 //y2=4.865
r86 (  24 25 ) resistor r=102.553 //w=0.094 //l=0.2 //layer=ply \
 //thickness=0.18 //x=2.555 //y=4.79 //x2=2.355 //y2=4.79
r87 (  23 39 ) resistor r=38.6777 //w=0.284 //l=0.198997 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.915 //x2=2.235 //y2=2.08
r88 (  22 37 ) resistor r=21.2976 //w=0.217 //l=0.0928709 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.27 //y2=1.375
r89 (  22 23 ) resistor r=238.436 //w=0.094 //l=0.465 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.45 //x2=2.31 //y2=1.915
r90 (  21 37 ) resistor r=39.0671 //w=0.217 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=1.22 //x2=2.27 //y2=1.375
r91 (  20 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.27 //y2=0.755
r92 (  20 21 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=2.31 //y=0.91 //x2=2.31 //y2=1.22
r93 (  15 30 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=1.375 //x2=1.825 //y2=1.375
r94 (  14 37 ) resistor r=11.4558 //w=0.217 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=1.375 //x2=2.27 //y2=1.375
r95 (  13 29 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=1.94 //y=0.755 //x2=1.825 //y2=0.755
r96 (  12 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=2.27 //y2=0.755
r97 (  12 13 ) resistor r=110.245 //w=0.094 //l=0.215 //layer=ply \
 //thickness=0.18 //x=2.155 //y=0.755 //x2=1.94 //y2=0.755
r98 (  11 30 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=1.22 //x2=1.825 //y2=1.375
r99 (  10 29 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.825 //y2=0.755
r100 (  10 11 ) resistor r=158.957 //w=0.094 //l=0.31 //layer=ply \
 //thickness=0.18 //x=1.785 //y=0.91 //x2=1.785 //y2=1.22
r101 (  9 26 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.63 //y=6.02 //x2=2.63 //y2=4.865
r102 (  8 35 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=2.19 //y=6.02 //x2=2.19 //y2=4.865
r103 (  7 14 ) resistor r=55.3787 //w=0.094 //l=0.108 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=2.155 //y2=1.375
r104 (  7 15 ) resistor r=54.866 //w=0.094 //l=0.107 //layer=ply \
 //thickness=0.18 //x=2.047 //y=1.375 //x2=1.94 //y2=1.375
r105 (  5 32 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=4.7 //x2=2.22 //y2=4.7
r106 (  2 39 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=2.08
r107 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=2.22 //y=2.08 //x2=2.22 //y2=4.7
ends PM_NAND3X1_PCELL\%noxref_4

subckt PM_NAND3X1_PCELL\%noxref_5 ( 1 5 9 13 17 35 )
c31 ( 35 0 ) capacitor c=0.0747858f //x=0.455 //y=0.375
c32 ( 17 0 ) capacitor c=0.0266691f //x=2.445 //y=1.59
c33 ( 13 0 ) capacitor c=0.0156939f //x=2.445 //y=0.54
c34 ( 9 0 ) capacitor c=0.00678203f //x=1.56 //y=0.625
c35 ( 5 0 ) capacitor c=0.0236189f //x=1.475 //y=1.59
c36 ( 1 0 ) capacitor c=0.0109947f //x=0.59 //y=1.505
r37 (  18 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=1.59 //x2=1.56 //y2=1.63
r38 (  18 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=1.59 //x2=2.045 //y2=1.59
r39 (  17 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=1.59 //x2=2.53 //y2=1.59
r40 (  17 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=1.59 //x2=2.045 //y2=1.59
r41 (  14 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.645 //y=0.54 //x2=1.56 //y2=0.5
r42 (  14 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.645 //y=0.54 //x2=2.045 //y2=0.54
r43 (  13 35 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.445 //y=0.54 //x2=2.53 //y2=0.54
r44 (  13 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=2.445 //y=0.54 //x2=2.045 //y2=0.54
r45 (  10 35 ) resistor r=1.40859 //w=0.34 //l=0.125 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=1.63
r46 (  10 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=1.56 //y=1.505 //x2=1.56 //y2=0.89
r47 (  9 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.5
r48 (  9 35 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=1.56 //y=0.625 //x2=1.56 //y2=0.89
r49 (  6 35 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=0.675 //y=1.59 //x2=0.59 //y2=1.63
r50 (  6 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=0.675 //y=1.59 //x2=1.075 //y2=1.59
r51 (  5 35 ) resistor r=5.4201 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=1.475 //y=1.59 //x2=1.56 //y2=1.63
r52 (  5 35 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=1.475 //y=1.59 //x2=1.075 //y2=1.59
r53 (  1 35 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=0.59 //y=1.505 //x2=0.59 //y2=1.63
r54 (  1 35 ) resistor r=42.0963 //w=0.187 //l=0.615 //layer=li \
 //thickness=0.1 //x=0.59 //y=1.505 //x2=0.59 //y2=0.89
ends PM_NAND3X1_PCELL\%noxref_5

subckt PM_NAND3X1_PCELL\%noxref_6 ( 2 7 8 9 13 14 15 20 22 25 26 28 29 34 )
c52 ( 34 0 ) capacitor c=0.0672371f //x=3.33 //y=4.7
c53 ( 29 0 ) capacitor c=0.0273931f //x=3.33 //y=1.915
c54 ( 28 0 ) capacitor c=0.0471168f //x=3.33 //y=2.08
c55 ( 26 0 ) capacitor c=0.0432517f //x=3.85 //y=1.26
c56 ( 25 0 ) capacitor c=0.0200379f //x=3.85 //y=0.915
c57 ( 22 0 ) capacitor c=0.0158629f //x=3.695 //y=1.415
c58 ( 20 0 ) capacitor c=0.0157803f //x=3.695 //y=0.76
c59 ( 15 0 ) capacitor c=0.0218028f //x=3.32 //y=1.57
c60 ( 14 0 ) capacitor c=0.0207459f //x=3.32 //y=1.26
c61 ( 13 0 ) capacitor c=0.0194308f //x=3.32 //y=0.915
c62 ( 9 0 ) capacitor c=0.158794f //x=3.51 //y=6.02
c63 ( 8 0 ) capacitor c=0.110114f //x=3.07 //y=6.02
c64 ( 2 0 ) capacitor c=0.096694f //x=3.33 //y=2.08
r65 (  28 29 ) resistor r=52.7279 //w=0.214 //l=0.165 //layer=ply \
 //thickness=0.18 //x=3.33 //y=2.08 //x2=3.33 //y2=1.915
r66 (  26 36 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=1.26 //x2=3.81 //y2=1.415
r67 (  25 35 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.81 //y2=0.76
r68 (  25 26 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.85 //y=0.915 //x2=3.85 //y2=1.26
r69 (  23 32 ) resistor r=10.701 //w=0.21 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=1.415 //x2=3.36 //y2=1.415
r70 (  22 36 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=1.415 //x2=3.81 //y2=1.415
r71 (  21 31 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.475 //y=0.76 //x2=3.36 //y2=0.76
r72 (  20 35 ) resistor r=5.52526 //w=0.168 //l=0.115 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.81 //y2=0.76
r73 (  20 21 ) resistor r=112.809 //w=0.094 //l=0.22 //layer=ply \
 //thickness=0.18 //x=3.695 //y=0.76 //x2=3.475 //y2=0.76
r74 (  17 34 ) resistor r=37.236 //w=0.233 //l=0.249199 //layer=ply \
 //thickness=0.18 //x=3.51 //y=4.865 //x2=3.33 //y2=4.7
r75 (  15 32 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.36 //y2=1.415
r76 (  15 29 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.57 //x2=3.32 //y2=1.915
r77 (  14 32 ) resistor r=39.5823 //w=0.21 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=1.26 //x2=3.36 //y2=1.415
r78 (  13 31 ) resistor r=45.1352 //w=0.168 //l=0.173853 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.36 //y2=0.76
r79 (  13 14 ) resistor r=176.904 //w=0.094 //l=0.345 //layer=ply \
 //thickness=0.18 //x=3.32 //y=0.915 //x2=3.32 //y2=1.26
r80 (  10 34 ) resistor r=53.7854 //w=0.233 //l=0.332415 //layer=ply \
 //thickness=0.18 //x=3.07 //y=4.865 //x2=3.33 //y2=4.7
r81 (  9 17 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.51 //y=6.02 //x2=3.51 //y2=4.865
r82 (  8 10 ) resistor r=592.245 //w=0.094 //l=1.155 //layer=ply \
 //thickness=0.18 //x=3.07 //y=6.02 //x2=3.07 //y2=4.865
r83 (  7 22 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.695 //y2=1.415
r84 (  7 23 ) resistor r=56.4043 //w=0.094 //l=0.11 //layer=ply \
 //thickness=0.18 //x=3.585 //y=1.415 //x2=3.475 //y2=1.415
r85 (  5 34 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=4.7 //x2=3.33 //y2=4.7
r86 (  2 28 ) resistor r=152 //w=0.17 //l=0.17 //layer=licon //count=1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=2.08
r87 (  2 5 ) resistor r=179.337 //w=0.187 //l=2.62 //layer=li //thickness=0.1 \
 //x=3.33 //y=2.08 //x2=3.33 //y2=4.7
ends PM_NAND3X1_PCELL\%noxref_6

subckt PM_NAND3X1_PCELL\%noxref_7 ( 7 8 15 23 29 30 32 33 34 35 37 38 39 )
c69 ( 39 0 ) capacitor c=0.023087f //x=3.145 //y=5.02
c70 ( 38 0 ) capacitor c=0.023519f //x=2.265 //y=5.02
c71 ( 37 0 ) capacitor c=0.0224735f //x=1.385 //y=5.02
c72 ( 35 0 ) capacitor c=0.00853354f //x=3.395 //y=0.915
c73 ( 34 0 ) capacitor c=0.0019954f //x=3.29 //y=5.155
c74 ( 33 0 ) capacitor c=0.00424403f //x=2.41 //y=5.155
c75 ( 32 0 ) capacitor c=0.135127f //x=4.07 //y=5.07
c76 ( 30 0 ) capacitor c=0.00777616f //x=3.67 //y=1.665
c77 ( 29 0 ) capacitor c=0.0191287f //x=3.985 //y=1.665
c78 ( 23 0 ) capacitor c=0.0371522f //x=3.985 //y=5.155
c79 ( 15 0 ) capacitor c=0.0266604f //x=3.205 //y=5.155
c80 ( 8 0 ) capacitor c=0.00549987f //x=1.615 //y=5.155
c81 ( 7 0 ) capacitor c=0.0226675f //x=2.325 //y=5.155
r82 (  31 32 ) resistor r=227.251 //w=0.187 //l=3.32 //layer=li \
 //thickness=0.1 //x=4.07 //y=1.75 //x2=4.07 //y2=5.07
r83 (  29 31 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=4.07 //y2=1.75
r84 (  29 30 ) resistor r=21.5615 //w=0.187 //l=0.315 //layer=li \
 //thickness=0.1 //x=3.985 //y=1.665 //x2=3.67 //y2=1.665
r85 (  25 30 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.585 //y=1.58 //x2=3.67 //y2=1.665
r86 (  25 35 ) resistor r=39.016 //w=0.187 //l=0.57 //layer=li //thickness=0.1 \
 //x=3.585 //y=1.58 //x2=3.585 //y2=1.01
r87 (  24 34 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.375 //y=5.155 //x2=3.29 //y2=5.155
r88 (  23 32 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=3.985 //y=5.155 //x2=4.07 //y2=5.07
r89 (  23 24 ) resistor r=41.754 //w=0.187 //l=0.61 //layer=li //thickness=0.1 \
 //x=3.985 //y=5.155 //x2=3.375 //y2=5.155
r90 (  17 34 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.155
r91 (  17 39 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=3.29 //y=5.24 //x2=3.29 //y2=5.725
r92 (  16 33 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.495 //y=5.155 //x2=2.41 //y2=5.155
r93 (  15 34 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.205 //y=5.155 //x2=3.29 //y2=5.155
r94 (  15 16 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li \
 //thickness=0.1 //x=3.205 //y=5.155 //x2=2.495 //y2=5.155
r95 (  9 33 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.41 //y=5.24 //x2=2.41 //y2=5.155
r96 (  9 38 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=2.41 //y=5.24 //x2=2.41 //y2=5.725
r97 (  7 33 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=2.325 //y=5.155 //x2=2.41 //y2=5.155
r98 (  7 8 ) resistor r=48.5989 //w=0.187 //l=0.71 //layer=li //thickness=0.1 \
 //x=2.325 //y=5.155 //x2=1.615 //y2=5.155
r99 (  1 8 ) resistor r=7.15173 //w=0.17 //l=0.120208 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.615 //y2=5.155
r100 (  1 37 ) resistor r=33.1979 //w=0.187 //l=0.485 //layer=li \
 //thickness=0.1 //x=1.53 //y=5.24 //x2=1.53 //y2=5.725
ends PM_NAND3X1_PCELL\%noxref_7

subckt PM_NAND3X1_PCELL\%noxref_8 ( 1 3 11 15 25 28 29 )
c41 ( 29 0 ) capacitor c=0.0457566f //x=2.965 //y=0.375
c42 ( 28 0 ) capacitor c=0.00467097f //x=1.86 //y=0.91
c43 ( 25 0 ) capacitor c=0.00156479f //x=3.1 //y=0.995
c44 ( 15 0 ) capacitor c=0.00737666f //x=4.07 //y=0.625
c45 ( 11 0 ) capacitor c=0.0152902f //x=3.985 //y=0.54
c46 ( 3 0 ) capacitor c=0.00718386f //x=3.1 //y=0.625
c47 ( 1 0 ) capacitor c=0.0279585f //x=3.015 //y=0.995
r48 (  15 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.5
r49 (  15 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li \
 //thickness=0.1 //x=4.07 //y=0.625 //x2=4.07 //y2=0.89
r50 (  12 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.185 //y=0.54 //x2=3.1 //y2=0.5
r51 (  12 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.185 //y=0.54 //x2=3.585 //y2=0.54
r52 (  11 29 ) resistor r=3.57586 //w=0.17 //l=0.103078 //layer=li \
 //thickness=0.1 //x=3.985 //y=0.54 //x2=4.07 //y2=0.5
r53 (  11 29 ) resistor r=27.3797 //w=0.187 //l=0.4 //layer=li //thickness=0.1 \
 //x=3.985 //y=0.54 //x2=3.585 //y2=0.54
r54 (  7 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=0.995
r55 (  7 29 ) resistor r=10.2674 //w=0.187 //l=0.15 //layer=li //thickness=0.1 \
 //x=3.1 //y=1.08 //x2=3.1 //y2=1.23
r56 (  4 25 ) resistor r=5.4201 //w=0.17 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.995
r57 (  4 29 ) resistor r=1.36898 //w=0.187 //l=0.02 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.91 //x2=3.1 //y2=0.89
r58 (  3 29 ) resistor r=3.57586 //w=0.17 //l=0.125 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.5
r59 (  3 29 ) resistor r=18.139 //w=0.187 //l=0.265 //layer=li //thickness=0.1 \
 //x=3.1 //y=0.625 //x2=3.1 //y2=0.89
r60 (  2 28 ) resistor r=0.751729 //w=0.17 //l=0.085 //layer=li \
 //thickness=0.1 //x=2.135 //y=0.995 //x2=2.05 //y2=0.995
r61 (  1 25 ) resistor r=1.40859 //w=0.34 //l=0.085 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=3.1 //y2=0.995
r62 (  1 2 ) resistor r=60.2353 //w=0.187 //l=0.88 //layer=li //thickness=0.1 \
 //x=3.015 //y=0.995 //x2=2.135 //y2=0.995
ends PM_NAND3X1_PCELL\%noxref_8

