magic
tech sky130A
magscale 1 2
timestamp 1669201029
<< nwell >>
rect -87 786 17181 1550
<< pwell >>
rect -34 -34 17128 544
<< nmos >>
rect 168 288 198 349
tri 198 288 214 304 sw
rect 362 296 392 349
tri 392 296 408 312 sw
rect 168 258 274 288
tri 274 258 304 288 sw
rect 362 266 468 296
tri 468 266 498 296 sw
rect 168 157 198 258
tri 198 242 214 258 nw
tri 258 242 274 258 ne
tri 198 157 214 173 sw
tri 258 157 274 173 se
rect 274 157 304 258
rect 362 165 392 266
tri 392 250 408 266 nw
tri 452 250 468 266 ne
tri 392 165 408 181 sw
tri 452 165 468 181 se
rect 468 165 498 266
tri 168 127 198 157 ne
rect 198 127 274 157
tri 274 127 304 157 nw
tri 362 135 392 165 ne
rect 392 135 468 165
tri 468 135 498 165 nw
rect 813 290 843 351
tri 843 290 859 306 sw
rect 1113 290 1143 351
rect 813 260 919 290
tri 919 260 949 290 sw
rect 813 159 843 260
tri 843 244 859 260 nw
tri 903 244 919 260 ne
tri 843 159 859 175 sw
tri 903 159 919 175 se
rect 919 159 949 260
tri 1008 260 1038 290 se
rect 1038 260 1143 290
rect 1008 166 1038 260
tri 1038 244 1054 260 nw
tri 1097 244 1113 260 ne
tri 1038 166 1054 182 sw
tri 1097 166 1113 182 se
rect 1113 166 1143 260
tri 813 129 843 159 ne
rect 843 129 919 159
tri 919 129 949 159 nw
tri 1008 136 1038 166 ne
rect 1038 136 1113 166
tri 1113 136 1143 166 nw
rect 1315 298 1345 351
tri 1345 298 1361 314 sw
rect 1315 268 1421 298
tri 1421 268 1451 298 sw
rect 1315 167 1345 268
tri 1345 252 1361 268 nw
tri 1405 252 1421 268 ne
tri 1345 167 1361 183 sw
tri 1405 167 1421 183 se
rect 1421 167 1451 268
tri 1315 137 1345 167 ne
rect 1345 137 1421 167
tri 1421 137 1451 167 nw
rect 1775 290 1805 351
tri 1805 290 1821 306 sw
rect 2075 290 2105 351
rect 1775 260 1881 290
tri 1881 260 1911 290 sw
rect 1775 159 1805 260
tri 1805 244 1821 260 nw
tri 1865 244 1881 260 ne
tri 1805 159 1821 175 sw
tri 1865 159 1881 175 se
rect 1881 159 1911 260
tri 1970 260 2000 290 se
rect 2000 260 2105 290
rect 1970 166 2000 260
tri 2000 244 2016 260 nw
tri 2059 244 2075 260 ne
tri 2000 166 2016 182 sw
tri 2059 166 2075 182 se
rect 2075 166 2105 260
tri 1775 129 1805 159 ne
rect 1805 129 1881 159
tri 1881 129 1911 159 nw
tri 1970 136 2000 166 ne
rect 2000 136 2075 166
tri 2075 136 2105 166 nw
rect 2277 298 2307 351
tri 2307 298 2323 314 sw
rect 2277 268 2383 298
tri 2383 268 2413 298 sw
rect 2277 167 2307 268
tri 2307 252 2323 268 nw
tri 2367 252 2383 268 ne
tri 2307 167 2323 183 sw
tri 2367 167 2383 183 se
rect 2383 167 2413 268
tri 2277 137 2307 167 ne
rect 2307 137 2383 167
tri 2383 137 2413 167 nw
rect 2758 288 2788 349
tri 2788 288 2804 304 sw
rect 2952 296 2982 349
tri 2982 296 2998 312 sw
rect 2758 258 2864 288
tri 2864 258 2894 288 sw
rect 2952 266 3058 296
tri 3058 266 3088 296 sw
rect 2758 157 2788 258
tri 2788 242 2804 258 nw
tri 2848 242 2864 258 ne
tri 2788 157 2804 173 sw
tri 2848 157 2864 173 se
rect 2864 157 2894 258
rect 2952 165 2982 266
tri 2982 250 2998 266 nw
tri 3042 250 3058 266 ne
tri 2982 165 2998 181 sw
tri 3042 165 3058 181 se
rect 3058 165 3088 266
tri 2758 127 2788 157 ne
rect 2788 127 2864 157
tri 2864 127 2894 157 nw
tri 2952 135 2982 165 ne
rect 2982 135 3058 165
tri 3058 135 3088 165 nw
rect 3424 288 3454 349
tri 3454 288 3470 304 sw
rect 3618 296 3648 349
tri 3648 296 3664 312 sw
rect 3424 258 3530 288
tri 3530 258 3560 288 sw
rect 3618 266 3724 296
tri 3724 266 3754 296 sw
rect 3424 157 3454 258
tri 3454 242 3470 258 nw
tri 3514 242 3530 258 ne
tri 3454 157 3470 173 sw
tri 3514 157 3530 173 se
rect 3530 157 3560 258
rect 3618 165 3648 266
tri 3648 250 3664 266 nw
tri 3708 250 3724 266 ne
tri 3648 165 3664 181 sw
tri 3708 165 3724 181 se
rect 3724 165 3754 266
tri 3424 127 3454 157 ne
rect 3454 127 3530 157
tri 3530 127 3560 157 nw
tri 3618 135 3648 165 ne
rect 3648 135 3724 165
tri 3724 135 3754 165 nw
rect 4069 290 4099 351
tri 4099 290 4115 306 sw
rect 4369 290 4399 351
rect 4069 260 4175 290
tri 4175 260 4205 290 sw
rect 4069 159 4099 260
tri 4099 244 4115 260 nw
tri 4159 244 4175 260 ne
tri 4099 159 4115 175 sw
tri 4159 159 4175 175 se
rect 4175 159 4205 260
tri 4264 260 4294 290 se
rect 4294 260 4399 290
rect 4264 166 4294 260
tri 4294 244 4310 260 nw
tri 4353 244 4369 260 ne
tri 4294 166 4310 182 sw
tri 4353 166 4369 182 se
rect 4369 166 4399 260
tri 4069 129 4099 159 ne
rect 4099 129 4175 159
tri 4175 129 4205 159 nw
tri 4264 136 4294 166 ne
rect 4294 136 4369 166
tri 4369 136 4399 166 nw
rect 4571 298 4601 351
tri 4601 298 4617 314 sw
rect 4571 268 4677 298
tri 4677 268 4707 298 sw
rect 4571 167 4601 268
tri 4601 252 4617 268 nw
tri 4661 252 4677 268 ne
tri 4601 167 4617 183 sw
tri 4661 167 4677 183 se
rect 4677 167 4707 268
tri 4571 137 4601 167 ne
rect 4601 137 4677 167
tri 4677 137 4707 167 nw
rect 5052 288 5082 349
tri 5082 288 5098 304 sw
rect 5246 296 5276 349
tri 5276 296 5292 312 sw
rect 5052 258 5158 288
tri 5158 258 5188 288 sw
rect 5246 266 5352 296
tri 5352 266 5382 296 sw
rect 5052 157 5082 258
tri 5082 242 5098 258 nw
tri 5142 242 5158 258 ne
tri 5082 157 5098 173 sw
tri 5142 157 5158 173 se
rect 5158 157 5188 258
rect 5246 165 5276 266
tri 5276 250 5292 266 nw
tri 5336 250 5352 266 ne
tri 5276 165 5292 181 sw
tri 5336 165 5352 181 se
rect 5352 165 5382 266
tri 5052 127 5082 157 ne
rect 5082 127 5158 157
tri 5158 127 5188 157 nw
tri 5246 135 5276 165 ne
rect 5276 135 5352 165
tri 5352 135 5382 165 nw
rect 5697 290 5727 351
tri 5727 290 5743 306 sw
rect 5997 290 6027 351
rect 5697 260 5803 290
tri 5803 260 5833 290 sw
rect 5697 159 5727 260
tri 5727 244 5743 260 nw
tri 5787 244 5803 260 ne
tri 5727 159 5743 175 sw
tri 5787 159 5803 175 se
rect 5803 159 5833 260
tri 5892 260 5922 290 se
rect 5922 260 6027 290
rect 5892 166 5922 260
tri 5922 244 5938 260 nw
tri 5981 244 5997 260 ne
tri 5922 166 5938 182 sw
tri 5981 166 5997 182 se
rect 5997 166 6027 260
tri 5697 129 5727 159 ne
rect 5727 129 5803 159
tri 5803 129 5833 159 nw
tri 5892 136 5922 166 ne
rect 5922 136 5997 166
tri 5997 136 6027 166 nw
rect 6199 298 6229 351
tri 6229 298 6245 314 sw
rect 6199 268 6305 298
tri 6305 268 6335 298 sw
rect 6199 167 6229 268
tri 6229 252 6245 268 nw
tri 6289 252 6305 268 ne
tri 6229 167 6245 183 sw
tri 6289 167 6305 183 se
rect 6305 167 6335 268
tri 6199 137 6229 167 ne
rect 6229 137 6305 167
tri 6305 137 6335 167 nw
rect 6659 290 6689 351
tri 6689 290 6705 306 sw
rect 6959 290 6989 351
rect 6659 260 6765 290
tri 6765 260 6795 290 sw
rect 6659 159 6689 260
tri 6689 244 6705 260 nw
tri 6749 244 6765 260 ne
tri 6689 159 6705 175 sw
tri 6749 159 6765 175 se
rect 6765 159 6795 260
tri 6854 260 6884 290 se
rect 6884 260 6989 290
rect 6854 166 6884 260
tri 6884 244 6900 260 nw
tri 6943 244 6959 260 ne
tri 6884 166 6900 182 sw
tri 6943 166 6959 182 se
rect 6959 166 6989 260
tri 6659 129 6689 159 ne
rect 6689 129 6765 159
tri 6765 129 6795 159 nw
tri 6854 136 6884 166 ne
rect 6884 136 6959 166
tri 6959 136 6989 166 nw
rect 7161 298 7191 351
tri 7191 298 7207 314 sw
rect 7161 268 7267 298
tri 7267 268 7297 298 sw
rect 7161 167 7191 268
tri 7191 252 7207 268 nw
tri 7251 252 7267 268 ne
tri 7191 167 7207 183 sw
tri 7251 167 7267 183 se
rect 7267 167 7297 268
tri 7161 137 7191 167 ne
rect 7191 137 7267 167
tri 7267 137 7297 167 nw
rect 7642 288 7672 349
tri 7672 288 7688 304 sw
rect 7836 296 7866 349
tri 7866 296 7882 312 sw
rect 7642 258 7748 288
tri 7748 258 7778 288 sw
rect 7836 266 7942 296
tri 7942 266 7972 296 sw
rect 7642 157 7672 258
tri 7672 242 7688 258 nw
tri 7732 242 7748 258 ne
tri 7672 157 7688 173 sw
tri 7732 157 7748 173 se
rect 7748 157 7778 258
rect 7836 165 7866 266
tri 7866 250 7882 266 nw
tri 7926 250 7942 266 ne
tri 7866 165 7882 181 sw
tri 7926 165 7942 181 se
rect 7942 165 7972 266
tri 7642 127 7672 157 ne
rect 7672 127 7748 157
tri 7748 127 7778 157 nw
tri 7836 135 7866 165 ne
rect 7866 135 7942 165
tri 7942 135 7972 165 nw
rect 8308 288 8338 349
tri 8338 288 8354 304 sw
rect 8502 296 8532 349
tri 8532 296 8548 312 sw
rect 8308 258 8414 288
tri 8414 258 8444 288 sw
rect 8502 266 8608 296
tri 8608 266 8638 296 sw
rect 8308 157 8338 258
tri 8338 242 8354 258 nw
tri 8398 242 8414 258 ne
tri 8338 157 8354 173 sw
tri 8398 157 8414 173 se
rect 8414 157 8444 258
rect 8502 165 8532 266
tri 8532 250 8548 266 nw
tri 8592 250 8608 266 ne
tri 8532 165 8548 181 sw
tri 8592 165 8608 181 se
rect 8608 165 8638 266
tri 8308 127 8338 157 ne
rect 8338 127 8414 157
tri 8414 127 8444 157 nw
tri 8502 135 8532 165 ne
rect 8532 135 8608 165
tri 8608 135 8638 165 nw
rect 8953 290 8983 351
tri 8983 290 8999 306 sw
rect 9253 290 9283 351
rect 8953 260 9059 290
tri 9059 260 9089 290 sw
rect 8953 159 8983 260
tri 8983 244 8999 260 nw
tri 9043 244 9059 260 ne
tri 8983 159 8999 175 sw
tri 9043 159 9059 175 se
rect 9059 159 9089 260
tri 9148 260 9178 290 se
rect 9178 260 9283 290
rect 9148 166 9178 260
tri 9178 244 9194 260 nw
tri 9237 244 9253 260 ne
tri 9178 166 9194 182 sw
tri 9237 166 9253 182 se
rect 9253 166 9283 260
tri 8953 129 8983 159 ne
rect 8983 129 9059 159
tri 9059 129 9089 159 nw
tri 9148 136 9178 166 ne
rect 9178 136 9253 166
tri 9253 136 9283 166 nw
rect 9455 298 9485 351
tri 9485 298 9501 314 sw
rect 9455 268 9561 298
tri 9561 268 9591 298 sw
rect 9455 167 9485 268
tri 9485 252 9501 268 nw
tri 9545 252 9561 268 ne
tri 9485 167 9501 183 sw
tri 9545 167 9561 183 se
rect 9561 167 9591 268
tri 9455 137 9485 167 ne
rect 9485 137 9561 167
tri 9561 137 9591 167 nw
rect 9936 288 9966 349
tri 9966 288 9982 304 sw
rect 10130 296 10160 349
tri 10160 296 10176 312 sw
rect 9936 258 10042 288
tri 10042 258 10072 288 sw
rect 10130 266 10236 296
tri 10236 266 10266 296 sw
rect 9936 157 9966 258
tri 9966 242 9982 258 nw
tri 10026 242 10042 258 ne
tri 9966 157 9982 173 sw
tri 10026 157 10042 173 se
rect 10042 157 10072 258
rect 10130 165 10160 266
tri 10160 250 10176 266 nw
tri 10220 250 10236 266 ne
tri 10160 165 10176 181 sw
tri 10220 165 10236 181 se
rect 10236 165 10266 266
tri 9936 127 9966 157 ne
rect 9966 127 10042 157
tri 10042 127 10072 157 nw
tri 10130 135 10160 165 ne
rect 10160 135 10236 165
tri 10236 135 10266 165 nw
rect 10581 290 10611 351
tri 10611 290 10627 306 sw
rect 10881 290 10911 351
rect 10581 260 10687 290
tri 10687 260 10717 290 sw
rect 10581 159 10611 260
tri 10611 244 10627 260 nw
tri 10671 244 10687 260 ne
tri 10611 159 10627 175 sw
tri 10671 159 10687 175 se
rect 10687 159 10717 260
tri 10776 260 10806 290 se
rect 10806 260 10911 290
rect 10776 166 10806 260
tri 10806 244 10822 260 nw
tri 10865 244 10881 260 ne
tri 10806 166 10822 182 sw
tri 10865 166 10881 182 se
rect 10881 166 10911 260
tri 10581 129 10611 159 ne
rect 10611 129 10687 159
tri 10687 129 10717 159 nw
tri 10776 136 10806 166 ne
rect 10806 136 10881 166
tri 10881 136 10911 166 nw
rect 11083 298 11113 351
tri 11113 298 11129 314 sw
rect 11083 268 11189 298
tri 11189 268 11219 298 sw
rect 11083 167 11113 268
tri 11113 252 11129 268 nw
tri 11173 252 11189 268 ne
tri 11113 167 11129 183 sw
tri 11173 167 11189 183 se
rect 11189 167 11219 268
tri 11083 137 11113 167 ne
rect 11113 137 11189 167
tri 11189 137 11219 167 nw
rect 11543 290 11573 351
tri 11573 290 11589 306 sw
rect 11843 290 11873 351
rect 11543 260 11649 290
tri 11649 260 11679 290 sw
rect 11543 159 11573 260
tri 11573 244 11589 260 nw
tri 11633 244 11649 260 ne
tri 11573 159 11589 175 sw
tri 11633 159 11649 175 se
rect 11649 159 11679 260
tri 11738 260 11768 290 se
rect 11768 260 11873 290
rect 11738 166 11768 260
tri 11768 244 11784 260 nw
tri 11827 244 11843 260 ne
tri 11768 166 11784 182 sw
tri 11827 166 11843 182 se
rect 11843 166 11873 260
tri 11543 129 11573 159 ne
rect 11573 129 11649 159
tri 11649 129 11679 159 nw
tri 11738 136 11768 166 ne
rect 11768 136 11843 166
tri 11843 136 11873 166 nw
rect 12045 298 12075 351
tri 12075 298 12091 314 sw
rect 12045 268 12151 298
tri 12151 268 12181 298 sw
rect 12045 167 12075 268
tri 12075 252 12091 268 nw
tri 12135 252 12151 268 ne
tri 12075 167 12091 183 sw
tri 12135 167 12151 183 se
rect 12151 167 12181 268
tri 12045 137 12075 167 ne
rect 12075 137 12151 167
tri 12151 137 12181 167 nw
rect 12526 288 12556 349
tri 12556 288 12572 304 sw
rect 12720 296 12750 349
tri 12750 296 12766 312 sw
rect 12526 258 12632 288
tri 12632 258 12662 288 sw
rect 12720 266 12826 296
tri 12826 266 12856 296 sw
rect 12526 157 12556 258
tri 12556 242 12572 258 nw
tri 12616 242 12632 258 ne
tri 12556 157 12572 173 sw
tri 12616 157 12632 173 se
rect 12632 157 12662 258
rect 12720 165 12750 266
tri 12750 250 12766 266 nw
tri 12810 250 12826 266 ne
tri 12750 165 12766 181 sw
tri 12810 165 12826 181 se
rect 12826 165 12856 266
tri 12526 127 12556 157 ne
rect 12556 127 12632 157
tri 12632 127 12662 157 nw
tri 12720 135 12750 165 ne
rect 12750 135 12826 165
tri 12826 135 12856 165 nw
rect 13192 288 13222 349
tri 13222 288 13238 304 sw
rect 13386 296 13416 349
tri 13416 296 13432 312 sw
rect 13192 258 13298 288
tri 13298 258 13328 288 sw
rect 13386 266 13492 296
tri 13492 266 13522 296 sw
rect 13192 157 13222 258
tri 13222 242 13238 258 nw
tri 13282 242 13298 258 ne
tri 13222 157 13238 173 sw
tri 13282 157 13298 173 se
rect 13298 157 13328 258
rect 13386 165 13416 266
tri 13416 250 13432 266 nw
tri 13476 250 13492 266 ne
tri 13416 165 13432 181 sw
tri 13476 165 13492 181 se
rect 13492 165 13522 266
tri 13192 127 13222 157 ne
rect 13222 127 13298 157
tri 13298 127 13328 157 nw
tri 13386 135 13416 165 ne
rect 13416 135 13492 165
tri 13492 135 13522 165 nw
rect 13837 290 13867 351
tri 13867 290 13883 306 sw
rect 14137 290 14167 351
rect 13837 260 13943 290
tri 13943 260 13973 290 sw
rect 13837 159 13867 260
tri 13867 244 13883 260 nw
tri 13927 244 13943 260 ne
tri 13867 159 13883 175 sw
tri 13927 159 13943 175 se
rect 13943 159 13973 260
tri 14032 260 14062 290 se
rect 14062 260 14167 290
rect 14032 166 14062 260
tri 14062 244 14078 260 nw
tri 14121 244 14137 260 ne
tri 14062 166 14078 182 sw
tri 14121 166 14137 182 se
rect 14137 166 14167 260
tri 13837 129 13867 159 ne
rect 13867 129 13943 159
tri 13943 129 13973 159 nw
tri 14032 136 14062 166 ne
rect 14062 136 14137 166
tri 14137 136 14167 166 nw
rect 14339 298 14369 351
tri 14369 298 14385 314 sw
rect 14339 268 14445 298
tri 14445 268 14475 298 sw
rect 14339 167 14369 268
tri 14369 252 14385 268 nw
tri 14429 252 14445 268 ne
tri 14369 167 14385 183 sw
tri 14429 167 14445 183 se
rect 14445 167 14475 268
tri 14339 137 14369 167 ne
rect 14369 137 14445 167
tri 14445 137 14475 167 nw
rect 14820 288 14850 349
tri 14850 288 14866 304 sw
rect 15014 296 15044 349
tri 15044 296 15060 312 sw
rect 14820 258 14926 288
tri 14926 258 14956 288 sw
rect 15014 266 15120 296
tri 15120 266 15150 296 sw
rect 14820 157 14850 258
tri 14850 242 14866 258 nw
tri 14910 242 14926 258 ne
tri 14850 157 14866 173 sw
tri 14910 157 14926 173 se
rect 14926 157 14956 258
rect 15014 165 15044 266
tri 15044 250 15060 266 nw
tri 15104 250 15120 266 ne
tri 15044 165 15060 181 sw
tri 15104 165 15120 181 se
rect 15120 165 15150 266
tri 14820 127 14850 157 ne
rect 14850 127 14926 157
tri 14926 127 14956 157 nw
tri 15014 135 15044 165 ne
rect 15044 135 15120 165
tri 15120 135 15150 165 nw
rect 15486 288 15516 349
tri 15516 288 15532 304 sw
tri 15770 296 15786 312 se
rect 15786 296 15816 349
rect 15486 258 15592 288
tri 15592 258 15622 288 sw
tri 15680 266 15710 296 se
rect 15710 266 15816 296
rect 15486 157 15516 258
tri 15516 242 15532 258 nw
tri 15576 242 15592 258 ne
tri 15516 157 15532 173 sw
tri 15576 157 15592 173 se
rect 15592 157 15622 258
rect 15680 165 15710 266
tri 15710 250 15726 266 nw
tri 15770 250 15786 266 ne
tri 15710 165 15726 181 sw
tri 15770 165 15786 181 se
rect 15786 165 15816 266
tri 15486 127 15516 157 ne
rect 15516 127 15592 157
tri 15592 127 15622 157 nw
tri 15680 135 15710 165 ne
rect 15710 135 15786 165
tri 15786 135 15816 165 nw
rect 16152 288 16182 349
tri 16182 288 16198 304 sw
rect 16346 296 16376 349
tri 16376 296 16392 312 sw
rect 16152 258 16258 288
tri 16258 258 16288 288 sw
rect 16346 266 16452 296
tri 16452 266 16482 296 sw
rect 16152 157 16182 258
tri 16182 242 16198 258 nw
tri 16242 242 16258 258 ne
tri 16182 157 16198 173 sw
tri 16242 157 16258 173 se
rect 16258 157 16288 258
rect 16346 251 16377 266
tri 16377 251 16392 266 nw
tri 16436 251 16451 266 ne
rect 16451 251 16482 266
rect 16346 165 16376 251
tri 16376 165 16392 181 sw
tri 16436 165 16452 181 se
rect 16452 165 16482 251
tri 16152 127 16182 157 ne
rect 16182 127 16258 157
tri 16258 127 16288 157 nw
tri 16346 135 16376 165 ne
rect 16376 135 16452 165
tri 16452 135 16482 165 nw
rect 16805 297 16835 350
tri 16835 297 16851 313 sw
rect 16805 267 16911 297
tri 16911 267 16941 297 sw
rect 16805 166 16835 267
tri 16835 251 16851 267 nw
tri 16895 251 16911 267 ne
tri 16835 166 16851 182 sw
tri 16895 166 16911 182 se
rect 16911 166 16941 267
tri 16805 136 16835 166 ne
rect 16835 136 16911 166
tri 16911 136 16941 166 nw
<< pmos >>
rect 187 1004 217 1404
rect 275 1004 305 1404
rect 363 1004 393 1404
rect 451 1004 481 1404
rect 913 1004 943 1404
rect 1001 1004 1031 1404
rect 1089 1004 1119 1404
rect 1177 1004 1207 1404
rect 1265 1004 1295 1404
rect 1353 1004 1383 1404
rect 1875 1004 1905 1404
rect 1963 1004 1993 1404
rect 2051 1004 2081 1404
rect 2139 1004 2169 1404
rect 2227 1004 2257 1404
rect 2315 1004 2345 1404
rect 2777 1004 2807 1404
rect 2865 1004 2895 1404
rect 2953 1004 2983 1404
rect 3041 1004 3071 1404
rect 3443 1004 3473 1404
rect 3531 1004 3561 1404
rect 3619 1004 3649 1404
rect 3707 1004 3737 1404
rect 4169 1004 4199 1404
rect 4257 1004 4287 1404
rect 4345 1004 4375 1404
rect 4433 1004 4463 1404
rect 4521 1004 4551 1404
rect 4609 1004 4639 1404
rect 5071 1004 5101 1404
rect 5159 1004 5189 1404
rect 5247 1004 5277 1404
rect 5335 1004 5365 1404
rect 5797 1004 5827 1404
rect 5885 1004 5915 1404
rect 5973 1004 6003 1404
rect 6061 1004 6091 1404
rect 6149 1004 6179 1404
rect 6237 1004 6267 1404
rect 6759 1004 6789 1404
rect 6847 1004 6877 1404
rect 6935 1004 6965 1404
rect 7023 1004 7053 1404
rect 7111 1004 7141 1404
rect 7199 1004 7229 1404
rect 7661 1004 7691 1404
rect 7749 1004 7779 1404
rect 7837 1004 7867 1404
rect 7925 1004 7955 1404
rect 8327 1004 8357 1404
rect 8415 1004 8445 1404
rect 8503 1004 8533 1404
rect 8591 1004 8621 1404
rect 9053 1004 9083 1404
rect 9141 1004 9171 1404
rect 9229 1004 9259 1404
rect 9317 1004 9347 1404
rect 9405 1004 9435 1404
rect 9493 1004 9523 1404
rect 9955 1004 9985 1404
rect 10043 1004 10073 1404
rect 10131 1004 10161 1404
rect 10219 1004 10249 1404
rect 10681 1004 10711 1404
rect 10769 1004 10799 1404
rect 10857 1004 10887 1404
rect 10945 1004 10975 1404
rect 11033 1004 11063 1404
rect 11121 1004 11151 1404
rect 11643 1004 11673 1404
rect 11731 1004 11761 1404
rect 11819 1004 11849 1404
rect 11907 1004 11937 1404
rect 11995 1004 12025 1404
rect 12083 1004 12113 1404
rect 12545 1004 12575 1404
rect 12633 1004 12663 1404
rect 12721 1004 12751 1404
rect 12809 1004 12839 1404
rect 13211 1004 13241 1404
rect 13299 1004 13329 1404
rect 13387 1004 13417 1404
rect 13475 1004 13505 1404
rect 13937 1004 13967 1404
rect 14025 1004 14055 1404
rect 14113 1004 14143 1404
rect 14201 1004 14231 1404
rect 14289 1004 14319 1404
rect 14377 1004 14407 1404
rect 14839 1005 14869 1405
rect 14927 1005 14957 1405
rect 15015 1005 15045 1405
rect 15103 1005 15133 1405
rect 15503 1005 15533 1405
rect 15591 1005 15621 1405
rect 15679 1005 15709 1405
rect 15767 1005 15797 1405
rect 16171 1005 16201 1405
rect 16259 1005 16289 1405
rect 16347 1005 16377 1405
rect 16435 1005 16465 1405
rect 16814 1004 16844 1404
rect 16902 1004 16932 1404
<< ndiff >>
rect 112 333 168 349
rect 112 299 122 333
rect 156 299 168 333
rect 112 261 168 299
rect 198 333 362 349
rect 198 304 219 333
tri 198 288 214 304 ne
rect 214 299 219 304
rect 253 299 316 333
rect 350 299 362 333
rect 214 288 362 299
rect 392 312 554 349
tri 392 296 408 312 ne
rect 408 296 554 312
rect 112 227 122 261
rect 156 227 168 261
tri 274 258 304 288 ne
rect 304 261 362 288
tri 468 266 498 296 ne
rect 112 193 168 227
rect 112 159 122 193
rect 156 159 168 193
rect 112 127 168 159
tri 198 242 214 258 se
rect 214 242 258 258
tri 258 242 274 258 sw
rect 198 208 274 242
rect 198 174 219 208
rect 253 174 274 208
rect 198 173 274 174
tri 198 157 214 173 ne
rect 214 157 258 173
tri 258 157 274 173 nw
rect 304 227 316 261
rect 350 227 362 261
rect 304 193 362 227
rect 304 159 316 193
rect 350 159 362 193
tri 392 250 408 266 se
rect 408 250 452 266
tri 452 250 468 266 sw
rect 392 217 468 250
rect 392 183 413 217
rect 447 183 468 217
rect 392 181 468 183
tri 392 165 408 181 ne
rect 408 165 452 181
tri 452 165 468 181 nw
rect 498 261 554 296
rect 498 227 510 261
rect 544 227 554 261
rect 498 193 554 227
tri 168 127 198 157 sw
tri 274 127 304 157 se
rect 304 135 362 159
tri 362 135 392 165 sw
tri 468 135 498 165 se
rect 498 159 510 193
rect 544 159 554 193
rect 498 135 554 159
rect 304 127 554 135
rect 112 123 554 127
rect 112 89 122 123
rect 156 89 316 123
rect 350 89 413 123
rect 447 89 510 123
rect 544 89 554 123
rect 112 73 554 89
rect 757 335 813 351
rect 757 301 767 335
rect 801 301 813 335
rect 757 263 813 301
rect 843 335 1113 351
rect 843 306 864 335
tri 843 290 859 306 ne
rect 859 301 864 306
rect 898 301 961 335
rect 995 301 1058 335
rect 1092 301 1113 335
rect 859 290 1113 301
rect 1143 335 1199 351
rect 1143 301 1155 335
rect 1189 301 1199 335
rect 757 229 767 263
rect 801 229 813 263
tri 919 260 949 290 ne
rect 949 263 1008 290
rect 757 195 813 229
rect 757 161 767 195
rect 801 161 813 195
rect 757 129 813 161
tri 843 244 859 260 se
rect 859 244 903 260
tri 903 244 919 260 sw
rect 843 210 919 244
rect 843 176 864 210
rect 898 176 919 210
rect 843 175 919 176
tri 843 159 859 175 ne
rect 859 159 903 175
tri 903 159 919 175 nw
rect 949 229 961 263
rect 995 229 1008 263
tri 1008 260 1038 290 nw
rect 949 195 1008 229
rect 949 161 961 195
rect 995 161 1008 195
tri 1038 244 1054 260 se
rect 1054 244 1097 260
tri 1097 244 1113 260 sw
rect 1038 216 1113 244
rect 1038 182 1059 216
rect 1093 182 1113 216
tri 1038 166 1054 182 ne
rect 1054 166 1097 182
tri 1097 166 1113 182 nw
tri 813 129 843 159 sw
tri 919 129 949 159 se
rect 949 136 1008 161
tri 1008 136 1038 166 sw
tri 1113 136 1143 166 se
rect 1143 136 1199 301
rect 949 129 1199 136
rect 757 125 1199 129
rect 757 91 767 125
rect 801 91 961 125
rect 995 91 1058 125
rect 1092 91 1155 125
rect 1189 91 1199 125
rect 757 75 1199 91
rect 1259 335 1315 351
rect 1259 301 1269 335
rect 1303 301 1315 335
rect 1259 263 1315 301
rect 1345 314 1507 351
tri 1345 298 1361 314 ne
rect 1361 298 1507 314
tri 1421 268 1451 298 ne
rect 1259 229 1269 263
rect 1303 229 1315 263
rect 1259 195 1315 229
rect 1259 161 1269 195
rect 1303 161 1315 195
tri 1345 252 1361 268 se
rect 1361 252 1405 268
tri 1405 252 1421 268 sw
rect 1345 219 1421 252
rect 1345 185 1366 219
rect 1400 185 1421 219
rect 1345 183 1421 185
tri 1345 167 1361 183 ne
rect 1361 167 1405 183
tri 1405 167 1421 183 nw
rect 1451 263 1507 298
rect 1451 229 1463 263
rect 1497 229 1507 263
rect 1451 195 1507 229
rect 1259 137 1315 161
tri 1315 137 1345 167 sw
tri 1421 137 1451 167 se
rect 1451 161 1463 195
rect 1497 161 1507 195
rect 1451 137 1507 161
rect 1259 125 1507 137
rect 1259 91 1269 125
rect 1303 91 1366 125
rect 1400 91 1463 125
rect 1497 91 1507 125
rect 1259 75 1507 91
rect 1719 335 1775 351
rect 1719 301 1729 335
rect 1763 301 1775 335
rect 1719 263 1775 301
rect 1805 335 2075 351
rect 1805 306 1826 335
tri 1805 290 1821 306 ne
rect 1821 301 1826 306
rect 1860 301 1923 335
rect 1957 301 2020 335
rect 2054 301 2075 335
rect 1821 290 2075 301
rect 2105 335 2161 351
rect 2105 301 2117 335
rect 2151 301 2161 335
rect 1719 229 1729 263
rect 1763 229 1775 263
tri 1881 260 1911 290 ne
rect 1911 263 1970 290
rect 1719 195 1775 229
rect 1719 161 1729 195
rect 1763 161 1775 195
rect 1719 129 1775 161
tri 1805 244 1821 260 se
rect 1821 244 1865 260
tri 1865 244 1881 260 sw
rect 1805 210 1881 244
rect 1805 176 1826 210
rect 1860 176 1881 210
rect 1805 175 1881 176
tri 1805 159 1821 175 ne
rect 1821 159 1865 175
tri 1865 159 1881 175 nw
rect 1911 229 1923 263
rect 1957 229 1970 263
tri 1970 260 2000 290 nw
rect 1911 195 1970 229
rect 1911 161 1923 195
rect 1957 161 1970 195
tri 2000 244 2016 260 se
rect 2016 244 2059 260
tri 2059 244 2075 260 sw
rect 2000 216 2075 244
rect 2000 182 2021 216
rect 2055 182 2075 216
tri 2000 166 2016 182 ne
rect 2016 166 2059 182
tri 2059 166 2075 182 nw
tri 1775 129 1805 159 sw
tri 1881 129 1911 159 se
rect 1911 136 1970 161
tri 1970 136 2000 166 sw
tri 2075 136 2105 166 se
rect 2105 136 2161 301
rect 1911 129 2161 136
rect 1719 125 2161 129
rect 1719 91 1729 125
rect 1763 91 1923 125
rect 1957 91 2020 125
rect 2054 91 2117 125
rect 2151 91 2161 125
rect 1719 75 2161 91
rect 2221 335 2277 351
rect 2221 301 2231 335
rect 2265 301 2277 335
rect 2221 263 2277 301
rect 2307 314 2469 351
tri 2307 298 2323 314 ne
rect 2323 298 2469 314
tri 2383 268 2413 298 ne
rect 2221 229 2231 263
rect 2265 229 2277 263
rect 2221 195 2277 229
rect 2221 161 2231 195
rect 2265 161 2277 195
tri 2307 252 2323 268 se
rect 2323 252 2367 268
tri 2367 252 2383 268 sw
rect 2307 219 2383 252
rect 2307 185 2328 219
rect 2362 185 2383 219
rect 2307 183 2383 185
tri 2307 167 2323 183 ne
rect 2323 167 2367 183
tri 2367 167 2383 183 nw
rect 2413 263 2469 298
rect 2413 229 2425 263
rect 2459 229 2469 263
rect 2413 195 2469 229
rect 2221 137 2277 161
tri 2277 137 2307 167 sw
tri 2383 137 2413 167 se
rect 2413 161 2425 195
rect 2459 161 2469 195
rect 2413 137 2469 161
rect 2221 125 2469 137
rect 2221 91 2231 125
rect 2265 91 2328 125
rect 2362 91 2425 125
rect 2459 91 2469 125
rect 2221 75 2469 91
rect 2702 333 2758 349
rect 2702 299 2712 333
rect 2746 299 2758 333
rect 2702 261 2758 299
rect 2788 333 2952 349
rect 2788 304 2809 333
tri 2788 288 2804 304 ne
rect 2804 299 2809 304
rect 2843 299 2906 333
rect 2940 299 2952 333
rect 2804 288 2952 299
rect 2982 312 3144 349
tri 2982 296 2998 312 ne
rect 2998 296 3144 312
rect 2702 227 2712 261
rect 2746 227 2758 261
tri 2864 258 2894 288 ne
rect 2894 261 2952 288
tri 3058 266 3088 296 ne
rect 2702 193 2758 227
rect 2702 159 2712 193
rect 2746 159 2758 193
rect 2702 127 2758 159
tri 2788 242 2804 258 se
rect 2804 242 2848 258
tri 2848 242 2864 258 sw
rect 2788 208 2864 242
rect 2788 174 2809 208
rect 2843 174 2864 208
rect 2788 173 2864 174
tri 2788 157 2804 173 ne
rect 2804 157 2848 173
tri 2848 157 2864 173 nw
rect 2894 227 2906 261
rect 2940 227 2952 261
rect 2894 193 2952 227
rect 2894 159 2906 193
rect 2940 159 2952 193
tri 2982 250 2998 266 se
rect 2998 250 3042 266
tri 3042 250 3058 266 sw
rect 2982 217 3058 250
rect 2982 183 3003 217
rect 3037 183 3058 217
rect 2982 181 3058 183
tri 2982 165 2998 181 ne
rect 2998 165 3042 181
tri 3042 165 3058 181 nw
rect 3088 261 3144 296
rect 3088 227 3100 261
rect 3134 227 3144 261
rect 3088 193 3144 227
tri 2758 127 2788 157 sw
tri 2864 127 2894 157 se
rect 2894 135 2952 159
tri 2952 135 2982 165 sw
tri 3058 135 3088 165 se
rect 3088 159 3100 193
rect 3134 159 3144 193
rect 3088 135 3144 159
rect 2894 127 3144 135
rect 2702 123 3144 127
rect 2702 89 2712 123
rect 2746 89 2906 123
rect 2940 89 3003 123
rect 3037 89 3100 123
rect 3134 89 3144 123
rect 2702 73 3144 89
rect 3368 333 3424 349
rect 3368 299 3378 333
rect 3412 299 3424 333
rect 3368 261 3424 299
rect 3454 333 3618 349
rect 3454 304 3475 333
tri 3454 288 3470 304 ne
rect 3470 299 3475 304
rect 3509 299 3572 333
rect 3606 299 3618 333
rect 3470 288 3618 299
rect 3648 312 3810 349
tri 3648 296 3664 312 ne
rect 3664 296 3810 312
rect 3368 227 3378 261
rect 3412 227 3424 261
tri 3530 258 3560 288 ne
rect 3560 261 3618 288
tri 3724 266 3754 296 ne
rect 3368 193 3424 227
rect 3368 159 3378 193
rect 3412 159 3424 193
rect 3368 127 3424 159
tri 3454 242 3470 258 se
rect 3470 242 3514 258
tri 3514 242 3530 258 sw
rect 3454 208 3530 242
rect 3454 174 3475 208
rect 3509 174 3530 208
rect 3454 173 3530 174
tri 3454 157 3470 173 ne
rect 3470 157 3514 173
tri 3514 157 3530 173 nw
rect 3560 227 3572 261
rect 3606 227 3618 261
rect 3560 193 3618 227
rect 3560 159 3572 193
rect 3606 159 3618 193
tri 3648 250 3664 266 se
rect 3664 250 3708 266
tri 3708 250 3724 266 sw
rect 3648 217 3724 250
rect 3648 183 3669 217
rect 3703 183 3724 217
rect 3648 181 3724 183
tri 3648 165 3664 181 ne
rect 3664 165 3708 181
tri 3708 165 3724 181 nw
rect 3754 261 3810 296
rect 3754 227 3766 261
rect 3800 227 3810 261
rect 3754 193 3810 227
tri 3424 127 3454 157 sw
tri 3530 127 3560 157 se
rect 3560 135 3618 159
tri 3618 135 3648 165 sw
tri 3724 135 3754 165 se
rect 3754 159 3766 193
rect 3800 159 3810 193
rect 3754 135 3810 159
rect 3560 127 3810 135
rect 3368 123 3810 127
rect 3368 89 3378 123
rect 3412 89 3572 123
rect 3606 89 3669 123
rect 3703 89 3766 123
rect 3800 89 3810 123
rect 3368 73 3810 89
rect 4013 335 4069 351
rect 4013 301 4023 335
rect 4057 301 4069 335
rect 4013 263 4069 301
rect 4099 335 4369 351
rect 4099 306 4120 335
tri 4099 290 4115 306 ne
rect 4115 301 4120 306
rect 4154 301 4217 335
rect 4251 301 4314 335
rect 4348 301 4369 335
rect 4115 290 4369 301
rect 4399 335 4455 351
rect 4399 301 4411 335
rect 4445 301 4455 335
rect 4013 229 4023 263
rect 4057 229 4069 263
tri 4175 260 4205 290 ne
rect 4205 263 4264 290
rect 4013 195 4069 229
rect 4013 161 4023 195
rect 4057 161 4069 195
rect 4013 129 4069 161
tri 4099 244 4115 260 se
rect 4115 244 4159 260
tri 4159 244 4175 260 sw
rect 4099 210 4175 244
rect 4099 176 4120 210
rect 4154 176 4175 210
rect 4099 175 4175 176
tri 4099 159 4115 175 ne
rect 4115 159 4159 175
tri 4159 159 4175 175 nw
rect 4205 229 4217 263
rect 4251 229 4264 263
tri 4264 260 4294 290 nw
rect 4205 195 4264 229
rect 4205 161 4217 195
rect 4251 161 4264 195
tri 4294 244 4310 260 se
rect 4310 244 4353 260
tri 4353 244 4369 260 sw
rect 4294 216 4369 244
rect 4294 182 4315 216
rect 4349 182 4369 216
tri 4294 166 4310 182 ne
rect 4310 166 4353 182
tri 4353 166 4369 182 nw
tri 4069 129 4099 159 sw
tri 4175 129 4205 159 se
rect 4205 136 4264 161
tri 4264 136 4294 166 sw
tri 4369 136 4399 166 se
rect 4399 136 4455 301
rect 4205 129 4455 136
rect 4013 125 4455 129
rect 4013 91 4023 125
rect 4057 91 4217 125
rect 4251 91 4314 125
rect 4348 91 4411 125
rect 4445 91 4455 125
rect 4013 75 4455 91
rect 4515 335 4571 351
rect 4515 301 4525 335
rect 4559 301 4571 335
rect 4515 263 4571 301
rect 4601 314 4763 351
tri 4601 298 4617 314 ne
rect 4617 298 4763 314
tri 4677 268 4707 298 ne
rect 4515 229 4525 263
rect 4559 229 4571 263
rect 4515 195 4571 229
rect 4515 161 4525 195
rect 4559 161 4571 195
tri 4601 252 4617 268 se
rect 4617 252 4661 268
tri 4661 252 4677 268 sw
rect 4601 219 4677 252
rect 4601 185 4622 219
rect 4656 185 4677 219
rect 4601 183 4677 185
tri 4601 167 4617 183 ne
rect 4617 167 4661 183
tri 4661 167 4677 183 nw
rect 4707 263 4763 298
rect 4707 229 4719 263
rect 4753 229 4763 263
rect 4707 195 4763 229
rect 4515 137 4571 161
tri 4571 137 4601 167 sw
tri 4677 137 4707 167 se
rect 4707 161 4719 195
rect 4753 161 4763 195
rect 4707 137 4763 161
rect 4515 125 4763 137
rect 4515 91 4525 125
rect 4559 91 4622 125
rect 4656 91 4719 125
rect 4753 91 4763 125
rect 4515 75 4763 91
rect 4996 333 5052 349
rect 4996 299 5006 333
rect 5040 299 5052 333
rect 4996 261 5052 299
rect 5082 333 5246 349
rect 5082 304 5103 333
tri 5082 288 5098 304 ne
rect 5098 299 5103 304
rect 5137 299 5200 333
rect 5234 299 5246 333
rect 5098 288 5246 299
rect 5276 312 5438 349
tri 5276 296 5292 312 ne
rect 5292 296 5438 312
rect 4996 227 5006 261
rect 5040 227 5052 261
tri 5158 258 5188 288 ne
rect 5188 261 5246 288
tri 5352 266 5382 296 ne
rect 4996 193 5052 227
rect 4996 159 5006 193
rect 5040 159 5052 193
rect 4996 127 5052 159
tri 5082 242 5098 258 se
rect 5098 242 5142 258
tri 5142 242 5158 258 sw
rect 5082 208 5158 242
rect 5082 174 5103 208
rect 5137 174 5158 208
rect 5082 173 5158 174
tri 5082 157 5098 173 ne
rect 5098 157 5142 173
tri 5142 157 5158 173 nw
rect 5188 227 5200 261
rect 5234 227 5246 261
rect 5188 193 5246 227
rect 5188 159 5200 193
rect 5234 159 5246 193
tri 5276 250 5292 266 se
rect 5292 250 5336 266
tri 5336 250 5352 266 sw
rect 5276 217 5352 250
rect 5276 183 5297 217
rect 5331 183 5352 217
rect 5276 181 5352 183
tri 5276 165 5292 181 ne
rect 5292 165 5336 181
tri 5336 165 5352 181 nw
rect 5382 261 5438 296
rect 5382 227 5394 261
rect 5428 227 5438 261
rect 5382 193 5438 227
tri 5052 127 5082 157 sw
tri 5158 127 5188 157 se
rect 5188 135 5246 159
tri 5246 135 5276 165 sw
tri 5352 135 5382 165 se
rect 5382 159 5394 193
rect 5428 159 5438 193
rect 5382 135 5438 159
rect 5188 127 5438 135
rect 4996 123 5438 127
rect 4996 89 5006 123
rect 5040 89 5200 123
rect 5234 89 5297 123
rect 5331 89 5394 123
rect 5428 89 5438 123
rect 4996 73 5438 89
rect 5641 335 5697 351
rect 5641 301 5651 335
rect 5685 301 5697 335
rect 5641 263 5697 301
rect 5727 335 5997 351
rect 5727 306 5748 335
tri 5727 290 5743 306 ne
rect 5743 301 5748 306
rect 5782 301 5845 335
rect 5879 301 5942 335
rect 5976 301 5997 335
rect 5743 290 5997 301
rect 6027 335 6083 351
rect 6027 301 6039 335
rect 6073 301 6083 335
rect 5641 229 5651 263
rect 5685 229 5697 263
tri 5803 260 5833 290 ne
rect 5833 263 5892 290
rect 5641 195 5697 229
rect 5641 161 5651 195
rect 5685 161 5697 195
rect 5641 129 5697 161
tri 5727 244 5743 260 se
rect 5743 244 5787 260
tri 5787 244 5803 260 sw
rect 5727 210 5803 244
rect 5727 176 5748 210
rect 5782 176 5803 210
rect 5727 175 5803 176
tri 5727 159 5743 175 ne
rect 5743 159 5787 175
tri 5787 159 5803 175 nw
rect 5833 229 5845 263
rect 5879 229 5892 263
tri 5892 260 5922 290 nw
rect 5833 195 5892 229
rect 5833 161 5845 195
rect 5879 161 5892 195
tri 5922 244 5938 260 se
rect 5938 244 5981 260
tri 5981 244 5997 260 sw
rect 5922 216 5997 244
rect 5922 182 5943 216
rect 5977 182 5997 216
tri 5922 166 5938 182 ne
rect 5938 166 5981 182
tri 5981 166 5997 182 nw
tri 5697 129 5727 159 sw
tri 5803 129 5833 159 se
rect 5833 136 5892 161
tri 5892 136 5922 166 sw
tri 5997 136 6027 166 se
rect 6027 136 6083 301
rect 5833 129 6083 136
rect 5641 125 6083 129
rect 5641 91 5651 125
rect 5685 91 5845 125
rect 5879 91 5942 125
rect 5976 91 6039 125
rect 6073 91 6083 125
rect 5641 75 6083 91
rect 6143 335 6199 351
rect 6143 301 6153 335
rect 6187 301 6199 335
rect 6143 263 6199 301
rect 6229 314 6391 351
tri 6229 298 6245 314 ne
rect 6245 298 6391 314
tri 6305 268 6335 298 ne
rect 6143 229 6153 263
rect 6187 229 6199 263
rect 6143 195 6199 229
rect 6143 161 6153 195
rect 6187 161 6199 195
tri 6229 252 6245 268 se
rect 6245 252 6289 268
tri 6289 252 6305 268 sw
rect 6229 219 6305 252
rect 6229 185 6250 219
rect 6284 185 6305 219
rect 6229 183 6305 185
tri 6229 167 6245 183 ne
rect 6245 167 6289 183
tri 6289 167 6305 183 nw
rect 6335 263 6391 298
rect 6335 229 6347 263
rect 6381 229 6391 263
rect 6335 195 6391 229
rect 6143 137 6199 161
tri 6199 137 6229 167 sw
tri 6305 137 6335 167 se
rect 6335 161 6347 195
rect 6381 161 6391 195
rect 6335 137 6391 161
rect 6143 125 6391 137
rect 6143 91 6153 125
rect 6187 91 6250 125
rect 6284 91 6347 125
rect 6381 91 6391 125
rect 6143 75 6391 91
rect 6603 335 6659 351
rect 6603 301 6613 335
rect 6647 301 6659 335
rect 6603 263 6659 301
rect 6689 335 6959 351
rect 6689 306 6710 335
tri 6689 290 6705 306 ne
rect 6705 301 6710 306
rect 6744 301 6807 335
rect 6841 301 6904 335
rect 6938 301 6959 335
rect 6705 290 6959 301
rect 6989 335 7045 351
rect 6989 301 7001 335
rect 7035 301 7045 335
rect 6603 229 6613 263
rect 6647 229 6659 263
tri 6765 260 6795 290 ne
rect 6795 263 6854 290
rect 6603 195 6659 229
rect 6603 161 6613 195
rect 6647 161 6659 195
rect 6603 129 6659 161
tri 6689 244 6705 260 se
rect 6705 244 6749 260
tri 6749 244 6765 260 sw
rect 6689 210 6765 244
rect 6689 176 6710 210
rect 6744 176 6765 210
rect 6689 175 6765 176
tri 6689 159 6705 175 ne
rect 6705 159 6749 175
tri 6749 159 6765 175 nw
rect 6795 229 6807 263
rect 6841 229 6854 263
tri 6854 260 6884 290 nw
rect 6795 195 6854 229
rect 6795 161 6807 195
rect 6841 161 6854 195
tri 6884 244 6900 260 se
rect 6900 244 6943 260
tri 6943 244 6959 260 sw
rect 6884 216 6959 244
rect 6884 182 6905 216
rect 6939 182 6959 216
tri 6884 166 6900 182 ne
rect 6900 166 6943 182
tri 6943 166 6959 182 nw
tri 6659 129 6689 159 sw
tri 6765 129 6795 159 se
rect 6795 136 6854 161
tri 6854 136 6884 166 sw
tri 6959 136 6989 166 se
rect 6989 136 7045 301
rect 6795 129 7045 136
rect 6603 125 7045 129
rect 6603 91 6613 125
rect 6647 91 6807 125
rect 6841 91 6904 125
rect 6938 91 7001 125
rect 7035 91 7045 125
rect 6603 75 7045 91
rect 7105 335 7161 351
rect 7105 301 7115 335
rect 7149 301 7161 335
rect 7105 263 7161 301
rect 7191 314 7353 351
tri 7191 298 7207 314 ne
rect 7207 298 7353 314
tri 7267 268 7297 298 ne
rect 7105 229 7115 263
rect 7149 229 7161 263
rect 7105 195 7161 229
rect 7105 161 7115 195
rect 7149 161 7161 195
tri 7191 252 7207 268 se
rect 7207 252 7251 268
tri 7251 252 7267 268 sw
rect 7191 219 7267 252
rect 7191 185 7212 219
rect 7246 185 7267 219
rect 7191 183 7267 185
tri 7191 167 7207 183 ne
rect 7207 167 7251 183
tri 7251 167 7267 183 nw
rect 7297 263 7353 298
rect 7297 229 7309 263
rect 7343 229 7353 263
rect 7297 195 7353 229
rect 7105 137 7161 161
tri 7161 137 7191 167 sw
tri 7267 137 7297 167 se
rect 7297 161 7309 195
rect 7343 161 7353 195
rect 7297 137 7353 161
rect 7105 125 7353 137
rect 7105 91 7115 125
rect 7149 91 7212 125
rect 7246 91 7309 125
rect 7343 91 7353 125
rect 7105 75 7353 91
rect 7586 333 7642 349
rect 7586 299 7596 333
rect 7630 299 7642 333
rect 7586 261 7642 299
rect 7672 333 7836 349
rect 7672 304 7693 333
tri 7672 288 7688 304 ne
rect 7688 299 7693 304
rect 7727 299 7790 333
rect 7824 299 7836 333
rect 7688 288 7836 299
rect 7866 312 8028 349
tri 7866 296 7882 312 ne
rect 7882 296 8028 312
rect 7586 227 7596 261
rect 7630 227 7642 261
tri 7748 258 7778 288 ne
rect 7778 261 7836 288
tri 7942 266 7972 296 ne
rect 7586 193 7642 227
rect 7586 159 7596 193
rect 7630 159 7642 193
rect 7586 127 7642 159
tri 7672 242 7688 258 se
rect 7688 242 7732 258
tri 7732 242 7748 258 sw
rect 7672 208 7748 242
rect 7672 174 7693 208
rect 7727 174 7748 208
rect 7672 173 7748 174
tri 7672 157 7688 173 ne
rect 7688 157 7732 173
tri 7732 157 7748 173 nw
rect 7778 227 7790 261
rect 7824 227 7836 261
rect 7778 193 7836 227
rect 7778 159 7790 193
rect 7824 159 7836 193
tri 7866 250 7882 266 se
rect 7882 250 7926 266
tri 7926 250 7942 266 sw
rect 7866 217 7942 250
rect 7866 183 7887 217
rect 7921 183 7942 217
rect 7866 181 7942 183
tri 7866 165 7882 181 ne
rect 7882 165 7926 181
tri 7926 165 7942 181 nw
rect 7972 261 8028 296
rect 7972 227 7984 261
rect 8018 227 8028 261
rect 7972 193 8028 227
tri 7642 127 7672 157 sw
tri 7748 127 7778 157 se
rect 7778 135 7836 159
tri 7836 135 7866 165 sw
tri 7942 135 7972 165 se
rect 7972 159 7984 193
rect 8018 159 8028 193
rect 7972 135 8028 159
rect 7778 127 8028 135
rect 7586 123 8028 127
rect 7586 89 7596 123
rect 7630 89 7790 123
rect 7824 89 7887 123
rect 7921 89 7984 123
rect 8018 89 8028 123
rect 7586 73 8028 89
rect 8252 333 8308 349
rect 8252 299 8262 333
rect 8296 299 8308 333
rect 8252 261 8308 299
rect 8338 333 8502 349
rect 8338 304 8359 333
tri 8338 288 8354 304 ne
rect 8354 299 8359 304
rect 8393 299 8456 333
rect 8490 299 8502 333
rect 8354 288 8502 299
rect 8532 312 8694 349
tri 8532 296 8548 312 ne
rect 8548 296 8694 312
rect 8252 227 8262 261
rect 8296 227 8308 261
tri 8414 258 8444 288 ne
rect 8444 261 8502 288
tri 8608 266 8638 296 ne
rect 8252 193 8308 227
rect 8252 159 8262 193
rect 8296 159 8308 193
rect 8252 127 8308 159
tri 8338 242 8354 258 se
rect 8354 242 8398 258
tri 8398 242 8414 258 sw
rect 8338 208 8414 242
rect 8338 174 8359 208
rect 8393 174 8414 208
rect 8338 173 8414 174
tri 8338 157 8354 173 ne
rect 8354 157 8398 173
tri 8398 157 8414 173 nw
rect 8444 227 8456 261
rect 8490 227 8502 261
rect 8444 193 8502 227
rect 8444 159 8456 193
rect 8490 159 8502 193
tri 8532 250 8548 266 se
rect 8548 250 8592 266
tri 8592 250 8608 266 sw
rect 8532 217 8608 250
rect 8532 183 8553 217
rect 8587 183 8608 217
rect 8532 181 8608 183
tri 8532 165 8548 181 ne
rect 8548 165 8592 181
tri 8592 165 8608 181 nw
rect 8638 261 8694 296
rect 8638 227 8650 261
rect 8684 227 8694 261
rect 8638 193 8694 227
tri 8308 127 8338 157 sw
tri 8414 127 8444 157 se
rect 8444 135 8502 159
tri 8502 135 8532 165 sw
tri 8608 135 8638 165 se
rect 8638 159 8650 193
rect 8684 159 8694 193
rect 8638 135 8694 159
rect 8444 127 8694 135
rect 8252 123 8694 127
rect 8252 89 8262 123
rect 8296 89 8456 123
rect 8490 89 8553 123
rect 8587 89 8650 123
rect 8684 89 8694 123
rect 8252 73 8694 89
rect 8897 335 8953 351
rect 8897 301 8907 335
rect 8941 301 8953 335
rect 8897 263 8953 301
rect 8983 335 9253 351
rect 8983 306 9004 335
tri 8983 290 8999 306 ne
rect 8999 301 9004 306
rect 9038 301 9101 335
rect 9135 301 9198 335
rect 9232 301 9253 335
rect 8999 290 9253 301
rect 9283 335 9339 351
rect 9283 301 9295 335
rect 9329 301 9339 335
rect 8897 229 8907 263
rect 8941 229 8953 263
tri 9059 260 9089 290 ne
rect 9089 263 9148 290
rect 8897 195 8953 229
rect 8897 161 8907 195
rect 8941 161 8953 195
rect 8897 129 8953 161
tri 8983 244 8999 260 se
rect 8999 244 9043 260
tri 9043 244 9059 260 sw
rect 8983 210 9059 244
rect 8983 176 9004 210
rect 9038 176 9059 210
rect 8983 175 9059 176
tri 8983 159 8999 175 ne
rect 8999 159 9043 175
tri 9043 159 9059 175 nw
rect 9089 229 9101 263
rect 9135 229 9148 263
tri 9148 260 9178 290 nw
rect 9089 195 9148 229
rect 9089 161 9101 195
rect 9135 161 9148 195
tri 9178 244 9194 260 se
rect 9194 244 9237 260
tri 9237 244 9253 260 sw
rect 9178 216 9253 244
rect 9178 182 9199 216
rect 9233 182 9253 216
tri 9178 166 9194 182 ne
rect 9194 166 9237 182
tri 9237 166 9253 182 nw
tri 8953 129 8983 159 sw
tri 9059 129 9089 159 se
rect 9089 136 9148 161
tri 9148 136 9178 166 sw
tri 9253 136 9283 166 se
rect 9283 136 9339 301
rect 9089 129 9339 136
rect 8897 125 9339 129
rect 8897 91 8907 125
rect 8941 91 9101 125
rect 9135 91 9198 125
rect 9232 91 9295 125
rect 9329 91 9339 125
rect 8897 75 9339 91
rect 9399 335 9455 351
rect 9399 301 9409 335
rect 9443 301 9455 335
rect 9399 263 9455 301
rect 9485 314 9647 351
tri 9485 298 9501 314 ne
rect 9501 298 9647 314
tri 9561 268 9591 298 ne
rect 9399 229 9409 263
rect 9443 229 9455 263
rect 9399 195 9455 229
rect 9399 161 9409 195
rect 9443 161 9455 195
tri 9485 252 9501 268 se
rect 9501 252 9545 268
tri 9545 252 9561 268 sw
rect 9485 219 9561 252
rect 9485 185 9506 219
rect 9540 185 9561 219
rect 9485 183 9561 185
tri 9485 167 9501 183 ne
rect 9501 167 9545 183
tri 9545 167 9561 183 nw
rect 9591 263 9647 298
rect 9591 229 9603 263
rect 9637 229 9647 263
rect 9591 195 9647 229
rect 9399 137 9455 161
tri 9455 137 9485 167 sw
tri 9561 137 9591 167 se
rect 9591 161 9603 195
rect 9637 161 9647 195
rect 9591 137 9647 161
rect 9399 125 9647 137
rect 9399 91 9409 125
rect 9443 91 9506 125
rect 9540 91 9603 125
rect 9637 91 9647 125
rect 9399 75 9647 91
rect 9880 333 9936 349
rect 9880 299 9890 333
rect 9924 299 9936 333
rect 9880 261 9936 299
rect 9966 333 10130 349
rect 9966 304 9987 333
tri 9966 288 9982 304 ne
rect 9982 299 9987 304
rect 10021 299 10084 333
rect 10118 299 10130 333
rect 9982 288 10130 299
rect 10160 312 10322 349
tri 10160 296 10176 312 ne
rect 10176 296 10322 312
rect 9880 227 9890 261
rect 9924 227 9936 261
tri 10042 258 10072 288 ne
rect 10072 261 10130 288
tri 10236 266 10266 296 ne
rect 9880 193 9936 227
rect 9880 159 9890 193
rect 9924 159 9936 193
rect 9880 127 9936 159
tri 9966 242 9982 258 se
rect 9982 242 10026 258
tri 10026 242 10042 258 sw
rect 9966 208 10042 242
rect 9966 174 9987 208
rect 10021 174 10042 208
rect 9966 173 10042 174
tri 9966 157 9982 173 ne
rect 9982 157 10026 173
tri 10026 157 10042 173 nw
rect 10072 227 10084 261
rect 10118 227 10130 261
rect 10072 193 10130 227
rect 10072 159 10084 193
rect 10118 159 10130 193
tri 10160 250 10176 266 se
rect 10176 250 10220 266
tri 10220 250 10236 266 sw
rect 10160 217 10236 250
rect 10160 183 10181 217
rect 10215 183 10236 217
rect 10160 181 10236 183
tri 10160 165 10176 181 ne
rect 10176 165 10220 181
tri 10220 165 10236 181 nw
rect 10266 261 10322 296
rect 10266 227 10278 261
rect 10312 227 10322 261
rect 10266 193 10322 227
tri 9936 127 9966 157 sw
tri 10042 127 10072 157 se
rect 10072 135 10130 159
tri 10130 135 10160 165 sw
tri 10236 135 10266 165 se
rect 10266 159 10278 193
rect 10312 159 10322 193
rect 10266 135 10322 159
rect 10072 127 10322 135
rect 9880 123 10322 127
rect 9880 89 9890 123
rect 9924 89 10084 123
rect 10118 89 10181 123
rect 10215 89 10278 123
rect 10312 89 10322 123
rect 9880 73 10322 89
rect 10525 335 10581 351
rect 10525 301 10535 335
rect 10569 301 10581 335
rect 10525 263 10581 301
rect 10611 335 10881 351
rect 10611 306 10632 335
tri 10611 290 10627 306 ne
rect 10627 301 10632 306
rect 10666 301 10729 335
rect 10763 301 10826 335
rect 10860 301 10881 335
rect 10627 290 10881 301
rect 10911 335 10967 351
rect 10911 301 10923 335
rect 10957 301 10967 335
rect 10525 229 10535 263
rect 10569 229 10581 263
tri 10687 260 10717 290 ne
rect 10717 263 10776 290
rect 10525 195 10581 229
rect 10525 161 10535 195
rect 10569 161 10581 195
rect 10525 129 10581 161
tri 10611 244 10627 260 se
rect 10627 244 10671 260
tri 10671 244 10687 260 sw
rect 10611 210 10687 244
rect 10611 176 10632 210
rect 10666 176 10687 210
rect 10611 175 10687 176
tri 10611 159 10627 175 ne
rect 10627 159 10671 175
tri 10671 159 10687 175 nw
rect 10717 229 10729 263
rect 10763 229 10776 263
tri 10776 260 10806 290 nw
rect 10717 195 10776 229
rect 10717 161 10729 195
rect 10763 161 10776 195
tri 10806 244 10822 260 se
rect 10822 244 10865 260
tri 10865 244 10881 260 sw
rect 10806 216 10881 244
rect 10806 182 10827 216
rect 10861 182 10881 216
tri 10806 166 10822 182 ne
rect 10822 166 10865 182
tri 10865 166 10881 182 nw
tri 10581 129 10611 159 sw
tri 10687 129 10717 159 se
rect 10717 136 10776 161
tri 10776 136 10806 166 sw
tri 10881 136 10911 166 se
rect 10911 136 10967 301
rect 10717 129 10967 136
rect 10525 125 10967 129
rect 10525 91 10535 125
rect 10569 91 10729 125
rect 10763 91 10826 125
rect 10860 91 10923 125
rect 10957 91 10967 125
rect 10525 75 10967 91
rect 11027 335 11083 351
rect 11027 301 11037 335
rect 11071 301 11083 335
rect 11027 263 11083 301
rect 11113 314 11275 351
tri 11113 298 11129 314 ne
rect 11129 298 11275 314
tri 11189 268 11219 298 ne
rect 11027 229 11037 263
rect 11071 229 11083 263
rect 11027 195 11083 229
rect 11027 161 11037 195
rect 11071 161 11083 195
tri 11113 252 11129 268 se
rect 11129 252 11173 268
tri 11173 252 11189 268 sw
rect 11113 219 11189 252
rect 11113 185 11134 219
rect 11168 185 11189 219
rect 11113 183 11189 185
tri 11113 167 11129 183 ne
rect 11129 167 11173 183
tri 11173 167 11189 183 nw
rect 11219 263 11275 298
rect 11219 229 11231 263
rect 11265 229 11275 263
rect 11219 195 11275 229
rect 11027 137 11083 161
tri 11083 137 11113 167 sw
tri 11189 137 11219 167 se
rect 11219 161 11231 195
rect 11265 161 11275 195
rect 11219 137 11275 161
rect 11027 125 11275 137
rect 11027 91 11037 125
rect 11071 91 11134 125
rect 11168 91 11231 125
rect 11265 91 11275 125
rect 11027 75 11275 91
rect 11487 335 11543 351
rect 11487 301 11497 335
rect 11531 301 11543 335
rect 11487 263 11543 301
rect 11573 335 11843 351
rect 11573 306 11594 335
tri 11573 290 11589 306 ne
rect 11589 301 11594 306
rect 11628 301 11691 335
rect 11725 301 11788 335
rect 11822 301 11843 335
rect 11589 290 11843 301
rect 11873 335 11929 351
rect 11873 301 11885 335
rect 11919 301 11929 335
rect 11487 229 11497 263
rect 11531 229 11543 263
tri 11649 260 11679 290 ne
rect 11679 263 11738 290
rect 11487 195 11543 229
rect 11487 161 11497 195
rect 11531 161 11543 195
rect 11487 129 11543 161
tri 11573 244 11589 260 se
rect 11589 244 11633 260
tri 11633 244 11649 260 sw
rect 11573 210 11649 244
rect 11573 176 11594 210
rect 11628 176 11649 210
rect 11573 175 11649 176
tri 11573 159 11589 175 ne
rect 11589 159 11633 175
tri 11633 159 11649 175 nw
rect 11679 229 11691 263
rect 11725 229 11738 263
tri 11738 260 11768 290 nw
rect 11679 195 11738 229
rect 11679 161 11691 195
rect 11725 161 11738 195
tri 11768 244 11784 260 se
rect 11784 244 11827 260
tri 11827 244 11843 260 sw
rect 11768 216 11843 244
rect 11768 182 11789 216
rect 11823 182 11843 216
tri 11768 166 11784 182 ne
rect 11784 166 11827 182
tri 11827 166 11843 182 nw
tri 11543 129 11573 159 sw
tri 11649 129 11679 159 se
rect 11679 136 11738 161
tri 11738 136 11768 166 sw
tri 11843 136 11873 166 se
rect 11873 136 11929 301
rect 11679 129 11929 136
rect 11487 125 11929 129
rect 11487 91 11497 125
rect 11531 91 11691 125
rect 11725 91 11788 125
rect 11822 91 11885 125
rect 11919 91 11929 125
rect 11487 75 11929 91
rect 11989 335 12045 351
rect 11989 301 11999 335
rect 12033 301 12045 335
rect 11989 263 12045 301
rect 12075 314 12237 351
tri 12075 298 12091 314 ne
rect 12091 298 12237 314
tri 12151 268 12181 298 ne
rect 11989 229 11999 263
rect 12033 229 12045 263
rect 11989 195 12045 229
rect 11989 161 11999 195
rect 12033 161 12045 195
tri 12075 252 12091 268 se
rect 12091 252 12135 268
tri 12135 252 12151 268 sw
rect 12075 219 12151 252
rect 12075 185 12096 219
rect 12130 185 12151 219
rect 12075 183 12151 185
tri 12075 167 12091 183 ne
rect 12091 167 12135 183
tri 12135 167 12151 183 nw
rect 12181 263 12237 298
rect 12181 229 12193 263
rect 12227 229 12237 263
rect 12181 195 12237 229
rect 11989 137 12045 161
tri 12045 137 12075 167 sw
tri 12151 137 12181 167 se
rect 12181 161 12193 195
rect 12227 161 12237 195
rect 12181 137 12237 161
rect 11989 125 12237 137
rect 11989 91 11999 125
rect 12033 91 12096 125
rect 12130 91 12193 125
rect 12227 91 12237 125
rect 11989 75 12237 91
rect 12470 333 12526 349
rect 12470 299 12480 333
rect 12514 299 12526 333
rect 12470 261 12526 299
rect 12556 333 12720 349
rect 12556 304 12577 333
tri 12556 288 12572 304 ne
rect 12572 299 12577 304
rect 12611 299 12674 333
rect 12708 299 12720 333
rect 12572 288 12720 299
rect 12750 312 12912 349
tri 12750 296 12766 312 ne
rect 12766 296 12912 312
rect 12470 227 12480 261
rect 12514 227 12526 261
tri 12632 258 12662 288 ne
rect 12662 261 12720 288
tri 12826 266 12856 296 ne
rect 12470 193 12526 227
rect 12470 159 12480 193
rect 12514 159 12526 193
rect 12470 127 12526 159
tri 12556 242 12572 258 se
rect 12572 242 12616 258
tri 12616 242 12632 258 sw
rect 12556 208 12632 242
rect 12556 174 12577 208
rect 12611 174 12632 208
rect 12556 173 12632 174
tri 12556 157 12572 173 ne
rect 12572 157 12616 173
tri 12616 157 12632 173 nw
rect 12662 227 12674 261
rect 12708 227 12720 261
rect 12662 193 12720 227
rect 12662 159 12674 193
rect 12708 159 12720 193
tri 12750 250 12766 266 se
rect 12766 250 12810 266
tri 12810 250 12826 266 sw
rect 12750 217 12826 250
rect 12750 183 12771 217
rect 12805 183 12826 217
rect 12750 181 12826 183
tri 12750 165 12766 181 ne
rect 12766 165 12810 181
tri 12810 165 12826 181 nw
rect 12856 261 12912 296
rect 12856 227 12868 261
rect 12902 227 12912 261
rect 12856 193 12912 227
tri 12526 127 12556 157 sw
tri 12632 127 12662 157 se
rect 12662 135 12720 159
tri 12720 135 12750 165 sw
tri 12826 135 12856 165 se
rect 12856 159 12868 193
rect 12902 159 12912 193
rect 12856 135 12912 159
rect 12662 127 12912 135
rect 12470 123 12912 127
rect 12470 89 12480 123
rect 12514 89 12674 123
rect 12708 89 12771 123
rect 12805 89 12868 123
rect 12902 89 12912 123
rect 12470 73 12912 89
rect 13136 333 13192 349
rect 13136 299 13146 333
rect 13180 299 13192 333
rect 13136 261 13192 299
rect 13222 333 13386 349
rect 13222 304 13243 333
tri 13222 288 13238 304 ne
rect 13238 299 13243 304
rect 13277 299 13340 333
rect 13374 299 13386 333
rect 13238 288 13386 299
rect 13416 312 13578 349
tri 13416 296 13432 312 ne
rect 13432 296 13578 312
rect 13136 227 13146 261
rect 13180 227 13192 261
tri 13298 258 13328 288 ne
rect 13328 261 13386 288
tri 13492 266 13522 296 ne
rect 13136 193 13192 227
rect 13136 159 13146 193
rect 13180 159 13192 193
rect 13136 127 13192 159
tri 13222 242 13238 258 se
rect 13238 242 13282 258
tri 13282 242 13298 258 sw
rect 13222 208 13298 242
rect 13222 174 13243 208
rect 13277 174 13298 208
rect 13222 173 13298 174
tri 13222 157 13238 173 ne
rect 13238 157 13282 173
tri 13282 157 13298 173 nw
rect 13328 227 13340 261
rect 13374 227 13386 261
rect 13328 193 13386 227
rect 13328 159 13340 193
rect 13374 159 13386 193
tri 13416 250 13432 266 se
rect 13432 250 13476 266
tri 13476 250 13492 266 sw
rect 13416 217 13492 250
rect 13416 183 13437 217
rect 13471 183 13492 217
rect 13416 181 13492 183
tri 13416 165 13432 181 ne
rect 13432 165 13476 181
tri 13476 165 13492 181 nw
rect 13522 261 13578 296
rect 13522 227 13534 261
rect 13568 227 13578 261
rect 13522 193 13578 227
tri 13192 127 13222 157 sw
tri 13298 127 13328 157 se
rect 13328 135 13386 159
tri 13386 135 13416 165 sw
tri 13492 135 13522 165 se
rect 13522 159 13534 193
rect 13568 159 13578 193
rect 13522 135 13578 159
rect 13328 127 13578 135
rect 13136 123 13578 127
rect 13136 89 13146 123
rect 13180 89 13340 123
rect 13374 89 13437 123
rect 13471 89 13534 123
rect 13568 89 13578 123
rect 13136 73 13578 89
rect 13781 335 13837 351
rect 13781 301 13791 335
rect 13825 301 13837 335
rect 13781 263 13837 301
rect 13867 335 14137 351
rect 13867 306 13888 335
tri 13867 290 13883 306 ne
rect 13883 301 13888 306
rect 13922 301 13985 335
rect 14019 301 14082 335
rect 14116 301 14137 335
rect 13883 290 14137 301
rect 14167 335 14223 351
rect 14167 301 14179 335
rect 14213 301 14223 335
rect 13781 229 13791 263
rect 13825 229 13837 263
tri 13943 260 13973 290 ne
rect 13973 263 14032 290
rect 13781 195 13837 229
rect 13781 161 13791 195
rect 13825 161 13837 195
rect 13781 129 13837 161
tri 13867 244 13883 260 se
rect 13883 244 13927 260
tri 13927 244 13943 260 sw
rect 13867 210 13943 244
rect 13867 176 13888 210
rect 13922 176 13943 210
rect 13867 175 13943 176
tri 13867 159 13883 175 ne
rect 13883 159 13927 175
tri 13927 159 13943 175 nw
rect 13973 229 13985 263
rect 14019 229 14032 263
tri 14032 260 14062 290 nw
rect 13973 195 14032 229
rect 13973 161 13985 195
rect 14019 161 14032 195
tri 14062 244 14078 260 se
rect 14078 244 14121 260
tri 14121 244 14137 260 sw
rect 14062 216 14137 244
rect 14062 182 14083 216
rect 14117 182 14137 216
tri 14062 166 14078 182 ne
rect 14078 166 14121 182
tri 14121 166 14137 182 nw
tri 13837 129 13867 159 sw
tri 13943 129 13973 159 se
rect 13973 136 14032 161
tri 14032 136 14062 166 sw
tri 14137 136 14167 166 se
rect 14167 136 14223 301
rect 13973 129 14223 136
rect 13781 125 14223 129
rect 13781 91 13791 125
rect 13825 91 13985 125
rect 14019 91 14082 125
rect 14116 91 14179 125
rect 14213 91 14223 125
rect 13781 75 14223 91
rect 14283 335 14339 351
rect 14283 301 14293 335
rect 14327 301 14339 335
rect 14283 263 14339 301
rect 14369 314 14531 351
tri 14369 298 14385 314 ne
rect 14385 298 14531 314
tri 14445 268 14475 298 ne
rect 14283 229 14293 263
rect 14327 229 14339 263
rect 14283 195 14339 229
rect 14283 161 14293 195
rect 14327 161 14339 195
tri 14369 252 14385 268 se
rect 14385 252 14429 268
tri 14429 252 14445 268 sw
rect 14369 219 14445 252
rect 14369 185 14390 219
rect 14424 185 14445 219
rect 14369 183 14445 185
tri 14369 167 14385 183 ne
rect 14385 167 14429 183
tri 14429 167 14445 183 nw
rect 14475 263 14531 298
rect 14475 229 14487 263
rect 14521 229 14531 263
rect 14475 195 14531 229
rect 14283 137 14339 161
tri 14339 137 14369 167 sw
tri 14445 137 14475 167 se
rect 14475 161 14487 195
rect 14521 161 14531 195
rect 14475 137 14531 161
rect 14283 125 14531 137
rect 14283 91 14293 125
rect 14327 91 14390 125
rect 14424 91 14487 125
rect 14521 91 14531 125
rect 14283 75 14531 91
rect 14764 333 14820 349
rect 14764 299 14774 333
rect 14808 299 14820 333
rect 14764 261 14820 299
rect 14850 333 15014 349
rect 14850 304 14871 333
tri 14850 288 14866 304 ne
rect 14866 299 14871 304
rect 14905 299 14968 333
rect 15002 299 15014 333
rect 14866 288 15014 299
rect 15044 333 15204 349
rect 15044 312 15162 333
tri 15044 296 15060 312 ne
rect 15060 299 15162 312
rect 15196 299 15204 333
rect 15060 296 15204 299
rect 14764 227 14774 261
rect 14808 227 14820 261
tri 14926 258 14956 288 ne
rect 14956 261 15014 288
tri 15120 266 15150 296 ne
rect 14764 193 14820 227
rect 14764 159 14774 193
rect 14808 159 14820 193
rect 14764 127 14820 159
tri 14850 242 14866 258 se
rect 14866 242 14910 258
tri 14910 242 14926 258 sw
rect 14850 208 14926 242
rect 14850 174 14871 208
rect 14905 174 14926 208
rect 14850 173 14926 174
tri 14850 157 14866 173 ne
rect 14866 157 14910 173
tri 14910 157 14926 173 nw
rect 14956 227 14968 261
rect 15002 227 15014 261
rect 14956 193 15014 227
rect 14956 159 14968 193
rect 15002 159 15014 193
tri 15044 250 15060 266 se
rect 15060 250 15104 266
tri 15104 250 15120 266 sw
rect 15044 217 15120 250
rect 15044 183 15064 217
rect 15098 183 15120 217
rect 15044 181 15120 183
tri 15044 165 15060 181 ne
rect 15060 165 15104 181
tri 15104 165 15120 181 nw
rect 15150 261 15204 296
rect 15150 227 15162 261
rect 15196 227 15204 261
rect 15150 193 15204 227
tri 14820 127 14850 157 sw
tri 14926 127 14956 157 se
rect 14956 135 15014 159
tri 15014 135 15044 165 sw
tri 15120 135 15150 165 se
rect 15150 159 15162 193
rect 15196 159 15204 193
rect 15150 135 15204 159
rect 14956 127 15204 135
rect 14764 123 15204 127
rect 14764 89 14774 123
rect 14808 89 14968 123
rect 15002 89 15064 123
rect 15098 89 15162 123
rect 15196 89 15204 123
rect 14764 73 15204 89
rect 15430 333 15486 349
rect 15430 299 15440 333
rect 15474 299 15486 333
rect 15430 261 15486 299
rect 15516 333 15786 349
rect 15516 304 15537 333
tri 15516 288 15532 304 ne
rect 15532 299 15537 304
rect 15571 299 15634 333
rect 15668 312 15786 333
rect 15668 299 15770 312
rect 15532 296 15770 299
tri 15770 296 15786 312 nw
rect 15816 333 15872 349
rect 15816 299 15828 333
rect 15862 299 15872 333
rect 15532 288 15680 296
rect 15430 227 15440 261
rect 15474 227 15486 261
tri 15592 258 15622 288 ne
rect 15622 261 15680 288
tri 15680 266 15710 296 nw
rect 15430 193 15486 227
rect 15430 159 15440 193
rect 15474 159 15486 193
rect 15430 127 15486 159
tri 15516 242 15532 258 se
rect 15532 242 15576 258
tri 15576 242 15592 258 sw
rect 15516 208 15592 242
rect 15516 174 15537 208
rect 15571 174 15592 208
rect 15516 173 15592 174
tri 15516 157 15532 173 ne
rect 15532 157 15576 173
tri 15576 157 15592 173 nw
rect 15622 227 15634 261
rect 15668 227 15680 261
rect 15622 193 15680 227
rect 15622 159 15634 193
rect 15668 159 15680 193
tri 15710 250 15726 266 se
rect 15726 250 15770 266
tri 15770 250 15786 266 sw
rect 15710 217 15786 250
rect 15710 183 15731 217
rect 15765 183 15786 217
rect 15710 181 15786 183
tri 15710 165 15726 181 ne
rect 15726 165 15770 181
tri 15770 165 15786 181 nw
rect 15816 261 15872 299
rect 15816 227 15828 261
rect 15862 227 15872 261
rect 15816 193 15872 227
tri 15486 127 15516 157 sw
tri 15592 127 15622 157 se
rect 15622 135 15680 159
tri 15680 135 15710 165 sw
tri 15786 135 15816 165 se
rect 15816 159 15828 193
rect 15862 159 15872 193
rect 15816 135 15872 159
rect 15622 127 15872 135
rect 15430 123 15872 127
rect 15430 89 15440 123
rect 15474 89 15634 123
rect 15668 89 15731 123
rect 15765 89 15828 123
rect 15862 89 15872 123
rect 15430 73 15872 89
rect 16096 333 16152 349
rect 16096 299 16106 333
rect 16140 299 16152 333
rect 16096 261 16152 299
rect 16182 333 16346 349
rect 16182 304 16203 333
tri 16182 288 16198 304 ne
rect 16198 299 16203 304
rect 16237 299 16300 333
rect 16334 299 16346 333
rect 16198 288 16346 299
rect 16376 312 16538 349
tri 16376 296 16392 312 ne
rect 16392 296 16538 312
rect 16096 227 16106 261
rect 16140 227 16152 261
tri 16258 258 16288 288 ne
rect 16288 261 16346 288
tri 16452 266 16482 296 ne
rect 16096 193 16152 227
rect 16096 159 16106 193
rect 16140 159 16152 193
rect 16096 127 16152 159
tri 16182 242 16198 258 se
rect 16198 242 16242 258
tri 16242 242 16258 258 sw
rect 16182 208 16258 242
rect 16182 174 16203 208
rect 16237 174 16258 208
rect 16182 173 16258 174
tri 16182 157 16198 173 ne
rect 16198 157 16242 173
tri 16242 157 16258 173 nw
rect 16288 227 16300 261
rect 16334 227 16346 261
tri 16377 251 16392 266 se
rect 16392 251 16436 266
tri 16436 251 16451 266 sw
rect 16482 261 16538 296
rect 16288 193 16346 227
rect 16288 159 16300 193
rect 16334 159 16346 193
rect 16376 217 16452 251
rect 16376 183 16397 217
rect 16431 183 16452 217
rect 16376 181 16452 183
tri 16376 165 16392 181 ne
rect 16392 165 16436 181
tri 16436 165 16452 181 nw
rect 16482 227 16494 261
rect 16528 227 16538 261
rect 16482 193 16538 227
tri 16152 127 16182 157 sw
tri 16258 127 16288 157 se
rect 16288 135 16346 159
tri 16346 135 16376 165 sw
tri 16452 135 16482 165 se
rect 16482 159 16494 193
rect 16528 159 16538 193
rect 16482 135 16538 159
rect 16288 127 16538 135
rect 16096 123 16538 127
rect 16096 89 16106 123
rect 16140 89 16300 123
rect 16334 89 16397 123
rect 16431 89 16494 123
rect 16528 89 16538 123
rect 16096 73 16538 89
rect 16749 334 16805 350
rect 16749 300 16759 334
rect 16793 300 16805 334
rect 16749 262 16805 300
rect 16835 334 16995 350
rect 16835 313 16953 334
tri 16835 297 16851 313 ne
rect 16851 300 16953 313
rect 16987 300 16995 334
rect 16851 297 16995 300
tri 16911 267 16941 297 ne
rect 16749 228 16759 262
rect 16793 228 16805 262
rect 16749 194 16805 228
rect 16749 160 16759 194
rect 16793 160 16805 194
tri 16835 251 16851 267 se
rect 16851 251 16895 267
tri 16895 251 16911 267 sw
rect 16835 218 16911 251
rect 16835 184 16855 218
rect 16889 184 16911 218
rect 16835 182 16911 184
tri 16835 166 16851 182 ne
rect 16851 166 16895 182
tri 16895 166 16911 182 nw
rect 16941 262 16995 297
rect 16941 228 16953 262
rect 16987 228 16995 262
rect 16941 194 16995 228
rect 16749 136 16805 160
tri 16805 136 16835 166 sw
tri 16911 136 16941 166 se
rect 16941 160 16953 194
rect 16987 160 16995 194
rect 16941 136 16995 160
rect 16749 124 16995 136
rect 16749 90 16759 124
rect 16793 90 16855 124
rect 16889 90 16953 124
rect 16987 90 16995 124
rect 16749 74 16995 90
<< pdiff >>
rect 131 1366 187 1404
rect 131 1332 141 1366
rect 175 1332 187 1366
rect 131 1298 187 1332
rect 131 1264 141 1298
rect 175 1264 187 1298
rect 131 1230 187 1264
rect 131 1196 141 1230
rect 175 1196 187 1230
rect 131 1162 187 1196
rect 131 1128 141 1162
rect 175 1128 187 1162
rect 131 1093 187 1128
rect 131 1059 141 1093
rect 175 1059 187 1093
rect 131 1004 187 1059
rect 217 1366 275 1404
rect 217 1332 229 1366
rect 263 1332 275 1366
rect 217 1298 275 1332
rect 217 1264 229 1298
rect 263 1264 275 1298
rect 217 1230 275 1264
rect 217 1196 229 1230
rect 263 1196 275 1230
rect 217 1162 275 1196
rect 217 1128 229 1162
rect 263 1128 275 1162
rect 217 1093 275 1128
rect 217 1059 229 1093
rect 263 1059 275 1093
rect 217 1004 275 1059
rect 305 1366 363 1404
rect 305 1332 317 1366
rect 351 1332 363 1366
rect 305 1298 363 1332
rect 305 1264 317 1298
rect 351 1264 363 1298
rect 305 1230 363 1264
rect 305 1196 317 1230
rect 351 1196 363 1230
rect 305 1162 363 1196
rect 305 1128 317 1162
rect 351 1128 363 1162
rect 305 1004 363 1128
rect 393 1366 451 1404
rect 393 1332 405 1366
rect 439 1332 451 1366
rect 393 1298 451 1332
rect 393 1264 405 1298
rect 439 1264 451 1298
rect 393 1230 451 1264
rect 393 1196 405 1230
rect 439 1196 451 1230
rect 393 1162 451 1196
rect 393 1128 405 1162
rect 439 1128 451 1162
rect 393 1093 451 1128
rect 393 1059 405 1093
rect 439 1059 451 1093
rect 393 1004 451 1059
rect 481 1366 535 1404
rect 481 1332 493 1366
rect 527 1332 535 1366
rect 481 1298 535 1332
rect 481 1264 493 1298
rect 527 1264 535 1298
rect 481 1230 535 1264
rect 481 1196 493 1230
rect 527 1196 535 1230
rect 481 1162 535 1196
rect 481 1128 493 1162
rect 527 1128 535 1162
rect 481 1004 535 1128
rect 857 1366 913 1404
rect 857 1332 867 1366
rect 901 1332 913 1366
rect 857 1298 913 1332
rect 857 1264 867 1298
rect 901 1264 913 1298
rect 857 1230 913 1264
rect 857 1196 867 1230
rect 901 1196 913 1230
rect 857 1162 913 1196
rect 857 1128 867 1162
rect 901 1128 913 1162
rect 857 1093 913 1128
rect 857 1059 867 1093
rect 901 1059 913 1093
rect 857 1004 913 1059
rect 943 1366 1001 1404
rect 943 1332 955 1366
rect 989 1332 1001 1366
rect 943 1298 1001 1332
rect 943 1264 955 1298
rect 989 1264 1001 1298
rect 943 1230 1001 1264
rect 943 1196 955 1230
rect 989 1196 1001 1230
rect 943 1162 1001 1196
rect 943 1128 955 1162
rect 989 1128 1001 1162
rect 943 1093 1001 1128
rect 943 1059 955 1093
rect 989 1059 1001 1093
rect 943 1004 1001 1059
rect 1031 1366 1089 1404
rect 1031 1332 1043 1366
rect 1077 1332 1089 1366
rect 1031 1298 1089 1332
rect 1031 1264 1043 1298
rect 1077 1264 1089 1298
rect 1031 1230 1089 1264
rect 1031 1196 1043 1230
rect 1077 1196 1089 1230
rect 1031 1162 1089 1196
rect 1031 1128 1043 1162
rect 1077 1128 1089 1162
rect 1031 1004 1089 1128
rect 1119 1366 1177 1404
rect 1119 1332 1131 1366
rect 1165 1332 1177 1366
rect 1119 1298 1177 1332
rect 1119 1264 1131 1298
rect 1165 1264 1177 1298
rect 1119 1230 1177 1264
rect 1119 1196 1131 1230
rect 1165 1196 1177 1230
rect 1119 1162 1177 1196
rect 1119 1128 1131 1162
rect 1165 1128 1177 1162
rect 1119 1093 1177 1128
rect 1119 1059 1131 1093
rect 1165 1059 1177 1093
rect 1119 1004 1177 1059
rect 1207 1366 1265 1404
rect 1207 1332 1219 1366
rect 1253 1332 1265 1366
rect 1207 1298 1265 1332
rect 1207 1264 1219 1298
rect 1253 1264 1265 1298
rect 1207 1230 1265 1264
rect 1207 1196 1219 1230
rect 1253 1196 1265 1230
rect 1207 1162 1265 1196
rect 1207 1128 1219 1162
rect 1253 1128 1265 1162
rect 1207 1004 1265 1128
rect 1295 1366 1353 1404
rect 1295 1332 1307 1366
rect 1341 1332 1353 1366
rect 1295 1298 1353 1332
rect 1295 1264 1307 1298
rect 1341 1264 1353 1298
rect 1295 1230 1353 1264
rect 1295 1196 1307 1230
rect 1341 1196 1353 1230
rect 1295 1162 1353 1196
rect 1295 1128 1307 1162
rect 1341 1128 1353 1162
rect 1295 1093 1353 1128
rect 1295 1059 1307 1093
rect 1341 1059 1353 1093
rect 1295 1004 1353 1059
rect 1383 1366 1437 1404
rect 1383 1332 1395 1366
rect 1429 1332 1437 1366
rect 1383 1298 1437 1332
rect 1383 1264 1395 1298
rect 1429 1264 1437 1298
rect 1383 1230 1437 1264
rect 1383 1196 1395 1230
rect 1429 1196 1437 1230
rect 1383 1162 1437 1196
rect 1383 1128 1395 1162
rect 1429 1128 1437 1162
rect 1383 1004 1437 1128
rect 1819 1366 1875 1404
rect 1819 1332 1829 1366
rect 1863 1332 1875 1366
rect 1819 1298 1875 1332
rect 1819 1264 1829 1298
rect 1863 1264 1875 1298
rect 1819 1230 1875 1264
rect 1819 1196 1829 1230
rect 1863 1196 1875 1230
rect 1819 1162 1875 1196
rect 1819 1128 1829 1162
rect 1863 1128 1875 1162
rect 1819 1093 1875 1128
rect 1819 1059 1829 1093
rect 1863 1059 1875 1093
rect 1819 1004 1875 1059
rect 1905 1366 1963 1404
rect 1905 1332 1917 1366
rect 1951 1332 1963 1366
rect 1905 1298 1963 1332
rect 1905 1264 1917 1298
rect 1951 1264 1963 1298
rect 1905 1230 1963 1264
rect 1905 1196 1917 1230
rect 1951 1196 1963 1230
rect 1905 1162 1963 1196
rect 1905 1128 1917 1162
rect 1951 1128 1963 1162
rect 1905 1093 1963 1128
rect 1905 1059 1917 1093
rect 1951 1059 1963 1093
rect 1905 1004 1963 1059
rect 1993 1366 2051 1404
rect 1993 1332 2005 1366
rect 2039 1332 2051 1366
rect 1993 1298 2051 1332
rect 1993 1264 2005 1298
rect 2039 1264 2051 1298
rect 1993 1230 2051 1264
rect 1993 1196 2005 1230
rect 2039 1196 2051 1230
rect 1993 1162 2051 1196
rect 1993 1128 2005 1162
rect 2039 1128 2051 1162
rect 1993 1004 2051 1128
rect 2081 1366 2139 1404
rect 2081 1332 2093 1366
rect 2127 1332 2139 1366
rect 2081 1298 2139 1332
rect 2081 1264 2093 1298
rect 2127 1264 2139 1298
rect 2081 1230 2139 1264
rect 2081 1196 2093 1230
rect 2127 1196 2139 1230
rect 2081 1162 2139 1196
rect 2081 1128 2093 1162
rect 2127 1128 2139 1162
rect 2081 1093 2139 1128
rect 2081 1059 2093 1093
rect 2127 1059 2139 1093
rect 2081 1004 2139 1059
rect 2169 1366 2227 1404
rect 2169 1332 2181 1366
rect 2215 1332 2227 1366
rect 2169 1298 2227 1332
rect 2169 1264 2181 1298
rect 2215 1264 2227 1298
rect 2169 1230 2227 1264
rect 2169 1196 2181 1230
rect 2215 1196 2227 1230
rect 2169 1162 2227 1196
rect 2169 1128 2181 1162
rect 2215 1128 2227 1162
rect 2169 1004 2227 1128
rect 2257 1366 2315 1404
rect 2257 1332 2269 1366
rect 2303 1332 2315 1366
rect 2257 1298 2315 1332
rect 2257 1264 2269 1298
rect 2303 1264 2315 1298
rect 2257 1230 2315 1264
rect 2257 1196 2269 1230
rect 2303 1196 2315 1230
rect 2257 1162 2315 1196
rect 2257 1128 2269 1162
rect 2303 1128 2315 1162
rect 2257 1093 2315 1128
rect 2257 1059 2269 1093
rect 2303 1059 2315 1093
rect 2257 1004 2315 1059
rect 2345 1366 2399 1404
rect 2345 1332 2357 1366
rect 2391 1332 2399 1366
rect 2345 1298 2399 1332
rect 2345 1264 2357 1298
rect 2391 1264 2399 1298
rect 2345 1230 2399 1264
rect 2345 1196 2357 1230
rect 2391 1196 2399 1230
rect 2345 1162 2399 1196
rect 2345 1128 2357 1162
rect 2391 1128 2399 1162
rect 2345 1004 2399 1128
rect 2721 1366 2777 1404
rect 2721 1332 2731 1366
rect 2765 1332 2777 1366
rect 2721 1298 2777 1332
rect 2721 1264 2731 1298
rect 2765 1264 2777 1298
rect 2721 1230 2777 1264
rect 2721 1196 2731 1230
rect 2765 1196 2777 1230
rect 2721 1162 2777 1196
rect 2721 1128 2731 1162
rect 2765 1128 2777 1162
rect 2721 1093 2777 1128
rect 2721 1059 2731 1093
rect 2765 1059 2777 1093
rect 2721 1004 2777 1059
rect 2807 1366 2865 1404
rect 2807 1332 2819 1366
rect 2853 1332 2865 1366
rect 2807 1298 2865 1332
rect 2807 1264 2819 1298
rect 2853 1264 2865 1298
rect 2807 1230 2865 1264
rect 2807 1196 2819 1230
rect 2853 1196 2865 1230
rect 2807 1162 2865 1196
rect 2807 1128 2819 1162
rect 2853 1128 2865 1162
rect 2807 1093 2865 1128
rect 2807 1059 2819 1093
rect 2853 1059 2865 1093
rect 2807 1004 2865 1059
rect 2895 1366 2953 1404
rect 2895 1332 2907 1366
rect 2941 1332 2953 1366
rect 2895 1298 2953 1332
rect 2895 1264 2907 1298
rect 2941 1264 2953 1298
rect 2895 1230 2953 1264
rect 2895 1196 2907 1230
rect 2941 1196 2953 1230
rect 2895 1162 2953 1196
rect 2895 1128 2907 1162
rect 2941 1128 2953 1162
rect 2895 1004 2953 1128
rect 2983 1366 3041 1404
rect 2983 1332 2995 1366
rect 3029 1332 3041 1366
rect 2983 1298 3041 1332
rect 2983 1264 2995 1298
rect 3029 1264 3041 1298
rect 2983 1230 3041 1264
rect 2983 1196 2995 1230
rect 3029 1196 3041 1230
rect 2983 1162 3041 1196
rect 2983 1128 2995 1162
rect 3029 1128 3041 1162
rect 2983 1093 3041 1128
rect 2983 1059 2995 1093
rect 3029 1059 3041 1093
rect 2983 1004 3041 1059
rect 3071 1366 3125 1404
rect 3071 1332 3083 1366
rect 3117 1332 3125 1366
rect 3071 1298 3125 1332
rect 3071 1264 3083 1298
rect 3117 1264 3125 1298
rect 3071 1230 3125 1264
rect 3071 1196 3083 1230
rect 3117 1196 3125 1230
rect 3071 1162 3125 1196
rect 3071 1128 3083 1162
rect 3117 1128 3125 1162
rect 3071 1004 3125 1128
rect 3387 1366 3443 1404
rect 3387 1332 3397 1366
rect 3431 1332 3443 1366
rect 3387 1298 3443 1332
rect 3387 1264 3397 1298
rect 3431 1264 3443 1298
rect 3387 1230 3443 1264
rect 3387 1196 3397 1230
rect 3431 1196 3443 1230
rect 3387 1162 3443 1196
rect 3387 1128 3397 1162
rect 3431 1128 3443 1162
rect 3387 1093 3443 1128
rect 3387 1059 3397 1093
rect 3431 1059 3443 1093
rect 3387 1004 3443 1059
rect 3473 1366 3531 1404
rect 3473 1332 3485 1366
rect 3519 1332 3531 1366
rect 3473 1298 3531 1332
rect 3473 1264 3485 1298
rect 3519 1264 3531 1298
rect 3473 1230 3531 1264
rect 3473 1196 3485 1230
rect 3519 1196 3531 1230
rect 3473 1162 3531 1196
rect 3473 1128 3485 1162
rect 3519 1128 3531 1162
rect 3473 1093 3531 1128
rect 3473 1059 3485 1093
rect 3519 1059 3531 1093
rect 3473 1004 3531 1059
rect 3561 1366 3619 1404
rect 3561 1332 3573 1366
rect 3607 1332 3619 1366
rect 3561 1298 3619 1332
rect 3561 1264 3573 1298
rect 3607 1264 3619 1298
rect 3561 1230 3619 1264
rect 3561 1196 3573 1230
rect 3607 1196 3619 1230
rect 3561 1162 3619 1196
rect 3561 1128 3573 1162
rect 3607 1128 3619 1162
rect 3561 1004 3619 1128
rect 3649 1366 3707 1404
rect 3649 1332 3661 1366
rect 3695 1332 3707 1366
rect 3649 1298 3707 1332
rect 3649 1264 3661 1298
rect 3695 1264 3707 1298
rect 3649 1230 3707 1264
rect 3649 1196 3661 1230
rect 3695 1196 3707 1230
rect 3649 1162 3707 1196
rect 3649 1128 3661 1162
rect 3695 1128 3707 1162
rect 3649 1093 3707 1128
rect 3649 1059 3661 1093
rect 3695 1059 3707 1093
rect 3649 1004 3707 1059
rect 3737 1366 3791 1404
rect 3737 1332 3749 1366
rect 3783 1332 3791 1366
rect 3737 1298 3791 1332
rect 3737 1264 3749 1298
rect 3783 1264 3791 1298
rect 3737 1230 3791 1264
rect 3737 1196 3749 1230
rect 3783 1196 3791 1230
rect 3737 1162 3791 1196
rect 3737 1128 3749 1162
rect 3783 1128 3791 1162
rect 3737 1004 3791 1128
rect 4113 1366 4169 1404
rect 4113 1332 4123 1366
rect 4157 1332 4169 1366
rect 4113 1298 4169 1332
rect 4113 1264 4123 1298
rect 4157 1264 4169 1298
rect 4113 1230 4169 1264
rect 4113 1196 4123 1230
rect 4157 1196 4169 1230
rect 4113 1162 4169 1196
rect 4113 1128 4123 1162
rect 4157 1128 4169 1162
rect 4113 1093 4169 1128
rect 4113 1059 4123 1093
rect 4157 1059 4169 1093
rect 4113 1004 4169 1059
rect 4199 1366 4257 1404
rect 4199 1332 4211 1366
rect 4245 1332 4257 1366
rect 4199 1298 4257 1332
rect 4199 1264 4211 1298
rect 4245 1264 4257 1298
rect 4199 1230 4257 1264
rect 4199 1196 4211 1230
rect 4245 1196 4257 1230
rect 4199 1162 4257 1196
rect 4199 1128 4211 1162
rect 4245 1128 4257 1162
rect 4199 1093 4257 1128
rect 4199 1059 4211 1093
rect 4245 1059 4257 1093
rect 4199 1004 4257 1059
rect 4287 1366 4345 1404
rect 4287 1332 4299 1366
rect 4333 1332 4345 1366
rect 4287 1298 4345 1332
rect 4287 1264 4299 1298
rect 4333 1264 4345 1298
rect 4287 1230 4345 1264
rect 4287 1196 4299 1230
rect 4333 1196 4345 1230
rect 4287 1162 4345 1196
rect 4287 1128 4299 1162
rect 4333 1128 4345 1162
rect 4287 1004 4345 1128
rect 4375 1366 4433 1404
rect 4375 1332 4387 1366
rect 4421 1332 4433 1366
rect 4375 1298 4433 1332
rect 4375 1264 4387 1298
rect 4421 1264 4433 1298
rect 4375 1230 4433 1264
rect 4375 1196 4387 1230
rect 4421 1196 4433 1230
rect 4375 1162 4433 1196
rect 4375 1128 4387 1162
rect 4421 1128 4433 1162
rect 4375 1093 4433 1128
rect 4375 1059 4387 1093
rect 4421 1059 4433 1093
rect 4375 1004 4433 1059
rect 4463 1366 4521 1404
rect 4463 1332 4475 1366
rect 4509 1332 4521 1366
rect 4463 1298 4521 1332
rect 4463 1264 4475 1298
rect 4509 1264 4521 1298
rect 4463 1230 4521 1264
rect 4463 1196 4475 1230
rect 4509 1196 4521 1230
rect 4463 1162 4521 1196
rect 4463 1128 4475 1162
rect 4509 1128 4521 1162
rect 4463 1004 4521 1128
rect 4551 1366 4609 1404
rect 4551 1332 4563 1366
rect 4597 1332 4609 1366
rect 4551 1298 4609 1332
rect 4551 1264 4563 1298
rect 4597 1264 4609 1298
rect 4551 1230 4609 1264
rect 4551 1196 4563 1230
rect 4597 1196 4609 1230
rect 4551 1162 4609 1196
rect 4551 1128 4563 1162
rect 4597 1128 4609 1162
rect 4551 1093 4609 1128
rect 4551 1059 4563 1093
rect 4597 1059 4609 1093
rect 4551 1004 4609 1059
rect 4639 1366 4693 1404
rect 4639 1332 4651 1366
rect 4685 1332 4693 1366
rect 4639 1298 4693 1332
rect 4639 1264 4651 1298
rect 4685 1264 4693 1298
rect 4639 1230 4693 1264
rect 4639 1196 4651 1230
rect 4685 1196 4693 1230
rect 4639 1162 4693 1196
rect 4639 1128 4651 1162
rect 4685 1128 4693 1162
rect 4639 1004 4693 1128
rect 5015 1366 5071 1404
rect 5015 1332 5025 1366
rect 5059 1332 5071 1366
rect 5015 1298 5071 1332
rect 5015 1264 5025 1298
rect 5059 1264 5071 1298
rect 5015 1230 5071 1264
rect 5015 1196 5025 1230
rect 5059 1196 5071 1230
rect 5015 1162 5071 1196
rect 5015 1128 5025 1162
rect 5059 1128 5071 1162
rect 5015 1093 5071 1128
rect 5015 1059 5025 1093
rect 5059 1059 5071 1093
rect 5015 1004 5071 1059
rect 5101 1366 5159 1404
rect 5101 1332 5113 1366
rect 5147 1332 5159 1366
rect 5101 1298 5159 1332
rect 5101 1264 5113 1298
rect 5147 1264 5159 1298
rect 5101 1230 5159 1264
rect 5101 1196 5113 1230
rect 5147 1196 5159 1230
rect 5101 1162 5159 1196
rect 5101 1128 5113 1162
rect 5147 1128 5159 1162
rect 5101 1093 5159 1128
rect 5101 1059 5113 1093
rect 5147 1059 5159 1093
rect 5101 1004 5159 1059
rect 5189 1366 5247 1404
rect 5189 1332 5201 1366
rect 5235 1332 5247 1366
rect 5189 1298 5247 1332
rect 5189 1264 5201 1298
rect 5235 1264 5247 1298
rect 5189 1230 5247 1264
rect 5189 1196 5201 1230
rect 5235 1196 5247 1230
rect 5189 1162 5247 1196
rect 5189 1128 5201 1162
rect 5235 1128 5247 1162
rect 5189 1004 5247 1128
rect 5277 1366 5335 1404
rect 5277 1332 5289 1366
rect 5323 1332 5335 1366
rect 5277 1298 5335 1332
rect 5277 1264 5289 1298
rect 5323 1264 5335 1298
rect 5277 1230 5335 1264
rect 5277 1196 5289 1230
rect 5323 1196 5335 1230
rect 5277 1162 5335 1196
rect 5277 1128 5289 1162
rect 5323 1128 5335 1162
rect 5277 1093 5335 1128
rect 5277 1059 5289 1093
rect 5323 1059 5335 1093
rect 5277 1004 5335 1059
rect 5365 1366 5419 1404
rect 5365 1332 5377 1366
rect 5411 1332 5419 1366
rect 5365 1298 5419 1332
rect 5365 1264 5377 1298
rect 5411 1264 5419 1298
rect 5365 1230 5419 1264
rect 5365 1196 5377 1230
rect 5411 1196 5419 1230
rect 5365 1162 5419 1196
rect 5365 1128 5377 1162
rect 5411 1128 5419 1162
rect 5365 1004 5419 1128
rect 5741 1366 5797 1404
rect 5741 1332 5751 1366
rect 5785 1332 5797 1366
rect 5741 1298 5797 1332
rect 5741 1264 5751 1298
rect 5785 1264 5797 1298
rect 5741 1230 5797 1264
rect 5741 1196 5751 1230
rect 5785 1196 5797 1230
rect 5741 1162 5797 1196
rect 5741 1128 5751 1162
rect 5785 1128 5797 1162
rect 5741 1093 5797 1128
rect 5741 1059 5751 1093
rect 5785 1059 5797 1093
rect 5741 1004 5797 1059
rect 5827 1366 5885 1404
rect 5827 1332 5839 1366
rect 5873 1332 5885 1366
rect 5827 1298 5885 1332
rect 5827 1264 5839 1298
rect 5873 1264 5885 1298
rect 5827 1230 5885 1264
rect 5827 1196 5839 1230
rect 5873 1196 5885 1230
rect 5827 1162 5885 1196
rect 5827 1128 5839 1162
rect 5873 1128 5885 1162
rect 5827 1093 5885 1128
rect 5827 1059 5839 1093
rect 5873 1059 5885 1093
rect 5827 1004 5885 1059
rect 5915 1366 5973 1404
rect 5915 1332 5927 1366
rect 5961 1332 5973 1366
rect 5915 1298 5973 1332
rect 5915 1264 5927 1298
rect 5961 1264 5973 1298
rect 5915 1230 5973 1264
rect 5915 1196 5927 1230
rect 5961 1196 5973 1230
rect 5915 1162 5973 1196
rect 5915 1128 5927 1162
rect 5961 1128 5973 1162
rect 5915 1004 5973 1128
rect 6003 1366 6061 1404
rect 6003 1332 6015 1366
rect 6049 1332 6061 1366
rect 6003 1298 6061 1332
rect 6003 1264 6015 1298
rect 6049 1264 6061 1298
rect 6003 1230 6061 1264
rect 6003 1196 6015 1230
rect 6049 1196 6061 1230
rect 6003 1162 6061 1196
rect 6003 1128 6015 1162
rect 6049 1128 6061 1162
rect 6003 1093 6061 1128
rect 6003 1059 6015 1093
rect 6049 1059 6061 1093
rect 6003 1004 6061 1059
rect 6091 1366 6149 1404
rect 6091 1332 6103 1366
rect 6137 1332 6149 1366
rect 6091 1298 6149 1332
rect 6091 1264 6103 1298
rect 6137 1264 6149 1298
rect 6091 1230 6149 1264
rect 6091 1196 6103 1230
rect 6137 1196 6149 1230
rect 6091 1162 6149 1196
rect 6091 1128 6103 1162
rect 6137 1128 6149 1162
rect 6091 1004 6149 1128
rect 6179 1366 6237 1404
rect 6179 1332 6191 1366
rect 6225 1332 6237 1366
rect 6179 1298 6237 1332
rect 6179 1264 6191 1298
rect 6225 1264 6237 1298
rect 6179 1230 6237 1264
rect 6179 1196 6191 1230
rect 6225 1196 6237 1230
rect 6179 1162 6237 1196
rect 6179 1128 6191 1162
rect 6225 1128 6237 1162
rect 6179 1093 6237 1128
rect 6179 1059 6191 1093
rect 6225 1059 6237 1093
rect 6179 1004 6237 1059
rect 6267 1366 6321 1404
rect 6267 1332 6279 1366
rect 6313 1332 6321 1366
rect 6267 1298 6321 1332
rect 6267 1264 6279 1298
rect 6313 1264 6321 1298
rect 6267 1230 6321 1264
rect 6267 1196 6279 1230
rect 6313 1196 6321 1230
rect 6267 1162 6321 1196
rect 6267 1128 6279 1162
rect 6313 1128 6321 1162
rect 6267 1004 6321 1128
rect 6703 1366 6759 1404
rect 6703 1332 6713 1366
rect 6747 1332 6759 1366
rect 6703 1298 6759 1332
rect 6703 1264 6713 1298
rect 6747 1264 6759 1298
rect 6703 1230 6759 1264
rect 6703 1196 6713 1230
rect 6747 1196 6759 1230
rect 6703 1162 6759 1196
rect 6703 1128 6713 1162
rect 6747 1128 6759 1162
rect 6703 1093 6759 1128
rect 6703 1059 6713 1093
rect 6747 1059 6759 1093
rect 6703 1004 6759 1059
rect 6789 1366 6847 1404
rect 6789 1332 6801 1366
rect 6835 1332 6847 1366
rect 6789 1298 6847 1332
rect 6789 1264 6801 1298
rect 6835 1264 6847 1298
rect 6789 1230 6847 1264
rect 6789 1196 6801 1230
rect 6835 1196 6847 1230
rect 6789 1162 6847 1196
rect 6789 1128 6801 1162
rect 6835 1128 6847 1162
rect 6789 1093 6847 1128
rect 6789 1059 6801 1093
rect 6835 1059 6847 1093
rect 6789 1004 6847 1059
rect 6877 1366 6935 1404
rect 6877 1332 6889 1366
rect 6923 1332 6935 1366
rect 6877 1298 6935 1332
rect 6877 1264 6889 1298
rect 6923 1264 6935 1298
rect 6877 1230 6935 1264
rect 6877 1196 6889 1230
rect 6923 1196 6935 1230
rect 6877 1162 6935 1196
rect 6877 1128 6889 1162
rect 6923 1128 6935 1162
rect 6877 1004 6935 1128
rect 6965 1366 7023 1404
rect 6965 1332 6977 1366
rect 7011 1332 7023 1366
rect 6965 1298 7023 1332
rect 6965 1264 6977 1298
rect 7011 1264 7023 1298
rect 6965 1230 7023 1264
rect 6965 1196 6977 1230
rect 7011 1196 7023 1230
rect 6965 1162 7023 1196
rect 6965 1128 6977 1162
rect 7011 1128 7023 1162
rect 6965 1093 7023 1128
rect 6965 1059 6977 1093
rect 7011 1059 7023 1093
rect 6965 1004 7023 1059
rect 7053 1366 7111 1404
rect 7053 1332 7065 1366
rect 7099 1332 7111 1366
rect 7053 1298 7111 1332
rect 7053 1264 7065 1298
rect 7099 1264 7111 1298
rect 7053 1230 7111 1264
rect 7053 1196 7065 1230
rect 7099 1196 7111 1230
rect 7053 1162 7111 1196
rect 7053 1128 7065 1162
rect 7099 1128 7111 1162
rect 7053 1004 7111 1128
rect 7141 1366 7199 1404
rect 7141 1332 7153 1366
rect 7187 1332 7199 1366
rect 7141 1298 7199 1332
rect 7141 1264 7153 1298
rect 7187 1264 7199 1298
rect 7141 1230 7199 1264
rect 7141 1196 7153 1230
rect 7187 1196 7199 1230
rect 7141 1162 7199 1196
rect 7141 1128 7153 1162
rect 7187 1128 7199 1162
rect 7141 1093 7199 1128
rect 7141 1059 7153 1093
rect 7187 1059 7199 1093
rect 7141 1004 7199 1059
rect 7229 1366 7283 1404
rect 7229 1332 7241 1366
rect 7275 1332 7283 1366
rect 7229 1298 7283 1332
rect 7229 1264 7241 1298
rect 7275 1264 7283 1298
rect 7229 1230 7283 1264
rect 7229 1196 7241 1230
rect 7275 1196 7283 1230
rect 7229 1162 7283 1196
rect 7229 1128 7241 1162
rect 7275 1128 7283 1162
rect 7229 1004 7283 1128
rect 7605 1366 7661 1404
rect 7605 1332 7615 1366
rect 7649 1332 7661 1366
rect 7605 1298 7661 1332
rect 7605 1264 7615 1298
rect 7649 1264 7661 1298
rect 7605 1230 7661 1264
rect 7605 1196 7615 1230
rect 7649 1196 7661 1230
rect 7605 1162 7661 1196
rect 7605 1128 7615 1162
rect 7649 1128 7661 1162
rect 7605 1093 7661 1128
rect 7605 1059 7615 1093
rect 7649 1059 7661 1093
rect 7605 1004 7661 1059
rect 7691 1366 7749 1404
rect 7691 1332 7703 1366
rect 7737 1332 7749 1366
rect 7691 1298 7749 1332
rect 7691 1264 7703 1298
rect 7737 1264 7749 1298
rect 7691 1230 7749 1264
rect 7691 1196 7703 1230
rect 7737 1196 7749 1230
rect 7691 1162 7749 1196
rect 7691 1128 7703 1162
rect 7737 1128 7749 1162
rect 7691 1093 7749 1128
rect 7691 1059 7703 1093
rect 7737 1059 7749 1093
rect 7691 1004 7749 1059
rect 7779 1366 7837 1404
rect 7779 1332 7791 1366
rect 7825 1332 7837 1366
rect 7779 1298 7837 1332
rect 7779 1264 7791 1298
rect 7825 1264 7837 1298
rect 7779 1230 7837 1264
rect 7779 1196 7791 1230
rect 7825 1196 7837 1230
rect 7779 1162 7837 1196
rect 7779 1128 7791 1162
rect 7825 1128 7837 1162
rect 7779 1004 7837 1128
rect 7867 1366 7925 1404
rect 7867 1332 7879 1366
rect 7913 1332 7925 1366
rect 7867 1298 7925 1332
rect 7867 1264 7879 1298
rect 7913 1264 7925 1298
rect 7867 1230 7925 1264
rect 7867 1196 7879 1230
rect 7913 1196 7925 1230
rect 7867 1162 7925 1196
rect 7867 1128 7879 1162
rect 7913 1128 7925 1162
rect 7867 1093 7925 1128
rect 7867 1059 7879 1093
rect 7913 1059 7925 1093
rect 7867 1004 7925 1059
rect 7955 1366 8009 1404
rect 7955 1332 7967 1366
rect 8001 1332 8009 1366
rect 7955 1298 8009 1332
rect 7955 1264 7967 1298
rect 8001 1264 8009 1298
rect 7955 1230 8009 1264
rect 7955 1196 7967 1230
rect 8001 1196 8009 1230
rect 7955 1162 8009 1196
rect 7955 1128 7967 1162
rect 8001 1128 8009 1162
rect 7955 1004 8009 1128
rect 8271 1366 8327 1404
rect 8271 1332 8281 1366
rect 8315 1332 8327 1366
rect 8271 1298 8327 1332
rect 8271 1264 8281 1298
rect 8315 1264 8327 1298
rect 8271 1230 8327 1264
rect 8271 1196 8281 1230
rect 8315 1196 8327 1230
rect 8271 1162 8327 1196
rect 8271 1128 8281 1162
rect 8315 1128 8327 1162
rect 8271 1093 8327 1128
rect 8271 1059 8281 1093
rect 8315 1059 8327 1093
rect 8271 1004 8327 1059
rect 8357 1366 8415 1404
rect 8357 1332 8369 1366
rect 8403 1332 8415 1366
rect 8357 1298 8415 1332
rect 8357 1264 8369 1298
rect 8403 1264 8415 1298
rect 8357 1230 8415 1264
rect 8357 1196 8369 1230
rect 8403 1196 8415 1230
rect 8357 1162 8415 1196
rect 8357 1128 8369 1162
rect 8403 1128 8415 1162
rect 8357 1093 8415 1128
rect 8357 1059 8369 1093
rect 8403 1059 8415 1093
rect 8357 1004 8415 1059
rect 8445 1366 8503 1404
rect 8445 1332 8457 1366
rect 8491 1332 8503 1366
rect 8445 1298 8503 1332
rect 8445 1264 8457 1298
rect 8491 1264 8503 1298
rect 8445 1230 8503 1264
rect 8445 1196 8457 1230
rect 8491 1196 8503 1230
rect 8445 1162 8503 1196
rect 8445 1128 8457 1162
rect 8491 1128 8503 1162
rect 8445 1004 8503 1128
rect 8533 1366 8591 1404
rect 8533 1332 8545 1366
rect 8579 1332 8591 1366
rect 8533 1298 8591 1332
rect 8533 1264 8545 1298
rect 8579 1264 8591 1298
rect 8533 1230 8591 1264
rect 8533 1196 8545 1230
rect 8579 1196 8591 1230
rect 8533 1162 8591 1196
rect 8533 1128 8545 1162
rect 8579 1128 8591 1162
rect 8533 1093 8591 1128
rect 8533 1059 8545 1093
rect 8579 1059 8591 1093
rect 8533 1004 8591 1059
rect 8621 1366 8675 1404
rect 8621 1332 8633 1366
rect 8667 1332 8675 1366
rect 8621 1298 8675 1332
rect 8621 1264 8633 1298
rect 8667 1264 8675 1298
rect 8621 1230 8675 1264
rect 8621 1196 8633 1230
rect 8667 1196 8675 1230
rect 8621 1162 8675 1196
rect 8621 1128 8633 1162
rect 8667 1128 8675 1162
rect 8621 1004 8675 1128
rect 8997 1366 9053 1404
rect 8997 1332 9007 1366
rect 9041 1332 9053 1366
rect 8997 1298 9053 1332
rect 8997 1264 9007 1298
rect 9041 1264 9053 1298
rect 8997 1230 9053 1264
rect 8997 1196 9007 1230
rect 9041 1196 9053 1230
rect 8997 1162 9053 1196
rect 8997 1128 9007 1162
rect 9041 1128 9053 1162
rect 8997 1093 9053 1128
rect 8997 1059 9007 1093
rect 9041 1059 9053 1093
rect 8997 1004 9053 1059
rect 9083 1366 9141 1404
rect 9083 1332 9095 1366
rect 9129 1332 9141 1366
rect 9083 1298 9141 1332
rect 9083 1264 9095 1298
rect 9129 1264 9141 1298
rect 9083 1230 9141 1264
rect 9083 1196 9095 1230
rect 9129 1196 9141 1230
rect 9083 1162 9141 1196
rect 9083 1128 9095 1162
rect 9129 1128 9141 1162
rect 9083 1093 9141 1128
rect 9083 1059 9095 1093
rect 9129 1059 9141 1093
rect 9083 1004 9141 1059
rect 9171 1366 9229 1404
rect 9171 1332 9183 1366
rect 9217 1332 9229 1366
rect 9171 1298 9229 1332
rect 9171 1264 9183 1298
rect 9217 1264 9229 1298
rect 9171 1230 9229 1264
rect 9171 1196 9183 1230
rect 9217 1196 9229 1230
rect 9171 1162 9229 1196
rect 9171 1128 9183 1162
rect 9217 1128 9229 1162
rect 9171 1004 9229 1128
rect 9259 1366 9317 1404
rect 9259 1332 9271 1366
rect 9305 1332 9317 1366
rect 9259 1298 9317 1332
rect 9259 1264 9271 1298
rect 9305 1264 9317 1298
rect 9259 1230 9317 1264
rect 9259 1196 9271 1230
rect 9305 1196 9317 1230
rect 9259 1162 9317 1196
rect 9259 1128 9271 1162
rect 9305 1128 9317 1162
rect 9259 1093 9317 1128
rect 9259 1059 9271 1093
rect 9305 1059 9317 1093
rect 9259 1004 9317 1059
rect 9347 1366 9405 1404
rect 9347 1332 9359 1366
rect 9393 1332 9405 1366
rect 9347 1298 9405 1332
rect 9347 1264 9359 1298
rect 9393 1264 9405 1298
rect 9347 1230 9405 1264
rect 9347 1196 9359 1230
rect 9393 1196 9405 1230
rect 9347 1162 9405 1196
rect 9347 1128 9359 1162
rect 9393 1128 9405 1162
rect 9347 1004 9405 1128
rect 9435 1366 9493 1404
rect 9435 1332 9447 1366
rect 9481 1332 9493 1366
rect 9435 1298 9493 1332
rect 9435 1264 9447 1298
rect 9481 1264 9493 1298
rect 9435 1230 9493 1264
rect 9435 1196 9447 1230
rect 9481 1196 9493 1230
rect 9435 1162 9493 1196
rect 9435 1128 9447 1162
rect 9481 1128 9493 1162
rect 9435 1093 9493 1128
rect 9435 1059 9447 1093
rect 9481 1059 9493 1093
rect 9435 1004 9493 1059
rect 9523 1366 9577 1404
rect 9523 1332 9535 1366
rect 9569 1332 9577 1366
rect 9523 1298 9577 1332
rect 9523 1264 9535 1298
rect 9569 1264 9577 1298
rect 9523 1230 9577 1264
rect 9523 1196 9535 1230
rect 9569 1196 9577 1230
rect 9523 1162 9577 1196
rect 9523 1128 9535 1162
rect 9569 1128 9577 1162
rect 9523 1004 9577 1128
rect 9899 1366 9955 1404
rect 9899 1332 9909 1366
rect 9943 1332 9955 1366
rect 9899 1298 9955 1332
rect 9899 1264 9909 1298
rect 9943 1264 9955 1298
rect 9899 1230 9955 1264
rect 9899 1196 9909 1230
rect 9943 1196 9955 1230
rect 9899 1162 9955 1196
rect 9899 1128 9909 1162
rect 9943 1128 9955 1162
rect 9899 1093 9955 1128
rect 9899 1059 9909 1093
rect 9943 1059 9955 1093
rect 9899 1004 9955 1059
rect 9985 1366 10043 1404
rect 9985 1332 9997 1366
rect 10031 1332 10043 1366
rect 9985 1298 10043 1332
rect 9985 1264 9997 1298
rect 10031 1264 10043 1298
rect 9985 1230 10043 1264
rect 9985 1196 9997 1230
rect 10031 1196 10043 1230
rect 9985 1162 10043 1196
rect 9985 1128 9997 1162
rect 10031 1128 10043 1162
rect 9985 1093 10043 1128
rect 9985 1059 9997 1093
rect 10031 1059 10043 1093
rect 9985 1004 10043 1059
rect 10073 1366 10131 1404
rect 10073 1332 10085 1366
rect 10119 1332 10131 1366
rect 10073 1298 10131 1332
rect 10073 1264 10085 1298
rect 10119 1264 10131 1298
rect 10073 1230 10131 1264
rect 10073 1196 10085 1230
rect 10119 1196 10131 1230
rect 10073 1162 10131 1196
rect 10073 1128 10085 1162
rect 10119 1128 10131 1162
rect 10073 1004 10131 1128
rect 10161 1366 10219 1404
rect 10161 1332 10173 1366
rect 10207 1332 10219 1366
rect 10161 1298 10219 1332
rect 10161 1264 10173 1298
rect 10207 1264 10219 1298
rect 10161 1230 10219 1264
rect 10161 1196 10173 1230
rect 10207 1196 10219 1230
rect 10161 1162 10219 1196
rect 10161 1128 10173 1162
rect 10207 1128 10219 1162
rect 10161 1093 10219 1128
rect 10161 1059 10173 1093
rect 10207 1059 10219 1093
rect 10161 1004 10219 1059
rect 10249 1366 10303 1404
rect 10249 1332 10261 1366
rect 10295 1332 10303 1366
rect 10249 1298 10303 1332
rect 10249 1264 10261 1298
rect 10295 1264 10303 1298
rect 10249 1230 10303 1264
rect 10249 1196 10261 1230
rect 10295 1196 10303 1230
rect 10249 1162 10303 1196
rect 10249 1128 10261 1162
rect 10295 1128 10303 1162
rect 10249 1004 10303 1128
rect 10625 1366 10681 1404
rect 10625 1332 10635 1366
rect 10669 1332 10681 1366
rect 10625 1298 10681 1332
rect 10625 1264 10635 1298
rect 10669 1264 10681 1298
rect 10625 1230 10681 1264
rect 10625 1196 10635 1230
rect 10669 1196 10681 1230
rect 10625 1162 10681 1196
rect 10625 1128 10635 1162
rect 10669 1128 10681 1162
rect 10625 1093 10681 1128
rect 10625 1059 10635 1093
rect 10669 1059 10681 1093
rect 10625 1004 10681 1059
rect 10711 1366 10769 1404
rect 10711 1332 10723 1366
rect 10757 1332 10769 1366
rect 10711 1298 10769 1332
rect 10711 1264 10723 1298
rect 10757 1264 10769 1298
rect 10711 1230 10769 1264
rect 10711 1196 10723 1230
rect 10757 1196 10769 1230
rect 10711 1162 10769 1196
rect 10711 1128 10723 1162
rect 10757 1128 10769 1162
rect 10711 1093 10769 1128
rect 10711 1059 10723 1093
rect 10757 1059 10769 1093
rect 10711 1004 10769 1059
rect 10799 1366 10857 1404
rect 10799 1332 10811 1366
rect 10845 1332 10857 1366
rect 10799 1298 10857 1332
rect 10799 1264 10811 1298
rect 10845 1264 10857 1298
rect 10799 1230 10857 1264
rect 10799 1196 10811 1230
rect 10845 1196 10857 1230
rect 10799 1162 10857 1196
rect 10799 1128 10811 1162
rect 10845 1128 10857 1162
rect 10799 1004 10857 1128
rect 10887 1366 10945 1404
rect 10887 1332 10899 1366
rect 10933 1332 10945 1366
rect 10887 1298 10945 1332
rect 10887 1264 10899 1298
rect 10933 1264 10945 1298
rect 10887 1230 10945 1264
rect 10887 1196 10899 1230
rect 10933 1196 10945 1230
rect 10887 1162 10945 1196
rect 10887 1128 10899 1162
rect 10933 1128 10945 1162
rect 10887 1093 10945 1128
rect 10887 1059 10899 1093
rect 10933 1059 10945 1093
rect 10887 1004 10945 1059
rect 10975 1366 11033 1404
rect 10975 1332 10987 1366
rect 11021 1332 11033 1366
rect 10975 1298 11033 1332
rect 10975 1264 10987 1298
rect 11021 1264 11033 1298
rect 10975 1230 11033 1264
rect 10975 1196 10987 1230
rect 11021 1196 11033 1230
rect 10975 1162 11033 1196
rect 10975 1128 10987 1162
rect 11021 1128 11033 1162
rect 10975 1004 11033 1128
rect 11063 1366 11121 1404
rect 11063 1332 11075 1366
rect 11109 1332 11121 1366
rect 11063 1298 11121 1332
rect 11063 1264 11075 1298
rect 11109 1264 11121 1298
rect 11063 1230 11121 1264
rect 11063 1196 11075 1230
rect 11109 1196 11121 1230
rect 11063 1162 11121 1196
rect 11063 1128 11075 1162
rect 11109 1128 11121 1162
rect 11063 1093 11121 1128
rect 11063 1059 11075 1093
rect 11109 1059 11121 1093
rect 11063 1004 11121 1059
rect 11151 1366 11205 1404
rect 11151 1332 11163 1366
rect 11197 1332 11205 1366
rect 11151 1298 11205 1332
rect 11151 1264 11163 1298
rect 11197 1264 11205 1298
rect 11151 1230 11205 1264
rect 11151 1196 11163 1230
rect 11197 1196 11205 1230
rect 11151 1162 11205 1196
rect 11151 1128 11163 1162
rect 11197 1128 11205 1162
rect 11151 1004 11205 1128
rect 11587 1366 11643 1404
rect 11587 1332 11597 1366
rect 11631 1332 11643 1366
rect 11587 1298 11643 1332
rect 11587 1264 11597 1298
rect 11631 1264 11643 1298
rect 11587 1230 11643 1264
rect 11587 1196 11597 1230
rect 11631 1196 11643 1230
rect 11587 1162 11643 1196
rect 11587 1128 11597 1162
rect 11631 1128 11643 1162
rect 11587 1093 11643 1128
rect 11587 1059 11597 1093
rect 11631 1059 11643 1093
rect 11587 1004 11643 1059
rect 11673 1366 11731 1404
rect 11673 1332 11685 1366
rect 11719 1332 11731 1366
rect 11673 1298 11731 1332
rect 11673 1264 11685 1298
rect 11719 1264 11731 1298
rect 11673 1230 11731 1264
rect 11673 1196 11685 1230
rect 11719 1196 11731 1230
rect 11673 1162 11731 1196
rect 11673 1128 11685 1162
rect 11719 1128 11731 1162
rect 11673 1093 11731 1128
rect 11673 1059 11685 1093
rect 11719 1059 11731 1093
rect 11673 1004 11731 1059
rect 11761 1366 11819 1404
rect 11761 1332 11773 1366
rect 11807 1332 11819 1366
rect 11761 1298 11819 1332
rect 11761 1264 11773 1298
rect 11807 1264 11819 1298
rect 11761 1230 11819 1264
rect 11761 1196 11773 1230
rect 11807 1196 11819 1230
rect 11761 1162 11819 1196
rect 11761 1128 11773 1162
rect 11807 1128 11819 1162
rect 11761 1004 11819 1128
rect 11849 1366 11907 1404
rect 11849 1332 11861 1366
rect 11895 1332 11907 1366
rect 11849 1298 11907 1332
rect 11849 1264 11861 1298
rect 11895 1264 11907 1298
rect 11849 1230 11907 1264
rect 11849 1196 11861 1230
rect 11895 1196 11907 1230
rect 11849 1162 11907 1196
rect 11849 1128 11861 1162
rect 11895 1128 11907 1162
rect 11849 1093 11907 1128
rect 11849 1059 11861 1093
rect 11895 1059 11907 1093
rect 11849 1004 11907 1059
rect 11937 1366 11995 1404
rect 11937 1332 11949 1366
rect 11983 1332 11995 1366
rect 11937 1298 11995 1332
rect 11937 1264 11949 1298
rect 11983 1264 11995 1298
rect 11937 1230 11995 1264
rect 11937 1196 11949 1230
rect 11983 1196 11995 1230
rect 11937 1162 11995 1196
rect 11937 1128 11949 1162
rect 11983 1128 11995 1162
rect 11937 1004 11995 1128
rect 12025 1366 12083 1404
rect 12025 1332 12037 1366
rect 12071 1332 12083 1366
rect 12025 1298 12083 1332
rect 12025 1264 12037 1298
rect 12071 1264 12083 1298
rect 12025 1230 12083 1264
rect 12025 1196 12037 1230
rect 12071 1196 12083 1230
rect 12025 1162 12083 1196
rect 12025 1128 12037 1162
rect 12071 1128 12083 1162
rect 12025 1093 12083 1128
rect 12025 1059 12037 1093
rect 12071 1059 12083 1093
rect 12025 1004 12083 1059
rect 12113 1366 12167 1404
rect 12113 1332 12125 1366
rect 12159 1332 12167 1366
rect 12113 1298 12167 1332
rect 12113 1264 12125 1298
rect 12159 1264 12167 1298
rect 12113 1230 12167 1264
rect 12113 1196 12125 1230
rect 12159 1196 12167 1230
rect 12113 1162 12167 1196
rect 12113 1128 12125 1162
rect 12159 1128 12167 1162
rect 12113 1004 12167 1128
rect 12489 1366 12545 1404
rect 12489 1332 12499 1366
rect 12533 1332 12545 1366
rect 12489 1298 12545 1332
rect 12489 1264 12499 1298
rect 12533 1264 12545 1298
rect 12489 1230 12545 1264
rect 12489 1196 12499 1230
rect 12533 1196 12545 1230
rect 12489 1162 12545 1196
rect 12489 1128 12499 1162
rect 12533 1128 12545 1162
rect 12489 1093 12545 1128
rect 12489 1059 12499 1093
rect 12533 1059 12545 1093
rect 12489 1004 12545 1059
rect 12575 1366 12633 1404
rect 12575 1332 12587 1366
rect 12621 1332 12633 1366
rect 12575 1298 12633 1332
rect 12575 1264 12587 1298
rect 12621 1264 12633 1298
rect 12575 1230 12633 1264
rect 12575 1196 12587 1230
rect 12621 1196 12633 1230
rect 12575 1162 12633 1196
rect 12575 1128 12587 1162
rect 12621 1128 12633 1162
rect 12575 1093 12633 1128
rect 12575 1059 12587 1093
rect 12621 1059 12633 1093
rect 12575 1004 12633 1059
rect 12663 1366 12721 1404
rect 12663 1332 12675 1366
rect 12709 1332 12721 1366
rect 12663 1298 12721 1332
rect 12663 1264 12675 1298
rect 12709 1264 12721 1298
rect 12663 1230 12721 1264
rect 12663 1196 12675 1230
rect 12709 1196 12721 1230
rect 12663 1162 12721 1196
rect 12663 1128 12675 1162
rect 12709 1128 12721 1162
rect 12663 1004 12721 1128
rect 12751 1366 12809 1404
rect 12751 1332 12763 1366
rect 12797 1332 12809 1366
rect 12751 1298 12809 1332
rect 12751 1264 12763 1298
rect 12797 1264 12809 1298
rect 12751 1230 12809 1264
rect 12751 1196 12763 1230
rect 12797 1196 12809 1230
rect 12751 1162 12809 1196
rect 12751 1128 12763 1162
rect 12797 1128 12809 1162
rect 12751 1093 12809 1128
rect 12751 1059 12763 1093
rect 12797 1059 12809 1093
rect 12751 1004 12809 1059
rect 12839 1366 12893 1404
rect 12839 1332 12851 1366
rect 12885 1332 12893 1366
rect 12839 1298 12893 1332
rect 12839 1264 12851 1298
rect 12885 1264 12893 1298
rect 12839 1230 12893 1264
rect 12839 1196 12851 1230
rect 12885 1196 12893 1230
rect 12839 1162 12893 1196
rect 12839 1128 12851 1162
rect 12885 1128 12893 1162
rect 12839 1004 12893 1128
rect 13155 1366 13211 1404
rect 13155 1332 13165 1366
rect 13199 1332 13211 1366
rect 13155 1298 13211 1332
rect 13155 1264 13165 1298
rect 13199 1264 13211 1298
rect 13155 1230 13211 1264
rect 13155 1196 13165 1230
rect 13199 1196 13211 1230
rect 13155 1162 13211 1196
rect 13155 1128 13165 1162
rect 13199 1128 13211 1162
rect 13155 1093 13211 1128
rect 13155 1059 13165 1093
rect 13199 1059 13211 1093
rect 13155 1004 13211 1059
rect 13241 1366 13299 1404
rect 13241 1332 13253 1366
rect 13287 1332 13299 1366
rect 13241 1298 13299 1332
rect 13241 1264 13253 1298
rect 13287 1264 13299 1298
rect 13241 1230 13299 1264
rect 13241 1196 13253 1230
rect 13287 1196 13299 1230
rect 13241 1162 13299 1196
rect 13241 1128 13253 1162
rect 13287 1128 13299 1162
rect 13241 1093 13299 1128
rect 13241 1059 13253 1093
rect 13287 1059 13299 1093
rect 13241 1004 13299 1059
rect 13329 1366 13387 1404
rect 13329 1332 13341 1366
rect 13375 1332 13387 1366
rect 13329 1298 13387 1332
rect 13329 1264 13341 1298
rect 13375 1264 13387 1298
rect 13329 1230 13387 1264
rect 13329 1196 13341 1230
rect 13375 1196 13387 1230
rect 13329 1162 13387 1196
rect 13329 1128 13341 1162
rect 13375 1128 13387 1162
rect 13329 1004 13387 1128
rect 13417 1366 13475 1404
rect 13417 1332 13429 1366
rect 13463 1332 13475 1366
rect 13417 1298 13475 1332
rect 13417 1264 13429 1298
rect 13463 1264 13475 1298
rect 13417 1230 13475 1264
rect 13417 1196 13429 1230
rect 13463 1196 13475 1230
rect 13417 1162 13475 1196
rect 13417 1128 13429 1162
rect 13463 1128 13475 1162
rect 13417 1093 13475 1128
rect 13417 1059 13429 1093
rect 13463 1059 13475 1093
rect 13417 1004 13475 1059
rect 13505 1366 13559 1404
rect 13505 1332 13517 1366
rect 13551 1332 13559 1366
rect 13505 1298 13559 1332
rect 13505 1264 13517 1298
rect 13551 1264 13559 1298
rect 13505 1230 13559 1264
rect 13505 1196 13517 1230
rect 13551 1196 13559 1230
rect 13505 1162 13559 1196
rect 13505 1128 13517 1162
rect 13551 1128 13559 1162
rect 13505 1004 13559 1128
rect 13881 1366 13937 1404
rect 13881 1332 13891 1366
rect 13925 1332 13937 1366
rect 13881 1298 13937 1332
rect 13881 1264 13891 1298
rect 13925 1264 13937 1298
rect 13881 1230 13937 1264
rect 13881 1196 13891 1230
rect 13925 1196 13937 1230
rect 13881 1162 13937 1196
rect 13881 1128 13891 1162
rect 13925 1128 13937 1162
rect 13881 1093 13937 1128
rect 13881 1059 13891 1093
rect 13925 1059 13937 1093
rect 13881 1004 13937 1059
rect 13967 1366 14025 1404
rect 13967 1332 13979 1366
rect 14013 1332 14025 1366
rect 13967 1298 14025 1332
rect 13967 1264 13979 1298
rect 14013 1264 14025 1298
rect 13967 1230 14025 1264
rect 13967 1196 13979 1230
rect 14013 1196 14025 1230
rect 13967 1162 14025 1196
rect 13967 1128 13979 1162
rect 14013 1128 14025 1162
rect 13967 1093 14025 1128
rect 13967 1059 13979 1093
rect 14013 1059 14025 1093
rect 13967 1004 14025 1059
rect 14055 1366 14113 1404
rect 14055 1332 14067 1366
rect 14101 1332 14113 1366
rect 14055 1298 14113 1332
rect 14055 1264 14067 1298
rect 14101 1264 14113 1298
rect 14055 1230 14113 1264
rect 14055 1196 14067 1230
rect 14101 1196 14113 1230
rect 14055 1162 14113 1196
rect 14055 1128 14067 1162
rect 14101 1128 14113 1162
rect 14055 1004 14113 1128
rect 14143 1366 14201 1404
rect 14143 1332 14155 1366
rect 14189 1332 14201 1366
rect 14143 1298 14201 1332
rect 14143 1264 14155 1298
rect 14189 1264 14201 1298
rect 14143 1230 14201 1264
rect 14143 1196 14155 1230
rect 14189 1196 14201 1230
rect 14143 1162 14201 1196
rect 14143 1128 14155 1162
rect 14189 1128 14201 1162
rect 14143 1093 14201 1128
rect 14143 1059 14155 1093
rect 14189 1059 14201 1093
rect 14143 1004 14201 1059
rect 14231 1366 14289 1404
rect 14231 1332 14243 1366
rect 14277 1332 14289 1366
rect 14231 1298 14289 1332
rect 14231 1264 14243 1298
rect 14277 1264 14289 1298
rect 14231 1230 14289 1264
rect 14231 1196 14243 1230
rect 14277 1196 14289 1230
rect 14231 1162 14289 1196
rect 14231 1128 14243 1162
rect 14277 1128 14289 1162
rect 14231 1004 14289 1128
rect 14319 1366 14377 1404
rect 14319 1332 14331 1366
rect 14365 1332 14377 1366
rect 14319 1298 14377 1332
rect 14319 1264 14331 1298
rect 14365 1264 14377 1298
rect 14319 1230 14377 1264
rect 14319 1196 14331 1230
rect 14365 1196 14377 1230
rect 14319 1162 14377 1196
rect 14319 1128 14331 1162
rect 14365 1128 14377 1162
rect 14319 1093 14377 1128
rect 14319 1059 14331 1093
rect 14365 1059 14377 1093
rect 14319 1004 14377 1059
rect 14407 1366 14461 1404
rect 14407 1332 14419 1366
rect 14453 1332 14461 1366
rect 14407 1298 14461 1332
rect 14407 1264 14419 1298
rect 14453 1264 14461 1298
rect 14407 1230 14461 1264
rect 14407 1196 14419 1230
rect 14453 1196 14461 1230
rect 14407 1162 14461 1196
rect 14407 1128 14419 1162
rect 14453 1128 14461 1162
rect 14407 1004 14461 1128
rect 14783 1365 14839 1405
rect 14783 1331 14793 1365
rect 14827 1331 14839 1365
rect 14783 1297 14839 1331
rect 14783 1263 14793 1297
rect 14827 1263 14839 1297
rect 14783 1229 14839 1263
rect 14783 1195 14793 1229
rect 14827 1195 14839 1229
rect 14783 1161 14839 1195
rect 14783 1127 14793 1161
rect 14827 1127 14839 1161
rect 14783 1093 14839 1127
rect 14783 1059 14793 1093
rect 14827 1059 14839 1093
rect 14783 1005 14839 1059
rect 14869 1365 14927 1405
rect 14869 1331 14881 1365
rect 14915 1331 14927 1365
rect 14869 1297 14927 1331
rect 14869 1263 14881 1297
rect 14915 1263 14927 1297
rect 14869 1229 14927 1263
rect 14869 1195 14881 1229
rect 14915 1195 14927 1229
rect 14869 1161 14927 1195
rect 14869 1127 14881 1161
rect 14915 1127 14927 1161
rect 14869 1093 14927 1127
rect 14869 1059 14881 1093
rect 14915 1059 14927 1093
rect 14869 1005 14927 1059
rect 14957 1365 15015 1405
rect 14957 1331 14969 1365
rect 15003 1331 15015 1365
rect 14957 1297 15015 1331
rect 14957 1263 14969 1297
rect 15003 1263 15015 1297
rect 14957 1229 15015 1263
rect 14957 1195 14969 1229
rect 15003 1195 15015 1229
rect 14957 1161 15015 1195
rect 14957 1127 14969 1161
rect 15003 1127 15015 1161
rect 14957 1005 15015 1127
rect 15045 1365 15103 1405
rect 15045 1331 15057 1365
rect 15091 1331 15103 1365
rect 15045 1297 15103 1331
rect 15045 1263 15057 1297
rect 15091 1263 15103 1297
rect 15045 1229 15103 1263
rect 15045 1195 15057 1229
rect 15091 1195 15103 1229
rect 15045 1161 15103 1195
rect 15045 1127 15057 1161
rect 15091 1127 15103 1161
rect 15045 1005 15103 1127
rect 15133 1365 15187 1405
rect 15133 1331 15145 1365
rect 15179 1331 15187 1365
rect 15133 1297 15187 1331
rect 15133 1263 15145 1297
rect 15179 1263 15187 1297
rect 15133 1229 15187 1263
rect 15133 1195 15145 1229
rect 15179 1195 15187 1229
rect 15133 1161 15187 1195
rect 15133 1127 15145 1161
rect 15179 1127 15187 1161
rect 15133 1093 15187 1127
rect 15133 1059 15145 1093
rect 15179 1059 15187 1093
rect 15133 1005 15187 1059
rect 15449 1365 15503 1405
rect 15449 1331 15457 1365
rect 15491 1331 15503 1365
rect 15449 1297 15503 1331
rect 15449 1263 15457 1297
rect 15491 1263 15503 1297
rect 15449 1229 15503 1263
rect 15449 1195 15457 1229
rect 15491 1195 15503 1229
rect 15449 1161 15503 1195
rect 15449 1127 15457 1161
rect 15491 1127 15503 1161
rect 15449 1005 15503 1127
rect 15533 1297 15591 1405
rect 15533 1263 15545 1297
rect 15579 1263 15591 1297
rect 15533 1229 15591 1263
rect 15533 1195 15545 1229
rect 15579 1195 15591 1229
rect 15533 1161 15591 1195
rect 15533 1127 15545 1161
rect 15579 1127 15591 1161
rect 15533 1093 15591 1127
rect 15533 1059 15545 1093
rect 15579 1059 15591 1093
rect 15533 1005 15591 1059
rect 15621 1365 15679 1405
rect 15621 1331 15633 1365
rect 15667 1331 15679 1365
rect 15621 1297 15679 1331
rect 15621 1263 15633 1297
rect 15667 1263 15679 1297
rect 15621 1229 15679 1263
rect 15621 1195 15633 1229
rect 15667 1195 15679 1229
rect 15621 1161 15679 1195
rect 15621 1127 15633 1161
rect 15667 1127 15679 1161
rect 15621 1005 15679 1127
rect 15709 1297 15767 1405
rect 15709 1263 15721 1297
rect 15755 1263 15767 1297
rect 15709 1229 15767 1263
rect 15709 1195 15721 1229
rect 15755 1195 15767 1229
rect 15709 1161 15767 1195
rect 15709 1127 15721 1161
rect 15755 1127 15767 1161
rect 15709 1005 15767 1127
rect 15797 1365 15853 1405
rect 15797 1331 15809 1365
rect 15843 1331 15853 1365
rect 15797 1297 15853 1331
rect 15797 1263 15809 1297
rect 15843 1263 15853 1297
rect 15797 1229 15853 1263
rect 15797 1195 15809 1229
rect 15843 1195 15853 1229
rect 15797 1161 15853 1195
rect 15797 1127 15809 1161
rect 15843 1127 15853 1161
rect 15797 1005 15853 1127
rect 16115 1365 16171 1405
rect 16115 1331 16125 1365
rect 16159 1331 16171 1365
rect 16115 1297 16171 1331
rect 16115 1263 16125 1297
rect 16159 1263 16171 1297
rect 16115 1229 16171 1263
rect 16115 1195 16125 1229
rect 16159 1195 16171 1229
rect 16115 1161 16171 1195
rect 16115 1127 16125 1161
rect 16159 1127 16171 1161
rect 16115 1005 16171 1127
rect 16201 1297 16259 1405
rect 16201 1263 16213 1297
rect 16247 1263 16259 1297
rect 16201 1229 16259 1263
rect 16201 1195 16213 1229
rect 16247 1195 16259 1229
rect 16201 1161 16259 1195
rect 16201 1127 16213 1161
rect 16247 1127 16259 1161
rect 16201 1093 16259 1127
rect 16201 1059 16213 1093
rect 16247 1059 16259 1093
rect 16201 1005 16259 1059
rect 16289 1365 16347 1405
rect 16289 1331 16301 1365
rect 16335 1331 16347 1365
rect 16289 1297 16347 1331
rect 16289 1263 16301 1297
rect 16335 1263 16347 1297
rect 16289 1229 16347 1263
rect 16289 1195 16301 1229
rect 16335 1195 16347 1229
rect 16289 1161 16347 1195
rect 16289 1127 16301 1161
rect 16335 1127 16347 1161
rect 16289 1005 16347 1127
rect 16377 1297 16435 1405
rect 16377 1263 16389 1297
rect 16423 1263 16435 1297
rect 16377 1229 16435 1263
rect 16377 1195 16389 1229
rect 16423 1195 16435 1229
rect 16377 1161 16435 1195
rect 16377 1127 16389 1161
rect 16423 1127 16435 1161
rect 16377 1093 16435 1127
rect 16377 1059 16389 1093
rect 16423 1059 16435 1093
rect 16377 1005 16435 1059
rect 16465 1365 16519 1405
rect 16465 1331 16477 1365
rect 16511 1331 16519 1365
rect 16465 1297 16519 1331
rect 16465 1263 16477 1297
rect 16511 1263 16519 1297
rect 16465 1229 16519 1263
rect 16465 1195 16477 1229
rect 16511 1195 16519 1229
rect 16465 1161 16519 1195
rect 16465 1127 16477 1161
rect 16511 1127 16519 1161
rect 16465 1005 16519 1127
rect 16758 1366 16814 1404
rect 16758 1332 16768 1366
rect 16802 1332 16814 1366
rect 16758 1298 16814 1332
rect 16758 1264 16768 1298
rect 16802 1264 16814 1298
rect 16758 1230 16814 1264
rect 16758 1196 16768 1230
rect 16802 1196 16814 1230
rect 16758 1162 16814 1196
rect 16758 1128 16768 1162
rect 16802 1128 16814 1162
rect 16758 1093 16814 1128
rect 16758 1059 16768 1093
rect 16802 1059 16814 1093
rect 16758 1004 16814 1059
rect 16844 1366 16902 1404
rect 16844 1332 16856 1366
rect 16890 1332 16902 1366
rect 16844 1298 16902 1332
rect 16844 1264 16856 1298
rect 16890 1264 16902 1298
rect 16844 1230 16902 1264
rect 16844 1196 16856 1230
rect 16890 1196 16902 1230
rect 16844 1162 16902 1196
rect 16844 1128 16856 1162
rect 16890 1128 16902 1162
rect 16844 1093 16902 1128
rect 16844 1059 16856 1093
rect 16890 1059 16902 1093
rect 16844 1004 16902 1059
rect 16932 1366 16986 1404
rect 16932 1332 16944 1366
rect 16978 1332 16986 1366
rect 16932 1298 16986 1332
rect 16932 1264 16944 1298
rect 16978 1264 16986 1298
rect 16932 1230 16986 1264
rect 16932 1196 16944 1230
rect 16978 1196 16986 1230
rect 16932 1162 16986 1196
rect 16932 1128 16944 1162
rect 16978 1128 16986 1162
rect 16932 1093 16986 1128
rect 16932 1059 16944 1093
rect 16978 1059 16986 1093
rect 16932 1004 16986 1059
<< ndiffc >>
rect 122 299 156 333
rect 219 299 253 333
rect 316 299 350 333
rect 122 227 156 261
rect 122 159 156 193
rect 219 174 253 208
rect 316 227 350 261
rect 316 159 350 193
rect 413 183 447 217
rect 510 227 544 261
rect 510 159 544 193
rect 122 89 156 123
rect 316 89 350 123
rect 413 89 447 123
rect 510 89 544 123
rect 767 301 801 335
rect 864 301 898 335
rect 961 301 995 335
rect 1058 301 1092 335
rect 1155 301 1189 335
rect 767 229 801 263
rect 767 161 801 195
rect 864 176 898 210
rect 961 229 995 263
rect 961 161 995 195
rect 1059 182 1093 216
rect 767 91 801 125
rect 961 91 995 125
rect 1058 91 1092 125
rect 1155 91 1189 125
rect 1269 301 1303 335
rect 1269 229 1303 263
rect 1269 161 1303 195
rect 1366 185 1400 219
rect 1463 229 1497 263
rect 1463 161 1497 195
rect 1269 91 1303 125
rect 1366 91 1400 125
rect 1463 91 1497 125
rect 1729 301 1763 335
rect 1826 301 1860 335
rect 1923 301 1957 335
rect 2020 301 2054 335
rect 2117 301 2151 335
rect 1729 229 1763 263
rect 1729 161 1763 195
rect 1826 176 1860 210
rect 1923 229 1957 263
rect 1923 161 1957 195
rect 2021 182 2055 216
rect 1729 91 1763 125
rect 1923 91 1957 125
rect 2020 91 2054 125
rect 2117 91 2151 125
rect 2231 301 2265 335
rect 2231 229 2265 263
rect 2231 161 2265 195
rect 2328 185 2362 219
rect 2425 229 2459 263
rect 2425 161 2459 195
rect 2231 91 2265 125
rect 2328 91 2362 125
rect 2425 91 2459 125
rect 2712 299 2746 333
rect 2809 299 2843 333
rect 2906 299 2940 333
rect 2712 227 2746 261
rect 2712 159 2746 193
rect 2809 174 2843 208
rect 2906 227 2940 261
rect 2906 159 2940 193
rect 3003 183 3037 217
rect 3100 227 3134 261
rect 3100 159 3134 193
rect 2712 89 2746 123
rect 2906 89 2940 123
rect 3003 89 3037 123
rect 3100 89 3134 123
rect 3378 299 3412 333
rect 3475 299 3509 333
rect 3572 299 3606 333
rect 3378 227 3412 261
rect 3378 159 3412 193
rect 3475 174 3509 208
rect 3572 227 3606 261
rect 3572 159 3606 193
rect 3669 183 3703 217
rect 3766 227 3800 261
rect 3766 159 3800 193
rect 3378 89 3412 123
rect 3572 89 3606 123
rect 3669 89 3703 123
rect 3766 89 3800 123
rect 4023 301 4057 335
rect 4120 301 4154 335
rect 4217 301 4251 335
rect 4314 301 4348 335
rect 4411 301 4445 335
rect 4023 229 4057 263
rect 4023 161 4057 195
rect 4120 176 4154 210
rect 4217 229 4251 263
rect 4217 161 4251 195
rect 4315 182 4349 216
rect 4023 91 4057 125
rect 4217 91 4251 125
rect 4314 91 4348 125
rect 4411 91 4445 125
rect 4525 301 4559 335
rect 4525 229 4559 263
rect 4525 161 4559 195
rect 4622 185 4656 219
rect 4719 229 4753 263
rect 4719 161 4753 195
rect 4525 91 4559 125
rect 4622 91 4656 125
rect 4719 91 4753 125
rect 5006 299 5040 333
rect 5103 299 5137 333
rect 5200 299 5234 333
rect 5006 227 5040 261
rect 5006 159 5040 193
rect 5103 174 5137 208
rect 5200 227 5234 261
rect 5200 159 5234 193
rect 5297 183 5331 217
rect 5394 227 5428 261
rect 5394 159 5428 193
rect 5006 89 5040 123
rect 5200 89 5234 123
rect 5297 89 5331 123
rect 5394 89 5428 123
rect 5651 301 5685 335
rect 5748 301 5782 335
rect 5845 301 5879 335
rect 5942 301 5976 335
rect 6039 301 6073 335
rect 5651 229 5685 263
rect 5651 161 5685 195
rect 5748 176 5782 210
rect 5845 229 5879 263
rect 5845 161 5879 195
rect 5943 182 5977 216
rect 5651 91 5685 125
rect 5845 91 5879 125
rect 5942 91 5976 125
rect 6039 91 6073 125
rect 6153 301 6187 335
rect 6153 229 6187 263
rect 6153 161 6187 195
rect 6250 185 6284 219
rect 6347 229 6381 263
rect 6347 161 6381 195
rect 6153 91 6187 125
rect 6250 91 6284 125
rect 6347 91 6381 125
rect 6613 301 6647 335
rect 6710 301 6744 335
rect 6807 301 6841 335
rect 6904 301 6938 335
rect 7001 301 7035 335
rect 6613 229 6647 263
rect 6613 161 6647 195
rect 6710 176 6744 210
rect 6807 229 6841 263
rect 6807 161 6841 195
rect 6905 182 6939 216
rect 6613 91 6647 125
rect 6807 91 6841 125
rect 6904 91 6938 125
rect 7001 91 7035 125
rect 7115 301 7149 335
rect 7115 229 7149 263
rect 7115 161 7149 195
rect 7212 185 7246 219
rect 7309 229 7343 263
rect 7309 161 7343 195
rect 7115 91 7149 125
rect 7212 91 7246 125
rect 7309 91 7343 125
rect 7596 299 7630 333
rect 7693 299 7727 333
rect 7790 299 7824 333
rect 7596 227 7630 261
rect 7596 159 7630 193
rect 7693 174 7727 208
rect 7790 227 7824 261
rect 7790 159 7824 193
rect 7887 183 7921 217
rect 7984 227 8018 261
rect 7984 159 8018 193
rect 7596 89 7630 123
rect 7790 89 7824 123
rect 7887 89 7921 123
rect 7984 89 8018 123
rect 8262 299 8296 333
rect 8359 299 8393 333
rect 8456 299 8490 333
rect 8262 227 8296 261
rect 8262 159 8296 193
rect 8359 174 8393 208
rect 8456 227 8490 261
rect 8456 159 8490 193
rect 8553 183 8587 217
rect 8650 227 8684 261
rect 8650 159 8684 193
rect 8262 89 8296 123
rect 8456 89 8490 123
rect 8553 89 8587 123
rect 8650 89 8684 123
rect 8907 301 8941 335
rect 9004 301 9038 335
rect 9101 301 9135 335
rect 9198 301 9232 335
rect 9295 301 9329 335
rect 8907 229 8941 263
rect 8907 161 8941 195
rect 9004 176 9038 210
rect 9101 229 9135 263
rect 9101 161 9135 195
rect 9199 182 9233 216
rect 8907 91 8941 125
rect 9101 91 9135 125
rect 9198 91 9232 125
rect 9295 91 9329 125
rect 9409 301 9443 335
rect 9409 229 9443 263
rect 9409 161 9443 195
rect 9506 185 9540 219
rect 9603 229 9637 263
rect 9603 161 9637 195
rect 9409 91 9443 125
rect 9506 91 9540 125
rect 9603 91 9637 125
rect 9890 299 9924 333
rect 9987 299 10021 333
rect 10084 299 10118 333
rect 9890 227 9924 261
rect 9890 159 9924 193
rect 9987 174 10021 208
rect 10084 227 10118 261
rect 10084 159 10118 193
rect 10181 183 10215 217
rect 10278 227 10312 261
rect 10278 159 10312 193
rect 9890 89 9924 123
rect 10084 89 10118 123
rect 10181 89 10215 123
rect 10278 89 10312 123
rect 10535 301 10569 335
rect 10632 301 10666 335
rect 10729 301 10763 335
rect 10826 301 10860 335
rect 10923 301 10957 335
rect 10535 229 10569 263
rect 10535 161 10569 195
rect 10632 176 10666 210
rect 10729 229 10763 263
rect 10729 161 10763 195
rect 10827 182 10861 216
rect 10535 91 10569 125
rect 10729 91 10763 125
rect 10826 91 10860 125
rect 10923 91 10957 125
rect 11037 301 11071 335
rect 11037 229 11071 263
rect 11037 161 11071 195
rect 11134 185 11168 219
rect 11231 229 11265 263
rect 11231 161 11265 195
rect 11037 91 11071 125
rect 11134 91 11168 125
rect 11231 91 11265 125
rect 11497 301 11531 335
rect 11594 301 11628 335
rect 11691 301 11725 335
rect 11788 301 11822 335
rect 11885 301 11919 335
rect 11497 229 11531 263
rect 11497 161 11531 195
rect 11594 176 11628 210
rect 11691 229 11725 263
rect 11691 161 11725 195
rect 11789 182 11823 216
rect 11497 91 11531 125
rect 11691 91 11725 125
rect 11788 91 11822 125
rect 11885 91 11919 125
rect 11999 301 12033 335
rect 11999 229 12033 263
rect 11999 161 12033 195
rect 12096 185 12130 219
rect 12193 229 12227 263
rect 12193 161 12227 195
rect 11999 91 12033 125
rect 12096 91 12130 125
rect 12193 91 12227 125
rect 12480 299 12514 333
rect 12577 299 12611 333
rect 12674 299 12708 333
rect 12480 227 12514 261
rect 12480 159 12514 193
rect 12577 174 12611 208
rect 12674 227 12708 261
rect 12674 159 12708 193
rect 12771 183 12805 217
rect 12868 227 12902 261
rect 12868 159 12902 193
rect 12480 89 12514 123
rect 12674 89 12708 123
rect 12771 89 12805 123
rect 12868 89 12902 123
rect 13146 299 13180 333
rect 13243 299 13277 333
rect 13340 299 13374 333
rect 13146 227 13180 261
rect 13146 159 13180 193
rect 13243 174 13277 208
rect 13340 227 13374 261
rect 13340 159 13374 193
rect 13437 183 13471 217
rect 13534 227 13568 261
rect 13534 159 13568 193
rect 13146 89 13180 123
rect 13340 89 13374 123
rect 13437 89 13471 123
rect 13534 89 13568 123
rect 13791 301 13825 335
rect 13888 301 13922 335
rect 13985 301 14019 335
rect 14082 301 14116 335
rect 14179 301 14213 335
rect 13791 229 13825 263
rect 13791 161 13825 195
rect 13888 176 13922 210
rect 13985 229 14019 263
rect 13985 161 14019 195
rect 14083 182 14117 216
rect 13791 91 13825 125
rect 13985 91 14019 125
rect 14082 91 14116 125
rect 14179 91 14213 125
rect 14293 301 14327 335
rect 14293 229 14327 263
rect 14293 161 14327 195
rect 14390 185 14424 219
rect 14487 229 14521 263
rect 14487 161 14521 195
rect 14293 91 14327 125
rect 14390 91 14424 125
rect 14487 91 14521 125
rect 14774 299 14808 333
rect 14871 299 14905 333
rect 14968 299 15002 333
rect 15162 299 15196 333
rect 14774 227 14808 261
rect 14774 159 14808 193
rect 14871 174 14905 208
rect 14968 227 15002 261
rect 14968 159 15002 193
rect 15064 183 15098 217
rect 15162 227 15196 261
rect 15162 159 15196 193
rect 14774 89 14808 123
rect 14968 89 15002 123
rect 15064 89 15098 123
rect 15162 89 15196 123
rect 15440 299 15474 333
rect 15537 299 15571 333
rect 15634 299 15668 333
rect 15828 299 15862 333
rect 15440 227 15474 261
rect 15440 159 15474 193
rect 15537 174 15571 208
rect 15634 227 15668 261
rect 15634 159 15668 193
rect 15731 183 15765 217
rect 15828 227 15862 261
rect 15828 159 15862 193
rect 15440 89 15474 123
rect 15634 89 15668 123
rect 15731 89 15765 123
rect 15828 89 15862 123
rect 16106 299 16140 333
rect 16203 299 16237 333
rect 16300 299 16334 333
rect 16106 227 16140 261
rect 16106 159 16140 193
rect 16203 174 16237 208
rect 16300 227 16334 261
rect 16300 159 16334 193
rect 16397 183 16431 217
rect 16494 227 16528 261
rect 16494 159 16528 193
rect 16106 89 16140 123
rect 16300 89 16334 123
rect 16397 89 16431 123
rect 16494 89 16528 123
rect 16759 300 16793 334
rect 16953 300 16987 334
rect 16759 228 16793 262
rect 16759 160 16793 194
rect 16855 184 16889 218
rect 16953 228 16987 262
rect 16953 160 16987 194
rect 16759 90 16793 124
rect 16855 90 16889 124
rect 16953 90 16987 124
<< pdiffc >>
rect 141 1332 175 1366
rect 141 1264 175 1298
rect 141 1196 175 1230
rect 141 1128 175 1162
rect 141 1059 175 1093
rect 229 1332 263 1366
rect 229 1264 263 1298
rect 229 1196 263 1230
rect 229 1128 263 1162
rect 229 1059 263 1093
rect 317 1332 351 1366
rect 317 1264 351 1298
rect 317 1196 351 1230
rect 317 1128 351 1162
rect 405 1332 439 1366
rect 405 1264 439 1298
rect 405 1196 439 1230
rect 405 1128 439 1162
rect 405 1059 439 1093
rect 493 1332 527 1366
rect 493 1264 527 1298
rect 493 1196 527 1230
rect 493 1128 527 1162
rect 867 1332 901 1366
rect 867 1264 901 1298
rect 867 1196 901 1230
rect 867 1128 901 1162
rect 867 1059 901 1093
rect 955 1332 989 1366
rect 955 1264 989 1298
rect 955 1196 989 1230
rect 955 1128 989 1162
rect 955 1059 989 1093
rect 1043 1332 1077 1366
rect 1043 1264 1077 1298
rect 1043 1196 1077 1230
rect 1043 1128 1077 1162
rect 1131 1332 1165 1366
rect 1131 1264 1165 1298
rect 1131 1196 1165 1230
rect 1131 1128 1165 1162
rect 1131 1059 1165 1093
rect 1219 1332 1253 1366
rect 1219 1264 1253 1298
rect 1219 1196 1253 1230
rect 1219 1128 1253 1162
rect 1307 1332 1341 1366
rect 1307 1264 1341 1298
rect 1307 1196 1341 1230
rect 1307 1128 1341 1162
rect 1307 1059 1341 1093
rect 1395 1332 1429 1366
rect 1395 1264 1429 1298
rect 1395 1196 1429 1230
rect 1395 1128 1429 1162
rect 1829 1332 1863 1366
rect 1829 1264 1863 1298
rect 1829 1196 1863 1230
rect 1829 1128 1863 1162
rect 1829 1059 1863 1093
rect 1917 1332 1951 1366
rect 1917 1264 1951 1298
rect 1917 1196 1951 1230
rect 1917 1128 1951 1162
rect 1917 1059 1951 1093
rect 2005 1332 2039 1366
rect 2005 1264 2039 1298
rect 2005 1196 2039 1230
rect 2005 1128 2039 1162
rect 2093 1332 2127 1366
rect 2093 1264 2127 1298
rect 2093 1196 2127 1230
rect 2093 1128 2127 1162
rect 2093 1059 2127 1093
rect 2181 1332 2215 1366
rect 2181 1264 2215 1298
rect 2181 1196 2215 1230
rect 2181 1128 2215 1162
rect 2269 1332 2303 1366
rect 2269 1264 2303 1298
rect 2269 1196 2303 1230
rect 2269 1128 2303 1162
rect 2269 1059 2303 1093
rect 2357 1332 2391 1366
rect 2357 1264 2391 1298
rect 2357 1196 2391 1230
rect 2357 1128 2391 1162
rect 2731 1332 2765 1366
rect 2731 1264 2765 1298
rect 2731 1196 2765 1230
rect 2731 1128 2765 1162
rect 2731 1059 2765 1093
rect 2819 1332 2853 1366
rect 2819 1264 2853 1298
rect 2819 1196 2853 1230
rect 2819 1128 2853 1162
rect 2819 1059 2853 1093
rect 2907 1332 2941 1366
rect 2907 1264 2941 1298
rect 2907 1196 2941 1230
rect 2907 1128 2941 1162
rect 2995 1332 3029 1366
rect 2995 1264 3029 1298
rect 2995 1196 3029 1230
rect 2995 1128 3029 1162
rect 2995 1059 3029 1093
rect 3083 1332 3117 1366
rect 3083 1264 3117 1298
rect 3083 1196 3117 1230
rect 3083 1128 3117 1162
rect 3397 1332 3431 1366
rect 3397 1264 3431 1298
rect 3397 1196 3431 1230
rect 3397 1128 3431 1162
rect 3397 1059 3431 1093
rect 3485 1332 3519 1366
rect 3485 1264 3519 1298
rect 3485 1196 3519 1230
rect 3485 1128 3519 1162
rect 3485 1059 3519 1093
rect 3573 1332 3607 1366
rect 3573 1264 3607 1298
rect 3573 1196 3607 1230
rect 3573 1128 3607 1162
rect 3661 1332 3695 1366
rect 3661 1264 3695 1298
rect 3661 1196 3695 1230
rect 3661 1128 3695 1162
rect 3661 1059 3695 1093
rect 3749 1332 3783 1366
rect 3749 1264 3783 1298
rect 3749 1196 3783 1230
rect 3749 1128 3783 1162
rect 4123 1332 4157 1366
rect 4123 1264 4157 1298
rect 4123 1196 4157 1230
rect 4123 1128 4157 1162
rect 4123 1059 4157 1093
rect 4211 1332 4245 1366
rect 4211 1264 4245 1298
rect 4211 1196 4245 1230
rect 4211 1128 4245 1162
rect 4211 1059 4245 1093
rect 4299 1332 4333 1366
rect 4299 1264 4333 1298
rect 4299 1196 4333 1230
rect 4299 1128 4333 1162
rect 4387 1332 4421 1366
rect 4387 1264 4421 1298
rect 4387 1196 4421 1230
rect 4387 1128 4421 1162
rect 4387 1059 4421 1093
rect 4475 1332 4509 1366
rect 4475 1264 4509 1298
rect 4475 1196 4509 1230
rect 4475 1128 4509 1162
rect 4563 1332 4597 1366
rect 4563 1264 4597 1298
rect 4563 1196 4597 1230
rect 4563 1128 4597 1162
rect 4563 1059 4597 1093
rect 4651 1332 4685 1366
rect 4651 1264 4685 1298
rect 4651 1196 4685 1230
rect 4651 1128 4685 1162
rect 5025 1332 5059 1366
rect 5025 1264 5059 1298
rect 5025 1196 5059 1230
rect 5025 1128 5059 1162
rect 5025 1059 5059 1093
rect 5113 1332 5147 1366
rect 5113 1264 5147 1298
rect 5113 1196 5147 1230
rect 5113 1128 5147 1162
rect 5113 1059 5147 1093
rect 5201 1332 5235 1366
rect 5201 1264 5235 1298
rect 5201 1196 5235 1230
rect 5201 1128 5235 1162
rect 5289 1332 5323 1366
rect 5289 1264 5323 1298
rect 5289 1196 5323 1230
rect 5289 1128 5323 1162
rect 5289 1059 5323 1093
rect 5377 1332 5411 1366
rect 5377 1264 5411 1298
rect 5377 1196 5411 1230
rect 5377 1128 5411 1162
rect 5751 1332 5785 1366
rect 5751 1264 5785 1298
rect 5751 1196 5785 1230
rect 5751 1128 5785 1162
rect 5751 1059 5785 1093
rect 5839 1332 5873 1366
rect 5839 1264 5873 1298
rect 5839 1196 5873 1230
rect 5839 1128 5873 1162
rect 5839 1059 5873 1093
rect 5927 1332 5961 1366
rect 5927 1264 5961 1298
rect 5927 1196 5961 1230
rect 5927 1128 5961 1162
rect 6015 1332 6049 1366
rect 6015 1264 6049 1298
rect 6015 1196 6049 1230
rect 6015 1128 6049 1162
rect 6015 1059 6049 1093
rect 6103 1332 6137 1366
rect 6103 1264 6137 1298
rect 6103 1196 6137 1230
rect 6103 1128 6137 1162
rect 6191 1332 6225 1366
rect 6191 1264 6225 1298
rect 6191 1196 6225 1230
rect 6191 1128 6225 1162
rect 6191 1059 6225 1093
rect 6279 1332 6313 1366
rect 6279 1264 6313 1298
rect 6279 1196 6313 1230
rect 6279 1128 6313 1162
rect 6713 1332 6747 1366
rect 6713 1264 6747 1298
rect 6713 1196 6747 1230
rect 6713 1128 6747 1162
rect 6713 1059 6747 1093
rect 6801 1332 6835 1366
rect 6801 1264 6835 1298
rect 6801 1196 6835 1230
rect 6801 1128 6835 1162
rect 6801 1059 6835 1093
rect 6889 1332 6923 1366
rect 6889 1264 6923 1298
rect 6889 1196 6923 1230
rect 6889 1128 6923 1162
rect 6977 1332 7011 1366
rect 6977 1264 7011 1298
rect 6977 1196 7011 1230
rect 6977 1128 7011 1162
rect 6977 1059 7011 1093
rect 7065 1332 7099 1366
rect 7065 1264 7099 1298
rect 7065 1196 7099 1230
rect 7065 1128 7099 1162
rect 7153 1332 7187 1366
rect 7153 1264 7187 1298
rect 7153 1196 7187 1230
rect 7153 1128 7187 1162
rect 7153 1059 7187 1093
rect 7241 1332 7275 1366
rect 7241 1264 7275 1298
rect 7241 1196 7275 1230
rect 7241 1128 7275 1162
rect 7615 1332 7649 1366
rect 7615 1264 7649 1298
rect 7615 1196 7649 1230
rect 7615 1128 7649 1162
rect 7615 1059 7649 1093
rect 7703 1332 7737 1366
rect 7703 1264 7737 1298
rect 7703 1196 7737 1230
rect 7703 1128 7737 1162
rect 7703 1059 7737 1093
rect 7791 1332 7825 1366
rect 7791 1264 7825 1298
rect 7791 1196 7825 1230
rect 7791 1128 7825 1162
rect 7879 1332 7913 1366
rect 7879 1264 7913 1298
rect 7879 1196 7913 1230
rect 7879 1128 7913 1162
rect 7879 1059 7913 1093
rect 7967 1332 8001 1366
rect 7967 1264 8001 1298
rect 7967 1196 8001 1230
rect 7967 1128 8001 1162
rect 8281 1332 8315 1366
rect 8281 1264 8315 1298
rect 8281 1196 8315 1230
rect 8281 1128 8315 1162
rect 8281 1059 8315 1093
rect 8369 1332 8403 1366
rect 8369 1264 8403 1298
rect 8369 1196 8403 1230
rect 8369 1128 8403 1162
rect 8369 1059 8403 1093
rect 8457 1332 8491 1366
rect 8457 1264 8491 1298
rect 8457 1196 8491 1230
rect 8457 1128 8491 1162
rect 8545 1332 8579 1366
rect 8545 1264 8579 1298
rect 8545 1196 8579 1230
rect 8545 1128 8579 1162
rect 8545 1059 8579 1093
rect 8633 1332 8667 1366
rect 8633 1264 8667 1298
rect 8633 1196 8667 1230
rect 8633 1128 8667 1162
rect 9007 1332 9041 1366
rect 9007 1264 9041 1298
rect 9007 1196 9041 1230
rect 9007 1128 9041 1162
rect 9007 1059 9041 1093
rect 9095 1332 9129 1366
rect 9095 1264 9129 1298
rect 9095 1196 9129 1230
rect 9095 1128 9129 1162
rect 9095 1059 9129 1093
rect 9183 1332 9217 1366
rect 9183 1264 9217 1298
rect 9183 1196 9217 1230
rect 9183 1128 9217 1162
rect 9271 1332 9305 1366
rect 9271 1264 9305 1298
rect 9271 1196 9305 1230
rect 9271 1128 9305 1162
rect 9271 1059 9305 1093
rect 9359 1332 9393 1366
rect 9359 1264 9393 1298
rect 9359 1196 9393 1230
rect 9359 1128 9393 1162
rect 9447 1332 9481 1366
rect 9447 1264 9481 1298
rect 9447 1196 9481 1230
rect 9447 1128 9481 1162
rect 9447 1059 9481 1093
rect 9535 1332 9569 1366
rect 9535 1264 9569 1298
rect 9535 1196 9569 1230
rect 9535 1128 9569 1162
rect 9909 1332 9943 1366
rect 9909 1264 9943 1298
rect 9909 1196 9943 1230
rect 9909 1128 9943 1162
rect 9909 1059 9943 1093
rect 9997 1332 10031 1366
rect 9997 1264 10031 1298
rect 9997 1196 10031 1230
rect 9997 1128 10031 1162
rect 9997 1059 10031 1093
rect 10085 1332 10119 1366
rect 10085 1264 10119 1298
rect 10085 1196 10119 1230
rect 10085 1128 10119 1162
rect 10173 1332 10207 1366
rect 10173 1264 10207 1298
rect 10173 1196 10207 1230
rect 10173 1128 10207 1162
rect 10173 1059 10207 1093
rect 10261 1332 10295 1366
rect 10261 1264 10295 1298
rect 10261 1196 10295 1230
rect 10261 1128 10295 1162
rect 10635 1332 10669 1366
rect 10635 1264 10669 1298
rect 10635 1196 10669 1230
rect 10635 1128 10669 1162
rect 10635 1059 10669 1093
rect 10723 1332 10757 1366
rect 10723 1264 10757 1298
rect 10723 1196 10757 1230
rect 10723 1128 10757 1162
rect 10723 1059 10757 1093
rect 10811 1332 10845 1366
rect 10811 1264 10845 1298
rect 10811 1196 10845 1230
rect 10811 1128 10845 1162
rect 10899 1332 10933 1366
rect 10899 1264 10933 1298
rect 10899 1196 10933 1230
rect 10899 1128 10933 1162
rect 10899 1059 10933 1093
rect 10987 1332 11021 1366
rect 10987 1264 11021 1298
rect 10987 1196 11021 1230
rect 10987 1128 11021 1162
rect 11075 1332 11109 1366
rect 11075 1264 11109 1298
rect 11075 1196 11109 1230
rect 11075 1128 11109 1162
rect 11075 1059 11109 1093
rect 11163 1332 11197 1366
rect 11163 1264 11197 1298
rect 11163 1196 11197 1230
rect 11163 1128 11197 1162
rect 11597 1332 11631 1366
rect 11597 1264 11631 1298
rect 11597 1196 11631 1230
rect 11597 1128 11631 1162
rect 11597 1059 11631 1093
rect 11685 1332 11719 1366
rect 11685 1264 11719 1298
rect 11685 1196 11719 1230
rect 11685 1128 11719 1162
rect 11685 1059 11719 1093
rect 11773 1332 11807 1366
rect 11773 1264 11807 1298
rect 11773 1196 11807 1230
rect 11773 1128 11807 1162
rect 11861 1332 11895 1366
rect 11861 1264 11895 1298
rect 11861 1196 11895 1230
rect 11861 1128 11895 1162
rect 11861 1059 11895 1093
rect 11949 1332 11983 1366
rect 11949 1264 11983 1298
rect 11949 1196 11983 1230
rect 11949 1128 11983 1162
rect 12037 1332 12071 1366
rect 12037 1264 12071 1298
rect 12037 1196 12071 1230
rect 12037 1128 12071 1162
rect 12037 1059 12071 1093
rect 12125 1332 12159 1366
rect 12125 1264 12159 1298
rect 12125 1196 12159 1230
rect 12125 1128 12159 1162
rect 12499 1332 12533 1366
rect 12499 1264 12533 1298
rect 12499 1196 12533 1230
rect 12499 1128 12533 1162
rect 12499 1059 12533 1093
rect 12587 1332 12621 1366
rect 12587 1264 12621 1298
rect 12587 1196 12621 1230
rect 12587 1128 12621 1162
rect 12587 1059 12621 1093
rect 12675 1332 12709 1366
rect 12675 1264 12709 1298
rect 12675 1196 12709 1230
rect 12675 1128 12709 1162
rect 12763 1332 12797 1366
rect 12763 1264 12797 1298
rect 12763 1196 12797 1230
rect 12763 1128 12797 1162
rect 12763 1059 12797 1093
rect 12851 1332 12885 1366
rect 12851 1264 12885 1298
rect 12851 1196 12885 1230
rect 12851 1128 12885 1162
rect 13165 1332 13199 1366
rect 13165 1264 13199 1298
rect 13165 1196 13199 1230
rect 13165 1128 13199 1162
rect 13165 1059 13199 1093
rect 13253 1332 13287 1366
rect 13253 1264 13287 1298
rect 13253 1196 13287 1230
rect 13253 1128 13287 1162
rect 13253 1059 13287 1093
rect 13341 1332 13375 1366
rect 13341 1264 13375 1298
rect 13341 1196 13375 1230
rect 13341 1128 13375 1162
rect 13429 1332 13463 1366
rect 13429 1264 13463 1298
rect 13429 1196 13463 1230
rect 13429 1128 13463 1162
rect 13429 1059 13463 1093
rect 13517 1332 13551 1366
rect 13517 1264 13551 1298
rect 13517 1196 13551 1230
rect 13517 1128 13551 1162
rect 13891 1332 13925 1366
rect 13891 1264 13925 1298
rect 13891 1196 13925 1230
rect 13891 1128 13925 1162
rect 13891 1059 13925 1093
rect 13979 1332 14013 1366
rect 13979 1264 14013 1298
rect 13979 1196 14013 1230
rect 13979 1128 14013 1162
rect 13979 1059 14013 1093
rect 14067 1332 14101 1366
rect 14067 1264 14101 1298
rect 14067 1196 14101 1230
rect 14067 1128 14101 1162
rect 14155 1332 14189 1366
rect 14155 1264 14189 1298
rect 14155 1196 14189 1230
rect 14155 1128 14189 1162
rect 14155 1059 14189 1093
rect 14243 1332 14277 1366
rect 14243 1264 14277 1298
rect 14243 1196 14277 1230
rect 14243 1128 14277 1162
rect 14331 1332 14365 1366
rect 14331 1264 14365 1298
rect 14331 1196 14365 1230
rect 14331 1128 14365 1162
rect 14331 1059 14365 1093
rect 14419 1332 14453 1366
rect 14419 1264 14453 1298
rect 14419 1196 14453 1230
rect 14419 1128 14453 1162
rect 14793 1331 14827 1365
rect 14793 1263 14827 1297
rect 14793 1195 14827 1229
rect 14793 1127 14827 1161
rect 14793 1059 14827 1093
rect 14881 1331 14915 1365
rect 14881 1263 14915 1297
rect 14881 1195 14915 1229
rect 14881 1127 14915 1161
rect 14881 1059 14915 1093
rect 14969 1331 15003 1365
rect 14969 1263 15003 1297
rect 14969 1195 15003 1229
rect 14969 1127 15003 1161
rect 15057 1331 15091 1365
rect 15057 1263 15091 1297
rect 15057 1195 15091 1229
rect 15057 1127 15091 1161
rect 15145 1331 15179 1365
rect 15145 1263 15179 1297
rect 15145 1195 15179 1229
rect 15145 1127 15179 1161
rect 15145 1059 15179 1093
rect 15457 1331 15491 1365
rect 15457 1263 15491 1297
rect 15457 1195 15491 1229
rect 15457 1127 15491 1161
rect 15545 1263 15579 1297
rect 15545 1195 15579 1229
rect 15545 1127 15579 1161
rect 15545 1059 15579 1093
rect 15633 1331 15667 1365
rect 15633 1263 15667 1297
rect 15633 1195 15667 1229
rect 15633 1127 15667 1161
rect 15721 1263 15755 1297
rect 15721 1195 15755 1229
rect 15721 1127 15755 1161
rect 15809 1331 15843 1365
rect 15809 1263 15843 1297
rect 15809 1195 15843 1229
rect 15809 1127 15843 1161
rect 16125 1331 16159 1365
rect 16125 1263 16159 1297
rect 16125 1195 16159 1229
rect 16125 1127 16159 1161
rect 16213 1263 16247 1297
rect 16213 1195 16247 1229
rect 16213 1127 16247 1161
rect 16213 1059 16247 1093
rect 16301 1331 16335 1365
rect 16301 1263 16335 1297
rect 16301 1195 16335 1229
rect 16301 1127 16335 1161
rect 16389 1263 16423 1297
rect 16389 1195 16423 1229
rect 16389 1127 16423 1161
rect 16389 1059 16423 1093
rect 16477 1331 16511 1365
rect 16477 1263 16511 1297
rect 16477 1195 16511 1229
rect 16477 1127 16511 1161
rect 16768 1332 16802 1366
rect 16768 1264 16802 1298
rect 16768 1196 16802 1230
rect 16768 1128 16802 1162
rect 16768 1059 16802 1093
rect 16856 1332 16890 1366
rect 16856 1264 16890 1298
rect 16856 1196 16890 1230
rect 16856 1128 16890 1162
rect 16856 1059 16890 1093
rect 16944 1332 16978 1366
rect 16944 1264 16978 1298
rect 16944 1196 16978 1230
rect 16944 1128 16978 1162
rect 16944 1059 16978 1093
<< psubdiff >>
rect -34 482 17128 544
rect -34 461 34 482
rect -34 427 -17 461
rect 17 427 34 461
rect 632 461 700 482
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect -34 313 34 353
rect 632 427 649 461
rect 683 427 700 461
rect 1594 461 1662 482
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 632 313 700 353
rect 1594 427 1611 461
rect 1645 427 1662 461
rect 2556 461 2624 482
rect 1594 387 1662 427
rect 1594 353 1611 387
rect 1645 353 1662 387
rect 632 279 649 313
rect 683 279 700 313
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect -34 17 34 57
rect 632 57 649 91
rect 683 57 700 91
rect 1594 313 1662 353
rect 2556 427 2573 461
rect 2607 427 2624 461
rect 3222 461 3290 482
rect 2556 387 2624 427
rect 2556 353 2573 387
rect 2607 353 2624 387
rect 1594 279 1611 313
rect 1645 279 1662 313
rect 1594 239 1662 279
rect 1594 205 1611 239
rect 1645 205 1662 239
rect 1594 165 1662 205
rect 1594 131 1611 165
rect 1645 131 1662 165
rect 1594 91 1662 131
rect 632 17 700 57
rect 1594 57 1611 91
rect 1645 57 1662 91
rect 2556 313 2624 353
rect 3222 427 3239 461
rect 3273 427 3290 461
rect 3888 461 3956 482
rect 3222 387 3290 427
rect 3222 353 3239 387
rect 3273 353 3290 387
rect 2556 279 2573 313
rect 2607 279 2624 313
rect 2556 239 2624 279
rect 2556 205 2573 239
rect 2607 205 2624 239
rect 2556 165 2624 205
rect 2556 131 2573 165
rect 2607 131 2624 165
rect 2556 91 2624 131
rect 1594 17 1662 57
rect 2556 57 2573 91
rect 2607 57 2624 91
rect 3222 313 3290 353
rect 3888 427 3905 461
rect 3939 427 3956 461
rect 4850 461 4918 482
rect 3888 387 3956 427
rect 3888 353 3905 387
rect 3939 353 3956 387
rect 3222 279 3239 313
rect 3273 279 3290 313
rect 3222 239 3290 279
rect 3222 205 3239 239
rect 3273 205 3290 239
rect 3222 165 3290 205
rect 3222 131 3239 165
rect 3273 131 3290 165
rect 3222 91 3290 131
rect 2556 17 2624 57
rect 3222 57 3239 91
rect 3273 57 3290 91
rect 3888 313 3956 353
rect 4850 427 4867 461
rect 4901 427 4918 461
rect 5516 461 5584 482
rect 4850 387 4918 427
rect 4850 353 4867 387
rect 4901 353 4918 387
rect 3888 279 3905 313
rect 3939 279 3956 313
rect 3888 239 3956 279
rect 3888 205 3905 239
rect 3939 205 3956 239
rect 3888 165 3956 205
rect 3888 131 3905 165
rect 3939 131 3956 165
rect 3888 91 3956 131
rect 3222 17 3290 57
rect 3888 57 3905 91
rect 3939 57 3956 91
rect 4850 313 4918 353
rect 5516 427 5533 461
rect 5567 427 5584 461
rect 6478 461 6546 482
rect 5516 387 5584 427
rect 5516 353 5533 387
rect 5567 353 5584 387
rect 4850 279 4867 313
rect 4901 279 4918 313
rect 4850 239 4918 279
rect 4850 205 4867 239
rect 4901 205 4918 239
rect 4850 165 4918 205
rect 4850 131 4867 165
rect 4901 131 4918 165
rect 4850 91 4918 131
rect 3888 17 3956 57
rect 4850 57 4867 91
rect 4901 57 4918 91
rect 5516 313 5584 353
rect 6478 427 6495 461
rect 6529 427 6546 461
rect 7440 461 7508 482
rect 6478 387 6546 427
rect 6478 353 6495 387
rect 6529 353 6546 387
rect 5516 279 5533 313
rect 5567 279 5584 313
rect 5516 239 5584 279
rect 5516 205 5533 239
rect 5567 205 5584 239
rect 5516 165 5584 205
rect 5516 131 5533 165
rect 5567 131 5584 165
rect 5516 91 5584 131
rect 4850 17 4918 57
rect 5516 57 5533 91
rect 5567 57 5584 91
rect 6478 313 6546 353
rect 7440 427 7457 461
rect 7491 427 7508 461
rect 8106 461 8174 482
rect 7440 387 7508 427
rect 7440 353 7457 387
rect 7491 353 7508 387
rect 6478 279 6495 313
rect 6529 279 6546 313
rect 6478 239 6546 279
rect 6478 205 6495 239
rect 6529 205 6546 239
rect 6478 165 6546 205
rect 6478 131 6495 165
rect 6529 131 6546 165
rect 6478 91 6546 131
rect 5516 17 5584 57
rect 6478 57 6495 91
rect 6529 57 6546 91
rect 7440 313 7508 353
rect 8106 427 8123 461
rect 8157 427 8174 461
rect 8772 461 8840 482
rect 8106 387 8174 427
rect 8106 353 8123 387
rect 8157 353 8174 387
rect 7440 279 7457 313
rect 7491 279 7508 313
rect 7440 239 7508 279
rect 7440 205 7457 239
rect 7491 205 7508 239
rect 7440 165 7508 205
rect 7440 131 7457 165
rect 7491 131 7508 165
rect 7440 91 7508 131
rect 6478 17 6546 57
rect 7440 57 7457 91
rect 7491 57 7508 91
rect 8106 313 8174 353
rect 8772 427 8789 461
rect 8823 427 8840 461
rect 9734 461 9802 482
rect 8772 387 8840 427
rect 8772 353 8789 387
rect 8823 353 8840 387
rect 8106 279 8123 313
rect 8157 279 8174 313
rect 8106 239 8174 279
rect 8106 205 8123 239
rect 8157 205 8174 239
rect 8106 165 8174 205
rect 8106 131 8123 165
rect 8157 131 8174 165
rect 8106 91 8174 131
rect 7440 17 7508 57
rect 8106 57 8123 91
rect 8157 57 8174 91
rect 8772 313 8840 353
rect 9734 427 9751 461
rect 9785 427 9802 461
rect 10400 461 10468 482
rect 9734 387 9802 427
rect 9734 353 9751 387
rect 9785 353 9802 387
rect 8772 279 8789 313
rect 8823 279 8840 313
rect 8772 239 8840 279
rect 8772 205 8789 239
rect 8823 205 8840 239
rect 8772 165 8840 205
rect 8772 131 8789 165
rect 8823 131 8840 165
rect 8772 91 8840 131
rect 8106 17 8174 57
rect 8772 57 8789 91
rect 8823 57 8840 91
rect 9734 313 9802 353
rect 10400 427 10417 461
rect 10451 427 10468 461
rect 11362 461 11430 482
rect 10400 387 10468 427
rect 10400 353 10417 387
rect 10451 353 10468 387
rect 9734 279 9751 313
rect 9785 279 9802 313
rect 9734 239 9802 279
rect 9734 205 9751 239
rect 9785 205 9802 239
rect 9734 165 9802 205
rect 9734 131 9751 165
rect 9785 131 9802 165
rect 9734 91 9802 131
rect 8772 17 8840 57
rect 9734 57 9751 91
rect 9785 57 9802 91
rect 10400 313 10468 353
rect 11362 427 11379 461
rect 11413 427 11430 461
rect 12324 461 12392 482
rect 11362 387 11430 427
rect 11362 353 11379 387
rect 11413 353 11430 387
rect 10400 279 10417 313
rect 10451 279 10468 313
rect 10400 239 10468 279
rect 10400 205 10417 239
rect 10451 205 10468 239
rect 10400 165 10468 205
rect 10400 131 10417 165
rect 10451 131 10468 165
rect 10400 91 10468 131
rect 9734 17 9802 57
rect 10400 57 10417 91
rect 10451 57 10468 91
rect 11362 313 11430 353
rect 12324 427 12341 461
rect 12375 427 12392 461
rect 12990 461 13058 482
rect 12324 387 12392 427
rect 12324 353 12341 387
rect 12375 353 12392 387
rect 11362 279 11379 313
rect 11413 279 11430 313
rect 11362 239 11430 279
rect 11362 205 11379 239
rect 11413 205 11430 239
rect 11362 165 11430 205
rect 11362 131 11379 165
rect 11413 131 11430 165
rect 11362 91 11430 131
rect 10400 17 10468 57
rect 11362 57 11379 91
rect 11413 57 11430 91
rect 12324 313 12392 353
rect 12990 427 13007 461
rect 13041 427 13058 461
rect 13656 461 13724 482
rect 12990 387 13058 427
rect 12990 353 13007 387
rect 13041 353 13058 387
rect 12324 279 12341 313
rect 12375 279 12392 313
rect 12324 239 12392 279
rect 12324 205 12341 239
rect 12375 205 12392 239
rect 12324 165 12392 205
rect 12324 131 12341 165
rect 12375 131 12392 165
rect 12324 91 12392 131
rect 11362 17 11430 57
rect 12324 57 12341 91
rect 12375 57 12392 91
rect 12990 313 13058 353
rect 13656 427 13673 461
rect 13707 427 13724 461
rect 14618 461 14686 482
rect 13656 387 13724 427
rect 13656 353 13673 387
rect 13707 353 13724 387
rect 12990 279 13007 313
rect 13041 279 13058 313
rect 12990 239 13058 279
rect 12990 205 13007 239
rect 13041 205 13058 239
rect 12990 165 13058 205
rect 12990 131 13007 165
rect 13041 131 13058 165
rect 12990 91 13058 131
rect 12324 17 12392 57
rect 12990 57 13007 91
rect 13041 57 13058 91
rect 13656 313 13724 353
rect 14618 427 14635 461
rect 14669 427 14686 461
rect 15284 461 15352 482
rect 14618 387 14686 427
rect 14618 353 14635 387
rect 14669 353 14686 387
rect 15284 427 15301 461
rect 15335 427 15352 461
rect 15950 461 16018 482
rect 15284 387 15352 427
rect 13656 279 13673 313
rect 13707 279 13724 313
rect 13656 239 13724 279
rect 13656 205 13673 239
rect 13707 205 13724 239
rect 13656 165 13724 205
rect 13656 131 13673 165
rect 13707 131 13724 165
rect 13656 91 13724 131
rect 12990 17 13058 57
rect 13656 57 13673 91
rect 13707 57 13724 91
rect 14618 313 14686 353
rect 15284 353 15301 387
rect 15335 353 15352 387
rect 14618 279 14635 313
rect 14669 279 14686 313
rect 14618 239 14686 279
rect 14618 205 14635 239
rect 14669 205 14686 239
rect 14618 165 14686 205
rect 14618 131 14635 165
rect 14669 131 14686 165
rect 14618 91 14686 131
rect 13656 17 13724 57
rect 14618 57 14635 91
rect 14669 57 14686 91
rect 15284 313 15352 353
rect 15950 427 15967 461
rect 16001 427 16018 461
rect 16616 461 16684 482
rect 15950 387 16018 427
rect 15950 353 15967 387
rect 16001 353 16018 387
rect 16616 427 16633 461
rect 16667 427 16684 461
rect 17060 461 17128 482
rect 16616 387 16684 427
rect 15284 279 15301 313
rect 15335 279 15352 313
rect 15284 239 15352 279
rect 15284 205 15301 239
rect 15335 205 15352 239
rect 15284 165 15352 205
rect 15284 131 15301 165
rect 15335 131 15352 165
rect 15284 91 15352 131
rect 14618 17 14686 57
rect 15284 57 15301 91
rect 15335 57 15352 91
rect 15950 313 16018 353
rect 16616 353 16633 387
rect 16667 353 16684 387
rect 17060 427 17077 461
rect 17111 427 17128 461
rect 15950 279 15967 313
rect 16001 279 16018 313
rect 15950 239 16018 279
rect 15950 205 15967 239
rect 16001 205 16018 239
rect 15950 165 16018 205
rect 15950 131 15967 165
rect 16001 131 16018 165
rect 15950 91 16018 131
rect 15284 17 15352 57
rect 15950 57 15967 91
rect 16001 57 16018 91
rect 16616 313 16684 353
rect 17060 387 17128 427
rect 17060 353 17077 387
rect 17111 353 17128 387
rect 16616 279 16633 313
rect 16667 279 16684 313
rect 16616 239 16684 279
rect 16616 205 16633 239
rect 16667 205 16684 239
rect 16616 165 16684 205
rect 16616 131 16633 165
rect 16667 131 16684 165
rect 16616 91 16684 131
rect 15950 17 16018 57
rect 16616 57 16633 91
rect 16667 57 16684 91
rect 17060 313 17128 353
rect 17060 279 17077 313
rect 17111 279 17128 313
rect 17060 239 17128 279
rect 17060 205 17077 239
rect 17111 205 17128 239
rect 17060 165 17128 205
rect 17060 131 17077 165
rect 17111 131 17128 165
rect 17060 91 17128 131
rect 16616 17 16684 57
rect 17060 57 17077 91
rect 17111 57 17128 91
rect 17060 17 17128 57
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5163 17
rect 5197 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5755 17
rect 5789 -17 5829 17
rect 5863 -17 5903 17
rect 5937 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6125 17
rect 6159 -17 6199 17
rect 6233 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6569 17
rect 6603 -17 6643 17
rect 6677 -17 6717 17
rect 6751 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7087 17
rect 7121 -17 7161 17
rect 7195 -17 7235 17
rect 7269 -17 7309 17
rect 7343 -17 7383 17
rect 7417 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7679 17
rect 7713 -17 7753 17
rect 7787 -17 7827 17
rect 7861 -17 7901 17
rect 7935 -17 7975 17
rect 8009 -17 8049 17
rect 8083 -17 8197 17
rect 8231 -17 8271 17
rect 8305 -17 8345 17
rect 8379 -17 8419 17
rect 8453 -17 8493 17
rect 8527 -17 8567 17
rect 8601 -17 8641 17
rect 8675 -17 8715 17
rect 8749 -17 8863 17
rect 8897 -17 8937 17
rect 8971 -17 9011 17
rect 9045 -17 9085 17
rect 9119 -17 9159 17
rect 9193 -17 9233 17
rect 9267 -17 9307 17
rect 9341 -17 9381 17
rect 9415 -17 9455 17
rect 9489 -17 9529 17
rect 9563 -17 9603 17
rect 9637 -17 9677 17
rect 9711 -17 9825 17
rect 9859 -17 9899 17
rect 9933 -17 9973 17
rect 10007 -17 10047 17
rect 10081 -17 10121 17
rect 10155 -17 10195 17
rect 10229 -17 10269 17
rect 10303 -17 10343 17
rect 10377 -17 10491 17
rect 10525 -17 10565 17
rect 10599 -17 10639 17
rect 10673 -17 10713 17
rect 10747 -17 10787 17
rect 10821 -17 10861 17
rect 10895 -17 10935 17
rect 10969 -17 11009 17
rect 11043 -17 11083 17
rect 11117 -17 11157 17
rect 11191 -17 11231 17
rect 11265 -17 11305 17
rect 11339 -17 11453 17
rect 11487 -17 11527 17
rect 11561 -17 11601 17
rect 11635 -17 11675 17
rect 11709 -17 11749 17
rect 11783 -17 11823 17
rect 11857 -17 11897 17
rect 11931 -17 11971 17
rect 12005 -17 12045 17
rect 12079 -17 12119 17
rect 12153 -17 12193 17
rect 12227 -17 12267 17
rect 12301 -17 12415 17
rect 12449 -17 12489 17
rect 12523 -17 12563 17
rect 12597 -17 12637 17
rect 12671 -17 12711 17
rect 12745 -17 12785 17
rect 12819 -17 12859 17
rect 12893 -17 12933 17
rect 12967 -17 13081 17
rect 13115 -17 13155 17
rect 13189 -17 13229 17
rect 13263 -17 13303 17
rect 13337 -17 13377 17
rect 13411 -17 13451 17
rect 13485 -17 13525 17
rect 13559 -17 13599 17
rect 13633 -17 13747 17
rect 13781 -17 13821 17
rect 13855 -17 13895 17
rect 13929 -17 13969 17
rect 14003 -17 14043 17
rect 14077 -17 14117 17
rect 14151 -17 14191 17
rect 14225 -17 14265 17
rect 14299 -17 14339 17
rect 14373 -17 14413 17
rect 14447 -17 14487 17
rect 14521 -17 14561 17
rect 14595 -17 14709 17
rect 14743 -17 14783 17
rect 14817 -17 14857 17
rect 14891 -17 14931 17
rect 14965 -17 15005 17
rect 15039 -17 15079 17
rect 15113 -17 15153 17
rect 15187 -17 15227 17
rect 15261 -17 15375 17
rect 15409 -17 15449 17
rect 15483 -17 15523 17
rect 15557 -17 15597 17
rect 15631 -17 15671 17
rect 15705 -17 15745 17
rect 15779 -17 15819 17
rect 15853 -17 15893 17
rect 15927 -17 16041 17
rect 16075 -17 16115 17
rect 16149 -17 16189 17
rect 16223 -17 16263 17
rect 16297 -17 16337 17
rect 16371 -17 16411 17
rect 16445 -17 16485 17
rect 16519 -17 16559 17
rect 16593 -17 16707 17
rect 16741 -17 16781 17
rect 16815 -17 16855 17
rect 16889 -17 16929 17
rect 16963 -17 17003 17
rect 17037 -17 17128 17
rect -34 -34 17128 -17
<< nsubdiff >>
rect -34 1497 17128 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5163 1497
rect 5197 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5755 1497
rect 5789 1463 5829 1497
rect 5863 1463 5903 1497
rect 5937 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6125 1497
rect 6159 1463 6199 1497
rect 6233 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6569 1497
rect 6603 1463 6643 1497
rect 6677 1463 6717 1497
rect 6751 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7087 1497
rect 7121 1463 7161 1497
rect 7195 1463 7235 1497
rect 7269 1463 7309 1497
rect 7343 1463 7383 1497
rect 7417 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7679 1497
rect 7713 1463 7753 1497
rect 7787 1463 7827 1497
rect 7861 1463 7901 1497
rect 7935 1463 7975 1497
rect 8009 1463 8049 1497
rect 8083 1463 8197 1497
rect 8231 1463 8271 1497
rect 8305 1463 8345 1497
rect 8379 1463 8419 1497
rect 8453 1463 8493 1497
rect 8527 1463 8567 1497
rect 8601 1463 8641 1497
rect 8675 1463 8715 1497
rect 8749 1463 8863 1497
rect 8897 1463 8937 1497
rect 8971 1463 9011 1497
rect 9045 1463 9085 1497
rect 9119 1463 9159 1497
rect 9193 1463 9233 1497
rect 9267 1463 9307 1497
rect 9341 1463 9381 1497
rect 9415 1463 9455 1497
rect 9489 1463 9529 1497
rect 9563 1463 9603 1497
rect 9637 1463 9677 1497
rect 9711 1463 9825 1497
rect 9859 1463 9899 1497
rect 9933 1463 9973 1497
rect 10007 1463 10047 1497
rect 10081 1463 10121 1497
rect 10155 1463 10195 1497
rect 10229 1463 10269 1497
rect 10303 1463 10343 1497
rect 10377 1463 10491 1497
rect 10525 1463 10565 1497
rect 10599 1463 10639 1497
rect 10673 1463 10713 1497
rect 10747 1463 10787 1497
rect 10821 1463 10861 1497
rect 10895 1463 10935 1497
rect 10969 1463 11009 1497
rect 11043 1463 11083 1497
rect 11117 1463 11157 1497
rect 11191 1463 11231 1497
rect 11265 1463 11305 1497
rect 11339 1463 11453 1497
rect 11487 1463 11527 1497
rect 11561 1463 11601 1497
rect 11635 1463 11675 1497
rect 11709 1463 11749 1497
rect 11783 1463 11823 1497
rect 11857 1463 11897 1497
rect 11931 1463 11971 1497
rect 12005 1463 12045 1497
rect 12079 1463 12119 1497
rect 12153 1463 12193 1497
rect 12227 1463 12267 1497
rect 12301 1463 12415 1497
rect 12449 1463 12489 1497
rect 12523 1463 12563 1497
rect 12597 1463 12637 1497
rect 12671 1463 12711 1497
rect 12745 1463 12785 1497
rect 12819 1463 12859 1497
rect 12893 1463 12933 1497
rect 12967 1463 13081 1497
rect 13115 1463 13155 1497
rect 13189 1463 13229 1497
rect 13263 1463 13303 1497
rect 13337 1463 13377 1497
rect 13411 1463 13451 1497
rect 13485 1463 13525 1497
rect 13559 1463 13599 1497
rect 13633 1463 13747 1497
rect 13781 1463 13821 1497
rect 13855 1463 13895 1497
rect 13929 1463 13969 1497
rect 14003 1463 14043 1497
rect 14077 1463 14117 1497
rect 14151 1463 14191 1497
rect 14225 1463 14265 1497
rect 14299 1463 14339 1497
rect 14373 1463 14413 1497
rect 14447 1463 14487 1497
rect 14521 1463 14561 1497
rect 14595 1463 14709 1497
rect 14743 1463 14783 1497
rect 14817 1463 14857 1497
rect 14891 1463 14931 1497
rect 14965 1463 15005 1497
rect 15039 1463 15079 1497
rect 15113 1463 15153 1497
rect 15187 1463 15227 1497
rect 15261 1463 15375 1497
rect 15409 1463 15449 1497
rect 15483 1463 15523 1497
rect 15557 1463 15597 1497
rect 15631 1463 15671 1497
rect 15705 1463 15745 1497
rect 15779 1463 15819 1497
rect 15853 1463 15893 1497
rect 15927 1463 16041 1497
rect 16075 1463 16115 1497
rect 16149 1463 16189 1497
rect 16223 1463 16263 1497
rect 16297 1463 16337 1497
rect 16371 1463 16411 1497
rect 16445 1463 16485 1497
rect 16519 1463 16559 1497
rect 16593 1463 16707 1497
rect 16741 1463 16781 1497
rect 16815 1463 16855 1497
rect 16889 1463 16929 1497
rect 16963 1463 17003 1497
rect 17037 1463 17128 1497
rect -34 1423 34 1463
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect 632 1423 700 1463
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect -34 979 34 1019
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 1594 1423 1662 1463
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect 632 979 700 1019
rect 1594 1389 1611 1423
rect 1645 1389 1662 1423
rect 2556 1423 2624 1463
rect 1594 1349 1662 1389
rect 1594 1315 1611 1349
rect 1645 1315 1662 1349
rect 1594 1275 1662 1315
rect 1594 1241 1611 1275
rect 1645 1241 1662 1275
rect 1594 1201 1662 1241
rect 1594 1167 1611 1201
rect 1645 1167 1662 1201
rect 1594 1127 1662 1167
rect 1594 1093 1611 1127
rect 1645 1093 1662 1127
rect 1594 1053 1662 1093
rect 1594 1019 1611 1053
rect 1645 1019 1662 1053
rect 632 945 649 979
rect 683 945 700 979
rect -34 871 -17 905
rect 17 884 34 905
rect 632 905 700 945
rect 1594 979 1662 1019
rect 2556 1389 2573 1423
rect 2607 1389 2624 1423
rect 3222 1423 3290 1463
rect 2556 1349 2624 1389
rect 2556 1315 2573 1349
rect 2607 1315 2624 1349
rect 2556 1275 2624 1315
rect 2556 1241 2573 1275
rect 2607 1241 2624 1275
rect 2556 1201 2624 1241
rect 2556 1167 2573 1201
rect 2607 1167 2624 1201
rect 2556 1127 2624 1167
rect 2556 1093 2573 1127
rect 2607 1093 2624 1127
rect 2556 1053 2624 1093
rect 2556 1019 2573 1053
rect 2607 1019 2624 1053
rect 1594 945 1611 979
rect 1645 945 1662 979
rect 632 884 649 905
rect 17 871 649 884
rect 683 884 700 905
rect 1594 905 1662 945
rect 2556 979 2624 1019
rect 3222 1389 3239 1423
rect 3273 1389 3290 1423
rect 3888 1423 3956 1463
rect 3222 1349 3290 1389
rect 3222 1315 3239 1349
rect 3273 1315 3290 1349
rect 3222 1275 3290 1315
rect 3222 1241 3239 1275
rect 3273 1241 3290 1275
rect 3222 1201 3290 1241
rect 3222 1167 3239 1201
rect 3273 1167 3290 1201
rect 3222 1127 3290 1167
rect 3222 1093 3239 1127
rect 3273 1093 3290 1127
rect 3222 1053 3290 1093
rect 3222 1019 3239 1053
rect 3273 1019 3290 1053
rect 2556 945 2573 979
rect 2607 945 2624 979
rect 1594 884 1611 905
rect 683 871 1611 884
rect 1645 884 1662 905
rect 2556 905 2624 945
rect 3222 979 3290 1019
rect 3888 1389 3905 1423
rect 3939 1389 3956 1423
rect 4850 1423 4918 1463
rect 3888 1349 3956 1389
rect 3888 1315 3905 1349
rect 3939 1315 3956 1349
rect 3888 1275 3956 1315
rect 3888 1241 3905 1275
rect 3939 1241 3956 1275
rect 3888 1201 3956 1241
rect 3888 1167 3905 1201
rect 3939 1167 3956 1201
rect 3888 1127 3956 1167
rect 3888 1093 3905 1127
rect 3939 1093 3956 1127
rect 3888 1053 3956 1093
rect 3888 1019 3905 1053
rect 3939 1019 3956 1053
rect 3222 945 3239 979
rect 3273 945 3290 979
rect 2556 884 2573 905
rect 1645 871 2573 884
rect 2607 884 2624 905
rect 3222 905 3290 945
rect 3888 979 3956 1019
rect 4850 1389 4867 1423
rect 4901 1389 4918 1423
rect 5516 1423 5584 1463
rect 4850 1349 4918 1389
rect 4850 1315 4867 1349
rect 4901 1315 4918 1349
rect 4850 1275 4918 1315
rect 4850 1241 4867 1275
rect 4901 1241 4918 1275
rect 4850 1201 4918 1241
rect 4850 1167 4867 1201
rect 4901 1167 4918 1201
rect 4850 1127 4918 1167
rect 4850 1093 4867 1127
rect 4901 1093 4918 1127
rect 4850 1053 4918 1093
rect 4850 1019 4867 1053
rect 4901 1019 4918 1053
rect 3888 945 3905 979
rect 3939 945 3956 979
rect 3222 884 3239 905
rect 2607 871 3239 884
rect 3273 884 3290 905
rect 3888 905 3956 945
rect 4850 979 4918 1019
rect 5516 1389 5533 1423
rect 5567 1389 5584 1423
rect 6478 1423 6546 1463
rect 5516 1349 5584 1389
rect 5516 1315 5533 1349
rect 5567 1315 5584 1349
rect 5516 1275 5584 1315
rect 5516 1241 5533 1275
rect 5567 1241 5584 1275
rect 5516 1201 5584 1241
rect 5516 1167 5533 1201
rect 5567 1167 5584 1201
rect 5516 1127 5584 1167
rect 5516 1093 5533 1127
rect 5567 1093 5584 1127
rect 5516 1053 5584 1093
rect 5516 1019 5533 1053
rect 5567 1019 5584 1053
rect 4850 945 4867 979
rect 4901 945 4918 979
rect 3888 884 3905 905
rect 3273 871 3905 884
rect 3939 884 3956 905
rect 4850 905 4918 945
rect 5516 979 5584 1019
rect 6478 1389 6495 1423
rect 6529 1389 6546 1423
rect 7440 1423 7508 1463
rect 6478 1349 6546 1389
rect 6478 1315 6495 1349
rect 6529 1315 6546 1349
rect 6478 1275 6546 1315
rect 6478 1241 6495 1275
rect 6529 1241 6546 1275
rect 6478 1201 6546 1241
rect 6478 1167 6495 1201
rect 6529 1167 6546 1201
rect 6478 1127 6546 1167
rect 6478 1093 6495 1127
rect 6529 1093 6546 1127
rect 6478 1053 6546 1093
rect 6478 1019 6495 1053
rect 6529 1019 6546 1053
rect 5516 945 5533 979
rect 5567 945 5584 979
rect 4850 884 4867 905
rect 3939 871 4867 884
rect 4901 884 4918 905
rect 5516 905 5584 945
rect 6478 979 6546 1019
rect 7440 1389 7457 1423
rect 7491 1389 7508 1423
rect 8106 1423 8174 1463
rect 7440 1349 7508 1389
rect 7440 1315 7457 1349
rect 7491 1315 7508 1349
rect 7440 1275 7508 1315
rect 7440 1241 7457 1275
rect 7491 1241 7508 1275
rect 7440 1201 7508 1241
rect 7440 1167 7457 1201
rect 7491 1167 7508 1201
rect 7440 1127 7508 1167
rect 7440 1093 7457 1127
rect 7491 1093 7508 1127
rect 7440 1053 7508 1093
rect 7440 1019 7457 1053
rect 7491 1019 7508 1053
rect 6478 945 6495 979
rect 6529 945 6546 979
rect 5516 884 5533 905
rect 4901 871 5533 884
rect 5567 884 5584 905
rect 6478 905 6546 945
rect 7440 979 7508 1019
rect 8106 1389 8123 1423
rect 8157 1389 8174 1423
rect 8772 1423 8840 1463
rect 8106 1349 8174 1389
rect 8106 1315 8123 1349
rect 8157 1315 8174 1349
rect 8106 1275 8174 1315
rect 8106 1241 8123 1275
rect 8157 1241 8174 1275
rect 8106 1201 8174 1241
rect 8106 1167 8123 1201
rect 8157 1167 8174 1201
rect 8106 1127 8174 1167
rect 8106 1093 8123 1127
rect 8157 1093 8174 1127
rect 8106 1053 8174 1093
rect 8106 1019 8123 1053
rect 8157 1019 8174 1053
rect 7440 945 7457 979
rect 7491 945 7508 979
rect 6478 884 6495 905
rect 5567 871 6495 884
rect 6529 884 6546 905
rect 7440 905 7508 945
rect 8106 979 8174 1019
rect 8772 1389 8789 1423
rect 8823 1389 8840 1423
rect 9734 1423 9802 1463
rect 8772 1349 8840 1389
rect 8772 1315 8789 1349
rect 8823 1315 8840 1349
rect 8772 1275 8840 1315
rect 8772 1241 8789 1275
rect 8823 1241 8840 1275
rect 8772 1201 8840 1241
rect 8772 1167 8789 1201
rect 8823 1167 8840 1201
rect 8772 1127 8840 1167
rect 8772 1093 8789 1127
rect 8823 1093 8840 1127
rect 8772 1053 8840 1093
rect 8772 1019 8789 1053
rect 8823 1019 8840 1053
rect 8106 945 8123 979
rect 8157 945 8174 979
rect 7440 884 7457 905
rect 6529 871 7457 884
rect 7491 884 7508 905
rect 8106 905 8174 945
rect 8772 979 8840 1019
rect 9734 1389 9751 1423
rect 9785 1389 9802 1423
rect 10400 1423 10468 1463
rect 9734 1349 9802 1389
rect 9734 1315 9751 1349
rect 9785 1315 9802 1349
rect 9734 1275 9802 1315
rect 9734 1241 9751 1275
rect 9785 1241 9802 1275
rect 9734 1201 9802 1241
rect 9734 1167 9751 1201
rect 9785 1167 9802 1201
rect 9734 1127 9802 1167
rect 9734 1093 9751 1127
rect 9785 1093 9802 1127
rect 9734 1053 9802 1093
rect 9734 1019 9751 1053
rect 9785 1019 9802 1053
rect 8772 945 8789 979
rect 8823 945 8840 979
rect 8106 884 8123 905
rect 7491 871 8123 884
rect 8157 884 8174 905
rect 8772 905 8840 945
rect 9734 979 9802 1019
rect 10400 1389 10417 1423
rect 10451 1389 10468 1423
rect 11362 1423 11430 1463
rect 10400 1349 10468 1389
rect 10400 1315 10417 1349
rect 10451 1315 10468 1349
rect 10400 1275 10468 1315
rect 10400 1241 10417 1275
rect 10451 1241 10468 1275
rect 10400 1201 10468 1241
rect 10400 1167 10417 1201
rect 10451 1167 10468 1201
rect 10400 1127 10468 1167
rect 10400 1093 10417 1127
rect 10451 1093 10468 1127
rect 10400 1053 10468 1093
rect 10400 1019 10417 1053
rect 10451 1019 10468 1053
rect 9734 945 9751 979
rect 9785 945 9802 979
rect 8772 884 8789 905
rect 8157 871 8789 884
rect 8823 884 8840 905
rect 9734 905 9802 945
rect 10400 979 10468 1019
rect 11362 1389 11379 1423
rect 11413 1389 11430 1423
rect 12324 1423 12392 1463
rect 11362 1349 11430 1389
rect 11362 1315 11379 1349
rect 11413 1315 11430 1349
rect 11362 1275 11430 1315
rect 11362 1241 11379 1275
rect 11413 1241 11430 1275
rect 11362 1201 11430 1241
rect 11362 1167 11379 1201
rect 11413 1167 11430 1201
rect 11362 1127 11430 1167
rect 11362 1093 11379 1127
rect 11413 1093 11430 1127
rect 11362 1053 11430 1093
rect 11362 1019 11379 1053
rect 11413 1019 11430 1053
rect 10400 945 10417 979
rect 10451 945 10468 979
rect 9734 884 9751 905
rect 8823 871 9751 884
rect 9785 884 9802 905
rect 10400 905 10468 945
rect 11362 979 11430 1019
rect 12324 1389 12341 1423
rect 12375 1389 12392 1423
rect 12990 1423 13058 1463
rect 12324 1349 12392 1389
rect 12324 1315 12341 1349
rect 12375 1315 12392 1349
rect 12324 1275 12392 1315
rect 12324 1241 12341 1275
rect 12375 1241 12392 1275
rect 12324 1201 12392 1241
rect 12324 1167 12341 1201
rect 12375 1167 12392 1201
rect 12324 1127 12392 1167
rect 12324 1093 12341 1127
rect 12375 1093 12392 1127
rect 12324 1053 12392 1093
rect 12324 1019 12341 1053
rect 12375 1019 12392 1053
rect 11362 945 11379 979
rect 11413 945 11430 979
rect 10400 884 10417 905
rect 9785 871 10417 884
rect 10451 884 10468 905
rect 11362 905 11430 945
rect 12324 979 12392 1019
rect 12990 1389 13007 1423
rect 13041 1389 13058 1423
rect 13656 1423 13724 1463
rect 12990 1349 13058 1389
rect 12990 1315 13007 1349
rect 13041 1315 13058 1349
rect 12990 1275 13058 1315
rect 12990 1241 13007 1275
rect 13041 1241 13058 1275
rect 12990 1201 13058 1241
rect 12990 1167 13007 1201
rect 13041 1167 13058 1201
rect 12990 1127 13058 1167
rect 12990 1093 13007 1127
rect 13041 1093 13058 1127
rect 12990 1053 13058 1093
rect 12990 1019 13007 1053
rect 13041 1019 13058 1053
rect 12324 945 12341 979
rect 12375 945 12392 979
rect 11362 884 11379 905
rect 10451 871 11379 884
rect 11413 884 11430 905
rect 12324 905 12392 945
rect 12990 979 13058 1019
rect 13656 1389 13673 1423
rect 13707 1389 13724 1423
rect 14618 1423 14686 1463
rect 13656 1349 13724 1389
rect 13656 1315 13673 1349
rect 13707 1315 13724 1349
rect 13656 1275 13724 1315
rect 13656 1241 13673 1275
rect 13707 1241 13724 1275
rect 13656 1201 13724 1241
rect 13656 1167 13673 1201
rect 13707 1167 13724 1201
rect 13656 1127 13724 1167
rect 13656 1093 13673 1127
rect 13707 1093 13724 1127
rect 13656 1053 13724 1093
rect 13656 1019 13673 1053
rect 13707 1019 13724 1053
rect 12990 945 13007 979
rect 13041 945 13058 979
rect 12324 884 12341 905
rect 11413 871 12341 884
rect 12375 884 12392 905
rect 12990 905 13058 945
rect 13656 979 13724 1019
rect 14618 1389 14635 1423
rect 14669 1389 14686 1423
rect 15284 1423 15352 1463
rect 14618 1349 14686 1389
rect 14618 1315 14635 1349
rect 14669 1315 14686 1349
rect 14618 1275 14686 1315
rect 14618 1241 14635 1275
rect 14669 1241 14686 1275
rect 14618 1201 14686 1241
rect 14618 1167 14635 1201
rect 14669 1167 14686 1201
rect 14618 1127 14686 1167
rect 14618 1093 14635 1127
rect 14669 1093 14686 1127
rect 14618 1053 14686 1093
rect 14618 1019 14635 1053
rect 14669 1019 14686 1053
rect 13656 945 13673 979
rect 13707 945 13724 979
rect 12990 884 13007 905
rect 12375 871 13007 884
rect 13041 884 13058 905
rect 13656 905 13724 945
rect 14618 979 14686 1019
rect 15284 1389 15301 1423
rect 15335 1389 15352 1423
rect 15950 1423 16018 1463
rect 16598 1459 16684 1463
rect 15284 1349 15352 1389
rect 15284 1315 15301 1349
rect 15335 1315 15352 1349
rect 15284 1275 15352 1315
rect 15284 1241 15301 1275
rect 15335 1241 15352 1275
rect 15284 1201 15352 1241
rect 15284 1167 15301 1201
rect 15335 1167 15352 1201
rect 15284 1127 15352 1167
rect 15284 1093 15301 1127
rect 15335 1093 15352 1127
rect 15284 1053 15352 1093
rect 15284 1019 15301 1053
rect 15335 1019 15352 1053
rect 14618 945 14635 979
rect 14669 945 14686 979
rect 13656 884 13673 905
rect 13041 871 13673 884
rect 13707 884 13724 905
rect 14618 905 14686 945
rect 15284 979 15352 1019
rect 15950 1389 15967 1423
rect 16001 1389 16018 1423
rect 16616 1423 16684 1459
rect 15950 1349 16018 1389
rect 15950 1315 15967 1349
rect 16001 1315 16018 1349
rect 15950 1275 16018 1315
rect 15950 1241 15967 1275
rect 16001 1241 16018 1275
rect 15950 1201 16018 1241
rect 15950 1167 15967 1201
rect 16001 1167 16018 1201
rect 15950 1127 16018 1167
rect 15950 1093 15967 1127
rect 16001 1093 16018 1127
rect 15950 1053 16018 1093
rect 15950 1019 15967 1053
rect 16001 1019 16018 1053
rect 15284 945 15301 979
rect 15335 945 15352 979
rect 14618 884 14635 905
rect 13707 871 14635 884
rect 14669 884 14686 905
rect 15284 905 15352 945
rect 15950 979 16018 1019
rect 16616 1389 16633 1423
rect 16667 1389 16684 1423
rect 17060 1423 17128 1463
rect 16616 1349 16684 1389
rect 16616 1315 16633 1349
rect 16667 1315 16684 1349
rect 16616 1275 16684 1315
rect 16616 1241 16633 1275
rect 16667 1241 16684 1275
rect 16616 1201 16684 1241
rect 16616 1167 16633 1201
rect 16667 1167 16684 1201
rect 16616 1127 16684 1167
rect 16616 1093 16633 1127
rect 16667 1093 16684 1127
rect 16616 1053 16684 1093
rect 16616 1019 16633 1053
rect 16667 1019 16684 1053
rect 15950 945 15967 979
rect 16001 945 16018 979
rect 15284 884 15301 905
rect 14669 871 15301 884
rect 15335 884 15352 905
rect 15950 905 16018 945
rect 16616 979 16684 1019
rect 17060 1389 17077 1423
rect 17111 1389 17128 1423
rect 17060 1349 17128 1389
rect 17060 1315 17077 1349
rect 17111 1315 17128 1349
rect 17060 1275 17128 1315
rect 17060 1241 17077 1275
rect 17111 1241 17128 1275
rect 17060 1201 17128 1241
rect 17060 1167 17077 1201
rect 17111 1167 17128 1201
rect 17060 1127 17128 1167
rect 17060 1093 17077 1127
rect 17111 1093 17128 1127
rect 17060 1053 17128 1093
rect 17060 1019 17077 1053
rect 17111 1019 17128 1053
rect 16616 945 16633 979
rect 16667 945 16684 979
rect 15950 884 15967 905
rect 15335 871 15967 884
rect 16001 884 16018 905
rect 16616 905 16684 945
rect 17060 979 17128 1019
rect 17060 945 17077 979
rect 17111 945 17128 979
rect 16616 884 16633 905
rect 16001 871 16633 884
rect 16667 884 16684 905
rect 17060 905 17128 945
rect 17060 884 17077 905
rect 16667 871 17077 884
rect 17111 871 17128 905
rect -34 822 17128 871
<< psubdiffcont >>
rect -17 427 17 461
rect -17 353 17 387
rect 649 427 683 461
rect 649 353 683 387
rect -17 279 17 313
rect -17 205 17 239
rect -17 131 17 165
rect -17 57 17 91
rect 1611 427 1645 461
rect 1611 353 1645 387
rect 649 279 683 313
rect 649 205 683 239
rect 649 131 683 165
rect 649 57 683 91
rect 2573 427 2607 461
rect 2573 353 2607 387
rect 1611 279 1645 313
rect 1611 205 1645 239
rect 1611 131 1645 165
rect 1611 57 1645 91
rect 3239 427 3273 461
rect 3239 353 3273 387
rect 2573 279 2607 313
rect 2573 205 2607 239
rect 2573 131 2607 165
rect 2573 57 2607 91
rect 3905 427 3939 461
rect 3905 353 3939 387
rect 3239 279 3273 313
rect 3239 205 3273 239
rect 3239 131 3273 165
rect 3239 57 3273 91
rect 4867 427 4901 461
rect 4867 353 4901 387
rect 3905 279 3939 313
rect 3905 205 3939 239
rect 3905 131 3939 165
rect 3905 57 3939 91
rect 5533 427 5567 461
rect 5533 353 5567 387
rect 4867 279 4901 313
rect 4867 205 4901 239
rect 4867 131 4901 165
rect 4867 57 4901 91
rect 6495 427 6529 461
rect 6495 353 6529 387
rect 5533 279 5567 313
rect 5533 205 5567 239
rect 5533 131 5567 165
rect 5533 57 5567 91
rect 7457 427 7491 461
rect 7457 353 7491 387
rect 6495 279 6529 313
rect 6495 205 6529 239
rect 6495 131 6529 165
rect 6495 57 6529 91
rect 8123 427 8157 461
rect 8123 353 8157 387
rect 7457 279 7491 313
rect 7457 205 7491 239
rect 7457 131 7491 165
rect 7457 57 7491 91
rect 8789 427 8823 461
rect 8789 353 8823 387
rect 8123 279 8157 313
rect 8123 205 8157 239
rect 8123 131 8157 165
rect 8123 57 8157 91
rect 9751 427 9785 461
rect 9751 353 9785 387
rect 8789 279 8823 313
rect 8789 205 8823 239
rect 8789 131 8823 165
rect 8789 57 8823 91
rect 10417 427 10451 461
rect 10417 353 10451 387
rect 9751 279 9785 313
rect 9751 205 9785 239
rect 9751 131 9785 165
rect 9751 57 9785 91
rect 11379 427 11413 461
rect 11379 353 11413 387
rect 10417 279 10451 313
rect 10417 205 10451 239
rect 10417 131 10451 165
rect 10417 57 10451 91
rect 12341 427 12375 461
rect 12341 353 12375 387
rect 11379 279 11413 313
rect 11379 205 11413 239
rect 11379 131 11413 165
rect 11379 57 11413 91
rect 13007 427 13041 461
rect 13007 353 13041 387
rect 12341 279 12375 313
rect 12341 205 12375 239
rect 12341 131 12375 165
rect 12341 57 12375 91
rect 13673 427 13707 461
rect 13673 353 13707 387
rect 13007 279 13041 313
rect 13007 205 13041 239
rect 13007 131 13041 165
rect 13007 57 13041 91
rect 14635 427 14669 461
rect 14635 353 14669 387
rect 15301 427 15335 461
rect 13673 279 13707 313
rect 13673 205 13707 239
rect 13673 131 13707 165
rect 13673 57 13707 91
rect 15301 353 15335 387
rect 14635 279 14669 313
rect 14635 205 14669 239
rect 14635 131 14669 165
rect 14635 57 14669 91
rect 15967 427 16001 461
rect 15967 353 16001 387
rect 16633 427 16667 461
rect 15301 279 15335 313
rect 15301 205 15335 239
rect 15301 131 15335 165
rect 15301 57 15335 91
rect 16633 353 16667 387
rect 17077 427 17111 461
rect 15967 279 16001 313
rect 15967 205 16001 239
rect 15967 131 16001 165
rect 15967 57 16001 91
rect 17077 353 17111 387
rect 16633 279 16667 313
rect 16633 205 16667 239
rect 16633 131 16667 165
rect 16633 57 16667 91
rect 17077 279 17111 313
rect 17077 205 17111 239
rect 17077 131 17111 165
rect 17077 57 17111 91
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4497 -17 4531 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4793 -17 4827 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5089 -17 5123 17
rect 5163 -17 5197 17
rect 5237 -17 5271 17
rect 5311 -17 5345 17
rect 5385 -17 5419 17
rect 5459 -17 5493 17
rect 5607 -17 5641 17
rect 5681 -17 5715 17
rect 5755 -17 5789 17
rect 5829 -17 5863 17
rect 5903 -17 5937 17
rect 5977 -17 6011 17
rect 6051 -17 6085 17
rect 6125 -17 6159 17
rect 6199 -17 6233 17
rect 6273 -17 6307 17
rect 6347 -17 6381 17
rect 6421 -17 6455 17
rect 6569 -17 6603 17
rect 6643 -17 6677 17
rect 6717 -17 6751 17
rect 6791 -17 6825 17
rect 6865 -17 6899 17
rect 6939 -17 6973 17
rect 7013 -17 7047 17
rect 7087 -17 7121 17
rect 7161 -17 7195 17
rect 7235 -17 7269 17
rect 7309 -17 7343 17
rect 7383 -17 7417 17
rect 7531 -17 7565 17
rect 7605 -17 7639 17
rect 7679 -17 7713 17
rect 7753 -17 7787 17
rect 7827 -17 7861 17
rect 7901 -17 7935 17
rect 7975 -17 8009 17
rect 8049 -17 8083 17
rect 8197 -17 8231 17
rect 8271 -17 8305 17
rect 8345 -17 8379 17
rect 8419 -17 8453 17
rect 8493 -17 8527 17
rect 8567 -17 8601 17
rect 8641 -17 8675 17
rect 8715 -17 8749 17
rect 8863 -17 8897 17
rect 8937 -17 8971 17
rect 9011 -17 9045 17
rect 9085 -17 9119 17
rect 9159 -17 9193 17
rect 9233 -17 9267 17
rect 9307 -17 9341 17
rect 9381 -17 9415 17
rect 9455 -17 9489 17
rect 9529 -17 9563 17
rect 9603 -17 9637 17
rect 9677 -17 9711 17
rect 9825 -17 9859 17
rect 9899 -17 9933 17
rect 9973 -17 10007 17
rect 10047 -17 10081 17
rect 10121 -17 10155 17
rect 10195 -17 10229 17
rect 10269 -17 10303 17
rect 10343 -17 10377 17
rect 10491 -17 10525 17
rect 10565 -17 10599 17
rect 10639 -17 10673 17
rect 10713 -17 10747 17
rect 10787 -17 10821 17
rect 10861 -17 10895 17
rect 10935 -17 10969 17
rect 11009 -17 11043 17
rect 11083 -17 11117 17
rect 11157 -17 11191 17
rect 11231 -17 11265 17
rect 11305 -17 11339 17
rect 11453 -17 11487 17
rect 11527 -17 11561 17
rect 11601 -17 11635 17
rect 11675 -17 11709 17
rect 11749 -17 11783 17
rect 11823 -17 11857 17
rect 11897 -17 11931 17
rect 11971 -17 12005 17
rect 12045 -17 12079 17
rect 12119 -17 12153 17
rect 12193 -17 12227 17
rect 12267 -17 12301 17
rect 12415 -17 12449 17
rect 12489 -17 12523 17
rect 12563 -17 12597 17
rect 12637 -17 12671 17
rect 12711 -17 12745 17
rect 12785 -17 12819 17
rect 12859 -17 12893 17
rect 12933 -17 12967 17
rect 13081 -17 13115 17
rect 13155 -17 13189 17
rect 13229 -17 13263 17
rect 13303 -17 13337 17
rect 13377 -17 13411 17
rect 13451 -17 13485 17
rect 13525 -17 13559 17
rect 13599 -17 13633 17
rect 13747 -17 13781 17
rect 13821 -17 13855 17
rect 13895 -17 13929 17
rect 13969 -17 14003 17
rect 14043 -17 14077 17
rect 14117 -17 14151 17
rect 14191 -17 14225 17
rect 14265 -17 14299 17
rect 14339 -17 14373 17
rect 14413 -17 14447 17
rect 14487 -17 14521 17
rect 14561 -17 14595 17
rect 14709 -17 14743 17
rect 14783 -17 14817 17
rect 14857 -17 14891 17
rect 14931 -17 14965 17
rect 15005 -17 15039 17
rect 15079 -17 15113 17
rect 15153 -17 15187 17
rect 15227 -17 15261 17
rect 15375 -17 15409 17
rect 15449 -17 15483 17
rect 15523 -17 15557 17
rect 15597 -17 15631 17
rect 15671 -17 15705 17
rect 15745 -17 15779 17
rect 15819 -17 15853 17
rect 15893 -17 15927 17
rect 16041 -17 16075 17
rect 16115 -17 16149 17
rect 16189 -17 16223 17
rect 16263 -17 16297 17
rect 16337 -17 16371 17
rect 16411 -17 16445 17
rect 16485 -17 16519 17
rect 16559 -17 16593 17
rect 16707 -17 16741 17
rect 16781 -17 16815 17
rect 16855 -17 16889 17
rect 16929 -17 16963 17
rect 17003 -17 17037 17
<< nsubdiffcont >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4497 1463 4531 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4793 1463 4827 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5089 1463 5123 1497
rect 5163 1463 5197 1497
rect 5237 1463 5271 1497
rect 5311 1463 5345 1497
rect 5385 1463 5419 1497
rect 5459 1463 5493 1497
rect 5607 1463 5641 1497
rect 5681 1463 5715 1497
rect 5755 1463 5789 1497
rect 5829 1463 5863 1497
rect 5903 1463 5937 1497
rect 5977 1463 6011 1497
rect 6051 1463 6085 1497
rect 6125 1463 6159 1497
rect 6199 1463 6233 1497
rect 6273 1463 6307 1497
rect 6347 1463 6381 1497
rect 6421 1463 6455 1497
rect 6569 1463 6603 1497
rect 6643 1463 6677 1497
rect 6717 1463 6751 1497
rect 6791 1463 6825 1497
rect 6865 1463 6899 1497
rect 6939 1463 6973 1497
rect 7013 1463 7047 1497
rect 7087 1463 7121 1497
rect 7161 1463 7195 1497
rect 7235 1463 7269 1497
rect 7309 1463 7343 1497
rect 7383 1463 7417 1497
rect 7531 1463 7565 1497
rect 7605 1463 7639 1497
rect 7679 1463 7713 1497
rect 7753 1463 7787 1497
rect 7827 1463 7861 1497
rect 7901 1463 7935 1497
rect 7975 1463 8009 1497
rect 8049 1463 8083 1497
rect 8197 1463 8231 1497
rect 8271 1463 8305 1497
rect 8345 1463 8379 1497
rect 8419 1463 8453 1497
rect 8493 1463 8527 1497
rect 8567 1463 8601 1497
rect 8641 1463 8675 1497
rect 8715 1463 8749 1497
rect 8863 1463 8897 1497
rect 8937 1463 8971 1497
rect 9011 1463 9045 1497
rect 9085 1463 9119 1497
rect 9159 1463 9193 1497
rect 9233 1463 9267 1497
rect 9307 1463 9341 1497
rect 9381 1463 9415 1497
rect 9455 1463 9489 1497
rect 9529 1463 9563 1497
rect 9603 1463 9637 1497
rect 9677 1463 9711 1497
rect 9825 1463 9859 1497
rect 9899 1463 9933 1497
rect 9973 1463 10007 1497
rect 10047 1463 10081 1497
rect 10121 1463 10155 1497
rect 10195 1463 10229 1497
rect 10269 1463 10303 1497
rect 10343 1463 10377 1497
rect 10491 1463 10525 1497
rect 10565 1463 10599 1497
rect 10639 1463 10673 1497
rect 10713 1463 10747 1497
rect 10787 1463 10821 1497
rect 10861 1463 10895 1497
rect 10935 1463 10969 1497
rect 11009 1463 11043 1497
rect 11083 1463 11117 1497
rect 11157 1463 11191 1497
rect 11231 1463 11265 1497
rect 11305 1463 11339 1497
rect 11453 1463 11487 1497
rect 11527 1463 11561 1497
rect 11601 1463 11635 1497
rect 11675 1463 11709 1497
rect 11749 1463 11783 1497
rect 11823 1463 11857 1497
rect 11897 1463 11931 1497
rect 11971 1463 12005 1497
rect 12045 1463 12079 1497
rect 12119 1463 12153 1497
rect 12193 1463 12227 1497
rect 12267 1463 12301 1497
rect 12415 1463 12449 1497
rect 12489 1463 12523 1497
rect 12563 1463 12597 1497
rect 12637 1463 12671 1497
rect 12711 1463 12745 1497
rect 12785 1463 12819 1497
rect 12859 1463 12893 1497
rect 12933 1463 12967 1497
rect 13081 1463 13115 1497
rect 13155 1463 13189 1497
rect 13229 1463 13263 1497
rect 13303 1463 13337 1497
rect 13377 1463 13411 1497
rect 13451 1463 13485 1497
rect 13525 1463 13559 1497
rect 13599 1463 13633 1497
rect 13747 1463 13781 1497
rect 13821 1463 13855 1497
rect 13895 1463 13929 1497
rect 13969 1463 14003 1497
rect 14043 1463 14077 1497
rect 14117 1463 14151 1497
rect 14191 1463 14225 1497
rect 14265 1463 14299 1497
rect 14339 1463 14373 1497
rect 14413 1463 14447 1497
rect 14487 1463 14521 1497
rect 14561 1463 14595 1497
rect 14709 1463 14743 1497
rect 14783 1463 14817 1497
rect 14857 1463 14891 1497
rect 14931 1463 14965 1497
rect 15005 1463 15039 1497
rect 15079 1463 15113 1497
rect 15153 1463 15187 1497
rect 15227 1463 15261 1497
rect 15375 1463 15409 1497
rect 15449 1463 15483 1497
rect 15523 1463 15557 1497
rect 15597 1463 15631 1497
rect 15671 1463 15705 1497
rect 15745 1463 15779 1497
rect 15819 1463 15853 1497
rect 15893 1463 15927 1497
rect 16041 1463 16075 1497
rect 16115 1463 16149 1497
rect 16189 1463 16223 1497
rect 16263 1463 16297 1497
rect 16337 1463 16371 1497
rect 16411 1463 16445 1497
rect 16485 1463 16519 1497
rect 16559 1463 16593 1497
rect 16707 1463 16741 1497
rect 16781 1463 16815 1497
rect 16855 1463 16889 1497
rect 16929 1463 16963 1497
rect 17003 1463 17037 1497
rect -17 1389 17 1423
rect -17 1315 17 1349
rect -17 1241 17 1275
rect -17 1167 17 1201
rect -17 1093 17 1127
rect -17 1019 17 1053
rect 649 1389 683 1423
rect 649 1315 683 1349
rect 649 1241 683 1275
rect 649 1167 683 1201
rect 649 1093 683 1127
rect 649 1019 683 1053
rect -17 945 17 979
rect 1611 1389 1645 1423
rect 1611 1315 1645 1349
rect 1611 1241 1645 1275
rect 1611 1167 1645 1201
rect 1611 1093 1645 1127
rect 1611 1019 1645 1053
rect 649 945 683 979
rect -17 871 17 905
rect 2573 1389 2607 1423
rect 2573 1315 2607 1349
rect 2573 1241 2607 1275
rect 2573 1167 2607 1201
rect 2573 1093 2607 1127
rect 2573 1019 2607 1053
rect 1611 945 1645 979
rect 649 871 683 905
rect 3239 1389 3273 1423
rect 3239 1315 3273 1349
rect 3239 1241 3273 1275
rect 3239 1167 3273 1201
rect 3239 1093 3273 1127
rect 3239 1019 3273 1053
rect 2573 945 2607 979
rect 1611 871 1645 905
rect 3905 1389 3939 1423
rect 3905 1315 3939 1349
rect 3905 1241 3939 1275
rect 3905 1167 3939 1201
rect 3905 1093 3939 1127
rect 3905 1019 3939 1053
rect 3239 945 3273 979
rect 2573 871 2607 905
rect 4867 1389 4901 1423
rect 4867 1315 4901 1349
rect 4867 1241 4901 1275
rect 4867 1167 4901 1201
rect 4867 1093 4901 1127
rect 4867 1019 4901 1053
rect 3905 945 3939 979
rect 3239 871 3273 905
rect 5533 1389 5567 1423
rect 5533 1315 5567 1349
rect 5533 1241 5567 1275
rect 5533 1167 5567 1201
rect 5533 1093 5567 1127
rect 5533 1019 5567 1053
rect 4867 945 4901 979
rect 3905 871 3939 905
rect 6495 1389 6529 1423
rect 6495 1315 6529 1349
rect 6495 1241 6529 1275
rect 6495 1167 6529 1201
rect 6495 1093 6529 1127
rect 6495 1019 6529 1053
rect 5533 945 5567 979
rect 4867 871 4901 905
rect 7457 1389 7491 1423
rect 7457 1315 7491 1349
rect 7457 1241 7491 1275
rect 7457 1167 7491 1201
rect 7457 1093 7491 1127
rect 7457 1019 7491 1053
rect 6495 945 6529 979
rect 5533 871 5567 905
rect 8123 1389 8157 1423
rect 8123 1315 8157 1349
rect 8123 1241 8157 1275
rect 8123 1167 8157 1201
rect 8123 1093 8157 1127
rect 8123 1019 8157 1053
rect 7457 945 7491 979
rect 6495 871 6529 905
rect 8789 1389 8823 1423
rect 8789 1315 8823 1349
rect 8789 1241 8823 1275
rect 8789 1167 8823 1201
rect 8789 1093 8823 1127
rect 8789 1019 8823 1053
rect 8123 945 8157 979
rect 7457 871 7491 905
rect 9751 1389 9785 1423
rect 9751 1315 9785 1349
rect 9751 1241 9785 1275
rect 9751 1167 9785 1201
rect 9751 1093 9785 1127
rect 9751 1019 9785 1053
rect 8789 945 8823 979
rect 8123 871 8157 905
rect 10417 1389 10451 1423
rect 10417 1315 10451 1349
rect 10417 1241 10451 1275
rect 10417 1167 10451 1201
rect 10417 1093 10451 1127
rect 10417 1019 10451 1053
rect 9751 945 9785 979
rect 8789 871 8823 905
rect 11379 1389 11413 1423
rect 11379 1315 11413 1349
rect 11379 1241 11413 1275
rect 11379 1167 11413 1201
rect 11379 1093 11413 1127
rect 11379 1019 11413 1053
rect 10417 945 10451 979
rect 9751 871 9785 905
rect 12341 1389 12375 1423
rect 12341 1315 12375 1349
rect 12341 1241 12375 1275
rect 12341 1167 12375 1201
rect 12341 1093 12375 1127
rect 12341 1019 12375 1053
rect 11379 945 11413 979
rect 10417 871 10451 905
rect 13007 1389 13041 1423
rect 13007 1315 13041 1349
rect 13007 1241 13041 1275
rect 13007 1167 13041 1201
rect 13007 1093 13041 1127
rect 13007 1019 13041 1053
rect 12341 945 12375 979
rect 11379 871 11413 905
rect 13673 1389 13707 1423
rect 13673 1315 13707 1349
rect 13673 1241 13707 1275
rect 13673 1167 13707 1201
rect 13673 1093 13707 1127
rect 13673 1019 13707 1053
rect 13007 945 13041 979
rect 12341 871 12375 905
rect 14635 1389 14669 1423
rect 14635 1315 14669 1349
rect 14635 1241 14669 1275
rect 14635 1167 14669 1201
rect 14635 1093 14669 1127
rect 14635 1019 14669 1053
rect 13673 945 13707 979
rect 13007 871 13041 905
rect 15301 1389 15335 1423
rect 15301 1315 15335 1349
rect 15301 1241 15335 1275
rect 15301 1167 15335 1201
rect 15301 1093 15335 1127
rect 15301 1019 15335 1053
rect 14635 945 14669 979
rect 13673 871 13707 905
rect 15967 1389 16001 1423
rect 15967 1315 16001 1349
rect 15967 1241 16001 1275
rect 15967 1167 16001 1201
rect 15967 1093 16001 1127
rect 15967 1019 16001 1053
rect 15301 945 15335 979
rect 14635 871 14669 905
rect 16633 1389 16667 1423
rect 16633 1315 16667 1349
rect 16633 1241 16667 1275
rect 16633 1167 16667 1201
rect 16633 1093 16667 1127
rect 16633 1019 16667 1053
rect 15967 945 16001 979
rect 15301 871 15335 905
rect 17077 1389 17111 1423
rect 17077 1315 17111 1349
rect 17077 1241 17111 1275
rect 17077 1167 17111 1201
rect 17077 1093 17111 1127
rect 17077 1019 17111 1053
rect 16633 945 16667 979
rect 15967 871 16001 905
rect 17077 945 17111 979
rect 16633 871 16667 905
rect 17077 871 17111 905
<< poly >>
rect 187 1404 217 1430
rect 275 1404 305 1430
rect 363 1404 393 1430
rect 451 1404 481 1430
rect 913 1404 943 1430
rect 1001 1404 1031 1430
rect 1089 1404 1119 1430
rect 1177 1404 1207 1430
rect 1265 1404 1295 1430
rect 1353 1404 1383 1430
rect 187 973 217 1004
rect 275 973 305 1004
rect 363 973 393 1004
rect 451 973 481 1004
rect 187 957 305 973
rect 187 943 205 957
rect 195 923 205 943
rect 239 943 305 957
rect 349 957 481 973
rect 239 923 249 943
rect 195 907 249 923
rect 349 923 359 957
rect 393 943 481 957
rect 1875 1404 1905 1430
rect 1963 1404 1993 1430
rect 2051 1404 2081 1430
rect 2139 1404 2169 1430
rect 2227 1404 2257 1430
rect 2315 1404 2345 1430
rect 913 973 943 1004
rect 1001 973 1031 1004
rect 1089 973 1119 1004
rect 1177 973 1207 1004
rect 393 923 403 943
rect 349 907 403 923
rect 861 957 1031 973
rect 861 923 871 957
rect 905 943 1031 957
rect 1083 957 1207 973
rect 905 923 915 943
rect 861 907 915 923
rect 1083 923 1093 957
rect 1127 943 1207 957
rect 1265 973 1295 1004
rect 1353 973 1383 1004
rect 1265 957 1383 973
rect 1265 943 1315 957
rect 1127 923 1137 943
rect 1083 907 1137 923
rect 1305 923 1315 943
rect 1349 943 1383 957
rect 2777 1404 2807 1430
rect 2865 1404 2895 1430
rect 2953 1404 2983 1430
rect 3041 1404 3071 1430
rect 1875 973 1905 1004
rect 1963 973 1993 1004
rect 2051 973 2081 1004
rect 2139 973 2169 1004
rect 1349 923 1359 943
rect 1305 907 1359 923
rect 1823 957 1993 973
rect 1823 923 1833 957
rect 1867 943 1993 957
rect 2045 957 2169 973
rect 1867 923 1877 943
rect 1823 907 1877 923
rect 2045 923 2055 957
rect 2089 943 2169 957
rect 2227 973 2257 1004
rect 2315 973 2345 1004
rect 2227 957 2345 973
rect 2227 943 2277 957
rect 2089 923 2099 943
rect 2045 907 2099 923
rect 2267 923 2277 943
rect 2311 943 2345 957
rect 3443 1404 3473 1430
rect 3531 1404 3561 1430
rect 3619 1404 3649 1430
rect 3707 1404 3737 1430
rect 2311 923 2321 943
rect 2267 907 2321 923
rect 2777 973 2807 1004
rect 2865 973 2895 1004
rect 2953 973 2983 1004
rect 3041 973 3071 1004
rect 2777 957 2895 973
rect 2777 943 2795 957
rect 2785 923 2795 943
rect 2829 943 2895 957
rect 2939 957 3071 973
rect 2829 923 2839 943
rect 2785 907 2839 923
rect 2939 923 2949 957
rect 2983 943 3071 957
rect 4169 1404 4199 1430
rect 4257 1404 4287 1430
rect 4345 1404 4375 1430
rect 4433 1404 4463 1430
rect 4521 1404 4551 1430
rect 4609 1404 4639 1430
rect 2983 923 2993 943
rect 2939 907 2993 923
rect 3443 973 3473 1004
rect 3531 973 3561 1004
rect 3619 973 3649 1004
rect 3707 973 3737 1004
rect 3443 957 3561 973
rect 3443 943 3461 957
rect 3451 923 3461 943
rect 3495 943 3561 957
rect 3605 957 3737 973
rect 3495 923 3505 943
rect 3451 907 3505 923
rect 3605 923 3615 957
rect 3649 943 3737 957
rect 5071 1404 5101 1430
rect 5159 1404 5189 1430
rect 5247 1404 5277 1430
rect 5335 1404 5365 1430
rect 4169 973 4199 1004
rect 4257 973 4287 1004
rect 4345 973 4375 1004
rect 4433 973 4463 1004
rect 3649 923 3659 943
rect 3605 907 3659 923
rect 4117 957 4287 973
rect 4117 923 4127 957
rect 4161 943 4287 957
rect 4339 957 4463 973
rect 4161 923 4171 943
rect 4117 907 4171 923
rect 4339 923 4349 957
rect 4383 943 4463 957
rect 4521 973 4551 1004
rect 4609 973 4639 1004
rect 4521 957 4639 973
rect 4521 943 4571 957
rect 4383 923 4393 943
rect 4339 907 4393 923
rect 4561 923 4571 943
rect 4605 943 4639 957
rect 5797 1404 5827 1430
rect 5885 1404 5915 1430
rect 5973 1404 6003 1430
rect 6061 1404 6091 1430
rect 6149 1404 6179 1430
rect 6237 1404 6267 1430
rect 4605 923 4615 943
rect 4561 907 4615 923
rect 5071 973 5101 1004
rect 5159 973 5189 1004
rect 5247 973 5277 1004
rect 5335 973 5365 1004
rect 5071 957 5189 973
rect 5071 943 5089 957
rect 5079 923 5089 943
rect 5123 943 5189 957
rect 5233 957 5365 973
rect 5123 923 5133 943
rect 5079 907 5133 923
rect 5233 923 5243 957
rect 5277 943 5365 957
rect 6759 1404 6789 1430
rect 6847 1404 6877 1430
rect 6935 1404 6965 1430
rect 7023 1404 7053 1430
rect 7111 1404 7141 1430
rect 7199 1404 7229 1430
rect 5797 973 5827 1004
rect 5885 973 5915 1004
rect 5973 973 6003 1004
rect 6061 973 6091 1004
rect 5277 923 5287 943
rect 5233 907 5287 923
rect 5745 957 5915 973
rect 5745 923 5755 957
rect 5789 943 5915 957
rect 5967 957 6091 973
rect 5789 923 5799 943
rect 5745 907 5799 923
rect 5967 923 5977 957
rect 6011 943 6091 957
rect 6149 973 6179 1004
rect 6237 973 6267 1004
rect 6149 957 6267 973
rect 6149 943 6199 957
rect 6011 923 6021 943
rect 5967 907 6021 923
rect 6189 923 6199 943
rect 6233 943 6267 957
rect 7661 1404 7691 1430
rect 7749 1404 7779 1430
rect 7837 1404 7867 1430
rect 7925 1404 7955 1430
rect 6759 973 6789 1004
rect 6847 973 6877 1004
rect 6935 973 6965 1004
rect 7023 973 7053 1004
rect 6233 923 6243 943
rect 6189 907 6243 923
rect 6707 957 6877 973
rect 6707 923 6717 957
rect 6751 943 6877 957
rect 6929 957 7053 973
rect 6751 923 6761 943
rect 6707 907 6761 923
rect 6929 923 6939 957
rect 6973 943 7053 957
rect 7111 973 7141 1004
rect 7199 973 7229 1004
rect 7111 957 7229 973
rect 7111 943 7161 957
rect 6973 923 6983 943
rect 6929 907 6983 923
rect 7151 923 7161 943
rect 7195 943 7229 957
rect 8327 1404 8357 1430
rect 8415 1404 8445 1430
rect 8503 1404 8533 1430
rect 8591 1404 8621 1430
rect 7195 923 7205 943
rect 7151 907 7205 923
rect 7661 973 7691 1004
rect 7749 973 7779 1004
rect 7837 973 7867 1004
rect 7925 973 7955 1004
rect 7661 957 7779 973
rect 7661 943 7679 957
rect 7669 923 7679 943
rect 7713 943 7779 957
rect 7823 957 7955 973
rect 7713 923 7723 943
rect 7669 907 7723 923
rect 7823 923 7833 957
rect 7867 943 7955 957
rect 9053 1404 9083 1430
rect 9141 1404 9171 1430
rect 9229 1404 9259 1430
rect 9317 1404 9347 1430
rect 9405 1404 9435 1430
rect 9493 1404 9523 1430
rect 7867 923 7877 943
rect 7823 907 7877 923
rect 8327 973 8357 1004
rect 8415 973 8445 1004
rect 8503 973 8533 1004
rect 8591 973 8621 1004
rect 8327 957 8445 973
rect 8327 943 8345 957
rect 8335 923 8345 943
rect 8379 943 8445 957
rect 8489 957 8621 973
rect 8379 923 8389 943
rect 8335 907 8389 923
rect 8489 923 8499 957
rect 8533 943 8621 957
rect 9955 1404 9985 1430
rect 10043 1404 10073 1430
rect 10131 1404 10161 1430
rect 10219 1404 10249 1430
rect 9053 973 9083 1004
rect 9141 973 9171 1004
rect 9229 973 9259 1004
rect 9317 973 9347 1004
rect 8533 923 8543 943
rect 8489 907 8543 923
rect 9001 957 9171 973
rect 9001 923 9011 957
rect 9045 943 9171 957
rect 9223 957 9347 973
rect 9045 923 9055 943
rect 9001 907 9055 923
rect 9223 923 9233 957
rect 9267 943 9347 957
rect 9405 973 9435 1004
rect 9493 973 9523 1004
rect 9405 957 9523 973
rect 9405 943 9455 957
rect 9267 923 9277 943
rect 9223 907 9277 923
rect 9445 923 9455 943
rect 9489 943 9523 957
rect 10681 1404 10711 1430
rect 10769 1404 10799 1430
rect 10857 1404 10887 1430
rect 10945 1404 10975 1430
rect 11033 1404 11063 1430
rect 11121 1404 11151 1430
rect 9489 923 9499 943
rect 9445 907 9499 923
rect 9955 973 9985 1004
rect 10043 973 10073 1004
rect 10131 973 10161 1004
rect 10219 973 10249 1004
rect 9955 957 10073 973
rect 9955 943 9973 957
rect 9963 923 9973 943
rect 10007 943 10073 957
rect 10117 957 10249 973
rect 10007 923 10017 943
rect 9963 907 10017 923
rect 10117 923 10127 957
rect 10161 943 10249 957
rect 11643 1404 11673 1430
rect 11731 1404 11761 1430
rect 11819 1404 11849 1430
rect 11907 1404 11937 1430
rect 11995 1404 12025 1430
rect 12083 1404 12113 1430
rect 10681 973 10711 1004
rect 10769 973 10799 1004
rect 10857 973 10887 1004
rect 10945 973 10975 1004
rect 10161 923 10171 943
rect 10117 907 10171 923
rect 10629 957 10799 973
rect 10629 923 10639 957
rect 10673 943 10799 957
rect 10851 957 10975 973
rect 10673 923 10683 943
rect 10629 907 10683 923
rect 10851 923 10861 957
rect 10895 943 10975 957
rect 11033 973 11063 1004
rect 11121 973 11151 1004
rect 11033 957 11151 973
rect 11033 943 11083 957
rect 10895 923 10905 943
rect 10851 907 10905 923
rect 11073 923 11083 943
rect 11117 943 11151 957
rect 12545 1404 12575 1430
rect 12633 1404 12663 1430
rect 12721 1404 12751 1430
rect 12809 1404 12839 1430
rect 11643 973 11673 1004
rect 11731 973 11761 1004
rect 11819 973 11849 1004
rect 11907 973 11937 1004
rect 11117 923 11127 943
rect 11073 907 11127 923
rect 11591 957 11761 973
rect 11591 923 11601 957
rect 11635 943 11761 957
rect 11813 957 11937 973
rect 11635 923 11645 943
rect 11591 907 11645 923
rect 11813 923 11823 957
rect 11857 943 11937 957
rect 11995 973 12025 1004
rect 12083 973 12113 1004
rect 11995 957 12113 973
rect 11995 943 12045 957
rect 11857 923 11867 943
rect 11813 907 11867 923
rect 12035 923 12045 943
rect 12079 943 12113 957
rect 13211 1404 13241 1430
rect 13299 1404 13329 1430
rect 13387 1404 13417 1430
rect 13475 1404 13505 1430
rect 12079 923 12089 943
rect 12035 907 12089 923
rect 12545 973 12575 1004
rect 12633 973 12663 1004
rect 12721 973 12751 1004
rect 12809 973 12839 1004
rect 12545 957 12663 973
rect 12545 943 12563 957
rect 12553 923 12563 943
rect 12597 943 12663 957
rect 12707 957 12839 973
rect 12597 923 12607 943
rect 12553 907 12607 923
rect 12707 923 12717 957
rect 12751 943 12839 957
rect 13937 1404 13967 1430
rect 14025 1404 14055 1430
rect 14113 1404 14143 1430
rect 14201 1404 14231 1430
rect 14289 1404 14319 1430
rect 14377 1404 14407 1430
rect 12751 923 12761 943
rect 12707 907 12761 923
rect 13211 973 13241 1004
rect 13299 973 13329 1004
rect 13387 973 13417 1004
rect 13475 973 13505 1004
rect 13211 957 13329 973
rect 13211 943 13229 957
rect 13219 923 13229 943
rect 13263 943 13329 957
rect 13373 957 13505 973
rect 13263 923 13273 943
rect 13219 907 13273 923
rect 13373 923 13383 957
rect 13417 943 13505 957
rect 14839 1405 14869 1431
rect 14927 1405 14957 1431
rect 15015 1405 15045 1431
rect 15103 1405 15133 1431
rect 13937 973 13967 1004
rect 14025 973 14055 1004
rect 14113 973 14143 1004
rect 14201 973 14231 1004
rect 13417 923 13427 943
rect 13373 907 13427 923
rect 13885 957 14055 973
rect 13885 923 13895 957
rect 13929 943 14055 957
rect 14107 957 14231 973
rect 13929 923 13939 943
rect 13885 907 13939 923
rect 14107 923 14117 957
rect 14151 943 14231 957
rect 14289 973 14319 1004
rect 14377 973 14407 1004
rect 14289 957 14407 973
rect 14289 943 14339 957
rect 14151 923 14161 943
rect 14107 907 14161 923
rect 14329 923 14339 943
rect 14373 943 14407 957
rect 15503 1405 15533 1431
rect 15591 1405 15621 1431
rect 15679 1405 15709 1431
rect 15767 1405 15797 1431
rect 14839 974 14869 1005
rect 14927 974 14957 1005
rect 15015 974 15045 1005
rect 15103 974 15133 1005
rect 14373 923 14383 943
rect 14329 907 14383 923
rect 14773 958 14957 974
rect 14773 924 14783 958
rect 14817 944 14957 958
rect 15003 958 15133 974
rect 14817 924 14827 944
rect 14773 908 14827 924
rect 15003 924 15013 958
rect 15047 944 15133 958
rect 16171 1405 16201 1431
rect 16259 1405 16289 1431
rect 16347 1405 16377 1431
rect 16435 1405 16465 1431
rect 15047 924 15057 944
rect 15003 908 15057 924
rect 15503 974 15533 1005
rect 15591 974 15621 1005
rect 15503 958 15621 974
rect 15503 944 15523 958
rect 15513 924 15523 944
rect 15557 944 15621 958
rect 15679 974 15709 1005
rect 15767 974 15797 1005
rect 16814 1404 16844 1430
rect 16902 1404 16932 1430
rect 15679 958 15863 974
rect 15679 944 15819 958
rect 15557 924 15567 944
rect 15513 908 15567 924
rect 15809 924 15819 944
rect 15853 924 15863 958
rect 15809 908 15863 924
rect 16171 974 16201 1005
rect 16259 974 16289 1005
rect 16347 974 16377 1005
rect 16435 974 16465 1005
rect 16105 958 16289 974
rect 16105 924 16115 958
rect 16149 944 16289 958
rect 16331 958 16465 974
rect 16149 924 16159 944
rect 16105 908 16159 924
rect 16331 924 16341 958
rect 16375 944 16465 958
rect 16814 973 16844 1004
rect 16902 973 16932 1004
rect 16375 924 16385 944
rect 16331 908 16385 924
rect 16771 957 16932 973
rect 16771 923 16781 957
rect 16815 943 16932 957
rect 16815 923 16825 943
rect 16771 907 16825 923
rect 195 433 249 449
rect 195 413 205 433
rect 168 399 205 413
rect 239 399 249 433
rect 168 383 249 399
rect 343 433 397 449
rect 343 399 353 433
rect 387 399 397 433
rect 343 383 397 399
rect 861 433 915 449
rect 861 413 871 433
rect 168 349 198 383
rect 362 349 392 383
rect 813 399 871 413
rect 905 399 915 433
rect 813 383 915 399
rect 1083 433 1137 449
rect 1083 399 1093 433
rect 1127 413 1137 433
rect 1305 433 1359 449
rect 1127 399 1143 413
rect 1083 383 1143 399
rect 1305 399 1315 433
rect 1349 399 1359 433
rect 1305 383 1359 399
rect 1823 433 1877 449
rect 1823 413 1833 433
rect 813 351 843 383
rect 1113 351 1143 383
rect 1315 351 1345 383
rect 1775 399 1833 413
rect 1867 399 1877 433
rect 1775 383 1877 399
rect 2045 433 2099 449
rect 2045 399 2055 433
rect 2089 413 2099 433
rect 2267 433 2321 449
rect 2089 399 2105 413
rect 2045 383 2105 399
rect 2267 399 2277 433
rect 2311 399 2321 433
rect 2267 383 2321 399
rect 2785 433 2839 449
rect 2785 413 2795 433
rect 1775 351 1805 383
rect 2075 351 2105 383
rect 2277 351 2307 383
rect 2758 399 2795 413
rect 2829 399 2839 433
rect 2758 383 2839 399
rect 2933 433 2987 449
rect 2933 399 2943 433
rect 2977 399 2987 433
rect 2933 383 2987 399
rect 3451 433 3505 449
rect 3451 413 3461 433
rect 2758 349 2788 383
rect 2952 349 2982 383
rect 3424 399 3461 413
rect 3495 399 3505 433
rect 3424 383 3505 399
rect 3599 433 3653 449
rect 3599 399 3609 433
rect 3643 399 3653 433
rect 3599 383 3653 399
rect 4117 433 4171 449
rect 4117 413 4127 433
rect 3424 349 3454 383
rect 3618 349 3648 383
rect 4069 399 4127 413
rect 4161 399 4171 433
rect 4069 383 4171 399
rect 4339 433 4393 449
rect 4339 399 4349 433
rect 4383 413 4393 433
rect 4561 433 4615 449
rect 4383 399 4399 413
rect 4339 383 4399 399
rect 4561 399 4571 433
rect 4605 399 4615 433
rect 4561 383 4615 399
rect 5079 433 5133 449
rect 5079 413 5089 433
rect 4069 351 4099 383
rect 4369 351 4399 383
rect 4571 351 4601 383
rect 5052 399 5089 413
rect 5123 399 5133 433
rect 5052 383 5133 399
rect 5227 433 5281 449
rect 5227 399 5237 433
rect 5271 399 5281 433
rect 5227 383 5281 399
rect 5745 433 5799 449
rect 5745 413 5755 433
rect 5052 349 5082 383
rect 5246 349 5276 383
rect 5697 399 5755 413
rect 5789 399 5799 433
rect 5697 383 5799 399
rect 5967 433 6021 449
rect 5967 399 5977 433
rect 6011 413 6021 433
rect 6189 433 6243 449
rect 6011 399 6027 413
rect 5967 383 6027 399
rect 6189 399 6199 433
rect 6233 399 6243 433
rect 6189 383 6243 399
rect 6707 433 6761 449
rect 6707 413 6717 433
rect 5697 351 5727 383
rect 5997 351 6027 383
rect 6199 351 6229 383
rect 6659 399 6717 413
rect 6751 399 6761 433
rect 6659 383 6761 399
rect 6929 433 6983 449
rect 6929 399 6939 433
rect 6973 413 6983 433
rect 7151 433 7205 449
rect 6973 399 6989 413
rect 6929 383 6989 399
rect 7151 399 7161 433
rect 7195 399 7205 433
rect 7151 383 7205 399
rect 7669 433 7723 449
rect 7669 413 7679 433
rect 6659 351 6689 383
rect 6959 351 6989 383
rect 7161 351 7191 383
rect 7642 399 7679 413
rect 7713 399 7723 433
rect 7642 383 7723 399
rect 7817 433 7871 449
rect 7817 399 7827 433
rect 7861 399 7871 433
rect 7817 383 7871 399
rect 8335 433 8389 449
rect 8335 413 8345 433
rect 7642 349 7672 383
rect 7836 349 7866 383
rect 8308 399 8345 413
rect 8379 399 8389 433
rect 8308 383 8389 399
rect 8483 433 8537 449
rect 8483 399 8493 433
rect 8527 399 8537 433
rect 8483 383 8537 399
rect 9001 433 9055 449
rect 9001 413 9011 433
rect 8308 349 8338 383
rect 8502 349 8532 383
rect 8953 399 9011 413
rect 9045 399 9055 433
rect 8953 383 9055 399
rect 9223 433 9277 449
rect 9223 399 9233 433
rect 9267 413 9277 433
rect 9445 433 9499 449
rect 9267 399 9283 413
rect 9223 383 9283 399
rect 9445 399 9455 433
rect 9489 399 9499 433
rect 9445 383 9499 399
rect 9963 433 10017 449
rect 9963 413 9973 433
rect 8953 351 8983 383
rect 9253 351 9283 383
rect 9455 351 9485 383
rect 9936 399 9973 413
rect 10007 399 10017 433
rect 9936 383 10017 399
rect 10111 433 10165 449
rect 10111 399 10121 433
rect 10155 399 10165 433
rect 10111 383 10165 399
rect 10629 433 10683 449
rect 10629 413 10639 433
rect 9936 349 9966 383
rect 10130 349 10160 383
rect 10581 399 10639 413
rect 10673 399 10683 433
rect 10581 383 10683 399
rect 10851 433 10905 449
rect 10851 399 10861 433
rect 10895 413 10905 433
rect 11073 433 11127 449
rect 10895 399 10911 413
rect 10851 383 10911 399
rect 11073 399 11083 433
rect 11117 399 11127 433
rect 11073 383 11127 399
rect 11591 433 11645 449
rect 11591 413 11601 433
rect 10581 351 10611 383
rect 10881 351 10911 383
rect 11083 351 11113 383
rect 11543 399 11601 413
rect 11635 399 11645 433
rect 11543 383 11645 399
rect 11813 433 11867 449
rect 11813 399 11823 433
rect 11857 413 11867 433
rect 12035 433 12089 449
rect 11857 399 11873 413
rect 11813 383 11873 399
rect 12035 399 12045 433
rect 12079 399 12089 433
rect 12035 383 12089 399
rect 12553 433 12607 449
rect 12553 413 12563 433
rect 11543 351 11573 383
rect 11843 351 11873 383
rect 12045 351 12075 383
rect 12526 399 12563 413
rect 12597 399 12607 433
rect 12526 383 12607 399
rect 12701 433 12755 449
rect 12701 399 12711 433
rect 12745 399 12755 433
rect 12701 383 12755 399
rect 13219 433 13273 449
rect 13219 413 13229 433
rect 12526 349 12556 383
rect 12720 349 12750 383
rect 13192 399 13229 413
rect 13263 399 13273 433
rect 13192 383 13273 399
rect 13367 433 13421 449
rect 13367 399 13377 433
rect 13411 399 13421 433
rect 13367 383 13421 399
rect 13885 433 13939 449
rect 13885 413 13895 433
rect 13192 349 13222 383
rect 13386 349 13416 383
rect 13837 399 13895 413
rect 13929 399 13939 433
rect 13837 383 13939 399
rect 14107 433 14161 449
rect 14107 399 14117 433
rect 14151 413 14161 433
rect 14329 433 14383 449
rect 14151 399 14167 413
rect 14107 383 14167 399
rect 14329 399 14339 433
rect 14373 399 14383 433
rect 14329 383 14383 399
rect 13837 351 13867 383
rect 14137 351 14167 383
rect 14339 351 14369 383
rect 14773 433 14827 449
rect 14773 399 14783 433
rect 14817 413 14827 433
rect 14995 433 15049 449
rect 14817 399 14850 413
rect 14773 383 14850 399
rect 14995 399 15005 433
rect 15039 399 15049 433
rect 14995 383 15049 399
rect 15513 433 15567 449
rect 15513 413 15523 433
rect 14820 349 14850 383
rect 15014 349 15044 383
rect 15486 399 15523 413
rect 15557 399 15567 433
rect 15809 433 15863 449
rect 15809 413 15819 433
rect 15486 383 15567 399
rect 15786 399 15819 413
rect 15853 399 15863 433
rect 15786 383 15863 399
rect 15486 349 15516 383
rect 15786 349 15816 383
rect 16105 433 16159 449
rect 16105 399 16115 433
rect 16149 413 16159 433
rect 16327 433 16381 449
rect 16149 399 16182 413
rect 16105 383 16182 399
rect 16327 399 16337 433
rect 16371 399 16381 433
rect 16327 383 16381 399
rect 16152 349 16182 383
rect 16346 349 16376 383
rect 16771 434 16825 450
rect 16771 400 16781 434
rect 16815 413 16825 434
rect 16815 400 16835 413
rect 16771 384 16835 400
rect 16805 350 16835 384
<< polycont >>
rect 205 923 239 957
rect 359 923 393 957
rect 871 923 905 957
rect 1093 923 1127 957
rect 1315 923 1349 957
rect 1833 923 1867 957
rect 2055 923 2089 957
rect 2277 923 2311 957
rect 2795 923 2829 957
rect 2949 923 2983 957
rect 3461 923 3495 957
rect 3615 923 3649 957
rect 4127 923 4161 957
rect 4349 923 4383 957
rect 4571 923 4605 957
rect 5089 923 5123 957
rect 5243 923 5277 957
rect 5755 923 5789 957
rect 5977 923 6011 957
rect 6199 923 6233 957
rect 6717 923 6751 957
rect 6939 923 6973 957
rect 7161 923 7195 957
rect 7679 923 7713 957
rect 7833 923 7867 957
rect 8345 923 8379 957
rect 8499 923 8533 957
rect 9011 923 9045 957
rect 9233 923 9267 957
rect 9455 923 9489 957
rect 9973 923 10007 957
rect 10127 923 10161 957
rect 10639 923 10673 957
rect 10861 923 10895 957
rect 11083 923 11117 957
rect 11601 923 11635 957
rect 11823 923 11857 957
rect 12045 923 12079 957
rect 12563 923 12597 957
rect 12717 923 12751 957
rect 13229 923 13263 957
rect 13383 923 13417 957
rect 13895 923 13929 957
rect 14117 923 14151 957
rect 14339 923 14373 957
rect 14783 924 14817 958
rect 15013 924 15047 958
rect 15523 924 15557 958
rect 15819 924 15853 958
rect 16115 924 16149 958
rect 16341 924 16375 958
rect 16781 923 16815 957
rect 205 399 239 433
rect 353 399 387 433
rect 871 399 905 433
rect 1093 399 1127 433
rect 1315 399 1349 433
rect 1833 399 1867 433
rect 2055 399 2089 433
rect 2277 399 2311 433
rect 2795 399 2829 433
rect 2943 399 2977 433
rect 3461 399 3495 433
rect 3609 399 3643 433
rect 4127 399 4161 433
rect 4349 399 4383 433
rect 4571 399 4605 433
rect 5089 399 5123 433
rect 5237 399 5271 433
rect 5755 399 5789 433
rect 5977 399 6011 433
rect 6199 399 6233 433
rect 6717 399 6751 433
rect 6939 399 6973 433
rect 7161 399 7195 433
rect 7679 399 7713 433
rect 7827 399 7861 433
rect 8345 399 8379 433
rect 8493 399 8527 433
rect 9011 399 9045 433
rect 9233 399 9267 433
rect 9455 399 9489 433
rect 9973 399 10007 433
rect 10121 399 10155 433
rect 10639 399 10673 433
rect 10861 399 10895 433
rect 11083 399 11117 433
rect 11601 399 11635 433
rect 11823 399 11857 433
rect 12045 399 12079 433
rect 12563 399 12597 433
rect 12711 399 12745 433
rect 13229 399 13263 433
rect 13377 399 13411 433
rect 13895 399 13929 433
rect 14117 399 14151 433
rect 14339 399 14373 433
rect 14783 399 14817 433
rect 15005 399 15039 433
rect 15523 399 15557 433
rect 15819 399 15853 433
rect 16115 399 16149 433
rect 16337 399 16371 433
rect 16781 400 16815 434
<< locali >>
rect -34 1497 17128 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5163 1497
rect 5197 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5755 1497
rect 5789 1463 5829 1497
rect 5863 1463 5903 1497
rect 5937 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6125 1497
rect 6159 1463 6199 1497
rect 6233 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6569 1497
rect 6603 1463 6643 1497
rect 6677 1463 6717 1497
rect 6751 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7087 1497
rect 7121 1463 7161 1497
rect 7195 1463 7235 1497
rect 7269 1463 7309 1497
rect 7343 1463 7383 1497
rect 7417 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7679 1497
rect 7713 1463 7753 1497
rect 7787 1463 7827 1497
rect 7861 1463 7901 1497
rect 7935 1463 7975 1497
rect 8009 1463 8049 1497
rect 8083 1463 8197 1497
rect 8231 1463 8271 1497
rect 8305 1463 8345 1497
rect 8379 1463 8419 1497
rect 8453 1463 8493 1497
rect 8527 1463 8567 1497
rect 8601 1463 8641 1497
rect 8675 1463 8715 1497
rect 8749 1463 8863 1497
rect 8897 1463 8937 1497
rect 8971 1463 9011 1497
rect 9045 1463 9085 1497
rect 9119 1463 9159 1497
rect 9193 1463 9233 1497
rect 9267 1463 9307 1497
rect 9341 1463 9381 1497
rect 9415 1463 9455 1497
rect 9489 1463 9529 1497
rect 9563 1463 9603 1497
rect 9637 1463 9677 1497
rect 9711 1463 9825 1497
rect 9859 1463 9899 1497
rect 9933 1463 9973 1497
rect 10007 1463 10047 1497
rect 10081 1463 10121 1497
rect 10155 1463 10195 1497
rect 10229 1463 10269 1497
rect 10303 1463 10343 1497
rect 10377 1463 10491 1497
rect 10525 1463 10565 1497
rect 10599 1463 10639 1497
rect 10673 1463 10713 1497
rect 10747 1463 10787 1497
rect 10821 1463 10861 1497
rect 10895 1463 10935 1497
rect 10969 1463 11009 1497
rect 11043 1463 11083 1497
rect 11117 1463 11157 1497
rect 11191 1463 11231 1497
rect 11265 1463 11305 1497
rect 11339 1463 11453 1497
rect 11487 1463 11527 1497
rect 11561 1463 11601 1497
rect 11635 1463 11675 1497
rect 11709 1463 11749 1497
rect 11783 1463 11823 1497
rect 11857 1463 11897 1497
rect 11931 1463 11971 1497
rect 12005 1463 12045 1497
rect 12079 1463 12119 1497
rect 12153 1463 12193 1497
rect 12227 1463 12267 1497
rect 12301 1463 12415 1497
rect 12449 1463 12489 1497
rect 12523 1463 12563 1497
rect 12597 1463 12637 1497
rect 12671 1463 12711 1497
rect 12745 1463 12785 1497
rect 12819 1463 12859 1497
rect 12893 1463 12933 1497
rect 12967 1463 13081 1497
rect 13115 1463 13155 1497
rect 13189 1463 13229 1497
rect 13263 1463 13303 1497
rect 13337 1463 13377 1497
rect 13411 1463 13451 1497
rect 13485 1463 13525 1497
rect 13559 1463 13599 1497
rect 13633 1463 13747 1497
rect 13781 1463 13821 1497
rect 13855 1463 13895 1497
rect 13929 1463 13969 1497
rect 14003 1463 14043 1497
rect 14077 1463 14117 1497
rect 14151 1463 14191 1497
rect 14225 1463 14265 1497
rect 14299 1463 14339 1497
rect 14373 1463 14413 1497
rect 14447 1463 14487 1497
rect 14521 1463 14561 1497
rect 14595 1463 14709 1497
rect 14743 1463 14783 1497
rect 14817 1463 14857 1497
rect 14891 1463 14931 1497
rect 14965 1463 15005 1497
rect 15039 1463 15079 1497
rect 15113 1463 15153 1497
rect 15187 1463 15227 1497
rect 15261 1463 15375 1497
rect 15409 1463 15449 1497
rect 15483 1463 15523 1497
rect 15557 1463 15597 1497
rect 15631 1463 15671 1497
rect 15705 1463 15745 1497
rect 15779 1463 15819 1497
rect 15853 1463 15893 1497
rect 15927 1463 16041 1497
rect 16075 1463 16115 1497
rect 16149 1463 16189 1497
rect 16223 1463 16263 1497
rect 16297 1463 16337 1497
rect 16371 1463 16411 1497
rect 16445 1463 16485 1497
rect 16519 1463 16559 1497
rect 16593 1463 16707 1497
rect 16741 1463 16781 1497
rect 16815 1463 16855 1497
rect 16889 1463 16929 1497
rect 16963 1463 17003 1497
rect 17037 1463 17128 1497
rect -34 1446 17128 1463
rect -34 1423 34 1446
rect -34 1389 -17 1423
rect 17 1389 34 1423
rect -34 1349 34 1389
rect -34 1315 -17 1349
rect 17 1315 34 1349
rect -34 1275 34 1315
rect -34 1241 -17 1275
rect 17 1241 34 1275
rect -34 1201 34 1241
rect -34 1167 -17 1201
rect 17 1167 34 1201
rect -34 1127 34 1167
rect -34 1093 -17 1127
rect 17 1093 34 1127
rect -34 1053 34 1093
rect -34 1019 -17 1053
rect 17 1019 34 1053
rect 141 1366 175 1446
rect 141 1298 175 1332
rect 141 1230 175 1264
rect 141 1162 175 1196
rect 141 1093 175 1128
rect 141 1027 175 1059
rect 229 1366 263 1404
rect 229 1298 263 1332
rect 229 1230 263 1264
rect 229 1162 263 1196
rect 229 1093 263 1128
rect 317 1366 351 1446
rect 317 1298 351 1332
rect 317 1230 351 1264
rect 317 1162 351 1196
rect 317 1111 351 1128
rect 405 1366 439 1404
rect 405 1298 439 1332
rect 405 1230 439 1264
rect 405 1162 439 1196
rect 229 1057 263 1059
rect 405 1093 439 1128
rect 493 1366 527 1446
rect 493 1298 527 1332
rect 493 1230 527 1264
rect 493 1162 527 1196
rect 493 1111 527 1128
rect 632 1423 700 1446
rect 632 1389 649 1423
rect 683 1389 700 1423
rect 632 1349 700 1389
rect 632 1315 649 1349
rect 683 1315 700 1349
rect 632 1275 700 1315
rect 632 1241 649 1275
rect 683 1241 700 1275
rect 632 1201 700 1241
rect 632 1167 649 1201
rect 683 1167 700 1201
rect 632 1127 700 1167
rect 405 1057 439 1059
rect 632 1093 649 1127
rect 683 1093 700 1127
rect 229 1023 535 1057
rect -34 979 34 1019
rect -34 945 -17 979
rect 17 945 34 979
rect -34 905 34 945
rect -34 871 -17 905
rect 17 871 34 905
rect -34 822 34 871
rect 205 957 239 973
rect 359 957 393 973
rect 205 609 239 923
rect -34 461 34 544
rect -34 427 -17 461
rect 17 427 34 461
rect -34 387 34 427
rect -34 353 -17 387
rect 17 353 34 387
rect 205 433 239 575
rect 205 383 239 399
rect 353 923 359 942
rect 353 907 393 923
rect 353 831 387 907
rect 353 433 387 797
rect 353 383 387 399
rect 501 535 535 1023
rect 632 1053 700 1093
rect 632 1019 649 1053
rect 683 1019 700 1053
rect 867 1366 901 1446
rect 867 1298 901 1332
rect 867 1230 901 1264
rect 867 1162 901 1196
rect 867 1093 901 1128
rect 867 1043 901 1059
rect 955 1366 989 1404
rect 955 1298 989 1332
rect 955 1230 989 1264
rect 955 1162 989 1196
rect 955 1093 989 1128
rect 1043 1366 1077 1446
rect 1043 1298 1077 1332
rect 1043 1230 1077 1264
rect 1043 1162 1077 1196
rect 1043 1111 1077 1128
rect 1131 1366 1165 1404
rect 1131 1298 1165 1332
rect 1131 1230 1165 1264
rect 1131 1162 1165 1196
rect 955 1048 989 1059
rect 1131 1093 1165 1128
rect 1219 1366 1253 1446
rect 1219 1298 1253 1332
rect 1219 1230 1253 1264
rect 1219 1162 1253 1196
rect 1219 1111 1253 1128
rect 1307 1366 1341 1404
rect 1307 1298 1341 1332
rect 1307 1230 1341 1264
rect 1307 1162 1341 1196
rect 1131 1048 1165 1059
rect 1307 1093 1341 1128
rect 1395 1366 1429 1446
rect 1395 1298 1429 1332
rect 1395 1230 1429 1264
rect 1395 1162 1429 1196
rect 1395 1111 1429 1128
rect 1594 1423 1662 1446
rect 1594 1389 1611 1423
rect 1645 1389 1662 1423
rect 1594 1349 1662 1389
rect 1594 1315 1611 1349
rect 1645 1315 1662 1349
rect 1594 1275 1662 1315
rect 1594 1241 1611 1275
rect 1645 1241 1662 1275
rect 1594 1201 1662 1241
rect 1594 1167 1611 1201
rect 1645 1167 1662 1201
rect 1594 1127 1662 1167
rect 1307 1048 1341 1059
rect 1594 1093 1611 1127
rect 1645 1093 1662 1127
rect 1594 1053 1662 1093
rect 632 979 700 1019
rect 955 1014 1497 1048
rect 632 945 649 979
rect 683 945 700 979
rect 632 905 700 945
rect 632 871 649 905
rect 683 871 700 905
rect 632 822 700 871
rect 871 957 905 973
rect -34 313 34 353
rect -34 279 -17 313
rect 17 279 34 313
rect -34 239 34 279
rect -34 205 -17 239
rect 17 205 34 239
rect -34 165 34 205
rect -34 131 -17 165
rect 17 131 34 165
rect -34 91 34 131
rect -34 57 -17 91
rect 17 57 34 91
rect 122 333 156 349
rect 316 333 350 349
rect 501 348 535 501
rect 156 299 219 333
rect 253 299 316 333
rect 122 261 156 299
rect 122 193 156 227
rect 316 261 350 299
rect 122 123 156 159
rect 122 73 156 89
rect 219 208 253 224
rect -34 34 34 57
rect 219 34 253 174
rect 316 193 350 227
rect 413 314 535 348
rect 632 461 700 544
rect 632 427 649 461
rect 683 427 700 461
rect 632 387 700 427
rect 632 353 649 387
rect 683 353 700 387
rect 871 534 905 923
rect 871 433 905 500
rect 871 383 905 399
rect 1093 957 1127 973
rect 1093 905 1127 923
rect 1093 433 1127 871
rect 1093 383 1127 399
rect 1315 957 1349 973
rect 1315 757 1349 923
rect 1463 847 1497 1014
rect 1462 831 1497 847
rect 1496 797 1497 831
rect 1594 1019 1611 1053
rect 1645 1019 1662 1053
rect 1829 1366 1863 1446
rect 1829 1298 1863 1332
rect 1829 1230 1863 1264
rect 1829 1162 1863 1196
rect 1829 1093 1863 1128
rect 1829 1043 1863 1059
rect 1917 1366 1951 1404
rect 1917 1298 1951 1332
rect 1917 1230 1951 1264
rect 1917 1162 1951 1196
rect 1917 1093 1951 1128
rect 2005 1366 2039 1446
rect 2005 1298 2039 1332
rect 2005 1230 2039 1264
rect 2005 1162 2039 1196
rect 2005 1111 2039 1128
rect 2093 1366 2127 1404
rect 2093 1298 2127 1332
rect 2093 1230 2127 1264
rect 2093 1162 2127 1196
rect 1917 1048 1951 1059
rect 2093 1093 2127 1128
rect 2181 1366 2215 1446
rect 2181 1298 2215 1332
rect 2181 1230 2215 1264
rect 2181 1162 2215 1196
rect 2181 1111 2215 1128
rect 2269 1366 2303 1404
rect 2269 1298 2303 1332
rect 2269 1230 2303 1264
rect 2269 1162 2303 1196
rect 2093 1048 2127 1059
rect 2269 1093 2303 1128
rect 2357 1366 2391 1446
rect 2357 1298 2391 1332
rect 2357 1230 2391 1264
rect 2357 1162 2391 1196
rect 2357 1111 2391 1128
rect 2556 1423 2624 1446
rect 2556 1389 2573 1423
rect 2607 1389 2624 1423
rect 2556 1349 2624 1389
rect 2556 1315 2573 1349
rect 2607 1315 2624 1349
rect 2556 1275 2624 1315
rect 2556 1241 2573 1275
rect 2607 1241 2624 1275
rect 2556 1201 2624 1241
rect 2556 1167 2573 1201
rect 2607 1167 2624 1201
rect 2556 1127 2624 1167
rect 2269 1048 2303 1059
rect 2556 1093 2573 1127
rect 2607 1093 2624 1127
rect 2556 1053 2624 1093
rect 1594 979 1662 1019
rect 1917 1014 2459 1048
rect 1594 945 1611 979
rect 1645 945 1662 979
rect 1594 905 1662 945
rect 1594 871 1611 905
rect 1645 871 1662 905
rect 1594 822 1662 871
rect 1833 957 1867 973
rect 1462 781 1497 797
rect 1315 433 1349 723
rect 1315 383 1349 399
rect 413 217 447 314
rect 632 313 700 353
rect 632 279 649 313
rect 683 279 700 313
rect 413 167 447 183
rect 510 261 544 277
rect 510 193 544 227
rect 316 123 350 159
rect 510 123 544 159
rect 350 89 413 123
rect 447 89 510 123
rect 316 73 350 89
rect 510 73 544 89
rect 632 239 700 279
rect 632 205 649 239
rect 683 205 700 239
rect 632 165 700 205
rect 632 131 649 165
rect 683 131 700 165
rect 632 91 700 131
rect 632 57 649 91
rect 683 57 700 91
rect 767 335 801 351
rect 961 335 995 351
rect 1155 335 1189 351
rect 801 301 864 335
rect 898 301 961 335
rect 995 301 1058 335
rect 1092 301 1155 335
rect 767 263 801 301
rect 767 195 801 229
rect 961 263 995 301
rect 1155 285 1189 301
rect 1269 335 1303 351
rect 1463 350 1497 781
rect 1269 263 1303 301
rect 767 125 801 161
rect 767 75 801 91
rect 864 210 898 226
rect 632 34 700 57
rect 864 34 898 176
rect 961 195 995 229
rect 1059 216 1093 232
rect 1269 216 1303 229
rect 1093 195 1303 216
rect 1093 182 1269 195
rect 1059 166 1093 182
rect 961 125 995 161
rect 1366 316 1497 350
rect 1594 461 1662 544
rect 1594 427 1611 461
rect 1645 427 1662 461
rect 1594 387 1662 427
rect 1594 353 1611 387
rect 1645 353 1662 387
rect 1833 535 1867 923
rect 1833 433 1867 501
rect 1833 383 1867 399
rect 2055 957 2089 973
rect 2055 461 2089 923
rect 2055 383 2089 399
rect 2277 957 2311 973
rect 2277 757 2311 923
rect 2277 433 2311 723
rect 2277 383 2311 399
rect 2425 535 2459 1014
rect 2556 1019 2573 1053
rect 2607 1019 2624 1053
rect 2731 1366 2765 1446
rect 2731 1298 2765 1332
rect 2731 1230 2765 1264
rect 2731 1162 2765 1196
rect 2731 1093 2765 1128
rect 2731 1027 2765 1059
rect 2819 1366 2853 1404
rect 2819 1298 2853 1332
rect 2819 1230 2853 1264
rect 2819 1162 2853 1196
rect 2819 1093 2853 1128
rect 2907 1366 2941 1446
rect 2907 1298 2941 1332
rect 2907 1230 2941 1264
rect 2907 1162 2941 1196
rect 2907 1111 2941 1128
rect 2995 1366 3029 1404
rect 2995 1298 3029 1332
rect 2995 1230 3029 1264
rect 2995 1162 3029 1196
rect 2819 1057 2853 1059
rect 2995 1093 3029 1128
rect 3083 1366 3117 1446
rect 3083 1298 3117 1332
rect 3083 1230 3117 1264
rect 3083 1162 3117 1196
rect 3083 1111 3117 1128
rect 3222 1423 3290 1446
rect 3222 1389 3239 1423
rect 3273 1389 3290 1423
rect 3222 1349 3290 1389
rect 3222 1315 3239 1349
rect 3273 1315 3290 1349
rect 3222 1275 3290 1315
rect 3222 1241 3239 1275
rect 3273 1241 3290 1275
rect 3222 1201 3290 1241
rect 3222 1167 3239 1201
rect 3273 1167 3290 1201
rect 3222 1127 3290 1167
rect 2995 1057 3029 1059
rect 3222 1093 3239 1127
rect 3273 1093 3290 1127
rect 2819 1023 3125 1057
rect 2556 979 2624 1019
rect 2556 945 2573 979
rect 2607 945 2624 979
rect 2556 905 2624 945
rect 2556 871 2573 905
rect 2607 871 2624 905
rect 2556 822 2624 871
rect 2795 957 2829 973
rect 2949 957 2983 973
rect 1366 219 1400 316
rect 1594 313 1662 353
rect 1594 279 1611 313
rect 1645 279 1662 313
rect 1366 169 1400 185
rect 1463 263 1497 279
rect 1463 195 1497 229
rect 1155 125 1189 141
rect 995 91 1058 125
rect 1092 91 1155 125
rect 961 75 995 91
rect 1155 75 1189 91
rect 1269 125 1303 161
rect 1463 125 1497 161
rect 1303 91 1366 125
rect 1400 91 1463 125
rect 1269 75 1303 91
rect 1463 75 1497 91
rect 1594 239 1662 279
rect 1594 205 1611 239
rect 1645 205 1662 239
rect 1594 165 1662 205
rect 1594 131 1611 165
rect 1645 131 1662 165
rect 1594 91 1662 131
rect 1594 57 1611 91
rect 1645 57 1662 91
rect 1729 335 1763 351
rect 1923 335 1957 351
rect 2117 335 2151 351
rect 1763 301 1826 335
rect 1860 301 1923 335
rect 1957 301 2020 335
rect 2054 301 2117 335
rect 1729 263 1763 301
rect 1729 195 1763 229
rect 1923 263 1957 301
rect 2117 285 2151 301
rect 2231 335 2265 351
rect 2425 350 2459 501
rect 2231 263 2265 301
rect 1729 125 1763 161
rect 1729 75 1763 91
rect 1826 210 1860 226
rect 1594 34 1662 57
rect 1826 34 1860 176
rect 1923 195 1957 229
rect 2021 216 2055 232
rect 2231 216 2265 229
rect 2055 195 2265 216
rect 2055 182 2231 195
rect 2021 166 2055 182
rect 1923 125 1957 161
rect 2328 316 2459 350
rect 2556 461 2624 544
rect 2556 427 2573 461
rect 2607 427 2624 461
rect 2556 387 2624 427
rect 2556 353 2573 387
rect 2607 353 2624 387
rect 2795 535 2829 923
rect 2795 433 2829 501
rect 2795 383 2829 399
rect 2943 923 2949 942
rect 2943 907 2983 923
rect 2943 905 2977 907
rect 2943 433 2977 871
rect 2943 383 2977 399
rect 3091 757 3125 1023
rect 3222 1053 3290 1093
rect 3222 1019 3239 1053
rect 3273 1019 3290 1053
rect 3397 1366 3431 1446
rect 3397 1298 3431 1332
rect 3397 1230 3431 1264
rect 3397 1162 3431 1196
rect 3397 1093 3431 1128
rect 3397 1027 3431 1059
rect 3485 1366 3519 1404
rect 3485 1298 3519 1332
rect 3485 1230 3519 1264
rect 3485 1162 3519 1196
rect 3485 1093 3519 1128
rect 3573 1366 3607 1446
rect 3573 1298 3607 1332
rect 3573 1230 3607 1264
rect 3573 1162 3607 1196
rect 3573 1111 3607 1128
rect 3661 1366 3695 1404
rect 3661 1298 3695 1332
rect 3661 1230 3695 1264
rect 3661 1162 3695 1196
rect 3485 1057 3519 1059
rect 3661 1093 3695 1128
rect 3749 1366 3783 1446
rect 3749 1298 3783 1332
rect 3749 1230 3783 1264
rect 3749 1162 3783 1196
rect 3749 1111 3783 1128
rect 3888 1423 3956 1446
rect 3888 1389 3905 1423
rect 3939 1389 3956 1423
rect 3888 1349 3956 1389
rect 3888 1315 3905 1349
rect 3939 1315 3956 1349
rect 3888 1275 3956 1315
rect 3888 1241 3905 1275
rect 3939 1241 3956 1275
rect 3888 1201 3956 1241
rect 3888 1167 3905 1201
rect 3939 1167 3956 1201
rect 3888 1127 3956 1167
rect 3661 1057 3695 1059
rect 3888 1093 3905 1127
rect 3939 1093 3956 1127
rect 3485 1023 3791 1057
rect 3222 979 3290 1019
rect 3222 945 3239 979
rect 3273 945 3290 979
rect 3222 905 3290 945
rect 3222 871 3239 905
rect 3273 871 3290 905
rect 3222 822 3290 871
rect 3461 957 3495 973
rect 3615 957 3649 973
rect 3461 831 3495 923
rect 2328 219 2362 316
rect 2556 313 2624 353
rect 2556 279 2573 313
rect 2607 279 2624 313
rect 2328 169 2362 185
rect 2425 263 2459 279
rect 2425 195 2459 229
rect 2117 125 2151 141
rect 1957 91 2020 125
rect 2054 91 2117 125
rect 1923 75 1957 91
rect 2117 75 2151 91
rect 2231 125 2265 161
rect 2425 125 2459 161
rect 2265 91 2328 125
rect 2362 91 2425 125
rect 2231 75 2265 91
rect 2425 75 2459 91
rect 2556 239 2624 279
rect 2556 205 2573 239
rect 2607 205 2624 239
rect 2556 165 2624 205
rect 2556 131 2573 165
rect 2607 131 2624 165
rect 2556 91 2624 131
rect 2556 57 2573 91
rect 2607 57 2624 91
rect 2712 333 2746 349
rect 2906 333 2940 349
rect 3091 348 3125 723
rect 2746 299 2809 333
rect 2843 299 2906 333
rect 2712 261 2746 299
rect 2712 193 2746 227
rect 2906 261 2940 299
rect 2712 123 2746 159
rect 2712 73 2746 89
rect 2809 208 2843 224
rect 2556 34 2624 57
rect 2809 34 2843 174
rect 2906 193 2940 227
rect 3003 314 3125 348
rect 3222 461 3290 544
rect 3222 427 3239 461
rect 3273 427 3290 461
rect 3222 387 3290 427
rect 3222 353 3239 387
rect 3273 353 3290 387
rect 3461 433 3495 797
rect 3461 383 3495 399
rect 3609 923 3615 942
rect 3609 907 3649 923
rect 3609 683 3643 907
rect 3609 433 3643 649
rect 3609 383 3643 399
rect 3757 831 3791 1023
rect 3888 1053 3956 1093
rect 3888 1019 3905 1053
rect 3939 1019 3956 1053
rect 4123 1366 4157 1446
rect 4123 1298 4157 1332
rect 4123 1230 4157 1264
rect 4123 1162 4157 1196
rect 4123 1093 4157 1128
rect 4123 1043 4157 1059
rect 4211 1366 4245 1404
rect 4211 1298 4245 1332
rect 4211 1230 4245 1264
rect 4211 1162 4245 1196
rect 4211 1093 4245 1128
rect 4299 1366 4333 1446
rect 4299 1298 4333 1332
rect 4299 1230 4333 1264
rect 4299 1162 4333 1196
rect 4299 1111 4333 1128
rect 4387 1366 4421 1404
rect 4387 1298 4421 1332
rect 4387 1230 4421 1264
rect 4387 1162 4421 1196
rect 4211 1048 4245 1059
rect 4387 1093 4421 1128
rect 4475 1366 4509 1446
rect 4475 1298 4509 1332
rect 4475 1230 4509 1264
rect 4475 1162 4509 1196
rect 4475 1111 4509 1128
rect 4563 1366 4597 1404
rect 4563 1298 4597 1332
rect 4563 1230 4597 1264
rect 4563 1162 4597 1196
rect 4387 1048 4421 1059
rect 4563 1093 4597 1128
rect 4651 1366 4685 1446
rect 4651 1298 4685 1332
rect 4651 1230 4685 1264
rect 4651 1162 4685 1196
rect 4651 1111 4685 1128
rect 4850 1423 4918 1446
rect 4850 1389 4867 1423
rect 4901 1389 4918 1423
rect 4850 1349 4918 1389
rect 4850 1315 4867 1349
rect 4901 1315 4918 1349
rect 4850 1275 4918 1315
rect 4850 1241 4867 1275
rect 4901 1241 4918 1275
rect 4850 1201 4918 1241
rect 4850 1167 4867 1201
rect 4901 1167 4918 1201
rect 4850 1127 4918 1167
rect 4563 1048 4597 1059
rect 4850 1093 4867 1127
rect 4901 1093 4918 1127
rect 4850 1053 4918 1093
rect 3888 979 3956 1019
rect 4211 1014 4753 1048
rect 3888 945 3905 979
rect 3939 945 3956 979
rect 3888 905 3956 945
rect 3888 871 3905 905
rect 3939 871 3956 905
rect 3888 822 3956 871
rect 4127 957 4161 973
rect 4127 831 4161 923
rect 3003 217 3037 314
rect 3222 313 3290 353
rect 3222 279 3239 313
rect 3273 279 3290 313
rect 3003 167 3037 183
rect 3100 261 3134 277
rect 3100 193 3134 227
rect 2906 123 2940 159
rect 3100 123 3134 159
rect 2940 89 3003 123
rect 3037 89 3100 123
rect 2906 73 2940 89
rect 3100 73 3134 89
rect 3222 239 3290 279
rect 3222 205 3239 239
rect 3273 205 3290 239
rect 3222 165 3290 205
rect 3222 131 3239 165
rect 3273 131 3290 165
rect 3222 91 3290 131
rect 3222 57 3239 91
rect 3273 57 3290 91
rect 3378 333 3412 349
rect 3572 333 3606 349
rect 3757 348 3791 797
rect 3412 299 3475 333
rect 3509 299 3572 333
rect 3378 261 3412 299
rect 3378 193 3412 227
rect 3572 261 3606 299
rect 3378 123 3412 159
rect 3378 73 3412 89
rect 3475 208 3509 224
rect 3222 34 3290 57
rect 3475 34 3509 174
rect 3572 193 3606 227
rect 3669 314 3791 348
rect 3888 461 3956 544
rect 3888 427 3905 461
rect 3939 427 3956 461
rect 3888 387 3956 427
rect 3888 353 3905 387
rect 3939 353 3956 387
rect 4127 433 4161 797
rect 4127 383 4161 399
rect 4349 957 4383 973
rect 4349 461 4383 923
rect 4349 383 4383 399
rect 4571 957 4605 973
rect 4571 757 4605 923
rect 4571 433 4605 723
rect 4571 383 4605 399
rect 4719 683 4753 1014
rect 4850 1019 4867 1053
rect 4901 1019 4918 1053
rect 5025 1366 5059 1446
rect 5025 1298 5059 1332
rect 5025 1230 5059 1264
rect 5025 1162 5059 1196
rect 5025 1093 5059 1128
rect 5025 1027 5059 1059
rect 5113 1366 5147 1404
rect 5113 1298 5147 1332
rect 5113 1230 5147 1264
rect 5113 1162 5147 1196
rect 5113 1093 5147 1128
rect 5201 1366 5235 1446
rect 5201 1298 5235 1332
rect 5201 1230 5235 1264
rect 5201 1162 5235 1196
rect 5201 1111 5235 1128
rect 5289 1366 5323 1404
rect 5289 1298 5323 1332
rect 5289 1230 5323 1264
rect 5289 1162 5323 1196
rect 5113 1057 5147 1059
rect 5289 1093 5323 1128
rect 5377 1366 5411 1446
rect 5377 1298 5411 1332
rect 5377 1230 5411 1264
rect 5377 1162 5411 1196
rect 5377 1111 5411 1128
rect 5516 1423 5584 1446
rect 5516 1389 5533 1423
rect 5567 1389 5584 1423
rect 5516 1349 5584 1389
rect 5516 1315 5533 1349
rect 5567 1315 5584 1349
rect 5516 1275 5584 1315
rect 5516 1241 5533 1275
rect 5567 1241 5584 1275
rect 5516 1201 5584 1241
rect 5516 1167 5533 1201
rect 5567 1167 5584 1201
rect 5516 1127 5584 1167
rect 5289 1057 5323 1059
rect 5516 1093 5533 1127
rect 5567 1093 5584 1127
rect 5113 1023 5419 1057
rect 4850 979 4918 1019
rect 4850 945 4867 979
rect 4901 945 4918 979
rect 4850 905 4918 945
rect 4850 871 4867 905
rect 4901 871 4918 905
rect 4850 822 4918 871
rect 5089 957 5123 973
rect 5243 957 5277 973
rect 3669 217 3703 314
rect 3888 313 3956 353
rect 3888 279 3905 313
rect 3939 279 3956 313
rect 3669 167 3703 183
rect 3766 261 3800 277
rect 3766 193 3800 227
rect 3572 123 3606 159
rect 3766 123 3800 159
rect 3606 89 3669 123
rect 3703 89 3766 123
rect 3572 73 3606 89
rect 3766 73 3800 89
rect 3888 239 3956 279
rect 3888 205 3905 239
rect 3939 205 3956 239
rect 3888 165 3956 205
rect 3888 131 3905 165
rect 3939 131 3956 165
rect 3888 91 3956 131
rect 3888 57 3905 91
rect 3939 57 3956 91
rect 4023 335 4057 351
rect 4217 335 4251 351
rect 4411 335 4445 351
rect 4057 301 4120 335
rect 4154 301 4217 335
rect 4251 301 4314 335
rect 4348 301 4411 335
rect 4023 263 4057 301
rect 4023 195 4057 229
rect 4217 263 4251 301
rect 4411 285 4445 301
rect 4525 335 4559 351
rect 4719 350 4753 649
rect 5089 609 5123 923
rect 4525 263 4559 301
rect 4023 125 4057 161
rect 4023 75 4057 91
rect 4120 210 4154 226
rect 3888 34 3956 57
rect 4120 34 4154 176
rect 4217 195 4251 229
rect 4315 216 4349 232
rect 4525 216 4559 229
rect 4349 195 4559 216
rect 4349 182 4525 195
rect 4315 166 4349 182
rect 4217 125 4251 161
rect 4622 316 4753 350
rect 4850 461 4918 544
rect 4850 427 4867 461
rect 4901 427 4918 461
rect 4850 387 4918 427
rect 4850 353 4867 387
rect 4901 353 4918 387
rect 5089 433 5123 575
rect 5089 383 5123 399
rect 5237 923 5243 942
rect 5237 907 5277 923
rect 5237 831 5271 907
rect 5237 433 5271 797
rect 5237 383 5271 399
rect 5385 535 5419 1023
rect 5516 1053 5584 1093
rect 5516 1019 5533 1053
rect 5567 1019 5584 1053
rect 5751 1366 5785 1446
rect 5751 1298 5785 1332
rect 5751 1230 5785 1264
rect 5751 1162 5785 1196
rect 5751 1093 5785 1128
rect 5751 1043 5785 1059
rect 5839 1366 5873 1404
rect 5839 1298 5873 1332
rect 5839 1230 5873 1264
rect 5839 1162 5873 1196
rect 5839 1093 5873 1128
rect 5927 1366 5961 1446
rect 5927 1298 5961 1332
rect 5927 1230 5961 1264
rect 5927 1162 5961 1196
rect 5927 1111 5961 1128
rect 6015 1366 6049 1404
rect 6015 1298 6049 1332
rect 6015 1230 6049 1264
rect 6015 1162 6049 1196
rect 5839 1048 5873 1059
rect 6015 1093 6049 1128
rect 6103 1366 6137 1446
rect 6103 1298 6137 1332
rect 6103 1230 6137 1264
rect 6103 1162 6137 1196
rect 6103 1111 6137 1128
rect 6191 1366 6225 1404
rect 6191 1298 6225 1332
rect 6191 1230 6225 1264
rect 6191 1162 6225 1196
rect 6015 1048 6049 1059
rect 6191 1093 6225 1128
rect 6279 1366 6313 1446
rect 6279 1298 6313 1332
rect 6279 1230 6313 1264
rect 6279 1162 6313 1196
rect 6279 1111 6313 1128
rect 6478 1423 6546 1446
rect 6478 1389 6495 1423
rect 6529 1389 6546 1423
rect 6478 1349 6546 1389
rect 6478 1315 6495 1349
rect 6529 1315 6546 1349
rect 6478 1275 6546 1315
rect 6478 1241 6495 1275
rect 6529 1241 6546 1275
rect 6478 1201 6546 1241
rect 6478 1167 6495 1201
rect 6529 1167 6546 1201
rect 6478 1127 6546 1167
rect 6191 1048 6225 1059
rect 6478 1093 6495 1127
rect 6529 1093 6546 1127
rect 6478 1053 6546 1093
rect 5516 979 5584 1019
rect 5839 1014 6381 1048
rect 5516 945 5533 979
rect 5567 945 5584 979
rect 5516 905 5584 945
rect 5516 871 5533 905
rect 5567 871 5584 905
rect 5516 822 5584 871
rect 5755 957 5789 973
rect 4622 219 4656 316
rect 4850 313 4918 353
rect 4850 279 4867 313
rect 4901 279 4918 313
rect 4622 169 4656 185
rect 4719 263 4753 279
rect 4719 195 4753 229
rect 4411 125 4445 141
rect 4251 91 4314 125
rect 4348 91 4411 125
rect 4217 75 4251 91
rect 4411 75 4445 91
rect 4525 125 4559 161
rect 4719 125 4753 161
rect 4559 91 4622 125
rect 4656 91 4719 125
rect 4525 75 4559 91
rect 4719 75 4753 91
rect 4850 239 4918 279
rect 4850 205 4867 239
rect 4901 205 4918 239
rect 4850 165 4918 205
rect 4850 131 4867 165
rect 4901 131 4918 165
rect 4850 91 4918 131
rect 4850 57 4867 91
rect 4901 57 4918 91
rect 5006 333 5040 349
rect 5200 333 5234 349
rect 5385 348 5419 501
rect 5040 299 5103 333
rect 5137 299 5200 333
rect 5006 261 5040 299
rect 5006 193 5040 227
rect 5200 261 5234 299
rect 5006 123 5040 159
rect 5006 73 5040 89
rect 5103 208 5137 224
rect 4850 34 4918 57
rect 5103 34 5137 174
rect 5200 193 5234 227
rect 5297 314 5419 348
rect 5516 461 5584 544
rect 5516 427 5533 461
rect 5567 427 5584 461
rect 5516 387 5584 427
rect 5516 353 5533 387
rect 5567 353 5584 387
rect 5755 534 5789 923
rect 5755 433 5789 500
rect 5755 383 5789 399
rect 5977 957 6011 973
rect 5977 905 6011 923
rect 5977 433 6011 871
rect 5977 383 6011 399
rect 6199 957 6233 973
rect 6199 757 6233 923
rect 6347 847 6381 1014
rect 6346 831 6381 847
rect 6380 797 6381 831
rect 6478 1019 6495 1053
rect 6529 1019 6546 1053
rect 6713 1366 6747 1446
rect 6713 1298 6747 1332
rect 6713 1230 6747 1264
rect 6713 1162 6747 1196
rect 6713 1093 6747 1128
rect 6713 1043 6747 1059
rect 6801 1366 6835 1404
rect 6801 1298 6835 1332
rect 6801 1230 6835 1264
rect 6801 1162 6835 1196
rect 6801 1093 6835 1128
rect 6889 1366 6923 1446
rect 6889 1298 6923 1332
rect 6889 1230 6923 1264
rect 6889 1162 6923 1196
rect 6889 1111 6923 1128
rect 6977 1366 7011 1404
rect 6977 1298 7011 1332
rect 6977 1230 7011 1264
rect 6977 1162 7011 1196
rect 6801 1048 6835 1059
rect 6977 1093 7011 1128
rect 7065 1366 7099 1446
rect 7065 1298 7099 1332
rect 7065 1230 7099 1264
rect 7065 1162 7099 1196
rect 7065 1111 7099 1128
rect 7153 1366 7187 1404
rect 7153 1298 7187 1332
rect 7153 1230 7187 1264
rect 7153 1162 7187 1196
rect 6977 1048 7011 1059
rect 7153 1093 7187 1128
rect 7241 1366 7275 1446
rect 7241 1298 7275 1332
rect 7241 1230 7275 1264
rect 7241 1162 7275 1196
rect 7241 1111 7275 1128
rect 7440 1423 7508 1446
rect 7440 1389 7457 1423
rect 7491 1389 7508 1423
rect 7440 1349 7508 1389
rect 7440 1315 7457 1349
rect 7491 1315 7508 1349
rect 7440 1275 7508 1315
rect 7440 1241 7457 1275
rect 7491 1241 7508 1275
rect 7440 1201 7508 1241
rect 7440 1167 7457 1201
rect 7491 1167 7508 1201
rect 7440 1127 7508 1167
rect 7153 1048 7187 1059
rect 7440 1093 7457 1127
rect 7491 1093 7508 1127
rect 7440 1053 7508 1093
rect 6478 979 6546 1019
rect 6801 1014 7343 1048
rect 6478 945 6495 979
rect 6529 945 6546 979
rect 6478 905 6546 945
rect 6478 871 6495 905
rect 6529 871 6546 905
rect 6478 822 6546 871
rect 6717 957 6751 973
rect 6346 781 6381 797
rect 6199 433 6233 723
rect 6199 383 6233 399
rect 5297 217 5331 314
rect 5516 313 5584 353
rect 5516 279 5533 313
rect 5567 279 5584 313
rect 5297 167 5331 183
rect 5394 261 5428 277
rect 5394 193 5428 227
rect 5200 123 5234 159
rect 5394 123 5428 159
rect 5234 89 5297 123
rect 5331 89 5394 123
rect 5200 73 5234 89
rect 5394 73 5428 89
rect 5516 239 5584 279
rect 5516 205 5533 239
rect 5567 205 5584 239
rect 5516 165 5584 205
rect 5516 131 5533 165
rect 5567 131 5584 165
rect 5516 91 5584 131
rect 5516 57 5533 91
rect 5567 57 5584 91
rect 5651 335 5685 351
rect 5845 335 5879 351
rect 6039 335 6073 351
rect 5685 301 5748 335
rect 5782 301 5845 335
rect 5879 301 5942 335
rect 5976 301 6039 335
rect 5651 263 5685 301
rect 5651 195 5685 229
rect 5845 263 5879 301
rect 6039 285 6073 301
rect 6153 335 6187 351
rect 6347 350 6381 781
rect 6153 263 6187 301
rect 5651 125 5685 161
rect 5651 75 5685 91
rect 5748 210 5782 226
rect 5516 34 5584 57
rect 5748 34 5782 176
rect 5845 195 5879 229
rect 5943 216 5977 232
rect 6153 216 6187 229
rect 5977 195 6187 216
rect 5977 182 6153 195
rect 5943 166 5977 182
rect 5845 125 5879 161
rect 6250 316 6381 350
rect 6478 461 6546 544
rect 6478 427 6495 461
rect 6529 427 6546 461
rect 6478 387 6546 427
rect 6478 353 6495 387
rect 6529 353 6546 387
rect 6717 535 6751 923
rect 6717 433 6751 501
rect 6717 383 6751 399
rect 6939 957 6973 973
rect 6939 461 6973 923
rect 6939 383 6973 399
rect 7161 957 7195 973
rect 7161 757 7195 923
rect 7161 433 7195 723
rect 7161 383 7195 399
rect 7309 535 7343 1014
rect 7440 1019 7457 1053
rect 7491 1019 7508 1053
rect 7615 1366 7649 1446
rect 7615 1298 7649 1332
rect 7615 1230 7649 1264
rect 7615 1162 7649 1196
rect 7615 1093 7649 1128
rect 7615 1027 7649 1059
rect 7703 1366 7737 1404
rect 7703 1298 7737 1332
rect 7703 1230 7737 1264
rect 7703 1162 7737 1196
rect 7703 1093 7737 1128
rect 7791 1366 7825 1446
rect 7791 1298 7825 1332
rect 7791 1230 7825 1264
rect 7791 1162 7825 1196
rect 7791 1111 7825 1128
rect 7879 1366 7913 1404
rect 7879 1298 7913 1332
rect 7879 1230 7913 1264
rect 7879 1162 7913 1196
rect 7703 1057 7737 1059
rect 7879 1093 7913 1128
rect 7967 1366 8001 1446
rect 7967 1298 8001 1332
rect 7967 1230 8001 1264
rect 7967 1162 8001 1196
rect 7967 1111 8001 1128
rect 8106 1423 8174 1446
rect 8106 1389 8123 1423
rect 8157 1389 8174 1423
rect 8106 1349 8174 1389
rect 8106 1315 8123 1349
rect 8157 1315 8174 1349
rect 8106 1275 8174 1315
rect 8106 1241 8123 1275
rect 8157 1241 8174 1275
rect 8106 1201 8174 1241
rect 8106 1167 8123 1201
rect 8157 1167 8174 1201
rect 8106 1127 8174 1167
rect 7879 1057 7913 1059
rect 8106 1093 8123 1127
rect 8157 1093 8174 1127
rect 7703 1023 8009 1057
rect 7440 979 7508 1019
rect 7440 945 7457 979
rect 7491 945 7508 979
rect 7440 905 7508 945
rect 7440 871 7457 905
rect 7491 871 7508 905
rect 7440 822 7508 871
rect 7679 957 7713 973
rect 7833 957 7867 973
rect 6250 219 6284 316
rect 6478 313 6546 353
rect 6478 279 6495 313
rect 6529 279 6546 313
rect 6250 169 6284 185
rect 6347 263 6381 279
rect 6347 195 6381 229
rect 6039 125 6073 141
rect 5879 91 5942 125
rect 5976 91 6039 125
rect 5845 75 5879 91
rect 6039 75 6073 91
rect 6153 125 6187 161
rect 6347 125 6381 161
rect 6187 91 6250 125
rect 6284 91 6347 125
rect 6153 75 6187 91
rect 6347 75 6381 91
rect 6478 239 6546 279
rect 6478 205 6495 239
rect 6529 205 6546 239
rect 6478 165 6546 205
rect 6478 131 6495 165
rect 6529 131 6546 165
rect 6478 91 6546 131
rect 6478 57 6495 91
rect 6529 57 6546 91
rect 6613 335 6647 351
rect 6807 335 6841 351
rect 7001 335 7035 351
rect 6647 301 6710 335
rect 6744 301 6807 335
rect 6841 301 6904 335
rect 6938 301 7001 335
rect 6613 263 6647 301
rect 6613 195 6647 229
rect 6807 263 6841 301
rect 7001 285 7035 301
rect 7115 335 7149 351
rect 7309 350 7343 501
rect 7115 263 7149 301
rect 6613 125 6647 161
rect 6613 75 6647 91
rect 6710 210 6744 226
rect 6478 34 6546 57
rect 6710 34 6744 176
rect 6807 195 6841 229
rect 6905 216 6939 232
rect 7115 216 7149 229
rect 6939 195 7149 216
rect 6939 182 7115 195
rect 6905 166 6939 182
rect 6807 125 6841 161
rect 7212 316 7343 350
rect 7440 461 7508 544
rect 7440 427 7457 461
rect 7491 427 7508 461
rect 7440 387 7508 427
rect 7440 353 7457 387
rect 7491 353 7508 387
rect 7679 535 7713 923
rect 7679 433 7713 501
rect 7679 383 7713 399
rect 7827 923 7833 942
rect 7827 907 7867 923
rect 7827 905 7861 907
rect 7827 433 7861 871
rect 7827 383 7861 399
rect 7975 757 8009 1023
rect 8106 1053 8174 1093
rect 8106 1019 8123 1053
rect 8157 1019 8174 1053
rect 8281 1366 8315 1446
rect 8281 1298 8315 1332
rect 8281 1230 8315 1264
rect 8281 1162 8315 1196
rect 8281 1093 8315 1128
rect 8281 1027 8315 1059
rect 8369 1366 8403 1404
rect 8369 1298 8403 1332
rect 8369 1230 8403 1264
rect 8369 1162 8403 1196
rect 8369 1093 8403 1128
rect 8457 1366 8491 1446
rect 8457 1298 8491 1332
rect 8457 1230 8491 1264
rect 8457 1162 8491 1196
rect 8457 1111 8491 1128
rect 8545 1366 8579 1404
rect 8545 1298 8579 1332
rect 8545 1230 8579 1264
rect 8545 1162 8579 1196
rect 8369 1057 8403 1059
rect 8545 1093 8579 1128
rect 8633 1366 8667 1446
rect 8633 1298 8667 1332
rect 8633 1230 8667 1264
rect 8633 1162 8667 1196
rect 8633 1111 8667 1128
rect 8772 1423 8840 1446
rect 8772 1389 8789 1423
rect 8823 1389 8840 1423
rect 8772 1349 8840 1389
rect 8772 1315 8789 1349
rect 8823 1315 8840 1349
rect 8772 1275 8840 1315
rect 8772 1241 8789 1275
rect 8823 1241 8840 1275
rect 8772 1201 8840 1241
rect 8772 1167 8789 1201
rect 8823 1167 8840 1201
rect 8772 1127 8840 1167
rect 8545 1057 8579 1059
rect 8772 1093 8789 1127
rect 8823 1093 8840 1127
rect 8369 1023 8675 1057
rect 8106 979 8174 1019
rect 8106 945 8123 979
rect 8157 945 8174 979
rect 8106 905 8174 945
rect 8106 871 8123 905
rect 8157 871 8174 905
rect 8106 822 8174 871
rect 8345 957 8379 973
rect 8499 957 8533 973
rect 8345 831 8379 923
rect 7212 219 7246 316
rect 7440 313 7508 353
rect 7440 279 7457 313
rect 7491 279 7508 313
rect 7212 169 7246 185
rect 7309 263 7343 279
rect 7309 195 7343 229
rect 7001 125 7035 141
rect 6841 91 6904 125
rect 6938 91 7001 125
rect 6807 75 6841 91
rect 7001 75 7035 91
rect 7115 125 7149 161
rect 7309 125 7343 161
rect 7149 91 7212 125
rect 7246 91 7309 125
rect 7115 75 7149 91
rect 7309 75 7343 91
rect 7440 239 7508 279
rect 7440 205 7457 239
rect 7491 205 7508 239
rect 7440 165 7508 205
rect 7440 131 7457 165
rect 7491 131 7508 165
rect 7440 91 7508 131
rect 7440 57 7457 91
rect 7491 57 7508 91
rect 7596 333 7630 349
rect 7790 333 7824 349
rect 7975 348 8009 723
rect 7630 299 7693 333
rect 7727 299 7790 333
rect 7596 261 7630 299
rect 7596 193 7630 227
rect 7790 261 7824 299
rect 7596 123 7630 159
rect 7596 73 7630 89
rect 7693 208 7727 224
rect 7440 34 7508 57
rect 7693 34 7727 174
rect 7790 193 7824 227
rect 7887 314 8009 348
rect 8106 461 8174 544
rect 8106 427 8123 461
rect 8157 427 8174 461
rect 8106 387 8174 427
rect 8106 353 8123 387
rect 8157 353 8174 387
rect 8345 433 8379 797
rect 8345 383 8379 399
rect 8493 923 8499 942
rect 8493 907 8533 923
rect 8493 831 8527 907
rect 8493 433 8527 797
rect 8493 383 8527 399
rect 8641 535 8675 1023
rect 8772 1053 8840 1093
rect 8772 1019 8789 1053
rect 8823 1019 8840 1053
rect 9007 1366 9041 1446
rect 9007 1298 9041 1332
rect 9007 1230 9041 1264
rect 9007 1162 9041 1196
rect 9007 1093 9041 1128
rect 9007 1043 9041 1059
rect 9095 1366 9129 1404
rect 9095 1298 9129 1332
rect 9095 1230 9129 1264
rect 9095 1162 9129 1196
rect 9095 1093 9129 1128
rect 9183 1366 9217 1446
rect 9183 1298 9217 1332
rect 9183 1230 9217 1264
rect 9183 1162 9217 1196
rect 9183 1111 9217 1128
rect 9271 1366 9305 1404
rect 9271 1298 9305 1332
rect 9271 1230 9305 1264
rect 9271 1162 9305 1196
rect 9095 1048 9129 1059
rect 9271 1093 9305 1128
rect 9359 1366 9393 1446
rect 9359 1298 9393 1332
rect 9359 1230 9393 1264
rect 9359 1162 9393 1196
rect 9359 1111 9393 1128
rect 9447 1366 9481 1404
rect 9447 1298 9481 1332
rect 9447 1230 9481 1264
rect 9447 1162 9481 1196
rect 9271 1048 9305 1059
rect 9447 1093 9481 1128
rect 9535 1366 9569 1446
rect 9535 1298 9569 1332
rect 9535 1230 9569 1264
rect 9535 1162 9569 1196
rect 9535 1111 9569 1128
rect 9734 1423 9802 1446
rect 9734 1389 9751 1423
rect 9785 1389 9802 1423
rect 9734 1349 9802 1389
rect 9734 1315 9751 1349
rect 9785 1315 9802 1349
rect 9734 1275 9802 1315
rect 9734 1241 9751 1275
rect 9785 1241 9802 1275
rect 9734 1201 9802 1241
rect 9734 1167 9751 1201
rect 9785 1167 9802 1201
rect 9734 1127 9802 1167
rect 9447 1048 9481 1059
rect 9734 1093 9751 1127
rect 9785 1093 9802 1127
rect 9734 1053 9802 1093
rect 8772 979 8840 1019
rect 9095 1014 9637 1048
rect 8772 945 8789 979
rect 8823 945 8840 979
rect 8772 905 8840 945
rect 8772 871 8789 905
rect 8823 871 8840 905
rect 8772 822 8840 871
rect 9011 957 9045 973
rect 7887 217 7921 314
rect 8106 313 8174 353
rect 8106 279 8123 313
rect 8157 279 8174 313
rect 7887 167 7921 183
rect 7984 261 8018 277
rect 7984 193 8018 227
rect 7790 123 7824 159
rect 7984 123 8018 159
rect 7824 89 7887 123
rect 7921 89 7984 123
rect 7790 73 7824 89
rect 7984 73 8018 89
rect 8106 239 8174 279
rect 8106 205 8123 239
rect 8157 205 8174 239
rect 8106 165 8174 205
rect 8106 131 8123 165
rect 8157 131 8174 165
rect 8106 91 8174 131
rect 8106 57 8123 91
rect 8157 57 8174 91
rect 8262 333 8296 349
rect 8456 333 8490 349
rect 8641 348 8675 501
rect 8296 299 8359 333
rect 8393 299 8456 333
rect 8262 261 8296 299
rect 8262 193 8296 227
rect 8456 261 8490 299
rect 8262 123 8296 159
rect 8262 73 8296 89
rect 8359 208 8393 224
rect 8106 34 8174 57
rect 8359 34 8393 174
rect 8456 193 8490 227
rect 8553 314 8675 348
rect 8772 461 8840 544
rect 8772 427 8789 461
rect 8823 427 8840 461
rect 8772 387 8840 427
rect 8772 353 8789 387
rect 8823 353 8840 387
rect 9011 535 9045 923
rect 9011 433 9045 501
rect 9011 383 9045 399
rect 9233 957 9267 973
rect 9233 461 9267 923
rect 9233 383 9267 399
rect 9455 957 9489 973
rect 9455 757 9489 923
rect 9455 433 9489 723
rect 9455 383 9489 399
rect 9603 831 9637 1014
rect 9734 1019 9751 1053
rect 9785 1019 9802 1053
rect 9909 1366 9943 1446
rect 9909 1298 9943 1332
rect 9909 1230 9943 1264
rect 9909 1162 9943 1196
rect 9909 1093 9943 1128
rect 9909 1027 9943 1059
rect 9997 1366 10031 1404
rect 9997 1298 10031 1332
rect 9997 1230 10031 1264
rect 9997 1162 10031 1196
rect 9997 1093 10031 1128
rect 10085 1366 10119 1446
rect 10085 1298 10119 1332
rect 10085 1230 10119 1264
rect 10085 1162 10119 1196
rect 10085 1111 10119 1128
rect 10173 1366 10207 1404
rect 10173 1298 10207 1332
rect 10173 1230 10207 1264
rect 10173 1162 10207 1196
rect 9997 1057 10031 1059
rect 10173 1093 10207 1128
rect 10261 1366 10295 1446
rect 10261 1298 10295 1332
rect 10261 1230 10295 1264
rect 10261 1162 10295 1196
rect 10261 1111 10295 1128
rect 10400 1423 10468 1446
rect 10400 1389 10417 1423
rect 10451 1389 10468 1423
rect 10400 1349 10468 1389
rect 10400 1315 10417 1349
rect 10451 1315 10468 1349
rect 10400 1275 10468 1315
rect 10400 1241 10417 1275
rect 10451 1241 10468 1275
rect 10400 1201 10468 1241
rect 10400 1167 10417 1201
rect 10451 1167 10468 1201
rect 10400 1127 10468 1167
rect 10173 1057 10207 1059
rect 10400 1093 10417 1127
rect 10451 1093 10468 1127
rect 9997 1023 10303 1057
rect 9734 979 9802 1019
rect 9734 945 9751 979
rect 9785 945 9802 979
rect 9734 905 9802 945
rect 9734 871 9751 905
rect 9785 871 9802 905
rect 9734 822 9802 871
rect 9973 957 10007 973
rect 10127 957 10161 973
rect 9603 535 9637 797
rect 9973 609 10007 923
rect 8553 217 8587 314
rect 8772 313 8840 353
rect 8772 279 8789 313
rect 8823 279 8840 313
rect 8553 167 8587 183
rect 8650 261 8684 277
rect 8650 193 8684 227
rect 8456 123 8490 159
rect 8650 123 8684 159
rect 8490 89 8553 123
rect 8587 89 8650 123
rect 8456 73 8490 89
rect 8650 73 8684 89
rect 8772 239 8840 279
rect 8772 205 8789 239
rect 8823 205 8840 239
rect 8772 165 8840 205
rect 8772 131 8789 165
rect 8823 131 8840 165
rect 8772 91 8840 131
rect 8772 57 8789 91
rect 8823 57 8840 91
rect 8907 335 8941 351
rect 9101 335 9135 351
rect 9295 335 9329 351
rect 8941 301 9004 335
rect 9038 301 9101 335
rect 9135 301 9198 335
rect 9232 301 9295 335
rect 8907 263 8941 301
rect 8907 195 8941 229
rect 9101 263 9135 301
rect 9295 285 9329 301
rect 9409 335 9443 351
rect 9603 350 9637 501
rect 9409 263 9443 301
rect 8907 125 8941 161
rect 8907 75 8941 91
rect 9004 210 9038 226
rect 8772 34 8840 57
rect 9004 34 9038 176
rect 9101 195 9135 229
rect 9199 216 9233 232
rect 9409 216 9443 229
rect 9233 195 9443 216
rect 9233 182 9409 195
rect 9199 166 9233 182
rect 9101 125 9135 161
rect 9506 316 9637 350
rect 9734 461 9802 544
rect 9734 427 9751 461
rect 9785 427 9802 461
rect 9734 387 9802 427
rect 9734 353 9751 387
rect 9785 353 9802 387
rect 9973 433 10007 575
rect 9973 383 10007 399
rect 10121 923 10127 942
rect 10121 907 10161 923
rect 10121 831 10155 907
rect 10121 433 10155 797
rect 10121 383 10155 399
rect 10269 535 10303 1023
rect 10400 1053 10468 1093
rect 10400 1019 10417 1053
rect 10451 1019 10468 1053
rect 10635 1366 10669 1446
rect 10635 1298 10669 1332
rect 10635 1230 10669 1264
rect 10635 1162 10669 1196
rect 10635 1093 10669 1128
rect 10635 1043 10669 1059
rect 10723 1366 10757 1404
rect 10723 1298 10757 1332
rect 10723 1230 10757 1264
rect 10723 1162 10757 1196
rect 10723 1093 10757 1128
rect 10811 1366 10845 1446
rect 10811 1298 10845 1332
rect 10811 1230 10845 1264
rect 10811 1162 10845 1196
rect 10811 1111 10845 1128
rect 10899 1366 10933 1404
rect 10899 1298 10933 1332
rect 10899 1230 10933 1264
rect 10899 1162 10933 1196
rect 10723 1048 10757 1059
rect 10899 1093 10933 1128
rect 10987 1366 11021 1446
rect 10987 1298 11021 1332
rect 10987 1230 11021 1264
rect 10987 1162 11021 1196
rect 10987 1111 11021 1128
rect 11075 1366 11109 1404
rect 11075 1298 11109 1332
rect 11075 1230 11109 1264
rect 11075 1162 11109 1196
rect 10899 1048 10933 1059
rect 11075 1093 11109 1128
rect 11163 1366 11197 1446
rect 11163 1298 11197 1332
rect 11163 1230 11197 1264
rect 11163 1162 11197 1196
rect 11163 1111 11197 1128
rect 11362 1423 11430 1446
rect 11362 1389 11379 1423
rect 11413 1389 11430 1423
rect 11362 1349 11430 1389
rect 11362 1315 11379 1349
rect 11413 1315 11430 1349
rect 11362 1275 11430 1315
rect 11362 1241 11379 1275
rect 11413 1241 11430 1275
rect 11362 1201 11430 1241
rect 11362 1167 11379 1201
rect 11413 1167 11430 1201
rect 11362 1127 11430 1167
rect 11075 1048 11109 1059
rect 11362 1093 11379 1127
rect 11413 1093 11430 1127
rect 11362 1053 11430 1093
rect 10400 979 10468 1019
rect 10723 1014 11265 1048
rect 10400 945 10417 979
rect 10451 945 10468 979
rect 10400 905 10468 945
rect 10400 871 10417 905
rect 10451 871 10468 905
rect 10400 822 10468 871
rect 10639 957 10673 973
rect 9506 219 9540 316
rect 9734 313 9802 353
rect 9734 279 9751 313
rect 9785 279 9802 313
rect 9506 169 9540 185
rect 9603 263 9637 279
rect 9603 195 9637 229
rect 9295 125 9329 141
rect 9135 91 9198 125
rect 9232 91 9295 125
rect 9101 75 9135 91
rect 9295 75 9329 91
rect 9409 125 9443 161
rect 9603 125 9637 161
rect 9443 91 9506 125
rect 9540 91 9603 125
rect 9409 75 9443 91
rect 9603 75 9637 91
rect 9734 239 9802 279
rect 9734 205 9751 239
rect 9785 205 9802 239
rect 9734 165 9802 205
rect 9734 131 9751 165
rect 9785 131 9802 165
rect 9734 91 9802 131
rect 9734 57 9751 91
rect 9785 57 9802 91
rect 9890 333 9924 349
rect 10084 333 10118 349
rect 10269 348 10303 501
rect 9924 299 9987 333
rect 10021 299 10084 333
rect 9890 261 9924 299
rect 9890 193 9924 227
rect 10084 261 10118 299
rect 9890 123 9924 159
rect 9890 73 9924 89
rect 9987 208 10021 224
rect 9734 34 9802 57
rect 9987 34 10021 174
rect 10084 193 10118 227
rect 10181 314 10303 348
rect 10400 461 10468 544
rect 10400 427 10417 461
rect 10451 427 10468 461
rect 10400 387 10468 427
rect 10400 353 10417 387
rect 10451 353 10468 387
rect 10639 534 10673 923
rect 10639 433 10673 500
rect 10639 383 10673 399
rect 10861 957 10895 973
rect 10861 905 10895 923
rect 10861 433 10895 871
rect 10861 383 10895 399
rect 11083 957 11117 973
rect 11083 757 11117 923
rect 11231 847 11265 1014
rect 11230 831 11265 847
rect 11264 797 11265 831
rect 11362 1019 11379 1053
rect 11413 1019 11430 1053
rect 11597 1366 11631 1446
rect 11597 1298 11631 1332
rect 11597 1230 11631 1264
rect 11597 1162 11631 1196
rect 11597 1093 11631 1128
rect 11597 1043 11631 1059
rect 11685 1366 11719 1404
rect 11685 1298 11719 1332
rect 11685 1230 11719 1264
rect 11685 1162 11719 1196
rect 11685 1093 11719 1128
rect 11773 1366 11807 1446
rect 11773 1298 11807 1332
rect 11773 1230 11807 1264
rect 11773 1162 11807 1196
rect 11773 1111 11807 1128
rect 11861 1366 11895 1404
rect 11861 1298 11895 1332
rect 11861 1230 11895 1264
rect 11861 1162 11895 1196
rect 11685 1048 11719 1059
rect 11861 1093 11895 1128
rect 11949 1366 11983 1446
rect 11949 1298 11983 1332
rect 11949 1230 11983 1264
rect 11949 1162 11983 1196
rect 11949 1111 11983 1128
rect 12037 1366 12071 1404
rect 12037 1298 12071 1332
rect 12037 1230 12071 1264
rect 12037 1162 12071 1196
rect 11861 1048 11895 1059
rect 12037 1093 12071 1128
rect 12125 1366 12159 1446
rect 12125 1298 12159 1332
rect 12125 1230 12159 1264
rect 12125 1162 12159 1196
rect 12125 1111 12159 1128
rect 12324 1423 12392 1446
rect 12324 1389 12341 1423
rect 12375 1389 12392 1423
rect 12324 1349 12392 1389
rect 12324 1315 12341 1349
rect 12375 1315 12392 1349
rect 12324 1275 12392 1315
rect 12324 1241 12341 1275
rect 12375 1241 12392 1275
rect 12324 1201 12392 1241
rect 12324 1167 12341 1201
rect 12375 1167 12392 1201
rect 12324 1127 12392 1167
rect 12037 1048 12071 1059
rect 12324 1093 12341 1127
rect 12375 1093 12392 1127
rect 12324 1053 12392 1093
rect 11362 979 11430 1019
rect 11685 1014 12227 1048
rect 11362 945 11379 979
rect 11413 945 11430 979
rect 11362 905 11430 945
rect 11362 871 11379 905
rect 11413 871 11430 905
rect 11362 822 11430 871
rect 11601 957 11635 973
rect 11230 781 11265 797
rect 11083 433 11117 723
rect 11083 383 11117 399
rect 10181 217 10215 314
rect 10400 313 10468 353
rect 10400 279 10417 313
rect 10451 279 10468 313
rect 10181 167 10215 183
rect 10278 261 10312 277
rect 10278 193 10312 227
rect 10084 123 10118 159
rect 10278 123 10312 159
rect 10118 89 10181 123
rect 10215 89 10278 123
rect 10084 73 10118 89
rect 10278 73 10312 89
rect 10400 239 10468 279
rect 10400 205 10417 239
rect 10451 205 10468 239
rect 10400 165 10468 205
rect 10400 131 10417 165
rect 10451 131 10468 165
rect 10400 91 10468 131
rect 10400 57 10417 91
rect 10451 57 10468 91
rect 10535 335 10569 351
rect 10729 335 10763 351
rect 10923 335 10957 351
rect 10569 301 10632 335
rect 10666 301 10729 335
rect 10763 301 10826 335
rect 10860 301 10923 335
rect 10535 263 10569 301
rect 10535 195 10569 229
rect 10729 263 10763 301
rect 10923 285 10957 301
rect 11037 335 11071 351
rect 11231 350 11265 781
rect 11037 263 11071 301
rect 10535 125 10569 161
rect 10535 75 10569 91
rect 10632 210 10666 226
rect 10400 34 10468 57
rect 10632 34 10666 176
rect 10729 195 10763 229
rect 10827 216 10861 232
rect 11037 216 11071 229
rect 10861 195 11071 216
rect 10861 182 11037 195
rect 10827 166 10861 182
rect 10729 125 10763 161
rect 11134 316 11265 350
rect 11362 461 11430 544
rect 11362 427 11379 461
rect 11413 427 11430 461
rect 11362 387 11430 427
rect 11362 353 11379 387
rect 11413 353 11430 387
rect 11601 535 11635 923
rect 11601 433 11635 501
rect 11601 383 11635 399
rect 11823 957 11857 973
rect 11823 461 11857 923
rect 11823 383 11857 399
rect 12045 957 12079 973
rect 12045 757 12079 923
rect 12045 433 12079 723
rect 12045 383 12079 399
rect 12193 535 12227 1014
rect 12324 1019 12341 1053
rect 12375 1019 12392 1053
rect 12499 1366 12533 1446
rect 12499 1298 12533 1332
rect 12499 1230 12533 1264
rect 12499 1162 12533 1196
rect 12499 1093 12533 1128
rect 12499 1027 12533 1059
rect 12587 1366 12621 1404
rect 12587 1298 12621 1332
rect 12587 1230 12621 1264
rect 12587 1162 12621 1196
rect 12587 1093 12621 1128
rect 12675 1366 12709 1446
rect 12675 1298 12709 1332
rect 12675 1230 12709 1264
rect 12675 1162 12709 1196
rect 12675 1111 12709 1128
rect 12763 1366 12797 1404
rect 12763 1298 12797 1332
rect 12763 1230 12797 1264
rect 12763 1162 12797 1196
rect 12587 1057 12621 1059
rect 12763 1093 12797 1128
rect 12851 1366 12885 1446
rect 12851 1298 12885 1332
rect 12851 1230 12885 1264
rect 12851 1162 12885 1196
rect 12851 1111 12885 1128
rect 12990 1423 13058 1446
rect 12990 1389 13007 1423
rect 13041 1389 13058 1423
rect 12990 1349 13058 1389
rect 12990 1315 13007 1349
rect 13041 1315 13058 1349
rect 12990 1275 13058 1315
rect 12990 1241 13007 1275
rect 13041 1241 13058 1275
rect 12990 1201 13058 1241
rect 12990 1167 13007 1201
rect 13041 1167 13058 1201
rect 12990 1127 13058 1167
rect 12763 1057 12797 1059
rect 12990 1093 13007 1127
rect 13041 1093 13058 1127
rect 12587 1023 12893 1057
rect 12324 979 12392 1019
rect 12324 945 12341 979
rect 12375 945 12392 979
rect 12324 905 12392 945
rect 12324 871 12341 905
rect 12375 871 12392 905
rect 12324 822 12392 871
rect 12563 957 12597 973
rect 12717 957 12751 973
rect 11134 219 11168 316
rect 11362 313 11430 353
rect 11362 279 11379 313
rect 11413 279 11430 313
rect 11134 169 11168 185
rect 11231 263 11265 279
rect 11231 195 11265 229
rect 10923 125 10957 141
rect 10763 91 10826 125
rect 10860 91 10923 125
rect 10729 75 10763 91
rect 10923 75 10957 91
rect 11037 125 11071 161
rect 11231 125 11265 161
rect 11071 91 11134 125
rect 11168 91 11231 125
rect 11037 75 11071 91
rect 11231 75 11265 91
rect 11362 239 11430 279
rect 11362 205 11379 239
rect 11413 205 11430 239
rect 11362 165 11430 205
rect 11362 131 11379 165
rect 11413 131 11430 165
rect 11362 91 11430 131
rect 11362 57 11379 91
rect 11413 57 11430 91
rect 11497 335 11531 351
rect 11691 335 11725 351
rect 11885 335 11919 351
rect 11531 301 11594 335
rect 11628 301 11691 335
rect 11725 301 11788 335
rect 11822 301 11885 335
rect 11497 263 11531 301
rect 11497 195 11531 229
rect 11691 263 11725 301
rect 11885 285 11919 301
rect 11999 335 12033 351
rect 12193 350 12227 501
rect 11999 263 12033 301
rect 11497 125 11531 161
rect 11497 75 11531 91
rect 11594 210 11628 226
rect 11362 34 11430 57
rect 11594 34 11628 176
rect 11691 195 11725 229
rect 11789 216 11823 232
rect 11999 216 12033 229
rect 11823 195 12033 216
rect 11823 182 11999 195
rect 11789 166 11823 182
rect 11691 125 11725 161
rect 12096 316 12227 350
rect 12324 461 12392 544
rect 12324 427 12341 461
rect 12375 427 12392 461
rect 12324 387 12392 427
rect 12324 353 12341 387
rect 12375 353 12392 387
rect 12563 535 12597 923
rect 12563 433 12597 501
rect 12563 383 12597 399
rect 12711 923 12717 942
rect 12711 907 12751 923
rect 12711 905 12745 907
rect 12711 433 12745 871
rect 12711 383 12745 399
rect 12859 757 12893 1023
rect 12990 1053 13058 1093
rect 12990 1019 13007 1053
rect 13041 1019 13058 1053
rect 13165 1366 13199 1446
rect 13165 1298 13199 1332
rect 13165 1230 13199 1264
rect 13165 1162 13199 1196
rect 13165 1093 13199 1128
rect 13165 1027 13199 1059
rect 13253 1366 13287 1404
rect 13253 1298 13287 1332
rect 13253 1230 13287 1264
rect 13253 1162 13287 1196
rect 13253 1093 13287 1128
rect 13341 1366 13375 1446
rect 13341 1298 13375 1332
rect 13341 1230 13375 1264
rect 13341 1162 13375 1196
rect 13341 1111 13375 1128
rect 13429 1366 13463 1404
rect 13429 1298 13463 1332
rect 13429 1230 13463 1264
rect 13429 1162 13463 1196
rect 13253 1057 13287 1059
rect 13429 1093 13463 1128
rect 13517 1366 13551 1446
rect 13517 1298 13551 1332
rect 13517 1230 13551 1264
rect 13517 1162 13551 1196
rect 13517 1111 13551 1128
rect 13656 1423 13724 1446
rect 13656 1389 13673 1423
rect 13707 1389 13724 1423
rect 13656 1349 13724 1389
rect 13656 1315 13673 1349
rect 13707 1315 13724 1349
rect 13656 1275 13724 1315
rect 13656 1241 13673 1275
rect 13707 1241 13724 1275
rect 13656 1201 13724 1241
rect 13656 1167 13673 1201
rect 13707 1167 13724 1201
rect 13656 1127 13724 1167
rect 13429 1057 13463 1059
rect 13656 1093 13673 1127
rect 13707 1093 13724 1127
rect 13253 1023 13559 1057
rect 12990 979 13058 1019
rect 12990 945 13007 979
rect 13041 945 13058 979
rect 13525 979 13559 1023
rect 12990 905 13058 945
rect 12990 871 13007 905
rect 13041 871 13058 905
rect 12990 822 13058 871
rect 13229 957 13263 973
rect 13383 957 13417 973
rect 13229 831 13263 923
rect 12096 219 12130 316
rect 12324 313 12392 353
rect 12324 279 12341 313
rect 12375 279 12392 313
rect 12096 169 12130 185
rect 12193 263 12227 279
rect 12193 195 12227 229
rect 11885 125 11919 141
rect 11725 91 11788 125
rect 11822 91 11885 125
rect 11691 75 11725 91
rect 11885 75 11919 91
rect 11999 125 12033 161
rect 12193 125 12227 161
rect 12033 91 12096 125
rect 12130 91 12193 125
rect 11999 75 12033 91
rect 12193 75 12227 91
rect 12324 239 12392 279
rect 12324 205 12341 239
rect 12375 205 12392 239
rect 12324 165 12392 205
rect 12324 131 12341 165
rect 12375 131 12392 165
rect 12324 91 12392 131
rect 12324 57 12341 91
rect 12375 57 12392 91
rect 12480 333 12514 349
rect 12674 333 12708 349
rect 12859 348 12893 723
rect 12514 299 12577 333
rect 12611 299 12674 333
rect 12480 261 12514 299
rect 12480 193 12514 227
rect 12674 261 12708 299
rect 12480 123 12514 159
rect 12480 73 12514 89
rect 12577 208 12611 224
rect 12324 34 12392 57
rect 12577 34 12611 174
rect 12674 193 12708 227
rect 12771 314 12893 348
rect 12990 461 13058 544
rect 12990 427 13007 461
rect 13041 427 13058 461
rect 12990 387 13058 427
rect 12990 353 13007 387
rect 13041 353 13058 387
rect 13229 433 13263 797
rect 13229 383 13263 399
rect 13377 923 13383 942
rect 13377 907 13417 923
rect 13377 905 13411 907
rect 13377 433 13411 871
rect 13377 383 13411 399
rect 12771 217 12805 314
rect 12990 313 13058 353
rect 12990 279 13007 313
rect 13041 279 13058 313
rect 12771 167 12805 183
rect 12868 261 12902 277
rect 12868 193 12902 227
rect 12674 123 12708 159
rect 12868 123 12902 159
rect 12708 89 12771 123
rect 12805 89 12868 123
rect 12674 73 12708 89
rect 12868 73 12902 89
rect 12990 239 13058 279
rect 12990 205 13007 239
rect 13041 205 13058 239
rect 12990 165 13058 205
rect 12990 131 13007 165
rect 13041 131 13058 165
rect 12990 91 13058 131
rect 12990 57 13007 91
rect 13041 57 13058 91
rect 13146 333 13180 349
rect 13340 333 13374 349
rect 13525 348 13559 945
rect 13656 1053 13724 1093
rect 13656 1019 13673 1053
rect 13707 1019 13724 1053
rect 13891 1366 13925 1446
rect 13891 1298 13925 1332
rect 13891 1230 13925 1264
rect 13891 1162 13925 1196
rect 13891 1093 13925 1128
rect 13891 1043 13925 1059
rect 13979 1366 14013 1404
rect 13979 1298 14013 1332
rect 13979 1230 14013 1264
rect 13979 1162 14013 1196
rect 13979 1093 14013 1128
rect 14067 1366 14101 1446
rect 14067 1298 14101 1332
rect 14067 1230 14101 1264
rect 14067 1162 14101 1196
rect 14067 1111 14101 1128
rect 14155 1366 14189 1404
rect 14155 1298 14189 1332
rect 14155 1230 14189 1264
rect 14155 1162 14189 1196
rect 13979 1048 14013 1059
rect 14155 1093 14189 1128
rect 14243 1366 14277 1446
rect 14243 1298 14277 1332
rect 14243 1230 14277 1264
rect 14243 1162 14277 1196
rect 14243 1111 14277 1128
rect 14331 1366 14365 1404
rect 14331 1298 14365 1332
rect 14331 1230 14365 1264
rect 14331 1162 14365 1196
rect 14155 1048 14189 1059
rect 14331 1093 14365 1128
rect 14419 1366 14453 1446
rect 14419 1298 14453 1332
rect 14419 1230 14453 1264
rect 14419 1162 14453 1196
rect 14419 1111 14453 1128
rect 14618 1423 14686 1446
rect 14618 1389 14635 1423
rect 14669 1389 14686 1423
rect 14618 1349 14686 1389
rect 14618 1315 14635 1349
rect 14669 1315 14686 1349
rect 14618 1275 14686 1315
rect 14618 1241 14635 1275
rect 14669 1241 14686 1275
rect 14618 1201 14686 1241
rect 14618 1167 14635 1201
rect 14669 1167 14686 1201
rect 14618 1127 14686 1167
rect 14331 1048 14365 1059
rect 14618 1093 14635 1127
rect 14669 1093 14686 1127
rect 14618 1053 14686 1093
rect 13656 979 13724 1019
rect 13979 1014 14521 1048
rect 13656 945 13673 979
rect 13707 945 13724 979
rect 13656 905 13724 945
rect 13656 871 13673 905
rect 13707 871 13724 905
rect 13656 822 13724 871
rect 13895 979 13929 995
rect 13180 299 13243 333
rect 13277 299 13340 333
rect 13146 261 13180 299
rect 13146 193 13180 227
rect 13340 261 13374 299
rect 13146 123 13180 159
rect 13146 73 13180 89
rect 13243 208 13277 224
rect 12990 34 13058 57
rect 13243 34 13277 174
rect 13340 193 13374 227
rect 13437 314 13559 348
rect 13656 461 13724 544
rect 13656 427 13673 461
rect 13707 427 13724 461
rect 13656 387 13724 427
rect 13656 353 13673 387
rect 13707 353 13724 387
rect 13895 433 13929 923
rect 13895 383 13929 399
rect 14117 957 14151 973
rect 14117 461 14151 923
rect 14117 383 14151 399
rect 14339 957 14373 973
rect 14339 757 14373 923
rect 14339 433 14373 723
rect 14339 383 14373 399
rect 14487 905 14521 1014
rect 13437 217 13471 314
rect 13656 313 13724 353
rect 13656 279 13673 313
rect 13707 279 13724 313
rect 13437 167 13471 183
rect 13534 261 13568 277
rect 13534 193 13568 227
rect 13340 123 13374 159
rect 13534 123 13568 159
rect 13374 89 13437 123
rect 13471 89 13534 123
rect 13340 73 13374 89
rect 13534 73 13568 89
rect 13656 239 13724 279
rect 13656 205 13673 239
rect 13707 205 13724 239
rect 13656 165 13724 205
rect 13656 131 13673 165
rect 13707 131 13724 165
rect 13656 91 13724 131
rect 13656 57 13673 91
rect 13707 57 13724 91
rect 13791 335 13825 351
rect 13985 335 14019 351
rect 14179 335 14213 351
rect 13825 301 13888 335
rect 13922 301 13985 335
rect 14019 301 14082 335
rect 14116 301 14179 335
rect 13791 263 13825 301
rect 13791 195 13825 229
rect 13985 263 14019 301
rect 14179 285 14213 301
rect 14293 335 14327 351
rect 14487 350 14521 871
rect 14618 1019 14635 1053
rect 14669 1019 14686 1053
rect 14793 1365 14827 1446
rect 14793 1297 14827 1331
rect 14793 1229 14827 1263
rect 14793 1161 14827 1195
rect 14793 1093 14827 1127
rect 14793 1025 14827 1059
rect 14881 1365 14917 1399
rect 14969 1365 15003 1446
rect 14881 1297 14915 1331
rect 14881 1229 14915 1263
rect 14881 1161 14915 1195
rect 14881 1093 14915 1127
rect 14969 1297 15003 1331
rect 14969 1229 15003 1263
rect 14969 1161 15003 1195
rect 14969 1111 15003 1127
rect 15057 1365 15091 1399
rect 15057 1297 15091 1331
rect 15057 1229 15091 1263
rect 15057 1161 15091 1195
rect 15057 1059 15091 1127
rect 14881 1025 15057 1059
rect 15145 1365 15179 1446
rect 15145 1297 15179 1331
rect 15145 1229 15179 1263
rect 15145 1161 15179 1195
rect 15145 1093 15179 1127
rect 15145 1025 15179 1059
rect 15284 1423 15352 1446
rect 15284 1389 15301 1423
rect 15335 1389 15352 1423
rect 15950 1423 16018 1446
rect 15284 1349 15352 1389
rect 15284 1315 15301 1349
rect 15335 1315 15352 1349
rect 15284 1275 15352 1315
rect 15284 1241 15301 1275
rect 15335 1241 15352 1275
rect 15284 1201 15352 1241
rect 15284 1167 15301 1201
rect 15335 1167 15352 1201
rect 15284 1127 15352 1167
rect 15284 1093 15301 1127
rect 15335 1093 15352 1127
rect 15284 1053 15352 1093
rect 14618 979 14686 1019
rect 15057 1009 15091 1025
rect 15284 1019 15301 1053
rect 15335 1019 15352 1053
rect 14618 945 14635 979
rect 14669 945 14686 979
rect 15284 979 15352 1019
rect 15457 1365 15843 1399
rect 15457 1297 15491 1331
rect 15457 1229 15491 1263
rect 15457 1161 15491 1195
rect 15457 1059 15491 1127
rect 15545 1297 15579 1313
rect 15545 1229 15579 1263
rect 15545 1161 15579 1195
rect 15545 1093 15579 1127
rect 15633 1297 15667 1331
rect 15633 1229 15667 1263
rect 15633 1161 15667 1195
rect 15633 1111 15667 1127
rect 15721 1297 15755 1313
rect 15721 1229 15755 1263
rect 15721 1161 15755 1195
rect 15721 1059 15755 1127
rect 15809 1297 15843 1331
rect 15809 1229 15843 1263
rect 15809 1161 15843 1195
rect 15809 1075 15843 1127
rect 15950 1389 15967 1423
rect 16001 1389 16018 1423
rect 16616 1423 16684 1446
rect 15950 1349 16018 1389
rect 15950 1315 15967 1349
rect 16001 1315 16018 1349
rect 15950 1275 16018 1315
rect 15950 1241 15967 1275
rect 16001 1241 16018 1275
rect 15950 1201 16018 1241
rect 15950 1167 15967 1201
rect 16001 1167 16018 1201
rect 15950 1127 16018 1167
rect 15950 1093 15967 1127
rect 16001 1093 16018 1127
rect 15545 1025 15721 1059
rect 15457 1009 15491 1025
rect 15721 1009 15755 1025
rect 15950 1053 16018 1093
rect 15950 1019 15967 1053
rect 16001 1019 16018 1053
rect 14618 905 14686 945
rect 14618 871 14635 905
rect 14669 871 14686 905
rect 14618 822 14686 871
rect 14783 958 14817 974
rect 15013 958 15047 974
rect 14783 905 14817 924
rect 14293 263 14327 301
rect 13791 125 13825 161
rect 13791 75 13825 91
rect 13888 210 13922 226
rect 13656 34 13724 57
rect 13888 34 13922 176
rect 13985 195 14019 229
rect 14083 216 14117 232
rect 14293 216 14327 229
rect 14117 195 14327 216
rect 14117 182 14293 195
rect 14083 166 14117 182
rect 13985 125 14019 161
rect 14390 316 14521 350
rect 14618 461 14686 544
rect 14618 427 14635 461
rect 14669 427 14686 461
rect 14618 387 14686 427
rect 14618 353 14635 387
rect 14669 353 14686 387
rect 14783 433 14817 871
rect 14783 383 14817 399
rect 15005 924 15013 942
rect 15005 908 15047 924
rect 15284 945 15301 979
rect 15335 945 15352 979
rect 15950 979 16018 1019
rect 16125 1365 16511 1399
rect 16125 1297 16159 1331
rect 16125 1229 16159 1263
rect 16125 1161 16159 1195
rect 16125 1059 16159 1127
rect 16213 1297 16247 1313
rect 16213 1229 16247 1263
rect 16213 1161 16247 1195
rect 16213 1093 16247 1127
rect 16301 1297 16335 1331
rect 16301 1229 16335 1263
rect 16301 1161 16335 1195
rect 16301 1111 16335 1127
rect 16389 1297 16423 1313
rect 16389 1229 16423 1263
rect 16389 1161 16423 1195
rect 16389 1093 16423 1127
rect 16477 1297 16511 1331
rect 16477 1229 16511 1263
rect 16477 1161 16511 1195
rect 16477 1111 16511 1127
rect 16616 1389 16633 1423
rect 16667 1389 16684 1423
rect 16616 1349 16684 1389
rect 16616 1315 16633 1349
rect 16667 1315 16684 1349
rect 16616 1275 16684 1315
rect 16616 1241 16633 1275
rect 16667 1241 16684 1275
rect 16616 1201 16684 1241
rect 16616 1167 16633 1201
rect 16667 1167 16684 1201
rect 16616 1127 16684 1167
rect 16616 1093 16633 1127
rect 16667 1093 16684 1127
rect 16213 1025 16519 1059
rect 16125 1009 16159 1025
rect 15005 831 15039 908
rect 15284 905 15352 945
rect 15284 871 15301 905
rect 15335 871 15352 905
rect 15284 822 15352 871
rect 15523 958 15557 974
rect 15523 905 15557 924
rect 15005 609 15039 797
rect 15005 433 15039 575
rect 15005 383 15039 399
rect 15284 461 15352 544
rect 15284 427 15301 461
rect 15335 427 15352 461
rect 15284 387 15352 427
rect 14390 219 14424 316
rect 14618 313 14686 353
rect 15284 353 15301 387
rect 15335 353 15352 387
rect 15523 433 15557 871
rect 15523 383 15557 399
rect 15819 958 15853 974
rect 15819 683 15853 924
rect 15950 945 15967 979
rect 16001 945 16018 979
rect 15950 905 16018 945
rect 15950 871 15967 905
rect 16001 871 16018 905
rect 15950 822 16018 871
rect 16115 958 16149 974
rect 15819 433 15853 649
rect 15819 383 15853 399
rect 15950 461 16018 544
rect 15950 427 15967 461
rect 16001 427 16018 461
rect 15950 387 16018 427
rect 14618 279 14635 313
rect 14669 279 14686 313
rect 14390 169 14424 185
rect 14487 263 14521 279
rect 14487 195 14521 229
rect 14179 125 14213 141
rect 14019 91 14082 125
rect 14116 91 14179 125
rect 13985 75 14019 91
rect 14179 75 14213 91
rect 14293 125 14327 161
rect 14487 125 14521 161
rect 14327 91 14390 125
rect 14424 91 14487 125
rect 14293 75 14327 91
rect 14487 75 14521 91
rect 14618 239 14686 279
rect 14618 205 14635 239
rect 14669 205 14686 239
rect 14618 165 14686 205
rect 14618 131 14635 165
rect 14669 131 14686 165
rect 14618 91 14686 131
rect 14618 57 14635 91
rect 14669 57 14686 91
rect 14774 333 14808 349
rect 14968 333 15002 349
rect 14808 299 14871 333
rect 14905 299 14968 333
rect 14774 261 14808 299
rect 14774 193 14808 227
rect 14968 261 15002 299
rect 15162 333 15196 349
rect 15065 253 15099 269
rect 14774 123 14808 159
rect 14774 73 14808 89
rect 14871 208 14905 224
rect 14618 34 14686 57
rect 14871 34 14905 174
rect 14968 193 15002 227
rect 15064 219 15065 234
rect 15064 217 15099 219
rect 15098 203 15099 217
rect 15162 261 15196 299
rect 15064 167 15098 183
rect 15162 193 15196 227
rect 14968 123 15002 159
rect 15162 123 15196 159
rect 15002 89 15064 123
rect 15098 89 15162 123
rect 14968 73 15002 89
rect 15162 73 15196 89
rect 15284 313 15352 353
rect 15950 353 15967 387
rect 16001 353 16018 387
rect 16115 433 16149 924
rect 16115 383 16149 399
rect 16337 958 16375 974
rect 16337 924 16341 958
rect 16337 908 16375 924
rect 16337 831 16371 908
rect 16337 433 16371 797
rect 16337 383 16371 399
rect 16485 831 16519 1025
rect 16616 1053 16684 1093
rect 16616 1019 16633 1053
rect 16667 1019 16684 1053
rect 16768 1366 16802 1446
rect 16768 1298 16802 1332
rect 16768 1230 16802 1264
rect 16768 1162 16802 1196
rect 16768 1093 16802 1128
rect 16768 1037 16802 1059
rect 16856 1366 16890 1404
rect 16856 1298 16890 1332
rect 16856 1230 16890 1264
rect 16856 1162 16890 1196
rect 16856 1093 16890 1128
rect 16616 979 16684 1019
rect 16616 945 16633 979
rect 16667 945 16684 979
rect 16616 905 16684 945
rect 16616 871 16633 905
rect 16667 871 16684 905
rect 16616 822 16684 871
rect 16781 957 16815 973
rect 16781 831 16815 923
rect 16856 933 16890 1059
rect 16944 1366 16978 1446
rect 16944 1298 16978 1332
rect 16944 1230 16978 1264
rect 16944 1162 16978 1196
rect 16944 1093 16978 1128
rect 16944 1037 16978 1059
rect 17060 1423 17128 1446
rect 17060 1389 17077 1423
rect 17111 1389 17128 1423
rect 17060 1349 17128 1389
rect 17060 1315 17077 1349
rect 17111 1315 17128 1349
rect 17060 1275 17128 1315
rect 17060 1241 17077 1275
rect 17111 1241 17128 1275
rect 17060 1201 17128 1241
rect 17060 1167 17077 1201
rect 17111 1167 17128 1201
rect 17060 1127 17128 1167
rect 17060 1093 17077 1127
rect 17111 1093 17128 1127
rect 17060 1053 17128 1093
rect 17060 1019 17077 1053
rect 17111 1019 17128 1053
rect 17060 979 17128 1019
rect 17060 945 17077 979
rect 17111 945 17128 979
rect 16856 899 16963 933
rect 15284 279 15301 313
rect 15335 279 15352 313
rect 15284 239 15352 279
rect 15284 205 15301 239
rect 15335 205 15352 239
rect 15284 165 15352 205
rect 15284 131 15301 165
rect 15335 131 15352 165
rect 15284 91 15352 131
rect 15284 57 15301 91
rect 15335 57 15352 91
rect 15440 333 15474 349
rect 15634 333 15668 349
rect 15474 299 15537 333
rect 15571 299 15634 333
rect 15440 261 15474 299
rect 15440 193 15474 227
rect 15634 261 15668 299
rect 15828 333 15862 349
rect 15440 123 15474 159
rect 15440 73 15474 89
rect 15537 208 15571 224
rect 15284 34 15352 57
rect 15537 34 15571 174
rect 15634 193 15668 227
rect 15731 253 15765 269
rect 15731 217 15765 219
rect 15731 167 15765 183
rect 15828 261 15862 299
rect 15828 193 15862 227
rect 15634 123 15668 159
rect 15828 123 15862 159
rect 15668 89 15731 123
rect 15765 89 15828 123
rect 15634 73 15668 89
rect 15828 73 15862 89
rect 15950 313 16018 353
rect 15950 279 15967 313
rect 16001 279 16018 313
rect 15950 239 16018 279
rect 15950 205 15967 239
rect 16001 205 16018 239
rect 15950 165 16018 205
rect 15950 131 15967 165
rect 16001 131 16018 165
rect 15950 91 16018 131
rect 15950 57 15967 91
rect 16001 57 16018 91
rect 16106 333 16140 349
rect 16300 333 16334 349
rect 16485 346 16519 797
rect 16140 299 16203 333
rect 16237 299 16300 333
rect 16106 261 16140 299
rect 16106 193 16140 227
rect 16300 261 16334 299
rect 16106 123 16140 159
rect 16106 73 16140 89
rect 16203 208 16237 224
rect 15950 34 16018 57
rect 16203 34 16237 174
rect 16300 193 16334 227
rect 16397 312 16519 346
rect 16616 461 16684 544
rect 16616 427 16633 461
rect 16667 427 16684 461
rect 16616 387 16684 427
rect 16616 353 16633 387
rect 16667 353 16684 387
rect 16781 434 16815 797
rect 16929 433 16963 899
rect 17060 905 17128 945
rect 17060 871 17077 905
rect 17111 871 17128 905
rect 17060 822 17128 871
rect 16781 384 16815 400
rect 16855 399 16963 433
rect 17060 461 17128 544
rect 17060 427 17077 461
rect 17111 427 17128 461
rect 16616 313 16684 353
rect 16397 253 16431 312
rect 16616 279 16633 313
rect 16667 279 16684 313
rect 16397 217 16431 219
rect 16397 167 16431 183
rect 16494 261 16528 278
rect 16494 193 16528 227
rect 16300 123 16334 159
rect 16494 123 16528 159
rect 16334 89 16397 123
rect 16431 89 16494 123
rect 16300 73 16334 89
rect 16494 73 16528 89
rect 16616 239 16684 279
rect 16616 205 16633 239
rect 16667 205 16684 239
rect 16616 165 16684 205
rect 16616 131 16633 165
rect 16667 131 16684 165
rect 16616 91 16684 131
rect 16616 57 16633 91
rect 16667 57 16684 91
rect 16616 34 16684 57
rect 16759 334 16793 350
rect 16759 262 16793 300
rect 16759 194 16793 228
rect 16855 218 16889 399
rect 17060 387 17128 427
rect 17060 353 17077 387
rect 17111 353 17128 387
rect 16855 168 16889 184
rect 16953 334 16987 350
rect 16953 262 16987 300
rect 16953 194 16987 228
rect 16759 124 16793 160
rect 16953 124 16987 160
rect 16793 90 16855 124
rect 16889 90 16953 124
rect 16759 34 16793 90
rect 16856 34 16890 90
rect 16953 34 16987 90
rect 17060 313 17128 353
rect 17060 279 17077 313
rect 17111 279 17128 313
rect 17060 239 17128 279
rect 17060 205 17077 239
rect 17111 205 17128 239
rect 17060 165 17128 205
rect 17060 131 17077 165
rect 17111 131 17128 165
rect 17060 91 17128 131
rect 17060 57 17077 91
rect 17111 57 17128 91
rect 17060 34 17128 57
rect -34 17 17128 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5163 17
rect 5197 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5755 17
rect 5789 -17 5829 17
rect 5863 -17 5903 17
rect 5937 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6125 17
rect 6159 -17 6199 17
rect 6233 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6569 17
rect 6603 -17 6643 17
rect 6677 -17 6717 17
rect 6751 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7087 17
rect 7121 -17 7161 17
rect 7195 -17 7235 17
rect 7269 -17 7309 17
rect 7343 -17 7383 17
rect 7417 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7679 17
rect 7713 -17 7753 17
rect 7787 -17 7827 17
rect 7861 -17 7901 17
rect 7935 -17 7975 17
rect 8009 -17 8049 17
rect 8083 -17 8197 17
rect 8231 -17 8271 17
rect 8305 -17 8345 17
rect 8379 -17 8419 17
rect 8453 -17 8493 17
rect 8527 -17 8567 17
rect 8601 -17 8641 17
rect 8675 -17 8715 17
rect 8749 -17 8863 17
rect 8897 -17 8937 17
rect 8971 -17 9011 17
rect 9045 -17 9085 17
rect 9119 -17 9159 17
rect 9193 -17 9233 17
rect 9267 -17 9307 17
rect 9341 -17 9381 17
rect 9415 -17 9455 17
rect 9489 -17 9529 17
rect 9563 -17 9603 17
rect 9637 -17 9677 17
rect 9711 -17 9825 17
rect 9859 -17 9899 17
rect 9933 -17 9973 17
rect 10007 -17 10047 17
rect 10081 -17 10121 17
rect 10155 -17 10195 17
rect 10229 -17 10269 17
rect 10303 -17 10343 17
rect 10377 -17 10491 17
rect 10525 -17 10565 17
rect 10599 -17 10639 17
rect 10673 -17 10713 17
rect 10747 -17 10787 17
rect 10821 -17 10861 17
rect 10895 -17 10935 17
rect 10969 -17 11009 17
rect 11043 -17 11083 17
rect 11117 -17 11157 17
rect 11191 -17 11231 17
rect 11265 -17 11305 17
rect 11339 -17 11453 17
rect 11487 -17 11527 17
rect 11561 -17 11601 17
rect 11635 -17 11675 17
rect 11709 -17 11749 17
rect 11783 -17 11823 17
rect 11857 -17 11897 17
rect 11931 -17 11971 17
rect 12005 -17 12045 17
rect 12079 -17 12119 17
rect 12153 -17 12193 17
rect 12227 -17 12267 17
rect 12301 -17 12415 17
rect 12449 -17 12489 17
rect 12523 -17 12563 17
rect 12597 -17 12637 17
rect 12671 -17 12711 17
rect 12745 -17 12785 17
rect 12819 -17 12859 17
rect 12893 -17 12933 17
rect 12967 -17 13081 17
rect 13115 -17 13155 17
rect 13189 -17 13229 17
rect 13263 -17 13303 17
rect 13337 -17 13377 17
rect 13411 -17 13451 17
rect 13485 -17 13525 17
rect 13559 -17 13599 17
rect 13633 -17 13747 17
rect 13781 -17 13821 17
rect 13855 -17 13895 17
rect 13929 -17 13969 17
rect 14003 -17 14043 17
rect 14077 -17 14117 17
rect 14151 -17 14191 17
rect 14225 -17 14265 17
rect 14299 -17 14339 17
rect 14373 -17 14413 17
rect 14447 -17 14487 17
rect 14521 -17 14561 17
rect 14595 -17 14709 17
rect 14743 -17 14783 17
rect 14817 -17 14857 17
rect 14891 -17 14931 17
rect 14965 -17 15005 17
rect 15039 -17 15079 17
rect 15113 -17 15153 17
rect 15187 -17 15227 17
rect 15261 -17 15375 17
rect 15409 -17 15449 17
rect 15483 -17 15523 17
rect 15557 -17 15597 17
rect 15631 -17 15671 17
rect 15705 -17 15745 17
rect 15779 -17 15819 17
rect 15853 -17 15893 17
rect 15927 -17 16041 17
rect 16075 -17 16115 17
rect 16149 -17 16189 17
rect 16223 -17 16263 17
rect 16297 -17 16337 17
rect 16371 -17 16411 17
rect 16445 -17 16485 17
rect 16519 -17 16559 17
rect 16593 -17 16707 17
rect 16741 -17 16781 17
rect 16815 -17 16855 17
rect 16889 -17 16929 17
rect 16963 -17 17003 17
rect 17037 -17 17128 17
rect -34 -34 17128 -17
<< viali >>
rect 57 1463 91 1497
rect 131 1463 165 1497
rect 205 1463 239 1497
rect 279 1463 313 1497
rect 353 1463 387 1497
rect 427 1463 461 1497
rect 501 1463 535 1497
rect 575 1463 609 1497
rect 723 1463 757 1497
rect 797 1463 831 1497
rect 871 1463 905 1497
rect 945 1463 979 1497
rect 1019 1463 1053 1497
rect 1093 1463 1127 1497
rect 1167 1463 1201 1497
rect 1241 1463 1275 1497
rect 1315 1463 1349 1497
rect 1389 1463 1423 1497
rect 1463 1463 1497 1497
rect 1537 1463 1571 1497
rect 1685 1463 1719 1497
rect 1759 1463 1793 1497
rect 1833 1463 1867 1497
rect 1907 1463 1941 1497
rect 1981 1463 2015 1497
rect 2055 1463 2089 1497
rect 2129 1463 2163 1497
rect 2203 1463 2237 1497
rect 2277 1463 2311 1497
rect 2351 1463 2385 1497
rect 2425 1463 2459 1497
rect 2499 1463 2533 1497
rect 2647 1463 2681 1497
rect 2721 1463 2755 1497
rect 2795 1463 2829 1497
rect 2869 1463 2903 1497
rect 2943 1463 2977 1497
rect 3017 1463 3051 1497
rect 3091 1463 3125 1497
rect 3165 1463 3199 1497
rect 3313 1463 3347 1497
rect 3387 1463 3421 1497
rect 3461 1463 3495 1497
rect 3535 1463 3569 1497
rect 3609 1463 3643 1497
rect 3683 1463 3717 1497
rect 3757 1463 3791 1497
rect 3831 1463 3865 1497
rect 3979 1463 4013 1497
rect 4053 1463 4087 1497
rect 4127 1463 4161 1497
rect 4201 1463 4235 1497
rect 4275 1463 4309 1497
rect 4349 1463 4383 1497
rect 4423 1463 4457 1497
rect 4497 1463 4531 1497
rect 4571 1463 4605 1497
rect 4645 1463 4679 1497
rect 4719 1463 4753 1497
rect 4793 1463 4827 1497
rect 4941 1463 4975 1497
rect 5015 1463 5049 1497
rect 5089 1463 5123 1497
rect 5163 1463 5197 1497
rect 5237 1463 5271 1497
rect 5311 1463 5345 1497
rect 5385 1463 5419 1497
rect 5459 1463 5493 1497
rect 5607 1463 5641 1497
rect 5681 1463 5715 1497
rect 5755 1463 5789 1497
rect 5829 1463 5863 1497
rect 5903 1463 5937 1497
rect 5977 1463 6011 1497
rect 6051 1463 6085 1497
rect 6125 1463 6159 1497
rect 6199 1463 6233 1497
rect 6273 1463 6307 1497
rect 6347 1463 6381 1497
rect 6421 1463 6455 1497
rect 6569 1463 6603 1497
rect 6643 1463 6677 1497
rect 6717 1463 6751 1497
rect 6791 1463 6825 1497
rect 6865 1463 6899 1497
rect 6939 1463 6973 1497
rect 7013 1463 7047 1497
rect 7087 1463 7121 1497
rect 7161 1463 7195 1497
rect 7235 1463 7269 1497
rect 7309 1463 7343 1497
rect 7383 1463 7417 1497
rect 7531 1463 7565 1497
rect 7605 1463 7639 1497
rect 7679 1463 7713 1497
rect 7753 1463 7787 1497
rect 7827 1463 7861 1497
rect 7901 1463 7935 1497
rect 7975 1463 8009 1497
rect 8049 1463 8083 1497
rect 8197 1463 8231 1497
rect 8271 1463 8305 1497
rect 8345 1463 8379 1497
rect 8419 1463 8453 1497
rect 8493 1463 8527 1497
rect 8567 1463 8601 1497
rect 8641 1463 8675 1497
rect 8715 1463 8749 1497
rect 8863 1463 8897 1497
rect 8937 1463 8971 1497
rect 9011 1463 9045 1497
rect 9085 1463 9119 1497
rect 9159 1463 9193 1497
rect 9233 1463 9267 1497
rect 9307 1463 9341 1497
rect 9381 1463 9415 1497
rect 9455 1463 9489 1497
rect 9529 1463 9563 1497
rect 9603 1463 9637 1497
rect 9677 1463 9711 1497
rect 9825 1463 9859 1497
rect 9899 1463 9933 1497
rect 9973 1463 10007 1497
rect 10047 1463 10081 1497
rect 10121 1463 10155 1497
rect 10195 1463 10229 1497
rect 10269 1463 10303 1497
rect 10343 1463 10377 1497
rect 10491 1463 10525 1497
rect 10565 1463 10599 1497
rect 10639 1463 10673 1497
rect 10713 1463 10747 1497
rect 10787 1463 10821 1497
rect 10861 1463 10895 1497
rect 10935 1463 10969 1497
rect 11009 1463 11043 1497
rect 11083 1463 11117 1497
rect 11157 1463 11191 1497
rect 11231 1463 11265 1497
rect 11305 1463 11339 1497
rect 11453 1463 11487 1497
rect 11527 1463 11561 1497
rect 11601 1463 11635 1497
rect 11675 1463 11709 1497
rect 11749 1463 11783 1497
rect 11823 1463 11857 1497
rect 11897 1463 11931 1497
rect 11971 1463 12005 1497
rect 12045 1463 12079 1497
rect 12119 1463 12153 1497
rect 12193 1463 12227 1497
rect 12267 1463 12301 1497
rect 12415 1463 12449 1497
rect 12489 1463 12523 1497
rect 12563 1463 12597 1497
rect 12637 1463 12671 1497
rect 12711 1463 12745 1497
rect 12785 1463 12819 1497
rect 12859 1463 12893 1497
rect 12933 1463 12967 1497
rect 13081 1463 13115 1497
rect 13155 1463 13189 1497
rect 13229 1463 13263 1497
rect 13303 1463 13337 1497
rect 13377 1463 13411 1497
rect 13451 1463 13485 1497
rect 13525 1463 13559 1497
rect 13599 1463 13633 1497
rect 13747 1463 13781 1497
rect 13821 1463 13855 1497
rect 13895 1463 13929 1497
rect 13969 1463 14003 1497
rect 14043 1463 14077 1497
rect 14117 1463 14151 1497
rect 14191 1463 14225 1497
rect 14265 1463 14299 1497
rect 14339 1463 14373 1497
rect 14413 1463 14447 1497
rect 14487 1463 14521 1497
rect 14561 1463 14595 1497
rect 14709 1463 14743 1497
rect 14783 1463 14817 1497
rect 14857 1463 14891 1497
rect 14931 1463 14965 1497
rect 15005 1463 15039 1497
rect 15079 1463 15113 1497
rect 15153 1463 15187 1497
rect 15227 1463 15261 1497
rect 15375 1463 15409 1497
rect 15449 1463 15483 1497
rect 15523 1463 15557 1497
rect 15597 1463 15631 1497
rect 15671 1463 15705 1497
rect 15745 1463 15779 1497
rect 15819 1463 15853 1497
rect 15893 1463 15927 1497
rect 16041 1463 16075 1497
rect 16115 1463 16149 1497
rect 16189 1463 16223 1497
rect 16263 1463 16297 1497
rect 16337 1463 16371 1497
rect 16411 1463 16445 1497
rect 16485 1463 16519 1497
rect 16559 1463 16593 1497
rect 16707 1463 16741 1497
rect 16781 1463 16815 1497
rect 16855 1463 16889 1497
rect 16929 1463 16963 1497
rect 17003 1463 17037 1497
rect 205 575 239 609
rect 353 797 387 831
rect 501 501 535 535
rect 871 500 905 534
rect 1093 871 1127 905
rect 1462 797 1496 831
rect 1315 723 1349 757
rect 1833 501 1867 535
rect 2055 433 2089 461
rect 2055 427 2089 433
rect 2277 723 2311 757
rect 2425 501 2459 535
rect 2795 501 2829 535
rect 2943 871 2977 905
rect 3091 723 3125 757
rect 3461 797 3495 831
rect 3609 649 3643 683
rect 3757 797 3791 831
rect 4127 797 4161 831
rect 4349 433 4383 461
rect 4349 427 4383 433
rect 4571 723 4605 757
rect 4719 649 4753 683
rect 5089 575 5123 609
rect 5237 797 5271 831
rect 5385 501 5419 535
rect 5755 500 5789 534
rect 5977 871 6011 905
rect 6346 797 6380 831
rect 6199 723 6233 757
rect 6717 501 6751 535
rect 6939 433 6973 461
rect 6939 427 6973 433
rect 7161 723 7195 757
rect 7309 501 7343 535
rect 7679 501 7713 535
rect 7827 871 7861 905
rect 7975 723 8009 757
rect 8345 797 8379 831
rect 8493 797 8527 831
rect 8641 501 8675 535
rect 9011 501 9045 535
rect 9233 433 9267 461
rect 9233 427 9267 433
rect 9455 723 9489 757
rect 9603 797 9637 831
rect 9973 575 10007 609
rect 9603 501 9637 535
rect 10121 797 10155 831
rect 10269 501 10303 535
rect 10639 500 10673 534
rect 10861 871 10895 905
rect 11230 797 11264 831
rect 11083 723 11117 757
rect 11601 501 11635 535
rect 11823 433 11857 461
rect 11823 427 11857 433
rect 12045 723 12079 757
rect 12193 501 12227 535
rect 12563 501 12597 535
rect 12711 871 12745 905
rect 12859 723 12893 757
rect 13229 797 13263 831
rect 13525 945 13559 979
rect 13377 871 13411 905
rect 13895 957 13929 979
rect 13895 945 13929 957
rect 14117 433 14151 461
rect 14117 427 14151 433
rect 14339 723 14373 757
rect 14487 871 14521 905
rect 15057 1025 15091 1059
rect 15457 1025 15491 1059
rect 15721 1025 15755 1059
rect 14783 871 14817 905
rect 16125 1025 16159 1059
rect 15005 797 15039 831
rect 15523 871 15557 905
rect 15005 575 15039 609
rect 15819 649 15853 683
rect 15819 399 15853 433
rect 15065 219 15099 253
rect 16115 399 16149 433
rect 16337 797 16371 831
rect 16485 797 16519 831
rect 15731 219 15765 253
rect 16781 797 16815 831
rect 16397 219 16431 253
rect 57 -17 91 17
rect 131 -17 165 17
rect 205 -17 239 17
rect 279 -17 313 17
rect 353 -17 387 17
rect 427 -17 461 17
rect 501 -17 535 17
rect 575 -17 609 17
rect 723 -17 757 17
rect 797 -17 831 17
rect 871 -17 905 17
rect 945 -17 979 17
rect 1019 -17 1053 17
rect 1093 -17 1127 17
rect 1167 -17 1201 17
rect 1241 -17 1275 17
rect 1315 -17 1349 17
rect 1389 -17 1423 17
rect 1463 -17 1497 17
rect 1537 -17 1571 17
rect 1685 -17 1719 17
rect 1759 -17 1793 17
rect 1833 -17 1867 17
rect 1907 -17 1941 17
rect 1981 -17 2015 17
rect 2055 -17 2089 17
rect 2129 -17 2163 17
rect 2203 -17 2237 17
rect 2277 -17 2311 17
rect 2351 -17 2385 17
rect 2425 -17 2459 17
rect 2499 -17 2533 17
rect 2647 -17 2681 17
rect 2721 -17 2755 17
rect 2795 -17 2829 17
rect 2869 -17 2903 17
rect 2943 -17 2977 17
rect 3017 -17 3051 17
rect 3091 -17 3125 17
rect 3165 -17 3199 17
rect 3313 -17 3347 17
rect 3387 -17 3421 17
rect 3461 -17 3495 17
rect 3535 -17 3569 17
rect 3609 -17 3643 17
rect 3683 -17 3717 17
rect 3757 -17 3791 17
rect 3831 -17 3865 17
rect 3979 -17 4013 17
rect 4053 -17 4087 17
rect 4127 -17 4161 17
rect 4201 -17 4235 17
rect 4275 -17 4309 17
rect 4349 -17 4383 17
rect 4423 -17 4457 17
rect 4497 -17 4531 17
rect 4571 -17 4605 17
rect 4645 -17 4679 17
rect 4719 -17 4753 17
rect 4793 -17 4827 17
rect 4941 -17 4975 17
rect 5015 -17 5049 17
rect 5089 -17 5123 17
rect 5163 -17 5197 17
rect 5237 -17 5271 17
rect 5311 -17 5345 17
rect 5385 -17 5419 17
rect 5459 -17 5493 17
rect 5607 -17 5641 17
rect 5681 -17 5715 17
rect 5755 -17 5789 17
rect 5829 -17 5863 17
rect 5903 -17 5937 17
rect 5977 -17 6011 17
rect 6051 -17 6085 17
rect 6125 -17 6159 17
rect 6199 -17 6233 17
rect 6273 -17 6307 17
rect 6347 -17 6381 17
rect 6421 -17 6455 17
rect 6569 -17 6603 17
rect 6643 -17 6677 17
rect 6717 -17 6751 17
rect 6791 -17 6825 17
rect 6865 -17 6899 17
rect 6939 -17 6973 17
rect 7013 -17 7047 17
rect 7087 -17 7121 17
rect 7161 -17 7195 17
rect 7235 -17 7269 17
rect 7309 -17 7343 17
rect 7383 -17 7417 17
rect 7531 -17 7565 17
rect 7605 -17 7639 17
rect 7679 -17 7713 17
rect 7753 -17 7787 17
rect 7827 -17 7861 17
rect 7901 -17 7935 17
rect 7975 -17 8009 17
rect 8049 -17 8083 17
rect 8197 -17 8231 17
rect 8271 -17 8305 17
rect 8345 -17 8379 17
rect 8419 -17 8453 17
rect 8493 -17 8527 17
rect 8567 -17 8601 17
rect 8641 -17 8675 17
rect 8715 -17 8749 17
rect 8863 -17 8897 17
rect 8937 -17 8971 17
rect 9011 -17 9045 17
rect 9085 -17 9119 17
rect 9159 -17 9193 17
rect 9233 -17 9267 17
rect 9307 -17 9341 17
rect 9381 -17 9415 17
rect 9455 -17 9489 17
rect 9529 -17 9563 17
rect 9603 -17 9637 17
rect 9677 -17 9711 17
rect 9825 -17 9859 17
rect 9899 -17 9933 17
rect 9973 -17 10007 17
rect 10047 -17 10081 17
rect 10121 -17 10155 17
rect 10195 -17 10229 17
rect 10269 -17 10303 17
rect 10343 -17 10377 17
rect 10491 -17 10525 17
rect 10565 -17 10599 17
rect 10639 -17 10673 17
rect 10713 -17 10747 17
rect 10787 -17 10821 17
rect 10861 -17 10895 17
rect 10935 -17 10969 17
rect 11009 -17 11043 17
rect 11083 -17 11117 17
rect 11157 -17 11191 17
rect 11231 -17 11265 17
rect 11305 -17 11339 17
rect 11453 -17 11487 17
rect 11527 -17 11561 17
rect 11601 -17 11635 17
rect 11675 -17 11709 17
rect 11749 -17 11783 17
rect 11823 -17 11857 17
rect 11897 -17 11931 17
rect 11971 -17 12005 17
rect 12045 -17 12079 17
rect 12119 -17 12153 17
rect 12193 -17 12227 17
rect 12267 -17 12301 17
rect 12415 -17 12449 17
rect 12489 -17 12523 17
rect 12563 -17 12597 17
rect 12637 -17 12671 17
rect 12711 -17 12745 17
rect 12785 -17 12819 17
rect 12859 -17 12893 17
rect 12933 -17 12967 17
rect 13081 -17 13115 17
rect 13155 -17 13189 17
rect 13229 -17 13263 17
rect 13303 -17 13337 17
rect 13377 -17 13411 17
rect 13451 -17 13485 17
rect 13525 -17 13559 17
rect 13599 -17 13633 17
rect 13747 -17 13781 17
rect 13821 -17 13855 17
rect 13895 -17 13929 17
rect 13969 -17 14003 17
rect 14043 -17 14077 17
rect 14117 -17 14151 17
rect 14191 -17 14225 17
rect 14265 -17 14299 17
rect 14339 -17 14373 17
rect 14413 -17 14447 17
rect 14487 -17 14521 17
rect 14561 -17 14595 17
rect 14709 -17 14743 17
rect 14783 -17 14817 17
rect 14857 -17 14891 17
rect 14931 -17 14965 17
rect 15005 -17 15039 17
rect 15079 -17 15113 17
rect 15153 -17 15187 17
rect 15227 -17 15261 17
rect 15375 -17 15409 17
rect 15449 -17 15483 17
rect 15523 -17 15557 17
rect 15597 -17 15631 17
rect 15671 -17 15705 17
rect 15745 -17 15779 17
rect 15819 -17 15853 17
rect 15893 -17 15927 17
rect 16041 -17 16075 17
rect 16115 -17 16149 17
rect 16189 -17 16223 17
rect 16263 -17 16297 17
rect 16337 -17 16371 17
rect 16411 -17 16445 17
rect 16485 -17 16519 17
rect 16559 -17 16593 17
rect 16707 -17 16741 17
rect 16781 -17 16815 17
rect 16855 -17 16889 17
rect 16929 -17 16963 17
rect 17003 -17 17037 17
<< metal1 >>
rect -34 1497 17128 1514
rect -34 1463 57 1497
rect 91 1463 131 1497
rect 165 1463 205 1497
rect 239 1463 279 1497
rect 313 1463 353 1497
rect 387 1463 427 1497
rect 461 1463 501 1497
rect 535 1463 575 1497
rect 609 1463 723 1497
rect 757 1463 797 1497
rect 831 1463 871 1497
rect 905 1463 945 1497
rect 979 1463 1019 1497
rect 1053 1463 1093 1497
rect 1127 1463 1167 1497
rect 1201 1463 1241 1497
rect 1275 1463 1315 1497
rect 1349 1463 1389 1497
rect 1423 1463 1463 1497
rect 1497 1463 1537 1497
rect 1571 1463 1685 1497
rect 1719 1463 1759 1497
rect 1793 1463 1833 1497
rect 1867 1463 1907 1497
rect 1941 1463 1981 1497
rect 2015 1463 2055 1497
rect 2089 1463 2129 1497
rect 2163 1463 2203 1497
rect 2237 1463 2277 1497
rect 2311 1463 2351 1497
rect 2385 1463 2425 1497
rect 2459 1463 2499 1497
rect 2533 1463 2647 1497
rect 2681 1463 2721 1497
rect 2755 1463 2795 1497
rect 2829 1463 2869 1497
rect 2903 1463 2943 1497
rect 2977 1463 3017 1497
rect 3051 1463 3091 1497
rect 3125 1463 3165 1497
rect 3199 1463 3313 1497
rect 3347 1463 3387 1497
rect 3421 1463 3461 1497
rect 3495 1463 3535 1497
rect 3569 1463 3609 1497
rect 3643 1463 3683 1497
rect 3717 1463 3757 1497
rect 3791 1463 3831 1497
rect 3865 1463 3979 1497
rect 4013 1463 4053 1497
rect 4087 1463 4127 1497
rect 4161 1463 4201 1497
rect 4235 1463 4275 1497
rect 4309 1463 4349 1497
rect 4383 1463 4423 1497
rect 4457 1463 4497 1497
rect 4531 1463 4571 1497
rect 4605 1463 4645 1497
rect 4679 1463 4719 1497
rect 4753 1463 4793 1497
rect 4827 1463 4941 1497
rect 4975 1463 5015 1497
rect 5049 1463 5089 1497
rect 5123 1463 5163 1497
rect 5197 1463 5237 1497
rect 5271 1463 5311 1497
rect 5345 1463 5385 1497
rect 5419 1463 5459 1497
rect 5493 1463 5607 1497
rect 5641 1463 5681 1497
rect 5715 1463 5755 1497
rect 5789 1463 5829 1497
rect 5863 1463 5903 1497
rect 5937 1463 5977 1497
rect 6011 1463 6051 1497
rect 6085 1463 6125 1497
rect 6159 1463 6199 1497
rect 6233 1463 6273 1497
rect 6307 1463 6347 1497
rect 6381 1463 6421 1497
rect 6455 1463 6569 1497
rect 6603 1463 6643 1497
rect 6677 1463 6717 1497
rect 6751 1463 6791 1497
rect 6825 1463 6865 1497
rect 6899 1463 6939 1497
rect 6973 1463 7013 1497
rect 7047 1463 7087 1497
rect 7121 1463 7161 1497
rect 7195 1463 7235 1497
rect 7269 1463 7309 1497
rect 7343 1463 7383 1497
rect 7417 1463 7531 1497
rect 7565 1463 7605 1497
rect 7639 1463 7679 1497
rect 7713 1463 7753 1497
rect 7787 1463 7827 1497
rect 7861 1463 7901 1497
rect 7935 1463 7975 1497
rect 8009 1463 8049 1497
rect 8083 1463 8197 1497
rect 8231 1463 8271 1497
rect 8305 1463 8345 1497
rect 8379 1463 8419 1497
rect 8453 1463 8493 1497
rect 8527 1463 8567 1497
rect 8601 1463 8641 1497
rect 8675 1463 8715 1497
rect 8749 1463 8863 1497
rect 8897 1463 8937 1497
rect 8971 1463 9011 1497
rect 9045 1463 9085 1497
rect 9119 1463 9159 1497
rect 9193 1463 9233 1497
rect 9267 1463 9307 1497
rect 9341 1463 9381 1497
rect 9415 1463 9455 1497
rect 9489 1463 9529 1497
rect 9563 1463 9603 1497
rect 9637 1463 9677 1497
rect 9711 1463 9825 1497
rect 9859 1463 9899 1497
rect 9933 1463 9973 1497
rect 10007 1463 10047 1497
rect 10081 1463 10121 1497
rect 10155 1463 10195 1497
rect 10229 1463 10269 1497
rect 10303 1463 10343 1497
rect 10377 1463 10491 1497
rect 10525 1463 10565 1497
rect 10599 1463 10639 1497
rect 10673 1463 10713 1497
rect 10747 1463 10787 1497
rect 10821 1463 10861 1497
rect 10895 1463 10935 1497
rect 10969 1463 11009 1497
rect 11043 1463 11083 1497
rect 11117 1463 11157 1497
rect 11191 1463 11231 1497
rect 11265 1463 11305 1497
rect 11339 1463 11453 1497
rect 11487 1463 11527 1497
rect 11561 1463 11601 1497
rect 11635 1463 11675 1497
rect 11709 1463 11749 1497
rect 11783 1463 11823 1497
rect 11857 1463 11897 1497
rect 11931 1463 11971 1497
rect 12005 1463 12045 1497
rect 12079 1463 12119 1497
rect 12153 1463 12193 1497
rect 12227 1463 12267 1497
rect 12301 1463 12415 1497
rect 12449 1463 12489 1497
rect 12523 1463 12563 1497
rect 12597 1463 12637 1497
rect 12671 1463 12711 1497
rect 12745 1463 12785 1497
rect 12819 1463 12859 1497
rect 12893 1463 12933 1497
rect 12967 1463 13081 1497
rect 13115 1463 13155 1497
rect 13189 1463 13229 1497
rect 13263 1463 13303 1497
rect 13337 1463 13377 1497
rect 13411 1463 13451 1497
rect 13485 1463 13525 1497
rect 13559 1463 13599 1497
rect 13633 1463 13747 1497
rect 13781 1463 13821 1497
rect 13855 1463 13895 1497
rect 13929 1463 13969 1497
rect 14003 1463 14043 1497
rect 14077 1463 14117 1497
rect 14151 1463 14191 1497
rect 14225 1463 14265 1497
rect 14299 1463 14339 1497
rect 14373 1463 14413 1497
rect 14447 1463 14487 1497
rect 14521 1463 14561 1497
rect 14595 1463 14709 1497
rect 14743 1463 14783 1497
rect 14817 1463 14857 1497
rect 14891 1463 14931 1497
rect 14965 1463 15005 1497
rect 15039 1463 15079 1497
rect 15113 1463 15153 1497
rect 15187 1463 15227 1497
rect 15261 1463 15375 1497
rect 15409 1463 15449 1497
rect 15483 1463 15523 1497
rect 15557 1463 15597 1497
rect 15631 1463 15671 1497
rect 15705 1463 15745 1497
rect 15779 1463 15819 1497
rect 15853 1463 15893 1497
rect 15927 1463 16041 1497
rect 16075 1463 16115 1497
rect 16149 1463 16189 1497
rect 16223 1463 16263 1497
rect 16297 1463 16337 1497
rect 16371 1463 16411 1497
rect 16445 1463 16485 1497
rect 16519 1463 16559 1497
rect 16593 1463 16707 1497
rect 16741 1463 16781 1497
rect 16815 1463 16855 1497
rect 16889 1463 16929 1497
rect 16963 1463 17003 1497
rect 17037 1463 17128 1497
rect -34 1446 17128 1463
rect 15051 1059 15097 1065
rect 15451 1059 15497 1065
rect 15715 1059 15761 1065
rect 16119 1059 16165 1065
rect 15045 1025 15057 1059
rect 15091 1025 15457 1059
rect 15491 1025 15503 1059
rect 15709 1025 15721 1059
rect 15755 1025 16125 1059
rect 16159 1025 16171 1059
rect 15051 1019 15097 1025
rect 15451 1019 15497 1025
rect 15715 1019 15761 1025
rect 16119 1019 16165 1025
rect 13519 979 13565 985
rect 13889 979 13935 985
rect 13513 945 13525 979
rect 13559 945 13895 979
rect 13929 945 13941 979
rect 13519 939 13565 945
rect 13889 939 13935 945
rect 1087 905 1133 911
rect 2937 905 2983 911
rect 5971 905 6017 911
rect 7821 905 7867 911
rect 10855 905 10901 911
rect 12705 905 12751 911
rect 13371 905 13417 911
rect 14481 905 14527 911
rect 14777 905 14823 911
rect 15517 905 15563 911
rect 1081 871 1093 905
rect 1127 871 2943 905
rect 2977 871 5977 905
rect 6011 871 7827 905
rect 7861 871 10861 905
rect 10895 871 12711 905
rect 12745 871 12757 905
rect 13365 871 13377 905
rect 13411 871 14487 905
rect 14521 871 14783 905
rect 14817 871 15523 905
rect 15557 871 15569 905
rect 1087 865 1133 871
rect 2937 865 2983 871
rect 5971 865 6017 871
rect 7821 865 7867 871
rect 10855 865 10901 871
rect 12705 865 12751 871
rect 13371 865 13417 871
rect 14481 865 14527 871
rect 14777 865 14823 871
rect 15517 865 15563 871
rect 347 831 393 837
rect 1456 831 1502 837
rect 3455 831 3501 837
rect 3751 831 3797 837
rect 4121 831 4167 837
rect 5231 831 5277 837
rect 6340 831 6386 837
rect 8339 831 8385 837
rect 8487 831 8533 837
rect 9597 831 9643 837
rect 10115 831 10161 837
rect 11224 831 11270 837
rect 13223 831 13269 837
rect 14999 831 15045 837
rect 16331 831 16377 837
rect 16479 831 16525 837
rect 16775 831 16821 837
rect 341 797 353 831
rect 387 797 1462 831
rect 1496 797 3461 831
rect 3495 797 3507 831
rect 3745 797 3757 831
rect 3791 797 4127 831
rect 4161 797 4173 831
rect 5225 797 5237 831
rect 5271 797 6346 831
rect 6380 797 8345 831
rect 8379 797 8391 831
rect 8481 797 8493 831
rect 8527 797 9603 831
rect 9637 797 9649 831
rect 10109 797 10121 831
rect 10155 797 11230 831
rect 11264 797 13229 831
rect 13263 797 13275 831
rect 14993 797 15005 831
rect 15039 797 16337 831
rect 16371 797 16383 831
rect 16473 797 16485 831
rect 16519 797 16781 831
rect 16815 797 16827 831
rect 347 791 393 797
rect 1456 791 1502 797
rect 3455 791 3501 797
rect 3751 791 3797 797
rect 4121 791 4167 797
rect 5231 791 5277 797
rect 6340 791 6386 797
rect 8339 791 8385 797
rect 8487 791 8533 797
rect 9597 791 9643 797
rect 10115 791 10161 797
rect 11224 791 11270 797
rect 13223 791 13269 797
rect 14999 791 15045 797
rect 16331 791 16377 797
rect 16479 791 16525 797
rect 16775 791 16821 797
rect 1309 757 1355 763
rect 2271 757 2317 763
rect 3085 757 3131 763
rect 4565 757 4611 763
rect 6193 757 6239 763
rect 7155 757 7201 763
rect 7969 757 8015 763
rect 9449 757 9495 763
rect 11077 757 11123 763
rect 12039 757 12085 763
rect 12853 757 12899 763
rect 14333 757 14379 763
rect 1303 723 1315 757
rect 1349 723 2277 757
rect 2311 723 3091 757
rect 3125 723 4571 757
rect 4605 723 4617 757
rect 6187 723 6199 757
rect 6233 723 7161 757
rect 7195 723 7975 757
rect 8009 723 9455 757
rect 9489 723 9501 757
rect 11071 723 11083 757
rect 11117 723 12045 757
rect 12079 723 12859 757
rect 12893 723 14339 757
rect 14373 723 14385 757
rect 1309 717 1355 723
rect 2271 717 2317 723
rect 3085 717 3131 723
rect 4565 717 4611 723
rect 6193 717 6239 723
rect 7155 717 7201 723
rect 7969 717 8015 723
rect 9449 717 9495 723
rect 11077 717 11123 723
rect 12039 717 12085 723
rect 12853 717 12899 723
rect 14333 717 14379 723
rect 3603 683 3649 689
rect 4713 683 4759 689
rect 15813 683 15859 689
rect 3597 649 3609 683
rect 3643 649 4719 683
rect 4753 649 15819 683
rect 15853 649 15865 683
rect 3603 643 3649 649
rect 4713 643 4759 649
rect 15813 643 15859 649
rect 199 609 245 615
rect 5083 609 5129 615
rect 9967 609 10013 615
rect 14999 609 15045 615
rect 193 575 205 609
rect 239 575 5089 609
rect 5123 575 9973 609
rect 10007 575 10019 609
rect 10121 575 15005 609
rect 15039 575 15051 609
rect 199 569 245 575
rect 5083 569 5129 575
rect 9967 569 10013 575
rect 495 535 541 541
rect 865 535 911 540
rect 1827 535 1873 541
rect 2419 535 2465 541
rect 2789 535 2835 541
rect 5379 535 5425 541
rect 5749 535 5795 540
rect 6711 535 6757 541
rect 7303 535 7349 541
rect 7673 535 7719 541
rect 8635 535 8681 541
rect 9005 535 9051 541
rect 9597 535 9643 541
rect 10121 535 10155 575
rect 14999 569 15045 575
rect 10263 535 10309 541
rect 10633 535 10679 540
rect 11595 535 11641 541
rect 12187 535 12233 541
rect 12557 535 12603 541
rect 489 501 501 535
rect 535 534 1833 535
rect 535 501 871 534
rect 495 495 541 501
rect 859 500 871 501
rect 905 501 1833 534
rect 1867 501 1879 535
rect 2413 501 2425 535
rect 2459 501 2795 535
rect 2829 501 2841 535
rect 5373 501 5385 535
rect 5419 534 6717 535
rect 5419 501 5755 534
rect 905 500 941 501
rect 865 494 911 500
rect 1827 495 1873 501
rect 2419 495 2465 501
rect 2789 495 2835 501
rect 5379 495 5425 501
rect 5743 500 5755 501
rect 5789 501 6717 534
rect 6751 501 6763 535
rect 7297 501 7309 535
rect 7343 501 7679 535
rect 7713 501 7725 535
rect 8629 501 8641 535
rect 8675 501 9011 535
rect 9045 501 9057 535
rect 9591 501 9603 535
rect 9637 501 10155 535
rect 10257 501 10269 535
rect 10303 534 11601 535
rect 10303 501 10639 534
rect 5789 500 5825 501
rect 5749 494 5795 500
rect 6711 495 6757 501
rect 7303 495 7349 501
rect 7673 495 7719 501
rect 8635 495 8681 501
rect 9005 495 9051 501
rect 9597 495 9643 501
rect 10263 495 10309 501
rect 10627 500 10639 501
rect 10673 501 11601 534
rect 11635 501 11647 535
rect 12181 501 12193 535
rect 12227 501 12563 535
rect 12597 501 12609 535
rect 10673 500 10709 501
rect 10633 494 10679 500
rect 11595 495 11641 501
rect 12187 495 12233 501
rect 12557 495 12603 501
rect 2049 461 2095 467
rect 4343 461 4389 467
rect 6933 461 6979 467
rect 9227 461 9273 467
rect 11817 461 11863 467
rect 14111 461 14157 467
rect 2043 427 2055 461
rect 2089 427 4349 461
rect 4383 427 6939 461
rect 6973 427 9233 461
rect 9267 427 11823 461
rect 11857 427 14117 461
rect 14151 427 14163 461
rect 15813 433 15859 439
rect 16109 433 16155 439
rect 2049 421 2095 427
rect 4343 421 4389 427
rect 6933 421 6979 427
rect 9227 421 9273 427
rect 11817 421 11863 427
rect 14111 421 14157 427
rect 15807 399 15819 433
rect 15853 399 16115 433
rect 16149 399 16161 433
rect 15813 393 15859 399
rect 16109 393 16155 399
rect 15059 253 15105 259
rect 15725 253 15771 259
rect 16391 253 16437 259
rect 15053 219 15065 253
rect 15099 219 15731 253
rect 15765 219 16397 253
rect 16431 219 16443 253
rect 15059 213 15105 219
rect 15725 213 15771 219
rect 16391 213 16437 219
rect -34 17 17128 34
rect -34 -17 57 17
rect 91 -17 131 17
rect 165 -17 205 17
rect 239 -17 279 17
rect 313 -17 353 17
rect 387 -17 427 17
rect 461 -17 501 17
rect 535 -17 575 17
rect 609 -17 723 17
rect 757 -17 797 17
rect 831 -17 871 17
rect 905 -17 945 17
rect 979 -17 1019 17
rect 1053 -17 1093 17
rect 1127 -17 1167 17
rect 1201 -17 1241 17
rect 1275 -17 1315 17
rect 1349 -17 1389 17
rect 1423 -17 1463 17
rect 1497 -17 1537 17
rect 1571 -17 1685 17
rect 1719 -17 1759 17
rect 1793 -17 1833 17
rect 1867 -17 1907 17
rect 1941 -17 1981 17
rect 2015 -17 2055 17
rect 2089 -17 2129 17
rect 2163 -17 2203 17
rect 2237 -17 2277 17
rect 2311 -17 2351 17
rect 2385 -17 2425 17
rect 2459 -17 2499 17
rect 2533 -17 2647 17
rect 2681 -17 2721 17
rect 2755 -17 2795 17
rect 2829 -17 2869 17
rect 2903 -17 2943 17
rect 2977 -17 3017 17
rect 3051 -17 3091 17
rect 3125 -17 3165 17
rect 3199 -17 3313 17
rect 3347 -17 3387 17
rect 3421 -17 3461 17
rect 3495 -17 3535 17
rect 3569 -17 3609 17
rect 3643 -17 3683 17
rect 3717 -17 3757 17
rect 3791 -17 3831 17
rect 3865 -17 3979 17
rect 4013 -17 4053 17
rect 4087 -17 4127 17
rect 4161 -17 4201 17
rect 4235 -17 4275 17
rect 4309 -17 4349 17
rect 4383 -17 4423 17
rect 4457 -17 4497 17
rect 4531 -17 4571 17
rect 4605 -17 4645 17
rect 4679 -17 4719 17
rect 4753 -17 4793 17
rect 4827 -17 4941 17
rect 4975 -17 5015 17
rect 5049 -17 5089 17
rect 5123 -17 5163 17
rect 5197 -17 5237 17
rect 5271 -17 5311 17
rect 5345 -17 5385 17
rect 5419 -17 5459 17
rect 5493 -17 5607 17
rect 5641 -17 5681 17
rect 5715 -17 5755 17
rect 5789 -17 5829 17
rect 5863 -17 5903 17
rect 5937 -17 5977 17
rect 6011 -17 6051 17
rect 6085 -17 6125 17
rect 6159 -17 6199 17
rect 6233 -17 6273 17
rect 6307 -17 6347 17
rect 6381 -17 6421 17
rect 6455 -17 6569 17
rect 6603 -17 6643 17
rect 6677 -17 6717 17
rect 6751 -17 6791 17
rect 6825 -17 6865 17
rect 6899 -17 6939 17
rect 6973 -17 7013 17
rect 7047 -17 7087 17
rect 7121 -17 7161 17
rect 7195 -17 7235 17
rect 7269 -17 7309 17
rect 7343 -17 7383 17
rect 7417 -17 7531 17
rect 7565 -17 7605 17
rect 7639 -17 7679 17
rect 7713 -17 7753 17
rect 7787 -17 7827 17
rect 7861 -17 7901 17
rect 7935 -17 7975 17
rect 8009 -17 8049 17
rect 8083 -17 8197 17
rect 8231 -17 8271 17
rect 8305 -17 8345 17
rect 8379 -17 8419 17
rect 8453 -17 8493 17
rect 8527 -17 8567 17
rect 8601 -17 8641 17
rect 8675 -17 8715 17
rect 8749 -17 8863 17
rect 8897 -17 8937 17
rect 8971 -17 9011 17
rect 9045 -17 9085 17
rect 9119 -17 9159 17
rect 9193 -17 9233 17
rect 9267 -17 9307 17
rect 9341 -17 9381 17
rect 9415 -17 9455 17
rect 9489 -17 9529 17
rect 9563 -17 9603 17
rect 9637 -17 9677 17
rect 9711 -17 9825 17
rect 9859 -17 9899 17
rect 9933 -17 9973 17
rect 10007 -17 10047 17
rect 10081 -17 10121 17
rect 10155 -17 10195 17
rect 10229 -17 10269 17
rect 10303 -17 10343 17
rect 10377 -17 10491 17
rect 10525 -17 10565 17
rect 10599 -17 10639 17
rect 10673 -17 10713 17
rect 10747 -17 10787 17
rect 10821 -17 10861 17
rect 10895 -17 10935 17
rect 10969 -17 11009 17
rect 11043 -17 11083 17
rect 11117 -17 11157 17
rect 11191 -17 11231 17
rect 11265 -17 11305 17
rect 11339 -17 11453 17
rect 11487 -17 11527 17
rect 11561 -17 11601 17
rect 11635 -17 11675 17
rect 11709 -17 11749 17
rect 11783 -17 11823 17
rect 11857 -17 11897 17
rect 11931 -17 11971 17
rect 12005 -17 12045 17
rect 12079 -17 12119 17
rect 12153 -17 12193 17
rect 12227 -17 12267 17
rect 12301 -17 12415 17
rect 12449 -17 12489 17
rect 12523 -17 12563 17
rect 12597 -17 12637 17
rect 12671 -17 12711 17
rect 12745 -17 12785 17
rect 12819 -17 12859 17
rect 12893 -17 12933 17
rect 12967 -17 13081 17
rect 13115 -17 13155 17
rect 13189 -17 13229 17
rect 13263 -17 13303 17
rect 13337 -17 13377 17
rect 13411 -17 13451 17
rect 13485 -17 13525 17
rect 13559 -17 13599 17
rect 13633 -17 13747 17
rect 13781 -17 13821 17
rect 13855 -17 13895 17
rect 13929 -17 13969 17
rect 14003 -17 14043 17
rect 14077 -17 14117 17
rect 14151 -17 14191 17
rect 14225 -17 14265 17
rect 14299 -17 14339 17
rect 14373 -17 14413 17
rect 14447 -17 14487 17
rect 14521 -17 14561 17
rect 14595 -17 14709 17
rect 14743 -17 14783 17
rect 14817 -17 14857 17
rect 14891 -17 14931 17
rect 14965 -17 15005 17
rect 15039 -17 15079 17
rect 15113 -17 15153 17
rect 15187 -17 15227 17
rect 15261 -17 15375 17
rect 15409 -17 15449 17
rect 15483 -17 15523 17
rect 15557 -17 15597 17
rect 15631 -17 15671 17
rect 15705 -17 15745 17
rect 15779 -17 15819 17
rect 15853 -17 15893 17
rect 15927 -17 16041 17
rect 16075 -17 16115 17
rect 16149 -17 16189 17
rect 16223 -17 16263 17
rect 16297 -17 16337 17
rect 16371 -17 16411 17
rect 16445 -17 16485 17
rect 16519 -17 16559 17
rect 16593 -17 16707 17
rect 16741 -17 16781 17
rect 16815 -17 16855 17
rect 16889 -17 16929 17
rect 16963 -17 17003 17
rect 17037 -17 17128 17
rect -34 -34 17128 -17
<< labels >>
rlabel metal1 16929 797 16963 831 1 Q
port 1 n
rlabel metal1 16929 723 16963 757 1 Q
port 2 n
rlabel metal1 16929 649 16963 683 1 Q
port 3 n
rlabel metal1 16929 575 16963 609 1 Q
port 4 n
rlabel metal1 16929 501 16963 535 1 Q
port 5 n
rlabel metal1 16929 427 16963 461 1 Q
port 6 n
rlabel metal1 16929 871 16963 905 1 Q
port 7 n
rlabel metal1 5089 575 5123 609 1 D
port 8 n
rlabel metal1 5089 501 5123 535 1 D
port 9 n
rlabel metal1 5089 723 5123 757 1 D
port 10 n
rlabel metal1 5089 797 5123 831 1 D
port 11 n
rlabel metal1 9973 575 10007 609 1 D
port 12 n
rlabel metal1 9973 723 10007 757 1 D
port 13 n
rlabel metal1 9973 797 10007 831 1 D
port 14 n
rlabel metal1 205 575 239 609 1 D
port 15 n
rlabel metal1 205 649 239 683 1 D
port 16 n
rlabel metal1 205 723 239 757 1 D
port 17 n
rlabel metal1 205 797 239 831 1 D
port 18 n
rlabel metal1 205 871 239 905 1 D
port 19 n
rlabel metal1 205 501 239 535 1 D
port 20 n
rlabel metal1 1093 871 1127 905 1 CLK
port 21 n
rlabel metal1 1093 723 1127 757 1 CLK
port 22 n
rlabel metal1 1093 649 1127 683 1 CLK
port 23 n
rlabel metal1 1093 427 1127 461 1 CLK
port 24 n
rlabel metal1 2943 649 2977 683 1 CLK
port 25 n
rlabel metal1 2943 871 2977 905 1 CLK
port 26 n
rlabel metal1 2943 501 2977 535 1 CLK
port 27 n
rlabel metal1 5977 871 6011 905 1 CLK
port 28 n
rlabel metal1 7827 871 7861 905 1 CLK
port 29 n
rlabel metal1 7827 501 7861 535 1 CLK
port 30 n
rlabel metal1 5977 723 6011 757 1 CLK
port 31 n
rlabel metal1 10861 871 10895 905 1 CLK
port 32 n
rlabel metal1 12711 871 12745 905 1 CLK
port 33 n
rlabel metal1 12711 501 12745 535 1 CLK
port 34 n
rlabel metal1 10861 723 10895 757 1 CLK
port 35 n
rlabel metal1 2055 427 2089 461 1 SN
port 36 n
rlabel metal1 2055 501 2089 535 1 SN
port 37 n
rlabel metal1 2055 649 2089 683 1 SN
port 38 n
rlabel metal1 4349 427 4383 461 1 SN
port 39 n
rlabel metal1 4349 501 4383 535 1 SN
port 40 n
rlabel metal1 4349 797 4383 831 1 SN
port 41 n
rlabel metal1 6939 427 6973 461 1 SN
port 42 n
rlabel metal1 11823 427 11857 461 1 SN
port 43 n
rlabel metal1 11823 501 11857 535 1 SN
port 44 n
rlabel metal1 14117 427 14151 461 1 SN
port 45 n
rlabel metal1 -34 1446 17128 1514 1 VPWR
port 46 n
rlabel metal1 -34 -34 17128 34 1 VGND
port 47 n
rlabel nwell 57 1463 91 1497 1 VPB
port 48 n
rlabel pwell 57 -17 91 17 1 VNB
port 49 n
<< end >>
